--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
LB3aUEj4hslbvCNFLuQqf4SdjU7urfbDcNq7i3j20nbC9SwBP24kdZi0AaoYzWWLh4WSEb3du7p9
LSd6OOnS3u8OGqCLGvXMnBxdixLMGd1XCS0KLIDA3B2t0CS84gWjwfEmJL/1uZIuBdUsTXzcKgUg
6ONcratiFmyp2hjxiMpuFrCDRrpGwTzWD0nvTwejh/q2WBnlTRWSHPANq/JoVjz3rW9mTCt1Rdy2
ONugjHssZmlps0iaTK3lOiSkdcy6Joj7OHbs2lJ8ecP3rg7gbK+iGE+Pd9yHVAxg6+VT4qLxY3iK
oNIGlIMMuHts+SCbgPyq/mYUG3iTejZbU7rcVw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="u6TC6SXH/xqgAw0HCBPIDUhK6hHALVlVZxPIgOmCaMA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
KORIwUlhacjYv7xF+kOkqMs4NGX+Do/I2Ffe+GUldW8z/p6Er/qn+iF2GobUhqNWISHZhaWm4DzJ
tvNE25QlZnzdIrhB75A9XTPaqAmsCzhnhqiuAPtWKFct9zkibgzyx5P93wvMWlfaW6OQJATEEY/g
e2qSZN6ExyUu/VFSKXFMneGMaIiF6t6X1peSubQKzBDNycA81FYTWMnXbRMqbl2/sPcva/7EopHW
T73l7iqu3CSYEzDqbDzWkdd/WQVYKytijPvlR3POiPkg3X29J1bD3Rd+ud0iDei6d8rj5ibACIRV
FcIa4N7WbrtqW6G4qpqotblVGbXbvYe3W9S9tw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="kFgjKRpsaovazxj+7ai6yH3o9+TUfwCJ23gfJXWcPPo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2208)
`protect data_block
5Dt8iIoW9E7INp1MKfoEIo13Qn8KDYhCB1QGD9SGSjwbrcM27v8T3JbY7mqUyHkJoEgC973Oeq7+
tGBJlyUvGJUL7ggAGGMyfH4DwbzU9xcKes71gan5nwp9ry91GzNeC76fR6WfMPyAWHi49AnPR9Y5
MnuHfQ1bm5rbztIutx7AMZqCfpZGmDBjD/fPz63dF2jGmZbLFOdMLd348dM2ytk0s6qpXf1mBvul
4gEh5ivC6nDYmEa9vNXbsG3HA0dJ6z8u1AxrRJOG3T18SrYBP+njfLQIDB/f61galO9cHxyEfWKX
nCbs7lCptjxoq0cHC02zaVA3smEESnRibt4sMzrkRupO7ce5a3tKR6/xAyG39ZGgE49HrSCnwCmZ
ehdlYM2v2B8y+sq3rOSgUtVMSprM2YCQQBc5Xz1yUU8MEex40upnv7nY1LWm0gXuixxiU/sd/BNF
BvnKgbkqPRuKb+2ZeIsgaWYfyRHAGdPWJq6OVHGhXBhzMC3Eg0nrE+YaMvM+LyQK2T21UAZfgzBh
LgimDzfni2a/wNDNupmHrFsjjXCS+Z5cDgLXazlODjzDAVyBNfFiGasPXV3TBhewfRcnr1mazyry
WYkumU+/wKDm86TfyVyoUGwKWdmanvHEFADJEx+Q8Ko3O+/61B3KkvCihtTjjT5NlTJH08GDLUFO
SZJcS8beSvITPt2yO8HohuLa/FDZgYk8IT7CDJScb1YOwFt1eQOaiY5PkwOBUUiTjZ94hLiyivio
FW7XN75mRPexwajXDjRiuzTfh9PgvOxc5KWSYmCprl9ICDXuSd29x9jlNmcCWpO8MnWH02Dhqayv
tg1uaz4byxx80TKtVg1K+0FoyD563e14Lbqb1CIpSq/Zghut96gcrrugxxKIw3H00UOGqNEFqND/
oV3rjdXNK9bVayQXm7BU0gMQiBHz0jbKnlwXqUN5mNt6JDJCBHLWmey123Z8M404+4jhzIW8pClK
gyJGJAxtJHhtmTqvGPUxJXt8r/xhGP93r4GLXvk/x/PBoQT2ez32Yd55tWePrxcJrvjWKye94Ft8
7VuIdqQKp9xIgwMv30BgjGhUuWG++JAAK5IUdDWhrNsnUmnErn3n+85G2tDjbOOBHQdpJlXRlWyu
XGdLZsz/dP1PhgogEjTqVKkf4c2DPIc41Q5Df8+IkR/yXVww4Q9olSRTW0YkK2/MOdmt0PgF5RUF
jzoK+JZYWeKvIXsqjrPhXije43+Gx2iK8RIqLKsb1ddxvKzqGhyezGHb8ikAzS68ntDZeyy8auE1
0r4u3pgcdf6dmFsBuQ/VH1snQn2Xev3mnVrNozwvrA+L9T0znpcjf9S0aSLdwAhGhtUrfEwM+9cw
bwUAC6Slvw0IQaNfWPTfxvBmzXjr4MIyEjI6dSZZe9Vu2ScP0WnxwkerRff3rgGODOq4RjZDkYdD
cbwF8Jl6SDz2FoQYOzWv4bCEoOmUyiC81WL3qzvVgpIGo8KJkt4b6EQKYvzaBvKuGbLKz2ZRyN4I
Feof4FMZb5n9G2ZGeHi6/7aay6wVqT41CymDfEBapyxTgP+mEctYICn9mdqszvIheGxijB+4Sj4w
pOwaCTgA7UxkjO8NW/VvMS5oMrg26j2U2yxD6ZNCKx6s2/Unekkn3j/i1ifzTtlQxXw7ztXCG8PO
8kvxHJTrBSr0O+EBzr2Haa1v60EG4z0YbdhCRX/aYo6K5XLfHYhUDzISf+rI610m+D+jgj8na5c1
jOc53mcc8bDM8VzvcWnWTjGGpWqcqT7N8PaMIMkAh9opagaJn5BhVbOvb72wkOjEstluzRyvgB8r
b6tal8TmcDRs5kYLBEUCV5zWaVMc1jiqe9DXr5VtdRhWWGWuCVbmCkGibLhwT2L202hzfxU9fcwN
IJs9WgWUAzi6sxOunnencmPgIJw6c0aaih/thBWFryDstRZ8DmnZ7jwvcjX+260CEvrWuTYIDWSM
mHRGz+UbQDZAiMboo4NWKgWPXrGbgt434z1toSa3ToH1acjdLJfSBjW3e/m7zL9n4IyU3XLlq9ow
vipXJ/tkynYojYdfFR9ua3CXpf2I/g+HCqO4MULpIQuOfJxoQCatoH9r8sw587CC0YSp4ZSmpiU6
edEUETUJVJCvego7wtdJJgtKORrDY1ebUgcp0zc8/uQV4JV4SCdefqvpnEaOgam6Zv90kkwzHoNi
fvgv+LmQVVse8fIJIZZshLwyIZjCFIlsSJPLbpv9FpW+uqlnS9dZDzOqLrFcOWNYSt39t82jrCqH
08GF+0bwvKD/RYCmRIvR5j9VMXZ3o9RzQnaKU+kAYFsgelWGvdsSnigXUDzhxcXhZxhzjR0Oz8iT
w2e9iJm1l3NqlaM9wBgJKBUlX/GwUC0ko6rwNNZ0FPrdfGokrjnZkNuU+yIl8EtH2lr+Bq3DInVU
AGXSrp9PG5leaRamTzauGRYnQ2eWDoiBapEEHFipw0NuiJaK0ElGjGBWH7x/I09yvP+IoZJxM3RV
uEwNuqY6CQ0w9xoLmrMkaVX37IY53PIg04yVwWii68bUKR4F5f5QnKA/cM3RlzltmZRmQxmsYgfN
r4q1ydwDcHfk6mPGPh9G2f73/J2hiiBlEAqVbl74KcemDKXEZKKMlQQdsk5A60uxv6TZpfyyUUUk
Q7aSzNTRBhZ7oH22xFKjy7dbKbddEtAc6O5tPlYKg3Jh3lCMIviHSRmCseHzlYE4ODpkCwRU48YQ
naYuY7QT3GAXdde23zmcwsyQqP/cKCUcsvXz3C0w64cvI7ecPIMnL7933vyby8hlPb+saZwsYYpD
MCkBkH/UbBDuJhJnnSI9FaU5b5xLstYOVFtb5gFMsWnizTGrYHYI8v4YcN1YxGdpMifq9KeREgHh
qamZg2T596GnsJc7hnRwkVylICe/TOCM8Y5S+BJ8C7DAy91Et14jVivV
`protect end_protected
