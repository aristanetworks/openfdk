--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Qbdj3ef+CFqEuSJrcwe6tO9ZHXNCDh5iNNaevZw7189S74xs0Od5MXu7mnZbR+ze8kH80rwADwlN
2omvHg/5QX/a0XDZq86YFo1XCGb+1nsk7FTiXBGN/S/cJLhSSdBqG353x/+6CRt26SLI1mHZdMtX
BYgW0UOtOJF1IHc2hZAkmR42JxOzElgnl9ZNdyZTPOWUoPV4pHhE3GDty/RP41Rf1QnDLhn+rSzZ
36OyCly6gSs9yD/p2Fqvkof2l1KGSd1Xy1JG5Dhp81BLvm4uD7NcTDUKQyQ+A9+dDmZlo+6FbCN4
Whk08iroN3NXdQwOaliLfLGeR4DJGa/b+mfLeQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="TtRpgfhpL2z56iGChUbcBM7Jrtb6DewKHFQanBsguuI="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
YuVd4BkgE812YXj9sQGiiiVgsY4w9SOgec/2iRtaxR/Tyc16lXcMHWCfSGnZVcdlWOwiXefFzKd6
tsdF7P4u7zOzKBK6svdUZqamnj/9WL23GebWR0InD5NYiLZ4jopq3ZRN0sAhMzO5bt5FWndCu2Ko
Sr0iS/7Nc89aVvXt5zpPTDeeSMVX9hCaDTSrrNn3xeYyfbOB0V5bAbKD7iRsIgWfILe3X8nsQJkP
t7IQ0Xm9tIpQHTRRejX1hcwgonTjx5JXvOClM49i5cqScYETAujzwPCX0CjtsZYGVX4gT0pHWHqC
VDED6pFNi90s7/npNk1MfnlVcWOUd6zhNq4a8g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="BhtPco56LtTKJ79VwR3n+TK3+Q/D1g9QqnwqMHH314E="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6608)
`protect data_block
H5iqpT/aHbBRL+BDAO9U9OLOLtPMrT0JO0JrWB+QzTWnOdSWa4nqh+2gHiwIIlhxzYaNhntRTdZP
xQveEgB5Nl+19L4PyECfha8+FQLBD/SR9vtKJ5obfzrd171H8PJukMsV7Cia6+0xhHUOwxy6Qd/V
A/DobBddre/moBNHMBp0yf0eMRSVxXztNtbmTBLmPXGq3YUBSF2FWrLFhwC6pa2dEz+SpUwJLOCZ
ELLN+KHD6jbgXPyJI41zmu7+0QxUHw+psHH/W09epf3a57L08uKg9vh06DuJ5t1p0n/5TJEFswTk
oDEdS1T07xDMzckRz7OVyx/ePwAZ7rp1BCPELCeF6EuH9cJshawf6aGcVl6A8pX7QGzAEWQgeASq
lcTRBjQqQAl4Sf0zVQ36zbH3hDaofxLcLWyAdZit724gfhQ3NGOsLRRZIhnyhvWNHwht+88o9oTS
3Eqy5uL43/R3xy8u7Evy+0y7F8Ykonh/k3zovSxwAS+ZAEoD/HIF+u1K0LpES2PFL7Kk7oj9hjNd
9xmChKgymsCv3xeXQb1UOpTYGAJMCaKe8NT9SeBtSUDjESt9dvaKqZI59A1lL2BI3kIfV7E7nqOH
vGEVWlK2j+Ifand9VyaU3FXV6PylWv9nhX01p+Kah9XZQd2LqXuh8+7V7L78Ct7ConkQDn5Dtxsm
NpHPETgsZN3HOiMPDvjrwBjGcWSniBQvz2fDlHXKlHTPgVs3N2pTvzCLxThLTZxq1plh728hVtKN
pWZFAp9ks4VX9U0iqyj7O/9V1Lu21kRuUX8OmadfUee91iqJJZ35E0v49FbcL3wXg6u+SHv8f0BM
XDLutBqs+qB6LfjV1HLdjvvxdJErePIgxt5FxMFSRvRI/EP3X5tVaYx6XlrBXQG8gJRkH9kw8FZB
GKrCNSBSkWOzgBSKXtOty+RdL/DnzkuZkxE0/qzWEF94XSUTwP82YZsrmG4fpeqhWdhWZ0+tYNOr
OpACpMM2sI2WuVeVEhVa3Mq/b4oXBXXxEpdiidM65gYzQ4/RwrmtzeFqOP8p1rDxiNc1w6/EURWR
2JHif+NhXzbxmWcVT2G3mgAQOhsNtvoFYntz4bVByRkRb8GKv5a8MvJ1hmv5A7BHV6VWcstuuiGq
Q10wT5vFTeGGGMRRR7z03gCm8HDkTDforurX+rbsjuqcDvpN7zAHRDRiVQ+DWbYJJnXy/ENwANHz
/+9ahO+1AMU0Zx+J9id8Y3yWimv5r9VNzlvvpARi4M4iwGDBn69HtZ5t2Dee7jKTc6i88y3gIkcw
vLD7o2NL6UVBbOujxzmry6Vj990z0KbNjOzersO9yWMNQPxkRk+0q9GMxO4EMMYXB/KDMcoBs8Ds
EBvzjUM5fzpUJK4e3qbQd1PAcoGYPWKoccjpG2QYI+KmfrbHzFN1mnlbKX89eN0rRFnX6dVqpQTi
qTZUwCP98QaroOkZzJo2SY0N7ZLEoW2T1ZN1/h0xDP1HFFA4P9CaVLcqVVdrPpT+phwYX09EZVx2
fhXgvArl2L8EsbaLu0vy0ppHAt9lSUTwXb5x49+tho9TCDF/rA8MYu449TH1AJiqbZDEuW8SjXzn
xLuPgifGMuOFtvzgpT57/x/UtABJBvpRnrcwcYZNhoxcE8YS+gQmUFoQvDs7pdRFw8bIx6AI6xuL
kHZmf8mYWuHK7CjNuMysB/V1RlRN9rpFnwPZaTP70kFUidBVeoL0rO0xELZSJ3uhRaKenOZmQVeX
OItjbQ4vBizo+4v3uYW9UozkcsOQvc1Wv5eg8wxCNIAOdAVkzRHwtSmndCHJzPYFcJRTn569KELM
ndVeVm/eIyIEdblUjMzSGEuyWmKZlLmoXfS+fvrgDvs603euYY2GiADLFomBJxGVbTzaq4pcbx7m
j4kJGv7xKO2rX7AtllRb0Wpq0Ujbep8SkFUVLUaXAVCjZbqwFtCvWQvQl97eNzrrUnd2lBQahJuK
TEnBXYV3mycWDS9bvhM1LjLFzxYZM7vizL8T90e5I+2MkP3GMScRL6ffDlprwAdawo9tS6Wg8LUk
QTzbz+qcQUclmEuGqfla0B3hphBztTorlpxm4SVBQz14EDei6eFcq6uRkAQp6obtXigDik5tYo+e
jdkO/6iS+MBVZ5gyZI1x2fHJpJyq2F3jeAmCkes9KTZ9giA332AYXp5bCHMELE8Q2Sf4pKUo0rwv
TVAUv8DDnHEyh/QFCFjXvB3meBLxlg4DjHgXmgJqjs75DGp/hDqvYs/2IJ5Lp/cjF3mLmPmjEBEm
bPa+glsAcJ29xqAMCZw5YMoreUGwuQ5jE7KZ26pcDRrHkcYtVgIyJETCVAmYGdVajLluUe6dpfUg
/91X8qxuddYjWu+BGiow5hG0tNvCPnR7fc3qsCdQDSKpk7mMCSX+GwQNx/Zy7IU8C5szDu3x4uU3
KQ4n8rIUYAp6AOWqLwq8lQutgfTPKeksYCzTakvfa5rkYAC6Xxss/IEZL/ALEAjLE4tqu6dXMDij
FWp5wlFggBwNeXHJlM0TSztot2Sum+4fsGmn4Rg7H6kkK1JL0cag2DCtxyR08jNILf/YPT9IWTty
kmTjCrGIR9t3tcpYD3qMKG1nEEM9BdpSmoaFqsAxsfD5DYw7CvXmkUtbJYatTaB8vo3LjqcUhp9V
/dms7lguuexDZSwHl5dPEtQirRiPFGXPQlAhTPmsQ/xzRsjYj8je65k9LbKDtm7a7JA/JBa05ced
EPU+J3vqTwWf3GzaLVGEQY+j29d1tbgVhjW+toVah7tokiD1wG0mq71kl0Wk+0/B1DR3JvxF7afV
rZhTxWXSEXvEYeR6Ju8Hg4b4Q3ZCnBWi8j71uzzoxtYCdmUn3PCJxNrmxed8ncvpDYXFX2P2oBey
SetgAL1QpDPcc9NWI5NXzfOXfs7gf8QPR/ZrmZBj94kjiYzhHqYDMGnr4lZ2NiZGiJ+DcZz5cAbt
nPmNCFzMXzQVxaTupDdujIvlhRL6IlFZ/qchCYTz/OdbCKLWCv9OSLei/lrO/3OUtuyIdfqJU4eC
2x3VoRN4wRvJu6xam4dQD+RkQRkgVW7nh1AFH+lxJFGzDUEZgg1BCPBuOuwwn4J3KW9iFiqbxuj8
tqv71VQD2r8lSppIzSNvnwnRRJVOM5J0Hj3TckvKD8+lr8bOudR5XzOx66hg46azm26FajzyubIt
LsVU52kKIcOeVmgHxvb4eaU2DTgfEXJI/cKXTlTdi5+daaMk1vOnYTbIxOyAF8sbKvg30/CpekUh
AnGMtD6Os4MrjI+za6thYfo0GRwvcJOa7wL877MFKf5QbCRKGMNJ5081oBoDkm0+INyTIA+QcA/O
gdN57xjXC11kI8OGRHKYeNVNeIjggBEpmxlffkYmo5PjY41rNPkHoSOm8GuyFk56BCEAE5UeHEb1
T7HgtLkwn+VAeXd2v3tgypB6tcQgWp/ukI3jMIkOHVsLXADsOPNmCX8PBSGYEgrnofxGY7PyjumW
9GBVM8HPkuRPEWHxQK3pp/DyOV+jMJf9xNhN4G4kDJXWF2+6OGNDiv0WeHokIS6YsP6F7+q1lg+1
SzKg8mcPDXKHwZ6ePxDk1NmA2CtEBOHVQZ0CpNmeqnc53t1/UzP3HHF6DhRbEwEt+YCnoifs0U9s
0FDARQX1rW2V7EVQY3shsP0A+P1pqdyUN5us0EkkdQOqcL4EcMBGF9W76gb8X0gWegOanCG67QXe
GtUFEw8DmMl9FuqBNb/EcMiJF0GJYObA8wTMrkIrdaXzarHFpMG6Trok9tYedQxWxyR9nqhdiSDE
U6vclBZkP5l6dTB81Exro4SvMyiTyhNFWWvunNPVK06XmNRvA6FdrmzFmsBzlLvt41BiR0Oj6bYZ
bJfDBFitQgwGyGR45SXJROZKzUe0BlzDOJuxhK3SQ/41iCQeuiZTLeGMlXyyt/MIRQ9pjneMEch2
j2V3cFCi4KfcykmY5RF/k5NMVa4q2P7OPyfksv5wDvhTIXNbzoLgo7I/9CbwFcVKMkA4V5NaInvi
uaFRVbYi2WzMYMs6Hw9+3bTx2KzM257m/TdPsaA2HTSaZGEWjjXAf/nqFVwA1k+jd3t7wIonZzPa
iDnkvyvsjUDh4Yq4p5GsGnNWMS4cxU3C78F9qFuK9/TJQH8LRf9OMFXsmJ6iyHeKuEnDar0Nq8V9
fPC4FrwST+oMSduk4GuuVf0Hh2vNDBLZSDuGDWLrT5g/xbQn6tCNE/KXKbmRPEH1TD0a3G8pZd+T
mh/uRx6Ud93HP8Dju2DLYrjiS8zq6C/BIhvvOQoiptbajxqoVb+zFgWWjDzxGQOA7H68n9JfPN8M
XOwKt1okNHy6BysmKF7WYq0urH508FdRfkiXC3HQafFQyZnopJPUIP3s87eQgOhAuJAceo8740ik
BACa8aVx99ZcC4LYjt1SZC4dHvRv6wbxTweDuweDH5P61ys7CqLtOUYsX7gwHWdG7HLtbUBrIlQs
zsiUYqWRjoZvKVhTRMzU0zUV34upfo4A26YF8ddSs/t2RzqIiOCiFxQneJ2ucXSElLCup75wSABI
xInegbc/+4U93LDQvGr2hFFFhKs3s1H074EUEd+oZ9Q5XdsDT+XJBdCLq1FocjLbX7FsxN81NYWy
RQZGhtPyiUZs0tMfFD/Qje2/3a6IB6GcA/JOlefJQ7sDe9jneu7TiYsPtUp1l3UiHLuS8CTd/j+M
8ECMKJeLJU+BHPduHqlOcFow5mpsEoAquBfMWn6DdbjvC0vtxXMdr5h7/wfgHqOZSBN58f2T+5L3
/BcN0CHzYeWatYhNGDH1NcpHNLxlfjjhUvWIuQjggB9YMYPV+TAn+7B9eZMN2BJ/piCsRYEXD8Dr
/Fu7z69smWK98IzWs7fcgwf3ZrcWJdi89vLgZJcQPTnFnxLbmpjK9ilySQe6nOtaj9z1vU8q/lVf
/LFlDU6/nnEkjoN/hCjzdUXMF1k6cMK/5/gRGKm68FNnV8SQgMuc+e15Vh7hKvqJ5jncJoXxRV6F
V8F7adNhx4F809GMausmnd9MRioSCyzyAjBfincdt/CIUMiQ3jC62RaEnuUIDxdeK0FRLySEx8lD
CpUqhyVb0GJ8q/On6PWv684yg69Pw68q3J/oQF03olemFMy8zINDHdWlrzKCTXtxozgaLAOEaJby
4fXjKp1EXDNB4sQpOl8D1ZpnSNHQHbQYPgV5+26IRsy75Eab/3ZrvoQPlUrfCu5eoEyZIv8W6uNb
wlXM5klnzJG5Q03Fx3X9ijJ0TbMyE2QWB+esyhCTAj6Pg0rmDGXfWWmNSjIaCTzPys+SHQ555zq3
S7iFkABJSBhWpywVA5LrFiIlkjcR6RY1Fszh+4DgAHqtIgc/w8rRSD6Cyj0imcodIjf012LIwfDO
pcHC32ts+Iq+HonAY+PBqLSBoCOiw8oYCEo8DrG3nC0CKW65Xy74iE0YescRO+03PCrnkv3IXAfV
N8cjN0aC0RxBVbP3D6Xc79bWeVFbuhaklZ9zr71YdYv4MrXQg0AgFfLhC2BlLJTVCAqvopZJnlRW
mfRIUaHhLWRLq3r52txhaYpWPPjrXxLzUb8sSRxu5cseH6FEKurNbtzEer5DV70VZ2pWqvWD7oJM
f6g7hQKEeuEH52ZxazYdUkdCDCGeCrgZ4CQEM7A1IO5rX+4wHs024KGD68Y1DasiQtzjd2ofE9RC
QRxpKkk2iKOZkD1JEvFqALHK54QcOxpiSjhgkmxzbzuvVQ90qrsOQcSRGwWM7RxmOgYkFGMsE16M
Ns5QLBHipGQxZZjCUhUCd1EAldjKcgknsiYgaQuDi4zKpxQRpcpwtd+e7htd60vtE3EZ9CI/WW7a
wxCjTnHHADREQFr6beIkQtJXXZ6v1NycFhrKvmFJF5ncIEA0apZLHsUxmwMMBiJ4rXz4hTMUFZYw
duQPaDp5mthzRKX7kwh9FkD1kHxFM2LBPq15kqQxMsl0TDSjVC+D8aGp37/Lxeb9T/cbmSgfpTe7
TapoAUgckDi8hN3jqt8hqbwzjvGy3g00kvnJLY8gfO+6HytrrkZV7ID9aUgN/6Q08RBrebvdqX1Z
cgC2FIFXHPeZKl2K10Ty2yGbSBdldyIXqMZeFdEP9qcbT+J2MHb7LRhSmFDR9lmEI5smV2HfiiG5
JWsL2Ep5h/Vo4ONNrx5Nln3saHsABAmZufZTEgNcF3HplAwjSH5vC8b7na48trArmYqSQcwuP9BN
Ap3V37K4MzIdbgvOHVvL56vurxZzcP+Y/U3hvdgXNDS/+NKqHIUtf9P7JKLuEANBb7JIDtERUGNe
jHB+IZjrfaAUzjTvjvzLyqnDzV2Ub7fsO9xe03QQHwqbH3IAOKfYhK4Yx+UmwOsftYMcO9O82fqq
HYbigaayxTvfmWIQZ+oAPmhN8KN6S3FFJJKJaowLmgw4qUCx0rH+OHClSLzPkMsvB09LCUdWeCCZ
ZPT6nbhcbpYMhZb0rLznecOQscf8netnQuTfihhB9s4m7GXh9ApATdsNmM4CVeTkXrwabSnER/wH
aCSWP45hwmagR6Sz2bUij93Exiz29vOYRgG/8RAn1yhTnXLQtv3lmFi+quedgwROwJXFnePc0iAI
bVoAsWl96/FNu2Su0SdDO4cLXRN/KFma/15lnb2yejdEJyO6zeln3uOzzoKSnzvecIVg1f2ULuCf
cKJFQN8795LL9JlTkzlZdvG1u6t8O46MMKeWMbxonxjL/zD6ffSF7LvZwi/r3HK4C1lbEGawRLsZ
IoQL6q+QZnVJ7IKimgN0P14A4jdDKz67AnUyGTVTqm7KvjtTNpOaPW82mILpUNq7gdd2NNh2cwB2
N5U4lG4wtAZKpZZntTvCHxIP+n4cSIneWwUYU64aesCy1O5tc4MUnVZDZlFsQNqMertTbwQRs/8h
Eb+TXODFEPjmaUa3Lel5VxONBnwG4tKqG4u5MMUMyhBceObV28AnOQr5kaGUa0XkV0N0L2yB/Qee
hABIalV3JedRejQimPOdPY14mn5o6IoIKOKudufk2CIbrlwQWNfYVG0aRNBQza/Qvm/LYbicOCN0
76I0Mtbp0fAl8S59pfsSue1zZ+D8NAXgR+Wei2oIAhFKP8DG0+yJBHMjBo0VFc13RrM12b9wTkC2
YdTsoVBFk6qLp0chgWSc0PIn6iN59xLirKDBSdJ+r5ZzlgopsEmt492CCvbhsIwrdsMgVY3Md27H
rocdA/bhMXoKLKm/4tpOi4peBYJXB8+d+PxCDCw0UjgMACqzwi6dp68i9N1/J6xj9DAFph9kEJcp
I3GmOnsMlBiCDIUSBwqwTvMGM9r8xDakUf8hEGwHS1JuqBWqgTMuVloK6tC1fpGPASwTyuZRgS8z
TI7N/KG0OY8Rm0/FnxYyYm68J47suU+FfQ1n7qNJHlESk/8IKertl0Cu1cXbuzaf0bwBJAudsCyM
t5AGWsoBqD1PoCzJOlHSdYfgfR1whtTBt7Jg7owrFfqpsfn6/28KN+YrQUothYoUggKFKYBSlUUV
vVLfvBONycpYCB1GnHaU8V4Vadj30lUWNlfHBl7t8sXzwIg/ZkG7Q5jwEhMeinuPIjoRwLMYBQHx
v1zrSGs7mxJkVOhz8iAGi6LVlJ2NQIMsqIP8zkSaW7GtbQio600TnmNn30BI4UKSrEsOyF81/0/h
rR3QA38IR8LNe9KpuK0x50vKoN9+b0Dhngoo9oE2zhgyMYfNJMbsMB1OsabWwEhL9YuWNshHnARw
RMWbdZJDbOWEwJaW3Dtzgq+dqqayo6byXHfZFFU/E79NESqfrslvwvmZgsbVwTbsuIxfQttL4sMC
EfJSqD9JSDeEjP4xumGJvkthhao8GF2PuvFomv3SyzVNuS9ZhmX5Mtnbo2jvKmDF/raBQjJZKTXF
3sSfOE5EEs8o0qyN9RgGVgypDcSE5Nn3h6PqVWidvhgeVTsCRdbaMLfUxxXF4sG8Ih9RmTWVnYBz
0nNZlQfJoRRlaSOHvMjmEDJSa/NUOI4w2RQWnVZYgD3oxsOTjHRxzf8W41tE6YqIL+K2kCDtZRFQ
7D7e/T2zCq/wY0ZKkFxfL8580RqV147hsZK3RUvf7AHl3QSYp9JgNaU2XUuBBc6rsxzFqZxIaX6k
JXU3Q92kuLAZZh8f+ncUKJFsM8CINUxRh2sczHTeUl9dHsRa2fjySaP5Uarn41aMLFITI7ZOs7pS
BYQFEynnFUJjX5LXpt/bZPlxFJ1soCtgZoQVArB5D3i9CQIc/OivtxJYXBnfyiyoJEYdvZDj6+XS
Gadh2omgSUtgmKdEGsAay+kicxca/eIoIV8iNbHM7QYDXCPRZDZDhVSxSZyEWhRZgM0bCTNXPz0u
f1d3cYQ5ViSFwL3ddCUhjMf0NpkusO0DPBO9aJ60VTussySygmehejir+0DLDhUXlkPakulDqmed
R3HC+aKNwrhl98T/OwMqGGyPvxQ+K1AE5rokyquYxXfzP8UbM6pXebXJauoD54kEo8tGSVouVNRz
w4fUvbP9BctorltqxXavA9sUAsk31BkxQkeZ0+44FnrqUGpK68YM1DSCalKw9tfBMD93i5c8jT2I
CvhSvO000JvC8u2XFYpA0M3FtP66sypBmBLDAwFdhj8UtvkZzn5OrIVrorlLO51lxAaxzNsOf089
xbLzw/Jw/8yDLZPHbJAyn/5HHgAylA9mgTHKeBCk3T10Z9vGy8hwUd2bCDQwA97VCzYn+6HSafdR
maKxZgl+81YcpyPgEenuN5qVTj2mVh7ITflVVpQpdmKsTWgQK3a2Tqf9/bwSi1pUg6HBPOg=
`protect end_protected
