--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
hTiD4N7mA96OaoSGjE/acjPt+HB2Ef1IO6brjw667UeGPj2N7YPKhecApq04rrBlMJVFay10L5RZ
xkqOPMWx8/emb/hMixZnogyiWicg3SRAczMCGuRM7rv7AFThmI/OeBE7xhV0eM3W9uidVQnioRBi
7+nOU0cEvr9ILKGl69VMmOiuw5+5hhyJH8h++m0gZHMSjOTF4orOypSnnC71IAGV0lMWfqlV8oXO
Octvbtq2ycaSkGq+EFY91OGYny8scTYad5GdkremxlZUDt4tby8pnHW6uFaSGsIkdGTGun2CUHUz
kiYblb/cbGXVinSAaoYbXkRYoUD/yukHnQnj6A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="V9ToAzewp+MbFwAxlHx2Lcyo21iev0WBVn6/Rh6D1JI="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
aYRiK98PSMfoACfMWalILAatmC5LmVCxnW80l0I9rVJx4sZFky6uDgaVhG2QhGsNrTOahryQFzVQ
21iKOWLKfiWLt5uo7fOu6gNd+uaCFK9+zmEudrb9+CXtr4tsHHPOyLem1/WnVqFbyaS8/DDWs2y3
hHPs+JXzaC+AzXxynlwu1PTp5Acqj6PZhcR9zoEDzI4seFyIFmi/VMtpAbpYhJQrJGlMRGIPp0HU
YRodidZBicjnWz//IwMen0eClFMb1nnugWP2m0RcrJuD5Fe7NWFwBOiwVeOIkqQm3fngaWv02NNS
8H2bzC0tLpZbac+GxCW7h5l1ffSjBu/uzRusiQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="KVuIPjTa950/RH7qFAuWteTt0AG5pvUPL2Yb8UbOrCY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10064)
`protect data_block
gh9/V37D/Y9rKoCmhQ49z9gHl97a1M1zc42qhKZJwpYxSpPERC+UfbUnFcNKHnO/tiKlGJCsddDB
NRllBQ7BLy/ybp3bgQjKabuO4BDENVjEQBG/Mqk6lQ1ES14W9QxB//7lTdXSYg6DmzxsxN0a8NEO
JMq6bSCTvYFPEKMs96+yPbpbSJ0W9YsR6mPBqORsFv8XfOuvguRk05BuXNq9VkQumQBix79XEYLH
RCWAoESYIc9kqbcRjFRCT8YZZBw8LoQNbcM4yALXIK2pHx9geEasIZqC+GzzOfwjnLasYeaNB+Iz
3QSBQoTBCYyM7AiE1Nq0qhZFiJX1nfPLJjUbTuiBUCJuhu/9vsE5X61uNoCNB5oLhm6daz57BQD1
Pv78QF6obSUSTMidVl224T37aBDZtZ18lprIba+Y6QJbOUPpv5kzTWugcOAYXcUkyNgZhta5OAT4
zyevMonb0D4MvL/epM7sadBhIc5Xe9DP3KJQ/5TdChODjrufT3cc8VMLthuvvJIhDBlaEYVJ+BEd
lqRs940Vf73HJrvm8yEWCKhLd69A+PYHP78iOKfayUJ/6RxLzee0sKQqgxnf3TWTM/ANa8pw8Zel
1e9E9aPRDDoSByjamofoZ1jk1LfompHjE+xajYYWU4nXTpTxEgrNwTKWHKzNGAeMsjX8dGwd7J4f
035sFELz1b0MIYQ71WWAF/41L1kfcsWUpM7WkparlpYXOCxDZLPWRbj5yXMtB+RPVK9wLdJBePY9
8yDKMyryrLe52E1DTmQbTwzMncjG70GWhJdJCTss07lYxnYCKFeqrcews+EOIOPPRDYR8w6VuwOV
7WS/t1fN3HQSODIMfZONIVKlvEkgMfGTS6Q0yqQyS80Sn9h9vdY9aWQ5Fw/wG4rloj2PDfkitCcW
k/g+T/96iuhTfMw1p9vw7cPLUscYjhK5i7Ni4VzXMkENjDTNhSg++QkCgGrqhlKRcaAZIZ6CtSVP
fCFvo9C1YfCgVcDoVO5U7GxsXcjtu7ZC8F/eL/wKHFxehjItjS74C+I48w0zdOQGST4qlWel9TS9
0Fncj5lpsB/QqJ5sYg2p408ooYkFdly4Dmprp3greOquDF7gYPGpfPdAglEqfMnCngjoTp8XZ3Kp
1ld9jPZdlRhZwkm8OQDUfhg/wrx0oZ8gkqL0nyaKQkRtzOVUZArRMV6Kvaf66oCmfrebzpN9yHFu
IOs8rfmMkFebOG9Yiv92nndjoXPub3wWSunccE98ncSU6Hz9PCcdUcU5rBzPF9paIZ1Kp1zI1Rne
JI3U85Be9gSVwaMis2X9btdNAcPEBQzX0UpN78IymnbJKNjT7c8Y0IFWUqR6gdNv6HjKAKoex+IF
zkoFmj0ucczaGzK7BsSchStl2BhPtMTHUKfQR6GqrZVMpfma8avxXo7MqJkKs0KMUK/jS/GO3ksd
G0/7dME83CbA/OPG/D8nHy5KuzFHwBGmcP0GE58Jz0R7D3bNeEhBeD3wMdL+045L3ikSkizZvXtc
dXks5ZInniMy9pIbOxArHvYGIat9138mzDFECks/9Z0IiWoldXCBuUKLehYtxnrfUfODzwCdZHz1
aXrfmS0ITfIUstQmbI1HEDEHrhy1bYDJmV5n6YKJaVRIFeHkLdTzz/fK0JWl3Ku52YYolIJJbww1
jzqesyS9ldItn64QrBXbWlwJD5fQDeqF/sjY4OBeg1Jc1OXWikAF/lAvNnMAoTLacENh6VzQPaCX
iEr3l5phvQ+5BiBcq4URpb1bdh4/WJwquHzVBQhv+dpFx2Me85RlnlLHO4VNxvHYIsIGk8DS1Ivk
Hj8AbCYOGdZs1usqgq3sYVb37hUX4nnPbT2xlkP+OtJcXISdgwk6BPNG8GixNrwwvIq6yfRAQkpK
EhgUngeN5OcL6XL//9+cOLUyXaltnbAVwHhfvn8vezA2FPI8t7nUnl3eSFNWxIHmRXjhDzBhHD1p
dkWZohQ1tq4V+eZItoS74xnhtFJnuwsva8UwMxbH96hSYLCalV9qZsK3w/RYIkcRTRY3FIpfzI4l
877lY21jTjX2wAbcr08bgSlBPl7mYOJGpbyx1PikNpt3OlhJQqH25PIFwn97/ntu2L1JQ5TZhmyb
SXNIH5T93H9cNILe48kz/vJHjaOPkAxJflN/f4vxOYJJ1TGFm6LF6XHNIPIb5LmDr67GcDgNVrJt
RfrqZw5u/hf0NT0QqhJ0r3sqeeeRx0K1x1Or1X9h+AsKy8/1+HoW3XJ+TiRKc625R6BmLfgh4oAt
f01h8dCYaEXxJSEt4FlVPtUVbcPnfzvHtjdQ49NVJ7M9UJop2+XWGuJErTgKcunByRln28YsOeYy
g2B3tdnpqtI6UAlqsurasOGTlwYoRioUSHVq1t0kSsCBR7aCnUnV9NdwzOd6tGfKLqhY23QbJY5r
he424eqFky2P4F5ImoNTxXICenAkbhZDxUeRywWmkfXE6kDAtCsFLztFsD0vlve0zItIRjmzugwK
WA7nnSVW7ecO2B3xTMc4eB29rMceyWntVk5DRsDE6lNbmVA9pk664HVpvUwcJl0rKFikHqxF7+cE
dg0bDy3vRFmup7gyhu1MTuXltR1tcfaP1heu+SHxep42K0uhyuhIwgXVZgYzY3iZKBerX3EeGdC0
6Ujq2P0SG6zV0lqF2PQE7HkIvxLOQo344AYyyUpZFfxf5VTERGUoslf51/mB54rskTzAlcxEcfiX
kRO2qmjM6/HWosJMDPulJ29g2CVq5HUtWT2tWtcIadP8i6KDkzZvLLwfW9inexS4Z973X+j1Z7JN
tU1TBszqk/LyCgNCzq78NjZpA+Zu1eetDfVPjQeA6dR+gVsLEokIZGJe3a7ocMZpM9tTQcfDF4Ja
+X4nGhXlEMlL0Xvm7OvRZL/oidiZ4dFE80LX8sNA1Sg7ukV6SM8tAnccnGZ7Srh6yebhAcmoBX2v
Rr46thpJ9nPNSaTj/0cwOoP0TO1qhNBIT5+YvhClV5c0vBqsEVgSVU0MvW/fsMyrdUPRFmPelikE
kXHPrkAh8E9rrR22ffg3Y8MYT1+iWxzSGtx0sex80DpTl5TLTq11+vjI/Cv1rvcNAih1JaexTlLK
99YpeOM+P42VaMDv4ZJO02WzyzcN7FkzBLyZj5M5scSQ0HMiHdL8xuoS3OX4cyNlHMfKMQm7GVDT
3haSn2eSntp0zDOn/YhBB48udbgzEkeHiLa1LZG6kQ7yRUbqOeE3QDZD7qwybE/uZ1QiYV1KmL3z
Pq/60jkPmDr8nrasdEwfXdyeCLPM/K0XBLdTtdYTC5F2lIlJeggvMqy54f6uKjNf+wbT78KRr2CE
PrjwBd4/Rgj8NEt5Wi82L15u8Ny8iMODu7Z8CAByZz8JoCe/Vo8cGD0xgdNgclVBj55mDjYBK/fW
cA9eUigF10zMFJgvPeAkM5nDdqxIPeFd3cnQbMSOSw+d20aF+85fKRkSo8Mo2nOQVKPzanEvgqRW
XLIezfyip18bXUlsR8b2JyIbcqmOks5YuH0vtV3Yh51CM1xfZZ/W3X46wfdaSP/zP8HDq07juMHV
UwkaFpNTlt2aN1DVL4cH1BigSyKM+JV50X0J4JDDHfjCoEaI59MkFfWxeh0y0806LvbzH0hW5MqN
w/X38vODc9q8jxfHwu4eFq+rj5tLamwAyxn72aDrbkmojX/mj/cDyReTsQHHXW9jJI5PDTATR2Hs
i64jO/90sE/ka86OOG4FefYpgf/KzG16cGWvL/cxLCN1SywXTGJk0qgRphhe3Spbqy4haTZekoZ0
m6Vu/tfj/E45DMvpkKJbuevFEvHBDoWGIl248MZHqJiR4/sgANOGdv23PHJFXqKmb+R3Et4CAANH
ozqlBZbgzjTtxQM2PGG3qwuPNZ5ozyS6sMmF2V2UPEIHyjxBoied/OXWx8Rn7qCMHJxx5Y0WOKuK
BvwUASOfhNgpaWWDhQwkj3Fo9BpOnFbs+3wOfApsYpRfpm5CP8qzNWMUK/MobL9dwEp6WKWMxYTi
J0w/jvbiwVr20aIuMT8E+TyYSs2bqAbJhRVCkaQOHuGu7zMQojJHGDcCK16Enm7JIOJj2J9Qii/9
24A0Jo3vRdq722ShGTW4RdanhHU+EBYabVQGNR4jXpOvJRxQ1ZXzNIQsXPZ5I0ReqJb1tR+IcPx5
3A7OGaq5l2yB7xq3g1eibJTWoLiU2bYNJMT2200qN2jSRv1v3wIgrtfak6dAHiesaRgD5LPSlf6E
Ms3rzF0pNbtwgUP7Qvh5i5+xyVlDzj5xQ3OYcMi8ofgpr2DK694I0//ivJ12GeBpNSytPEvIhXtc
ZfrUZJ9bw9dzy3TBEN7HaA56P1kKz3+0Rq+p0+60wzOXM3mHXQo2DQ44ZsaO3lZKNOaJD0px/Y0F
kXHBFmgK6vpJN75nEMXtlTXGRx5KhWLtoImtumTzD4zs3Tjhtoji1WpPeZfWeYWk5IUkh8MZts0n
ErR2N4DQ4NZTawVs/kLdL8+RlitZ9jLSOOf/4D/Jx6f5ouHeJla7YXtTHZUorBcAkR8prY2bQnGn
W4aounjLccU0mvo2hAF9kpAbi3rmxmxfBxw7br9UbTk4ttqeIW8+cCJYeMHoPnQ2OVLhueDWVUHe
uB6AGZKZvNts63mx9/juIN7+zt3lwbqz5Wj/0qTJc6h9eAsio3klNBWlEC5FH0q2SMmp7OOzFI66
kfYIK6UuMajPUeJQjF4KKP3GzVY5Hwr8r1FUUQb3db2TBZsXFupmndOaGPeRGak7iINnjjMrWxet
ZhUv2iUNppzq5WvxAqOAwkAe872sExf1PKLklLJ3c3cu96Eqz36iLpKU/agitQtv+GtYAew06RKg
o9E5f5PLa8xU0QLVNGYXVlbmtU48zVqQTQWAdeFOWN0fHcSttwIBwKnhBME+APSda6H7dEu/A45S
AITS+1yJtVK0owdBXoGZ2F85XXVJMN7Mxd+/pvBI6IREEB+lM5lvsRu9bqPsPlgorG4D9Pco+n/i
TkGnsLuyX8wJf2Z4MZ0ydHBR8r0HJXasvbkwKjLWjdFQWzfRiywqKneZcbK8hsNeh3VX4u9xCEOw
8TaDqEJKaMl+axXzxj9ly+pP5Y5g1kG2rraBaoq2rthgkvIF8O+3rLBJBFUKmD+WRiNso8sYkt++
XXSpogz/k+V4e0y56fokRYJNUTgPMdfi0wvlEKuS5tEki0JWzdDQt7ABlnrDJeDL9VkIZiHhvANV
Vs9gNCKe977fgDFfIAoHc56jIAZu9J7SIC2wDmMFP5HqtfI3dk4/YSq9owpzLrmuUm9QsprCpeNL
V75Pxap0eENn/S9MSS/mqW88wXL13ZrSA319SYeDgDbtr4efJ326JilypTtWbmTEsBIXpc3MtdDI
3nWzWvhP5SrHwKbXv8/O4u7Teg6WxEoNqS+b7EHhjDj/YrLNeKD35m4E2CEGBw9M+IYQdXnAgGGF
MXPmTY+ULHpqAErotlmHavEItsMKOSbkDMExNbwMg+KcgWHQ9KtykaGqVi36wNc19UlEODhmd6x8
ZyE/eT38jOZSuZQHIQW7UFQLa11bVFRp8xY8uQan4W6EoojN/8jv4ECN854oocSyiOV6bMOlk8Rv
+86m51AEL04f37l7JKZXmVyemOvH5O0Q9ooe0WapLuTnFtpi+rcKalSxb5aA94a5Xid0+7TRE19l
dIXoLRTol8x0BfooBChR0aEc5DQNt5O7riaY191UX7a9kbPjh917chCh1w6+0YNKZuJdZnGQk5dU
wBSV7GSY7DvgAKc8jpq/RqyRY4pKtUTfQBmW7nh4PVn4PCsbsC/uunGLQdi2lzLc0jDtSOUkomBW
g8msYkOxio7+4VrWrrbX5wBq7SRganrJCCeMZ3p9NgNnJJPyEgaAdOfj02qe7oBg5aAPFL3v52AL
uB0O/h0KT3GWS1Qbb+3vWvCt/7AihkUuvrtNiVHco63n4AQL2coPdMWFcCsxTr9yxfRXsqNvr2jx
tVZ6elVjwASGxD4r7leBqc4gQDvVRCSstaaEN7epZU2rsXcS+vcIfVX3TLIkIN1p9mjNnT6zZ77f
gcNIZFxYa7xLrrPwdna8DNh6FvCBYd82yG1kURA1woDQEvt47hj78fYKBQCTI665KxilnLc4mpbZ
GFyXrnYI8DTXBjYUgcLPAPYZU0kKbItGOnFWNWrPPIOAZdoWMt9wOs/fpBH3OPgFc+N3lfh2J9rt
tkXuOVPcOGSa5woyeFE+yGejoYY7x6OUfaK1FaBJY9h5VfxeQDka9LIJltWZ8oEpDHcVYvLY2IW+
8klN8kLRzng9T+O78l/hAbPCEb9s0jjRFSvf1Zt0QDwtUT5pI8OAX9i2ACeMWB1gzNKWokm8eLIi
CBWGnVpDgxr0tUCqm53pOTsiDDKyYb9u7jQ8EWgI83f+dByBs0Ly2LJtRmEjNPHFNK91h4bZKreF
4arUaA3yco6Ftz7QGNBVDuYYy68tEhpZZN+2gEQ4e7LpcXSelINEtLbm72ESFdMQj+xod9DUTztd
nciQZr82OEsMkxGFCHN2bpNzW0AQHNf4csb/tTZ7uQLLBUu9EoLzskmK5Upv5DmNkwTeYdvYZKSP
h3HVZGVH8+HEu9XPHq9yi0a+Y1oYM6Lgo97yF9AOLukT0NvY+/MtOPZeXBz1AWhzB3rum4bjzkxz
i6PKe5b0qvRp5HzIkbU2rZyemGW34XlI06ZHr8T3H3TxW1zVf69rBs58qC+uy9M7ipkbqbuJYBS8
z/QDqBqjSBIfSe/uNC2ksTyB/ikJNmfMBznsIIgsxcFFVTiwZ+67rgaVpwsLrA2Dnhbyy1Xa5UwB
EOsJCFbOoZMc+/1+evFI+c428WAEql/S15EDgAJ4hAkDnxja+ecZ89UjSGVe0yLjqoPzjLaWNN6c
/5yI5w7nkfuDxwuFBaOmafiljA4rCxuvhi7lU1V88ngPLPRHYuim/Z6yTI+WUV28HJgwP9uNUscz
hIpJS8U2xsEyUFrSy9eHaoeJEiXeG81lHquKT/HxZEAgXJB4BFarOw7rW/0iCUp6CxxwLQXuaMxG
rV9qIQspUEHhi5lYRDNN/WcdyRUm35FhmG88vyLHZF0gaXfdbrFt6DQJ/sq/L75aR0AV4ufRblWa
r0XbBYrNWBn5CWjF8WY/zU1WqqSNE4DE8Pfks6iXKZwWMwrwLkULzYhUxBg6fmcSagG8++OGxF1j
BtozJcFD6EgL/GSUzPXB9Hf3J6wQvBLf6YxEgX8bwGe5rFAKEzNe9q9VfztSWUkym7cH2pl6Ontm
wlhn2joCNS3pNa1Qg06MQoi7BYCDCH8KRDcqYGKzneTQjdSPhk/55dfzeZRj0lY4FgjM99ngAoqR
6c3uUdypmqn7VBvX42zFG+FTaaPa+JNm3pIyDfYrgkcNrmPAHKw1MzcZ4fYtYy7jnhqeRZlRXY9i
KXXs7KKEsylUs/4pAtB7s5CFrNtp+cku4VyHluSSsXKfe661eoAqg5Rd2h59OW5aXq9vAU1P1Iqq
g7J4U+Ha/TY8XGTqNjyhyPveQsyaZ8jd5ofLIbaoH6goZwX2u8EtiOh2108eMBsmNr/DzV6A+xWX
zWzHKF/YrkaGEy3kcYUXLV8K/GJFBlALyhoNZ3hbWIDkJIRIiRsyqcucoHItN2yDm3vXkSRY4KxI
mhVNuXSgdlWu9OTq/OZrC+xNzRZLFHVPxp85s2U3NkjQ5BIrZEUzxtWE6LWUMTZcBUuot65e8hUk
t2W39q4NsOS6uwqU0yB6ksbrx881P89ltVbqrJbOdNeprX7j4LbpdpyIhGMQnpTqCiYwCfNgy7wI
x9G0UHEd30ThyMYGqDjkCKjshHBBHpLC1zvtcCLqUOnNJEwzie3SfIvFT8y5Zk2vT2wURJtzn1VS
Qxl/q9FKDXkTzxRzCK4msoMi74UNOVJTBg09Re20Id9K0G8G7SIBcGp7TujHszOO06Y6MX0j2ivu
nHxq4OmTtD8cQeTCgddLEuAdppXvDFTFHCuSQeXb6YpaMEKD2fTTwMqIaOJthvGlGUDpzGW5a9qD
xFSxJi8BM/UzDGMPpy+QkoX1hSpbSvhJA9/zwY+TMo2je3yeMCuvsc9KKF0lNomFwCT3+VsCyWQX
73hcoN1e7UUAQkkIGlQx8XTwnbRFcAnsWDkSuIHcVio9hw0HRk6MfnbeXJ5JT4wlh10dHQSdA+PJ
dde142mLELLlkumQ0Y5QO0P4Jy27ZExQuTHS/i5cC3pfHQus+gQZHOGl7TW456Ku/H+9N4TY3PMS
v2U4FGGHBlg/uLR978XUNkyCFJrHxlsnPz0Py19gSyXGqJjDt2AV7ZHWxW6V8bJEvOA3LTV7gMZF
bs15tq74/TqXtmneuUYbaRt1zTvbGIOO23xR5L3e3WyWJ5+jPwI9lmNN4nkHkGUF3lxEA3XwCrez
LBPJUJiICalAC11xyt5+A0BH+y4vT2692xyXpmGcNMvyzz4mAHRDfwcTa+E6RMo1jJTx5JgKuASY
46gdb1QWulxq+WvuomaWAbc5lLAod7TZCJOJJSu2IcleXAUW/mha9lPD99I/WeERG/wKuCqNm4hS
rTMKUMv1hbiu8WGOjlDqn6cxdnAAq3TZUl/IFptRWDl5ZnRf1SABknXEy0u0NByrLqKaE3vaYlvo
lTWQySit4ujcgHFFigaz4mA/uF70LVxb8cZa/5r35BLGNwx6jO3YyrOhVt8FdHr7AJbPGjp6R98Y
utRMAFMajiojN+09BgDOqIWIyWCY5DHmcqo5VqsOjoUXw4Yr6AE72i+jfWj+8GKo4FgyFkJBmyDF
akg+0oweO/UPXa/rLfO6ifpv37hzZSqpqHe9MhRWlm8TMMbwQ8eWtU9FDSxTk2rD8ZnndcL2z23q
TNiP7dKOfO9WVLpWbeXgX6zNMpj8Kvn/MH+q8H+exzHsRDN1cwopzQC44BRO+CgLQQTy62lsPK+G
4FGIo5iRZx0rRa9hdTETOn6gIuBqSbQ45UP+Te14IR394qnn0M6iDeHcAcyC2y8QNUPuM1aODGOZ
O+O2+OogLbSYNN/ZWiCwniWM9Gf69ovWuwtXrzkE1C/Q/Ih5vC9n1OF34pe9qMrkET3HzqDzBykt
Me7FyOWkT59fAVHggk0r2SeAV1ItMEsdHzaQyYUQ3TlhPI2UnXIjxPo2ooY0clIIzkPWX8tcWWUz
POAd8Ygy/5pbJETMjY2BAY4Oc8svPMQL+rpZqhoxifp1mKgH8jzwC4sdRzrr6N2GqMyz3OEuLlh8
iPwULilebnOJb3VvPQsTlxvoWlB8qz09HAdyAt+zRmoCAZRHRw/HIwQ3sqGTazLL+S+CqLt5TE14
Of5kpDI8a0ZcYdmKKYDgKk2vzyGZMK6nNQxixdoeVUyAWxLkUbdkE9XjV8ICg4gVpBw1ni7u6L6S
hXMOafsdrXvhMtSNJwb+5YuQEIXZ02IP+w5Y6pO+Es0aoTqv/QHfmC49rWy3z0woBOP1y3qSo9kX
LLBclrx1re5FvitEcnInXvFj3B1R/a+Pnzmr6eezQGn7B9atLZlXJvTb0RbyO6uwylnLHnhOWC41
njFt3uWosV7xBRiTRhrzGk9Fl/U59BmgpC3TZjo6mnYsDsJ/lfzbTw7zzYzDackS2PIvsnL5ij6z
3oCdkQZ0EBTEHDSOXsznojQUtvRddVF3noNFwJbTa3kABSO8zCzcyoMpAtl1a+J2Gq9SGtapjLZA
oHPScp8wPlZVSS9IEiX6W4rSxAc7evANhUwIo3ickOgt8reNzv93ARnEeWar/a3n9vc473wbagDp
FgPuNiHSyVxC+dZnGkXXtEIEzPrQRAUIBwz4z+U4HowXMa4ofiEWOMjeASH2x02E2bOAuaS1Pazn
0dvyIruji/pI0um/aZYDsIUSkvmRkstzRK9P7mqGt1Z7Zgz73QUofTrJanhu+P/tsi/BUsEpz37X
hbKdZvN4yw5L77TWpIL9xNlw7NLcwC+na2gIshLzusTo7+hjVW04t1y26mm9fvynSzg0N3uW0CtA
Xttcoz43avqjmsfCou9mbYGN3FghnVn7YvCL4cc5jyjdyLXpsCuYSGoxvscPz9DklIjcj57JDIj5
eDMxgCKbNKaVSmJ81IqIpFBPVOkowCubxcjDqTMTAIfTHrkQ9KdMjqBE1NyJ+3+Q+LbA5uc1KhEr
rA4+f2pEwnuwvIJZkvcmxqvW+YFV/PEBS9tTS4vY2zoml/pzAFtKjBiQZIt2hs2sMgczXH7Rh45Y
iLQw3Xq8sQxVeFrUlVeE2ftXnHobiGSvqrh+2a5UecYAo2S5hHGFB8KXgDSrjF0DD/w0Tgcdwb0E
cUFmD1NNLUV6aBCMRyGVw7dY7tUPAbgxErlgL2dgvftaUaNcQshb4D7FnWrQPf5+L9gWFbBS1eLH
cdiPBGIgAff8kNLYvtbIlZ9mesUaP7cmgWw9kEAvKEBw8IDTggk8daAIwtNrt9QoTu0Y4oDzMl5n
cgOZpJcrSoVTEiRMZeIa2xQ4g0R3vaWcXQmW0Rr88AeeFKszsthCeXQwnanlTAgGmgy//FGlk0Is
4hkLfjxF4MpuDMj0zqvyYwEBb6DP3nkqu8iWFQSTKC8PG1KrczviPUjgrZWeIuY+6nE49D7Tu+Rv
jFdBpoOKFSHNCH6iEPCPkHP3fqJ7D4OyBVhqdfv1Dxkm1CMCPwH49Vk8/6rCRHDfNrwUtTgeQN/1
awXWWAb3+0zwUS4Iqxe64vKf1revoOOegAqQ9TbHmalDyqNxaBCBEwfUs6w2yiRe2MznCUNt8fQu
caXFnjmKe2pn8mU5RXez1cHjgxf2157rAevqzdFIh2nYWnYd2ba43vM9suYoRD6XPE1uOIlgPer8
u1s+BFgdPd7jGoXcBkdaAuyuuQ6nc/1uke/NZJxemlml44rhnYchju7CUOUu/dLT6xnkpDQSSz/5
W09P/I/saHp9Rvi32w2lxkZKrYvDKo1iweaP06wn38acSsTApBYRy6WJsI8KD3b15ZMwBl3h044t
QawBeKOiGvZigmd5kmErg/GukThrdjv7ECuO5xEG2uYv3kOkTuye96o4ul38ozKrb83sOrKN5UHw
odfWmXXgLJ2mvm50THSJwzrtDNfeDo2pCWxVsUZn7kBQ6CqSqhV++oC+pKKSYQuMaxsuMCyjIshS
EBzidyUtKlWWClodwQXW76Jqi5ew9O2YeCVrJjSchADVCTXnbpcqy0Gj88EUqAxeCENXbzxfkfw7
5q3L6DjppClYeVUCvzAD/0xv4vFZzX+hwu2LLJ4ggiKeSBipSbcTkwSUtxjsLJ+OGhftuo21fywF
6OdnOGLi0Tav/uraBYRF/RBfOZC29ROTaRzxg8ekBhBy9Q8nCspXzu1pF82dCOrUH+p/Pqwn7Wnq
cedyHY31uUMgm59/vCBetPJx86pp3yV6+09NLIedGBWCdnaZ+VfSsiOtK3Gs5gvbCWw0z1XGKB0T
iAayrnAxyUNmKpAjF9rKXZChvFOyZrBqDLN8dAPzJo/O6Jx8e/hFXUzbuUgFfxC/UBAXwQEaKo1c
g47hJhgbHSdX09d5Hv8YKJ6g9LlSPJx76ENjq9p0cKvBmJ530Hw+39hDK8mwx2mjJ2dowjdRMba0
rXEkJdw0o34qPT1jj7nUInHR5OZi1kEFTHe8A+Kqv9RIMyiCCRY4M268mFEUf2/SvX12gNcBDTWx
Evn5//ig4bKHuhu8jqaSTEqUxsMyp4b7soTKDXP2ip7aUES2vK78aDBblC8Igh7uUXDUWphFT4SW
yMPhrLc6YZvvAj2Jtgeq3oUp0mPEElywA06yoJBsFW5CW247SUca58rWQ52tkOFfS5iOe6lw4nKR
g3aoAe2Peck+s7rZJLWV+swu2vbP8WWMDmuF8yuvKU0VZNNuYZwVS9MHidkRjguebcoSWeRdARb0
3GIaUgSpbrut62NlVd9XU7/xZz5QHVqDN2LJZS4qZprx5JcFCGpjwrT1YG0+I9Qk40V5eQjw9kHA
P2zgHcBHwppbRA6CyQuJwkX7SSu0PEgFdm/2tCJzvy+vJ4iP9QUzO+bSBEq9naAx9V1G8rkB6hWw
IzdsEESTgylvsAsociyWEup+c081vRFiMl4Vrj6tKUGrkMcA0Zhvk7ezhwqkDYZvZVdR421XWsWd
h2HlQ2UDtG0oE8qVXBdv6UyK6GdQIhlfIkbh3SZKuV83yaNt0PBx0Qm8ccvqtQ+Qrc/ACH8kMWoB
5tP5wBZCeY3nBFzt4boqlEElxX2kMOkRYfvMUCcUtEPUQGe0S0GDR3rtFy0jum7o8Da4NyHu66E4
kVgF3NL8cz4f3nz95ALnuj5w2t+B8jDc5hfPLtcszhkrbEYrtyohqoseHFQNnaJQOtdQX15cROZu
IsEzK7Rnkyxgvp1WQUDrrEmUEbb9Xs5GPwajskItw/sauJ7hD0gLVT1TtEu95GtMwHIOY6F3phQs
0Re10sXHx9dRa6wfQ6ZrUtLoU/E4qa4uCh7x/NbG+bSuC3nSppfbvVXewA1d9I3qsoskUiYk/QTB
wVkpIBTQ5lK/Ibdy7b0yGRVhGN5VCVn9CoaxenOal7Y0sDWniW5BQSwVTUtJUsqN1I+FgYJhJLix
5Z5jRCJ5pLupYKp7hodcX52l7O4sGVEfpSD9YB47TpfD08TDcgYe6obytcmZ3IgceBOWOHtnriy2
P6XaDrDqp9yer9Cb7LTap9K8+qDAjChpeL8IzTWl7AZBhTzWIEJdve1/1n5Iuz4Wy+1kqWuLiHL6
LOOghJVWez3pBLJkbsNbm67hlK/jVejhEAJPBFY6OkXwWbakHpMWHwMFH/nFcVo1CXe9qrY5cTEA
qFOMprtjXJdMNkTSFu0Ys/sYoWrq529qFe3I0sSQfIZ3PVtBlqA9/Vke44elmiKiV/iyT9yZ9zUJ
YrloLpoO4iLnXl/RbXf5Vyv1Ur0k1wbYX8m2AlNbt2MmBhuUehG8VxxEMsPQPKAe/wheGrP0ns7g
FC6MNT18Ie4I5OWvoacG3mwMlHOJzsNCWVEC93HrSW5oBJmxrt+gPi9BoZguDThR/rVJAwLNET9+
1NhxiXcmyKWLul/j4ryHXfofAfL2RJG8NZRxNkjZODb5XQuFUsSvyOH9h1eY2IGxvkvYIl7AFxMv
2uZmsl7GFdQruUxm2bmLeBA5uwuHeGF4nHY0uEOrBMbAN4UKVlGOqMY7EDlLTGjG4HyuCFx9pZKR
fUqvscIHcUqIF1mBzWTpx57BVOhILWAINcPaJpipUtxmQUJDyF5VhSeSS9b6MV1VIwhlqUMx45O3
qGAySxsSkHLVrL51ujDk9fMb0yo/V4tKo68e4LwmuzaxmboP8UiFOypjd3++cllAXEsYXHhFi6Du
G63Ds1hWhEKWxW/fxMdTtnbBoiACg+/7XB23Y1FoHy4=
`protect end_protected
