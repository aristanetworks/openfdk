--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
jx885FhsJ6RG3/aDHTtOHDVbMBRNbdVAIxToyl/Hdvj3trwHnH/rLlQWb9LAUHpGv74ethJcpZVh
mvGjR2b9tlVtZY/HAnvcwXvHo/QbpShV0Qv7mrg9mBLn9mbAjCOOzLGvLPBO+o55H3hy+uUSI7P9
l5kLHOqHsqV9qlNOwfanwZUk0CxcEJjAotnuIRvSFr5mxymyvEiwkEXntV7ueDs9sRXZ36TWKu33
BkitdADtwM/nsFjnAVhnkq4uKSycFSQiqD2RjvQAGLeEiB6Hezv96jm81xi1QoKvy7j8xG8PJS/G
k8MYUSz/BBhvD+lzr4mmw+LXE6OWo9yyMonMSA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="XziLppClRThsLCTTls+BXaPDeqMV5v9ivnrUICVuX0s="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
jmlvH8tePQZ/6OkOFUodsAq35h8Y4r6Udmj9D04Ruxu2HEhHz01J7PMAbPVqlCB3Ep6Z0ExKtCMd
X0m8abYbkxyoIW3dybjwWqACXn+gSlbwFEpQEKISV53dtqNkeRgez1SlaWLzmcxNvWqgJnYA0CO+
74oLLffXnrpvKBTUOFuyLWluz4j948QS4tXDtzJTWaMpiSI0YJGqm9Ibv4K7B53zkZavddwVsNni
kCWNyrS2N6ods7si0O5JvO6uzv2EciSN9jNIpvYePeyaYQ62rkQiEtFc4breDrwwWvmMY7Nj9boi
03fm28684ZxSoSiMv4C8vCrilglxCgQ+JJvFpQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="wCLL0+6HSX31MyVZUROhMFCp3K21P05yfC/pt8ygcpM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10048)
`protect data_block
KNQcZCxTrO0bisYixTVRENGRku/F9j+zNhalzv9umW91OpjsKNpRd/KSZHJyBT3dapWvXIOpv2m4
qxab2sAV6lxsomI26Ut0pONRgK35r19MV5SH9wxGtUIdsj4huyNfRkywOiOybct+Bgp8UGHexp6D
LXSF5+RkCcd4iPY3FOQ19XqzfXY63l8FpFXwPjTYB1s5nzQSfHp906HFvNVRKQM76emf2+U3dPPe
FhS06S1wopTXWqgBahHKTjvyA1rcuKuTTbvn/nYcAnqG7XQmT2WHABYwGkKLKSrKcQ8zsc6WhQaS
1z8lO7s6K0eT4z4eSsHXxndFLZdsAgyspot57ZAOabU+cjU0WqNYmGyv2G4Yajawng7alHJuYHaP
qbneR30xylQ0e8uJHgccPZV2bNs73dJdQzSBmGrwZhu+KyE/mJJmbGcV5vVfF2gBOCtKn4S4pDu1
7EPOc71F1+ET3hfVseMTs/hAhGqjOmoo7qdI9k8Fn43S6EG/QRnN0rPW1KLqqYl42PhSkR7vydVv
/KSlKUIQPmeOHibAlaZdtleqeJRmTAYq45e4nG17YoDgMek84cqBNiuRtlDxRkzmPffURTF4drDB
PHJd7m+IRxKUvdGN1YqXA/lC5p1XBgZuJwOx3cEwliN0fiBnMGvAw1IdVEmh3hv4ZyBLp3fwrfbf
rQc6RAuzT+m17hQWjOLLh9wB56HF2g2t+XGU9Vy4nDiyXKYyoP3vrtZvQIPxuJuTqYd6wxi0Ixeh
RoHv2mKs4Ki/Z/mSRPuqvq7BUVIFrginpqpJFRmo4iFED5UMkIwlI4Del0EoN2E+8rDZ9J4GGLsc
wm99R9nlR40bBU3AQLYmQ+XEh9JPGhbcdokB7dWtpIHSEHsSPe7EVz08dm4vvVTknnqI8ZCDDgHR
8FO2uwa1mcUmFR8aVShzca4x262BGvibmosZPjjw/oF+5Kg9KJXiNec5IbcgmMeqJ1WlQDrpddxj
F84qVOmFmqm7Z/QzpinLZoPuud+wQAvZ+CTZxiifZkbVTUczzZRk98D82zMfUowNtVEOGAl8niWe
yd1zow0bWLp6PJbO4h8ZpP/ZHA+t3Gqo4QpDJDKdtM2vaT+vbfelUozjWC8jFyieQalTFeq64IaY
H3lFmAq/mXN1D3yT0If6FyQ63AS+rvo4oVEX0rJdPkfPg9KT+X/nrBThpE5OpHTxglp0Eo/ssiIS
aYujgaGLfeORE5I0BUQuiztbsEv1ST79UJaIX+d8e8sfWkDLCEqgTzugxcJ2/i7SpN0uOA+hJsUt
reR463Dq4Kzk5ttuKaGgIu4UTv/H23Gh9kHIChyYNvKq93405ZaVJusFkgWpD8B4OYrPVwaPggN/
xsyyoU4fZv/7tOfTP1NeEmtp2nfhsFGd43qiR+VBuo5nDQQRTixLIG52seHAkL9zipdJYiIBaize
1mtyyX2WDzMChLBrwV9AhwxhgKnEHFQOCeAJVKVXCPsPXeRkGWxE1svcWInkpsuCeRPPz/Q7DPEw
U1XmeMWGujbVQGWeZefd/nH9R89vxKoG5Gtj7Dem6pDhnqokBwAlQBou0MXi1vxOHoCymziI2r/A
KHRXGzFerwUoWU0KL0TZYo9TY+fx2PYEwPac7NmR6oAsofk10bSw2N3+p3qW7qOJ4qFE9sVbsEOD
JmUfgILpuX1xsvk6sR7V9OUTzF7VvZ66BiGnW9TtpBJmVDdTE9Oc1n3Jfe6ABiK72vs1VwJQ4R1H
zofzGB6lmr9r3dsP4leWuJe4kffyu7e76LhSarKsvDBdJtW4qv0QPGvi1byIb2IWS/d4enS4kSMW
0+kdijfh520ZdyO9byYPStdGaqErE1Becy21fDMfiuD/2i4Z9jC3dyUap4oSwcYhmm0cKPrxxgET
ighLVIowM8PkKobPBGWnYqCU6MK9fyxiMTEr2uAz0VWghoXoi/uIfluIz7fyM+XbhumoUX640UU8
jkKiOp5SdT4e5/kW9OJvs6XktqPTJROU5f764V5B29Nnqv43BVwfdg7bCKlCJ4XEsxZiM/8aPsDL
VmlMKW/YvE9aVD2dVe2yifxraM4VspwP/v29UPjQspuuBHcKGWQnpFIpnX+dV9V2GGQRMizdFMWe
ISYXhWCJJiNMZ1s3BxViwgZQNxMhHsSPHzn3lQB/gH9jBKY7PET02gIYRdEHCf7ifP53XBCuVyQI
L8ttFOyDDuuJl4iLTzTdt3a16GCFdLTW9CDeFO+aYzqQNWDxeORRSC4RhfRuBMM9tb2TbD7G8ONq
mz4HJWywOwwH0/84vcoYGby/YfXXhgEHXalaDLPA1Mji2tELMsYXLZrTjzwLFSGHmqS9jXQeGJ3H
l2QHomfj2+uriJx2S6H6/z9Szdyp9AKSSkqTrN3le1WHzvxbdGQP/kYlLj91vDf2HU/K3Yn8/Nm3
PRr1yQnxHufZ8cxf39Oaztp30SBmkLf1eI6vl9+RkceHMXrgu+Jm67q/5cq8j7gevJFU8BOJCWgL
6KSebDMq6op3Z+ygCt5+OjQV0l7/9bLVN9e9OmPM6ZZxEaurttPgA5tSzC+iY+0QuCl1ATmDTRE4
sPaVYbBDQJD/ar+KJrSkBvzHVwjTlufo0PUl/c9eC9fiDen2oRNrLsYqNUkiBrYgurkrJn6TLsrr
sUrtpEnIU60G3jFUYAexeBeFT4RpRRGqM80ERWJ+PS8K+SQcWpXRmCJD+FqvB5cYOsSOiZvyVqq3
33Aa59E/t+ryP3COUlzEawh/u0sw7eHrnExTdbuIFn5yynXkQEl4LZhFBRvtCXes7U8lQuBnpSx8
2dQSA+GZ5PewZbP5ex+jdCA3tFBLAQQaHjyFNiwwAsYHLZDgU/Mep4jbOt84iunL2jziFhtiKGoh
pxCod5P8PqQEo87ABICejZK5k3WAqjpVazBzhdaT+yeYPXvrdgOslgeE0VuNxcF3Btktrh1ilR6z
5zAk2Yh1Ul/daLX5XJbA9kc8s19ckCWSFHTFbQwOcg7EkvI7Naji00taOESeVxfPWz9OssZEkBOa
Ji323okVgnq0hEiQnM096IoUdaSukmL20OAVgjypo3/E8FeupLrxoaxwjfnQe5AUHXVhz1/9q/cC
dXmSFnr6Rp2A2VZ4ekC3TdPn4KHWcCR15lfcn+hw+jodxKa3sIwBbeW2eE8eK/PeGfnzNt1WKzb7
gbPtkBiGDp7jIgy9z8Vz60sLqdErgoxjFy7eyqG3kWQmqOLN2KuZMQ9PlnZBPwOIIJeO4TiNO3pp
Xwnj9dNq8sGtwDmiSUNwV36MCqmIuzbOO6boSTOkD39vn60Bv+4jemf7VdXV9p5tDwngQaNx14SL
eZrV4/kEbXh221wUzHP30Qu2mlO1CrcUM5KiXZgm9AGYCy9m5xFbNgj0HjK5ah3BvszvV9vQxaRV
u/t8mhtX5KBS1I+GZLxtZ2fdiJSksGi1iFvL+tl+eStv5uUM4KTx7R1guqKvPD/r8M6mP9CoOd/W
pDj0zaDHBds6k6Ypqx60ZjbCi9X2bXCwV2X3nsNYe+YyQAiofTPPEPW14x/o5dVbTCqhsC6CFrdZ
CTp3iKduzvVOx+7GuAcS7doicV8TAD6Y5KV8UXqRAF7RFo5+cX8E0FLsi2o7wF0cJ0mN/RpVJU/0
1DQGRinWk28RiH9ZpJ7CtRz1ojih1l3HPykaKgXrPFjfdZrlE8IMesepqJRAc93YSNr/PRl51z9l
K3pgKRGBikP3SaH3pxBJUjBPe9e4JKWNLtFX3OrBTFV8vY1h69PqnLfzYYuPcOLJi11RmFsEJvaZ
oo9BZZeoY1oHEMpslLWXtgOFliRb/5bPfOgBRA9fSn2gsiazr32dOHlRk7gXocOTAoSwsQniSTSW
zbWn3Yp19WB73ChQOUpR8ue3N9eoELV7p8sjbSSYjQdUszeOlG3yh6X8I4cz3YIyESnJoqwcOhd/
ZklqDpnd7WzZN94RnncdBaDGMHW4AXGjERhSeFxqxotr2c/7nN5RzflRqjjcBedgHyg7GdFWZy+P
15EyV6NKFOKLgArRW9P2MUMrUkg0pDmDX+PErVrAIPJF/Nmwqpes5MjiREgSEesbnuMLbmAW1KPl
ZMLXH3pi36/vU+FPOwtpBWHwGEw3wnPzY0mmixltABxH2lDQjFXo3VzisbwHg3lOy6yKlBXq+o2q
GNmY73MA6k5RldutIgnzObZDpXui9uHFIu2zl6mBEXwQ/eW/U6GnS+EhPxLR6Q2QsuBBw81Sf0/V
Lhngz5JQ/HMMN9n9j+p+Hlpp7Li8arSv0pKZH5uV57V2heDtQG69H6Fu3Hn4zjRj3CcR2gYqyEtF
a8BDzKdlTdsgVYVet09RFl3+wvUUJRzpdLDqihcHaFl1AQJfsQYtONKecYoEBDTUnuTsa66whBWY
ZCRhufvBDZGsUAeXt5m5a2f7z+nkJoVguqn2KIxFDYhM7N6PqZNHjnQGTFJIVrm7wO5ny3TuU29r
N54oUckXm8hFbYYOWwq2a7LAt364dYrTzFdbKDKKalRXsju0tTvKiBMfNXlpTHyxdki+0Da5yPrO
3LtbE236K8jRvEPhksAcU/1oldbfZXIwDx2caZub8/Rugpe1QLCMMU8wmQgL1E13Fbx1F0T+nMV6
snSFqvgC/Cg3yLs9kLfsbKAPwMPwo1pw/OAzlwKZDvXAzrUrLb7PqgABCzfQLMbp+f8vuncH3SEz
IYqpVYbDKQpJ8TTgRW5BbFftkRxEpL2OP0PdBmPnU/1lPUBGVMlNZXYSQxIbYOWosxW9A/70G7Q3
x7BFR3Pur1izspFAk3XFghVQ8g0SNsb0Fo2RgsWUldv9caZlbRqkjUB3z1X0F2SefzmIZoAJKhHr
jRx/dsUIt9OfB8+c9orXkHS+pybkK2hAoo8Y4DgC6VXl3ZI767JPOr6ZRFXsRpprq/JNDghKaRl3
uWR06ne+Obu4zDCfF/378E+DvNsHasb1ulzpfkn51jK3FL6nAz0KV6mrj3jz9CrdIysCFZNWSrDu
t7hu9yJqvCY7Hva5/Wh5HvMQYBGPmaY/orEitHHYRDELftqKcpu5WhVkQDa34MgzuCmU7iEDHfJ3
y16lldTJguAFuNEgFobj1C5T+lWtO4nkeKWr0UAY7GTYpc97gFDrEyVJmHdHSnb8lF/RvBAkwnOh
Uy7n7wkZkJlYKSwgujguHUQNI3JgAllku1kMGLRy4/U5IhYt8ax43u26dBdVvJ7W45X1R7OaFjs2
OdsYogLiKPrZWgbuH2xbwWNWxWa9gyDDckAsceIPPhQ5i4wweSWbUeGhCl/wRaGIjC3W/AHTu86I
kYw2bwdinOGC+fh4yPz8IKVFhps+QYk3TJXQ5miKnDoQwXsZpEzD8TIJX8TtRSpM8p1UnGayKWMj
wW2ii+XEoha5K50ShUMeHwyjdu/RIvJKsiXX03e6CaCNooQAXGWymXUDQ52Yb1Ci8rUMtLmA58ym
3thuMejZmdk1Sqmr5ZYZ+2hmBRUsggfXrgDlPWyw0aG2uyFlmLSUJGQ/M7M5SqCwgVHAzIL4LMBG
GeHTSGcT+CmHMtyorwXJKC3Ixk1F0cdBI6feTYgadFMvMukfq5SGba60+Ohtv2IjcaUInUYDXYz1
OKyjG0B/IeQf3JiVeO8WcbCq8ZPPdftCYHfHl2WQaQOkE/GTOSGx0qVZlWsPyn9zy3vC6sLeRLop
nUlAFZtgXKlBlvvsnQ1t4Z7g1EnHqxTFTjbwkD9f6jAjphUEl4DaqN9+ANBG8DSyXtWsqy7YGk/q
Fr/0yuamfRa4cEdR6mO4JazmJo+2CUK9Ry3wArQOsEd8mjc155VfREXtnSpyqoMTYMvtu9VxMgAY
1CjQtlpsHn+2q+4kd9MMiPZPXgwP8HJ7PuRbKsN8bPIDGchtwQYHozsqEyDO2s2cI9pTu/+9oGJf
//kbQZbK+zid1Y/8SYMJX/ZxOgRHWoP8/eIJ0EyIV45yV85YmzCbXemEbQZ0rcXNDwXOvVjoshNg
//KFW8EcSMv8tTkA9UzdEN6ch1qPIz3Isq5jrmluR9LJvZl1bkv9uBqktCpi1EHC7jdKJp5hUHTh
wRqSxn5S3EZch2QvrG7VAedNe9xe4L2FxF8oSTs6C2OaYt5ZQ3dfXGv/e0LBQVyomLyUXt6PlXcr
cOlBxwIpSssDiOJv9gO3fZJdir3VmjXz+8yktT8Rw8jG+NoF7BMrVY2siVKo+Ek4HXkcbM+z3sLR
vGfdL1zGbHpuzXoD1AL+oDd6+k8QG2oqdmdbXYxSTBob7FQek/9LcKmMsu11bUnO5+QbbnXU4yAz
7vH++vZuwPzi8g9eh7nSDucn+eu34KRekm/SfqdwCgYvJ6B8hIxYZ0e8TH5STKsp0W1Vb2LxLvKJ
4fwaGxjs3eQWHlUiQDiSLWgaRWTq6/NQqWpuOI8LZ+C/GLiDO6JFQ0CgB3AD0nA8LCwWb/gGS3HZ
O347GHpp90ydJAWObINlZilenB9GmabVpVgP1HCCXjeDsNPSopC+e5pcS9aZL+ndLlnGy0B+G9tI
6oPgcWyWbh82GsUJMZWjOw6XIdEbFV4QY/gmcf4rqjjU0+uahLQEBMUCi0ZYdJEJQGEdmhwdvLcC
Oka1B/8YpSWzkLaPV4QMGjR72tsEqOIYa6JMGZWaN7sd5nh09kKPsn3Ji34s5o0tuCtkrTJXg2Vv
TuhiJHN4JCzzlLKUQ9e6wIJNUxwQxx/rvVf9GdW0cIDqNmWj5Z5iSeLF7DUzWqez6loi88ORpLUD
Dab9ul3bcD+0QyHjkgV4PMSBE2/XNX5C2AIff2iqKUODe6R8TOkNFw62YUdN+LhM+aiWtkSaiMYj
Z0f4l9hE3Ns08PCnBKlfPo96v1Fz4zO0Apwez2K+vWbxgOoNaV41vg6Fnj4AP2U4KTHaOv5guIo1
nJT16cKdIj3stKY+cOZxq/g2nbZg0vu0Ex7tiDKDG1B+ICZb1AWir5LeArae28FHMVpUCS/zR6ua
Az1uOx71BEBS69SKs5aEsC6aRCqVViAzYSs7uRCi7jMYrfp7GqDDHizXhUb9P42w1UPv5RvuhyWR
DZ+bJ/Vfpf8J5jitjFT77lUvFKNJQVS1zpsY01PItSWbWY22bOAeWR3CCOfvG+7FYNsh7ln9j9YZ
MnIj2uxVrD435aR6pwI6PPQOQcBe+k+YVuoJzEHRpit7CU3sniwKU/8WUUPXIngtYbJxuUCbGqJA
TUWbuOegL9MGSv3O3haFQuCRS2PmMshztDcngeB7jryXAI1Rcinmmye7jJoG8g6Y3XkFjE0xecxI
1JDHZQnwlOJGiVQ0htn4XoCd4A9ytiGMgS49CjLrV0izM/NB3zW4e9v+7MFIpbrUOVJ6yaMWaqfj
8KZa6xeJGzfp5ORuf8CC0/EnHoR7/vgTXXPR9K9JeqeRVODpsw4MKzGjoSKcw+otuqqLIceDNoEM
ya43SPDKUkf0yXTQ38a9CVBA7ish5BKlnaFixYzehZYCer6d9yLnwfxVVtVXdqqJ8ect9TMM9+PG
RKqVBhcGwZhcha7erN/fzopa7FFnDc2fVYiwsLnrf4UZx/XBGNKo9dTqielAlYyL4RBOiuGemm2h
wGAcDUbCs/bYH9aGzzII980Pn1nLiijsEOTlvU/FWye+9Xz8Vw+Lg9vubpitlMb/g1+R+imH8C57
bVNmzlZS0S6MQk1zNDKOT7KtJwX7F3lPhVvePkwIDhJrZNYY+zV7qgQqhHba9UKQpoWDG9ePEYLn
bu1ukM/LDX5q8IYEkVMk5zOj63TjwvV1uCUMwVghJa8cW/pMK5VXLYtfhBYcb2fUqzGowOftsC+r
4pXMYUXip8yvoPZ17+MJ5cc9lEkjsiPOArRBG1TJ7CnchhoLYG2Y+zUe4nk/vcFr6ZFLRCOUrBsK
DN50sm34ThQpMTZZ2U4yqP5ZM7BdNTK6lE0VlEFmIjK0BNxt38ZIv+SB+YpSuC+knyxqg9Ncs04y
WlMhFSVQrxbkuwMBJx//nFZMUJmuaokKobctsjhVDeZT0gnFrAaJj6s4tS6Nlao5H2awEZD8rn2h
LH7HRnCGEpGuRxQK//Iwrz+XO1/M2/uKggElCbP5X13lyNuFzAZax+xUMf8q601vDw7w/1PIcpfb
0Le96h8k8kUEwCuyvCaLx5LUWlmmJFAoPJiUwozuVxOJ2TRYdpmBwdOIrn7I/54M6YtF1KYEbOcp
KZGzsp1tSl316QQDwbRAueYPycI6zanuLAUszPSpB98AGrV0Q96YvyyUeqbpdvEb8uPGHzhbg50g
WykwAEYcq4CMt79JKsSe1Lh6wG8yt9OdRXTg100IQk370aoP3yePuI8qfIkKqGFTYhpMYP78oy5X
u4LQ9Qlo8ijb2CH3Dh05INugdSEm8vtM/5+/L/yaycnMsmulrlM9Hdq2lVkkMccba0hfCrSmt0aL
PS7XG38ncmGUFGhNJd7VWDQCoFRTkyBfdraoyWPhQ3MJp7/mzhhrG+jcKozfcvuIJmjvtopoQarY
ebiz3dd0MUS0HkBWhT68hcvHFgh3RfsuPlaF46aGhQf5RsDEmUCSvg7oxB6J6v7Nm6vkLbXPoLMD
oWwLu4gu4iIANRcwGcp1NT3Sg/ktmAROUQ1ftpEwF1HdXq3bmKSw+9+b8B2WLZ35Ez5jpj9uFKkM
EeCjpJ3RFSJamzNvCyRmf/0v3lRX2oRH4jTWtGVKDWLiEDvsFuifO7dmCZXbJNFnmApfw4kcrHe0
UQa9IqDcL83t6htkUvo5BHS6RrebUhFbUXQeooICcE6ubHMPDFzPLZD189ZbHBJiuXNJErOuXm9e
KrteHVbuerbAP5E12AFyjNy9ZkRV8gu90xvxtUnj9JzjyTG7BDubxdMNohukqR3LxRxfa8jfVd1P
l+0s99EPdW+AegeY9D58zBpOrZkpXab6ewNpeJGQ4h5NUjb1CIbhXnTtwy7WkPxxNWVOY64hcuGo
4cv90OFVOMjGekk6PnGPq3Tr9CBvaiwJejfWN7AWykrWRbLyYrlTNXcstkqBi15lNA4ifsz9UDLt
/zWwHwI/+LmFZMDtWM7PcSV3h6iqniEs1MvxghiJVrTI1H3Uo+qR8TEMISDshDKqIlanSWe25Fde
CApn5vMsMbWllffHoeneIERgi7GYKPzsfTU4LhPvUp6dYkCWS+blJcHOaCi6Zz1q3tBJId842bjt
tBVIauF1FzSCAeyzx+lSmXt7o368OSN3aYDBRrDyMThqRglvMRS5q+a2d4/uZcv46zneM1qxI6xh
bpNVc/YtvpaD9QoLP/f+26RCDNR2s3Q7q/Qz4agCum4T+d62jOOH0RswzTDqVNR/GNgD6ZGqivUI
2xXBmeijmy6u+QHayRGMjrO9yYDEigk2Ts23qMweSOUWRhH64vrkBEDXEu8tnIzAHR2hH52fd4XN
Q26wJ4JD9LrfE4wMiJbJ7XYu+o1l+4NH0cQjYSaCDuxJPq6uJl4r1zVAWpVSgZt9Vu3Hwuc7Y0E2
6DHTUGSWfseASyoX93+sQNFdAAAvCOdd9XLtUJIxuoXq8ZeVUh+eH+KS9Mz0nT2UCHEafEvYQpdR
6cAgWRua4PO3/vNQcCnuJz2IUjZOC4jdtazqO7R16eEiOuA8n83e6fOdDzMbjXNwvizTi/zBtb1H
vmlp/x4YaE/8TtNkIRpllQnJRahdHMi1OEJNfowDZ6XbIOuxenoXbj+2TzfovxJWh7pBmcN1OJW/
XzBib2DDek4tXSDNv2LJzs9ueqnZ1nvoQnnHtWbEgsy9lVw+nqTaGMR28IvDdBjXB9S2W6JgzGrP
fF4CeellAC1BYUEKjVqE7GEFBYTboYZDFTPttKaOu7VoCEVHjOFA/US62ghhBcN9hrndZZiA+D5M
uNi4z5nz+JsSJlibokfPe93Mqm+1rgxkfbVDOGv2cDdQk8fVkg3any6gvDwXdGAWyuHZpGWSCzub
hkVPqjupuLtn2LTaKdU/W8n1PysydyuMGy+2nrmK9FFOeSVZPA+bqVAqj0B07QHZd/3m55geQCK5
KZJPPRRFOyMDBnlpzCcYxNFfuWY8oEKYyJ6GuMDPeqSXeDQwTKHnbbRvqc7m/IA5MeJozKFBIQLR
bdhTHecZy6O1cFqk1AbMUzUkPYZL1h5wV8JC+3XZO6zLaamnydhMEvX0ZuNoSmFh0zWzhA1Vlqba
F9mU+qOz8R5RtNsFuo4zyYytwVeGtBnsS7ZrLnv9yoKnhut9sVjEFo/fJDA1qEsNys2WdANC5JzE
3O341wnMLLgKmR51jRKci8ZzIWFHRgwvcchyPE1rXb33JARXe/cxCEm9q4TjnAPf2i8zWGttlA/5
nS4XSvoPfDJjyLuTodW32/TkAevv/oM58Kn+8FCYaqdQaH4tUpFEEljp4tTNFj0n2uAXDekUPrlU
vRyxxKjnBEegahjBeWfVLxI8Bc0p3/dAjQuxMnRHQGIP0jv5dOR1bTflK1qcbAET1pHNHjNzgWTi
Y2jhbvmnGwAl0E6+52ei3djvBLQljj2A1XOuKftJNba54JzBwTtHh5CQLk5uty0h6MWQDDwQgz6V
ECVFGcdw5ZT8gCyE4s/l3/77w4IQ5rVQA1nIDKTUoJ242N40z+54j9Hpuzp125sG9GInqNjC2sUg
nFSEGJtNhk17FYZ11fAzzMIBVdniV4uGXKeEcI5EeItN1QTPK72LSIczsBAy7/5tR7gfDr1up3Cy
xevmrAzmeKsEVRlZZhfwN02F617/hKJjRDWlZTCusOeWFv43JdWu/oW+9ZkHPWx4x/NtE2bz+nxs
E5v79Gv/KaixRlpejGbkNiDqIa2YNJP6cadlHU8Yd5QoSRzYxqZaiGOpTtdm6UUXsEAlceAUwxHi
P+qNRYBB9+Uh5hyaFA8dmMbz1vxnfc0XeMLso62ZqwrPrOH3mmgSceyUzZddX7dVhe7WtugBPuRN
kMTelAXXvm7CjSon0+c57EOqexuzaNccpyPfMkgiRpVvN6Tc54uJBiFvq9XbA80N0tHM0XRRVZ4b
URFc0UtY+ok+wUbYInDHcHP6ZH8opElWkf/hskW41LaJmeClZayMdJEFQV8K7JbqNhh0toF/J5xh
4NOcWwKffWH72unblD0tKuD47rBI/dUykEsuOO627jTweS4ISmSJlzxYNo61FnlROQepLtzSuEFu
TgR6fKAd3BeXdLOZMyLwqCTngJ6G4VLRr+kb7w6wG/PWMIVG022Ee2ujgF3Djw/CH0t1ZVBNDGva
3t/32af7JtZPwUGF0BrVGlQW922SKLL9MtLTZf9GCnr7kECKB7s5eU9482qJnTo72J+J6frTKC6d
Djw6VGJCsiBM+NB7il2mSULBH6Aj7ysJQbdmLrcydyqREHIsIuP5yAGHQmthtN7i2gE+9hZ0BFqp
+AHmgmsdZ5YHeyqzT9dXhR2QKB6Zv7nk/zHMQlRJuhFPq+UbxgMcdGXI7i0np1y5FyAh5NpVS6JA
8SHAXIS1cEbEQNi+N4Ben1u6OorPdnbkc2tvkWHuNgiNzJZhTC3a045Gem63qWm938+mNE/AO8Nu
98mpPl1WxOjC201v1W8H84nAk7cQHOsOE2uiplPzCW5aXEYN6Gh54iXlMDkiCnBSbVqpC2n//qdS
D8fPwgEo/eh0C2CUx7uWnzPzmU6lntb5F1Qj84BeNx+K0wF5ggbu/qKv1zwru0axYpbcUZRf2FsW
rMtG2vaLDabELm2UxjO4pRF/yViokmvja4mZR87VKuu/zCUrLyGNJccYx31TmFxmNQ7ojSlCsU99
g/Ghg8bPhcHTvuXYj6LuQCye8rEVT45yVvx6jSPMI6UbWml4Ou5xKdplOQ7iSQ2EpEzjqp2j3mGq
px0WynWifhCHJsMglmriPtclJZPTtXVpXY8M5046bk5RlZhk/hcSC0zS5Nb4tcC2G056dOa8E3vj
O6FFaW1b09qBI9vwtgX2/yf0mrY2jgYPj6udstDHKPW3IFGq8vIr+kjf0UCtXpRFXJVPqmYSOqyh
SdIh3H/aFQg91CGIvV1vzOQ+EdOeiQ1s+UWq5FvgjR85uQrwGZx3g71xWbL8yCOu1yAEFx+8UCCo
Ha4t0cZ7g+0ztwmpjes1Is2Sg9b5C3F7XWhi0F0eln3BzfezhkAJOG1Lnha8/vtY9R0CBU/SAFkU
YL0y+BipnpmJhSFX/Jx5e/2RvY7DL93xa6cvOiI3I58Bj4ApgEZbbMkKB+F86BLdm+dC/AYEIa+C
PcnWGL5D1BIpGADVjfIhzis6Egv7XQ6mPGkwj0KoPNsOerXN5vLRN6NyUA9RsXGNboEOxb15xDnS
U1OgdwiX8tyRfOLTuUwrcAo0NUl5xDCS/kFb/7kPGxCKvCIR1BaITOJAcd4kKMM35NItsKX0BQZU
p2uRh7xpydfcrfSG7qF6WNSYl7+cGSKM8yGo1BRvr3FsbnfvIm0hyXJTLcaYeoRYzyf0PkFApzH7
T2u6dB1aQkhXI9s5/tJ8HSPHGKHR4wDNpcLx/E3Lgzz1cGP3m2zfog9R4Cone5Fh/dmNoGiPpFlI
xprk6U0CtZYx7jYKInPHMgQhzQl2GCXVk7nVwoHm2EEtgX7k/d6c3STQ+Dyrx35Rd8AOAPRDTysC
I1STH/6Ed1CResSe6CtFdifFf5yZjPOyiNlKSDbrTwCxrE+msFWcLcr7M8EDw20jhA7bpFgYdRIF
1bP8BMDtDJppSP64BOjHU9l0h35VM7OPam0CJb75dejy8ZAlGDckzwmjVIUqpIh/Byhvw8MnVQIW
qUV3kpZEGhMCJ8Zf3GaAKuXh/4OlqMyXEeykFSh64kwgcbgUSX9HD5Pt7Up4IwDyQbv96kWUISUu
KZ1o88560ZAUQ+p1H8Cb94ASJcNzrEYTOLmdQHAbLuLCvJkJQzZjL+KXKNwNRWdcHhupTf7YnDG9
KIVVhdl6QBjqNClizfL+lxbovh2/1LgsjteW9UbIt6MJiAtWZ92ijy6Cm9WH5lfHwO2adXfG37Ek
gIRBHukZzaPLWk6yEwNZHFdv7TaO6gUxjn0VcxgRi83kWU6Pb8+lYaJNFNx+HoRJ7xa8NlvUVdHr
xk4/I/sHkKMiAei/2N/K5phVUH5P20MY2Nx55NgFxf9mcG0AzDTvK3ECrBvf4tn0bAtTM7I62ugV
3f5LrWs/grgVuDHxGUX5PKbBwpUB822jtxUj8oDwcTtZPR+UWLwNgFb1bZkbIrwJi4RuaIfGKuSK
G33JTuzJt0jJ/5wV7BnsGXEgWwCnU2ytzUU2E1LF4npzz9iksX2phJmfH6DClJrUWG1eCiEeMoMc
hEhhW4I5ndNbwBIWPw9wAFbu4vEH1LnXwLWsVCHmAZd/IaLDFnQfnGXbX1IBJNxx0t4rzi4gHa67
aUitqlPS3wF/ChsOyCJCIA==
`protect end_protected
