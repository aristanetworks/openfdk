--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
f9ldgtJrURHtBvlMakRySvoV/MpTA2DvDy5NarA6z2uxWnreGOfTLXchVKeSY5RbtxQhLB9vV6/H
mtMcHZbcby6wBZiCTe0Zd8w8+P+yemssPnluszXjwtNLkTuH1cUv38sdy4F6RzZ7n9L8Tu0w3epP
ARPBsHhJi4U435x13A21EJymGXxdbQeBqVvgXfWYir0QLr1rzAuluUNwx9ziyxuGE+1sp4kpzoO1
AwXDmBQ7bwRxogBJGFbQhEqg9Lh+N9LZrwOOtVVnNRUshG5egIEEIAbXB8JAPo4OEd2aZrxv89sL
k42owbxU33ohKxnYgWLZqXKReRpr+153+9Jgyg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="MniEttaNvMxMXYOqHQMgfPWWJ1WrSyeykmG381/WYmA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
UpADyk9o7wAQhO0ZivcpDvjO/HkLfkCSzC642l8CDUCogHWWulf7aif1hHeRwUE/tFONONPtN9p0
GA0WOtCbgErk9oPwnIaUk5g0Kj1u24stP3NizN5h8Jgb9UJAndXiii1SjBn9fsdZzEVwOkY48VD4
xU5gJmvClQJG7vJlFcXO+wkiHYCFzu9Fe6wp3eSFScs6HXnfnZ8uE0u2Q320alzkjUXIVPwiDuW1
uqeEXuvBT3hpbzEzEcZI6BYX9xW3NbP3lrebRt+JE9g0Mk6IsLyKRQaBFs/Inor4W+psx+wAGqIh
X7HrrnIX+pPrLaxm4zC7jCWBivzxEvcX6Cuy9g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Y9ucQ8IE+FkDZddEfyyoHvhkt+Qrn/C9uDgLsPjFSlU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12336)
`protect data_block
Zm1augp9qD9mxajYgQyDGVLBx7Krv/SgFVk1XYBINhJDK6//LO5K4ZoJfp0TWWNan5pi351m9Q7u
z+8z7bAiaGqjPCV7m6o1kwStZWaChOTCkX5zQO5qV28lkgmY0cx3A6/4eLzc8V8PlXJweznGKQ++
KJuSysRlaqggcbN1rX20gs+e3yy1qMHwEezKy8HupyF8wEZoHjZimN8MIO7GiTjr5r4nN6rfH0se
sN/Ubn35UgVd6hfairEpV1q/I2hEeVcSueNkrLlJQEyv94Ie7K4zkh1gzDdfoa/JT75KYPYYZEoS
2s7KEkpLKa4YO7gdgfZvvM+RQD43o7lMfgqnrd1BxXnpDpXoC2pvMy1jvGnv85/8X7zET6M60T5k
/LnAQBw5R2pLO9pkgnDXSEDVQfBe+3MY5PAFNi+qiueTH/ZCe9YoPyT+7+Hp8HXXPB15K6YlvlKS
EhjD4I13p12uXXBy1QlQNxkVcLKxacnkZex0SPlyFJnBQ8U+SnpNJyytUpe1AdT3TcmxbatoxXB6
sDdgutODPTAqL6tQrBZDo73xS7FTvhQt5iwmCXjZGXW1mMgMMP5F0wCXd5URMEztzz7ZfIPpu75h
0Lk8KpRrp7+PPV5JUacEavQFfpF7UsCa9yYAETDKjbb7eWukOLkgDuxgysuHz2Yz2LNCvpuHRsTv
Vza/h9XxVbcXDmN0rVv5pb96KtfYZbRm3pSAAeXKkFWAspBfe+Q/4nphLL8Say65urROlfoXNb8G
XYt2K3QcqwaQoXAyqeErrXVK3tr6OHup53OUyAyqTK0MvvRvXUdx8OAZiPVfF6kZ2KyXcN3/NJKI
RMbPmOGqmIn1A2dcr8Gq/80PKBtAQH30NDOvkVx3buAlhXttdKjAB7yXwx7ovc5xaqbJKTU5tXHw
OfOLRAivIPmjo/aJ0fS9mUUtP3zmjlRtqa3KwTKGrFv6Bb1rafuh9NhvvYQzmqOVoMk88vvGdimx
TsJmKU1iiGcQfoMq6UN59yFjGKNhHj13aTIeJUmGZ75+fOuPuC8/NVm4oq55Do0Q437PKex8JX/1
zAcLZR1S7AxpNCDJtM6U7dyu1BttkpWpO6Q9+/q5L+eDlZiE//6fAEficSP4In+2rg35gO6brGAq
T65yUYjWPYqBu5VUIaUeG9BBwe3RrEAUaLt8blAy1sH73ArwkHf1Sd1baHFB6PQpO4jXP+9l50Wx
ogxDCb+Os2eK5qAnPxoCZ8M+unYMq3DV+E3aNo9HnWkWhwqu8nn9PkWY6vtkgrRCpVBEmfeRNuG1
rklMjjlti6cg1P5h1XdxMyLIjZLEAXr7yVy0moV0NTYBKI73zj9hSdNeWbJkCRSPifxOsxzBrG+m
7Ce8vWY7f/uyedJBspjQ2GCAgL+fsz8VZ+NrYe5kDspaNqYIMSfvkbYBeydSlkmsApzYG6ddBm+o
4Teo759iJ0YzMA78XLVpz4jViilpIdDE9/il+Hi+s1sxnn+PvVW4/LoInJJWGdvERMCUywFF5hPE
Tx6UB3TiU8OQV6/lccn0tdyEDMtIbIy4EXrYXcsWoNDNWs1PeYNpsVYiC62ml5tDlMyohhgzKXuZ
Adur6AEURxK7+U1obm+UGUrYKBJSewtvjH9BXBo40TAOAYymyGHQtlvYZIR+W/OrgoK7h1SBrGkF
bci6TZmx3kyYc+mLCDI0VcFvtQIi+lq6N6bFvr4P+bM73mJNDqzx2GMBlPTCtF2d/Cev2fyaOF/E
kRPUXRtBXqAwuWQyZE8Wqnk3D5c0UbU1VLrW/FOI0Y84JtIkZwlFfkZkpXo323sDQgE7cUagmWSL
GPyZA2qYWu1MeyXZ2JIvetErSfHQQjSH7VQgCAoPrOx/cMKzGxoWTHTajnztSE2dwCIoe3SBaE+T
22Mc67TZxP8qIPmS6rynyvZDG3vlX4ft9oAqcJ+/sINIArQ0FSOW4hlYbbHX4J36Yk6Oka+kPGFp
ruOEUiGIyqKhadoJYEy5VjjC4MGGNAMHuu/iXd6I+Dw1lYXC0ffj/moFI0FOQZxv9w2BKh2ypO0C
f56u5wca2pbflwtakb8ms5pEDmAP2ZugQeOVrQBKosVHOgIy9blniH6NLV2Dia10S9Apv3mqny1i
Vdd9LSlID/KMYKmHAoYOQFstLwoZlSdIScQzIzcPc8CuxVS/5WIkaSLZbwuHehLFJb4O5HrOI5Ao
Q0v7pkAqsXvzH0sIEIzvYzSnjFA00oQK7HkkSsNzwvd8SmyEqTC0BhAu2qpQtl+bciJBe0ra8NM/
nBnjeiRdJpCohG/+EsIXDzvqCB/w40DqoJ8ng2ULYxPPjgaORhmjE+tag48U+/DIlIfZFhyd/vA0
cyYP0vl8mhhH8yidOCorduEYXlesycwGrZl7sGcuBsIDnNodKu5NQCyKgxb9k6y6cQf8OpIdkEhm
rkTyEjVkzaDnGCVFyDH1+J0MU91S0omHQMowMFB7iv7DP9joxJle9gKx/EjxUPGD2fnvu0LItlT/
jSWdSrXFQFqNhiIewoU6toGlm38VQPE0RX0nW2gB76Adi6oD4enm8d0DhgRtpi4HYbfiKGLweIu7
kSqxycwRQqjoxNelfC3bPbkOHtOJlHpfZwpzDM+eXHyVB4078hPvsAA6gNywqOOGNf7IXvwpU3gF
sY48UsqBRdUVAA6eZteYKQ8Zsr3Av277+sghWiBrZmprg9khLLZR5U5ji1FzOF1UL6jInQ1zz6i0
9vyg9cOqiZ08jqTCmrDidJu56bdrKqWv0YyyjY7jnf/cS7Cv/y4ziNshSQUUO5+KTjogtODRklsh
g7j7cDnodTv9S3oPpACNjGASkljcCXhKomLB95lh4PT5m6inp9yzZtmGIk4+zMCM/MwtEQHdjHPl
sTqeEmGJFsqB0Wg5M0kEW6IkxstSRzHPsqhVeIupAaipnc2oQngnS7I5hhXoVS9Qpqfqps8gbW2f
41qQq4TcRtUDkU5KqBL9xahsJnn/nnrf1FsJ9Q+Nf2s7HbykegdHQrRPfazmoC/Thd5q9fR2zbFP
83XForswvMy6BDv+wFwvmFt/ENDchHH09EoBKcM28xPQFX5rjaG/eGbqDcZxDe0NIyO7bZGPCnBq
hnWm3zQGDNfSlTTKkMuQRwMyitatuR3cSMw8B0hi8dBChmbv1hQWEr8sQ6/lHK75zeAHetoEypqw
hnBxmL7dKQCDbbiBdyKTBmquVQg+cqEUntACS1kT/mnt/sEuByDSkxt+nfsaDAnFnNcqcGrHtVyt
iUWDpTtYo7QyjQ1K65014JCgGM86prm5jVuLXQ3RekJuSZyq6ciuuZIo5fcYDh9GtGUWNMkF4MAx
tRp8ViXqSKXLlwiUP51N2FN4dzUB5fHMhSOnzn3kDw64weo/+tQFLEHBmSMyFuhdc3155JaFy2Yl
dFUwXZDtkvhfe+Ti0ryO4jr+XUTzo5COlYjpx9g9R4wkbuhC7sKkwU1WBgnsvaSmyLVOW67Rs7V7
AbcJMbb5pu7E4nSgKs0lFdHEZjHU0gUzblajOFp5tTixDc6md4+oVw1i5U2HQunq+y2WyiTECHuy
dLOKpIh5QkLqRMqzsZb4oXd1mS/wRXFFHi++BVIHfNwa6pbz927dMTmKxINfkPGRekBpjPd/wYuo
H3UnDz62ZGE8rbrIKwh/04T/ktgK5U7veMyof1tJzAsz9sfrBEZSn0woNaCfAeSA5zfv+T+4gKEb
rc+DX+CE7JU6G1lgaoLSl/LPYhA/p08qSZM7Nl+jAe8+B0icxUuPyijcjxw+Fn1VWbmTIPpHmcZh
ue0aYukRRLU0+EuMcI/wbZSr8SXnMlBjDmVYQuQgFHyPkSKmbPQFzeRcglrhTr7a25267lc0oKgr
rYTtvP+NStTxvuSWWAS5RKquRy5LdfvF9X39c0d5HlONQAzRAIdOgxtG38d6jVEYjMERiJgqe4JT
qK1lVTNWd0kR0YNiPeJNlYNuWrRlij+7M+gZ4bldXvVVUHcdgSz5FxFsmqmomUClU1rsvFm8RuQW
53JYFF5TAC5HoyAxCNjfvCYXnoIGzsBaLiR2zDUBwpguq7lB2hLnjJTovdkRtDIR4EUTfkZz8S+w
Oz9dcOWXT8c8Q/7f3jyzI8OP+WNbvz+CCOnJJZxW949jE6nuwluvlqVURnoHwjmWUqpTyULQ3qQ1
5qjCfUEs3mBd36Z5Dtw/5dxoZFjWhTs2yjCymK4taoB50RBjdFtAhBEWIvdNQtRlCvOiPv9Gvywg
aW0PHuD476fH9Ylm+kWp19DDKe6o8tRQwDeB+RXOfEFUlCxskUc8lA45pEyMcj7t6bCZHhjt23IC
12ZYfwn+s3MIPrrXmLANi7x1IrIXqtpaVHoPtQkG6kjEzMZbJ3RLNVHeCmOh4co+jYsbe1aq30IX
+kuQA/8UXHVXFO6+53YUwJVXWkmpFG5VUZJQgvewgptDw22JS8TzGw4AQWMsYwyZIx4A7wk7HdDC
DhCpzBX3PVgXo44MOUe7BoFhOZSXsuqgomfrJWlbSla1K35uAYy77zuHNtvbnDc6MKfLKKdxXQOX
OnBWZKQfItH2b4XEVe2MarRCIkmB/la5J7AeCIvvFc0yAQP9/giR/o5MGxA+qfk3Vf9Y57IFYJwE
JXD0ZJBeJ7SYHpcAZ3h6ppHf2nIHbkB5GuJL9VxlRqfcspwNeO/L3R3vyW8yufwi1/EXWwydUNGt
bMuGQ6cU3e9UjboxuyNwXF6duUkATI/nkTQLAzV/485DewbjfBWNTavwmTjzghZCcs5LvxNpfFhI
+p5K4viWdjs/8ZOS8a9hlfD+uLCfxweR1Fgp61hN2w/Ut0wSxv8GUXYxcnuIcEjq1t6MmsvB79Os
0J2aYi2gAtTkEsYrRAKttdIw5nZvrINO03jZYn3SJI5tEwk/e1HwDiq4r1YIxenJ3ItgGZrbKALa
F7eEePLujssPV0JvDx3CMhjR5lJOVHHpVtSFcmoN3kFehVqWagLD6knMtUtrlPciA0j0TXGHpjiN
aUtJ+yYF6G1Soxgl2bYk6KqWtOjlB/dXGKet9cBBeDWRAdpgCITQO+Gptxs92Uz6h4tpVl2YsdB6
h3A5VtxPyhk2g1BXWPSUG5c92lVpNB6SFWWA+ybfDLxaFLGj7hljszyb6a8HBf+ozoS4bvEaMzzj
n++wu0LWb56gi+b5e8Xum9j86XsxohVLkTcsXd25EHlvWN0TDyevdsZVq6vSTPQYiuvZ4oJmcx6W
f9KX9H4ONzr7uuG7E+55MXzZh8CDGuQM1MVZ8DA98HYu5tPxhgMmz0l+SPsQZAIhpxnJy4bY8lDJ
Ru8/R0cpzo3HGOy9tePpLPEzgjvXBpWHjoxPpnxUTCbA1Lpq9OlTfYbBubjl+boOFJ8VR/PVwqTL
oNXbJAuB/pi82I7tME9Ha4j3UqHnTDm90NPY7xNviXhLREHaMRmz+g5vrmRnsNqD8ZX5Z8PgqsOW
ar3Tv4rjhP3yxgHDcVcNuGIPzHEBZu60zPiNQIbwXziriXhqECHOXTTpXFTuQM2DiDLU94G4HH/W
10N31Fl3mGkt+00e6d3bKCl2beGIhkUN1++mokELWzw2JaLad3nmpRJEtsK3nZKmxJFyFTHBbWR+
IRTjuTAhOt0xIUMXe45+bc79UdZNbi42/ExTJUB4DaufSh4skHx59srwLhBzqnqMQfiZUHkaUNQP
XhduxN6e1PcSVG40yZCxxIuVLPoAlRUorqbM682LtT8l1GrZlGWptrh9qhQsdGBvECHPMjQptvqY
FRuHPA6VXZasufTL1G7eeU2mL0v8fD1+GMNW5wKcKWORLLo/CPA0v7/9OzoHeCX61BXJQvLPVjeG
Vp1CioJmaA3x/a36Y78AUvUWEhATIgBF6tMuPBBfBqqpOgkcJNFApxs/AEknpqwdF960BT5Qjb+6
zDnV8ikG9j3NFYM04NsbaB4vvL9pShATWoTLw3HKEvfVme0houKZoC52Z4BPG//6EY8BaAZNPSku
1EdeRiFosbqvg3uDuKnLzun37VyRBQf8y9HxeRnRiMK1FTTBfkmO5aadyboPosgwi/YgmquAA0it
zkAZhxHaqAHxfw/3RH9UgpzDp55rl44YrJaMlrZsSL6MBkISNDJWphp7eM8Eta9H88ecLA7WJhqo
y5oKASTSoZiB9P5oHu1DSYy9z0Znex/1VAIFOq//DVCaUG4KyTyABTPsstHhjVkDheAsDGRpmBwA
B1ueZcC6E8CWbGS+d22UH/IDKW1M38Mn1lTuhgO4JnjcvNkLdOlNcdLrvrTXjjfveFp2L2J9L7hC
ZhH4tgfPb0V4LeaJgEKFadVvs5ddCpv5RjcnxW0EeeevPbIMWr0vMIrPqrcP/Iztg1A6qde5Ajal
Yp2ADp6nPmBhFIYkU4g/s/lDetLp8gWsQytRJIs6VOBUDnbUIcVcQj43PnQcFvdXQMc1e+u86KTu
lilQR4YFPzXJn6RUy3GoCb2NLX7dUNgS3TlgYlAEjAFpPb9/w0izq2/6ijcgyHvwuBZ/I/aUQF4B
t94rw8W4s20UeOn0/uRKzQZUm6OQV2xnAnsBifxejZDgGv03Ihy20XYXdreCrjJPQ/EadCVLnBtz
RWEqc6w3YqYq5cAz4wRutnirEOwnPlSTQuGKIdSBhupd2VvZvdr1aGTPNOsxSiFXm3Cil+JsDIlM
MntJ+d4WFRZAdaDnDBmintYrtJe0HnwhIzhSiz54nb3Lm5axyGgteFPB+hf0nDIzpET1dwA0KazU
78b96WuB9+CDUtOD5oODW3Jn9qFh/JUQ5ibSbdGLNuDl3KxsxYiGp3I2oanyjW4pNPuYJ79adRfq
lPvTUqFmbOaVo0Cwo0an36nBSTQ56jhtmY/Xq+Q98N3SvHlA+cJNV/Oe7KlsLoGyWUYoTfmJzLgr
9ie5H+IpkNbEFaSmJUxUtVOVHR5jx28QiHWZvQERIy63bnyHutBZl8sSqAv+2EPxqwwINi/y5edf
SwUQG7SXKBbJUdTMZNXbLiUVGP8QCn/7KeWv1V4DIsATEH0Dg9I7FqdntoWGP8Y3bNETnEj0rKk7
wmKyWzCYcgPogxtCCmaqIOdl3JAJWFT8bz6eE3sZZ4rKYkx2Xi/vp/LDKzYopG1Smcf3hGZ7ghzf
yXq/uXA51tbu1N4vJA7Bp8TucnJ0sEcDCnu9KOj3Phan5e0YhC/Gyknnc+BOwOpSp70nCU3M7xaY
xUeA9ruRovpMhiW8cFCW3vrfZzs9slOWqDqQmhSeF6lsubBCeDFwIUSxS46mjYG4pR+Wa6sVm+dh
RJPwXNZaCmi/i8cHGPnlkxJN9cOXYuGKAUjovSElCWRZzxk0HzIAF7hwTFdOAFNE0a/WdYqb/iDN
I9/NsyPzZoIJgKGSbnptABTzL5lf7aeRiWWTF8qXg1vh58+BTHvssvZAkkafannPVOPkbHcNsY+x
b3KBnkmSP483iY1m4sVZ2xLM3yZUs8NXwAyOEqa3Gb5bIPjudUQH3xfUw5nDML0wa91fs/eSbFZn
AMwyhAC3kx0A+X5noLiz3N6nH+pa17mwQPZyFD8R4viev1hP0OMlZ7/zIdRKgV4MTcp2CrxQVqLJ
0Wmv2B5Cc1NFXHcL1Bs93j9GMkVnFRYrKQFWLkLdJ/zYZDxUviI8m+g6DpvMrIZ7mh1InQ/W+IUK
ZN57X/jLaiptoMahBI6Ur+wz6fE3XmqyRwwjHLk57+6Gt6W/O7cFJo4nT6WbB+oDk8kfTUl4UIEL
F73dx0IAzseLcRlj41QMw76GSesJ/szMKCYW3F4k4DffGttkCyVmRD0PWnnCCORWwzn2ckh55YXG
oYOihqLZojpvvorBSYPucWhM4RyCvp2IyCeHeotOVoRre/lGpkh4ERTVq10aI9dXOy/hhNlVbko9
nUlD1kVTnNXwJOYaMIbZNRn6aWA6lRGZMIY7dNW7UmNITquQ5uRSER9VYHSGcoXqUeDuu63K5FfZ
nRiyo73DT0Qyx9eCcrG7PTXccScgP9sxIBo2kjrcfpY3Q5HiON26l2gLwkJPxlt8E6lsnSMLuHdk
iGRa+k49pqzt2JYWQUji2nGg9yGuaB0pHB1n8jee86RhDzuySxQm+9iPPYJh7dlBwF6ECWolVCB8
BUtJmrVOK735bHkjpsJtgI1he1gMpb0mySjMU1Brv1thpwtifBprdcvcaL8OgPdLjgz7UTBqlJsh
njA59Om51EkYp369fb6/3raGFj5mAhopBJgYQ8PnDPaI8a8sD4ob7RkvjegwXlnNKKKAWuTHDrUh
LJ2z71LvKO2APcPYv5JMZPllmJM/MVEbVVhWY0fS2frUwkDaFMLnMbnfTvEentwzA/R1AE+dAog5
a89ufFRQgKA4FMmWOLcr3wIkUIT2EQyC6XIG6hxFDfdCEhlQT6uLel0cCSGSAAnagJ9sj7KrxuSt
cyCiDmBmK8yv+VatRTiGFU2io4Xga6ZBIKAvYCl/6uG22xIe7mTcD8FjfkL2f03WuMG3gDNUExJe
2CxRNvncZlNT78z8+rQ1b3gZecGwdIxg8bwEHHPbQ7xdt+W2yP9v5GdWH20P35uSmFy/Nyxl6cEW
sEzyRtiOgUdD8xbeM6EaoiNadFwAYkyQnn1Qtaa3sBhzVTuHKZOaYRs3cQUPQTGVJ0ZPbezVNy91
vGRqwj0kqaXHCelqC9XLvTayXkgpCndNYNXbBw6tMe+BspZpoNIEqCDVlOSFdsT44GnhhP4feks9
1FEmCAClr8N4Gr8Sihubg6h6fCR02v3RKa53XXLGWTontmxmxSrE6/3FpUAvT90Bgjvoi1x4RmI0
m4Ibrj/VXoD1Cd24VRV3uHAGe5Owj0MgRX+JyNQGxeDsNm7+lYucAuRUqhjjpAgCW6aQZlu/6ZGB
KcnoExeWBzPPIFXLqD+43sBRSftJYyDN8q30roQ970hAV5FruCfjnMUw0aqaR4T8zDvaaD/Jnjo/
yImKey8bn+TameXw6t3kShI6w7j4A0QqgZjL4088F2GwMptFvVXL5lIt9pF34/a8qgDxgiNjyNXj
EY++N+aDjl0jRttcuBCKWH0GMzuGVzDpTwP9w2r16hwONDYmRc8SykTsX6//ZwzuiK6zkp3l0y9d
ZQUdf7KmE2uwISfaO/QeiEZUq7dbQBHEuPgdrseHDkrE6XuCWt7XArD9oQUWLGkgToEbsSq86G2b
yD0mpgHQrpu4wkZWkRJ7JwRNpeKVgGREd/8Xsv3r/zg8q9hN5rCGvHkCCBB90q09NmTBIaSdsAD4
HZiWSFF2c6TVwFy6RultuWZphDxDgWnRyKrFoEffCCJeBhQWr061nnimBQMJoL9rkd8AACQpBksq
idYQIqT+iqCn7dV1xshyG/M/tQ4GvM4I2cE2ifGY/VGIeHmY86+ZxnEAj6+vqoFiEVvl+CcUfflZ
Siz+cH5O0pURQgioRYD5AvqT7fP3sztdrScafw/qs5LQegWVS0XYu6kaLlu8+kX5IVkkamrFKflC
kG58uMRkpRUql1DATYMTp7V0l4vtOuLLlxs+tD/11uegR9qovofE/bzxQQa7om+b/Y5YiyQh7BBO
qaFinfFjabnsy4DiB/hFSifUre9IT8UpneM3a1NzMnlqifCoS9mXQPAErV49Kvrmagu4gokU++If
PTZ0h5gw3rrR2ZfeNIYyhQPcJiR4G6kDwSd+kriap84no1nBfVA/wU07lVvx8QZYJXH32Tv+ZhzX
djmdTU0vWvE0QTPWNVTx1G1uHVeNfMPVJxWPtwXuFO22wO3t809J4RfPoqxelnsmJ2LZw+Sh3E8N
l60aMvC9jvihDxDZ1TBjG/t9P9yzmtteY5g1N6C4uIzrYOI+veZwWxOcIl8xRvJ0Qn6Du1C5au/i
NjIJNmIvBI7X98iac3AcA8q7NVIK4anquygtJNHkc+96seFd+V2rb8AeI5uw08dk89AMjozDHQ57
oAsNIJ0LanNjqWDRhh1IJ9rzwifpjecQ2z4k1Zn71HzS0S4FnB6XRup3X5gSMx/eSAn/zTq8W6/5
LsyuqrvcL1Upav6e4oyjNmgzSEKI/0ytPscNFVYSSoYpyc6nLVVY/bZD2Q2JhSwLT6U7VjcwIPkh
Bcj4wy7mKraqUxri3WcRHIKS+8H7tSuExAhCDOFe4HPB8hXzYcB4idxw68AvAxDg+X1KS7W6Sy+9
rVFdfjO4T+UiwFl22VcUnZYGZbfPEhHZaZZzmSx2KkTuGbeAiRRKshvs0nU6SQuKUJbW+99k+nTX
aBVQVveEadC2EjONc6+WlBZdssxtX6+ODp1qGLhwolslU0OVMJ5tUFqp0dvJkT8Bi6heinviAIoq
TkOkkz8o/5h5Zq8A1Ca1IUJW5DL5cRhwgw4Sj2mDjjs+PDaR94lVnjoXmnm5KU1LB5DU1BuK4tMd
GXf6Wx0GguRbP+MKlWr+fv6Do/o5gZvwwHT/mRf2C0iDX4RFWZQVrqGllgOeg57vXp35qPkDE3c6
Z11B+39LH4ZGndargy+5/SlvwTwBFU6Kd2ql5r78TGuWUyYxQIYnQkxlbZismJjEaufzME2yXrv/
da9TlaX0X+XSkpgJwmWptxFi+iaNDs/Q9PJ5425IgbYDX8NGNE0HPRwmg9axbERAHX/6KPm4M5GA
hSnV+IBVgs2KMuF9TdwkzGnWoWSwpZIjS+eoCm2ug3Tt1VrbADzFs/iasjydwCHbOcoV2CGVIcjY
VAY+XIO4SVYmdLzQcq6pWvqHELshSzLjhZYaZsSqLnBflbzo/tjvW83d68V68AybfHL39zdAKawu
zsMkmBhSTczQPF1uykH7dxDo45+syQcltZt/Xx2XlqcxR9jGNOxJ1ntdrvLY/DH18gJl4jMlE+HV
ME+rZkGT748IsYK/RK+5dujzsLZ6oRzSu4ShSPwOaI3q7hsJwNYqU8RDH34plHUapK39bTTl32bJ
OwqRnsJnyEJzcG5YiFzzyrDoXNEGGs63ruWU4gJpOK9lkHk34zYyBnkctQIxcXOq86TWVCw6t6xY
0Mh90HTdgsaDpco67Y1S3aXGgCqx3vNJALDtrPyFwqvtE3QPhT/M9FLTB2zubEAO++qoV+xPgS7Q
jJiJrJbfCLqGbkWa85Pur8PXYzjkwYsp9UZczYRpIwpOCo+dZ24KISNh1wH640pyBEBVe2yNMRJi
WJm+jB0dlPT1XYmQGXhUsAKEUdrbBspoKhwB3dVKXgklLtq8iH4kgZHXdMlaKjjErr+Fdb2BiIoi
I70YwMOx1Q/FsnzkerYxe3uijHG5mEyBNA5QVgIns0EjCfz00choMBqhjEfwzfgw3IkF1uOwb5Dn
3eR9FhLwMEJKu2j6M07jwjV+xVje/WCzRh8jW29ice+URvXsNsw2q7PlTulwJQlAFbSpIij0JubP
y/QgAPiykpLQ8Bx1RgVYKUULfuIYZK1OaqjRJSI9Nr1pSx3YnkIW60A6I7eycWtZPa32xdJSB21i
dTWfrLbGiKkwRSu/u/ZHvBVipWbCtUaYovHvhpGuBT3CNpA3s1inejrccbbM8Qk3gI1sd3DUmhpd
FMZ/UFMA4NzGbtk2cdN2tmJuZ/QrJaPtiR2yFIEWsAeBnMCDZ5gyffeDyNLnsMVmSankEfQ7srbl
bkgu/iSyGcy3S+4m/LcCdPMa5t0DYB4wbuW/JPmp/zgGufYZjsYGc1q7JHMLpvYm2pqKf6wVU6EG
yOYzSq8eRcEILvBZurnmScDvoPiwcXdtM87hrhOwT4p/4WFx+GhL3N48hPrQVd1IPfjQFlHVZqV5
2skWVLvychW11YEFt2xhynfCojduR+LAZ3dbUdXWrHpFf2Cg/xT80vJgVjE1OftmZ/8OMkw72TSj
6azMgNoFWnby3TWdts79+mXYwnE7DFEBvzqmZSL9s5HU7qIso5enfI/K+AcVoCo3kX+NAR6SkI+K
NuGYw1qRD4LmIVDB7R/DWGGcfs98isMALUUQhg8KUOcd6TZGS7hn+Q8kAOlw/6NwPWg2Hj8Xq7Mr
VT7ci71LB4H+aquqfmKU3bpkHogEWucv9fQugT3J73myAl2wSZQLIvAwwRjcWC2qkpUcPiq5lWOo
zc8TmncjW25b40A2KR2/tWQZITbZ85x5CysdIFoeFTy2bwdg4wydz4UxCwHtc4kX3OnsDenBWulz
5KYqO0Q01RuyqqEGFlwQZtIkVDgday6UEZD7yp2BR8VKAHfSKDmLZfp6OwhfNk3lQ6J2TBO+I/Mg
4mCHtpHwW4mcFwy0ijH8ifgFMEmEb7yLoSAp3qM7AxjLneOP6pFcMmEGNQDfeowFyQulfnkImCl9
30K/XJpFt49dn2whwAkO2R1Qv6JeIt4ky0qQ/gts1Lf1PjUsoDqTTDZm8GtGsZ29Vhqp4LJ8Bzls
cLggGbOMeej5hRBwjYddmZcHjpapcaDQynKU5yTWxF0Cy4ISG0u/L8j6aL5ufgzHXq7xwIZSl/N8
Nh2Gfdc32hCvMzVJ8BX07PLRadvZKYgFYk1Sz8LT87czv0J7rjzSZbxKaGupAK41kg0gxiYLLAss
RqBiTSUTHiFPDtKIPKuFC+rr4U9p3o19snFAAX0EYKW1Ce2t8rzAgwhxRE4XKryqFGIOVhPKMspG
AIaglGC70x8lDFry+CqNjfPOXsFGSoQrOh8fSp8oEQSL6kg2Z2+S02c0moSRlu6r3waVcBJ9FG0r
Yfu6ULlvlLjiEF5Yqp0MsQV8F5jzlx5tsZv6Ayo82+n+Uf183+xsuEOn432tDArVf8NcB2+BOpwX
sczymG2NqQO3qMZelEAh4iKWVTIWa1m3kskyDupjv75VsUMwPBK6IdSdHI1d+p0ljW2LKYzMaDjP
5b5KbpfD4M/0JtxS3jqC9gl16+Z1Hk9JASmY+anSX5ed72XPcp9togMzr+jAjJ7J9cPaj9mKXvxQ
GHJGs07QjKg6Mtrf7cJD8iYeiou37X8ZZRgh8wSB0RynvNJsd/0nBeMO3dEmQ3iFnEopULRmC8OA
5G086AN45aAULIZ7yoye4y/P3B6q1WbovV3hbEsDOwCHc4UCYyXaMFO1d85VUdqBzgsJBblZwwgp
laTwEFUhHgDPWOdPOeNpwNBpfAYvXUSJOnYZzcO+QPyGMGBn5Ah2ZhDNvw7UM4k6AC2dM7cjl3Lb
9HZBaRSHi1UWH9upqAXFQa8x6+LqIpSEfPf7l3Bdn1cNxvHhVuLaaELZFqtd9Qlsck2LUDgDGFbC
uZhB7Ud1K17XBepwOCVg1p8CQEVSHMQos7juvGa4ACcWXsLa0kkBzKC9v6+g/ZRKlBZbFuNyQVd0
9KhXqTSkGFxP0w03WRUHgrNvo0IggCQjS/WlETHuNfYA1fCaYgavCO1Azzj8ZjXSfgCh/LjpeyeK
Ibil1BN86QFeBIyvcqpcLmzD6wIWnSsU9DHAejBhNBe9UDJzpZDsWdgi4GUfNtKG7uI2NKl6loXD
xKTOk2dZqAhu9CJ/Nkx5FtYBa5IgI2km3T8e1LkfLVLSLarbDBoC3FRuP1ifsWyjuktO8XgWMFrq
1q0bu1luAr4X+CE5A3H/7gfIf0h+W7v/f2LUTVoZJIEEnPlIR5h70TlLqCFXzri68bPj9TTBP9L9
0yTkd+Lw2sIz9vMsmw/mczkjpvlBfEgSOMmQDDIzNR+JznP7b+OmrCPdVErtlkGtyg5nCW+53GqA
L/zdhnuzG4s5hWXSXtoVpc7eGpLzUWe2aIo/R1cCNg5notIMRSTuZRpZmIZDvT0FW0td0D/g4LrM
A40FfiC8CWNyXBhvcASNSRXBIogXHD/c2C0sjSYjanc1o0Upf1B5oc6QLeQt/q4vr2mHWGX2EkS5
OK5nppVv5fc+4yqpXgNeDc/hVzBgONGNGv3klSNhWNn+9rg/zKBhdgxc5dhimtkxZYgHbzbg8hFU
2d/uAkA3Rbs0jYQpgQS4/5qBC+oNfexxrWR81+Z3Mve+f6m5/9NcF52bR6c3wL44i/lryqrg/bRZ
b7C1xiiGgpuCGDgNmihL9EUS06bfkjIZzmC3yRTKzGg6no8hRU/5BrsnZD5X5v6mnzx7LClMG3yj
FmBGNFH5OExxoJvYZXeeVW2DHXUR+1a7zIFEjHdE5EGkYJU146cKQqc8urlJeFQ5n87zd6xML2WC
1b0wplxdnRHriTn7TQuZKQBtsgNedgZBOIY50PRU6W7t2MVARtl4C/jPhD7qEgz3nr4QkGsWII8I
sLXI+x+H2Su8WeqF1KFb23RP+RkgDxVBgVjLIjPIa1AgCGJgAkhzIGeYGKPtlVM5CkvbmTNpiC0F
cMNy+AXPYv9oTWb74RoUaAjlrosbkObwSQPj8p7MsnDinaSpdyGQSPrBH0MmULDNJ6cCfYuOl9vd
otkWqh+rSbi7baTT21v3vinkCCn+7XRqxSfXrgt/vYQwHFcnNjHvYGpVjtOa6u2OmCKv3nJat18j
/v+pM345WqTearZ+A7rS9jCzSNoAwbCL8O6W7L6nll/aYvaIZYddKStn/RtUNMqW2ggdZ2CRXYDd
WcZ7T9vnVTCxFpCv/2AKlX63i18F7LmS+pb5tgdY3rDw7ieN+fP6du6YWhW1hk95eNLJZuHctYbJ
JZ+VybbUNH4vw8oP6b3a6kEPfgSbvcZJHZ1+H0wSx1lAY2kDpkZLoDEI8H3QaybDnGrdivjw9uWu
LlI2fqas++ivsAVeqErNCeJUSRZ4FKJ+/ndKz6SWorPA6T5GXJd7rxkjYiE0LoqWV4pflTloVaEW
E6mkzkyYnDA8E97ykpxNd+sOIg9uspF5np06YvWlTBeKCWIMipQA+BAem9rFgYYEVHA+QjEp+Y7u
qIpUAE5whFjFk/w01SJXMMlcY4C0KF4KTEloO59XzoXV6aXzeTSYWRP9K7ELacLWa467WQALwdea
B7e3Yc8zm8qJ5KLSo2iMfBNi7RKja1oUju2nEbMXNHfe+Nf3N+3pdIBeBwQ4Hn6R3+V6MLf+gX4J
GvuqdiyvZ0/K35BwDTaQymZgeFVPmGcNnVPIFVBEXY6UZmkETUXRHur/oAJhJPVfUs7rLHTLyILM
ZA4kp90WNxvQkL3wtnn3qEQkAU7vTAwrMlLT1PZBKL6Aq67xtvWn2hdrnE8wau3V7lzYX19gDkuY
8W6qfSuFQHHN0WTfZ3hivC5vOVKoOYT71SsdAP49xGZCz3HQCKMeFcBMA6JS6RyadImISf31Xqnr
SWTrCiPot8RoMqF0I0vM/9e0kj+wfsLhEG6+IvM7tR/iYxlQFIq05+jeapQc9cEkzlnqZ2AA0AbH
hWdditCnKdsFYs9WT2bGLYYuLn46Oq5zpScqhUnEvKtFbmcOnkhY1JrG0r99mCCQmEyzBooBzxjm
OmVZgO8wZVADsKlSaxTV/x2LHl/tekQJDVVI/ODVmXbplJR3wipYc/YVy2N7dVp/kp54l878HJAU
ZKU+0AB1eqjgNVgPNx75Cnzz8AcCY9YwiD0j8S7ino+RcN+IvUHG4/m4mvSuIUNdfpl1etQn74Dx
TRT12jm8xJs3T2LJwvHItcSmXAMMO1c3ZX5UlFIN8v4TlauxuuCDECcE8rMzh3QVyvy0tVHP06NN
b57y5Xlsu5OE3MD4VPuof1t2vVp+H6UAHop6JeAx4SjfoHzzTfq4/gcKM2b4ROuJl72MsVinm7J2
4MHHE9MpVIdoTmvJ3VKA1+2MkSXGtlOXqvX3FlI3hHSUEv0vsZBRLyzA60sICuyooUucc1ActkuP
8x/F7cqOntP6Y5plmogc3tzw+aGfV35ebMAphY+aprwLqLCOEZOqQiSRRA/adEJ4WWKa7rGhC94O
C4Zs7sJ9Vs0J/8y4JDg8fmMXD400YBKy6o9YsxJjif8P6AxiEMCXUHiWWo9vfkfO3mZK84O0oZCI
jAVjpeEGHVp2pKAQgNoxoDydxztQH0CmfigN5Bo06imnjAxQfextXNGHDjYLu42eTLP7D96hGOoC
VT3zcORQHJOMdJhL+AKxStvPzh9dCcuPuTBTZEdpBPFKchicyEGByz8PM3XbOjOY0Mi5YvB1F5cN
vJaxws2dpPU6hgJ4hkRV1HLdupBuXMM4ngpnQZIp48BgUOCNE7jIby+auiCDdogS3w4JwwcCrMeo
a8yECcLYXDTTUf0dd4/gCoaFIFR1Yh0JKPHQsrGaUvMwrdv2c7SFJAzAz2UrvpwHXVqrejUi+pQF
9h1fk+m9wWPxAkG/b7IiY1Zrg8l+B9lgQ3MAGuY9tdz5QSIAtiW586S2Ar5ZsylwEIEwmCdezlaR
T/V9u8xzeHiwHEAcPSUzkpJYnrPG8zqUNzx9/6p+zM5zr1RUmWAc8y9eru8NCp8yn+aSzqESrttM
5d348nUm5zVsu790Qr8tFa9dD8JeyS1WyeWlchhMwWfh4zqOcTRP3MpklzvVC4pXRBp6WM/ZdUSj
NLfxqmhwTJe7k4agmE8X/WYfOwXodTtc
`protect end_protected
