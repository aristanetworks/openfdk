--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
R3hf6QhMYWplPIyVzmYs8abKmTI/Mh6mSopaO4PpjMjPdXeiYLk8grE0aUbIATnl1LyKNT0obfhz
2f2of+R7w+tf0SSIhCkcZrnnfhYbEHu4rndNZYEqIPo/cgRymilMapqwpONgaic/b9uoWbmtdJMR
SVxGektUk69vB2QTiO4uDn6MV2D7rPPIApFP5Z0aWz0dyOTJtkqulzjKsrysnRAVKIeybcW0hx67
EMqZYoVEb0I0mPHoHtTDoDTOx0deJEa2lX+fXrfcZg0GtAxSD8WCsW+/C/qWI0swiVrTDPM/f4FI
VE5bNZNS+RcZO4lNAWRvAUyKFiQEXpZg4Bwd3g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="5V3EUj7eaCscr6EhllGkEyxaeQN2CD3rxtYJUJB+NDg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
R+ZFK4/vSKoZkXRehjqFzzWfU8Gy3Zljbtz4XsMtdWex8V0lI4kyrZNHEi9anh3B4pPcGinIpelK
z9JR8QC3JBcM5uornaBD2yjs4IPrSxjoLDJGAxmp/PVd8p2pueBO1WXjzahPFoyVUucN5c7Whxpg
WZ7zZ01p0tmTyvpKVD047y6hEEVdUs3yx1LnZOOzDk87dDxDf+YAdw2Gpi+qV/0j017z7Zx8g+Nu
p5OIjRHzb+LUQo8MaWQSNn6dS48vqMRX848yILUmPWb/dafbWZapcaiPkFVu0AUTOjwgVrBt6EsX
pFoMPh2H0hRAbBAPZz82haJhcncfjbgoajntlw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="m3v+THawiBKTutIBCTeJgEtkf4mR+bVI+YVVRDS0+lA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`protect data_block
3q0tBJtUmPsUPgdDSK83bvFxTQNEiDUMp1eXmBdyx+OSlt0xGq3xujedm/O6Md45Torp0L4l6hmx
otlRE2oQXyMWf0h7d+Y+X7i/ZSljFY9albCIX2FRfy2UOinln3hfsu+dYT1MGR2sBng4zredSv5g
74KWc6G12qjSC/ZlZo42sdaeVjT270rHMcomIwYKQc9rQiyo+84DyNIKQreD4fSfV15hSStQE20B
hSy0FBXDOMNJK3IbdKv/XTeJc9lnhqwR3l+8ImkKwfB7aUDg3SVWRx2Q27Eu4tjmEKR0WZwPFYNG
bZkJHNdn0HMK60kW9i/hs59F5TWc4TI/V4pCXg/96Qnf/2msAngtl+mRfPp0FYY8BaNq0EsQx0GF
3nY09LqqvwLAW6pm4L9p3NIepzYJgAF3lGmPXMQJftmroDvY+lq50Hs/s0DKd59Je4fql1QU2qHq
QhvIpgNQP0Yts2HkFuAWIPeFSoY4l51tMeZuFVTKb68/WvUPPyhIzLEpUIUu/2tXpwER2w2Ik/bf
+BEYk93Jznvznl+jNDSMvVZAARUuDym/tzGkV/fNbBWotrn40evT7riDdZMimObY+H/7mituTrW7
I3PttWVqcey1zZd0V8cnG9xg1ALBDxcFoEdgN68GpVgUv6EA5tzHQ4l3m1qW26+bKDszt/Kw9ECM
KPaVvnBW4dggiDYh4zPTbLlHHMJ5PqEz1iiw7zv8xMRlTfenLi5zHW025qbQSzch8k9DBvRZoAkK
9mN2r+ZZC1kgNL7bLxTkLLxeliTV63GxqU1Vy99461Avpow6oQTUIcUjTxPhJe9sDW6s6F0RaW5l
BHqSi9yiukpkNk5ASPUija/jtw/YlJV+WjC6t6ImzEL5/AVx9hjTLOxJQhWYmteimU86pO4vVkw7
OGs/fRzjk8nDkySS1IkjbENYECstmRN3VD8eYWzQvdm9d1ZV46VQodzRfIS4AAsuqgYR2s9vvFx8
EbverJT5lt+/GLD2nQ540ZN0T9v29gJu47kpSXI1yrx0zW0SUK7KPPRUWKPnSNE/6QEEHBR1e5BY
SWzOR4SoDX6fQ5SyfFpFILgWgw/HvnQ+8m6Ca+bIm4xXNx8997uICFs2Jjki8M/ckb3pLulBEoRD
ncP6NgFpMHaIV1AeeRYp+VAg5bHv5dDL7545IzxDe04qlLEHfULymIsiZOHiceupNMi4/R6+XNvE
yEKvW1UBN19YWuvdjPTGsVmoXpLgp8oEiF4cReGKFeQsGISkWr8PLjYC05Ckq6T83IuhLVAvzzyO
9K18o7fdb/HwHCMUtSMKAqxELPIElFEANuLZ6phvbwY9OH43OaFqzoG+l4aAxd6iiHuLX+v9RUiC
Z+ouQLDd5mBC1qkVTNxXl3f69JYgpC1okthdrDtkMRRgUjED6FBsy+Q0BHISKMhiTT7K6Q80qs6N
q9v/WXU2fHa2ujFSWYAwLpdH5YH/oR1jM8iHQKcBMas0BSjSQpO7qraXis7GasvGD/e0kWcGq/5o
lesP8cGfPWFrIjUhvd6++B0sEBxQnJZhbkzLa5H6+FZnjF8Jh0ffVxbargBtlJJtHIaCeN2rTF4n
V2h6cM2J5rDGHiJDjXdIdMWev64fVQsM+nielFH/CeviWn1Dyh7PeP5zysja8HLvHdhTY+M8BW3M
lo99O9Ty2IssuS/CHqpwzmIFH7C8RTqWCnetKkiacz5RcQ5P44Gi0fWRl6YMSqeHmSmecDknnqim
NIT3dG1P1QQO5E44Yg3LlUKkXQo9XcRK/5zxuJ6r8BFLHL/rnxPovqeVnOBmWCgQOJ5Wm9v/unl2
75YMfFiQ6NLbFdgqpa1rP36zDnV78dnZZwAjmoJx3CvBNcLvGPa5S2NucLiRfG5XRsCY99DV8APS
BMIm9E97LhHrRpG3x4rdKHirC6KlH43VafkklM9nDPf5aB4QSMXEnv+xXGGIH+MeK76/lr6zr+mF
GeyA1l78zTAorEjlwFKMnyJk8uX1ZPq4XzPbGjHtG7SLgwec4dbGIOcsu76Qvk4gz0bT4iMPrqTK
WLWzRSfaeyO1lEs33FqikdOqBs2R6ZBLWoPfe4AnVR5jW6zk/GXdnNhsutDf0QM2YEMrJOXjfbLx
PGBcOibRZx096tzoIoGIZ3nlqdYQroSmClFSYvx/nHmqd4MZvzEDsDLfFn1S6dsbW91nmh2BTtXf
BJAFlsDI2ykK0cbSjrAa3WayocthhtsAAzqDn9IoB4je45qdi1eyTR9y80njZys2e4jOAnHyvhh/
UZteHl+IIrP5Asps2w8nO9OKCiw+kXy1krnv2hFGOe/ywOoWvixPUcQ0H4Dn9NOhIwMc9sWCmgbT
o8IhIHpxrWFi/2qpKp2O8Evg+jCsVlnU2GIZ1TzyMYUCAeKrXbTSHmiOS3qRBHxk9mSGqp9RsX/1
Hiz8r6RwSBTFhgLyfqb7XxhgDKMQYhsk/MeFlzwHrI8FGD+7SSy8RtgVMqb42m+FNyea5++dEzZj
qzwRWVJfmdmugHFTkCP0Rzyau6JUZhAoYUmhm2EY1eCgAKzsohBAxOSSQ3xUQ5EhVu+CxGuyhpLt
s5ng1VKcmZVBunLnJbmm+MWEDmmunPLl6juAIwIUw/6jX9XmvnrJq1bZmQadN9h4604fYolNLhgN
oy7GTpF5EFfwqRSQxwamjlJyo2CDxYJ6mPFrUwwMgoyMEmVXyBdS++50LdOLjZ4ny4b4JvIfQ1/K
crek3W43W7ug5Lp+Mg9Ts1/UlTl8vBPwI7h3yh6ExDsYlFExntKU0t8p0I+xNuhBvnLSUqRSqh0u
r+nCriQDGie3xvWQMLTMgv/1OCBRuoiGHHIZBAmTkwC+ajqPV8f6HaJpHId2bxMOiQn8R4DJnSXU
ZL4igQUZsYHIwKFWK5SOPgO5VqXNDaGFkY3F0NVsN75hnMc39/TQeURwJlObb2rPOptT5LqkPYXJ
Q9oTD4n3pO7FGNr4fDZFm5hZczZtBZku8A7VtpNvPjOfidIaA0AxFJ6eO8H77klWDvp/F2rJo7gD
bnj69AFt4HsXCpYjRO/8eFuQJ1XJTofD9Dy/+YfOVVsjjVQsumEsb8OSWu8pt19bHtIWO/YHmcp5
dt/+7cR7TEFj6pwWyMwU2MeDr2ptrVURwZJwqp42zhnDuWiFiu9FTIXHM5+x1kWUBOib58GSrO1R
9FdXP2HSYKXhp0npnQmIdQbc/1u/NlIWBuegP8zNiiIDbkaad0apQttxf+8u4W5D2QFU5JDRO2pg
jBNMHJKOR8F8+Qti9Z2EbUtd7QPSqQHt3W83xjmVvQhY3qxvnbuVB/CQusR0HR5VXgeTA+9A7qdb
6eGCfwdTaDopNkX1t2U2sLNFRCwRQpDhP3yuNL4+FECFMTnVuPiiMWdqQ7iB8Qqax5dXSKLPM98d
HSZXvtVm8t2/L8MsSY9LSEmxExLrvwT433BK07bwB9GJOSdte3pr7TUQ5QA819z2F98mf47OTInb
A16xzZmqUHtv9UVC1w3ldXBp5hU7Ria2MY2qSWZaPTOX4OtQBs4fx5LiNMHYJwofspsKn9A21+qd
NMwHHPGGuGcM/sZpPrI2geH+sv4BLqzWDWk2eQm7LjHIK9kwVFGkXBgQto147u/5u0GquTmgEQYq
Vj1XM3C8hHAfBW5vZ1f6MfzZL67fuk7KtrqxfC/CYHKb1ydb2uGwF939iBrQ2AKE/+Rw9mjdt1q/
BuqcNT7c7IVVaUMjTmjQjeD6cwmkfgVle9WHHokoGGdG3Nn5NzRvP1Cvyqcqg57lm12IYX5p3b/L
PUg2IenKYAWDULPXUZz5aEUjCtw7bjMvsEdACDBx7gIxeXw+3y4ciGqqVvaoWUTr3vqrKiUp9DEH
rrrL2+wbhxlszokQVERuwWjYJbiJZ0riiM+dK5TpHbX/3BlZfJ0TRdbkVD8OUwlsi9sdKg2tRlVB
4OOzIxPgmn8s8CW5/I0BJEJJeZ9xGa1kcj85wc+nzZymTeLKT3uNa1BIVbeSIotKFNR5Zng7m6Q6
CQYgpMkvOP3bLQ/WcGhIAq3yWOhs/nH6bbn7u2vJ6FmoE2UlWWJHDLU52xBoTfROkYxJ7xzUreQJ
l3eJitgLrxGMkLbAfR8pBOdQy26aAOugm8NORW8iyfGRElKVsB0HlP1ay5pkRyZJugtI2SAWXoPI
eF90mX34zAQyhYv+drqCZSEhUxJpRVaE4DuXnvIa3IVV
`protect end_protected
