--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   duplicate
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
daZuXD94Gnm/K7fasWOmH2e1bv0CnMKlsJRfWDfq5gTqXFZj0oms0sP2uWxdPI6qNOSHQSTw4S8j
+drXzrhOm50Mz3Gnn31l2RfMjJIuNc29yCcniqr1lJNSZcxo2t4nsqny2c+UrqgioRQfNPVcc1Hz
qMyvsohFFz3l9ZtPW5EjNPGbvBhCb/cogxwqKFGyKtBPhZAt8J28KT2W3LIhqTFgsAg0SV5io//t
+cqxtjQDQ06D/2CVqCuUo+ou8p8aDt7Mh60V9MLgkPoH6h3gFDjiWoMm3gsZomXPwL7JjSCs+fe8
YNewcQ8WpusmemIUCCqu4IB/BCvdbKmE1HpdCA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="lcEq3hHqgmduNT8tr1/nyK+ewxXc7/XN8THbfINt2VE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
lPChJEvffF0e+4vjgS6UyFvDnuX9KTg5nWaT5yXymRRagffaeJcpdyZcI68aEvIKlYPJ87FF3Qct
FCWJwoOrE0XWd9KQJwetI70zngJue6/0YgTCeBzmZNJ8iBy5a8/hPDwYQLsMRG4cfSNkth+f5xC3
dr9YLME1FiXpQIBKbLn9coaOYvgD4NUzyifSQvOaoTyJcKY2YHx18kZf9dTDS+qz/GwRXT7yG2o0
MpMX5wrzqGV9UfZlABzLUcNRGMex5q+VcIJwwy//Z288u+u7sN9ootWGzSg42QRT4urvS/Djbrif
CLMqwIa7qQtkRt35c6/oRuRdoz17vnebeQfIvQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="HM8O9jSm1KUsB5iDyd8ZWx0lcFX4xoVsCGSW/NwCqeY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22480)
`protect data_block
ToaCTlGe1G4k1wGsETJmBJwSAbH+n7vRhiMPm1vDmWmc/aP73kxWeHHHk4+HmrppISm5eyg8Ve+z
lxmh14MQMWwGJBliU0QxcRZl1VPanuYeczubIN3sAacZSKH8dekYBQfPkA3H8Tt4jBpXVdjo32fL
JVY4UCDaDzQF1/gGVzz8kYP6yuEd1Gi/KHrxKSu6UXlmtmvByTFFg+KayR9TGfavwNWLpBeFQ2N9
XeaS2afqQIgotd7A4GEj14c0iuORodIxyhNsoUoeJhLc1m6RO1DPjFtwWXbqdKzv+RecKjEZLZNX
fwcbME23uxeGMS2vB6u6fHxS4Q8T4wV/cx/6jksY2gPl62p3gw3lNLp/ynFLI1MhGtRUchXMxJMI
0OeLkiw2ZAEp57sJQ+cWTdVMTW3fhTm6PxXBlzs5vOmuoc/BJ07uOQrTcN98ZLEnCUUfv0TmmTBp
j/x1NBgBaYgnGyZb/dvWKk4qDFah2yt+N1GAND8bbULCrYISYWA6qxYLDvidmA4kpnn/oQ7gt6Qv
0CNqT63/HVcBxlayWHUZkjawhbp+w2+bF+wrNaFwUi/oXKBGSNaE/jrl7DPrsMbgTbwFnIVobR2e
DEfi0vWO5PwmeXKrQmRo/XwiIV0jWg7Xu6+/XEsVQsOsJvgLT/ELzyMloVitQjss01xtovwwaVYF
D9n41L7SjXVLPWtLo8HI4dIm/K+H/YuqcJSLshKq1jXzBorO0vPlyfB+pJwWULFtDEMrRIluOO+A
v2D+mFW2lEzJ5OSSgg+v2ol10k5345ye3nVstcdbwVVQqSlVkG2H/1ONV/s/zaP3M4USSR1lLv4h
ubHCMs5/iI+htm1xu0E1aC2UOsLiKq5gbpMQ94yzym42hLaRKSa4xzcZrF0L/rKAfE1DH2ZOF+RK
LXaQ5zkRSTfwclRr7GgzWRAbXlUHBu3lm2BOBT7VPd0w/M6bntPiRUhhs7w2j5YeEuAWqZD7mNpD
CEVQAFzz3Y59ipmLy962IdOneZfLpoF5erEjnf/LS5A7/TZBTc0CwyPrpe7sffHprbLkWRw9gB4G
KS2dn5rv6SXHCSSk10jNfSQQ9TBQble5Rwt21spfd6x2bH9tsi9IdbOk75yvmAGR2MnmRpl9hDWN
MXgNyDomc51bmhJaMsO1bv57G42dnsEQzn4/21rCy7FIDriqPc6MzcXI/OChoN/LMBG2cBwtcPfJ
+ycN/rZXFm44SyvWDZ6BKHOwgGKJ/WJztd0EioMgzwPp3kUbukiDqjuN5H53MZPlHnbzernf7Jln
LEDqcmwM6PFNN7JnJAxByKDDt734swbtUPsooFaV+hbjyFuUC6JLFXk6HuG6hvMLEW6M2zSZvoQa
ogIs/z56ZW6d37eHfsYzTr2MRtPH6T4kwPizRP1tspvWlas6IcCsHJ7hOiepnia/DGgZedJZNhkz
/gBKgtBn/kWK9lJr5AO0q8cGcu6USUU5fsjMumzIRuYNndyqZIKU8WlPc5sngZlPyfrUC+Ne+rjC
8lB4QDCdsZOQb1hIkaZFzKIOEHylkVpyMQwfG5KSp4meCk1R0EVePS+Mbw/p63mXCLbEHEdyzigw
QLY3xOnHcPaiHt8gzSj9o0xGiYXrJ4yzd3gVlKP4876tzZwJ/IQgmoIm1SJmcFk2QcJzP4loOpWm
6/KDmRgBOidrEbKewSrFHhdLh/caeLQZJXOsnBCUnLpat+FQ0k0aOUUyVtMa6J510sMYBjY5ZH5E
KWmebmIBX0f/Pgm7shZsooIyUKJOBOq1WO6Uk06AyNejIYgHNPj1f6kDgqN7uhpqBl0JivjlJ0mS
gk0mLbascld/oEH68W/EJqSPAcbsdZv6kabqjapRnIQDUk9KS+RA73VdKEAYm0mS3/HMJ5ABxMsm
DLsIbseyTYWvpDO1d8Oa6e6BL2KGW8vwTw0gV0LZ2BSqRh6ScB0XdrfwLZdOyMzbI1KZYuyoX1Lw
nsbJe9nSe5077eiRxKQz71pjewc33yxRTmZLTxyYbYOBhz5enlhqWnQHAs3ouThod4DvAjM4sS8D
YwShIB3Qo0MrP0gb5/DR3MlSdqtksBsXAuWbq0zG6i8MT1yoadEor2QhxdcHI8JJkJIM9KGkPAq3
5Z/uhDgnw/2bkYNZ//NjRwX7uajh3rqIx82nxxFYSZyZK+x6Zf4NYvUagfy9vuVNMRp1OQPfDFsx
fjIHil9wJWsRAXNt65Wknx40MFolTO6QvlkmTHL0PqMP27392hKppIZkv2d+0thcGMVHa3671q64
Ka4PJHZVZ3sD+7BupK55zdc86On7/jnZdHCHsFhe98NXTJ9x56SV/o4Z+MgoGIvCKbFn8quwrdv3
0P4JDowkel5tEObuEdFoWQc+iy/LlZKL1wQ6oDRd21ekOVnanBqmtLYC3Oi+zLYTZxHLpzsze/9O
DV6CnsFS7a0SvSQltkmbbxtVez/I1HDYn2YQPtUgn96I+9IGKEuaYauWvsYO7/qhAxwJknqGTeYu
5jIJ+YhY9defyCa6OvvTcBUeY5hDpFIpexFkmCjxSp17QWDZTg50gT4AvjGMx0L1CgHLm61aJOxw
AACZ9b5snMzzyaSWx+HUXacpWR2G12Dj2eRqXhAFqWXqtPPZhboz5bSf0a8qBBUZHqIYJipE3BjG
d9/oXnK0AChFjBwSML/g47RkZHQdpsB/Bqdm7hLAPb5cthuPotgNXp5LJm6wWHXVnXu4Uwixcyfr
pkmQOROfwmulrSGPnqx2IJUkZenG9EXBU4A5OShj5vSGQtASSqD1l2rRnZuC/Cv4P9yIh6y9DiFg
KbNFC0FVJ8MGlGCdH6K/2+cnGdGS3aTzKip75+EoPyXbnzMP5Rkb4BSK9lphl0wACZDwTN9SLEgo
ns3L8idvqEsxChh35R3afbwNocTW3l711VNEpgn8a0alcCam/tEUtjvsVkjwd4dtCbzSkzxdrsrr
iximLkrnnbow/3J8D/xJPnoQb/zytZaG7JVZiA2OVlcHGyq+QdrwAu/v1dNFArcWefO6yay3gWAL
DPqCet3bZNmKYW/B5HgWvnfL9jG1dzFOZDt2+uErAgAnd1//EvlNF69GfChKM+yebRCmXNOzMo6Q
buMMNcaFuxeTtyKRzelDxo22nmoDIjhmFK7QNwNr/jZ2PDQdeNmNCTld9n7cn+q2WO0T+8u/BW6Q
QkqWSsq5GlQFGqBFhIuH5lXA0ny3g1SD1oXLeOwXnz0OrBBRxsQph9J2IM24pvcE+qLU2cXjbA8B
jgni83lto1YFLn1YfIode0+1h1yOIj9KoP536eDrYmWFk0PSRIw+oTP6sP7S5f0JHOJeOVYDMj/A
lrOA8dTX88An1TOJfEgtJ3dqyaZdqpp+yOJMzFp3aIG0mF3LoLGuRTx3yg4wdPvgQkc9ZjYY7ja0
xUyxwj+jO8wUnFN2npEcxiq5xtmJHZQW2fnjLeCfmfM/FbZ8qHTRVFeOXhpHPKBjKZ3NrRi/srqE
EmUx20K1STkKEmLBP6i7vIBuzRc3guZ+D6TCd9c0BPSrttjJS5il3qpiESMJ2IN+vUsSacOv9002
tLHPmqbYBckJWeZ+JWbM6TxV8pANy7vezgNC0WoBYxrP/yVPcKebLkzd73CsX+l1jFN7g06q2Ef8
9SBbQGT6aIMrj+DZcTJCYtYB7F1+4dFQXw79zIJciP20nwYPY7KpSq89oaNxA3Hqc/zlwQH/tLgh
YG7HGrerik8Od3HKXCdb5TUWalCW3tEJc39jA1jVYIR8MSp9ORQGwBz+cru0rYPsuOmszegazpni
jc1oovNwGq1XOaDDRED/qRff6gfWrsrb/hIqf4s2bAFP8P3TFtex+LIuulaCBrPCXccJbrey5iDG
WekMY6dd09piW0r6AlAQgIrXvz3pjIKK/qlltr/kioDoyh+ibBQG5TMR8Ut8/Ze2GZtNDwVWYSyH
Ll44SCV65DrHgn/rssJSqD3IyenySodvP6ZtJ03JxL6xsMB4BtHRkOcTSdf4a/pvXIEnEvg0Y0d1
Y/TB/1Gw5WPUNz1cgqjZw69O5w0ZQWe1E/tj5D4lHqAvfTt/sji8eHm5Z2wq7sqcb4aU4y2sLVf8
xkFHFT724UdinYwbkbJwshAEIfWCnYh9zfcAAC4Q+5Ds40Q4mhO4f3druhXsDJ3E77jDiMo3y8cr
SREhkHmcHs/LLqWytmYfIopaJv0Qrj5AfHYMmS2NyzuS6DkkpRDYUCEWbLygDDJnqmhYnx/6E73/
cHF2Cv2+sVLawxPYAPJ5t1mgT6TA0YDozQ+q/ykEiTeK2Hho/PwPYMO8v5gVTreERMOhSy3tQ1ol
9hFpElAi/rpehCeMFE9bJeluuFDhEg01RNZAgve4rPM+PxphbK2ywqEdInXmY8KAoBJaXwSXADDl
Hhs0Hauxp8M4SD9MXoJJCJQ4hNNr/aTnPOkN0lDcOqym9eAN49UX9LPZpko/A7RUY166Ci2TmW0V
BuuBPNpi6XMKP4ACzfnjLpnSTA2u2mGv5VOkRBoNgDN/shauO2l/1u1mMG8EDeGeljYjNm1Y7Qnt
cX90nsHPH5EiwgHNE9CciJt8cQAY5eGY6qr/46QPGlF+u+MS2MhfMQjeiF+xkPYNvZrch9XY/4Uw
YHr8uRvXYdQR55BqA904uxJMAjlcy5CYb0op4AYy2RCDq382auEL9yURSqG5Ym0cTym20l5aDhKv
Gy85ONb61sRc6nyuOQ6Q8/ykIN2u1fi/k9YIH10iT8b4VTTPaVKFxTl3bg6Cl++fXQrAWnIm9ffj
Xt6YW4SZbvNh8/YcVrHHf39Ow+SPvMGb+ZdZpFKg8pzA/rz5rLUyJtRwgv1LT14wcD75qqHC9kHO
d+jejwcrkN6btqJP12Of2vOo0JOd6cVY7voBYM9ewLedEfwS/IxarwoHMzsoB+JcF6Ps87qr/Gg1
HLwGgbkCkKx9TQPwPaFeovGDuf3gMiBaj2lMfhjZKqzRSLG2ejWD28pcM2DpXwIDPz30zoExU2wI
fjjAdzjdPzhkWrzH9bAih25b30be5D5uTpW5SFZ541z2HId8fKHDO/48QHeftuBPz8nfWl+chQnf
1DGxhTuH9GORRDGHEfnd7pk0Nm+py0Eu7qXxKZ/DfJy/PnrsXv7o9j+WDtg+edPc5VvnA3V799SS
fBNkX7ms0bxlf60URJeY2lJdEcHHSsLuX09MF1YWG3JYtWnHxvNf+aFlDWsI2FeU7QEWfYGccMdB
7ygdeL12q8a7GTVGfalFB5bL7ZAAGtuMJw+sRewAugeQ/PRFa1aZXjbR6iWyhPtZGEuNUJTYGC5g
64t2MQT2GSPGhv1qcRfyTI9aixgE8dUE5VhvNzcv4eWBD1LvJORsAcITHU6XkgN4A4JLgAs9dhkc
NaF3lXUGQtPuxiDITvpX8GZC2r9Pk3CI7Sx+tJHxAYT/DvcLPfnCHnJL5U9HP0ON62MkfmP/1Cbp
rwCzHW8s/H+pRAJduCV742rQgyKBiLeeGDtSL+LH61PkmPtbuUiCRHCEYNrrWHkskCTvNBFn/fnr
VnvNtAiFs6w8BTOJ0rvA5NWNqYK6fM1Og1vPV+R8Dx8012dz/4xBc5LxhAFwtWtkRaKsNc/wY9O4
2L5HzQqs+WWKpeD95i6Gt+HmfdYSw+gzCeIqJ/i3NsuggIJsKxJDVQcWPJSKcnSvfTTCU6Po6CQC
Tj+zlBzs4re9w2Z0NTTSyxGaIj2lxWIjZIrkicsvZGLpa8r4xk1pj7YpdBY863qMkHEx2o2TFxo7
Sldz+uVpfd9JKgZGeHpu1gWS3zuo7vMie0TNiuRL8LcDaxQbKI/1Iur5thbLZNmMBsHkaxGgpDVW
+IfZBrtvURBR8WjTPsiPXaRmn0cX7857jQnDyzdcTaN+DbAB8ICD4PErnms/sUgvbfxWoHJ/+/dI
iJDOpdhevUZngVKvQi0PJdItCuL+HLEUgAcE9ALkHr1CUwklFeRhtgDIWbC6c3VHGHssX+24/IeM
usz2KwrFlh8hCDtMI+AGVl7ZHAu7fInd5U+ynCHWIB/YlOzGYRfOevIq4i7Cz5Wo/Kjk8++9V81+
/T19IQqNHOScH/DNUIbfNrQWOvg7GG1WTraZP9sbBr7Y44BXKpSewH/NKcVNXkcC2G2U7JGpSScb
avCKRDDzyL0YMYWmSFQMHj/veUw1/jHc8z69m5sNJ/ni3DkaGBDlkejj+wfbO3L+oFfAUi38aVRg
Q5RGIcnmxKfkSP6NAaNczv9DPrIyZGDGDatUpGru/UpEg0g2JMHcHSwE2tCvFf7y1E9GL9UpYrSo
feXu1vox2q5NvJOKmTmIUjJqoQTSocs3m9iswXmYNlEF8KpAGakRHHTOPY1Huiu5ikimBeP5SaaD
HxhFXrNH01YLmFjXMuKZJm9zlpta84I2srQqpDdhy/pwFCtvIS2oOfMTjypmkGd+bMSYY158wPy2
e17dtQOGexXizhRni44MLErShTMLsFmF3eO5hxcxeXkl8zeG30BrII7HqZX8lX0yD9fcVbMC/Mt7
A33SsQza097J/e3Oe6S33bztDOv6emnGD4QLKclwX0KjhQzkagPXTOEJL/whxWJjqb/Iq941UhUV
5GGUfoU+4ywYOaGsu+T13ESUow6ZoyXAk9YWdqGKvrfai7hi3aKzs4gCKrJJmQe3QkQt+CVO1bGN
v9EBOdKUw5RzhKHcct5SAVgmte2OTqUMUd/Wd1hZaGMY81QkHbkdZank6yNycyXjZUi5EAoheCnY
tY92qdFTdZ7Ec7watK/3Lby3cXyujpc3KYtCJeV9UK+B4893jAO0AyTgVJBFp1qT3WmQtqqkQh6Y
lepj3/amkUJQaDuoTNYdHGeAFlAOvv7OV1/owY3vC0J6MdzVsMd9X/XdLeu7oJJGPwsI7doH4/d1
T4OPtwHp+is+pempLzT4mQtrt1HuIkkto19Xbq65rkP9K5Y5/2+lZB1Mvbi3ZEzcsp/uhYRnM32x
Y1mbeZ2b38Eyl6V6qYPPnUoEHnB4Mz3RcMMp5albMhOlEhk+DFmQMAtWaUju6LU4KItCKk7Sphal
NUNeQP/LG2fs8LFWHqt29PU9aSieJZa03IOrFQolJbafGlbg7xOwCqlqlUvKBibXYi811Zu/M4cW
zDjoRvrWditeCxLrIf5cG2qX90H0r0BaHU8hAYQg9/9NhwlwJtEQGsfHI6YKq4toNP0skNSFnxyk
kUIX2IwmjsVgjU9rBVKjP9SqZO0FijF5d87F4LRhAQzT+mfJM7rjfKjB+x+hfQzoLaGTluiKI3MI
WOYnQzaHIh3qdk1HqvEn4GpHnpLc4lSTHnOW1H012WXpfOf8pH4ej0alc0zi3zOzP+tkRKzRVUnC
YO/rF8sDAYgwRQc01+++UBLH6kMJavh6a53pvPY2T8iGJe2zSHQFsPDFGnkhaSHKoTc/9uG5LYxH
plRDvH6ltDo3IVCE+sSR1d3yF/uQCBeA+NwvP+18SKcUE5Tzsc8q+aKu7IxNFhv3vRIgcYM1jxHL
9HRk+GUwiK6rHDGhjFuOWMJT9pzR3c1/gr9FDpb0zHX7OsUcCdzPBiKn+h0eLRWmJQp/jZytlQ3H
bbsvyARji8zH0SSAiCbbpBJ5GIPQCZ/VOvkRD73e8X1zzOZotfFniu2nDTLik1J6vnwCqkHZ7rQd
2d1JtmigOgktsKttA3FpwD1z9vTIcQx6t1DZzG1L9CEZYrhX5NFnrWomiB+9+O1wo20vnlfz+/vc
lNctKEhQKE+nTXFAbEN1/Hy8Ua/S6I2N8QkDujE4kbCVXsFHBos7DCWX2LrolcHrGVg0/Pr9sdL+
YdLMaBKeKxTBTtiXiHEcd3FH6S485r6o+v3Q/gu87DiSEk2QRj2RzVGSRDXXuS/JiVbA7X58BDOx
95e7QrBb8KZGVn2RERV/WQbNF+ocKBowg8pQ6kzzSLSMRunx6X2WFj7Ta+oKjn3ZOEmlSsP5VuTg
EzIDYBiqNwS9zqYdMZxqjRFIGiJyplhjQhODYalBo2AmSn7bd/GS3YJo6pUSqRjYqw1HNZqUBlW9
idh7H6c3HQTXb6DBLTE31t8p0xHkGa0uP21xDX+S2cohKbVVjrWDEsKEddGzNrxA/Yl2e0UgxIRd
/Mcz9y6qPvOd68P6XxKaZmMeN1wRxNjAHPhU1Nh+1zeo4S0zaXV+7LtFHwecbRzFj9xRA1+R2OXF
FUFb3wd01sAcFhTiwZAUuD80I8Za0Q2p9b5bZeaA/AjXTrVJLWXeHSuzbMcPTnUzQb5ykLHVdMJo
YBtnWc9Kz7jSMwEEQlIuESBEMK8dO5pROz2xJ0Hg8mO1yvJ3ECL7kXxfVXsYOJEOF8b3nuQciZaA
jQTKTrAN6/KLGZURKvvYCi/AnX9jfSKZ7YR5kqtkbPma7ZyWtcpZs6dd+lZd8m43FVpIgsDa1FfC
CxTyxL4vl20s7kmfC93lZrv8e3yd3Z6oVg7WXNPQ9OfJSQ1nf7gi6ISpFN2LQWTkBJlu/SWsICNk
mfxsfdnFAbLAayvK8PXStLCPyTOK4nP7OhsglD7vlY4dWz4VuXcU0MdIWwATT1LFNE9zsQTLfgQp
KYKe9Erd2YwLeocwxOMzLo2XJYTH6uqUPYpnUkdsqZaXMrt52sEY7vwr+lveXoYA+gIuNeHyMYxp
QYj0DH2CSG7jGluIR/qePB3QoAD2qgVuRY+avysO1Cg4wWRFPK1hmyvF0WGtBFTERZvDcROen1wP
yGlA1WjhUaBf/pRdCcn0dzom3EYn8yGFFL4/C06qzohwg1dI/HFjyltOXA9vQdZM3C17+7xgEj1G
bRiigA7ANhGkwjc6Cc1WsVImPwl+CUz7WM/DmGm9Mk4AB3IbT6dfrBP9RhkrkMAHVcVHLCDF4dTj
D7SP+6vDNKI9d8wteYEbQmkf9GVtT9mOo+2jmGU3qX9iCMmXFdOwxy6cyhofzQcukY4qsco63Itq
L5HDLyZDjDB2wO6pHIV7FwpzZyL99kIdeSCowVGqvQ0jBb+AZ8avTtvnWRrVeQfTFDLev3ctWalD
fNHPP55DWYfTCoNBuIJj2UaKtmP7ND6I+N1H1SzV6gX/H89OIaRg2rjA2AmXd6zWX+bAVzb3f6MA
cPWSnPZLOIuFUZb8u0KUeChKtvPGkKz8HKGDBbq83DuzCgMDXCyV0gDtzee6ozN0pMehDLT6YUD8
i21Mlr08eDPAqNEsPcgx79bp2zpeRTGSK4pD9JHGu3ElWU0txO/rZA/bPXCzP8+XcQVEt5eo6rKp
NmtL7OUoj8XQhLb4BchrUHzJFNtKVf29RAjckgFhDZ11HCKIHV4JOts1KyPPoYGmUekCSRfETdbL
7F00LGqeVjKLOBtzCEI+wAIuAVhIS0KfIlabMwGoyZDpmuN74zR2WdPkKJI9A399mi/ynPzRpr8z
T90QXSpVN2d9HNNaWUpN0JsaWQ7wY+yrKAMMfYwSfjWp0ArP5YnIY1c8dqaavMUZZLGQdqr7yn/s
kyjbJdBphl5X2noxXZDjbbn2os3/IozLoRGkHO1A1l1l/ODB8pzWUwKcMw12CywUU/BYOfYGxKNt
/8/EXzSixyCUTMdHGRtLK1GXCPITcx+BhYBhknkPl/kVLMSPlYKVverVHFCL+pyU58e3ZM/McG8R
IXq7XC5RMDgWQy1Az6AyyZPumyUgspanTfkvOHLyR+B+0ZW9B31TiZ+bi1kO6aQ9Ntn9IkJ3uzTV
bh9IfkfcVx1q8KW29AHZBQckWiuGyLXWqY8Oyq9zIMaAP6Oxk7ovdr53Y25kPljvxsNRW4Ehr26o
liWNFCWNewljdJtpFzVNbvhxVEHxyPZ/AdD9+shKNSWGu+Ag2X6H0eMzvUhjg3KrBw9erfuoOOco
Uql9IxZuh8pnNp1i0YExJtKdnc/BtmAmKibQtO9BHXvUbN9a/mWcdB45LwIw/vcK/f8/DfCTSVPU
pJVWF238VQiqr1HIF//LcpTKBwv2TNjFXJDhuzhLvy0PRBtR6japMrvmWryNZQgSLog+VvAhRZgj
CJqSXS5wz1fkInFSROzFwCtM8QsBDZ3LfXiUDnvoyrpCmbzwRrgPHFP5ROiyzWco4PuP4+Bta5kj
0Cn+VoWGb5Y2jD78H4QvYc1w941NwLaWvg975nyzZtcSITRjS3ZYR9g2qOo2Ojagg4y5FLGa3bGD
7e3IQbqNH4x67c8GBuGH8F1TwyZGxQiOgKamIKcULQl3SFO5tehOHXf1hJOkjW9TF14qrp9z5VV8
yacleIlO/8SbFaTp2DlILMhxK5iI0eLz0jY8SVHvO4H5YUtsjP6qC3x9lGp7IHS3ihnGqJinAnjc
+eWKzUFyEVX5IWKgzcJW6+nbVVM9/3mhytpWmaigOIS4X1JQ89Z49GbcYaHYZd0nN4fW+mjbnC6t
iDDR2x/YQYHa74DKbCr86wNpWcphLcz64Il26yYVdDgCzOFSDhzWqiUWyTFEG5LdbUSF4OFolWto
jSpRD75Eex5NrnZ+Xi+ax2FGQiAuhPWr0JmAyffVXrAzzSYMCnSDB79O3ellenibySG0EWtjLLBU
L9PO7EuSAGgGGsnTYWXtuxZJiaMMyGGnpUGPpqLqVATk8g0GRy8AUFFBxl+Ly7bs4TATN40s3Y+N
AlxMxu/N8k15215r7WZgzjfMmPgP5IlAUw6KruJAd63KtHEm/HdOsMLoeK7t1smP5U9a1gFjtEke
3j4XXh27YQ8l7Txja27dt5WFfwxpnW68qGy4cJloTvebwVkpBr73l95KFv8w92FKDVny6/bapU4q
JwjPreZ7hSKHU93fu5xHF2pqjwqtRuYkSHE2xrPDq6ljcfh3kddo6CiQ8kHkVxilcYbEf3Qr5YL9
uQp7bcVW/jc1rEq+J5i6JtgiDykIfKkHHPQjz8YUuWSx6qOj4/VWOSEZdwxsK6yO2+C2c5+lHSof
KqRngoHgkFeCG9IbKOC+DuWQjKO+rv6g/jQ4UOEQx61f9UROD9RCFj0QuyZ4qHpij11mGsNOTeXQ
KnSRNXGxBAsfogkJzcQenoawawumGdxxJYbZXbZ/RLe7mQz1Kw9vGdIlc8OulWCGyQSpfrzCZH2U
wYYobHE9gsqx+7l8FB4H9F/LsYcoU4WC0X5UtIJE0urDh5Z+v3y8uiY7q3upKrIre2+qwWQiQ+4j
Ge4Jixt4ZZBJ88ecuDoJzVx+FSxdjntdE9nSxSuSJKAV1wxq8ZxaXHKb/sS8QgOa/tmiU6SkoA92
1F8Vd0tP0pVxH7zDKC3uZPU1K83AMPOR4TpmJlDZZgaTFt1NBt1H+amIdwEPNKLArsNaXNij1jb8
kQgjwiP8g5ry4+fzZ+NilHQT/h54KuwGe3SBDwHGZSJKKCo77ZPnP8Kn6WyoV1aRaWq5Tq7ZxWd7
zZVs5kql00Nth6TqhVaIZV10hmqp4uL6SVwnSjcNlomde2n/7RhXywBdUgbov6u8xoCtthNpuJ8j
YnrqYjC6WQJiTNpyf0/9rtd1NzhvuvTUF84EUA6gHrjxSF8NwPK+oUJW7ZuKPVk2f2geC0jTT57K
ujF+AtCfLVUOo5TM421viUe1YQ6gsKoFEZMtvadF+2XcmWE6j0fMDfE/0sAmLQGd566UGlDdFsYO
MU+YzMpgxlqDoOYuIDYgbpXPtfI2C4ZAKYSZnMzH0hq0mKNmLb359AvUxTXM08O+aX2FgHTtVTWp
jUDAoG4q0RcFwWbJoDq1zV5tA/AvPd7gSzwFWC7Yx6bps213wrI6sEAiAQ2FkbYfDzA/+MeWQ/8g
bx6PYAsuOo+5DaHITlwILZwXjbUbrvnOYovERBX++vuDp9pfnCDVCHII/J57oZJdf+TB3MKLHu+6
QR5vkHOC6SCoo3PMqNGujO4Af5t0sitkNO7iRLOrLG0pKk9yD1rLcieQhnmpxx7CZdFD3Q+vFXXY
l4rc8QTisfHgEC436FTECbFYzEeB4xlSp7lTz34g0O6r5UfiZve+nIyKO5ma+vgmBdl6ue5Ts1Oz
U/eV+84SZ0w8xK0W/vI1L21BVRJ0ac5BnYdxAErbQb8Ws4xbfBPewi1rRGyE8HPAZN19R7vlTJxA
cuTvvfsp37yoXQOiJhLd5eblNdH9QuPgfQqFrTKAcMO4x+XtWlCIS8QNjtMiHFvJkmLh/1SyMsqN
vEZVXK4wGcZP51m152uHVr5aRJI149kLmCq9TfV8nheZ5yIhASud1FpkoIOBDPO+tpcAtUUxJLGI
IA9Ddlp6YNRai8DXkadpA9FHgun27aWSQJw1Qp0ac/JXFaIl/c6ae6RtSJpUNDdtzTBgajSdUhEJ
uPta74laBGRUjbgkL36GSn6g63Ni4Gk8VFSuT95zX79PRkeIk6nPVoomEUX0Pnuq4cTlcl0RZ7HG
2O1hTgo3tA99W+K0NAe4h+VcQGeGoVd5pJctuTcrSB8egqoQVZP9ciF2gYZDPkfa7UQkezSbS/yo
DiNJMeRAd2f11A9FqJo3qrE4vfHpKEpxV0OQG87Wmipw2UVAzO6O2kmlmLnmnPdnYjd1Uu/XEzL5
1rjUa76rdigzKkm2wnpNISae4b/1ZbccG3uJfYQ1NKx45GsWo3Ip9RWtWM7jnLWuEx8j5spM4KpC
FryvVlL3lFPVALCJMJDPTX7CVbRJxxWXpoEoyPXbvlcDCMbLEy7tYWa386Gn3oQnpyspvsDgyNE7
0I8yC7eW9Hg2alTer2JfenpmJoJXggOCWznR3QSv9f9v8WXR3BjcvIgJmbDqO21G3RuBvEcIFC1H
dPSjdkB7qFoBGmeBIyxJTmvzcSJOLXtgnVyzrnY8OXlF2hvHXncUTwd8DekfbEP4zkAn60Ouz67S
1zLNMiW0TyOFUY2x445b5VOG+m8Ez0cxz+ZOsqddGiDhmPsY4s1sTBigOkcIunkVY/CpHaxdgHD0
kbSxezGYw4QsqQLciGkkB7FKr9wNSxfFxxfD5YLBm6UxmbZtxqGciRXgp6dub65AqkCLCB3zzua0
Z1lfPhgbq0wvkN1EqgAYBEpd28nfmM3AoMFjkE9r2p3nT5Bm/hj0WVx+yKp+pvWLiygl4WzP6F+o
4neeMPQw8ikRAhT7h7OyX/uBPknFsECMNTnz/fG2x7N0LAn9DSISrwF145T/95qe5t2qOTIsOEHD
qsdA5hsR0P/D5x4pLXFDPzRyeDxiZDiSO09+UlliA3VhmV0bKdZAmaxdn/ucj+t9c+1anwr0Ad+v
6PsA0bRuz+1+g2qUphf61ee3WX1HdRuCXKZhb99ZPh2UtoNmMUtPpisqvogZ0F44CZOrLAWfVLja
2aKXn89sNoAytX8Ixqf9sk67WrKiVCPSbscm0JaCBuwwhrnDzF4m457QmgvVQKEwNH7U1TD+7527
Bwm0IKf/YoRqcNWJjK66bO8KD5kGKk6i59HQH6g5WXQHJXyJBeH0hVWIfZ/zRzZTmiHcTaAWNbNh
+WKMMKL0tUaXrbV4gZDJb3+cPvqgSxJ1E8oOUQKRPja0nHjBCsjWQ+8XKeiMBEr9XDefNHYjWIh9
b8JgsBTIweSVPgGxd8rlnRVPn8Hh6ko25go5bvt68fV1eCPactpz6xDHK+XP3PLc5dxKEp7llCne
9pKb70HHKOh25vmz7b711UPa4RdlYTOJkNN/Z2iA74hnyMjQ+b6objpSHCm7ZNFcSiSj1g0MQWWl
f8gqg7GBblMTjg7tSHfiDD1OEXcbjy7HCfzR9nfL+RktF3hC1R3+uNyh81dgiopu/jw/1DPpawZo
fvadbenchLUqQzQbTP1CXQxB1g5b9mSgbOx21eMceIjh6lGilgEnPek5Yei9uC1jONjn9hk5PShe
1s4wpWd2gU2nKD8bXAPjIDH1DPXQ4hJZ+g51Nt++5VmgOr16zTQQ8WESMFqDjANonu9EebsbjThr
5PyRDGh4ajWs71cKO4sXwEZAwRrRXrm3gWGBk4+9r6jB2V/N/rpEPieaHYyCgD1fmTBvnhCl/+vV
WX9DC6q4MKhe+vAa8H45PY4WgGlIDNUUPzWG0QgZVIFajD0Ypr2op+lFMGH4jXSzfFEqsLe7LPYL
OfiCXywC+ERoCUGgQHTmUiQbEJgCggg9uQ1rAmsQr+WU1hOTJ1VWD6eWhVMyeZUceqNjSuWY7XvO
C1nTJSYY3CyvXXmFJTlPlLD+RDp9ZnKrAqE6AEK0yr37Ogo7DFWcWz35z3RoPTCFOIUAvvdLhZdh
gR4bwJUULjzAeT7uP9ebRsAb2Td5RtJNLMYJy+tVl2CmuyMf9Nt4UPaC4339paw+T4R7QsNXiCHW
3uAC9B2MEmG851zfA47mNCRCgNm5FzfvaC48XQZ/fpqkB/pzBO5mdPc8/BuOMwslr5MfSv9ggKvg
XwlbG7um9CCGYzH4EFZAaFRRt6ADLYX9zJGIYUi7phnCnntBT2evpRQb1uwMrJ8V4jK0Tm5DNj49
z3QeOfeaV8wD4P2mKEfkS1BOkECmEV+rGmiCTfvlLoEhYQLFyL0hiIrH7uhp9SjbGs0hawzOhNVh
5Q50TngX+K0xDkx5fICOLP8xAFXhxxMEURfwLpoidoNBfPnOxq8PRVi1BMcvyNUSi4kckSH+Xd87
daqYwI3WR7PAKrT20kcKJKa26T56nfkplSD14rXSRHu9xqpsleFk+zVPIFCA3w3Qy+3bRd+3DDQ2
pt5mY1I4P5l+VkDpU40zmK3GPhcPaR2cDB0R19Py92LWbi2eJQK2NYbt1PTIpFa4yLVuFQg6c5kI
B0E4z3r/2eDGiItoNgOjuqF4innfu+9RZ60dhmj+S550jxznhUNjKh4JHX8g6U03Sawx7NwrEyKv
anaFzbV9+E2e/QWFJ9POCihftdlY4qJI2pG9AaFI1in6Ci1Y8u74jo+nWQ7T1ZsiKySLuglDLysW
7LN2DFgOpOLGJTYllPVg3lm/ehPx94T2OF8Y1cSdNKJJ8N1rddw2pgqnp24krGO5H5WIYM/FHlRT
/hFDlcE3hSxq/Q7JmVM0r6mgAREEK4KWfFUn+Am9P4cyUyzSDD9LuhbfklspmLYJdTEvIPFwrDeW
ad0SkCjSeUhKc7khqJk5VXYH1E1O4Y0k2t0h+NGwArqIN2MjfxIrLKJxxqK1TxKocV3DWQTB1Vre
o4NoCWDSJ+YslDt9dO/5mMynhuEFC/a7eLhm1Q653UWqy7X37irn1Z5WK10hXQF8dABKGCEbq473
F3YUmU3YdH8I7gictapXpsEaBFPi5O4EeXQp4qND9slQXefmP2a6xqZPK+G0m+ikwfHw2WNoYNZZ
IysE2+7mQE4uUgTdOZOaSnfLN+1G0h33+0VLyGhFd/1xhaud0QsmXfkrDpSsGCBaizJmRaWvGbHR
VBkaXsr93h/4t6PV7whw/yVTDbc+M9KH7dWYxxx3YYRTja9ljcFC30qAIMqXY8toieUMyMjmfHvo
Z0XE8oyJhPzVuSrDGIcveRDZ2eNA7J3qe8+7bDmN3gpKHKXGOxfMoeHKL6VN0466GhmRfrnDV9JI
youPSHThKJzXGceZRFcxg0pAi0axe0rEgaRv9svMb48hBtP6rbKD1ZrAdCkFtaXiNZ07SH+V8Mhg
Dy/oXr7YecRmWjqrdKJnoUxJmoogWEaM+mODIz2Wf1+Or1Hmzzyh1rsNqhofI+R4j17qaUE1ugn/
MwdtuhTrDamH7ymvDjmlj1KI92CXQISiUyax3g3gSVYeZ7rwct4CE77EnnhZrZzmB3ATJokUrJuF
UZRBCszQGt3eV6Feflr+6WAhMiAIb45IrxeLgRX68vt2800+fkp/VUsNFgakHpmpctLYsRr5tzWw
jYyQaCU19xKjWOKnNHoWT5Jt8MFS/+CgFNC/E1g52ObBiD8XrmWifZzOvijOWa9BEJwB4LDmq3Mj
f0ayiIc1ZTw/I/lJuDgU2lRjEbpyUKMYHp9JfBFLz8faIoe9iFvJMXf1jCti7tiFfB+HhdXNYkE4
vuSOX8v5FCtcl8mgJeMO2F+OVPhgno+PvVEpO60V4qg+6R6l66P6bnBJjAPvV2NHTtQiJG7Acp46
9yJRFRjPVw0+oZHD731fQE8R+ZrnMYCebeZV+Yb0FvKflp3U5NM6CXdxRANX4NeCOS0fCsIx0l0v
TsbXTs6n5mK0PhWlZ6SMtcGeF0mUCB6lijzYlwXb20ZlY2eHrvdukdQm4IBKQWPAoThn4MB4PzBG
gua/BuenYPfGbxuzFMJyxDCr9sp5jTtz3Gz9DCcMT3EnYcd/fmoarA92UrCy4f/kmMLk/dnfLrkx
CGMJYgeRQVCReInkF3lmdnRxXw73sPJbkKabe3e+Jn7WRQGGjDfvHUzML/3g+BVR+TmMxuU6DwH3
+pEGQasx5zzE4Txwj60GihO33ltlGAbULrEVQuvpHUM1l3t8p748p6A9JVWuNByUJo7wm5SYOgja
RVojCpDULTlRJN/3k7xMoPpSa2SvUjH5agjzii6OSkbCTrBCV7DPBM3Sg/E8ebJTcZWYfdv/WfFm
RrigtBhT/YUqQlrIMbIfd1b7Fdpvu+6zPysFdzbPJ5p0lNsMmVvZ8zM8NM1uMA5rjbY3WstH3hjL
HAIZnkVU0jKknRvVXVee4MoeQpIkBt4WyQgnIqnDKm1qaVriVLqAK6nH2Q3JzBUsCGfM9bX641GK
2J3gNCrwkqBJFX9YnOO4ZTtY0Pb8KR9IlrjD6FSxqwSbVmNk/ySU1j7cnmin6Rd+vUqCknCnKTLy
V2S2aCuYdp9IlcxQbdmg6aaIi+LT4t0LnYf6sPFC+zpNfIDi8rZI9aULWkf5mru0mQQ2cZ2fg/qq
eWBPeGZ7Gel9lVbGQ1ii37bQ1Ok2ppIv9eqyLyscY+MuAQCrQEda34Dze9+ZkPNx6mXXS5dzij+5
bqUmcTK7nr4b5D5g6BzdYt4a8kdCIcTRu+fWp7PPSKBDdUHB+JWQ4sb2bhAFEThrm64GcImaXh1r
84RrEIggYy+Nz9pUz7WI86jLK/dI/ecZbIsku/RE6E9fUEBGw5OmmdP/LfIg4sc2o/BOBWYrzHif
dERastFyGMU0A/J2zlQ8ScEhfBc2F9Q+gORakMffHwzuofQ4SGSMDtSdFyPbqAn6ZDlVmQpnBrfq
9BtXnfYlMa9DsiqNNXzp8ezieDYdqiv7PfEeakL1X7DHNwJ0nWsIDOEFhLS6BpqiGvtErTdmGlAy
LptVtOV1bTU+yyq+WfesOrPnzDcgTAR1hdhngBknthnwnLfrGlwd6bS2zEmq6uwDcIBfT32JDh9W
4oObfcnB37KVJJBrkV08s28AUod47ShHHufIG842v1UBbxoNbSs7kncYmLXPwDJW7K1d7/ZavJP+
P8gh7dbfp+uyVbfsKmJ7FJL6Glx9KGgenavzcGBY/aUzeCX/vtzFcosaxEYPkHOGJPewv1LvZbk3
BYxsmPnSSRYIKQW9eYKMGS3ijSL9Nr4uhcDEgmnhWGYaSamoTdkAsxvBSFgvx4pUfaysdQab3QF4
aXwGW72o28n0j6cqjdxViNKAZLOxjf4cK3N443zx0NAimDNEtshErGhc7XSUzjqwJigGhAXmsuil
hoqMh+RYex6FUOANKsnke9TD1RXXkn/bfaQxKZXyyPmToczJfOuHXwzN7rAal/Tj+4yqQdtowqUi
R+nlkj4mzmGZyKXxGr/gQ9KEbmxpw0XP9sbS/PSj061enLt3MwttPYX6/sPJc+VcJgkUoSFYjQ2N
1IKn4YdFLc+ykP06IlI2lCdI/SFsiS80YqvG/AacarIS130dRUGz9OSBwjOFXGn32LxMovRl/Nej
xrQ9cfSE1EeK85eYBxhnbQ4PmPZXW5luEqsENnxtjA0VyZBSC6ld0SuOzxy6u5/L9gKYQJV1jbTF
O3W9FgI4AXe8guquox+UuSNiP98vvX86I4fJfxklGDUg2ERsK0nqg8kq2iD4cxJ5I8Dm5mSM9UE8
xbY0kdocLDHG56R9HdxO3ZrELUnj+7hrUDVHF9CWtsLhanQ6DYdPkAZ7DCH3drJ0ZBkJQ1C56Vv+
IOz3vs7HDyV4T9Vjd5alHchOJUrfhMhurFhBxWQ0SAxhPQqONMaNygOqmgXK3dffPjES2K1V9oN6
X3ciO/aJCiP1FvgpRPsTlQlaDX+DD7h9a2EUrG6QJtvRoFtY57xrUzOHWpfASUYKvNGmUYldvnLt
mW34yZTMBzJicPrjkXcjVIKtksr2k4ofq/JXO5OdglFZf9KxAX5nPZ1ADezKltxDXEX1ces9HJow
ajsytmD88LjQ6jB0PAq3rrW54Qncv0Z634pU6xPpBHt7Clz4Hl2D4ok4vxar7M14s6Rkrk688WPI
IGogvoDv46eqlwIKdA4A4cboCJ4ORAO5knn82yoohVpiskwWwWmFrImqxGaVf03Gsltg38cUDi6r
0bHuDVGyIY7Ug0VzLLiH4hL5hEy9oHz5jPDeXR5zt1wnNUi0PakPKC8E8Xrb8ZzGIeZFGWPBL/xi
vVBPcdWMKSNtIW3Sxv+cqPl6QMXN7SOwznwh4wJFiacgrc0UqciALrvofTwi1MfRIA8IVkcXi/ru
rp9O70Gtb/0fY0L17DB7gTQ5831pSDcSZVEpwC6rkSV9qOTPdZeiBlD65EW1GxuLR75BURc11Ook
FByDz2Li29YjbstnhyqonrLcUt26krKU0QEcNL5tFxUWjYyX9oaLVkR/GyQ1dYceLUl8jBsg3780
FIhcZDnjnjZCsXrWFJOEf38qj9RbXn4b7TpTdxYsahSaO8T3L7tK6hoUzjPgzbAn5820jJshG0Oa
/d4lshLaO4n54p+V7VWCONQY6kyjHITUls5SdwFFDc7XadhO6tnlIwCCQpBycytcyWwSwW9Dm5bO
1uCgmOWzTZcFCMDqWVRU9rN7VNuUPESfgoV8h1sfw3dnvmsVAi9ueyb9q5IvDErJsN7x02/vT+/q
0TQjF1QbVy+sYckIXK6XrTdKtqr9+srCj0RDf5oXLV9yn7KLTnjSh73kwqPgtSlRVMOb5rWsinMG
qtpFAygkxJ9s2E1I6Gix34NEupbNwy7Fzzvzlap4wHH19+oDFEcTJRsI5PT2caw01m+EfdGXCueR
5ONy3qB6SUmcQSe/CWsR2R7G8kNUfgoO0BbxE35hmzSLxntCONz8VmuRhjpFfyd+HHqPrk/dzARE
mQq5GxVg3l2pRiPgpFZYwnUaVlWAZT5ZFSAtukim8gftZMFcfgzej7C8j7NUL7yOc9/FmMYPjati
21GJe9qAlC5qjuS4xSwWFeGBsDDMnfWRlkX5jyiPEN6ShYRWeJ5DvGBeOM237zdY/w2r+/Xorm23
vFvpAKMBTImYrfSoJZ0iRZPyKhxYd+HXnGZWpXKz3WrIEJ8ypPSyZylA6sB/EB9FLpdCu7wyZSRI
5vOyGXluy2tqHWnBp6omFmhAdq8O2g/nrUG48vMF4dafabJi9xhFBjDIpchKDXVSHGCy8HdjY/uL
TY6zNCrtGSwmJW12CDl28I9ufXY+1O7FZelldp2jO4hQXqTGMgzXGG0B4Qn/+rbS+Xfzse8tF54/
LR7cZqEQbRWThOUxvGNowqdbc4VGuU+P7u1ttUm3aIwky2HQDfVp5ZkuaXX6bJI5jfeUk2/29quW
ueCLbN/sSgWXXJ+Byg5b9SZxZlY4L9KwEU5dbD5GT1IREG8szM+xXrg6lxG05I6T/sp6l2/1LymP
YWLr9dUF4+0BtcG8dTMYfZDGpqB9Ieb0kPdbxOVt4yff2gHX0NkT5LpzPR9SeBYjSovTHqMxOk+G
nkISKUkLqyTyD4pao+cYxS+YZLtGSlE9JQvHnAj5YTHftlzfecCSNi2RVvvQmMzYAMBvKw4f1Meo
CViWP2JcrXxutq1b5Q1M7q2QH9a41Iga2xERc4rV9ROjjOSDdoAK+5jWEJnkxhzZXrSktVnWWQlK
uGGLTaICurqtlUmrAyQNj2Nq3WoiyZYOS3NkRug6jYdPoQ8GIjcPHW+UMdSMQJfqFVRSmdWqYo08
0Cwa5ZJtEwKLB7Y3u0/AfsALWFrEV6AHG9uFdI+LC+EOFMpBl08oESaV30EF5U0gvkvN+Ge13JlE
xti6PRN9JMt4prbj67Vv0XWRc3NUZF4YizpyrHJlrCYghKYO170VKdfghICo7wFrE1v5H57ZCoUj
L/uNANKNYc/DpQx0xK09q8KKQSSO9kS19efj26QoqToGtfrv8PoWJIDRxNIq0ckBiENVPaoZBZve
SHYdn/o3DNyQxG/4ijmYmZ60jgt1N6nlxocAgw6FalWqOqh6Vo55qV54gIuspbvzzeKvUCBfB42N
vo/+DttjTKZDZw8+9BisgwJm9pNfnycd0b9tK+bVLLf4YZ5IoSefCaiFdYbgUZPAVpgSh4eGMJWW
JvZ0oieB6thMJIrq3P6M+L9Pgztt6N/vtcPGNvIE9mFqBdNcJzxeJ+d8IknGLWaUQ4v2PdH/YR2G
dRManFpANdVlDVX8ctKbXGuyG+XFYE6KgmIyvzuWM0LdQQnNc6KjX61865+eazmVin9PPpctMeyu
MqUPhnwkQxpjUE5zCA59xaKbVmnXA/PpdEEUA+5S9BAeHJ6UUfBzXYdEhhUQ4qqELNduxE26hoOZ
UFa1yhOvgmAfjBEKLG/VUZEWGCiloWV7gyCTrqCAmHxMbweZp1BE5zOpfDzGIEwjgLkVx/H7GqU2
W00yxml3KhUU/U3XN94x9FvKPXz0eR2qMe+8QpGejkKdCZ4P2dyGrM3NI26BRuBFUVdbQhoWpReb
dPDdWuEr019vsaOiDCHfZI1fWk4HnQGpuux0opdYpYa+8MbPasNECqYlwYfqNYk0zNtJETiNZPA0
fQdcDemaU/PA4dMrcvyivbr9K9fTPRk5axaOJoN7ksvhic7fK02lHIr+0dicXMsP92vylsKRxMHm
pVPQljjtPwQsl5ty6BcmyS3V265nl7Vt+QabxQk1ZMfcF5j9OCq11/0g2/FPwL4cgZZk6SeieDpy
9/YtgIz5HE4w6si8zcy9JnWvEZ3M7flRf9LBodk8d4MofDXRNjdLDRTZIHqlE+bjKhncboouNeus
fbmQoemcJkBsdeL3lraH1Q0CFF5gWbiiza5r080WPiIQldEkza7j/H58mvBRt4gxdL0xhl14I30e
VOHcNUXvyotDiAX+OgoX1wnFGAaECPFKDArw3eglxXyHRxP8eNydNxF6A1Qu51vHuSM8dVqvzTwo
bUyF5CXIcGbHNWFpuUlKSbGk0npyYvafji3xozauIXhGJ9ENEG0/TMiZ5AhTvUqO2Cwj2OaDF0BA
GjgvB0mpOfqsB01/q5eRc9DRXAya0Upk4ws25pqkHfEuAG3Z0Z8lQZaHpWd1sWMjTTN8GVeh8ei7
dKmCbVhk7i7Js9Rr8ZnNh4Hs1b9z46aR1h5V8WuZC1buxTD1UfJc8skLJX4NUvbfRgOvmvdRP8NO
wED9t92CdOSx8cwZG7wjNw3QehSpVQ5LCHgBRh9AZLnsteJ1jrGZR6k4JgonpAepZcYOP6GI/E9N
3maTnBZh0NaJUxGCQ+DzNzUbFgXd3UwbKX1taxEi4t3mXA3+r2AWR+qg3IM0dKhViUeKeLqEgP8A
6ISIPY5P0JhbQkTp2EHty5ybC5a3aPht2qEsEn3jXm3+EYnyA1ZYesT0Cg7iMsRpiYN1mw4MxejH
fqOcYAgfsSfJW5XAWzyPufb63Y0m/EG8btEZ6god3QfbmW1Xvv/ResnWgii9vtjkXeVeKgUZJ4zA
dtEeGQlVWb89I/a8HpTHgudJJXE4Dw8NYUf/avJ1vOMvkp8ARJAanInQ38xGtIO60rMPegzIyJz/
uaWijll1HgE8NBXLnMlTTnDUklzwQ/hwyVinAJxH1Mu73gQlqtYnrSvebszdpFfDqd7k8YAvEvTT
n2vEIrZcJU4S4TwLvLQQSCZrWFutKU3S7yNjGxKsqqhnpqTWGrCqSCYNn8LKNqrIkoHUXiykcNY/
/ecWBXsi0tclBDF0XeH6P2WvZV2Ans9O2+20LYW6OmUul4c2hTnB7WTR5hT71gwlhZeHXH7SxBvT
dPuoIIPACkJ9DrVcsgxFDjK3WZ/GzMLQkmfK2QzehhDvs/lGPuF0BizbH+8Qd8/AgUHij2Y/PUik
LDMUYzDpjRkQVMhWOtMstdPWInST0AyByX8BSB6HF9nsw30CrO/Du3uKoC6hWzWR5sy/vuygJtIw
tTGPEt1p1y+hCkxTalK/IQatlQ+o8t3s+9pwk+nKOWr7aRbaXPIbSNyS5NRH4ByVG42xGpT+HJBV
ZqFXFrwdsub8Elf0idl+KPRUXy+/IJhNjmyHjHT50AUY3LyHTkdlkBls9vaELd6kaRH3XGOy6HWI
JNu4JfmHHINIs7o0sjPFnp4pv5Vx0es71xxpXgsLR120rnJrB4AJZfUfWVf48aCt1hxd42xbbn7l
LhKGBo4/1Iuy29xh83qxlBGkPSQJC5TkalpGXkeWBkoAKQ4aAkJqVOvjr+Y+ZiHnYn3fbArH4KN2
TRFjir+ceQ272CJ224IJef3gs9sMnsnqY1zbEpkWyWOx4F3o8lx0sufcpTgC9gP4cCWb0SaJQmb3
uY3RAnsVKyxZlxu8OxWuc3Asa+BazLzbOLRHJLJT3uZErgqf9DTogdT2TWuzwucoe3rCs3K83DzS
j0349/f01a3ZM4Tv/ogFgNuNgtQpqIGt+fMa+T9TobK1IFN+FrIAB4lZnK6D0JdvmKNiTzPRo5pU
9vRwQ1nqUu4QiflJsc5bpAOh8whee48+EDrzYs8amZy6xbFymcAvbvgB+1GyrRKZoWhb04k/II5A
JlYMl/VKf3QudTVlLt0+cuZ1eu/dkRbMf5zc2sMzQvAufUzSJ+mfJTLgk3mjspJCqR5yLbitiR1M
L23zNFX44ZqRABA1TkjriI6/YXJ6a8AKLzSIPJi0XtJ1CqJpeNNSjYhwwcqZZpCeIDLeLWQZcYAL
3w080CsyWkXkoziPIlaAXpZILFAQeSNRw6YPGckC4aQflH6VfEuMcGtTzNx23KslPBpoKrNDLEgv
YMHO6iHE53ddItjKZ3EbCeN/3XP9Ooy0N9aiilKoD7+FXoVi8pl0rjzeWFyeZQI10nrN0eQKGWrX
YcZLozKRAxdNmOryC2OOydqh8hEKex+7QR0oFyz+SYYZ6TaVoY67aAT0DDdLLp7FE5exKWV33Oaf
2Tvd5NzRzM3Os7XtWqI+SSAqOFAWOUh2QmODckCaeSmZLBS99qBeZyi+m5JswgG93KPO5CsBTGF5
HYofXxsvxFFfBqORdtkn4QbAMJflz+I36Ti8a8JaRtACi/P1MlouNLrrLbTB+f8ZpULRhWO9ecyr
AB+VTK2kiHNFhZGcaK99jYi7qqlohtw5Pl0yODaXhT7HQNfyL3TYiqFiGl5bhG70xFyU4IzXfjXt
k+HP+pOa5276W6BvJCSvYNCSYfVqllJevUyyktwGHPwFd9wvq1xUUC5WYpKeqdCZ05LUtU8UreF5
RbsfWDsQuUXU0gHv5JUDGRf3O8YbL2HSeCiYw4nnvMsJrirIRb6SmvkVC5xRqmGfazMg221bWv05
hdQGjTeHHPxjcZ/IEilUNpTEZ1bB5aLfsmCJuegNj2AW3IiAvKVJj4IJ5eC7UeyQzBx8jcvgc8ct
YkS40tIaJyc3aJPBMtJlu92g98pIpvJCqXKB6S6M4YhZT/9JmGG7c0O5TGCvjKajnynDb49buxBW
ATzDwer3c/LB+6GnDkomcaryDZK5W6s24pPvOiBDbtJ9yLjwQ5yhhpk1awUwXKxonsuAzqDa/SaH
evE6Zrw0lWM6oedj6rOwvRXHH1hZPr6NdCiupQsRg2ubl/9rJ0t22d+Lv0ZY6ziTEsVvkmjFVFRv
SETHAH6XkMAr88PZKHKlFSTJgENXSaBgUorkcAmMMKJxQALuszUMVZSdlEOCaYnuRaccGDTpd7Xa
hEncPnsxUe79jn8zXluX8JocaIXQd9CFBiJAQQalIKN8VGAnpm40uPe9L7mEGezFzPVWg/38I8ho
bSVEiUPIY0MphlbRMM6wWNYOe4x/XY6lOdlLk2yIlxzNrIchu9+PrkZ688UqgWTSUpetMV2Zq8Ww
RI4dMwh28WZBwLW8brxeGZ+Ev7+orGISgF/AkDGHnM6rYxuKw95IusNSUftb84aIxcA+wmtuit0t
79u04VcFS2Drd/QVfksPd8n7K5o4ULqQgeBQFM9l08tTAHzZ3OocerjY0NRt4zct1d4fckS7cLEv
bTsSm+wWR2C+Ux04h6EqQacOJl7y7ybPFVI/cbqurAhE9fxtnORq7AcYoTIPhiNHtj9MHXN+Jagc
QTuxMiavvPCa3sVtn6kQG13htpd3RSdHTEty4PmmPUePQleKmfnEziwDJm2wb0mKEKlbBJpaaWKu
oGDTVp8+IFbkzjorfIoBJxf1fVx93KsNzx/kPdlniyWjpacNixE4UB04/DuHRr4pEAAwTYfmokOY
Poh4cVF6gwXcjwCVJRXieVEMs+hQdPAUAlX9c3cEoab2cFcEg3uLlIiSFEIEXfCjdw872kQd7ycp
sJjfPFknFZhjOyHqJtbwk2Zly+nqU/jTZ4ZLcb3OXKrqP22hy16317tBB8bT/9JM+eWE3nCEZZO5
IYbaHoP8idJVFeLvhbVujD1ETcTs3dcUCPk9jOkrBGehDnzGynD29jIReG7vz5/MfLgfbX6LMYMp
NJum2GLZy/Kqjx+CQnmSbkwc09GiIxi7LootQcM6WOBjpTfjP1aN9Sy9BxU+6JDMaomXVwEkYJlf
vOghfNX8ufnc4PHKaQixK3r+PUNX1goasbKj004N/Ji0kFGp37347Ttd/O2GleW/sCvizf3whdQJ
OTBqXRWzVEhEbGwOtVV/jKuQIph4Dc8QDGWu4YofDeOAFWFJKm/mz9q8kpgv+DuyCem/MNYJBclj
rERU+kuMTzJoCMHVvUpqUPxSdR6OcBKKA5ypSq6B+7xq3vs/2Z+HZig9kVp4qS4aXFAJhtQdNfBR
lA+PSz7VMz+Yzu5ZRebC+0zwz9mywzkx1Y8tzb1DN5eWjZphavT+4Qk6YJb8zSGhUWwnFuLLLyYa
MnUDW3soWMfC9cBP3AF2jiBu1T0CM2C37Nvn7aj6csB9u320Q43UPF2O4mfAdhX/zYDjQCS1VbNP
xPDh/SWqGzbUCNXIdu6YWTJEuwJodNOEoO55x9zNWFQHxizWw+kT6j+5MUbTa8keDlhM10z6JbLD
KU1z5KVMZkWMs+cuzLmFM26vC1RIwplP2cCv1/ZmDikcaEUx3aPpZEEGhReplILTn/Ei0mHrycei
8zEDjZQ+gsdjPvl4+eSI1ZS9K4zPUmqduQp7iuVt4An3I8iJ2oOxyqal/n2DeN2zPyGiYUezhxjy
C8YAWuxY0UsCclShb/OKmLyjgikY6rvhRr04hl3emf8KMRyFpYFh/WNW0pxHpGN9BmaC/z/2O82j
C2MkAG9RQLJOgHHr/RYIsoLbtBB/zmyPdZe8GvlqA5Mpabci/BfeNqhIEeUwHJDinAS089U86Enm
qIhJ/UynN62qsVbrxo3ZMNbGdlD3C/7xUgLLHiEK9bsy6/22+NUO1pLOyDNG4e75cCsoaRD2o6w2
Wlm2B8AfZNOhHudC+bfnU8wKgFflrnNiWhkc+A7aCJeTQIc8fxp5a+uUGSOv0HgWQPnFryfbZ/ys
GQo4lNRIT7ykZ2ZjBTNr/fTAzhUC4U8pLC5lZhPByfFleFNIyiKlfvZQoveqMw5854S3JZ9hhubH
mX7EIztJac4xGYLIU3S5LwWDztMZlY0/IYMiKJe/B7vkW43XMHrZZ+mqUabXiFDonsGuWJznIXTY
YZdhrWAfjfNaChU3XNMnTOwjmuIY+GxBO83XRmyzLmT3etJ5fWA9bvvPYmmuqr+hpm2nzPE9nIF0
rTSKULKrXPiLViIr9NmnFuVfgOMvJpc41EVSdEcN0kbAAtJyRyR3pPMqgLqAgVz7M25ewWRb69DZ
NR9eI26CP6nrUUyekJ2lgz3BBrOnZrNkiYIS8AdMRqvMgtTRKDUqeCe7jl/T78QXDHJu9O1utA8P
viWWPvKXYNRsahBc+v8Ui5KBed905QMVqG7++PtDMOHGFFxXAoftJShi+/03yuooJtrLETl+UVze
0HwGvBQ5lCNx41Q7ASIN8HcYYfFRuNmROaV6vXAGFB/m/gJUuwJnP2IhKpXMWN0w7NmPbDObQf43
uRVAs845jggAKEeE8Zu2MiGYU498/qd10JN/vzGxUJ23CmHiHcX5W+vLp6mX9Bqkxq25zE3Xo88M
8UdSs+FQ0ybakulLNLdiTTaJ+U47V/1GOj4FaQgEkaxeE3MtcNmBqQgwH0O1kfD8I43V9u/15LqW
Kj6rfmD/Mk9QcqBzfo+P/w+SaHPBoeEJ0Q2jd+gJaNz05gz11hXAvgd/S1UQzF+cKTG57H5ktUIL
gnMpwkx6BhLGn1JZurTiNnpeAnutMx1PDXvEJd8CJSvKCtHUrH8QfhPYgme/L1079R+1l34V8Vq5
0e+4oNlDuhPKg9WoiOTPtqCtRjNTHSPO/kPaWPMQ75opz1ESp2aJne2QdHTj4UQ7lNDTqJKzbpte
HofOMf/KqJwUNtRGt9/A/dYq5Fc1kdYLPIUbMqnFh91QVglvjbtwKD5NGCIItoDldAVLCh5W5vWX
nxbRD4p8viQRuXt8iUwaHQWFjzDSDVrgbUxf/ftUCpUGQv3pya5970jPKqqBLG5mcFz4C54aqLnF
njyom30oddzlWhtOHcDK3la+yscseYOLB+CYn4W6kzYiXUPxnvyC1pVSXfLrjtAUihl70mmTPSJ9
9ecO+d+BmM9C6bbffOHA3ob5fsm2z72LjHeObKFjo3tV4OQyM2oU2sMuVbazf1C5PzHGh6RHECZe
cGlqLnsBW6L5rpIzYapqqVCt2vjxP18ShoHyeeBKoiU96LsRpw/5aUV5wR5Jf7GIYAeSvtcTvkva
dUaiwNlRiKd7SqcAfgHuRB11z9TreOphaBZzDtM2aupZllpnSMAXIkKlAFSgCMtdnXtDwrbpI1bs
Pa7NcwZ3K2VOQakdjTRESSpa+dQp5IwNBb3w5jHvMzOUrkliXkSnPH7omZL0iYaLyolQFNX4t0iA
OZC+RMJJR9dYnj4bvEB9stgA2DGRVxfLI/o4GbeSvaZsdGIgzn08dS+HbDcFaaK/XLicvMlQtu3L
1HY1AY66WUybGmp9j1l+O7nqSLExMEzeYK3RKZzueclEi3jPP0BwddebVtiHcEsg7sJ2mee845Ez
9E0mrQeyKPSjjSyrhL55XoeTR6v4tfqhQTy0G4tVheJUHFjyCTCIsXpHU12tdYQpLPr8pVSkssc6
0ngCJOXhWlsRm2zB1lIIOP8K3popaHO54VobJZmOxmskuwOelJvM7kkqu/tOQ3xk2XXqjI2AM9hx
RyzHzhRfkdCEhTl2VVEmOAOwBEIBE2M13YV9awe4s/zgKavPCAAYxW4D+LX1SDeLbLyXgyOzU7z/
hn/qOOkx1JB+OTcyDV2AbNAaGrcHqOfTqgEywmWYnB4B4qX7IruWbbIpIdzRHlfVxLfGT0inklEH
vBhwXWmzwuqqeNYAcxJGPQQZ2wMbjW7OYbY28jv2t74h9B1E6tLGLrhfKRR5JezAU5vX981kFPD3
bcQzdd82SRobCrhnrZ3WHJzASC+rJ3+ffGUEoXMayz+ttIL807I3vGKL/Mhu0QTbJFDnOqk1b1m1
8Xfu6QMoged5wUPgxEUxAaDtsAXyT/ZCK5aBmLlZup/bMQ4gCYQN/Wx0FRE1enku4KYRQQqfBfU9
Ypw4Dm7aMe6XsoHRby2cmczFRRtLbdMNgdALjs+ze48dw1++kX9alsKNfhRvRdSry497svwDEQNa
++q3UkVuL+6kbpoTTvX2uSdBM9ac1fqc9IEsuK4WWBK9EmTsRnYWGe0cNeu5/oJJ/3lLQQCCNatE
mLLYNJXCXRfH2rNMgnwkCv7CsNJTSzzqWCoL3qST6nrH/5CgELMpK9ZiTmQe4JIGLacaSAMYoAVK
ZIymLSVip5Liidqe6jgABNHnGyCTCbjGj2fv9L+nToZr6xqXzWer0MbosHUDvH6ojp5Er8dQb32I
ww7IwHB6Z42roBzX/KGU+EU2FE2uV3yJVts6yVcaThPfalMKHytNf9Pg8/IwCUvLt2nsjEuXiocO
Ul3jDNwrO0uIQFUejeRc7d4ntt0ctu7bP6V4djF1vJ+IsXWJSlQqcOXy85IVqgsQW9wRwmnjCP1Q
zQSPtuKKOvfRAa7J2jDW4WhG+pvJR3YzAsfbL2+cZeL6lqFvvuggyapjsLyXNGOTwIG8cnsGHHj+
S4LG/15DX6RV/BhyXM84mORlF6E8t4L/9/0DlGFn6/yuwVrbNg5aNYFB0iRK5aXVa3gmHUCgSHa5
te+60RTAmDR40oG/aHnWu7tvLIBr4Cw60K/wyWVy+V91IIJfxxGLgzZ5Z+OO8KXuQbcGeTBxzElp
ZlpzqfdMb//ioEHnZCXPR62bu4rTjIxT79plwlYx+9qxWc/1saZ+nRjLlahOcaaQiYp0jLAh98jM
X8D/gpVmRzmOIWGhMvzP+cEtNOk6fhVkUSrN/m5TiJc3PtdV1WC4gddKtCFae5yKGBak3mTID+mO
BjCUd7GhWtfFE0FcwJPaf6Ma0ddk5jkdJB77ePxVJ+4GANz1StG8pV7W82Avvz5Bk8KPd2aYcvUZ
d9d8re9FOpTDrnRR31qUePlVDuKC6qHd2GziFZPubCjZ4mk+QUm6qYZnF1a9qMMcr4ppwtSkaEcZ
U59NBt3WP+CbBJJKz0SymIWEd5UQNc90xl8Ek4miumnQm77MZ+kDEla0/5arGhHWoqHakmvwfnf8
o9zTPoyi0rYTZ1dD+U6xqvsqHbnaDJAP0Yyv+GmVrY+D0a2pAyORSrOyXCAKxmWCA79YcuQ8xDqe
I30p5fwztV8hHXWynZsd3qD6rEdIxMW5bVgzvvoTbCt8oIXnJf3cagIPu6GNAf9s3J9CJhLPpCZ6
J7g5CLPC8sjHfRyXVt4DE2Ls4Oct2W5bISOIzNLfCqWexg3Vt0l//4BRB+VKKYpBeooqPO3qBoWp
ULV6o2hyAjj6l3crzYojNIXbw/ykn3jfzyo9d34mvhZRSLOW62koJ71n2SfBe9jME+E8niBnfQGC
uQMt1lxtd3hhZpUapM+HtWDZjcF1jY+v1GGkn0i58irBUJ3PACP/e+tE4iXlrYNPJzbWEwf1CtEk
6DaKWowfYHU3oiomvOHo6GQvzmEudyCmwfUkPsnNULx0JIpxLI5f6cey+PJnLZSRjBeaTFPpo2AF
BL7/W89CQkc1HHTGDWAorfnJrJzwKxeIQw5e6+EiggFnA7GvGkKeu1DfddpKLNJ1RtxWQC4xDo0b
yPmjxLY1nfVgUb+5XZQGqWdevXWB/al1jJHzP6N7CMqijjK8VQ2174DW2f9KtcRABs+LCfzXE9U8
6qHGcJaNU7uvOYlWC+Z0eH968jNnAmVAKYtmLwy8JWQHLX8QvNkpGF2LNCo8ZdeeOmU9QsasGCoC
FWHIqNOn4wFIqb3SvuJNUzOzzSU10Df8lSCkdGVgfqh5VHDanewRvpVRYco94CEgieDs9entpkop
9HkXu3f1woq7PsSEN23uytRE/N3EDvySxrpdprSKQv6PnhBh35BFdfEz4McJiB7ua21YmeI6O8X2
O9vrfGMD3hB58m6rv7qAOX7qL/NUX9zI/EmSIcTGdd9MpkFBD5HtT/gAUDMDr4dSIAr1ZMar7TSF
AYyhYMf5RwLdd7PUxobm2CU3jKgVIuf2aYkSdApSDmaxcPU5AAGKXuWq8Z2SXUjSmm50upyq+eY/
hzZCk3fwr2i950X0WQfpEezPYvvOifdY6zmpA+ggMXjWqiGNwxOmogJeZ3EHwiA3sEGycv4mJsU7
/ZsLybfLoHuf7+uO/235nKxP2mCZHA==
`protect end_protected
