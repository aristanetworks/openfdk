--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
cKNBlPjiCrFnCvOhXd/45g2EKmXj24X89BDDyo2GiG+gd+H/LfCA/Sp2hhdEMUJYKl7A7VypYe4o
PCzcgFs+a8/jWLfBF/6Tlxo9lup3Nf/0ez7VnvHXShfOx7fXLUeQc8P7FasPHi3Fcko70YKTiXXa
mBtUyH+j8Vi6/ThUoB9xwzNTP/K5JlnypDdsHpQUfFFDVY+G1rlaDuOUVEORUjPjEonH2I+mMga8
Xo7fIK0NQocFDKGM2NVlbIUVSoCCh/Wxhzr0sYifTPGhoR/zggD9Lc7WWLON7sgDZBKv1AdGX/+F
aV+BnzOUTqPimSVNTOKjalPSoZestgtvVegHuw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Mv+Mc6N/94xgkMY6/40QS5AwuM2GUh1jIsKl1ScRCKA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
B8bwSSfDLiFccM1glNJxjO0xxwRj9kfaUIW3ddo2kIve0g7Ugo1ZIID7CyuqfPeUTZxuS0Vzdu/o
Vjm3geQVr0UK70PvlEZ9pLeT98unzqV1BfExzXsDqnLN/q7hIYtCLCzGAD4Km+xawO8yrcd7ubCe
2jXxsu/byDvDR03oyqU3UsssxjvaEG6CAoBSLfB686XJaDbYLgK09XuSPtQRhl5VRsL3v2dT7CI9
HusqkawCYqXi2SMHnWkjI8pchZKXAIWbGPPJpnZuA9420TYhwGuTjNWp0d3BQvO2HAKyZwq+8dn7
Y+R5/Ac+hkM7rRi0FZ+QXnIblbJB5MwmB1iuhg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="y4YDFc2+u3SC/A0RvypYR2c75Mi9Zdkt85LxzEsdzpQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33904)
`protect data_block
/ZfRLaNjYxB3lBbRiCwdijKZa/6x7ddGiZrE2y+IsluUwGJr1XeEFvup2V8ZL6pq7uqqYezpEUc5
+CL7i2MeIj0MZAnCHXbw7iKNSQCb3kntCYDl5V8RlFCH6diP0St6gFnWHqJwvIpueoTf/KgCMjK6
mhS+zcvjPD5NP92hHqfme5PEWdKrfMov8rj3brtJA6rwHGKNbDD+9zmpCzvSc05JylmOK7WSvNTk
77ruCEvSLss1vkVaZeBGAhHvUwbNkZk5uPta4LUXG2KEmHBz6CkUXAcvCGS1qd3FfuF2UfMHd2wW
XPc+8UH1zHzLPEDDfaYTyNgpeMwF5Bu5fnLGVUtVOHt5gMBU/ial3ujsHmfhbYVp2iSG3yj2v7kv
pr7d45g5akNk2ZM0JVQgmDDgXqMFU/u5RVIlBw84lJxkSdwh/80aEpWIIbtDDc6vhiIkekIDbEPN
W/M46lUTPlkuVixfotMv4mx8m35pMsKDo/9IezVcH4iLywv9rPRwIUiYQkJP32gDSMHrkwfnSaV0
kzbonDv8nDtc/lwG3R/+KPTbiczTFm2g2Duo8IFcQrLg6GEB2zUVIvWrz589bET2ZsFBtQG4dlmc
vN83IcnTKf3ym/XZSBtdnL4cHsmrFU5PEEYn2bH7nTMmC+zG9Rt9jwXCmAYWavPo5YV+F2Gs6qbE
AF3Zh27AoRiPNgeCGFXypPe/66uwpanRV280KeHcefDbYm36WlYip9BtOVVowM9fOrhtCnfvdaUX
D6aqOnhX2qsEyn3OaC91j4Gy618lUxcTuj6Hz2Vv7C9cmJn+TAlTc0gCjMfS1VHD9k5biEbwX24m
jq5c88OLcyTvcEcklrY9rJgdllQwnBhcZmjz3vtHa/OTrydr+ZgaM8bxYrUeE9dgNFn9xMLua649
W/KzTgMVIxbuw8C9Z7/YGDmRM9h8fD3JV2l52ADjNFs6HuUXXW1p6h2caOhAxx3flM5ygHLA3MiQ
KM1DDrANS14YokQtA+U823f4zqeAJPHCUDjdduyzI27VvgMsZVZc6M0KeY8g22bb5lKxkeSiKIeF
ZSRkbRdib+V7fenNg5LJWvCaD/sqTA6NO8Fv0keJS0Ls/vfeNhOuOVNj7nzu4u6SsbsWPaI8mwDe
RVwV3Bagz1BFb6mtrOuQpa+fCLQ5CMz4nfRWH0DTb1N6WVu03r+4pYKVVILGrokWP9Z98tyIASXM
Ku663y3rcuGSOezL/YLezZiS1Dfj+xPWOSUeEnHIMnxlCkfeRGq1qOdpHLvufBKZju6xl3SKfGLZ
8v/PWHmqpWHZ+13Hm1GX6TDFiaViuTrbO3m442ANYhH5FQc5C0svzq7p8aJBnPow1/+ypMdENo5G
Qca8onbCJtHuQBluWrHgTZH0H0Lk9uTZY5VJeU3V+0rSzk+iJ8Sjwjrm0i/D2L6rSriwY4F2FjDX
ft89Rz5nkMLsM5IbKNlNVj6c1EBSabJYmv2Bz3XTlOyx/+ayBVjodSRraNfO28+sRvxMIzArk50x
3HAIpXm8C4Rj/7VecQMP0tYdfONBsufhUsN8u97zf7syr66igFhUnhQ8QPCE2+T38TuXf73a6PKX
7wcZO24rs2uyRNW63UlO3OaJOmxSjg3z5wuppMbzRxNHWNco+bwwdBWxMrxgIuXdER0RaZZnYho/
RP7fbHusjo4c2INgW/Qqg4gvkBcLmwXbcnH9rVoUdt7VRMHXWMnNNIJus1C4TgOnFGhXJ8MWby1Y
87fGaC2Qy/01vb88adADyY6FXcCup3WKMnM2fAPNt++PDKfkNu7b0sCvQrDnGbRDXNMR0WIQIrDx
Ki1+/WKliePG5MljEkvR9XXT9rM5ZCE11L0P3AZCKivCNQdI7m8abUcqzY9o4bQH4ACbqeWFz3UP
ZfzY6ZbXG0lgJ8qY5Qvrz6/PaEQB2zZfDqds/s8BQxmKrWbQtm9dXxZ5CuH0ExYLE4Num9qu/Let
M4TsU9vNsyazVG9ej3kDzaFotDwFuNbENMAMsAjpdBvSyCCPO8OQq33hQ6ZkEhX56olMBdq8+AGP
P6wSw0E60vgPlh8agZKEJbhxcVnrh7jgoaB8QfvXxyVzZUp/4tVYWOGaioRw71mpmKr6Evwmf0e7
zVUFGDEdIuffGRYRozQ1Vl0nRKdj7br0VYfBn5z/92fpXZe8HEeHeJAOEh0huC/JzskknrQYctit
5O10b8DwpZzqj4Jfgbn4OXzjyBFtvxxH9+qoG5Zb/rHhVuhD0ZebyNlHn1FVVSmhyZX1Z6eCuBRC
iJIJkz6XDbNNmmk24TcHRDzBvLE3WB+ZeMDR3i1aukWSkTcLUVhLfq8lG2YxP3EospVGkimCod0k
Tq9aZ0LGd0JIfaubsjydHlYiLYiV2oeR5UiT1deFcFdmzAv+EZYorir8zx5Uia3Ahu73kXeBlL8G
Y9NGa5ruyKZJ6kdQE79wz1E713lYAKqUuBFjupJBQqZ6PeFRhwS7iURI5D1/XvUkMGqu1NNO2HTx
qaSSlN0M29hGN/mPsiTVRivBQqxiXaBOI0Bnih3hdqpFrIKFlty8Orj/2gYMlbBEGo7RSPMHdyqr
OrX4Nia2xI5Yo92jwqZxJmqzrWS+qILiP19eMa4K8k9eGn8P3L1H7OM5Tb4luqnm/zSSQsOoKIQJ
lWL7yQ6E5ZyTKFKhwP8qh/2n8w1HuY5M8zla4MjYr/0tWQ1S6ZRS40GzhuYLJEf8B92NJj4kFaTz
W2K4aJbosh7nz/ZT0QexpJ9E8+wICytM9+c0qDt77X3O9TbrZAw15BRkBtJ6Fv8hXT2lwHrYu56S
F1XyIwdpRK3PpsMy63Rb0BmAVLOObbZHLvvY3ootDfGHNjbmw6Vh1hzFJrzpbwyUOnToZXCYUwHs
8cJXddoxqsRH2DxtIvQAUZ4lCTs04n80TmYk2ewNc8bXHrajBmKplc+/U5OC1PyPm9I8biu+mcpd
lZreKayrMzA6TwthvRDvFB9KAJHvSbxtLEF5gi3v5UE5RhosMdGCmnxxO+ICAO925NeXWUfJz6CC
FwBYa86H/TZNFgnwVfUQw5E5jllRMpinaKn6QvJ2RnQYPfq7SuMFPtx9wlggavO2fia+Y+NsqJ3P
QUdZRVXSxfU3F/cfve0uPnblWn9aRTO4U5Mp6wec+P7rg6Ys2vQ8XyGOf666G5ymTKKh3tB8FfLz
EYKesTQUrlQyAluxQpxDXPQfiJ2xnGz3+DidA2kx2zwJOzHuIsAlyiB/zfEWUodyW82WeC5zHw7I
cHoHRkcesebD9O3VGcj5IHsu2APWideS88EuqHD37fHq0Xx0FwKKySvMh3FsJsqdkyShNBSCxzLZ
cfS+yMBMs8MnNzkdEzeMINucf/6936JMDW65fp1C4U6dxXlfaXNHTSJFNUWJkNmymjqvMJlsUHQL
QKnZVQ/T2upo8zJVLTld4g0TyxrOz/NhLKhzHOkt1ue1QFSvsL4E7ht4cSVQecGnbeAScwZq6n4L
L4pl0Wb1HIAljFzFFLQczdW0npbFzRdZMbcySP+75KF05uoH+VHDzSMOvCkVZ9N3MMyvyymgrfFs
b9meNZ7B8svV8ZVbU/Sxi8vob/tNeD68cOpgF2HG9knx1zS2UVVXmPvC38thmOywbShO3vYLVfeV
nKbpTjLIOb6VDmvFAisJ6820zxwQmzx518stVDvXLI9GjZQ3FaoIqYB7U1+yHzCawEnqlYO5uNId
i8xXTgcTrkk+UeR+z/lbKK8levbtPeS4ubwXNIy5yHfxD4cLNUboV8A71/oUSgUOBs4TyNdWMPTA
mbXRl/AsdPj83WdDj2hkfl2HGuPHfgqJDCuLwGI7vTjCgyj7ikRD4Pcu40Ax6Zfr2vKgLo//fYM1
uGdWGL53tqj7fh4BlKvdiNHlQocGOxfYD6s8UlCsEdxTwUVuwgOwi96JunHeshFPqAIaWUAbX3ME
3MFzw3W7M5Jj1iWl4Scns1pREs+cKWrQWUlMs3UffFuc0ZkFBfB9+3HrdHpfZiXg3E8mLpomXdN0
SEaQmFKWi4rZrmNtcS8+AknR6H1JwXFWKV/9Ab7Q+Ko4nmCwfDJdeAJiMBXLPlk75YftM0MJwM77
sEd0VKmz6mgSp4Dkh0wwti9uW4b+zIh/S4neccjKtvTqLUmz5xkom6Vb2pAEM/M2pam+eBC8g3ar
wcztIovnTlvNQlapbjly8uWgA2hpocSExHVhMNoDtyURAjGyFKWYH0b1KzCrZkCjVeqM22UdkUKE
CRAaQmdXv06vlcRHnK0bN2sDwWDAvbV89LZvjC6owsxBhQaNpMPalM8TuYovlZkpNo3ro5n/RQSm
4p07O6kzkdHzm52aEJwU+2tHWxAe0XY44oHvPbg8drlCL1W9ryeg62odXu7vcqj+LpI8niUWYzZY
Ad1Spzq36pDva4GBf5au9LC1+6P7/4CKxEZy1FO1U3i37EAMSr+wLCR579t0htyeay7Tmx+n9alf
JKsak8fSNHaCxInHeBmgPXExvLZzIKXjHFIEMlfMf3CQ9CO8NrILiXYTxkmagAMrDCJ6RdIPDQPo
hjjUlBnr5Ll4LDYW7PsTpHZaa8eETvojOU+g/3ybwpcCL58YRCbBkmLtZQYxL8Be4dGmRT9a8nLL
/FxHV6/p03JmlJ2KjioaptNeCzsRRIxA3tu9skRhaaQBuGatujmDvbnUkt6Rpy273SP7mYR8ncy2
rxNsmGOjR62izgwH0MAw2Bn/WorjajSi0AJq/05VwoeXPqBkSDdv9pmVnuavRIRiLim13+qkTWi/
vBbEKKHir+T7ibGuP+A34GHFZsfSIaxFZ1zk0vVdrEp1Tv0ghUmfeQFkA6DL4tYwM4AvWrbYDgXM
a84gfGHZhyS5ARDHmGNSR3MaQCcdHYZ7VE397YyWSp8cHV/JRq+jakhcx5P8j+Ju0Ty91VaOY3EH
m9i+YqwgrMHBqufGJGyqvKEO3v1jXNpJqPgZey8DcdZLa5JSjs0qnng1OSUKQCL/vLPrmzI9FXBW
F18rdmV5en3qbnwsmawHYRW9vQBp7MUBngO16RSejlPhY/ebMG2sFyGq/5WPxvZIf7kagpijEO2S
v1Iew81n5t6XGOVLMEsDuYRMHLXPwdRLCWO9sVGO47CwovrtiRsHoYL3y/r2sDmo1ZMJf7QOkMxb
jbMQbe/ZHOo5QXdDN3jt773uSH7e4CI1yYBbJQgeFyNMwbWhlf59k1LOfFL5Wa4bkPpMCx9+sTiO
Xy1+36a1PrRdLVIfTAfpbMt4bWY5u+0efcpt8ZypX3EM/Q1b1mBsHruAhLXg3HlDVlsfkydC3Dsu
2jI0DiWt+m7p3qKqDMsAhv476SYzjIH3wRyOJGZYPbAgYFwDiWCL8011CKqAgL5gAKX7ckdMl2x4
2NzzT7HIWuyReJ8IjTQxSvVxIl3Mr10WINl9bzI24bOP5zw2dR+iN4rDCthhKf1+DDULJBjF/fJY
kBrzDyBVjVdElRjXC8gzEO6GpAFmhgKUrv5JG7GOUI937/PdKpHnac/9M2QjnY1SuXpgSMbwZRoZ
7VtcY4WA1sK2WJ4Su3HzXWu4tmFx6rPyWf7v5Bzv5L0wIoYLjOt4J41gFrF/QrCobHpsCc0yvyaD
kAxpd2yMrFCdrD1cV0ZkTu0Dro6PZZaOTBKNIGi5oOG2kd9ncGxH0chVzCEjo5ZI1rXk+DL7Gg04
nlDbDA0mBP6b19g8ypK7rFJEzk1sa6Zg+44GLXJH3quGV+xcpmz3/3fCPKFoEKg7dDcP2lJkOOAX
mwLCsbIcrmvHf7oYDwa3zawIRD3y8VG1cBHwc7o9OdeeoCdjkKf7Kz+4n1VHUJgyKlxsAeQK+dhq
9esfTb8u0Z6Ed1Qg9FG7MdY4qFi9yKldMWXso8VTHS7+45aCE30UXaiZb+BqWU2P3AWYEo8gPrfg
abCH5X6I1Mn0gorQp5AZWTsozfde7rVdeIYGbLI5WefLM6CSNNs8FLiDSd3eL1qcG44qapRPFDLo
aSfVEyu2dKZ3bVfAYzKmP8FxGrIgpQt+J32oAmOjs5b97sQqH8cXbfPSt+6sJyMJLITZGO3d394m
2rczFaixU7J5UPPU8o9N6lCzJ3bwZTUuRhcOhDKIb018yQSoXmEJsjmFft0fwxE/9/8e7bbc65Ec
r/eFuWOdfsFRviodWKX2TmLAx6c93nd/pwM+XirIAtA7I0+EWCYycnIYuYnJq58bLS2eo6cLIXg0
7id9EAlCTXfmejbDIZN/muJKTit0V2U2KYBrhTwrOsg6lzUMb+ExeMOkcHF+0WiPM7SaAW/H8/HF
1spI6ApDb1+CbmQx/kqh0K8Qcel4wW37ACjg0aRrHyjlQ17NydYUmtzWIkNu+d5VGqL/6R+Q+4BM
SaJtS23gtKSpYGNC01GW+GeMeAyw5BKdZY6CyF1tWF1VGHoKxmi2CvX4oxguueSh0vw4svQGKby1
hb5viYuizfETHc+5LV1AU/Tb5xEroDfJ4qwGWanV7NC6cwPW8007UuA4canrh6GBKVtPQtyohaJ7
n7E+dcXKMmFlSLKjVKWP42qxGw+5dcXJXR/uLrrR+/8e22OLGj8uB9ivLqTu5YsyWzxUu9FyFirz
RWrrpl2QXJx/wUHW9sOFXBqj8PokC6WcyM/uoaOYo+LWwqnyhzjaO/pFgV77yKr28gcEl/wvRobI
Y76gIgL34b3J7nYXN6g1Rff74lUAEkd+UTC0BMOa4Juat0FhZh7H3Rv9dF+oR0T2BlSICO1/Nw30
xKCeofg2G/0C2EI2vj3kYkLIQVo11oXmUdaSI8qDO2Yct34v3IK0aW1/E5zQT3rAB4STWlo8aa45
3HVq+UWVZEkVO3LKzfaeuApRu19peC6uYeIrak2l0aI+W63anuz4QScsBUeGhKtor8vvogHKmCYg
SudIHq4ubrHg8JLahSl5xE/ieSCzaOaBa2t2iAPb1oHnjQ8ukkEtoomRfOajKlk/zQp9uGQ3kWr9
3WNB/oxROexG+oj5KbapKnBePsUIA9lC4eW8qRPqCnoEVlC3qSgcHGmCs1AvbbLcLWGVzNERDgkk
GAUdLiH5NNEk+ZRyZ8lkzClGo/lIOFtsSjoTBfqxSDiuaVkQLuF50zlpfPncMkSulLP6Tx1y+Yvr
+EAeieYiR+AI8Yu/9rcrDMAfYH0MojF0xmfOBuP9n+Q3yQUrvPjVcmqZBF6DfkwrY3GhlhWcLpAC
UXv10iNy5LGCKCshUkpOaTDvl+E6snqk8HM+2W5YnfwuJuQxlu15xm0DZWOakoCSU+bN/TGIAkkg
ymHJxVEA8AsqEH92oBTNqbhtLGTkAOPR1mXvlxVVXGDNfd2p/Z8hTBMuYt7PIIii3QfrfVnxbmst
wZ9qlDK6pPb0cG/FrH7xOdGiKVoVOdwT3AghmtQAHLFJe7/TgBZPzEhQU+IGLjmHCF3grBQyVQE9
bfoanEXmcvY7JVqv+wCMnzC5l3qe0OSijSAbv/LL5nss5x1rucWHU8Vez+JgkMmUCoXhPXAipXb9
3i/xdMMKrnKdimNLne2kQTVsZz2/9B3TWXK0gb6ApsC0nbh2ybha/m3XgxN5oKGRDvXdBjQwPMmJ
bYwEB1KVZY8Styq584dx/Ec0GKRaSCPl3OcsmJIlQRVhYd0WfvOCSJD/mUkiG762oF4ss1DJ40Gz
7Rok6BzVIMuytuR/fK65ZrugJPa0eFmHUSCx22MGUYPloaiYQjKrpsGeliJo8hAGRIix3GwFiIt7
5kaNWWYZZTgW3Io6aw0da1Wtm8MH0v4k63i2WCX/aBLnjQk7phS2E29UYQBFhcdolvvzwpBCIB4R
sVOD+vok7EBHdHZrscnTplOXv12DZ2+N/7TcLopCPGNgDPNohQBPKf2n1dTcOX9mAVaJlxa9zfYp
ZD7ZsuJkcZrwibe2cI+uDiCnhDn6MzocKWCOsWFTIgWKXNkHTOhkLnuq2KBrxC9y5uD8IYT+2SBA
BtgxHpzgxGnyAhp36rf5e3io/2oEXUqL7qaw26hJuIXV6nKjC3i0uf78GmSvt1iHRGe5+VvTR4m5
RIgS+NaH0pyONvIyYNAnuV2DfFqdlfNlOfxxooi1tt2ZHpvyhLi3zSdSdRGZ/oqTBbacc6/l8kks
UTQcdvhlJsWEE6Ux8fV3aiQ2evByEAKriFU4pU98BzDi/LARkGVQMqeMxjWzQksy65sAzzOvelgH
npz6DVXeefs3svIpk2LShVdgzo7xS6edsHWmADWbZMY8hn+qhxVLyEVx6EYkyKEy//nwRMF9t7jH
9xkqYWqce4oQSXWqcxMk3hSQFDwXPjro8OmPh2VOVL5RYK+csQljEVnIlaU/vOVcnX0vbRkW9B+a
m3OvlqH1puFyYGAmXqzqs0kv4k0nKaN6vDcmiqRBQ9NOTGUHmgPmIW/4vWv46cW8x8rsl9wNdeFC
aEGBftcmL5aFjNvTIuD0NR4fTMO3Ww+yTPdhBDQmX3rQZXy7UBfk9fGhV//17HZB93TVQ7r1iyOE
IF/GzrydKJh8VOCvrV2aZXfMNKTyoLEWAy9zQvRybiXiYsUDC5oeNHk37c0Nr2fgIK1xgVe5gAeD
kMeL5Bg8qGt/7FnPXalaVAXk9WesSn7WRP5N7AlrIGZ1yttrxDTN1gA9U64b9A9hwgZyndQS76iW
7RF03OJX8uaWD0o5/rHLY8evtRe2hADAlv07DDAPWyI8ws7/2O4OV95Cu3eWQYsRQFi3Gn1u/6N4
PnbxdLo30xwV3HEPWnKbmI/izUwENTawozAN6td+sg7EUn+u+n6zdBmJj8pBk5oI1EAhblUDSEPs
wWdzw9n3nAlkQFJVLKnx+A2+PmpQRmLLweNbsMweDGpaHrTetix3hv3iXK/h7Tjwa/iBCOw+UlsR
lziFQyoVWbiwCwhSMo4l7R6fqEXkqiVmVGbeyfyB7ioSzy8MdC6a92AQgb/ncaaOyKeYnJfgai3i
FZG91whUpb3zWgDi5ptjnZPuBRmpO4q7RbAolioV/bxnMlfanskp5b4zSbL4dg5ZSjVoFGHQMIXX
Gaf/uS6tKz6EaS/DeyVNl179f/esKVaUf8QSqOQ1s8yKjaza+sL4blHgzOttHfzjp7sM9qe3cZyi
C4U9YB6FpLdiAPZhwx0vVLBwQ4R3IR4yTSo3XGlIa4XOtZYFoO2DneF7k5LTjr3U3xlSFvnWDwdW
932rLLpfABbcL2zUlP1vjC82tMjqCElpXDzF+VfAb0FPE3eI8AH4Fc3o7mCdmEaOis7fx0euEjkP
LpfZ5zJpXWQrClov/gbSwAc3SVrCiEUwG/6KiL+7aH4KDYNTZAuzfHxGiwJgciHW6fJDi9xQTE4j
kMmXD6uFhsLDd2hW3rhOGqoGUVTkWP56rBs1t4sfA8tRk8RKpDbp0+ho1uggXNIpc6G/EpTuQwVQ
SaOyYXoRscJ2QLWMGrTD6zIh8YonyjMQezKG+cImOpCJuJZBWU71tMBhm9jUce32Ev0X8A6RjQZC
kP4VfCWszK27hX3wuYnQXn982pY1Y9S9+tMqTGZ2wcUFQA9NtYtXqEcLAyJfpeyd3KuBAsLTe5b2
FGGLfcbQNFoEPYWSCNcDHV+zfkfxjcerBB7as6WR0jQxD9hFxgyqyOjqFLTaWVQmxSxZFk4g2dwj
aUxpdoEmfJmRY/c/FYi1lZR0WIvv7Pjfpz8yEm6PGSipfpxRxDsyvRRJhG+ky8joy+I7k8I9ILm5
eUx14B/LJHPtkaQHaFPWXLxdEnbTRL/u1COWqsetQrossWSkdUmTxdp06hhOKSbEJOfbdLzkRgWk
OTXy6gkGVkQNU0ZZg/mQzaT8q4KqdQUD4wWbRwUY1aRnobFDnmMDTvXdlneUE4kVzjbI0rCTGtUw
Q/yKnRh9/XIafE1/GB9pKDWu/cVS/t6xvJcloAPwu1BWTej2a2KKRCKNHhiJSu8OONeyG5PZoFo4
r6K6iT43LXnDhLxRqyYt/8FMdtRAnLxkKecNXywwFnKOv6sqjquCF3j3ht03ih7ZWxHVcGXdUc+E
2KPqmv+wc5qEdXRKph+X0KNfg1oXXvDCjIICn7e/qU5E/ORwsR/IxVEMBU0yAW1s1DcSi3VyUXy3
T5yxYsPTdidluQ7rwuDsohvuQOPcFyJ7eavjmVw2QqJXa+FVKmfZnlWp1/D+HOyUQTEHG6oB0o1Z
d0kEHeWqWDVtl77+nF8AF0MMh51+oDt9Znq6kem/PWixx6v1l5qqJM1x4twKPF3y83iVhSiXX9c2
bbTMHUcuSKf8zKQRGC+GH7I7IFvEcmThN0Xtwzy80ei+nwsS2LLimlOhS521J6t9W6y6K2+i8EWw
BWMo1E2A+u2BvcLHdvjDiUHahznaLsntzMF8z8YSTCGIy+iBDemxwnv+L0hN2egHWwWeD0zvuUyz
64YnzP9hnFsHOTXpndS2thli7yBuS0a9u5ejFz9mTiChh9EBxLVpynU1byoSxn004bWwvLXvRfSG
m1kgXvhI6UsL4/NrTm7uApye8juJ/aGbpxXdp/Y38VEIfOYpW8TfRmfoavu21vfrXWqcIP63X/Eq
8Q8jQcIYO27tL9ZKk/tkiGxcOqverzicD/v1/7UVUn9VqjBqdNd5e3oLCgX49SFVrmGsqsX7A1VU
6NpEt15GyBNAnMZMadOKv049ZZfElTnFS/lQyhdRsxHA1sYSfVDwxIcB/TCQ14qrHPtLPNH102Sl
cZhwzbwutA9bS0m+khK8Q0zCer1h4o0PVyFjLSCyojVIxu1XJ9Q6J4qP8GR7KWDeBNg1d69gzB33
jTWeS9I4SRB5uTL+p4o4yx8tnj0wedyHt0crPMUqPXUsdtspY1fKuYsqxPGscM8Miv+/T3xSvkVh
N9jcLEBSQlCvPAOefP8Q7ij2HiKdi163YccRwUt5fLYJXED1FWdj4xaMXeELJd1i+OG+Yh3A6B04
HeGZKdxH4dIM+0wXGHF6hNG7+Vs+wyraNlaqbGOyGo4GoJCukRvfZoOumTUAv+H0O8ofKeLLF/bX
+N1hC4sbHW6FcnkTWQoYUBlILr7fOdufWUtmpadlZn3/Bs8WK4EXWRnaWEbWaLG3N+NBtBFTFuql
REAVf2fehJN+pxlHwMYt9+Pcknvbobdp+Zi1qqGxcxp0QIASsNXlTvn4ityZkacOwSll6cHD/GGn
XZTHGVAf7IhQfmoyqce2Fh02SK7iMTjajp7j+Od5cY+/BQmmV+ibWBAbpPKGqd6xi02jdhdPuEXo
D3yMbCC6ek1h8BYyl03tj+TK/AWaoj9uWzOr8BDxER2f/R2HMLSRlsEYG2b9TmxtAH4SzH3uPMh6
fI7B9dIS1pl2LWx+eoG7z8ArqVmAxEEXP8z3WtrinOd7c/nu4z2e9NnJB7zkeuhe/7SB5eRrk6NT
SPVqEpaCkgcsUdNYofeIQAD3PAa3SJQt7u9GxNerciHiC2rzFCsracMjn3B6NHfWr6OwSrmWe7/G
jdk/6PTD1jJQgh8kZF6SVh160ihUeJ48YIF/8Q88kb05UFhurdaUGXc6c8LRIZclMhMwKFDmkNsL
X+rR5AL1WvB13P94p3hn+OfWHlqanV1aHzQMlRP5dpByGBY2QQ1VD4wu8mmQYXTA2eJjadYh20YO
qPGEWM75nwFVtOykrDwRCHiMnLUap+Z4tGFQ/RE8ushwy031egkccGl1mHbX8msl0gpZvcWVqW4b
Z2ydlgNCgc02kRljMiDoK60LtPWjMFJap/ghGO/Xg3zhI+RYwK+iKPokw/t0ZV9SuVfQ8LUw6W2k
11Hu3uxRWutD10EHyhvEq6SE2xCheW/4vcDydR61VR8MV2n6646ADQL1Ftv3FFQObzXD48z8vZ+D
5Qtv86cwj4WH/yhUk+0ILT9A90Hn+9Ssp7rpG82mhF7nXFBwYdEtm3tqP1/x8SSAa8DBq+IEY43b
/F9XVKib9tLuPRKmgqnZHqFTgkOJR2D7JOh8lRkogv6Igi/IbwVS67xmXrIN6A32DDzBmsSe8BAJ
3In5GMSNcbDiYv2rGbJGQuvac9rxr0xSOWSG2FFnsrC1spBFZVokSbiJQjABzrbV5XM8dPGGlPxQ
ztiQLwTsVs8fTLgZ/cYKkUMiSDp/5btw+z4x3W7iU+agbHeVYNRY/NK3FZiH/gKD1S1tHLjzb5Lj
koPoeObysP8nD/OFKCY88Uecw3cPVujdzUYQl83rCfkb0RnC7/dTSYQTbihjofACh4a9f7PSUDMI
ZTrAx3k48PZW2l50L+HJQnhPc8vmYRBlMlFpzStz/tAFtGthptZSsd0Hh7iOJv/kZCvuVtWkS4fZ
KDEFkw6l3Gox1yhPIzwAbviYCwTW5EwpsnZ5iao3SEJ8DCcyOnKPYo45szj+WvHKfAc9cPHxUNHq
hC76J98gGDUwGKYstzNihxo9z5q1QEI7bc7oStU1jSkaKvlK6IV/SXO+8HOkuUAQCbS7hLI1FfFh
2Cg9mYm4sM74gUUcNqdzq4lb1JGySKfPaorFtQeq32ZWO3nIojZkZwU33aFMFgSk9RTniPoRglRb
CGcahQvtGgeOvxbU173EoFmJp/mezvX35bWlDOh5ZFgc3Hd/8G2VKSQk0Cyshhn6oQDHXveydiWk
7afLHPRtQBxuNM1qC9lYMCPucwSjk1XXZJSlphskEY/O8XqqG1X/k8f1uKW3IKAJo76+DDL5Y5C+
tkfO9qixg3W3HhzTrUFHiQmfptvVz74dInryzSNzYuh5ttFNrrGTIVkkWQwQc+dIFjcvRlZVuQ0z
4PLpAyMi17Q6PzS7gtNEoRU+Dg0E2jIukhAqTRP6k2OSoaVQEesvkv2jNwnnY499vugrVVl2wxUX
EIlyzy6rDKjKjOxVtUdmp7jS6wpb4AJWYDrK3gJLNolnmOk7cI8IBnKIYFdadUfLYqF1pQqDNzWh
BS8WjlHlQ1HpAW5YKIsgjQpLmxHNegza0tmElFAVBoM1WOpQOMgVE7CTH5k+VEzWzXhiOBgVISEm
1L9A006OnxDyjzVVklIng5rSpyWqMKPU/3I0IUFOm3FkmyTopsKuz2YBWtmK0fCL2F/GFJkr8q+x
3qjsbCMkHjtOcyfpT4GcykypoO/CfMssZK0jZ2L5udkpL0H7IJ6Xm1un0+XQ+FQgXKFv1cct5AA8
273B6kktSUdV2TZZRnOMd2aSxmXFkqX6lx9HU039kAh0qVwURogImK1FUTzuPAiby3ZcL7gAMLWN
CvgkfNkFx8vyDLQFxFjyyGnP93YzdDAhoFco6poDLL6t1WxNiv2mAW4U8/fE/F8PUEEVjq2M2QyZ
24ac4BHNeeObaJJarZNNonYOeuEu9ymJjGAAgf5j5Lsbi8fLCDrfGLqHETv+brCOTNch1zILAg6a
nhSahxgQpJrJ07Xk/cjOv1zV442vHDo0iQHqtE0IbfajiYG+ZepIDuMWM7DfM55IHIeFSjpBmznh
Cul0I7JXtWbYCCMtgytKi31rMQjAdN0r29v2ejhc8Cup7ojwomizMFs7yUbM/6Vs8ioynS2/vXwq
TENpSnCwzCw0rCchjqxL6ybCnNJ9yBWMesaRqbbDZZKkeW5GoZBw5leToXua9cpl8wmrDg24D9fA
bN9p0XpflRetG0VNc4Nt2HrCi0RZNlTjN0PyTjgbE9nB+kxQcChcfhVvHvIbDdVuh2lQ0HSID9wP
fAxs1KRa07jftPFlJAlx8ITUnfkt4tRosMhCStHLNvu04DQWzdl6+O0ls0MstbwApw3872kHtsyv
vAEyNdGhB9WqkMHWIxcJgNRySn+A7pDD7Z8Q7CyPkTlrdKD4r/wux8kEqhLjH99t1mKdvVLR2Yk8
tJhoCYRe4FGnGeI7nC3KksgbW2aUr8yJA2bC/ttEr4sAGZW3O5JD1YCoKInUDGhEonxfYRzMRkW9
wIVytEkPS709JHkt0qYOHIoWkULbLNALSZiUs6FOOoKB6ABR3MG5Cqj3SAyB9rbP9LToKm8ReFcY
8ZRSjNRSrJ13B9FePZbNQ4VN8VTlqbDrQ6WCLOglub230jXntuQ9MYKEoQ+4MYMWJpwaH9bp2yy9
ezAL0hB71eZQZg4yxdPoxCTfXyQvGUpMVG2Wkg01VR0jmd/ppbf+St0CEhS3VwhH7+7yUnQ6vhsG
vDxpSwQH5GXpHrR58LqMAOsj63WzOnwGIcRTzPoAPEW1lK3fX+pQKOeYvz1aEgB73rMoN8dyta4M
9s9JaQ+Xiy5h45XNzfC5+1S+/JMobgPsuxzo3t2xAmY4gvehLF4o1h1qnAJ5z3s53Y7VZDTgLIJg
+QlykdQP0qMGyMrZGsmihJoAMERmqULA7iU1Hhnu9MFxhubuKCVxWL6WSe2fn8rw7troNVSuknvB
/QtYibDkX8gBZlMXqtXVJjVJjdV9QDi+/mocpbyZzubv9UOYxxnd5xU1gk87zJL8jtQTEISxikHg
MJd6s9YhGHwKATU6f/XCgV6r6jrA0fZ/NudNnbdPSNx/XbLhR9GOODunoKfcBW+X4gWCYn0URId6
MzV8nsiYD08NX1a2EMoq68l3r7HxIgtCEAudbbCSggmin6W3CwT9NgcUiTFda+WY/bcObHLf1Djc
mRcunSBOFdFNI5nU/agHa2Zq2sz6g5DDg+Ykmnxbbi2YyikJC9OhROz6VFuGBcqqTI8VVD/Fawqg
tdlOcnHvRhBNfHPqjGhcZ9A2qacJUFjxxHkVNNDwSdNSIktHb+me9gSsB0F9yxp3eiZYjJOT8D8P
mw24UW90p9Y8xX/JrgqNgPMhTHO1aqUUZh91VfmUvaUF2EpW82wLIxePJUtcNum4v1q9exPBea10
u7Lwng7mF3dqoJgMi5jQcqaI6HrsKKYe11Q6HRXGb0AGjgU9ZqKBALEHuVIJLwzyQL4yqu/e24Ll
P6zypSiwBDdYgTVO8Astty2EDLvvvWtuTozMT8Z8TS5jTH0xUh8oI+YrRGPtiRyPyiHZQOaAduwf
u0BX/69nq3yFB/O2YUXz/szEFTFEopDCYQuBF9empoQbGi2Tqg3OjL9cjy0qObIqpyISH/SYRKCE
B4cGoa7lBvPwq7MIe2sjt+bI5phdKeQPX7RgL1OYyVF5Po+XBJZZzA5yBeHhepDOj2rsGTmE+YED
qtlVAGtUB2jYgZP8pCLbbr2xd0ixCMFdA6dPcq1vUn0Hz+GTSogLXpMVVkmm6GHekCVsE+7zQksd
HGQ7vt6rqDzZJTgcfejTRwHC6kRt2GL9VDOlnPlnvcnVg0Hf0T+k3yAQv9W7S00CDWUeHwQCStxJ
f0xitTovsphWsQWxVnua2vXmIaMp4/82PhbjyZz0aCef7jC1vX+zs9lwuTq6qFCwdRI4WFGEUxEk
Pl2dbvLoFybnSSEhWMhSi7+uEdtNb+2dCFPqyf5oolO+64Rc3cjNXOwK/oauuO1vvck6OoWwgMys
vn5Q47Bt8UnR6WZZ48Boy06IgJwVPA29Jc2+OT0IE7F7gm1lLwCFKe7Ew4r54MVbpKZ517yjl/zL
tHqxgblmoqslJrCthihvGkHGfvO6IEGiJcwYxiAft/+61Rcr0G2r7oC+69d9ga73LORtHu+2Tqge
NCz1XGFitnj8bWO9Y5BQCQ3tPq8GRjwymxAigEzOYGcFXnAfexvEu6KOLl0Prn0soQjuSCDsaHld
aKWSegb5EH4ZHguYHjBEnW8DXOtgx0IcoUbhejVOwGR3qMJWKzLGyaFVw6FBD1pr96Iu7CZBENeK
WbwVtc3uDBLGzw5Hm9urU9O59LFofdpmR7wsG0yoem7RTcUwo0/YDk+sAXuvNd79q7Nl0gXZxtXp
G3rQ2iIwKt7nhci0y9ovIE+IlwXVzThRJV9juyuiyUtJ997+HWiMLmODPm+bFVOyQYn2RBN30EF8
lM5kIXTj6Is4yjjE+//XTXEeAyJAtlPPkLaB3FJ7/IVXj/565Qdmw6ppfOOC1L//VMcQ/xTwc7bL
3NchF2DDAESDbPTuuwW003H+dLxlnziUtBtVYHcyUwAgluh/BuKhWwhyK6u2hRbrdGXdsSLicd1K
YGEQGIrYlaNp9cMx73UX91oceR18tE6B7UsQwxUyuYCEB4yvvyEekMOdUVHKlmaNRTiFkwpnDBWr
sRQbePA3I35CKruMq+tvM8r70AK23EMCbA6HA+qRpDyaC4ppUoHdiwno360MokUcR7YMDsWGrhiH
UdOvVDUjpJUTDGVeyz8aXovvHLqEMf30JR26FsNTBJBvpo7xzFl0keNsyiP+DIaosH9dqspe+QMa
zGJ0n4OMj2/JpOo8GBUXR4PTHmZyOHmuISFMgJKxKLbC+3SmBl/U0/GFB6EJ+AHlt8wr9YMkJ+qS
2XKkmxpTmXZahbKfAciRMzOuDhVOt1/RR2caINUTdmEdrnJoyN/nG5n3bAbpLD1h5APj87OfKwA/
lXFTGo1tMCvgY0PFD87dOM84WaTPe5VBNsCXF5GfKSSnTGtHUegKo7gZKMIgW2ePvsewRXRY3S2f
qAPjkaGmczMGkF+OVZayj3gEz8SD/fMbVnATaf56FexxrKi61TPOoALpDxPplVY1sLjVGJz7hVnS
YddxfLvTiQ3nbQufBOrxITsspNEswWr0lLu8TusoJsfm1GNbFE6P8TE+CJ6VXneHXw0lIj+jS13M
+sEQ92qvfjekCz3SPGNlYoW/l/vLqdaht8P/E6Ke8ynubDbfCcyLiy0KXtoiMCp4qT5nJyOyz5n2
HjBf4K9/oYVG16wcF3ye/s9Y6M1zduvJ5t0VP3vRaFuCpcW7oQhrMpHqFwVM9VHfTfPli330Rv66
Au8pr1JpB/Fwa1ZSC5Z08O2pEBa0G51lB6weoY7MB1W9KXFaz0+GjB7ayEtXFigvXrHIqVrFVzaJ
u0jq3vQv5mr2EG2XJLbPmo1KH8IhuicTpkBfZ/Gp0KAeA6U+I+pD2H2USV1xqHET3wuBl68Fe81n
djSXqdJ7Dqp7nH+zcJvKBkz7NOJeQwTZjf8u9lhHZmNCAzbJ5kiElsuu2CYo+TN3baOQtDiiCv1k
IeLzBIkwHHBiinHUjlC/z1EageJULzbVEEabXSvDMTG2l8tOM+tFIg+bp+6fh+JiLmZCq9yFxSt5
wFjet4J9tAkXjxqjFEv5k5H6nUm/PBR7kRYjsmfQOy78e5GWIthx7gf9HvUQUbECC49XOf3YneJ+
rZ+b0lFA+Ps/Kkp5MSfVXGRfkVqNCTwHCZCMYh4x/Llg+eYqNX//JRhz2i+g+VOiHvc+BwCGmdDE
MZdwRKxcG3q5sDD2RaisF4p+WlTHmBqb2/StddSYBz9lX3cvTjfsHpGbCdqCJamte9FcU0TvQ/RD
B1cFrp3CDiRut+KK9BQm/FVAnGD6Crw3oImMrYv/4o9svq+cIeg+trN0r/MLjg6G/g3VgzC2oSiB
XPo6S25EO4i/ImgiWUiBnqfGwr7cwuzkTYNI5c0xGHlIqHSpmwKp0h3bnS4b8qW+7PYJzgQSTJC0
u5j9IAze1OEvEvGY+aQVGyC3f5acL5bIDolp399vlfIHuNZS5crdP3ZsWcGeOgl+1w+ZjrDWCDZu
dsO8Z5yzdG2bQA6iFx0ipCNJ8QMHdAmooUsd4Ql5A2ZeiqAN13eW7kamJ3AfphSCb61eZKJWcPTO
jEo0Ey0axATN2xbhWXdQEYNbsAtedR8y7JTuZPETyUMOks59+FGuCqFecrsvw/t+6ipet30mezVh
NLE1+bSFAAUZC27mahlCCZGOk6PIPExDkQLNTfAEvH5SuOzFDfhsoZmmf0ldur4fvwC/lDBDkKz+
7zntoQUGCIIV8MxRtltKl1LcXQlUb/FYb7uGQ32hS3WveBxPFVCHrMhYex+iMwxymDqxTKVFG6MR
EnQdNTBXbGXOY+nccD2FsGKLRejoqJlnbhnzKdC9Jlxm96qOcl3I/u4UuzwvDpguRG3TRmgxbmcF
ZAJROFK8ZMlXTkHh0HgWDQdBjPUPKTyvSKVZjsXRQPZ7SwVZ9+NAONks23xnaAbxjYlyz/ls2VTO
odMyRj8p8USsWxSmq57+aLjsE37OazgX4U4HUnvrZvSU0DdHml10Yxy+XDUDWofveTqYx26x1q3n
sznoJQcr6F+atBInupKGKMBRHzEFwC4rlqT0lVZiTZuxt/VUF1nYvOogHo6FpIhscsiNeiWWDDE8
kcQ+7PAl/Z8vESY2I2sj8rypPywbhiBUSbpTRKlJqhzlwoG61efa381nE6eKnbxXPRdtZnqlPxM8
ua16qR+BQjZ9U5QjTP1nGpnltHEZCiMZD7ejmpqlsMnKNYFNrI8KsgALmwQWd4S+yAbE96Bw48Y+
y0noa1bykuBTzE5l5iff/g+QIRQZf+Y9lydQSF1N1y8lnyjhMD+Y9v0efkTazmTQbe2Le6uCZN1L
Dj54vMlSAHDXi1mgHDCoPDk8+y+nq70aKkIvYdpheS/loEcnjqs+U1icP5DgcRObyEv1NbnfwvZ5
5aHt0ROU/dQVMzI6t2GsJkDC5NHgn9AkXeNGCcW7gsQnj51BV9GxfLN7npjzKnK/jS0vZeWGcJBS
DdB7FUR0XV+v+/ekzmraSLxcgw5VJMS9YWckYSldLqDUDDh4TRyMXJuelCMnUjU7iH9hQ9Nasw/X
K32MgzDHs5hew7MwK3xk6LyQ+pMM64I89okIIisD7qJUVrs1uOqdn+adAEj23f7ZjmFJ4Rxbl06i
hphEuX1VppkcaBylpAx1swIlgkINFmtGBWZjZV4en8E/2NHadPo4otVUXSTb7Ct5MF082XTMurxL
4hGCSqltY3QUoOEPvykquOJI4SoR1N4o0OPNUqlDD6qr1e0GaSnQ8onmK84GlRNoXKYIqDSSXwV9
Uonr2+YMVbu+PACri6pB40Mj2todVximiZAykp7tsBAcITsoJAKD98s661K6OfJ0XECroj02Fn8b
Tqi1aTJa4nzO/G98P1g9FxxYm1IN3sbIJVd+LEXZgMq0ELtRCGE2KX6VbevaRHfigM08S5yWlafw
DUSlfmNMx/z3VzonBRYG8kT56i1pfxPLjki0ZFg7rkpNGWdWny2UdeIE1p40gc03jCLxa8FjmWxH
3u27ABU+UVkY1kWOy0CgbqAWD8oDmyLsdJ2m/7jd4DCVEhKtkz24z1S15cHWTjJdmDEEMyRf2cEG
JGrdKYP9CXWzfrlCh9r26Kf5N1hhBKxDQTYlDWMO0gq9TU1M0AHHMz97N4xWIcZ/repM6z0vDnjf
jwC8t0o1Tccfs5a2NecRRlbtwWLF0+O9JNPK9emiJeAGjXnmsXAnZQwZmTufcbmcCr2vib//TZhr
Fj7UlF5HO69x3z9l+KFrC77k5VkMpSghPBnGPAWtg3u9SY6r+GO/fJKBD/UTlwAS8zC2SE0jlOLc
RLwiEvgzXRMYuecpQnpd4ZVMxowDufUNMZhdKbEu4FBAxtQ56EMxxt5BV5vGdOZLAFJSBVD4RU8p
FivIMG9jnZ2BpfqDNbrtgDk+SPx76GE059UthEAyKO0pDmKBZ++WdmblPfIJ9DwotmcfHd8jMBmg
b6WKoE0EY5FERf3hteDbkM69LuDr5CZTGx7g16XRB07CQxSUVnBuqNqad2xPtZEL64tiBl2EQT/4
ZEl7gB3vobO6goaPPbtpGCiLpp4gBlQvGJUBYD4wmeDtLRIhiTUrYC2FvHxcD7kvTdQTuMh2ejsq
pHY0TYXp/3cGdM3Rdmd0/uF18TkHAXARaUg4gG0ygDxw8L9peBAsuYRsH9O2QevBqdSXxJpW2E6O
HXC+7tldAiojBgicbgeBD8WETNa8FehloGzAE9nLI9/fAgv6360DBeM8Tlq8ujLiAI2SInA8Z8jn
5ZA7uq1MAPnIyMsrFb5zatvid/Q2j/4991vTlR40w3REAGemA5OKd5LopssixeKAl9CgBpoNLK08
7YNLqVWtpJpDznFRNUslt/uN56ErovjIGi14naMAUj4vYCtHV7jWcVZJt2JcWRQvSLTW+IYsfZPH
rErMHNNeAipUCuayi6GeiHN+kKSo77wsFURdqDXNevXnQXkPhIQR+r6lUEljznM+TrmO1NpVwSDT
oC4nAzOCBnLA/HzdtEjPWISZAv7EKNtEKCEgSOpO7EbcdvzqWW3zUoBSFSbgrYkesVm97a4RXWgL
4mpAyKhtjxzNeQ8Aj54htqubmsjDcUlt7A3L3C/otYg8KXAYylIIAYY6n1wpy4seriyK8G5l8QdM
MpwXwFB1+E3hQERuOOuLTrwiRFglRodmEeyD8QwEObdZ4b0za0WnyTzyAvtFo5o/LPHTRysGKReU
D8a7rS2KSZs9Uj/KQvyFdPktzL85zCZTesmVYSQdnHPJaHF/+TZ6U/X4yUsS0K574TT4jNNFM4Q1
J0Yt78EiqYIGd+2dBSlXNq51GvKiGXC5o/1gCvj4QJH5ynV9fYNHK/1F75sZZ/LpFqGwM8086Usr
It+bNSeWLmxoiRE60X3ORFlkSIowYFH6Op0nEfYTz9SfYLCetXS5gs+89oIeKMJbC6eo+f6LrYKi
14hg62iA4TyMioeUXjZga9+KejjLvillQ6tyLXJa39fuR9IIe3b6MQqyOTkN+lcyjGdKXf0CU2YU
Pf4QnzMVlqnnyp9+XFz6cEOVyKyXr2oOuU0E4v4vpRV+oggC+vZs1XS8Vo/UBZNcqDGpdMlshNe5
EUakBmCp4UAuPGgfnp3USoVKQ4A4qxjZelAChTFRX21ilJEChndhqRjyuIIFl22lYtizdQ7rAr4K
5gLv6oFOxwAL2KkgNX6D9lB/ATQGFcSg9KJPi+4ossd6Ikfnyalmr59UgfvgdkEhjEV3wYgJftu6
hbQviS/Q0jnDkMqX3tmdy/1bhuIja8W5hJIEkpwtGMyAapTwQDwo63EFzyw3XCGNixusvBxw98Yj
WWxAo1qAQSXutIn+/hNqPjAf/EZkIRYIqmVBHz1QM6ocwFIy/GVbegUemoEKh8jqQbnEIPIXfXX0
fLzGWEgZJYT5oJWGqe10fKVEa2jPZyugHtmV061G/SU/LYxmBTXF8s0Bwm3iaMT33YgdaVrUa98L
JsVS2VxQSHw2OUm5WBMnfIa5QBjsv2NrA+ilow5ft0bRSUizymM/pdpKy9z7wV/afnqXL6/INMzq
u7zd/vFzJ1qComlSvTzaWSl4BxtAPhze2jUFv5wC9Z6F0aZiVm5HTK9SPwI4nzpzavAhT7GFI6z4
7iWFwWVjpkzbmMx/7ZwD0Z7Ippn6SaTOykwcVK8e0+9u+F7vjRJGyD0uuNx5ey1JEsth5+92uu+C
YH823MQYog6btXEQyxp4xB/7BMwkl+DJeeqwAASnODmnKa0WUSmohDGclw1n0wdHegMWIDvqx4HI
950zX7GHLjMIC4Dfv2LeqSF4kmveKhGLJ5j0k9I7HDQMMxpiLYd6CG9eNqh1nzQiCjIFfICTpOi0
2ZmckBmRgKtPnl8RSNSNMKqDwyV+Xfc1A3pFNu6M7geM5BxYF9baLSl6+EeeWlHoHWq4Ds3kFTbL
BYVhzaYeoTvIRg3vBjLRhNWpNCNOfhVtPbp5ln6fx2n0zfthcQ5XZeSj6tDhjg4Ll3g/IoCRw/fO
DBFipk9wdfozc6rUKEVaG5qQcwhm7FkG70h+C9xUSyYtniRA+QEhokps7WtHQXJSDSkFrB1AV+p/
cQNbNkPU6ImKywoblzdwKqK3MwQhmV5/6mkGPekWuJYsCULRcaAS3n3hSfz2xgqw/oZ1K2UlCyed
Q9JyY63LhrYP1tp88syF2QNKUviz9Cj0YWr9tQ6H7uG+xbeaHpNm0HxbUGGjKMs8d2CuPmaUk28r
E7GRqOjFEedSK15e0UEEBnQ31ltHKtfURxzHXNfkgiV2jY5UxbAcQ/6xTaiyVGUMWatVCO+YUq/5
p2b61aKHW6fKiarqxWQt+kmRu7FXEjXYsFyorgmzck2eGKQs1dIN2aj66RcjlfoKKhkLeriDdv3I
yvJiuoTYVXRVzd8NKyDDNqb7OocYLEqyyL/Dv9QB2Wu/Kl8QPgaeQxf9iWLxEfYRnLXHKaiOH5Qr
hdeixLABz6nIW1xX02AM3lKYWmshzlvZYTDjzNC/8WmnRJav4LNQvVqK3OUGCF/R+DQLh40jyJEz
6w9hFXUROAzC8yP5JNq7oFNwU4ns7Bd24+Ca2DF42OE4cwD2xaawjkeSjG7QcpIzeDa+wVY4GvHI
ds0/lrLxRF4yB/RcZi8SZnAe2zNpnnfVu2RYXuncgaV44YgVrYKYs/VoOXyAu//f6iwjTsyhB0xs
zyNaGQRotUFPBF9ILjZObiVUr5ER9LW6qgxT6jUgknQGAwMMYNJKx6075iWSEorNsEDEqEYo822S
H3yIwMQ+yktYNai4tIiZ3Zhs3CMhKu2U7HcL/D2y5Q2wE//qlGsMf5lJbRNHyqUKMaOAmiIdZMkW
OYzhPsenAGiQWSeVP8j+8Y5/D/nMGbxFx9psJjRsky1HbclR3Lc6He2I178YEOuJW/p8cf9T6rm+
/VLozG0gcLS0T/OVQcYZzgYBQ/Q4o7Y9uD/O/kVBuf6T5pCcmHvzJG3sJymUPXR4401Q7ODyCC0x
14m/4k5W3ygoB3jgFGcsQESHvDQUMNbOG4G2giVyHQ1gxfn5k/aaoU8EOzE7R3Df3fj7P+Kz3gSH
zrbE+amE8oPjs9hO2N4Xt6z6b5WDXSWoHmxFCwrCiTU4IQxGG0cERgvASRx4j+fJ5qn9wxMe5h27
DP28GdDFyI14qqkHu27eErTBli+w5kVnMHcb7nqI7na8tOnL5PQQfnF196+M5f/V1Sp9p3j3SX0P
eM6jz8nPowEhUUPKKvCpKR8Y9PolBWNnPEsTaODj+Klb1nZeSlbxVRPMtJ3EAWZeGZtr0exrR/IJ
Fw9Obh9l5kgs4LMhADi6RQAXofcK3ALDlELxPmr4JNCVseAr/eVdPjoSIqY1mKsdA9fiphraT7XC
cDNURaJFvXpPOKW2RZ6nlG/SAIK70Oaf0Lk2QB16yKtOsWi5iwfDNpefLY4lbM1dGqsm8oj3yOMk
zr8sAX7upzqqanTu3KeJnv3h1g75OTfsEwSSXSMijSp0wC9S4Nu/wZ2wqyfLeI0BIQbOU5Q3bqE0
uM/9BKVFwB/ZLIr8xOlgkMX4Zw7Gk7yj1BSEzEoSca+nVX0ZXqzu5nJGp+j6Zs/ytafmommoOLIS
tbm3NsuBQZVW/rr1SVall3plkZlhzZt52OM7oi9b6f0jF8zm7NOcDbvKPd8739PYWVBsSdUDGImK
lsastYdo6u45moKKK1kyyzuZoLsqwI4fpmlGkSVRSHjG0Dy6jOKC/0l1NVr767uvhE+hZAct10aL
/naB5I1hDSeOzONVDI9a8nRIVqKoQ5fl8fnli3xh1ske1b2OKz56c94qC1//fmGZZyTyagSrb/iN
KDvxIgSPRA9uq2o8FpZuAdEWEBajfS1w6m392u/aJy/jN5dYG0G0cJ6TM/EQAQzue1gYypiQSlVm
MfoxJBUFZIpu4K9cECfPLcUYEYRIPG5SW5856lhLYww1Rckp/zDVfeelu61gt1ZamgzMZcEaysZx
kgBnow0WsgG6Sswd8UX3E9P/XXQOJB8e5PKTrKoUr5gcJqMrxk35s+aKpzlSJqyywrtyUfnJDb0E
7x+y3id1mpDu4nBiBNLhPRM/9w7HeYTUchZpoimQpbIpOVA5bikYqwGhLK+j1IFN1ew/ABiwJgKW
P/rZkpyFPebcvN9ONRolgyODUPaZMUuB0TQTc3PCeLbU9i3TKvXCiBRlssgEJUR5UBNmJZTCQY/I
DJsbEoKulDuiSswU+G0YraWtZR+vtW6ZIrSVrgm9afj2vbPEKdwE23kH/QUjC16rBW4LTZDbRgnP
+XRkkc2my8QeGZe07iT99SQPEeWwL7GUAe2hvWLSs30f0svj2GecVKeey6dKL5TbclsBg7gnTgsb
xRXQlzFfQFCITZyOO/XIKU5McMRFkvYv4e6VotdS+EcNUYIVhMfpmZtxLPiArBx1P945EhbwkLKr
U9gz9AXQ78y7xawdFwp2YWbVtZzrBoR5inWaXSJfc0D8sD1ZBVBD96siQmA5HA7cUBUs3uJdcfz5
2lfC8OwOTFTP/W4OUSG8g39H+gcC5n2swWZiIgeZohHBZJAwZXDFUpHuapfidCvPy5WumoPqS2on
llxvjyYl2KtaJoMiAcNSrARO+aNrD2Xf/b2gOzv3F/ItlwFIWMFNM/nsFZl3y2ZGN+27a2eMk9JG
Wzck/ZhccLoxlB/sjy31c/A3MduhAu9zqvz6zyybXpTGEU9vPL0Y6Pfpuv/eJyhpzAhQ9GrLo1CT
lsWYg3WT+cfzmKNQrL+Y70RYAyPFNtV0rVANqbImDgmFiqIRkg85VNWdjeyR+HiYvvNTM4L/4lQ9
0v5SuKFMepDjAmkYMmKfOWHFnYV5poV6kZ0N0aczFfoHIWtgYTAVSRIBW9JWJAjyIXGD1wY18zTJ
u3hsZuA8UGGSZnnwHs/8IV3R4lIm0km12W3dT2RCj8i/PYOFE1bJRGyS6WqXBd26YhLOoJ81WGE7
oiqdSHqLwyWTA8vvCG9zNiNIi8R3M/W1niBSZYAAYQ8sB2MVD9lya9HMcfYslQ5vF0BTBlQlCuxi
hpggdzmjHVwUMndOrrvQE1jps0Q3S1zOn+vyTqHvdfy52swY5n0Y/vjM+FkD4oIu44J51LdgwE3N
nZeZZPchy3raC6VQBgsMbKViVzv+WVWeCyxTHuQdOCyOgdhhXa7UrGJ/R9AQqgzZkqEUPdBr9/Lk
pIkZLKqBXyJ1TKJuzkCJarx0f6/WuXeKHXLv8RXCgn5jU1jgBsMcBqb5VSNOANPktE11IZgsieZy
qj/aTDlOrChubhnGOUe2YO83/e907dw72cSefWPh7C1dKI+CGtyJ4HZ3GG3l9+2bzQwmBP5LSKKU
USntq2o2UTcSZ3SS4dYr5CHvfBNbu1wLFja2znhud27xwkXym5Ks0HTqBc72wj1WzVvWLInlpB8e
zJmnq9E1P7PWRdJjVuNrl3ql4lzGbn5Prqf7hrytv43HLLcBbvuOJZQxbhLBoybeGGu5y1B1qd9W
7C/KJBr1x0+TJyvG+Xlbie+yXZNjdRxvE0/wm6DgC4gE+dqn5D1t4B1PYu5gEBdAMaMaJExngF3W
dtots4t/pg6Mrx5AGal+ARur8Kfpi92JrLKKcsSlwLSidXn8ZWIML6mWhu1WDhB5ASOkdhkOH/pc
0MbSnVSoeDm5HKgAMf+EQX1h4q3xAit4kR+plxri8gp4toEkHS1Y1auabTIMdSsVTHle+IuvuuU2
CuMuhwdBdFjvk45BCNjuPIbeCHV2946ZwyBTMW5ngOkEbxgmiDOEoZPswGNmKPPwtC4NhjMNLqIB
nZx1v4CytGy2j0a2BXFsdVMJd/ZUQfP7AYd0btnq+l8usYeWPds+f1UYiBiWQTpF9aKniyVTDNNf
pnVDMxj//T70q0EWBBc8vIzl9sjFHxFWdRcTicI8Kj1PL0wTYdAR9/0X8LMDSHwCSVFlrVO91hmF
Xx61o74xyuM8fk1gmn9H+yRBQXN32xbWf0EF8e+lA5hjTAUb341u96msuCFBPZqmvMInKTkKWDhY
R7uXdiLlcOqR8cTEmgZZKpeqZ5ZU0BzwI7q9weeRJY3mBmhNsWDmsq6kmeDzR50jtE2yVaMEHuoM
rU2o3n8Hdx5hdtf7+lg3vo3n3AJiwBZInIYq/qNCU4jIgBjLzH6b4lSpNNslaNrgbSiQ6WUqWW6T
1yoZKO1PqaufD9BJX2VNHeCPOg5pzycAUkGVfmVhSjUVZUjgZaW6IGoXfO+2prjru1o7ssVfStUv
r6hZlbNNpRLKM6qQiPjWdnf6EcwMX/MHBaAQAX9kYVggtSFbJlQ4kD2yIJZvgyrpvcHK4aKFByfQ
gOMABUJwkE+0/sLp5ShpSP7CS3Gu9cb0/8FJCgZR/f001E0HILYesT3xOix47m40mCI4EnbSeRSB
PLWDcoXGsDfFkpqasA8JW7lkF/pd7aef8i2UWPc5dBgv/siWur46y2qRbrw0SM825CqY0vlMh0h8
S/rXzxU2VJZWa6VMfHD15XvkHMSe8zgGokx5XlzM3lbgj2wqPHF4DI/V5OtteSbhRlGkZwnQD/2M
ytNVzkGKLmwgEIBGJ2epJkrEBw0/SYZNv22kAnJL9JXAn/g6drj/QDoDRX97erE4TpR5D5bkv8q2
KgwsCQtI5/HRPJV5dvbzVJYIiCWoLtN1q7Zvf3U8eZrbm16ZNuybdisMEQFiwKh3OnYtAZktrTnL
0EZtWLB1yVW0swhFxIoT2pcRlXS9S+DxGrToCYydr1RPShGPIcZjvxyhuqWGDPQSpzt8b/k9Qp9E
fOcj6dmx6YcY+jDlsNVcu528m3w4j6ISUOu1ofrQb/z7txwzpoEjstlwSrnLHLJky7jAlLXrhLtL
klzy0Nhfj3jJ8pCohaxEja5FIAtnh3dEvNl7nXd5YwpmNg0lN5vLtC0dhQLwuozG8WKMH2ATtT8k
uKcWaqyMn6i3qF7iCvzuTWlvDT1afCzU2BDu4DrKaEZwxhwNLOM/sk6bf+0r3S59t2oprmGn2FDb
W3S4YRn0dE3SEK2FBe+o9FPN/ALXzFXZpaQjXpWaldSw1VLuWDCvm3Y59E1rZiVmus+P2CRpxVJg
lT1mkZ2baCfgWhyDSNxydeIEcUbGPRWnhnhBNIaUzMPpgCTIrQANaa0onS8ICxqer3LDe9jvJOQ1
0DkOKRRxbFgFw55KbupGtzx3DYTWft7Va7TAmIeEbm/GbAeN1wjE62aLFGYJYnDWBFR0vEE6eu9O
JV6YdcnfM9qPOqukiVRmPm5TyMutWQ1MiPtm4eBGyDbmcZoEIBAbp+ZRpoi1GqryZnOOhM7hCA3c
rAmQXugvenF4i9HeKw8J6eofB/dT61By0sgf/6Ydffwwrv82yxiH9zpwRschDAilN+JLE7gaxdFa
GyYLx7YqjB6Lc9AttJ72CHDNm6alusmtluaiqimzPaIuP8hxtWyrw8X/AvqZMkxWS/nx7NH0YV2T
zLmNi7or1KPWr8mDiVliOYBC0Is4HLkwvnJqdxHVC+CZpyC8Yq9zL8BklU3B4AEdaQ/ity1ofyEP
pLypKLYoOw+/Ng+co3LR6f6/FPuM7vSSEmhiFq2NvmQaFFmc+BX/lj8LdtTXjpwVjysNRXr+Qqnq
7URgsamc7FV+CzVwUb7EL8Q96mKMq3HEOm3eqmiMlAJ1u8lFAHmn+q1lzSfY8SrppCcoc98FwZy6
NXkyH7Zh5NOAanTUD4MTasATPfSpUBRMQHqrTUUse5b1SLie/GuspAtMgrGbLkHd4vO1d03bxIjq
hdX3MaCCj9rRDfYLxRsxJcnw+tKDD8894GJrsK82Ox1lG1iLGDGRMeMq6oCELhMrk8E+cnMcgOor
YNTn7dNGz22k1xAY8ePrHWEZzXlrvo4YvfMiSt3gmiSK4iOEWVfGb6M7vJRATXuDdE/UrGd6Ua18
MwFm7pKr5401LcaWKvJUYNAqz97/n4aJ5n3sZFC/CMEQmmIqkcjfib2gd/ChwWV5wO6Tnpusa3oI
RS65rs1cVv7Vtah/9zMx+60qSrrxXDVWRgr9v7KcwaIbwZjGctbBGFyND0aCbX9Wm77LIASbc5ar
68KuO8rwaNt7ot8jcR5DfHIHM0qDCQ64PCvTVkcyveZjFHi/KanKOBNzaGUgSlFvpnWZPXomgqTQ
uroPZC4HWhiEk0alC/suH23bz8HbqKbFPnBA84qiaNe6Zagzzqb6YmJa65L4TAK9Xhdh/JVXAZor
2IyU8ytfgiok3f401Z5H3XME0B+0RYdWJlEt8xcrhy++AJgjC70CcAtiol2DY7KRjQW3WfK1lfyb
+j+PaNZrg7zQXuA/mkKxO2C4EOPpubaPkl5r/5LuQfMIOolOowjlGtrFCdsxA5JpKCt1Kca0215O
GB0Q2lNbKQORe6Qwjw/xSp+RvhBZjwjT41avdwuYsJ5/DVudmsYgXyc2r0lsfIs6ue1jkOiIqVSR
d41VrscXdDlE9WHf7kB5WRWwPFjgPP92F5VG/ortIMGPuPD7rTo82MhDw68Z+IpaZTVnVYbQ0eIe
2GzAvYL+AhlqVoNo5c+YSUPEo/3soxvrT/U6KjbFbNyQUdcD1BtuHEAC5XwtQ9futfpSrBZzJcFZ
Q7vqpYisUIJh/jNFw72Sta0bhTjFmB9skv3KqIxf4HUfx6G3Nfl4RxpqIoEP9b/dmJMj3QVJJmbU
qpp93YRiG14jQx8SZqbeCVJHNu0paIjdUUQR+APzuUpS9xiEF9013UTKyFqsHKVpmq+m4n5qb7uk
5Q7uOTDoBoEhvlhx8q48bHKhokJ2cSpDhfAXMp9X0FYVmws6xHzJPZiZnnC3CdMJQh8/81j9PQvo
yiLrKGGC+Y0H4wym0MxngiOcknPPNEzqj+Ih2alqPGEhg0j1LRs+QNKflbiwL9k4tIWw9nvbWhEw
796z3oqoqdI/2zl/TiLZrG0rgwCyR3ZtxLEEDOTd0bHHr/zvaI9qH7KL/wbYj5FSw7LYz5h15W1b
AvWTv4oGa9tutTIrG8tviTWGXTlVKoRxb0ftX+i3kDLtb2oI8nBo6BwG56sWKYt+sFjq0lKx0yKu
4MCwVbedLPBkJ4c84MokRHs6OfJDjjC7bPyKF0+t5sRMmWoq4S+LR2xX+BmHNIyJEltRGLNtxyWp
Qr3+inItwJ4UNVSYsBVxQnoCDOQaiT+/WUlgLBx5AM+gHXfO2LTyPOD3Nq45U0GTxEBD1m0txrAo
k6pJAOVM9ebnso8UhzWxeK/wpJesOcIsXjZBL6dfoS5f5J7jmeMXj/WmyVWUu0c5STSawqhztP3P
FNEaAn+iQSyEY3ZUZDdGisvR07Kd24S8gkebznnGefwQQsUMFreORwViSoyBuQvn9UiG87cp1MrP
tyOUHmeLEGmif2zV7SPLE8xUO6RS02hcrrCgmfUtI5aOQeZGffGAHq2d7B5GsrmZOhHaR7pFlsj7
sBUhl8Oq8dAYI3I2y3ru47F+qMA7m4LyFzF93GZqwkT2CpwZ+G0k1wA19jTYjcgw3/+p2jwUZAg9
EpWxjUlaKqF9C8i+P8V8+u5IcdyHVcsRk9LOU6tADnOjgOWet9OPoiEzDh8QtlM+djPVKaqHrKcd
D7UGGHYAh75qT8gECN1yTXuALoDvUGjxkhX3fRKoRRkb5dou2rb45uopj4tnFe0Jn95Qgy3QY+mV
hBwu3pIsi7lX6tnBQe9bQ1WFaMQGk+TgHRElYWcan3r6WKuf+rAemGHUCHf3p9Qet7ST1gegOigh
ZI8ghaQxzdDqkz/3o6GkK8IVxUPd1htAv+kMwrvZ5LxRF8OTidG5VC9l6QijJiqKwRpD1Tjdpmn4
br2yOj6K5aF8zib/XM45nN1XvWW0z/Ex/v5GODd2su0dClASD/yvfVJVcmhuqyYFHu1qp/aC3La8
NcOMMyStLGM7BpvlogfTP4lheB0MbOjtyFjztM2GjEa5kG6pZ02TgE3Su+69ZVAkIXGdb/K0d7l/
yud16mYnVKAzWcl30Iahn6MKvdcwj9DRihwhplBehXsj0TsW0/+BlCjUz14ctwFDjNcssEU0I3Mi
DnBjrQNBAZqPEIE4ystVg6H5xTAxn+9x3S2A0oDEFXrDl7Pe8oRm27cqHSCGUc2JKjRx8tU6ov6/
3Bop9+cj5jZnS0grIM50WHjSt577Wi+KKYCpLuBab65dH3zw7opRQUNZ50rNShT2m1QrZfH8JN/U
vlfrkoxPONIEkimYFN9EQRLKq5MGvxO4ww5aMObGj4qfC00Q2rTDEh8bPqg/ovPOXjDvzc9z8Qb3
ItTcXCluATuo5yCpm3fT9PHf8GJsH7hs8LnKqCM9lbAggUxx09Gp3cqjyabVF+McqU3EP7L7/mLX
B2xiA7Vrok8UHxS/JkiFOvg8/hlfRx+KfXM6BkcIC1EfEEn+Y9yDNoFOsPgL5XVCFlLeFB0jLeFR
rMGpTy5CF/9QkRuq3ILCABwJmfNWaCIRP9hBYK1pplSqzCQ5NqvtUC7tbki8530ZwyGPXv2BeMb6
J8sCaWOMNU2Rwv/mdZ4itAClQ3HD5apwDy7Y8l69nl9hbWwmufl0LdPekYCzJKFdYRh6qZ4sVuVt
wJ6VTyTnnyRrfqE6K5WuY9bqfuoJk+jcqd6OB7WE5+OJ6ZvwF+5x9eyQBuNrez3Qd6IVU5s+aaZh
1LR7lt1wXd60SUgtr7jbkMwx1DgsZiIzFhDdFM8ZawUXAtqRboGnvGlfab5j5MaFoHCIDB36/w94
v6Nc+cZjktt214oKBvDJfxARdNkXuZ4VkQ9aL7xMWvxthR8e+spBd1ssFrd+a+wgvFjBYGDx4GeU
OH1ozNxXHWAUdbSCT64wklRAAojqlGOzJBzZuWKmtrrinoKhMDD/wleGAk98he6ZRKlP87mHNC1x
GLvS92Dhic6bspWS2z7q7cEgwGXdBIwe0TOTQwr180RUN8vCeHXA8gRs3FI1LxvzAM6EPT2BMl69
p/iQs+XoheyOd2yhMiPLOnhbgL9jlhUEHusulk2gFyQdHlUlXRyJt5czigGAqwAzbpHhmMWIOL+B
dzkylyxWsx/lhYFO0+ypElzU21vY2ls2v1sTTx9SU93BwPcB45PU3EVPHJ/xjBoOo9ujQUBLweMi
qJz4KLHIjBCN/jDW5Fr9l23MTAbtAQ0cn5UQ/fjrY4rn7ZrnbDoXy7DHAVcJFzFU5VGKq+AzHawH
fM0qZVXvo+efSyKfYT36G5vTAC4VmE/mRpoYqdTMcDiMU9yufF4ZqoN9gVYtAZN9Fnci4bUrtE8R
t3QJbdMZjJ7Mw3FadZwoQpv4zfsxv+QpNJqEjeU56/SuVPX3XXt+N6my7fpCN78c+vFQjGa8f44i
uwW8pdKBP5qDBTJN2R8JhsZfOPyaCmDMiVIGwrXw3jTZT1KJmpKZBuN0ulOr5JdQNb+Hv36qKctu
qEzLBKeV/VvsCm1gJIS84IpyeKrw92fVA0+TWIpC+sMqmJ7aAYsQZI3hDunoJY56u4nMNXdeA8xl
RtHVOOQ79MstUVg/CoSTbSUnDc28HuKXTQA48rbeDNJOGd9jcOAw/M8MAC540+2HYLRKDWDovNAb
COoVMQIAmy6NCk35x6/wcFX5+/cS8AdoW8kmkh04hSnsKx5yt7RNuoXj8X+gxeyKejHskk6Dyshe
8lpKEBZvgJxmkvq3Qd2uDF/dAReNpnTNy9pLJaHmopqSqOayL0HjN4rn7kwW66h8E/DX8DASzS6B
5rhpw+xcaQsRdw36x8lAlisPyvmYbb8Uy2ochlCnGDjg++Qr8GzZ5M/5NPK8+Kx2Op5Yp0++KH5X
zQ0RVdin4HgM7P5nIWdzXn5Wpf8iOYgzT5T/gBrnWkZN0WmhJabKmq9YWiTXJofihVu06fYZezO3
1ZR9c3eyHR+wxDmhtnrwd7c0SqnWZizIRscsfcXbHbDHPcVNBrPNIJng04F2pjUjum/lX7zE2f3z
rpFCr/rGNas3a7UWcLtmhO2a9ZlKFPDWmUJBghsc+j6Nn56iUF/OIH432K7UcKr481H50R9P+e/M
eGwOZlumYV+O5fwpn6ysRGmIsOKrjF/gzrWfkH1ztHuLes/FSmT6KBkaZB9yX4xZpevQ7e6+cGX6
XSFrEQm0/DAX/fDNX4fJsljAGM34/d3iK8DPnYcAKPCt8ZFdtmLONgPn0ZdDHwItGFaMq2D3t+Fa
Su+2LV/5q6CZY+2KFy5cOuLGQ01Bo3Qmix4dzKyHCdRifid0CSePprYzCdD9jbdCQjdX29xtuUQY
eX0vNltZYA+AZYB5ARo2Zj+i43l0Ib1GomVTsX3f3V+1xe4OMdcdLpD3Mo0eMZMGhwPZDmgjrzdu
Dnpgj6ZSEzK/rhn4jySFyJd6rxitGkUIZ2h7i/nGbAoLJ+dR9qmrHUSiRhI5xK+vderzmhKeKNyO
4TCGq17gmHAUMFkrppMWs+HsszLSPdIWNCaRd2x1XlIBZzKLfEtxuKQQo+jjpo/1Dsf3tcq4Rtav
JKCat9t+tMJNO1M5CrGTdezlyLHDTRig2ido07vFuEjdhJVCvttEKp+urVskW2D9w9a7Pwd724qK
ZB2fRKZOJBawoeOCI8dl+bRplSJp3vY4We13I1VbXOOBLemLO7toVdAP7tetoIBUqlcPBCI6a6J1
pYL5Qz1FCKYwLe9MFmJhbpSJv9fAKdmq6fWBgv0dUq4VhD7GyiB8ASHhE19cZn0MaDZucAX6sy70
AlF/kPW7ullw43Zr3/dwxuAVmBfmWnRco2xfLeBUx1a1MsD7SxkrGDG/wJBK5l4/904608mVvfQt
hmGmvY4degYFQoCXxoenbG847VXyq4BHnOdNY5saOwMNh6sMZDGKxhjuoFvkxRx+huG1SttJjmEO
9X/YD7r9KiqOHZVzqBRcL/xObCaU6H9gO/OHt8p2IVbhm8WG+w/2pB9cxkVX4Nxee4oeAyMcuFjw
BCt8T74/1vZIBfRC304Tzrah2NGJjan+VS7zvqYznRm/SDFkuZ94H9KWz2oHC6JDOyLCgHJ/23qB
REgWNC3NRAiHPSNNWyJGvJzHr4ivzKhp/0TS1vlqlAGGh4eOBeuAXyhjxqRwnnwbvfVGZt7TKkav
4inKdELxYU5T5Q4Iz0/gjTU96J9FXxrKYqCXHuV9Vl5glYg/62/6MD7FdncHfxE5HjsI4whs7Cvh
Na9RhpUECgc92ovORncTrnByv2bclMzTvC4LFh6wIy7mg2O6FqcN5i4d1xa4yUFqLdK3u4JaJMja
JTpRjlnWiIdBDkswSz4tTk+4oJjxTRK9uIGBtEkkPfEOJMOdz28zt7KApCkkqVvBF+5lBIBPvuRV
kRxuw49Xq0O9oC6uT28SpjFMwjn5LP8j8zO/7lL8KUeBP60Ci1tE4Y27XBsGzVHSrrUldyVYiYf2
HxldHSYg5zDWJQBMDUHh5o0il39bbuUxzQ/XFH8WCcxcae0e/XyvtrGGe9T4NtFTojFA/F3kLWs8
e9D85gxgWP90Rriw/TGutiEVctBq/GCJGsZuJ4BnaqVH5GGaCCBjzkdpWuH4d5h+fuvpsnJ6iMqW
gz09JuRaAg6Ce1MHHWz1EnQTcwQPVERps5cabczNSqQzVHCtG6nqAOuiBrdK+mvFXTxErE3X3nDH
FvLYfAf8plyFeSPJZCiu0CP/98MuYPxLmqOTcRph0SJjsJPx51iGndJVGO/M6ZBsc4HqgP+udLVu
ic56Z9r7D/VdWmkhabQ/1d8UGGbDE4dFzaRGhxC9GEOoqHWcJ8HoTEAXNMTHwDJV60mjCnfew2mF
5UwJa9VO/wRVRaMAygmpfOSOHUaOlOUkVM6FVgkm7NVoqLSjJF8uwoPucmMaodopHRJY8xQULEub
lJRN/YbXNAn9IQEHBxt9MQdq1d2L6ImEJ75BqV8dWBOYdrtF1Y8nPq6OxsglUGIINEPsDs+s/BPv
6d+E5Ll4eVXFBvzMhJeDns6j/966BpRIhGRrgcaNCtRJRKoTY6qmYhiw8etKCBTlyWU1deMksAMd
H/YADGfnfmIKtGwbJLiKNAbpvT3Op1Zo7nUT7Ilv9TjN80uDlN3fra2s7fCXHsS6FkJ3JZHajkL0
5GtEEgvu8x2g5LPsPK3E8isUWGYhPj4Z1Dz8uBZIiUlYjHNaIVhgshfP9UhtsOeSkIFVhbPF+Md4
0HGZbzR+ZYgwf2m5kaAm/noE8ogpoSwNKUdFYry+7RCcyWgVDs1ZXq0HEIpXYFvXNcuC+maWbRWP
6IHzG9KYr4hQYLh2gQ4okY2jY9WkmBlHsYhflAoYR1yUtdrCW5JRJq3fkWL1lRSZklwufoDabAHc
aY39kuDWTNHImyQhK7Rk7V44v/l0Muf1VVVfaDfrtvaAARwNf/2+rD/zX1sDLht3DThA/YxwWKZE
PpnSAbT9WCkWsq2EtU4VYsJVMkViIkxJ8bfXww+MugR17ZhnhBoYn6FimlYSUBmlgxkVlrZ4xnly
Fd/qPFH8dpQCu0V9kMvJcE2GHjZk0iapUQuSFwHPbNBfbgy24UGCinMIskAYwKDk8kD1gvQKbqyG
ohIU1N1LwW5gqNVRSWVbGdOY61tXBug1xkxiigodhjuXpPsxr1fENJ+BilgRN92ZOFlBaomMO15q
6ROEPJbSRiAutzCZ0Pcff6fMKZZO84kTf09MLWy5fdsXQdnXzLKYHsW8Uo00QWQ68mBbmpxUYW+t
AHO6JA1YbIt3khTTEBUFlJXaM7ktapIHWAdDBjLvrGqOQXLmBzfJxD1MjaLkXPoVzZNkjNqVOGdf
Wc1D1pw2rkV/VaofEYeL3/KaBMYLNI5lRJlzro8tG+1j5O8GeamOt7Gau7AuSriWPoJ2Sn+pZBvr
JGh8xpM+y6/Aw6GK0tzTy1c/vOKoWcbd3QRdyK4JQLx2xAzhQ5d5S1J+NuHNjwfEErVOi+jB7kPJ
wiYrc+zuk6Lo/6pzr4S+3xUga1GzBVIcPmns7WWxiMhM4Yn+yP5AYyZ4xXJSC6ctQC9UmPjNz9WI
uoGTKBitf7o7GBSmAMgmP5+hP/273Ljg1EO9d0lPbNP8QXUAY16kSzQvw4Ve1/l4t7wnvSt7i3bm
gIu/l2bqKxkxyawx6JlbpqAdwPWetWErp6hx1kak7CgKAyxMspPQ1bTD0LREZu60EFi+V4jNLEci
5HaHKkaBSptHUY27TXdM2ZAPVYtrgZvhhyk2lTxf+XZKTg/hy2pF7fYulCmI162jti3/etqokTFH
LJDGogp4mE+zi5mFefocXW4X+lT27Ll7JqDgnNNwIiU6dEbRiDM/A9RNidz5gVe6HIh3C3VmS+iS
GCWX3txhLXMHWXUxFFmPZIMMa2aop3Xoz4y5uWst6tmn63L6cLdzen4chrkc+vfkjTR5QUVrsVvU
ux+Vmk04thuHXEn106DfbFfeJ4YALbFknAwkw0lBcb6Wbc8REgmatfpOBrQcLxgQ2jFcljpS6pZ/
uK4UKfYD2Hl7fmqZnUd1nvRmHOJ12zznvoZFutSAyZduShykReHzPkr7M+J8uQ9Fg15YUvu5Cvf6
DFZuYXtIH5dLG3ollQ1C8VchWtIEcuoNK/V3Gv0mSVyJL2mgxV5tu9QTgZ+HV5U35er7tJM07n9i
HinrcJONN1GRqyqZzI1eZxMDzzp5vuNxS4MK1TLufOJPwgUjQh7zH0BY2hc3Xzmh90wWTEtfTdSe
8yncxCAmSLq0k0nDgM5CymhzrYtOua7RjmbNXQguX3UHl9VsuwKvTk1y/VIJGtEiC62M1SgFQEB6
+TVo1A4f2Mh28P32qGJHnHCg8oNAZ4zWQsSWNfuquaFlasJCcEM18KNUqGl5YOxPQJlo/0d1kKXC
J0LTmeRILXJl2HWnU/WQE8tvXxDjvVIiKITeBSxbndfHxrC+jcaGUWglyKsKwmly1c52+iuaTkyI
Jw1T5UY9JBdn+Xi0/E731o6BpIzNxK1yhvjN3WK/UBIYRiKbzpt3fQTtPJ7nIm8lWkAo6musNEc+
n7aCF+Y8v6F4hR0BPVYAft+i4h1PpubCI5cyzeb2tymRsJTJtrWyjYGlADoZ6KVPng9mgzCujYXw
GXCmCqFbe1y1u2ekDjuem5GpTK7aa+pFi/6EjSdOsW88HoG73SQN/EckNnhhcOWdKX4Kx8wZEn9h
JU6CyU/f979RBwcBPggXKPszsVmlP+YOoHMuSDoyDWp4Ax49QVmcCCPrzWfzPMs980OM1fxJSJ18
sUQghAknzEU24fkHWKL89O7qucUNbcVQ8aK9Ys71l4vxxTmEQHpQBeckps5nbli4nvII7C25pLpH
an1FUPCYzXS8wxsyPuqVju6HtzyZg7lbFsX3pm4mHSzXZCkvsxkK0GBxpfUEyX8A9TGJcQbJuoI4
P+vXYZa1ugR7CeoyqcwgZMGHdeuewaTvxAmlPCNU7GfYRKsPWW2dD0EY8/K0YGuDP58Xv0TthpY9
ldxKc5COnq5wEGl5ThE2vBXGM83jfuAiSHkpDYTsyU3l8Z+hZOrY2oUxXCZOh/hYrjCYGKj92ok3
0MPnYh0PMkzSbmYOnAr+fJBhoaktmcvefvh7krB90FJSqCeAfO5FBFWMz8buCyAxQRro1rRv7J0l
hJGp9qEDGUQ3l6CWTdr6qvbjPkoT9L89W5FF4UZzvLeCBAGOQcK+Tt6ayymcJAO16V1OwOKSapA7
kMcIdZNr7wp0u3NmK9XMPbzp0mdUHujo3watSo1pBKGfWCU97DMbKcrvTnhDLCDkNB8jK8kFeXjp
/AHxfePWmtbZI6Amp32wh62WOe97oWVYmACFjPLfAJZdmcn6H4JWaybFh/IIu66qGyoUEkTLTHAl
zLtKpnfx3oHzltK46LcDWsA4Ef2Dg7eJPMQ9jUvddez1CLbkNsEjlBtjOgKc3O+pIUdXUsot43HR
MYYWNZJMZgZAA5A3pEdQ9AtetJ8W9OxJxUDUiM5xZ+w+mg5N8Y++CWxwHKi9r5RNcVRl6GYO95HB
2oj3kJY/zczi+sVlodEVjMMzSOfOFKmHxDM9mZLHzrDTMiyZIZMtvf2MqsF5DyTeWGUCdXUFlHeW
Zt8UlHF6dSIkwZmdH/B7ZtPiRTeGJj/W7QiAg2aoc852tfbtxr9Io8DfIV8dJt1QstUwrKI4vQjb
hmLLOu21075kAa9xvzg0Z/qeaCD+cxC1joQZ1KQdkhSAZZP4ZlbgpHWj5QyuOLi1w6vsCVpeBEIK
x/oDDp432rqUouItbzR37nveTE2QlCaCXEPSj2grBLjCyYDAZykU4MPeVB9rsYM7ULFtit01XdRu
FSP1a/1JbJE50WL2182l65W9ezjo/esf6rjai/NvRRnijXSQ+lU0rmQhtRRG3//JFXYRmaMFPsI/
sVeH8VF9U4g/iJVxvhNvMHhgC5u/s4XZdi0G75wDptSN172zCZlASVpqr5eSf+W848zGCWEwO8ht
rdQFTMKwNOk3HJAEZr94Vm4NUjKBR2E1WXy9Tn39qcsYYd1Ogcnk5YRuzzhCWPiK97byhKBrZsjm
PVn5aMx9RxbzPUNjller2YF3JIA8vz5tBaMtJqErvcQ2Uz2YSHMAqJNTIV6UU51DCy65Be/gBGR5
/vnDGTMqh2rgT1IisP3U2hgMmfj5XF0ZBEuUI+0jFXrdCMZPdPDc0oPu9Pvz4yyj1oc0pz92b8En
WTh42PC6U1NezKTBNGO+YgycNuFt+KMoPpwiC3mx3eq0j2+XXpjGXxsvRXVunl3RK5HvgTpn4npM
7Deuk8PQ9dAtAP0Ub/QKVDDz2ZMaVKmSTtceULj72vtOjKDDvWMRSjlEr46xVCM8jQFV0NQrfPG7
z/ZIkRfcjeMP2asefly0wg+QLkfMMcrexyTicraDYVV6jL/DSUkyNuLuHskx+ugmyfPntFLIiokC
Rg7RroOmJch/iQS3SAMw6BBLAUeV3JcDElpoSGc8068cYmDi43EE9PaYvKVOa/765VXl3uxRnaPX
v0v/ny88b2sswjnID8FA+h/V6OMQH7lFWTMCsTpmhbr71n6VS7HkzreCoQQCgs/Bhm9AKK8+XVIO
x0voNr0Hssgz798A2GX/idvHpNHnJwu5BtER72kF2wi0BojSCg4LkpEv0JexL9X3g7BMPr3HtQtp
D+ML40OjIyRXDFfeCH9XuoIacV5Ce5bXH2fmYnw9SHVzvpNwtp8z/6LGqxyRN7zl9zZ85Tv9GrvI
gV3MI9KYRlKOoWc4t3pRbZk3tUuybDGiuhIjJFwEBfHKb4P/TxhKn0dLVJiBeCOFV0+VtnrX06T5
LdtetumEG0pvhojVeyzHWWmg2GbIyWia2IuFg8u0yrp8hBiYIfXb9ZLNARyJyqCdUDBM7Xi+QPqP
JTneGvRvp4R24X6qul+bZnxWp/5w2RTrcy5EbodNVfuiONTdilgSVB7QZbL1w6tpSe2H4t6WSdfh
/yjhhyClvwDQeUVgviWzjkpSyYuAcQxVCjg+3Epmu4rSFqlIATxgpmxlvGdMuONfDRgwGBL/HpI/
RI2PQ8Ke62mKwC46z1xfhcAQACE3WiSgKngOUH5WxdPyLfk2P/GVslquurfN+G4Gdi/AP8IingZA
xuIAmyzylHLNYJ6RIds3nZuoVgbZi5XPMnseYHbIWHMu1l1teH3VWShMTtKE8n+g0gdEFpkdNh/l
HNBJTTu/6JjufuJAPfShWQHN4TOwPOdHjeXuyOKCDVxvf9vZMIKueOFkNVtbzbzrDZ3dRlJYOasP
Nfq877GoA/2CcAjeHOR+1957P0pxGDCUVKakN5Bh1ggcHt+ng8UZ5BMJpVCo+JD6j/IuBjlOdlEC
41OpQfQ+gWT+nz0ZKRCVmq7xl44AzL2z91q5dgurEp9T/3I2sd1F4q3c/zej6mIrmgU1/0QPUH6f
54DBgAqon90+z8PHJbRfIysEOZn/aAfByl0V9RO5wPmulg3mXlFeUsfah5l6jKMfDW3t8BzqwR8y
YVPYHh1H8ueF04fHpuZMdTq2B7p5tx478SuBl4LNnjFAT9ZCbCp1YBXQVran9TFkEZ4vtpEXChjR
3NkI2hENjwYznCsYg3ar3GUIXw93Ut8NSKy/O+zaUiUdkqsjvY51vNeMc07Xtdorr5nLeybiJ4AT
G378W89yeBIXO9QJV5AZgHbjzNcz66MIFdiNPGRzA/TDq4LGn45RE04xzgFmmYC24Fk/ESdnTd8c
5m7kPHNQLsEHaHKrIe8ubOvqlcrAb0asGbMeULaDXX+AwjW8JvuHbHtNOp5mTmp+ftm4CtjH2Mw9
RGbZlC0y8aggUVbdXBkD8F2aSFbhNfKERKMJZJHzE2s2xwx+RBSpn063TZycFq+EqFhkj9zN8VX2
fi+w0aEZI0Z5eC86gudd0X+7AdLzcGd9QfjmWFwgsGOjN34kc1jo1hUWQR3eQHgv8CPyNL+JvoUw
mjBFc51byH4uZKp4HP5iMqbV/Xbw1B2yTor1tFZRaDVZ9/bX4FOZWxaJ/LG+pz63fQcdDy96CmRO
t9lF7wgNIes0QwJ/644NBtrWWn0N52SCBlBZF4isLCSC+osbIke/YVWS+4R3RD01Y5HKBd2AKxu+
Vi/88KEetu+5p+wNLLkOh3pMa5bzL52s4SGbekJs1KwM2vbqIsrKc4LFvfBF+kGyIMo+sxvDwWYk
JiDZ+onRaXN6fymdowuac6Pj8EqMmgZT1FyRe5MV4PDZCtmZmu/+Upa13GOMGhjs51qipcDJWq3m
41Vd3iiIVTyIoNafpzSZQjd9ETSdKArwuErt1ymiKNzS1Ji2OSISLFL7+HLE1+d3sjIezNTxCQuv
sVFM7U1+0dTFnqTKavTeNUS7q5Ikq0IrQlY1MycL0zi06XK36S8z2mZSfTTM1LOBUQZz+g3QfRp7
guPLGsse+7NtRYNaBBhouNoFFw8IF19Vj357+rVyZl9ORW73bD1ZQK/GINtKh1n6NGjWJoGrWXde
WjI1WRKjphR74kcLMQb9myye30flvOzb3dCQjBsK2aNZthD7VDDQ9dy70ABfZYXc1qWGSVXco89S
hJU/G94Vmknhzb6XldPhbRg4+9Sg7FR+YV3/127UdofAWFms27D9xUEwUcENlzY3ndnmVHWIUbdU
MU7U33Ut4ZS8zaZjVIsZ09YYmaFHrso8qX9MYoin9iL/CawZd7S/MIuTE9MRw6R6gKOsKAMYjimt
/SU/y0chhyQh2ra3EBjpY0/UhhSMp1Wk0fABHrdpT7IVVKXHZgWfzBw53Qa3NAqq94agdtVVlAU7
u+FOmfZjCkpZTtT3ozrrkqu8sIted+mNJTEALTWKL+zWBe2EnV1K1c1GUNyFrpHuXF8UdNY0UtTz
g668ZXzz4YXErfivt/s7yWO0GGBftWA2zMnWbOti+KCptBjGZteuyp8HDC53aY9w8Qk3iWqXuK0B
zejxc9JgkjqWcWfRk574r9oK//d0azicmRl3kcpL3OEprPlNA2fMQH88KBqtmD79mbDaKRj6TZNN
uLLNV8WVbQcW3BVNIsXuMdlp4vI3BUmDmyeBvlokwFQd+7OoJ0OB0QBl4c0m/SHC1ohjDUV3Zmqh
3L3R2HJ5Njbrd7A2nFJHjokxksVin1CaXvunnxOXlpM96LzuhXGdRetTZQkJli1PaF8Crl7z0hZR
jinwBMm+iST0yMeQk2bDX2XfF9TxFSGYp2x7T+l/6UiyDLqT1O5si5DLeEftrEYtDLA873WMSXWU
da6VebkSOz+yDgWWyuvppFtIzEBob22Mm+fQLICugFWFwTIE9mYZxt8c62EpWYyF7A8DMl3S73LI
vfpAkVqk6/BloqFY3QLceN8eBJ3jxurWrOVS6CNCET1HENlVmy9ZxecDPREueKCrp2+H+Lw0uUn1
xtjz6s8N6gyyPcNLLLbSmS8LhuIXOuVGB4YUBOks2w+FxzTX6orB3WSLn3DKbtUVIiuaX+vJQGC2
dlPPrSEQSIC0irVUgoZN8mQ66qQHsAQOk4UIdGhsX0Dd2PyExC4KUzmVw8r99oExTaZXwJTTyCSr
SUoj0OBAPDx/FoSz0WLcpYpMwrBvRHDT77ZD/M0uU6lz6U0t/vAFhSMfJSvt0TwmIoh5ANCJydQ4
ZZNdbCuMmxd7/ey8ErjSxohy89Rhv5Zk5R6RuLo+AqZLuRt72aQH8PEqA5HAg2lJv6GIYKnpKOXL
6ypy9VSh56tw+BGAp+CKlVq1l2JQyZjZSMOVMoLx5qmh0mur2sujOhb2+MJ12MwNWyT7uzuE1Q6d
Q1LHbxrfO74gMO2OzYynS+hDt+SUWN2qk+1nZfF1J+73ltKxQJf86Hr32xrjcqy0aVk8UnSJB4dv
UcrSWPC+BXh2Z6lvkcdx7B0JV3ceF/EF3rgTkSaKBWskFhz8uzKStnhkU4DQoD/C19H+g2oO0rce
/cMbVg66ejXT+6SNq8S7h/rrl67LajJ8V/C6DjsTpIApsuyqOowu3uHseLIROV3fkv774O3eTMsy
FNE4zX77XO+LckRKQ2WW03sZp87529+1coy6HILlghV5skMqUF/JF13qHZWM/tpA0DcOjCyYOSzU
W8Yn5xybhjEOmETvio1KsU9SU5w1HcD2iF6aVj3IJH/oWpA87obrOsMpF9l5O5OxilhDqzaZL/IC
vIoPLfQ5+yOy6Yw/jThzaSl2B/CD0B3L4dgWCBFFnZuuYDG2yAAEBL5U7mo8FTPf5TTW/SgMcJdL
IWNz4MBGQuT0cRDXJ2lBOlaPAtAiKWEcIazlbVUvkLz60FftVfSHUq2nVeXC6pfArGikAV/n66oy
QfvWv/jnxkdyqF6r2efKJAgsXnLwlG8A2iTMije57/Cctvj8SiVQNL1TUJuiPHeBIDnA+QVo3fjQ
euh8JUPDncFihtZD6sd3y/gJcehXBFbW/ooHs94V2nkvAKwlmSKhc3OkSi8ElnUACeFI0L5hoPBw
t9ExXmmCMumITkwqS3ssi7h4/HVB8wWfPXHCCoP7MPsLPBFqFLetVWe6jI3x5u6f4dOf3OAa35kK
4H1YmFf8cpDfBZCJds7LjIg3FcjWG4M0de9I8bfVAu3ynIG3VCeTBAPGECfbWRZqVuff66penjUm
r02qN+uggOcuVOXQp/qz8O8GT9HvSKhIijdvyCXyO5keXVJJfXzw4gVw7FA6541Ibn+gMlhepaGY
fWgqgo5ewLouhCMWuI67Q6+qCoOhzLWbH+Rsyx1517xbV6gVxflULhXvLstxPojtPG2hrV3tLPUJ
iyBcESCYaQGP3Of0mkuKph0+7ZgU3EAvfG5t9rtLrPaZaMqZWscESFr/eJiQ96duJ85QRmZbZTH9
om+eThNziXoIzf956D1DXnyACnLJDW3onfrcSCnDwwgQvbe6d0AWg5UhE1Q5Zxx0LsjHI0p42BTA
9sx8ZBrvVPLFaqfYiSGgr6P3HG/tiJsbCbscWl2jztmRlCdeatMlHNcz3WNgdaQB0lMe/tm/CCmz
f2FIbH0UAYXaozV26TNOyaywUe/BpPW+0a04KCxNaPivDwFv+m6n+KPxRdULt+T65P6hLV1+YJVL
XFlopNj3/e4Ss2gTusnbY3WvtO8mR2hyKZ1rdasqcQX27N2xHPOYxTldQ0m9i2uouaA+AUPe1j64
orATCJWmbuyzMXFPArjCpTsShk+TDxwHAX0/lYnQnibAKjz4xGdSkb7LWLlteQpso07kf3pnYHUe
x+grWtMUUV00VB4C7UbmPcx3ZIMkixdEflkgAx0YaqPEoe8Chg+efzqIxT+ZmF8N0H6aH2YDPyMP
4LjsYeHtH9L0Rc1wOUxaj0Prw2J99zgqS+MQLDoZ5pn3G4UMXpOi5YUwR1Z0jyVP2EdRR/Pk1LgP
zO4qYRJy3nlscGnoTCoOgSn3QFMN3vqtGYxY19R17c/ZJNTBEOaKrRaRVyUhYUAqNAn7o05+kORq
mX2zvt6DTkzfiitec/FrhXRh6/xqKkyUqe5er9Zfy3qcLLR1V+KWXd5lIqb1VGAN3h19mfHHoD3A
809Z8X3e44zvI/3xD7lhLE/Ry82evPUCjjRnRMGhuXl49Ck2jPAETCz5w1vdofYfoVct9U0NjtiO
wnK/zmy4lnasXyC7c+95Z7WatcMdS7IEVQXzXcuJ+LHzzwDx5mDiDEKVNQxjuTKsXnYkn2as7Oik
51DqbF4mQiloVGcfCNaUn9mqUiqq5RadcTq1/86zrTIUWOKvbmc7iCl0OEPbmGL7WjhpvgxkPhbe
+uejLtquTV/LyFJXKjiWYImmsYYvzF3BFsfvqhJg2qtuEYK7VG3RXARbGB9ocUc3IxV+wuPJpYrU
bX59MXMrKK+T7ganm1eJVwtm9dS56UCdNJIT+iVoiblwJS1Ii7EMK1eHdiduIATrNBms7VdU25f1
5Fyk1T0091R8J+Y0sVHGtHZ5jrdGYNZhhla6LWhNzeiKcLiUK24fLk0kUjTf7yrkaVJqlaYvzx+n
QpKDyDpwGalsR+FT7D+/+s5vRiWewjxnNzfwzLDgjM2VN2RNWMqog27TND4ODvthYkRDjyqTkfKE
qwJONWd1b5bvrtDrK9pO9o2gjBDPMQCBo/ANVp3fPiPQw9bujiFO7wbwwp6PFgePXLRzMlaTvFL6
9MUw9hv6T6ySmPePwSAq35raTibOMFv/7XxZSl5X3n9Q0cV8j164gIiH39TXKa/yMI0JiDdqpUjH
ZtCsApHXGXqVFl8Z/S7FD7o8Suc86Fh1bfIw6wu8aiYPRnxEe81DpZ+vOeSygo8/UAZOeBewNRXM
lwkVUc5vWV9Knn2f08plM9EsHWmRLwpNoPG3LcckjIFyoastcQeAgGtu66fOPYqPaV27OCVXKWHl
P3qtKwV3A9Pgs3pragMlB++vs3mSZ9csZInpH4inXf53qYelooZ9qcBXRhCZJDKdN0K+PIO17Vxr
qxRH/w7+zALgpRQGVmivEW05kOhUIKUXHt5kk+eXRLmP2gM/h2H9v4j7WKHJjSVOB0Ajbrm1z2k9
IIxaiQD8nPaAsrcHwuGyA8UlaYXp8YNLPsWH1xqE1I3+yM685PZhY9nq7UYmQSv9BKsj2yBecIld
VdOC2gwz8nOO0KIkedl3Gmns6WAjKo7xl0TuqzZT5UyZ9a+WTVWHpd4hPQFnkMLFSe8Cpd1uSONK
WCd5UaxakXBtS2Iq8NW/7pjTRyXsljwynL6jKqxTkwYs4hA4NdtL24ZPYLRvTTeljDLjYPrSDhoc
IeRqF+j3MSGBO8yCf2JjW+Zy0Xnv/+RUSUQvViB3JaAtuqDMJaI8RLfoKS5UCTsVpswYkUTNWdmm
3iC0lK4fkKKiVYDgedKh7PfDceJXgmG2QSWgs2Ky2dJFtUn+NQuwk6In3VfPVFxDaleTdRqHG7zK
ptSqag+djLN1Cc/cGXUfmAevUALa2XHGCQNH9UCG4rJ4GEh4IXlJGXQE/ioNYkKaH67aB548cOhR
saHVsCbCFO5GST7eKqjFk6iPGPfEbxLlJ1hc4AmMhq4v0H8JLC4Udez9qHx2HWyVinX5KMvK1InI
Q9YDQl8Ts7UgMfxaLUCfzanxCRDG2KZetHgnuzldddgh/e611pNWIVO7jKBUon5I2YoLPqO78Si6
efEIMNSRl4IJ0pLMobPqNBJ++0JTecu9BjtquD7BFMCtbb+vSqQ5/1m5rm0ZGJ4v1t8VuID+t094
v3mIM4W8WztYht3Bms7YcMOa5nN8wCV9PS6zkFg17+fZZcvOMwAKfrjG83vJH++hx+HWBKrgpKR2
a4isXon8mxfDgG/3mBVczlYtb3jFoE1yP13VvHW1Fr7d0Frc9gMkDq6Hjz5Q4GepufX2mEYwZOun
XgxLlS3PiRDLgIp5j1KhMqYR2eIvTKL6WOwjyAwDeprZocnHXip1Lkq502zt4ILy0Neq5ueFm2QV
xqpKRiJHu3HQ2yJe74XojnWeCJLNb+0TU2Yw9J4TbMuSdeRMGgpgIat+WCOWZ8mwM5kcGcctrtkb
eMYT+QaIFEFHGu/FZz8TG2P3/xGQtxY5+HA+a3wyPuwdacRvcHPpJ4zgHx8VdLsxycHkcrUxvoiB
1g2Z4gzIQ/Ex9Eft7n0ajdw+/PbYiBqZywp0SsoQjwrpjRjIBNwtq+996wVgEcoC+ZtyoUStKQCh
OtkB8i8MJ4Ck2sGjTvvFMdq9BVIFqyBLQBhRjJZsU5LaUVFD6QnaqwzWxYPh4HMU1kbfbtEQn8ce
DcwAHhDuoUii87a2WVAoW80wcLO91QYym8KzJ9wCSyYIVLDW+xGtgyrJAv9imC1T9FavkvvifqUY
FQNubkEJ6+xchAg6NxYxUp84XrRufzwq9NUmuHsqhlJlrZ/lBB4+8e3Q2Y9WjQaap6ksr6kWFMzg
8fNb6eQ9L2+qz9XOiFABJ1+tNjRmq10eTqG+YG1sQtdtWOj1rZ26IQLz7tHCXIMucuDZP4EuYHk6
xfbhxdZEQYKicEbENGGOeFmI0S97zGRK9Ux8icMBHSMsjG3TMA+g8rCxcDqW+fUeaiTiyRmCMa7M
MoGbGs9ni6rdGPGo9rwScUYc62VWkbzSHCtxBcz56UhEPeIfGDRZb87Ym0WGu7kTIG6YKEG9I+bp
ZjPkFT0BEBEf50bO94QinHS+MwWwor/tcabQNYNANgWDHLpg5Eg5OggToS/3dA==
`protect end_protected
