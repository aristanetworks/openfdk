--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Mpbjqm6x3tKY/blXyrCD8Z3t4XwDBTLLLxNpgyhiym8/9DfTcPohs6GsQrmFuEM7J9X4vq5+DmVV
FNZSRrW3FoRVsHt0aWjCcnIeccmijiutfVnliy7lzTVV9J0/CXIL+c6s3g7g/eeBI0aWgGKxv7+p
z/LSXhcOmqO+3J7UoVLBzCbK57eaezRDv/hPnikweYdp0MuOZD0apbgIDiVLbSfuZNM29s/QvjpK
RJ3CJ4d62aa4Epgmd59NcvnAhNGlNPW2jDblwdxYlLHx/4xH58QsyKpcrObqkOI43jF+Gd+VkDYo
+O1YMHH6TNFuH6fMBDykxAWbiIxgYym9G2N30A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="mDys1KoudjE03SrCQtpimugp8cMb+6nm7kz0gH74b8U="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
EHkJY/dTETIWUIDylpSOHPa6Hc8WNXG27DVdN50GACh4uIH2eSDosI16FzcI1kmtku0c2RdtJuq6
1PVhH+5NavagKmVJB5wvTUntQezaPNVJvTKrL722M26evs87SIjTkvhoujPZ7jCaEMOHn0DYMyqP
eucEDqlnqnlyhf9EoDgiym1ON9bKSevE79hjaXzPfj8efSg1ciy0AavCivLrO0/rSAXkTJ6As1TH
QzQaDLLJHvbbiSNFjvXVLs7kW7hi/oUNNjDdr2cd8N+oI9hqKpfPQ+NglR1Ua9tZc2FFbh2+9nQC
8LpASltbSymQVL5ZYBjkzWikPfjsY5RY6jqQ2g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="bX5ZnEp0YSlxZCoWapoGc97vtQFdueHv4la/PHwNUrQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7280)
`protect data_block
i/gs81aIRblUkIueEMDRonv0ZsSa8tJqRDmt3y+bnaxb/E4gELkO2fVy+fcNh8GwmHsOvnikrmC9
IOHLZUT7dStIGt7qydRLbt3IhbS+hgNbDlwyUlZCrkztt6VczrnLXd6YZV/ENt1g2lqFSpPK0iS/
S7qDstxX0nXFzyjXcmHBjgMffYyrcVsBz/IPYdAdVHFttCuQFfgXSgtCrPmw+7ApSPsmOUpcWab2
RIo1tPYp14dqAh6wgQ+SbYlkRj0+SY1zYw0x7M1J5TtoBExthrukLr3bII8N2figtR9ExyPcSsDs
ei6rIdhZNgdjfyQ08k6u5o5JcwjoyGvyd9WzkjD5YzV6rrErpoT5USgnCI/5AQkYIbEP/ldRSkB3
wFRhz9fSGMcFdlWpY+7gEYGt8sSLfatAQ1m+Yjw1pYVT/XpdTgFLP+POdhPt6ItiTS7TleDUjjsb
5aXPenZ5ZTjxZuezYxPiybxbPHwdhETIy12qgZuvk0K1Q1N7X7jIxVEAkKmnudtXV23/F96A/eO1
iRkJH+4ByrlhgDkLQjFIL1/R+5cr2gUzqcd4R6DkG5CAv6tmncN3wfyJGrIvA2TwK7pD/uAoryyU
orcGXZJzpTod97D0z3a2j9UmG5vremDpQcpUMROHOab6IapWLbQ1Gz7iVGNpn10IfCbP6aQUyMC1
oVJPC2RVVL6ennpr7ik4GV3/Dt+z5kEM0X0Q+T+FPmZYoSobnWfOsreFTGtkAEMjlQHQ9IMWPwJg
/wN5LG3NurgiISRyWl4J2rFwziFQXp+aEfifu5L3xNKUfrzYhhPsm/nN2Y543Jc0vaKJfhukqTTt
+x73I3/TAdwMlwSk2oX6lszdhmK06jBNTAUBqpVy4Kwhsk6ugl8t3hob3nAbP0pI5h/Ok8zLdOmS
+M7VX4e76nB2kgcmugYmnci/ntz1uWxY8Ss7n9DZP9Zxlt1JsTEjzSjlK1y5HPjeaOy+7+HKwZYq
YQ5Q9468YM5FgC6CabQIg/znSRNEM6slHVRuSXjHqqudmgkznfgPRDm6OqgiGwFS6zm7dQWgf+Wd
yIydnmPLYXIPS6kIdLEkuLo9Jv8EwY9x4r6S0+FyRfF7/zmqmU8s33mxzJC7cTPydd+UP8Fhw/S2
E8RgWvQhdX7QlHbIsuJyeDA88OWd9kD2QnGBbiqpkqS3nWCjOi3N54mlmfT/Ou+p57pEkvU5dzIG
0IWYp+fT1i62FtrazV0df+WLCqG7wvuyFi9oERaE9DeMVi4xAtNUhn96wp+K2XrOp2+CTUEnrhM6
gsPEshTfkS2xGTy1v0JYQV0wwHTuppYmwrJCIhuyaBG74b7hlyauYw2+B3s5LsMrVL7p2PNgJAcd
0zM5k2V0K8lU824TUEZ1Ucd6wEhjhjP3GuCXuAuURBtcCjHUM0ZzWZjc256ipNuWd/OjM839a6VR
GL04NAFE57bHfezYOHaw1ikJ0ZKkOSfAaQ16eceF68ivKgJpIb+ezx7T0AyIVhpBSKfMzzmWsbEZ
X5Rjk4ZFfNwVgrjUfghRdqN7B+BOeMwQeZn6mX07BF8QazCjNeX/n+thgiLl37wT7LRudH1LoS4J
voBSkYseE1/33dwQ3XNhPj9Luu+Ww7E9q5aaOCGEr3Ws3vW3WO3MEB5JYh/egik5O9+b3105alms
6AtCE1OgTivE+ThBeF139z4f2cexjgcI75Aqo1/sTKoa5wd3fvJ7F2vzuBMDnW+u5KKksrvPPBAV
HLe2438yrqwCf9rA7lTBnR4ZvjivYIpdI/GqjpI71WBi4ehOSr4ri1vya/DD5DHCkVu1fcRLybNl
uRF1YNXazskoWZZyZcfXmB/zD1bc1KIciSrnwOnUUt98GFU4kU3Uqf6skOyQE2kIQNmYZAC17a/0
JtWAiIzqpYMRX8THhamBqAgSducmSwcnnXfsmBltGRLZQQGaXxQoVHk5GYnDzkcy6obWAWe7xOoD
x4uupqJx5wSxOCnMa6/JV0xxz7qlz+wL6aJ9MfXkBXQ33cwB/ItfrptqAsLr2i1JQtIMVq4rT7iF
a71ndtvM+dptYWrK2rAnYpAbNIMz7JGTZFVBlbq4tZvKRkDhwKYEEClPlGkI8kTQZaqeO8KB9tQD
ZEUZY9Xz8KRajp5ow+iSjzIB4C7jEqQW2G7Vj3kFLMZMJlz/gh04RB7QR+jymtemxBFNZZQ596Da
ykWC5bCt48bm/5XCL86OQj0k64GIfZyoGTi9/DNOySHCCwDL/5pFPyT28J5D6fBMDhGu1ws4otXk
0RP6v85ha4GhztTpkEOm4NBlD7zLvzBVs9BnrqVDeGppyFDGoJRQS3TTY9kgyHPBSQben4n10xky
3bMcu+ZvbIu47Or+qq4PCAaMb6AB/H54t/ttPacpeQA2l85e3YGmewA0kPNsz3vYUSpNdhWAMSAl
bQJx05YYSHOAQ7PtnEp5phw749xpfGCA2ObNM6ODTdBIUcogLPoHT92ReN9rOTOuXiH3zF9oJgMf
dUW7a7B7hoN1/EoUWASMt3GPaOQB04r0/ILpd9EaVTlPyNlRO3ifXoWPaMuKQBbbAjtMlubIsvtJ
Q4Er18vbTqT/RZnMISITPLwsDLBb8HAoxC40YBjHmX/H/NyDdGfENbcNtiWVVJ8RXd1HeX3NcLP2
M2Zzma03suKoiAn7ZkoQ81MXJ+VntbHvhsxIDZKARXxqhk5eD6TEu53ye221/GNh2cUwufIuFtzB
4GtUc83g8obKYhq7NZGdHxqBz46oiM/fznWoKX/GHXSpH6VFzy2dSmQO0g7aT+lsW85/NrMENQcc
ai6W6W3hBqiEM+onzgQygD2E74cblQH9i4nTbp22lKNjLsm+0lGtDpB7bwwLsMBld4uf82YMLvZJ
7nM4SyfF+dIe8zcyM28iimzCT9G+1KNx+hPVh/Jq+vV/V/nms1HLDen4XX8vC0mdr7sPLtn8dSyO
RxdntU+HscCMeIOqn+RFGPoOD//cFYEDv2wPkQQZ1Or+f1KoH1thd0NkS0KXBg+BfQp/hMzattEa
s6FyjaZ8hQVkxAeoLj9NAm4uQbJ5qwIZZQgjjMlyMxQLk0Ttm4D6s2HaPkuUhWzjYXOkP2D04wAg
xT57gbmwt9ZjBbDx+ER+cNvdc0cl1YtIl4B4K/lkOuUFolDSQ9jDM0GAtlLbzoGCg9UAQuo5FnpC
5a71NXRpMs5nmPX96dytITfAcdCJUK1iz7Ie4KyWs/HD+L7V5Vsu7qOyrW6j3v5HmpWaS5gRqkjq
xtx63xOuo757pizg+7Zr8r4WL1LNkmOdyLmIm1Ml86+tszXRBptr16GEEEB9t8pcZr/K3+Q7lJkJ
GRfXFI8bn7Pi8D8vlMlPeyHDu7Ifcqu1dYJrsICwKLbwHRUGEjI56KrWNbHSfA3mPhVpvFnss1Tj
lD3OxP+3VQCfszIKwtqMu6Zd4Tv/mxSnobyDzuALB3N1WnNCQxJnu9p4azilYEYqAOn3bT0iRlIt
u8ihzC22fGmcNaK6kbWwV18JJqI1rDKGSXwMgQuhXUYVCUMGNrmAKJVbgv1Vz96jZnZuGlw5Xkyl
NwvFdXt0KHavrj8/SnXdu8uJqdteuPP2x1VUkPbKCXyw9VHdXntgdN4rTzVvcodiPjYu+lrF4/4h
WCjDy+WORWPRhBb+8ND8N9SdaRMaziTxShchi6yZu2MAGblpk6wntu5LwfLWZd37mqPUI+YA7SVf
fHC4WED3iHOwrfjMASAdqXkiLbsp/QjFGIpEQFro45JR8GN/bsywfgAjwI0tuc2hWb5nPQnkiyij
/M9VeBJXe9xFUEBcwxP8rAadSKxESQM4ItIdC4mM+JhUrenO+xlgcq5C5VDZUcbsfpzjA0ciQKX/
9X2vw72X1UsQqTpbKGywrWUVqYcJBMliN8lcDlQAoAefTS306MjbBNTkM33PDjJgHbgNKPr2QYp/
+uQs5H/bfpq+ASqRZgNK0qQIt7Oz+8NszIkmyw7+AKPHNJvfGJsjzXMh+Shd+EnOBNTmfT23hoN5
q3xTO4gqGT2PJJFJ9tq9920mylL1joG5Ulw4IvClzELkhxtIlZMwibQtdQK/TBVB2b7TxBwhbuJj
xgjkVvtoOXfgFXA5Frq2tf7UhUCVMiRFbyEqd7bzGFaB8L6QUfLZo89ChYosa7kilupYfVt59N1w
APLNPPA9HD1YVP9dnwsz/TMGWdM6np3J3XlSSIhoet/zhm8+LKWYqhHaOh/LBGBSveansKTNWhtF
DA3oUOM+RPAzRY/7b5Y+GRbq4bzs5VVO8IiAhOiDIza6UG1/trYZlhoC6ZDwmzzkQRLCNW/LrIDC
+roQi+9cX6ne1/Czbwr5qvp2ah3NNtPJ5WBFVy4T+3Y9yGrkOHZZltdU/+4TstXvZXJMENIJRKpz
awr3ZodW+hHP+JGySuF8UHUtlf7IzQSNyhwN/abhazqVrWqWUIL9EoE12xzH9Ywh3jNJdaNud1pv
PNB9dJxghIEFnr0UHEnUBLaQykDxGHHyMy7ao8SvEh5O+v4rvSirCyIkI4PAEc0SUjeT2Js44lO8
pg/ciiC6RLJfyyF52Xb7CG6q0QnvBHWPVarEiG8S4GQRJRISNnstkjYyaYIw3qKknkhsr2OhXLSx
HJYglYy1HogiKab0Fs1gCHgMg5Mqrz0QUFAPtRo0wVldyx9CydwBtAYXt8ZmRzw9BmxF/djfsGSD
liFyzq4OvhAcuIQAaJWAhhIRru5Rbm6xqkMME95cX8PFIpQ2w7H+LBXymKR/S8HQscxFsgTJU30j
FUzNbgJBPFxj2sGffruSdYNjqyWWq8xcitWq8/iepfOS1f29RELfZRPM26ioOVrhev4HZOjaR+//
tdMMqTOHECKr3N1IsmLv0GzjW0ET2q8fBktAdSmaLqhdN5glz1yefJNCjKXQoG/xBOZX+nIF/8+5
ORCDizUQQhZnaAawXhXyula2ZzZI5Hqt0i2yRI8N+RrjHldTpllhXv08TrTVdCDEhO2A2F+tDKXJ
TbdA7AKs74GZNkobC+ffTYAGiIPLdc6TYwbN1DrA57lJXORufVh19fQbBQwjob20h5eExePdJPS2
57/SWpqAow+uGEq63cm1UGRZyB1KtE0uY3OVugyRsXF7r0LDI89ozRn+euGsl4AqCc8i9fP4CMxO
22UI8MoJM8vtnCC/wo9YbQ7riKvXKUnK96T3tZ9BXVxvg2A+FQ3RukF8B1PQ8vaQLxF+t/KnfN6i
F3CB1M8ikTNM3syDXLI72Pc+WvljhGyAmKelif2wSkkTWHCx6UlEKFTtYKYhErVKA+OZKimWxgkm
1wewA2wRAl3SuddePwkdj4XgpNXZ6hvXR9AwTQAoHdjoRCZiJsAHr7JWyj/GoEhfi3r0KJznsEjW
wtoWC/33sq3152Kcs5mWokF2dQLr2RZlEiSWch975270L8JOIOzs6a8dRCIRMIcD8Fpqt/FVwC8l
Pkl0EQ6W3cCTriQ8Msn8LcI/vQtU0zw4FjBulgDCcLON1CHzkDTbV5fYUcyxPr+EMclo5LxdySP2
1Npt5y0dEUBOAlFl10y7qQGGhebZ8ILCO240dtoHFnhr8qy51jBDzfzAbFCe+u9ky6OOS+QxLQ/7
2YrGpAp92VGCTV4OfzPDx7XWer/llk/ePx8MNziNagX07ZpDuVXcEAgLA3bzB0QQKL9iRC0et/Nr
uIgdPUb93aFyEARYvx9yH9/9wp857cKnx0e9nsSKgWSQqKKYrXksJq+BGQvqDxZlv15+c3LmPeUT
S4wjXqJq9JZhwhHKnFem6JJejElqjP/A7mYLdzMaQK5TTXCoO/ZEfxNz+3+LRMZ0nmNbsfk+vw7r
CXoCmrxnHl9XtMzgXP4I9YDkuPo6Yg5NiHiKRmvUOD+XIjmRu54m+8bYk7W/sZWGhBoRwXf0mxYe
pVK56iJfZ96I3JNdq7lJB7z92/FXWq1wZLcWZXFqfncIDZBiul0VlpOwP1hQmwgsfGTXrs3t4hwz
dw/wqRNq+wOWLFkV9iw1cpjzhcIN8CBdZNSMdgBNJV9c0IxnD9cXAhi7CscC5+gn02aAjipbVvAk
euA0cTe8z8djDOfhiHMQBzYW3N8a+mdlm2YZmHujxuMR/M/i0Y8v8JRpazY9BnxNZodvvQVl/QLr
JBl2/JDSAWo+I5ej1DDD+mljfLe3TbOqnT1o4YZDjlMod11mLuFjE2UUejO301j6CbUAB+wqag2l
PAL5QlDkTPMujN+lIbgP+RqfD6dQm8QWr8w+nwnZ/eV/9iU8KD3NfbvlQ+OgsU9xSaXyW710OvTx
hTwEsFFMj5x18/7cnejsHlgPFeS4LvyUAqSIox9JkiQzHwICsnz5Wbk0iy5vsgHQu6cxG8t3Iign
8/cKX6BaZ5Nk2tsc2WYSF1GMyrVMt5SFNuKPhhj2LLcSOxUAMk98scz22vU+O2ZgNtkWQ2B92Y8R
tT8fZ6vNfb75YBr553AmTuqqJ9H6A1RCj8Vk1e4brU84Ft3+BZJZX37le8ICT+K/J7BW1voAd6Zz
H7gGvbXhUCdU+jjnUEZazt1IvRScXMBwkb9Efnf3Ir8eerqQSxzp++2EsyA8tb6ANQky5RKcYizH
TvcRblK2LAv9UpUA0D0EOa+f8jU57AGJAM6I5Gx+Kubx8w/0aLHzMUayuxYfeaZVjrQtBVfq/Nra
ZhzECvFVCcKyLN33OAQk8d4CirZhauiLUY6Oh8V8+8Yg/rJgCyKpbQxE+85WbabKSkEsA4wOw75p
RO8UymbLPg3dzZD+qp163mx06v2Bg9Y6+idH9DDjwcyRDBDww0EcVcPDNg1dcC5ubTWYu/jfPShA
cXA5g4BV6RjKHlWTt1s2YuE8bZImKJamFLZBgbvduvPngpunffx8UJCpRxkfLm12CwomjoMwSpW0
daRcvGv16/rwwfzVHAHPSlHz5B9PvwxKASIe0z/+ZrNskPOrPSp7wUF9tl5wkthYEyUGHUwz93Yg
XUUp4L7BBCdRJMmgCCinddowazK8O4KkreeJNW9E2aG5jYKa9hod/EmQhxCr/FxukO4xoheNrrdN
nhtIKdFK7IIh0Q6rhIDksy1vva78bA7LUTgLC4JEFylT+HDTCmn5ShxZcvnPi7NahTKfskQFAdsV
zpxfR9r4ULRcungl5CDAjpwTHY2GthnlYDrKWlmRZK9bPeWPThZzAABH5o+HXgVN3pWbZW0l8Jqc
Es+r0GT5Qwjf+Q/ZHCnixp9TOFXA+Ih9C4jzoT0GR06OFTKsm/6KJ/7kju7Kvb4oEnoBKwwixhIp
P4ZaZ7r9RqYkJfRvKnSccsinoawZ+wZm+lhdMzmlxRbu2yNJyGeDGPtI+fQ281G98c/8t5WX93JZ
iMazOnuM5dtm3IOq9hJ4VyuG7BodpgF7h050nWmTCcxWf6W4PzeEHfd+S4zKrwvGN3IrYARC67XC
njcCPIltJoATZb1HwKdd9Eewnpt/ABZuyMkym0j2R87aomURa+4N8TsHlXnyPWQ8xYar+VxMYcw3
hahzJ+zzcPiZXEoCGphs5ACOLSLAVycfsiinqNKwSbq7avOW9j4OrJ/CJ1lgWqyaIMsveNVhB9sY
SKAyCkYhLm/8Jroc6J54ULc6DayhP82SQ0jH+5DcqCG40WJ/ESHoRt2ie8H3YC7JFSfQlCfzw/8Y
/vW4/uBW9q+f1pDC0GqBzUaRAjVY/WfZFVmHTW18330kmHNYgfGo4KIAc1V1Z81mFcrMU2TuW4Kt
mWlGnDWTRR5/mY1V0YvRZQcuf3UZ4XnlNz5gwjtvErC53DsRdmBD5oj86FVuL7bMr9MFkmRNDm7k
uSa53tWNAz/6FbIdGE92K0fmHNszjhzv5TtvcmimYtCu4MhZ9bLTOYjuJiNWFT4SNaHju8GZIHdL
V8H02QxRRhY1B3XaLs0qtv+g1NczxEzyvK8TsPTsE8RpPA0dW3vxLraCKDE3rIw7h1qgYdO4tpkM
crONWNahvYhQ9PlrANeDcbiKoJ2oltDAsYjVXCx9BegCzsH2NZCB5B1KS7jr6d9BApRxdiAz+6yN
tewMsJkLNEnOmrw8Olyos7VyggY3eAQylhomoKHS1aPGzDD3zQsgIihATASGJNN2Hq+vKbk97N8d
HTJEPACXdRycIvH6lbUx9gU2yxC0EKGau+lyTrx2KOY6Inpajbi8eDiivXfX15JadpVlUl5ouAIM
zMHlKKfu/gKi3c/jpO721yu9UMWDpjYuRkINWWkfQFYdqv25S3FDa1/6ZcrAI7YeAdounzkR68hI
YgpnSI2nm1Mfa3eEtd/AFjDyaT9F4RwMhAQ+TfBYoU/Kx6c8P40lOjmnbv25YGeRRMk5c0xfXeXX
iT5xmkb2SJ27hz4s3Glsa9Iqygr5nCAmpKORiJ8LY36piZFO6kMEbf7l1JcGQx0YqAG7spTtzQvl
0RZLiWRtCMTa++mVZ2oNjBZlsgVwFpbx/Fg7rcR2uQCe7nMe4JgHG30hzPoveS+V3s/nC05Jr9bE
u9DYrFEQOgv20YhcGgYtA0VfTPFW2Suc/cbjepJmRmGR/TU44lDmK7GdsKakYntHu0rJiYOjUxa+
SuDN0/knNkdeNVPrBcA49X2576xh4RG7zlEx8XUqcLYb3bPTj3MisRPvk+ZHX88MHKuByzB0rBKs
Nto2dzWcgfl/GYbcGNONY4Ih+B3XaO8PgzcZSQMlfUenqjwldIypfvsnAR4XR+oSupc5vwEfDULF
e698ls12IsULEongRv2VNvCYyxVAciFQMfm1uN5WJwDMyc35gr3mpx6sR5VQMMhrYeK4Cq2SK9U6
TjuGZol24zBaN78ZLUtJ7RDeannDUM86PxxRBVrNelO0GuE9nbXf1R6Un7oB4VZq6T6DL6lWXDfA
KBJFVPaea4xMOm75YiNRJ/vDGRWycYloI4GvyxjvXnJsJOVcnqZYCwlLUzMnJnJ9UILCnEjuT+86
0Lmsae8ikZxYwav05xRTLbINz/2ZWaK8bGkhCMdrlOTYwRatFx87lmiJdlaGMQ9nhQjwgEi/9KbR
9FWnPpPcCdmK3vW8E8lC+XOhFpCR8ZyotxWwIeb/ILSRTb8oYU99v+a3k4kr6B9mmiXt/NemjC08
Ut/bJKsVJvyTJBJoBj0GYth1Ov2RcYZA7CxsO5UPN6BAlCSUcjr50/e4GUKtzVmHPu+2SesYXgWn
IR9tpfm1Ifytl7firKeQKjMtXjd1oCh/eE8500muM+i0NAZPVrm18hE3MXKWzzMEu2VTJ0C1Q8hQ
BHcZGpfLgr3L6WdbEd+NNesCN9t3Y+GrUN1NFtMj9GSE2aUUhY1C3KeaWFAuclXGwRQ56AwOUyWr
kuUfAgSyGQRluaotKutOOnrlqXaFE+vqZswc97FUfTLJbth1Ra6TFn4eChn+zfd+/zpUSPKzlmmp
MQNdS+9/ImLdfb7a7WD1DS8FWiENoIYSB7/6C+PqiE+VmGLSIHqgpwEZG6vlfpfvvkj3c2HNXtyT
EuNtIPw2dXTcXnsmgGi84c42bnH8aLg4V9EEIi82ZegheAKrygDCTic9CqQUrlT4E9j9UKaKEdZe
pten6ZDqhYymnS9X8cgURHI4WQ8vvYEZEZRL+OGSD7/DRxvdzjW1GSWT9X9nhayIPiLqUgT2jSHg
/fvRBUu34617+vn8QVif/hotaKxS3AnpSR35uQggHrBrYwvr1qo1Hl0=
`protect end_protected
