--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
aHmE86jdfWLbwjzluBJ93LCJGT/IskbKLB0mVpSaa1euJ9gtkHY7fKf2CZEeejc3DKmz5+jPZ5Z6
XgBzBNQ+b7tJBeKISWqOVeyitqtgXuDNsYACZ8LQnbrFvnHh+BOEtg40Hkr9kbRrKCHQDicVZ43o
TKdG5kJr2PfnCGaIWDa5a/IYlSHLj29O67aXxIFBC0/bU2gETp3fkzo90S05B6Fkj7q6NlYGrM3c
WlxA9Lt/7D+0+zg2OP/u0qPEScwa4K++W6UhpSaEKtapjV4iixPYL7TQtWE4Ut5ZlzYPzBKvnpfG
5ZgFEuwCWjv/5BtKuCqJv1f0v/BcY3T+7heLGA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Yut9vqKU+YqlkYQF82nP0y0ZI40khRlq3iXwuJ+KKmE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
IEbKhgZ7VOQ+dwBBHPku4/YRCEVKMVub5bmueYcdYjwgMnoc2g1KULu6TGCYtCaI94H8UPgSb3EW
eGN1itlz88M3L8q9WbgOKPUFVw99Tm3GVXSZU4V//Tb3QNdRH2qrY44uVLGbQ9mkYa2ERKwqoni6
qANoEZUfHxRnSTKYHChNBV/UsC87ocUqgrD3ATONfa7G26nRSdDnwQ79x8H0hADuMPRMaVF1ORYy
QrymCRD3KbNoEIz++n1AnqIkdNeVxBKNy4nSMtNKEgeUcQVzM1r069GXDmTa2LsYlArLc5Pu02/5
yuG/SAj9ujBkI1lTy1m2KVVuPChGjilWGHTkAw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="//HuwZPNHbgbEQYIJEhWHcJDA79RbcLebyOa0zct/pU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4512)
`protect data_block
NNOXknLHx5a2SEZb4SLivdaHfD7X960pbTxw2XLtTI0kHOh6jNvkHbFzluRZmQ9VhWKZQbJ/rcn8
Bir/7iVu+HxHslGkGnx7IzcuTd6SWXamqLqW2HFJE9Hl0jZ4dwigB0/JkoCkQ0zYyrkfVDR3cyv3
mxTZ06Ss8sLfBcPtqwtTKCnvruQn48c8CYG4OoyULOxbH62QxsKDcMZ5Tyvlkrvz2BZf0Ookf9fD
qC45UjtnaQ8PlpN4kYGEt+WbYWEjyAxk7VCmkzhU+V2722ns/NL/p/jwNhA0Mi9W7zxi82vo0rQJ
OcxLDRuKzT/0Te3daxLVsBv6O9Xix7gochArVsJIMCIHg3+Z49iVXn6qZ/Sj1Pws3po+xd0PU6S6
gPVageks9ccuHp4xRZ/gqsra0phgSJLCHgO9/4h6leePTjVKW48M+B/Y5azpDBFk8FgqnnHH2stt
YmvQIc8c1I8rdjuEvXTwGT0Vkp9VVc3vE+K2ldL/HdMJr+Cu9Zlobux4ahudPlp9cuGsDFiCbqn4
LjvM9kN2ZOwYDdMz4EWtUFPB6fZlqUlN7mOLjlmeNcQTC6U2CyXLIQraog+3lVn+IDn5anXp5aJO
M5+SWRG7hJcjT4BjeEtZGN+zwJIbkMxyiQjq9nRjCiXGwVyQqMmmo5GlaowpVZrJTjHPczcYxix+
3jYezdHqzLDg2eFNcgWUmAF1J4ZUdeuJYXQBSB/RgKfYHgKFwBlPi7QPAomUGUB8o+1WJhVdjsoa
YHse1kG/zphgJr2dHDwL2Xa3k/p1yfLuNrlQCbN2JJepOhMAW8Z5n73x6K6gHdzzfiibnIp1CoWf
N8BgDBM496+NuPb0LUFev75tr013jn1axJsIXLgwzarc+vYzW6wWCrzdC2ixKJndfmYsGYB0P6O5
gX/YZ6MHJbRFt6HC349aZa/NFrY4V43UYMevnuGtEPT1MrrDizEt0tSLSMBt8wSVnkz1pe7OGrmN
VbBkQ9zcuLLczslH8PudtFCab96TMwWzKq7scalu7Io4Sa88zWdLMpsQHP3dputHZbeTzGg+n20Y
5ocLLNy/Kd579LNzm14zrXrDBWa1XYS3HBmS550SVkF1n3PZzRxlRA/Qz/4SuT2JRtNNwkrXEViP
sQ7Y5ihci1nwbVznvuEn6qYYHnq9Kz4Hidp4IgutT8/da0LaBz7k1YxSOiIGwd/oeXeesHPd4xkr
ia+RSC8jjXXi159a0bavf3QEyF8xEj04boXva+70/B7CsWS/lDpfFhgmqr/2jOyNHfxCL3XxxYy9
JuMmCG1lANYYFaBECJMzFBhDu4NYTGnLoZn3wkTEYMSOdMjigrUsdzDr+vut04Einv9EFmZhWBkp
rIJBgjpnfifU2XcDfcerZn/SC0+t0wawEY+TjYzjS/3CYPSmgxMvSgiTaW3DNvTjmagdADp0PqB7
kWmU7lOnVQEKpRhPsdC8thoBpzyP3Hm0VsNTZ3RdK0kJLgzUZGAuoxF/i2kXZqbewNKLTF7BYIKm
GWZ1Dgdq45QVKzvd34Bccdz7EMbqdfjipmS12Yq+bUvAZEJ8sGIoC15WuDAN1o1UErL+AcbQueSc
gUtJT81QPJuEMZ0i5th4EiZGw3PTWmZlBc8n25XaLAvjynj4h/v+mRw0P2nMDRkZjV4n/tCh1E6o
AdGh9wZ0EXlTpVZUrXNxHDTYMcCSNR144fP62DkzXDfojl8YrdTM6o0hVqykY6RfsH8u30WmWjEZ
KpSUJypWF8XLceKUfj5vP23FJhg6mFrz7Wz+tcUWeZ6bdPCj+celTMX1ZkK4LUygRRAQ52TjtaRp
ZKDud1RS4DPN6aFkrS2QZ/PgY0jk/jwr7UPgnYiODxvFvoXLaJkk6h3qLiGNU8i1TUK+4QHkKsUT
wXEbVCPCAdWW5Un0JJuw2JpM/dB5dWq82QZF+MBcUJrad1mBXrvk3PTm50QrfVHy7zgwA3CV/KD4
o2EJ9U8OsMm5niZ371xvkse+NyRmJTh9eCLx6XOf98UPAvflNtWE6grRGDa//2kHQUOBeHfdtVcl
kB2jWRatZaGCHndrZAJrSw2ZaJSEV/4GgczbxXTYNEhv2irR+43YhhpqJg6rpqUv0G2G+7God5Eg
B7ffqdLWvU+Wmcf6Mm09QV+KeEz1I+XK+sBEq3XzuRGs+h2BdX2Ya3kLtB9HxFpb/yrs4qZyrYCP
slbL9GfzK8eWji9n1ZnbpwLa2OUbIGNUCqbFjAPqsed1vMI3To4e9Hrxju9iLiEaASsB+h1QTmaC
4w3bGcpAFuIdMuux8RnH22h0S5cNze7fbPdapEynoJ3Gc4HDSI3KMTtyHgJKMq1pk9thPfMg1gdS
yz1V6q3UD8Sz8hFx+theng3frJqEf4l89ePNafY4Df5vQP90SIPStAtyD7V4SMGoIfgoQ4adKwr/
Vs2+i4fpnkzdbWUN1ep/EEGGa0MQQD/Golq2WuF+hckW1+cVcCfZPsMJrb8rHsDkE/rVKhac+VwH
49T4Y8gwxq2na6QmI7R7vaIiiTaos4QOZeF8jy0BtlmVMRSw5gVBPPp3042yXkM9+5MEmYG0emyX
zwtnU8yGxlUXAp6acNTZnERxXaUla3x8wCHDAKOoJ+F4a5X9YjOjZbpJI0Z3vTQZ0VR9LCSouPun
iJdtovhTT/ThZyiTWt47KT9nAuby8KS9U/KYzWnJpfsp+RfxE+q/RIuVLVqai2I7hrCkorOxd49S
jUhpNiwWb+GweW+ktUD4KKUHYA54uip4ltc0hVBsRSDKhVX230d3Wj5McDSb5Bua4ovicvXxobtP
Ertn6UfmJ1gRxcfifv0jny3dwrQ5ACNoEO7H+URH9lPjB5DTIu1gfAg/3waT9+UH4TenvMn3+7oL
7iHDwAXRItsixRV+9KqJTnSJaVWeXRhQd7mjLLCa3BVYxsCJF8YoV1XdKVAqmhhSqMIS0lr/jQrA
QeZPoOlp0FsK2IJAfW2Aw220VHlkWl94RsefeAWLaThlXqRhny6SyrB0RUAw2A/wzuIEyMFOnXGG
CRhKuutEUH+0gE+TFRoY71ugjrYRt9OpaedrnayVL/dSDZJrPu0zKUjkpTF2YrPwK1N7E4XRWAyj
5mfwPKaKrMifF4EcItW/WL4vxgYcDVzzsqeeSV0y9/v0wBP+8IbwhMq8QUJ9jTwC7terGsKdB+vL
bf62o7Vl+cBPeZk9+DiCvTPtTtYmN0Q83NvskBZTgnVUCvAS7jK9J7nW50O9gdps9ZqsCHFqEupM
JXebhOXRT1lzeBd1rn9T8dn9waQXu33nziRAyhBSPEPIHdd9YganL5xv4tTOKmQ2rOU/VDWX9XhL
wqQIjk2tKzHztF/hmn1Xt2JctJWV+WpyhTo2U76DbW6M61nJHJrxnW5uDSskI3ACGKqGLFgCF1AF
FrWdQ07w3Rgqh81FUiL6IG02pK0Dsnli2MjgNrQVAvP4RNhM+dyF+AKzHFuN6hhsuRhufMQ9Sl0+
2rR2Efb1fkPm50mRZkGDvgQ/86EByJjCd2wQRMK/OAIXkh/FGRM5t0ZwbboFUXzrnXcxvNcjId8C
NMHgOrdurrQRWKqZaGvgqazKlcGgkGNP2AyRpzTkXuv1DfgLPLFkv0VTyE3uZB+n7iNhvR+nkTzN
izOaz65z7mRyA17f+fa0FvQ+PKKwqGZMbnt0K8AoJ7l6725QfeUg1ysvgxKWw8BP+awZaHUHBqOa
Ji9+1ZGq/QDQweKD5TSH7G4D6rxxx3vs3lnsg+DbVVzqXyMuJYSDpW5VtsWfWQheLdep3mlmtEWH
Vwnb81k4hKxAKzUJNH6I1unAK9GH25kNa2rSmvrdqJwNDxEZdpUfnSfmNGRDH/tGKsOmRxs2bYj5
N2N0lh9VLO2gG4L3BK5wFOM2OHgMGm9eQX4RTyGdp20qINnycKQGQPS4NeJPs5i5UhgqZ+xKiC1u
ASSxRPsAmg7zC0SOD8KXDy3pHo46CsQ0lU2yCLc4DRmsn9AZaneMIbHWE0B1lMWzSoBN1bL/nEXO
UxedJ0tsW3IhNTlBPTwxaTx/4SQPy2eJTinLW13DSd4EtiDg5BEep1wy6TFvhhLU7/HpEp7Bh6Vc
RSpCsdVGvA7SMwiWvadPuBZAhBEMu1DkpcFoCc1GDfZrDow8c1oFpXX7s1PZiZTtK6qNDBllBAj1
qbPxfQ/8+zNZ1RKN+VQaKaP/jHTBgQl6IsafMGeWUCVNwCJmnkvH0UxGwnLFTYDYP0zPaEY3C+dG
pM7K2gsOEjdiHKujyOxrrVe1fAUiSgeNoCNZolu0z7Nbj3NA7H45x+psIgFEy4QJJ6DZJV+q/4he
Jv408uXD7WZcFJr3aIU4F6u9QyoA4RYgKn9cM+473o/X2ldgTikWeD6/RkWWX5XZTidR1lTUHm0E
zbzMnvZd44ghECooaBOOf2++G1awbvY4DVtyQPJuQp0pT1okACqzU6TbM6/gFQFSbenBx47gXeZy
Ip6hLvGrHAqBnVKxGsH7ILst9P8ImzZvpqDqT32N0i6BZcMXStC0vHkP6utvUevs4No7DLJDBfmf
8JlZzN2XvAD/xDX0609XSB2VfSJwl/brrpBSOOZeyqEvYvR63CePpaJTzNxBxH4X95NdQYVvzV8w
XLiEZ42iJi2JHYNpO5hmYh5QFc59x/KyBm202C/TQhQqzipCQyjVsHBmWcnSq8G99sxdzr7U3j6m
ZlaiTzPfWr4vKy4c+a+TONC6eo1X6gFPSv8fKgG9HJNNtHuOFK94IMUDkory1mh1uNKJkpzez/wU
EYhGvciHqUTNHBiMb7RyjMOzghnZ2dFIUj4iustyTcDrXAXlRQvNAXKD7fm0LicPJTYksNadLx+w
4I4yQ6fVH9O5l9y6ZJa3Q6O5u6QQ8Pwlkx8XCaGNZHrynrGDUoYOscLtV7yROILYU0+yMFiD+m+y
tiV0vWg7xufMf83vGyD786bcfZsuHlg0dZVvlc2hf0M3mNznApOJolxqYMtfnj/dK5cSEI/ksRK/
vAWdLgC287lf6bOd9IW3WHS7d0zprOYRsny6CPQq+nTJDvYfBBIkWWQ89H5NuYjr1o2wDarAV6h/
kd3iEorDgaCLqZ660ILHSOgcrPlURQhvheDTWmzetV3B8sVMxcb46wumziU20fPFFtPRXXOMsati
4Cyw6l9s2fCKM2OWArC0hRRjt0CMMECAYUn/V8rZsZwMMikKTGB0JO6MGdekDqYCFBnjTSZaFesS
7dEUetBlqtGuLCrY4UkavBiTYa6ngLCGmuqn1u9IR2/OsrQtduaZ8tpU8Y2x24e6VUHLHlAiuy2A
6YqvAjXb/ZxsH1viAIgdP0++KUyR2Ocg8ZHCjWBlyzppLFMR8uFeKT/nfnsOfejurHzvAw35OsQv
RDr5kDF8aL9nN2+h9RMIVc70p04o4fyMU84YdyZzhFbu5EGQ/vrVR0XeechNzWcEy7i0YOhUCCrG
K7B6iPWFi26PUbSAhX5Z5ke8Bgq5Qpru4+tmxSwQyfPkJXWA5jB5zKnzdjMKrK6dv63ZeIvo3Yg+
MKQNJzoJhIkvUjfyCboO1WIPakpQ5siqjX1uG0aWQISodO4lvKb1+ZQgITWb6QHMmcEc94lMk2gB
vAe0D3AVKOv3thvo8Ye2Fpp6keoMuM0zNaa4GPlu83UeR6Qe1EoC5dTwGbN4+13NAFqiBaWumAhj
Zqdsnocwrkt9TOZod5v6sjC+xLb7Q9wzaTzXW4EER2eFMApjYrOCF+LcAk6kfDS4GIAeqgrH38fc
PFA0gi2ky45mCGrNYnj9l59SS4kQVZ9xp+rYIQvokW51RfNDqxsbGv8pG6jXacVQ0ptDqJnTlRFR
6Phz1MIGSo+DiFtRB4IiRX+7NbNdTeEUDBL2HCYyluCiVR2J1uwfCP7XOssci9bsrAqPzzuFAeea
5Qw6jR6t3rgMjHfadYC+sTAu+YokXAQarLhgikTM9zKSV5QITpQat3CKM5kosl+TMY+pbxUjUWJV
PkhVl1e6hDFX
`protect end_protected
