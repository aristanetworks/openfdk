--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
iucYP2l2zh1kinqD5eSYX3JXZrF8Xxf31NUCqlnNTHaCbocmKC4eF4PdtD9HttizBO4J37UsCxHo
8qsDwbXNgN/cbq2fZgl8noMEwoy+0bQSabY5IfiVgsXF0uklkRgiaHP9n9gxoEysfsIZS0Pd9sr2
KPsCKoyucujQA/3yh5UlTjqEa5h4og61iWwk1CF0HcAHEYtTOEJLkW1nNRgwmLvtaqtNFEAGUjgI
CGR5JcF3dZFRIEpRKI43WlBDeE/0zrFFrhipSFjoNZDiaiGK4imTP7mtgrMJsR1M1SjxxuBGptEP
S7UblbAXxVcEzvM166BYkjcMIjzxkFWAtIc2BQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="+23tTkZ6r34eQKLh8JdhotqiG7EiJqZ9jd1aNOXPEE0="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
fwf5jZgCjAETnaVEZ7xCviOH3uJ7eyFzahRFej8fW4ZP5zG7lTjJ+IkZfYHlykyrM76XujelubZI
J0r/bN7xqKRFqN3NM97WUYSbbizYBIv/tTrkEtouaf4rxCQ2KVc78iPDN6mmuKvo1RHlaz6uJGnL
6Ivlh9dtkGH69GtjMqtau1m1YGOtIYK2B/BXxw35iSLn2mAKu7o++W7ztojh9/WTxv5mMccN90NN
fKUeJ1J+gsNzZ/6Y4J2sjv3byey9cbUijq1CzLdeVFAwOCFe3ugHuXxzZssALm3lHm8M9iYc+ctM
ZunuKVIUOyYRzxAEc3AWj7KxidmtziLLtHZVPQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="gRrkwJzbSpHLV65pW6pJRNxdQGEujWQqyhGUlZwmlPQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2512)
`protect data_block
eDXOHNJiVm7boR7QZR/hWvWXx7F1njcMtoVIb2Eh9hYL2m/1Ods5VWE8abURO3pdwGRl4qMq2y9z
AxHOrCA8lF3KuhW2oIbNonYFgDacZQbsCaOa8a3rcIsq5br3lvjo3HuaoDLosWly200MQYTqaO/l
4xZPcyxlxtTIb8tIk1xpNNeTopghWbJqGVVFRVXNljo8EURa3Cw+3BKicduHERxcYy1Rz/eRbnYV
q5+YPqdo5wKpWENTqMbqUjS/LszEEUiDcUTGJlMa3OfQCSt5rex/n4TNydu3wiqGOISZKQGcROXk
SUmykN1awfLrTa8NVSQ9S9GMMCDBDIuYrPVpulNlTg1+n1mS+KKw1FTcXvwE2UNigostGTSPR6Kx
IlpUODOOpw49Y9xsKIqB+dGm5faWS9aKa8WMlNPVWVfM80j+4+f5bUEe48+suX3gvchiE5u0WJ5k
M+Zeeeou+VbLvhKMZTEXAq9SDOgngmtlWBBVFtwy2jEyeDLBef9EgBBcNldzx8VOd0iKRYR01XbW
U65fi1JWTumyk7nTOkL7YM5MgfykzjIOwqkxF4nFMay6k+PpH2/3/0uTDZFzuqOwdEDg8WZJg1l3
vKIoOBbb4OlcShZuRWGmfbP82WErfd3FwiLVBBnD9YXe5BJtViecCGQrp5tpa4YbdufCzT9E6Ktd
w46kiydYLmKiIq/Lul3mr/D8uXtb53bslJEObMgBs+8yJ5jqB37X+O/W7Fh1FUMYNzUKBqxm9f0x
ckY4xovSgiDnxnUUuRQuURIiyc4axb4vRuANmHWtL48BvZBDJzF4SDE5araksrHPtg6y9hCsjIpZ
ebpt1DWwEhO6HKY9Nj58lQxNkwc8ydzb8X9A33nu+aptT4fN5kuOuHP3AGswy9Y6/khPHoIhCYkz
dtkRm+JiBUqivPcdNBKQxhFH/kxDiyVmew4pl5zUx/2Qg8zV3QxTlLUvepaHLnBwqUyfOMqQZfW2
9OrqqGV9F9ZPeMpi9kbasLPwyKGp24G9mo2rETdB0Y+M5CG7VZ17vFaPuBeXJjxpbvb/gwRmgLUp
WRqdZaw0itFBem3YNp1y3ejT1sxh5Zc8ZcleqnOVqBaIRuZ9voUk2b3zpfqh0Y3mMeMcNho8FsKm
83MsoUdjgQW/Ralqk72VqZQ6te3hfL1RYDGaT3msZgL+/l3lGG4r5WkfKOnfBkT/dM/z6T7fpxjr
xuHja/oIdroc3DZg5P95Rlq/s5IXDU3Zud9iqgi2cJRjOAHsdIhPjGuOExH418OBFvmOC3K/dgoq
aFDfe2gzMcnk91Pnk7mReb5YdMewxzGfKyja0RMZ4plOvt2+f5HxckfoNFYR6/obLCzfYPbJy5B6
Rv664bjjAqA0dpK69VbeAAD2Su2Ox5PYNxKzBNL1LDEY5itae48d726D2kOqx4HpbSCewNp7aDtA
pv29tc5errEg8yZrFTjtGhEwh6w8SyyqJtzQ4PPr9K06HNM5WP4aShQNI6AQO3nD8j5Lzd4y30DZ
NjqcB3BQHJ8eHf8b6UsnuDTOjI+iuRBMm58r0O+5FZO/1VFiddfWgdNNuAL+7Qv6uKsju9AHer7M
wM+Q4IEFMu+4gpk38cIJCG1/A1xhDFrgnnr2ngQ5LhLKuKVqS1oxUvqFSzTMrmHRsEAsHHX4ox0g
3oqYzBFk9xiKI3oNtbpB/ThgoJdUd3xZTiWTSZvXZg7VhFj9qV04SGa+B18t/8eYrG1kfqb3y82l
tEdsVffDuOqBRUQvwc9XhAtN2wb2EOxhd2rzMW6wWCbM+v8w1aCToxYBuo8cVlwouAbx5UL9Tjy2
Q/7eSXuhA2WFx9UtmMyeA+PEKVlvOr9wAY/w06gh8o9mCGoL4LBJ9lLRnK1idDcZZRbZF9hX7aj4
Y7Q0+kJ64ZOQBFyG/0xtkDGcuvvfK7OqXDGUQhwTTZxISLoGBC8FUuLmyquifp1ohYdz7rW4Ruf/
mNQ1mlCvzrSgYWdov/6fyKGQpOqw2o6UgkVDMLEEfP5OwhI61UlUxh8DaDrhhlDq0oYIO4oIREyF
onKJkiGhpGBueHKTKr8ov04vP/bV0Z/vkgTvGyJIlgM8oxrg9Q5732aC33Pg0jLCV2pq94LVV2tC
hXC7SI6Bq2UvUBl8KWcM6Y5n+1E4fXnGQg4naJVrxpTf1PZSN0ezri1iViIxJsEZjnwmE8UFYxMA
+nm1PgyZflgxbjHsRlJg1/II/ceR9MAfm2VamV6Esiv/l2wRtgR77WBsbKv8ub/OQek+xaMgDoqP
WSovDRUgFhYf7mBZqJkoH02Xut2HD9jqwUcz1447MHdSVmJxy6KuhcSPZwsOUlbw+ZLp6wyyS3FX
6KnYK12wwj9Sr031AKBnQ2IUWLd8gcq98IHWgrlEWEs8XOXwcLbytMjLn+AW/mDkZ+UoXLYP6JH5
ZkA2/Mh+UIae0oCvwxoA5LhaKMRwiULTnn0jGuoqmhQd9/s1Qms0vkWD54ko5nCOnv2AAmcEYY7v
F+y3nSSREiU5AMl5mW0NSJ06pHkj6+SYWIsO15VxhxRpwlsQX8juCsMGlZU0jGZ3ZSYlw2ZK1tRh
eqI19VBQwhhhygM544FxxM4hMPeYlV0q6SRO9tUsYMhTGLKK1Mj7aZkfXEEx0rf5Gl4cWcyxjdb9
zJX1LccQm1PUqnu5PXxCWCQite9+0I3ZsP6LUjwqb4mnSYfkO+oqJYeNY2rG/7QO59pxh9Xgnc5j
5lthLDKAXJrPq7Zg89U1wcPlJfDAHpsukpTtIAgwQ6yp1Izm4UysTa4IYkt7ecF5hlZAsPuusXIV
FwUnnIACzERKImmpJ8TTVad/SLaT5f4apsSZZDw8MlrBY9S5OAiu15LjqIBI7NN9nMapzuwtRgP6
zyzsfHHlkVsIktsanO41JlwEvWz+7bCg5/B2qaIuImnSSAEqL6L4C/MaOP8pYRTgM7UwJWxVkx8c
rQmPJ6vE9l5NbUR+03He8pxnKQeMzK+I3+JafOMn0WaJHeU3K399aF6JOJ6qSxIwAC64F4ztkyqk
cxf6yb5y5ELJVVflcBFcaejM36a9QzwXsSRB3BOVBcTgQQNkamJGxqsDGdvnbG7H/gCm20avlXz2
jBtIhRfv9SE7hRzLI6i6rMHXDxQ9/3wTYhBqTDMM+Pt5Lp4sxrisljJ5nXcW4Vfnvmyp/CIYGzhc
v65fMAov0AB0ioda67Xg2Y+G1jTan8nf5B26/a5Ry5Jkipmh0zjIj3bComEFzyCv37ixnwq/Qirv
H6lo8wPKzAsR/kcS8/IeVDuGAF6/Vryprr5QuHl5P6fxIlU0NLYLxqJ+gLLzUwsyki3kI4KjbcIE
M874aQ==
`protect end_protected
