--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
WU0Sghsar1J1rCEF7R1mlZ7+TCMzZI+ss8BzzXRJCOcrmAldB/X+yN0y/wUP8WNie3b+N5CzYxC4
S2PdxQBL4DFm0nte07ASFNWHXMXKRwbjPy626JPwT7Tf/n7bMp6ZEautO9J4KhQ+2gs5AhIz3A0G
MUDFwyWlQT3ytAT8NEte3g6fzazcnaLDPs4l+D+/m3w5f+cmNvEwlSZ+CCi/R7m/XjK8WhlZsQsa
MhUPQQ5gi10wtAPz/0W2406JbvCuIBehYzykXzeQJbwKvmjf/jH8wW81djcmmtYHwvqG+WdO8E8Q
0aBxKUFy1BSABo4MwzkUlhxf3b/nXRsyw+UyRw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="w4WTXo36BlGahsRX4ZCpVJfzdWYivJxLmwlBEqYY8+4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
hapAsaWFmxC3k+rrSz1Y1NU7ZFAMn0dUjqAjdJxt1G+t0E2mL0FB3rTUtdtcGnfXU6HKxhapAnCF
NWnutjAdeLTPvJOCqvFkgLvsSXnr8uq4Nmv1J/r84cDAKTKs94fUDgvsZrWAtQ05Wf9QQTLId3RU
9xS9Hb3s8q55Nqd29Lnm0wQm3QWUH0JMC5LuIt488R99P+je/mhCOCxYm4L37O7Av9cV8B9XcE6B
GxgYGS0nPZtPDgWQQueqxVsfXSOtx7OTXFt5NI09jr3e69TT73bPYCV2KUDR2BrDZPNgQBwdZMZq
dd1VWqZwM4WZWFNWh7V2pTN0NjG7RdieaQV+sQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="/Up6kQCGIRfumEJ1Ax1C+NI9z6+1TXo4RYPoAxDLWdU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 38816)
`protect data_block
rk9Ut9imGHukTq57IMIP7z1nUWLaMYO5icNp757HrLc7yO2MHw85gqkHLYaPrxk22K6BtOi3m3Z+
lge5e3Eq3fPptbmtuI0Z/N2yrvXsQ4LcnrdPUcjJRN5oQVcNJs3TU//4q/1XmYAMC1wFP1DdKyyc
H76lTsBzGl6Vp5GW5A9DFiUI5g9Q056uWWTXU4Dn+XC1KC/iYDQRAE4lBh1VQayRXoh8vCBLQB0U
orz8mgslXe3SlQbZyiSmd+PrVqSbsfd60H+fggnbrGYuoJkPjAvHmEVgAWL2ttVr5DwLo8poDjcY
GGenOLM4TDg6eJ0lAWZFqlSFb+9FQhTbkp4UwYUXbEsQQXyCvPFb9xGOaHoYeFyAk0x0odASyRl8
rxwEO3sF6u8qO/nWCd3OjsyCrNcaM5gJQnIo7PDM8ihLc/AWMDICd+j9g0WRRFXVY3YxlRwSuZGx
bTx/2PjcPAt3KHM5qyux3WftxF2SGKIUws2rORh0v6vxeWLLJFHZbI66COBq9fspFT/ByYs1FHiG
qiowQYnKsf9NWdrQHjZ7uBfPQ0YxCipoj+akGvUlTHDQuta6NhcOjMDd603H10GlvH/g7AwaI0yU
o4nrtv4mxHdTHU9ctTws/g2F3PPyTYq3cvxATnVWQnbmOZQRJttJZ4GXNPhK3zudDAaciuvxFSCA
wq3QDPG1evaIKOT9VuvtX+lvl8pmb2sHHpVp1uKG+1qmnXa9H38l+/u5wxYhiwLjnsoL4H7ioXjc
ZwGaQeK4gf+bCw7CG+8ezzDArj7fziUN0tY/vfiScMtkT1RryTJUxb3YXn2fY0DxDCzhFj+D8FiU
rjTrrvTMmARAvI5SpB4RI05dnCk3QzfnYshME0KCBCMhajrDrv42yY6R2ouTG6Ubn+StfnYzN6NU
zvm8eXeUoWLbfvuuQvWksthrHwrIb7RYK1mBWrKH5iytws+Wyj3X2tKLqEIopvFLukMh8o3gbKwk
tRNhG8dgiDOC7qIjA/AGeYm6/Lbr1lEBERWimALSiedEH9TwXDx9GnVl005jlmY46WfwRfX9JFoI
XV/EDqubElwkXkPZBiD/rK8ALD3sml280DJN3v+J/0s7C8OA/U+wEX1Tb3n9ORR1erCmWenFbgLM
KU2mnkuSGsuqqdAgyANdRm/tX74sZfckZSFgmZas2wTua/ix07DaAY32HnYCMemJfSgugubfKQDb
1Cgd5tYkPFGgl9vuzoTTLbZiSM4b6/Q9hOMWIZ6dVot3EhXEcZlxan+8yf2OiE77SNHzOtbLcY8x
kwGzDrJfKxR4ONPvAMEIVHserddf6Go6LVBLRCXvMNepwCBQrH7/76XCb4V5aDQbHLjEJhJKym6r
WU6YRHg2ZbWVveUX9sjKQKtEsG9imYn3g/khgdnsp3w5QXeZbLi9UubeTN0PrBh1IZyEKNmV8pR8
UcxjRb9AviQ7E9Yklg3K/84ItnQnUe8XoLGo6q54n+ZvH1qiJFLkZF8THlOLJq8GsCWbUB4c8YR6
uFQE3tJUO5cS7+MtTqD11B+zLRXPR+elx0i2OHsvWLdzqfEZZ/TR9tm6yiQzphDa9MJt/8uC6WiZ
R0ATk7xZRqnDXLbQ32qCg7eiPCfSkjmxzKLfpTe+/8MibXa3MG1HvwPoBiz5T6aYvrQivd1sOL0z
D94S5k0wCnCXDTkaKeXGzEYghOYOHyw2kCfIwp1+n5VSxjl6ra7MY9BT7+mrdTmjWdovwavn7Noy
YypBFKe5mVmUfaptOj/5CsOL+TZNEoHnYKkjK3q7e715kCqd1sgSKjqZPzVQVAlU1ocW1br4AUyj
Ti6pifmKJsFM2c84NgEsZtZYzqY/Cs5FQgGBoIy7PPPXI/RrbFAbzMOHO5cOVVovtZ/VyRonn9rK
30KjC/j/68k1jjvUggxc+5iaZKa7EUCldHzhze5scnZUD6c8jLpQ0R8PxEBukajkAAZAgKfwUQlW
EXjWq/IzyWajrBqB6DFXFodWVsFDd8gKduHFvBMjpXf5Bj94oKMajmvpbiKVi2ykkHlHUA7ZrKPm
FrQbu+0qIPWTV3/jckgS6oDxioOnGOsVgqRobj18yCcGNudINpRhVV6pQj/owWzh1hlgNDjJozuB
KyrJCdXJSPMLKEM7KuQ59HhC4MQ1mKAsgyr5vpr9S1GenBnlt6JvWY5gJql92EXe5fu62/bPr6el
eDsNUcpd8HP4vDy6bXtRsY2hKqI5ZysJoAdCQEudg5ySRKXgTMy1bOHWIdi3VvI6xWyZ2Inq49oH
zIDWXaZ/HHNW2nNDvp2g4C70/FaZKZhSBgAl6QK7sXx7dyseGoGdgM2ude1Ce34OxRlW7oO2BNoM
2XBU3iKH4ulzGxYxottctw20uie/H8r0ACfbwnchw/f86vTuegKqvAv053uGouvToz4aInWKflyd
+4B5kn6tE0/pDODH0qLeYEGvNn1bnxMX/g5w4M3+gXAEqzTUsGMgOHDCKT+MZKs4YmjaNy1PjC/y
X9Ou3Iwcmm5LfMr+y0Nap7SEGEc24gGVKSkFtK6efF/h83KCRShpebrGBkrybNp25NEidaEOMZOj
+YO3zOSa76rJHpHhoBQte5WIf90GzWRKi87j1bzQBwP5vrt/HnMDzKmVcuCCE4AEU763MerAO98X
lvU8bSD8xttrtSMEjBAAOBRbE1z1cIl5N4CteauAdxg9GioEVbR/B9PnxYerHAQiQTo4e5TWYWJJ
GzXmQrDXPFKPLjkHt3td077Oe4/ZfyMPKtb7HY1Rxoq8HyzuWzwx9KRK6ZYf18+clnB8KkS0VmLS
FQNByEJG0eBSnese7bTI7HRvkACKYV1FNOc6NpP6jX9ZHwIl4wgb0FSM1WuOqgfSN2CMlqzsqvkL
c0QVS7JG9DGKVJQBC9d2C46KKuI11tO8FYlU3qF1CrMelPwtC62pF/nE6AGfYd0pfSHkBLa3/QY8
HuoTBptXJYfeK/bxz2egBzgWJNP9PRixxCLnvqe2rtYjT92UzXFqXBEOPvVC0bdcuv/li9IKYHHW
zVFc4c+GQE/sI4xvKW6mwb/Uz0a+ueLfWnTjgePKKrtpg+b5g1ht+JgYbcA+BVvboknlTW9tYmfr
OVo+Zn+qrTlI4LfegDpeYLHVegO0Z2aYJJuxdqkQozPlvwf1vyd0jqCssCBTJyFLgYi4WqSsUeWI
2RDO3kyFdzLuQwnpDBNp1e+wbJiqEJEtdyUJw4y1nWvgd441uHKFO2kbKEvi+CyB6XDJ8xwHXpNG
zK7vSioKAHasaXAT/C+44Xg2YTudjctFGzOv2EAiGn/mU07PzyvjwtqHOp+VRnU/T/hqjuVXIaL8
9dgY8c2WNi0t7fdU3cANEfzhdzUlqQ5zVjJL0yAg4DjnB63XZElMvGSM97xYiG0DHd+i9/+EaeOT
hLFZiF+Dg7E7LJmUtWJVW3R3kiqyu+TwJ3U6gL/vNpqqdjUrBlk6rRPEyYuOVSutQuUYcEIW+YrT
Fp1KOuZLy3ZAj+qF03zk4+2q/u1XsebDro6ejPBApUJvhbgcx9JFAqVJTfYeXUfAT0P079lImKdw
XBfgKpiphmDgT2VzPaRzyU3ZyldrmuIlvexVTlIOZnzxGhlhWRGfpqb8khqkEA9KXkB96IDBs7ac
RwXFbfHRIkuWTvL1PkajLXilOomF2VyR23RrZ+0zosyTrUtxfZkf/SENe1pE1J/ALH6+oVe4WzAE
yx/e+2wyUhHr5ujyAlV3Vir+G0tMUTWsMtd18/+q8aY3i32d9FgjDQACwpZM2yUaWAD83rvpoJJS
MOILpwahtm6hbYUAG+Y7AH4ouKds+3Gi8CMtVaiWN8ZWbYMSJj/m7F0uWulFtv0EOtYvWIMTNEpR
vMCvKWedcULXHACcnGKpSx8YESe8k0BfBAaS8FL59ozzhbuvkaOccRLPZYYGkWWFN5vh3XfNeTVH
xHshGSuEhJhVaroQdjDw8m4tOC9NRapPDkc/aP3XZPN62c6rHfrMdQPZwEzT+nN+nP6xr9Ra9WcC
wVBPWwNArZ903VHI0K97s7SBso61+D6zNuKe19y+F6TscT8lW6TAjxtNEBa6DkoqVjSAj/zZqha8
lwe0bxyAt8HJNzc+HpSIbLCEpbIgV67rv1ypWXU2sleQfNgXGKzOTLJMNOmBxQmJI9hU9B2kUuf7
MUEi0RvtILOxGNlxLjLrYRZBAp0unKgPSw/fgjIMnU0j07SMGJlHP82jkYrktDumA2YUGkNJbJpB
rMwQAVCS4qUb935HQfR/2JzJB1vh3aMJwUF2Sut0+fVLXdtHYuli0xSO99c6vrPuyz/60Jqw2YE2
/TcIOK99n4uEMri0sru1x0JN3hZ+OYaOIPFc9ZoL7byI0HhfHmO8g6vo5dmoePSM/IZ3iMmKPbF1
Pm57zsrWeBMKOEm+Kgt1s9nr/+mtc403dNX7M/3kMw599dGttolskf7P9tSs64rQwpzxZMDMwB3q
+XN4k6UOBRkxPabaYpWDa4SrDmZqKaIM3G66WOb5LyZC8eg7Rn/S2J1vwnYmlNO2ocS44NnOW9LH
lqI9p5PmA+751RzjwqCyIFkRYkhpspFiGQPibhoyLfsVLXIpHvH5UhdrfIKvA5KgN3S3WvXEnUk1
sJgtxJLLX5lnvKpuFFedd0AG8vdh97fWEsGHl8rwxFL0GNsaQtQGqJltaEdOqGMzr/4a3BBcV6bI
cdfcH7TDwNtGMb1BzL6CXQm7dSsKa+KfBGorIQDI/hr+BVeTOTdwneCQrg77Qkij+nPKjuGowdbe
Z0WLNBV+pKKUldMGthTp2N9RLrR5hS2hU/NHhmCsn9eNOUdQNi/vYqSMIrrbjQnv7Uh7epFs7Gxr
ZTLiwm1aW+jvzcKvwEDUM9kpW7Z9dGzrdePyUn2dzc162ET/uf0ttnm7nfAa2WXp0kABf1fEwq3v
IIIaRQaOJhDjFraR7WRYDB0PGW0HDbiVARFVShC3OLwxL8tHsOVD7Spkjc7uhuw8Osiw+xQEIYei
cxjd7vsshC+jryNeJJPUyjhvesCkbMHXViRFSNQOvj/SsP25LjYxpCarRc9G7riGD7ZwSRhOTExd
nNM+3ocPL6eN5sCckl04qwMtwHtLvpbhdFUqDm4oqU/Pe25zLBp2PO3JW+ErMAmRGDRb+X6xC/UL
cEwzJolEUy6Fyw7b+01KAYxw6DHciojecPmkWVM3AjY9Zw06kXHYctmA83p9TUr7/8Q6N7Z/Nrlo
OUZnDf0A0mqLFjE1vwqeVGQs41AhWnwapfs/xb/3ADM0MFrgLp8kuf4cgxPS3jU7cWgkEmoPEUmT
78r7qxeC8L5VbOD4eEerQA7Vc/PFNOmnoveJO1mut2/dtYsWrygkaLM9t16ec7o4MrRCNUmJMIYA
/u5YqaI884u3mK31pZ5Wj30Grgu5tsQFJ4fOi/9K+YRnma1gsSq+q+EO4UIfXGUpebikcWageWbl
Ad70tqd1PmeVRWKtVZT+tsFdVFuFe583/rbxROdlH+Sn1vudSgK8MiiJT3p1j4j9bYjs+KVtqTZk
skf+LHNJ2u+SoDcick7+yffooS1qbisl7pS7TiEqX0nW7q0warsIj5s51gUfRjeVmEyv7pupfrMi
FVyF9iadkCrA2AvKaZr/7VPCh9xTmJYb/s/HPeflN09vXONzaL/2RK5SZJo4Y61bfpaGPEekHEjI
zBFqVueW1u5SWNujbdzYIZYP0mfmUZrmejIFBNCddqvgTSHv/EM5dhsyBR9d0hV3y9FLGHRkvvSb
yAV+Uup6KuOwWF42yWK9I1piWFewd5WEZlpWCSygpsOS8tgwOGM16ZLh3PRHThFzDaagXZVhqlKL
6tFCWhEml68GVNeCbHrMWtPmVgYfbnGa5uvwFEPnP+t3KrVwDWSVbX/KGlW6mnGYrAZjUfQutnQw
CvcK6rkhkrqpqz+iKFgmezOHqN8USEida+h2kgnxP8Sn68neufMSWjMFXAxPd2W6jX4oAkXWOixZ
EASf0bR7aNdee405mQzDf1Yv4Ucc0B5wnDFfeP3F4K5Jhg91ynKpGXZ4sALxQ8HWrZquuUCE2QcY
Sr11V0L2OnlBREhOqphYdgiBQsrDF1OaD6bdg9yCBx2K+pRBOcgwOzjDbhh3HaYUappz8TUeaYo7
y9GFBXtsWt5muKnmT97GWc5ykPlm2yv7kwR5YJ718iBxI3ugay33S5fawUbttGJERyrajruZ8Eu8
oTdtornVsBFKzIri8E1xDwZpHVLRWt8odu1pHM52V1DNRM/ti6Ap46XE5g5U8rM/9ZmY9AKYxu52
NurDwr8Fjuvllev0YoGYP3xfMBbpbbl2kFfXMfm2WKFhrvPHe4O9frYOnU0x6cQmOm1iVDklfMpm
eDf9KFzLsIu6RtuUWca3nghSXofgs/Qyiap30A7MHEyAAX2OxZWe+t1TLocYI2ZIvmQOUBLdwQXu
eckc9RVC4FxfkKJxJ5QKatLNjjeyZxJb/gl5tMkbJHB9ZulL6vvoBlFRj9ioG7k2oNjSeKz9Yw+D
44EyXCRj2Uk41+iECVKEH6jxQxlxRhkou2PAsgTE3ildsB23AE2GcKFPyvvn+/FAJ9uFfCn50kgF
kV+dbh/U4iRtQ8Xv+bNx254Y5lw+cV2kc7LzGv+6q305OIUmZ6UyonWgZn5oLYd1+WnK0iDwtbDj
JrKlwlgh0lvoo+bWaGxbShKVZIfdDrKhuf9rI7v9kPdJHfXXlactfJmc29+MKr5aEbIEXD4Z24ra
XMA6nb5+mX28v/SRvuvUAtMe28aBh8MJAME9VT0odR0ungVqvUOxLvqun2XBDeZhBTXtbBBiAbfK
IS9lFGv8Np+/f31QadYOp/DjyWyTgjkKYfrDAayoYLgitRNZcJZ5uLVqlugvGMHowrvq8W2hIulQ
iNroZEikY2APUAI7oFPqv2XVDYFRzRdmNMvKZ5k+P8/a7vSK0ubaNnkZAPtERciXkUEbCAPDKg5o
QAXdjTgQwgQ5krZ3u4QQIl+1yF8bMVTpbH1Sx1fKzue4adUafGL1XkG3qOoDqmJLxli0Mqlsp/D2
Nr0nZdork1KPn80fnQOiHOVrfrDAErGuazeT29k5b2ltbFVtE6RWtvdQvCJNkaH1kz37QJzHQpLA
tKXHzGEaaES4eEahp9S0l5xWsCd/L/P0gZLnch0LL5DpMHo+4IrL8OJGPGKIEL2zPPZ5yP+pjYdu
deg+zN3N2DGxRoiYx10ce6C2IsLM237d50gEGaPzDaVVANZe7T7X4CtDG6nopDZnNFZOn/7S7Sxl
oYvDVBkY1XzrmmR2Kc8A5G2I4nJRlA9W7eGaG+xlDGkPP/wifQs75X854UM4XZ+iQjNq6sIDL1RG
p73iduHHMjVR462agSPckezUxMeDDPXWIj71Z1O1gATJlCDMY+LbXmIAGZ1AlVGHO1KMX6nHCNwX
ZVab2n8+t6Vv0Mcda8MCY3sIMsDrHfvH532bkC9Sv07FpPyVt5AKbcdftG73kWaIgwfsy4uozth3
uAjQbOGgz8r3nc/kPU2Z+RGMkOd4twhavhBowi+NgEfUlM71FAzS2Q5kWOB4RqWEh/FfZPn2W5Oe
HQEfGAbyEZyUUIXyPNC8XtH+PYufWpLzGkBDmSFseXZNdmBI2jmv7VG2jwHbOwfkrm0WemaQHt0o
hvAjfN5SpCh4QLqpP+NDf7At/dReFlglTzzH+y58t05e3bInzGpUpzpqooqHqrq4UPt9ed12915n
t6GCK79+4ywMdj3IkMP/KozkbwMn+dDHRiipFEZ88bOY89c5nykS25frhGxY9X69kYKGShilrjzq
DpF0pP17HMvvG7uwEvgEkR3HwEApKcAuKh1t5s5vgsl3Smw+JaQHOb516aYHhXyTupcrlDpfQBuK
Fcjr0R/PcYyk3veSfLDxRr5x4749cl3L2eyMQMbt6tHf2nvw4GUSgtLAgOIW4nA+rgy3Xz0ttKvs
HZYBU2pTafusYgTMokF3+souy3qq2GCq/i6IwLRqeDz/DbL/zPkuOAWlnpJKp6/KItslP5i7HPsZ
gmuXpw1U6jz14OLAH5HYXNfHJ7rd8hy3LfPh1j4epg3YPqPpwEMYeWVWRs7UvKr3MryWS1WAYRNX
D9k6idt8Fz0yPJH6CNGosGfZ3x1J9LbcDWFW8ngpDobr7bQ18wH1p0NyrnC5Prqrpegu/ti35gzp
8OV0ksPZuiwzYGLZ06gE9YLsA3atiFR56S548xSi+IoaK3TdJgaN5Yn35cuY7hqF/sfCqAGPALXL
7J8b2FmZJ1+2DMWibyNwwZkhCOSMdImhjlvFRRACS65HHgARQx1cWRVEvKEzKMV0+NVLhXMHaW4S
WQV+0rGB7ovnIN9+JeeXMNDrtf2/OxEiyuoCqPffal5C5kHOyIY1Njv7Ar7rXzhQ9t9YYQ3uKsOT
j7lc5h1yshkPVo0k5OIsNxWSptzmkUjaXTKejldTFgD5MQiu2A1zNPtqOUvtr/O3WftcorvHOXQG
/XKgTB8IObcQXmHHVbGsVhBEPdA3ctGhL8mf0gpKJ09SHXYHEMXcrbwoo+y96PbEemn811pqJs1f
hpCg1uYRyCHtmaaRXFaBPuaXwp65Q8jacT8oLODGFGcvg1kq2kcIkb91fupPtvXxqD9MIQ0rf/Dq
p7HeuWDu9zMs5Rslz+qfCyIbFN3kRtJGnk1fHhcfdU2TtK6sS88VHoaf2FNTqrItECsrH0TKCr+F
4VRssE8FeAH4EDoJM8TFGh8q61C9ibSc7eAN8QStJ3QIJvJv2I8UWkIV6PIRzic7CZINiOG4m9yn
+r0cJFhURdsGRTh38FJG0yosgN4wbbFpnmo3YWBEq4xkisRiD4ZlxhOHxBiv9raYaloXohSBYVsW
9M7oxUsMg1rEQHEYZh3267KFkT8SZgn07yr/dP8fdfUhkaXBuXlrHYMqp8hlqF47eyeXTQogy1xJ
LKGkO3sYDCMGoKpfhmgHtjjaGp1WXXjkxqhBLwpFieVairZU+JIG/E8jMOOQIaMzXEv2sZGCOCS6
kvXZ3GILlV60Dsk6FnZ7zIUKaUNOZpidDpYMHwlBHkBQx+e1IRxO0vd6Bw77hrGtxw0DE4Ukk4Qk
lor2qKzrlS+7fsmeirJbPxDdmVjlpJqIES6x2oci2a1K1NhIzY+NOgLNgxuhWnLw9VPeTYuJHN1O
GXnUMy3Rwv0VoLGowpBsTfBgm2gVGBTWZpbueaFrQ4KsC5yPzE4rlavuWUP8t2nrzxG1NWNzqL2c
KYMv32u9670OofvkBiOAPaNVtGSmauVpWeP2oeiIsR11q+RNPhlyftcjR6aj4PiuF1GxCBFBQ9n8
dIKF0vPiTgdz9b7MTWZpPU8SBpRKcLx/FR9vvjV8SAdqm4UQsqTtBU+3wpc7WIHahfwiB6Kc+1Gp
Og9pQfacoTx91Ownh8eggLwVrfJYE3w+1QNiRQ13U8I33SJKMrH8KCdyv0aRvJh5VTtT4HawRqXa
1H2dyGvF4sz8KAwfyx1D9pFDrEuzgVHQMNc2yEvXXy2rTjizDAUKUCbXxjw7GgM2HJbLMHEkP4ZG
4w4e3TrZnKpePjA70r+9169vdYILWAZBPvk/I42Zs2KjWYxnFWao6XoJTxDkTuknBDfFTsvqNPDT
ThUcArjU5W4NjV4g1vhd4d9ZkhnZazu/yz+LhIEQkUbFbg7aS2TOCxYzmEPGlsoMYkTRlLXJPOBk
E+cC66+pLDm7qq9xlnXHDwX5RO54Q1IqDf2vHgw7CHQTj/E5PS51eku8fAbsO+N8ugHGoWZpqbTE
p/lXv2KK6MjxUqo7otgVCzP4XySBezB5S5CY7hUAdKxVKQhTKLQ86BVJY5M6j5ntz4MP1RW8LpIP
8bNCp0JLC7PVPqQUPpBGvH95+vBRpJmLrNRyKk/9e4C7AcmjDB/UqH/WtH5b5qzDyfUYUGI3JLxD
xomRUe8ntnzZKz3Lm2EuhFvZcO0o1BAjTxGMWG662PwWoT9BuEzZcLawlRp8QtSXtcwGXIsIJg8T
fhBMjbW5Ky3XngoHG5kWBN+/kHpl+MVyr5J7FPwZ2JUpy4qLYq6QqZZXEmTxHpJT4ykLBCjLIyc1
ochlVUWIJevn2l44Yo6e2dcC8zarr92LEMi591vJxGWQq3fpTGNc0KbYEkerooDS57W7cOjATOK/
qwA2h6qTtwxHfpfmM06UzwoWxszlTaB+YpAaqgXpbi8blIO3kJNnQruutwBjGOqPboCRSeFU/JJ+
Y+rWpzpb/6mL/B7i/yFhrefpmHbUMPGV1c0VsprJY+unLMqjGPfTo9wdQdeU3BK2rOoCgHch2ZAw
9XoqpyAMJ6Fp8LYHE4SlF0PLB1j2xZCfX6z8mm9heRrXmP9Wld6bhElrPPR66TQ34YtKCpLepgCt
SM9TNvBFHn33vShqj+uj0YxE/57B6DUvcw4ql6XI8frwyRjAD9mtpnDfLjJxB5By5l63Vrp7f/y3
zvUo8tOO9BfJt9O+zSd/sMfKv+73fPbM6k5vAgcgeMs8TBTxn9HytU+2s4G6mveaUjY+2AhYIP/0
1Vx543DvYA977/DzbTu6Q4Ihq/6j0U6IGGIQjmu8bHSluxkAWOVuFW95AJOIHq7D85aI4f+EZaBF
UorpSpcejfANv70bOSyIXtJ7wc1Lh67upkK/EAibc0WhL6DelpibDZCHCRMf2v71rXmAnFx0BvSV
2Lyb618/fGFpD9T6rQorGhXbWnVWsiRXntJ3R0Qzm/sa39xvjVAhdahnYyTjgrAmmsne1S2lBL1/
rAdNB4y3JB5WPY4pAnH95A27oDflRmeiPhLD/2dnBtm0Ty+S0WPEguRqrHs374cF4yc1lj/XPqCy
s/NCzOp8LdGl55hx4iWeCwE1hSEiDfGBvchMK2eITWMq9rw1phMW/X+zRIk5IwZxgO9VI/wTfoG+
+V09I77lEBR8acy61xt1hGsYpfYkBbTBQblgaPGNcoRvPn8eq2cZ7V4GNM00/dJmwUUdnFtRABfj
lqNV1LTtccduVylMIFsEW4Bs1jTNfssHjwki/i5qaxMiIEPZwBsIh7qslIFQO7R+ohpjfbKwEkkZ
jsGFtwax9IIQBklOBIGn4p498TCXj95yiYJF/rFsKZxChvxfu0B3H5CM0npLueyRzDH45CxUgLwn
9ez2xxXsfHkSrsut5YxjFoNtPFFgkPoDDXb4iewc9kaI64JVAO95AXuBgIpvPkvY3vP2ASPPREG3
FPSv5WIsT4EZxLjkz8eRbNOYMqXeoh2Zn3cIGflHe2J+fzpD2vhoVq1oCOQb8nxMxqUC5Z50xGRf
aG+CZ6EKeMw8fVU/X14tImlah1uMwdqTD7MXK5X4nLmspzXy7nEcwf1LihYhK56pkckDLnBwPZzW
R4NVGZrwrVTMOfRV/dUr8OD4OUE5hen90xypRHl4hjxttQbEM8Q5MgUuw4jaLhXzIxnx4CLp+0Zw
MmXnZF5mgdLg2TX2mgyOxh98jVa2O4TTh9aJ+PLzWuQi6mOalfskwK4cp6VqBZtmIZf1jxrIPwZH
66C3tnbwZwh2fN3wZ3nhgZp+WxV4BUCLmAidJDJ5GP78bVnX7D/PBEzQv7SfTbXUmvCEyMfYfHmf
DEhG/UvUS34C2/Aisv4uBr5vv9HiMCgJKuJttVE27/MQN1pgmSJIaBoIfsGFhokheWoChDbJpXOE
7TPD9ba0SDjaPdB+WdnwlsTZmntevon/l3dWwIgzKyG6JhHpbv6QQvyELho9ik4CJKWW9AM0IQ94
pfwP9EH/GcF8kVb//w0cho09zcENFHzsNFY25yxN3kB+UEXNxnYrIO/2vqmKLtMYVb64bspPvINF
Ujcn7LTxClQ8C0rxP+B0fePHERHMiSHbK1iryfSodH0BJv8m8DKUL6szONrZLFOCJ54KKwouoRKp
D3sMVgVf3M6X/G5Swgzx0khO/5MN6N4K+U4GwydjZTL+FzJotuEiv5odEjSG0N3YB5twUEMAFlWL
DS2kDaXb9b7bHKGkWg3Ywcmy6xaAN/DdHBrYVMQjTIq8o1fMFRQyyT7xHJWMHIXbYcHireUintYO
3Kpr4sEhwgcDzt+Q+cNFAPxKGeH815r87sTrmJ0jiJcblOVQx+9UHB8BVXMICKCTK8xI6Pf/gk+1
sFQSDhEZW4uLExTDIGwaHgxczlJkGpVUoZzTkKq0AATL0CizpjFvsEuJPX/OL9MBxR+GLpB/juLh
WA6fsq7zK/hP944G6VyidWV42XC8EDfucM/UuyD+AK1kJb83ExYizS3SujGEQFe98u5/yNH9qnOa
fGMPsNsVWZzZKwo6Dy0TvZShk4iJVVEpU55LThFdowX2O/KIExYJFjx/UTfl3oFwziRAyAwrvhBe
JvNDDgD5JaWiEaGZe5P9KWD4immpUpcTDQ7ktySNP4cMHXZqFR3oNCo9PNw3AubmEYaROahTDXtO
+VM3T5I0Ndl1GAql6NKx3VGzbUcKSShFzSdJafwrdP6p289Vqj7wiHez8I3zMN9x0SYatPGddNwT
+cHepN+ZVgi30mdzY5pXVnfaQFsRKi+DyBld9TfvaxvIujs+HdlBtzJ7WBAaJv3hw6x7mwhN/TmG
Z8yBosVkAYQZhaCc8cSCRPhnKwZQbJqwIUxum1JfkC60+Xuxt+wC2JbICm/JarV9djUgSuH3EZia
1m1Q0JCBJyKUAWqzmPzXuj/qgMgkRgCaddlKz7MTIohkRGnjrRKyOBv7sQf92KpujSuCyCW5FKoZ
fMixOvAbICit9f93dOc3C/AeCOsAoDQo1q68WGl2rZbo20beQw3G75HDzQ44MJ2EbgYa0m2aBfOl
472DSz1F3ITKKoNnF8LEMb/RFWn43KrCdlekIeWGG29DZlehf9yR6vwGxAwwCJ9DGlSD72yHQM8V
F4cgtOyBTkAadSLmMWHYYSLOerlRlelSwiUFrLsfCHpFbjVewKlmxfJ4rzKhuSysiFRr7fC/EP1y
1OQ6adjViHc8+yr0pLlJGeXNp2/9fKPBno3XJU9lcpdiRX7T8BsMOOZ3kgyj4wfh+9oZpmwoFB9w
hjDPVFTWyyqSjhRP355XNTumc1joxHEHS4/tSjO2c6IZyCEdqubkjkRh01CIwAAcPjXcZBVcEPpq
LYZr/4WJgLSYR34gMRPkOpbtNCj36PpPsg8UwH9Db3tnqfUixCi7zvOz7H6Ovkpz29GZ7uXgCc2a
bWcgnNCyBiZX1xBYjwlLdyIRgrpFbMWQaxLe52CNVPtD0cs3PClQgLaSeNNhsm67d3kefeFUEqvC
BIu6JsjeoMIZkUI8wHYoefm9PObnE8+HF6G43dHWNDH2xqskwmr27w5LqoBZhtnaKt9tqLPOalI9
QqjJd5ZC5aQue2DM9qbocKCsXLuGyPnRnG2+Ocg4absAQeHB1PTowROGMOEFpsSgbcgRx6fwx4tB
Cy8MuEMNFwgHbU0imlCAzIWNeyimrPtafXe7YrZXwZDsUAAioTl4+lw5DQDmjmkZd+/7DOk6FXjO
yjcx5GUknPKLyxdPFC7VsIbH41tEbDrMC/Dd7mW8+9fH9VMwE/AwSQ51xzF0gJaxtg2uLJCboHu+
krkyMxINtypxUPaOncOSLOk1lhrZMHwm+QGOLzR1xlah0ulpCZakHomOpU8nfw5OH2fV2aoj+lX2
phGiBn58z6ZQvhityvp6ebK/CYygW5pm3pOWSM+wLgmYtb4zUYxnt62IOMJjlFe+EFa3WC/Kc/o/
7XuJBpwwg2EHxnh9OnkKIwJ0fvV9DHhf3DFkv1y/OtBLdnC2TjOv2tf85xr76DP7j6FLFT7qsgsb
i0UoDj1kUK65BxuEqb4tXr7R9d8S/uyhB2vkKFLzMM4ENEXy0Zc9IZrdPsz7aT9WZ7h/cSVinNh+
yJGVVKrXygioKxBHLImXYC3rFMBRC34s2/Z12clAjTu+e/5NSmxufM1wwZlIOfbBnp4m17lmq+rP
XI5BHCRI2lCNdHmbT7utv4eTroWlKS01NQi7Mu9kX7ebSEXfKuH9aN278mwFDYV06xpOu4IROBtE
fUP7wVH++gHJUtOVJmUq+zZZe02M8z4kF8ytYPUoX6FmMy3DQilqAg5o/w4owTe1kP6y6YvTfZme
wY5bQYP9YEvN6mv4FAxPPRYmmHzHR79KneSJleurkhM3OszzknYc3d6q2/QOV45XumE3syaO6UUi
0KjrFK6WuhiNAa6bBf8yT/IkWnJnoZ5DQg9S525ZQO+zSJIBkafGJg8gtZR3DvgqaxJY+FYb5EZg
/qsF9qCPR7TKrBHL8bDQqSwhjauXZJKNERXR5A8cnVJZy/JdmiSYyDYnZByquaNh9u2X2MmBIvEC
DNhh5CP6L6+fLa2CFo9FfztiR3aWqmMkzifYuvCi4eH/BpORq5umczCuAep8bJhu32Z8tn8QCHa0
qOwtKNmdNwgusQRU3bIqcUVySlAzQ3BUyk5YYBEMybEE7tioUCb05HUM+QeiPnFtGzy9+oip+Nwg
XNEO6T8pPwkjPFGa5RyrB7nkBdz5yDmsoCljgMwOgTnwk3MAGXvJkhqHd1aDTfcNW7cdXLpEEWk9
p6wQgegvHfRV6yNIQopZnURbH13ZIeyOobQO9IHfp/VBOpFLnNRPPTMRiw8kQN3TgYbJYH247Zba
iOWSSXC76H95d4Gx+L91uV9Hh24LWdiXbdDTWOED338y5DKI6aXRAxPv3gyXrwRc0Ej4SGF7y6SR
NhmUpo/Rrva2AutDBMFljNxKfBB7EDtpTS2eEImp164q/xjMb16qCbXUBUhHCgTt65bdOvHUtabf
5ORtffnbdeYbaml+9VsFkfSE1sYz3lggOQO/PzXXNQtRLR71VKnEqbiw7hx5Hx/QVZBpimJFDIqp
ORK1XjSnxrIHhp9GIpp5pBFfLFUzYWIpPz8laajTQD3BT3AcpVtneAp34uFgct80YyWGGe6Se/vy
WalkKA8kYQho1weropqh/NDTnl88jvz2lIbBbXnvL+MxBHlIiP9Upb5emj4pLfPy9G/1Ac9lTrUW
TKNMRis+/Ceb3hH79n83qoQfeFQ0ugX59ORW2uOWrruqOVaJ9wmFRz68kJcLpsTiRIdJ7QWzG02c
bPRJTluqEgSQlRvDqC/e+kTj6NC2yf5HIyvjBQQHzfGzdOB6jcWZyfC6jjTlW90MsCukQCwps08c
9XmRCwL9AH8N1bIstYnjeooAsRVLh6gcFZm/WvVuOSE0SLWHWSZrOnpYkxk1/y5wpziIhEDmFL8D
yuTlRcnrfFGD2SXdbivxQLR1a5iw/VmnSZSSfqiyU+GzSGxgaVeMCljwn6cb0S2chvKvg/qtnPCk
AtnU0mUYZrQw5P+jQnx4TtXrdCCmtDfhsD9qor2ismoFtxNvtbPvyxEwbLI1uLTvIXZC3rDYO4Gk
DhUeCIKgVujI3w/MM+KCL52Ybl09uFr4SebWu6vx4ldzxJisP/J1pwN3V7vVOFpAX1Yse8wMw46v
8kXfvEyibWBs195d/NCTAvI7zDu845tHFc7ssqir8c6cs3LaGYqgBDAfFTppDcFGrqPpUksAzFkk
dEDegYTCjh5332Li3eP1Xp68o93EhlrknAg7EQC6/O1da0S4aJhwdybe+NZPKsT7+9+Efo6w1DQC
zxus/b1Ir5dFjJxFFPEJNBzUYaNhnVofNM+BNyTFN13EDBS2LhB465kRleAoyRocNg5mN0kT2Z+A
pjNMb45luRTIBAP9ZYomJWYAzkot6mamSl1w8Ip2dlCfXAYiPRYFJXkq0uz+TUIBAk9IJuPpqoRf
+aIDYOlT/eKkDyvLBOo5WBz7k1PMSmySSM7iZJ21dA6q1ApJ0b5kf9dmkZfOLa+1F/nR3tiGjSdR
g05i0BYt6UhjqnlhZn0Ze+adsRcY0jm7Hu9Dp9oBCZk9kls1ScGnS71rnL24Ca10SuSLzw9yzjVS
/8RKj+CQE76kT+PXeytgC8v4hQ5+79WCaPkau5EMdvGj/4cPZR7AoNuXwClapfZ0dSRUVYZV5Uyx
IW9xC1gjRirTtp7uNhzlHBs1LV4g6Q+a7RtdpNzGjxp0r45YQHydpnQh2kbM3JANHtfi7rOB58E5
j/yaBYo/OsqxvilZ8sqf3eb3b1h3jUYWzvG95PD8u1RlaaraNZJHq+tMNmuGt+1S8+7z5f5FFiD7
vrPQO513b4fGvjY5cAIUHpR27nOH7cuIGqK748SFUt1XSoM4wU4B8E3CdQ0cyrJn4gGxlXhDItyS
d9z2R9vMDRpUQExMc6siImV5KZMHThEYe/7xcbcIjroCImZWQ0llIYjUGWsiG9mBU1YHclTdWCnc
0J2x1fs2doTjlB9lvnKO97Cn1xB71otMZwdplipwjURxIdHH90e7goDIqkFBhkE6L2MBfTpZvRhX
Wdln2SgPkNMgdt5Y0MjMglJiNoLQ7HEiU4Z6S4dhS4keLS/d2oGH04yvAxfm0XXqyp+V0WOLnfDt
6OoAr2aJvrjYlLmce7gsAAQhroK2smgMd41PmY2RSPhk3oIyWcC+gomsCwEjPoalaekIxQuFrK7O
kek1V1a2abeBLrhFuUQkQFgTTOYYRrbBEl7LidBC7x99kudZylnA21gPAEngtxNxrchzEGXgXpGh
TiH5x1jbbiTeVyJnJgtV2VglfZ0ThNjfCnWEFKjOP250upHWFfwUNy+r7OsJExe13BYnAvhQyxNz
vHUoNvWLCDYQEl4X0CmpNZPY4l3P8l6aiBlXLayiDTokjdP2Uu/FZAdgMFI2SzAyTgS0sSpC49u2
lBGXGtnMl9o1RWcXdim57YopqWyK7erWBXCgFujQ8OnRYjoTh3AJg8OW6O5A/66NyRz40TtmvciV
r+5sbOYbqKo8SPefn5QvwHrSD37NRTbgQpLwu37jB56ZnAt4SdbN1YyhdGXMgZjDmcrsc1jAXibQ
novLJb2e1DQpWDTFo8Lia1IrRQpnrVM9GD0Mayxztd8BJtxt32saMMQwJM05Rfl322jJis6CgrDq
i/uznhronRdQ1tRt6E7J4LSJmLrMnDLETbwvVr6Udcax4ht0VeaxY2QTwA2JsIIwfSlEgpSJXhxD
zszU97FF6jlwIW864rXuZQI7UYG/74n9Czb0Nyno1LzFVCPsIEkevPaHIwCyvlBg9mZTeh/c+eVM
6wrmIHk0MaLh35RAmIkH+78EwVJXSHEnJRZuqMsSMjslg2o2QK6Kn7NODUQtsMFYJxhLbYrnvODz
NmVAluvJqPNJY8sAGQ4PaLmcUOmygaUU3i9SRSxtrwEZYurpedGHzkEIzejv6lj/zZNOHDHjzOjd
d46QkVQWaVW8wyAZhaGxKv8KWrPav3phYRP+66yO5bwCy9M3wqziMI7EXurtWggUNPCzM89/qe1h
gygFvkJEMzq5YtT6bryeAzyHyUqyyXCkU+QBhpX5lz19FLgjSdJMTnF2ysXJhSkC/xppNpKN1XOK
p0j7shjcOqwHFJmlCXSysK/sDl+AR+KEhku1l2Qe0aA9Dtk6OMHmWEQsKBCQU1bMDn5i7zujKY/9
aMTMs7aRFdvKmH967sx5gTOXhTWFYCZR32nZzO/RPBneXmejkzlCHd6PbrbplTpB4X+GKCV2+A2p
TuDHinBCT9zujljjJCwTq0CRkJ5T8cSesJC0zPawXr+22uRROJdD16fttIxkwjGbPWEYrn90zNcV
jS5NnAHINyiaKs/HbfPy9nI5gBvGcZ92IlltzO8knfGFsutws/sMhJE+6u2RoilX39PtiDC6l+ZC
JQN0GlHzcR446/ojw2664a3aN/PL8xcXrPwlLe9Qxxnwqr6e1+rATqaJSDov3YhnPwLdNoJZ5ftW
kfG7cLQpCNl0zgR5q2L7cm+Wtjw0wOPT9UbYaL0kl9MfiT9buLWHuQy5DienSGgc4+cajWEuKHwB
RlLBipgGlQsLOSMxRKyhUBzqru7A1ankqYhTYBZC9yXF9meplyzHRepWP7xpT1N9inaS0s07Qloo
+/7QgsBRYN5CLURYOoeX8vundypRAMC7SuIyNcZpoJq6pRFrdhjxAsjQHEfeqgANOp2rDNrB2dm9
Jkiu3X7EZzKUbOqQA7xE5I8mUgMjqocHq02pVC55XPqzrt7nbLASym+DDQPQcJTr1HPII9LPya+p
i0DWfwgOIcQkndwve1GRVPA60sCffHvM3TLj/qbyNlcEI/4b0EFrhtOWJbMZZoRi9e5LpRFwM2sx
6z5cZapsYc5olpL9d7xPEjcdF9rQabIwZwgkc+/iBINRi4V+OA4FGwllCQo/yIBkOcrX3PAd7+l8
D18CV+uuydNqp94+e84B9m+rMOQ2jzLpfdXoyppYlrLZIUVJQl0Ju+HfzGQu9yYEK7q9r52ZwPMA
FXph46RojoR0m8AHDZ0ZnTjLgATKxyVwd12RLWacRas07OCOYyhYTXj/XEeCrfCDggDVnP7G/zFu
huat071QDea6OTXqJqCcoslziuVS9joQC9fHTVyuQOikMfLZEyU4OeZTHwHVOyU7DCI0w55S2k54
i7b5PBd06kg9BXAkR6Xph8srBrmEZov7W/wMhlXWUAbkuYYmd6Q2qDe5XjdNHVbPWRcZ3vBuYxQ7
uOZFsy+KxjPSMr6SZq6UXHabJrLstxerJAHmQ/qzSPfa00HNnrkHIsaMEtsvvpQkRBKNEcrQBFNn
K0bUZY035Y25pQrJLcAdmQicqkvCH4CKBfy9Z8c55yxA47h55bxImfa2J2iK3BpVndK/vjj4qPdj
Nhu5SfXq2NU5lDI9/U7eMStwHnnCoK1LIdPbNCgl17rfw3S8MCbbL62HXZYTo7+6VrSvUJ6QXXnu
l8RrDdzjSn2PRjQiufEGTe0BmifgTW6dbeYymMV0JTqhUOA9KptqnvZfb82maA2H59rDBGeXijYZ
WZcaxJlH2L1D3kx4aQtWNvZPBmMmDcPu/uSazjQl3PbJGFrvsVE8OJbkxTNFcUv3druIyLx3JnRt
A86eezjSWaOFmipSa22xPiYJNcpofUaXBdZTHg5b9YZFHf1X4gHWHS/1gyptGA/JQIrD7ApoRY1J
A28ibm8xT4hfSTiK1baTz8MP7yfWnruUMkM43TlTrUDj3+EdBBALFxHZlW1hyMKC5QrjLFsUiA7m
XoVNJAM8VA0YvnhLCjuHI/9qEVZuFYiWlF3gUCw/fDLJSGTQpcCYD/ISSXJ8Czpf+Wi43kwNEecG
3usiaN5uRcOIPYNkMyYDPcnh24d+iFX5FSu+5XmWOIADgIzLrZCdP3H6ktG8IqXDMBsDxgiFtAHL
vDFPv/yrPeZQRN9hmNuLtYl9IbpmCG0MEzD3AkDuS/rNjH3lX2D2ShPr51CMiFyx1Dzwlelk+YUD
AKg9AQavC+fv1xicbuo4FRxHcpaj7KMuyYxWgJ18bRsjFIzUiXYFVZFO4swth9AmKAQzYSetnEwh
Bb+imYUHzuUuDqH4GX5KrzSrOiF54pV5BrNaj2jcgE+90Fboqv9eebcBGSd4UZtJt+fkPw4bI8q4
2BcJzN7BWd+D+9m2ttDVISwn/2wBPMl/NT1kcjwBcg2azRHaLDmoFHmsbmeUs1z+t/74jRKDQ/eM
kTkGgNJxmnnqBYqZ8924v+1DRhgwZjY7GDk2M5bpQGtBmZ8mQ4cnBG46/UZAfkT3CyHI0DPdTxR0
lNgiWhanL8w63GW75HFe8CaWLh6kzxL+EpG+Np2Dm+gee7hJcodmeeGc2c9L5V0Sr2eioZetoTpq
95S2tus8rKkCdGyZWz6Rjwmrm8qVlAmilQ9MSTDWhWyAHTp2ElNqWML52Wuf+BI5ztH7UZEvIKk0
2JYvYH/9/8bWFdy9LASOeEsNV9UW+XSn9DQz6aEH5MbNpMzpTd1h08EBF1mi2qL0OOSP7+5uikNH
wQ3JLydmjOZ8zyP4Qu1kYyXRvBqh2BiBrJaMUXIG+9fGmEfbCaV8DLtS+44KvABCVYLk/SEXrBgi
EXq7XWDWEYnirzz2JYuEaarpPVrKdGy8Zl6OV+3VVBLj4WhbcnkN+FtqdXtTbdb/9+VS0bwUE5Wj
x10dRCaGzsnPx3Pvg1NY3gQAVp/TbeIK/L7nYT8+/m775oVWaGcPVzp3Vr6HTrej7ujTTuul2SsT
CFcFIRyRhdv/eP4QoY+mY07oS+DOQ7/y43ZWRpq59qDUe8CB7B+ts0BSU2qS8DX7ALTWPpYTY7QH
dSSP++5Czvj2fP9xSBMrBLa/6FbP15LxIbcpmEmKsS8zKvJTkUYuE+c1tbpNUPo50Nz3EiJWpb5e
7iqNh2tUVJPIHUf5Um4/0yRY/eUCzd3ZZoQeXj2tPHtLVs0AIvjikeA5bcijpc6wouXUXNVOyF1e
u0t2UKiI5UgEHPrRj6C93o9osozCN3fCmhkLIf44nhexWpDMzu7CefG/aG+1u7GGW+U/iiCnwYPG
LQq9z71goeTycJff3sywTZuTmC+0UCxhejYay0u+wC4uVmryOk838PgE1KsegyIUfIo0w/W/rSP4
6ICsvSMXSRVU3As0QRwDj/ZDtIeyCNAz5li8scT/91Ux1/3beRN0KqZlVx6Ah6790EfAA/lpyF5S
GcY7JAgEjL5VPsnP3DPNSaCJqnDQqRWoRWSrOvjVfccYbIYwZldlEi7CBwniFOfH4zkLhAt1v6La
a+DX4IODSWbjP+yvaX4JoqmCpvqM5rOFc75Q88q+S4/NsBxNiD0N2shsEppaoWh9eZs5cIYXzonx
aUow1eCoyZtArmDFtWWCqbYT9idET4rtBMlRnPmMyxwy5TfB1nvYc2k4yqGY4W13BYVQAeWI6UJ5
TK9rZLWujuGRWTfSsRrgIyRqmbIMXi3tSM6XLyp8iGmA+16vkCzJEja2pnuvWG4yW4QIRke3Xgo0
aXD/VJiZkIbIN0CPQr2y+0yrI8KywozQ2b/1dCmQGfRcyJNVav9dUi3ngjXEmhEvrOmSKXXTrQxL
T6QYwKb+zJfldg64rCi7eAl5GUdViVrlTg4X0zHliRCWToNd0uAdgLNzhvX1wtgXaZkw6fc388n+
JD+8hN97dOTNBmzdhS0juBf0UXe3xpBFUnC54YJhZN6pAS0Pid007C6Y/izDakur2B7/39YCgj7r
SsV8Sb/igUgOQtwxWKySrQ0usdfo08y17DbAEthpJMKms76K5o/q/FrlWPJ0t7Ayi3BBkp1W3Hz7
b7lGWIpi3t/6D/SUMNHXQ2EHKWQmEGXKbUCcQd0gco4esUNSUz+fXGgrYIHF5p2O8lM//RZS83LN
7c2e5sIxS4xdSj28bqmtnPizy0PobCRBnBfVFmqW1JVvPqJ8J2371+nIPjOKeE0lVjr+1yDn8p4f
z6RnLsAXD+AauorymCJs8L5iJ0h3DF2UqK/btXB/iypLG9rK7uPvHi0uW+pkm/PSwyE2rpfDkTXd
0wn/KlIfZ9kxNcs3d6QEnPRN728EozgKmgKGwurQZ4vfIISLL648SlqELEi8Ou8KwEPqxSMnfzo9
IswqiG2NCEwRbsJL8CR10ihi2dykCx2CnG8VeLVMdQSNphV2heZmpzI8G1UJDfaefJ0YilXLvpaY
hk+GUqgp1to61BT/JURFYIPecCstXdPs4CtWryy0Tm+l2X9SdH365F7EaiyLN5aTDGExg4NnbbXP
whI33qQGfwnEteAo/ybFWeGKDJCnh8Xk8Lm9jtfoYGISxMvDSEWjUqH3RmVySTuIW/iBEKJAHmMq
evHjI0ZJJgyeuluGFQbnJUm3C1w4jTHz3ZvOYxAdgXzXOzJk/cIJce+r2L9rRmgFQy/S7AtmCVLj
FEjaSLu6cSvMpg9nFift8sO4aGQWLQbxgvaB8dpILJzkLQNdHHfqQF9GE4M3aPWPIgAiWrb2Z1Rq
OzgLnEmsvwHkUbi3Se1OjQL5jHvU8C7z0HbaMA/irWg428ytrlZWhoBqnAKkagApqn7r7U3PEmgB
DIct2DxJtCi8pxScRJMZtFMPvEyBixsnH2Klst/4OE2IpHjnfEwmUXk9VAoYB/mxC3bcr074/oKL
LVpiCPE53t7jGfNy1NROiQnucsHRDxNUOyhRY70JaPT7ABjNKxQkavWnae22afj2OY9yQ40ZjzRX
XQvKAlOTvPvlZ0QrTNYcY2PuvV8abb0bMMZVZuQwBzReAc+sayEjAJGDJLgMJ0TLoO0s2JoLpECz
k0iSQ0NY2QsizRubJOEDHgaLPwKKnLp/FnNkcrQ6E3fgaCtClGtv19JoCcxEdUJFt9LGZ7e0mO3W
0kPf/Q+gHO0W7j5P5+WYPHM4aDtaGxbBAchb+l7qmf9dJEkMXJMGHO9/adDT4a56Ccb5W+h2yQl3
9XehZcNXlGYXkmArLShlWpbYhoIW2EmpaKc+YizJY86LG1kQATqdfg2CV3mDSPvA1c9CVZqTJp3O
ZacIt5eTrNrcB5QbHXRmPkSxy8KbNprwLeUs7LrH/4JEosFABxZls13EJl0YotrF2cEC5AxfEkVf
jgfjOiAUhpVSXt1CzGOcQkSIkIa8hbEA9NC61e0fTtsT8DImPlQz4Y9hceSI3GdmD/F/a7MeCUjl
1Oomf3hyZorKR6oCanykQdhGzlXAGb55s18BDVRDlKWgEv4njE1uhS2WGVoKJF4YCOCRh3fPqbyA
NaF4UBqyLoNZkIGN9NSj178I6G5zETaYjlEswS1QilFd2ua7MiQhd8xr+CaZTrjG7OgrJtbksvg4
1HExUWW4WBKarxWltnPiCT8SW/XTAJV8CmTrPdQ8llmsV8FSPOPSWC4mWX6kQoe/z3HllGhFBxwF
KUfOxPFGlzDSjYJkQ+CKE/mgsIo76GRdKLKoJ4HDVewmOB3qDiUT4CeHsh23LElnuTg9MojmNRVK
v0rKzqrvBtjgQvGnYgmj1WAVJ8yXAGBl7EZp4gl4ikS9tNAuPOwr+MBRanhqMWRMP5NjOfKsJtD/
KwcDijq44MJUmqJpE18ErlQepfEr8ekX1KDQH0cwyeiwTsofXo4wL+BBrxlnpwTuJLksKgsTSNZF
rqWsIJTnbvVXEpX5dWHV8fIKTUmEilAiOENt9XdKbPzCxIZ/yQ+bK2kVfObW49v4ot0q0xLusEMc
YmjY8LZnoLP5p6pE8MEEZKkl4726QOgmOLMvLJd+Xx201pNOn+ilkkYplvXv7JOlUIfD5O2PAqc9
0LleCpkk423bkBA1u3VMlpypEQMTaDw0g9uSK//2miq25wgniaHCmgilqvUjuvYoYtTXV/x+Ua9F
YkWwcWSRnFBcS2q05zmqqtEi+KomdjcoHtjUiorU8WXboN85so3A4TwEyvdQlmQzi3GyRy7sv5hK
CD/CvRgxsoJ/KVuPDoB1JYwNcwGBogId2OxNj7TDqbcsS5sjnH8T5Hi2nZlL9Tur/tJ9n/CIa7/r
r6VsPoaAYA8xczBUReqBm7HarDsAnf7gBqSa040bi6ZFCFT0495SPXId2ttw4LBL/aybTKhFBQnE
NQsxG/uxJDNrTCHrOC+ixAzDouSXOpIUJT9Ahhma6N/x02ct546fZeDTU86qB651/9MJrw1+/uL9
L5Lt5O0+lKMHvSOMsM3sd+3CkRBmAI0VPt1KO3M8LijBD5e+hp/QpGbCcHwDEWbIo+0UC1P3WHSV
Z3Fr4CNtJGniWFatQ7qX8vy3lQQoURKPd+RF5G075CWfcvfKcfIdddUJZ94DD0EL5b09GihsOYwE
V6GoSneubfgnotbn+nGTNth6tJXqe8BE+w4ccUpRdQFbQpTyxOmKIcGJndKiYepTKIztiWFD1nWT
B57amYWPMPq+kEG7+j6ji7KiQ+YGaiyixWfGje4EWi9MJzktOQYDRfqHkGhPwuVtclZt2doRnmHg
0FQ4DBbfEW0kvpKC1BdUvGV5kj2EEBeqrZRlz1mW5tcFwY6zgw5hbh8oPg/U2hbsYVHYX4d+aKGM
yujbjESsYUo+v0BqujA3pQyDCDVdP9CY0UrhPmtnYIjQNitPBz2Y43jxrF+hSVn0CPL9SxTejk67
ICpqU5HGvWpccYPt2Y6pxNIAZIOLfsz8gPybACr4eEI1PytZIcVPfCr9vTTtUDPmSDNsKiTnLS9N
aIpK7hHo4n8MR4++G3aAz4wFTDKZHtm6mz/2LKjBNefP4gOcWXjTxqK9hns47aFg0LespwEmYWnD
GtHa+KJ7OmPyJvfcMBbGGNr/nvhwH/TX+qsmzIwbQHAj/E4fxK967FrMoQrU0IiOnP+McWEIaYCz
2e9hdhbHT3jHkN7+5eBRpaRaoLgD0zsxW9r44c92OYQWEsLTfOHxUIvvxcwvlrWA25nPaNgEIkB1
16H6IagWNC50DuUijbyrtskF+2kAhVGHGBYes6sbYx2neenO6kvlBZeCfvnGHs/m1PjS4THl8OqG
yK/LIJ+KZJ578IFOq+kPPWR65jILoZL20zYXg4PKbxjcJ89cOw4iXa7ip3YTcz0T5K+CBds+SZsD
kXnZeq315zPoVcUfqVjck+8pYE7AJGMt+PyYs33O4GaUHkprvAVAOWenbeoQInUXpcTJCqLHpu4+
dAlrpbbSdmYoycEH8m65h9RR/K68h2kqldTSDfFmEewrrPW+Ft2zP7jVYe0a3cJCCpqN8Harsnxa
dXG6grxtg58EdUmRIdqGaDb9QpLRMKu3qhAdQROvbMdyDB9fdt/KxHRhqeK0SzyczD9CdJ2oGeLW
4UMrdisxIXr0NKJY/MFsPQYrN3hr+L55Ioh1VK/DqouIr4rDcwOzGI2CBETRiw78mtZTgHI58FOR
rnc6XcL7BZvEnh1KEwMGqTjd8HAlWZG6aMLNEDibNdJNurd3ISX6iEYenwdZZojIvVyP3+Upjvx9
LnhzKdwwlCRp1tQLIlCluYWH5UhkY/STVY4oNZXqsZ0nIALeH7rLsuWF0mJMkJyCMe0E0/KuIBM/
akckmhwujrQVV7yy1qUD8FFrt1TybbF2M68K+x/Z1WBEy5jeUHZ5OLDVt5fJha+2uLUuKXKXbAUl
4ohjj3UTta5UAAZzIWJp3VMu3aBRa9saDJlmwXRfTdrn8ecFr0W5v/j4FisezjLuALlVaHbm+k58
Ef59Wx6cR/cyHdi9+8/ejKq89Vqlm1VKdh/Xwxp6k9EGBDssDa3WIQDxDKtHVzXoajUB6Vz+sU3D
1or6QRjKcXB6BKjJ4ZEFyS3MX7fmSv28raC11L0FaGpy4gasbY376FyYf+l10GOqMoIKnzG5CoZG
kDChIYr4lDZZberj4HcSfRTP5nAnLMG+fguTrwzZA1nLWy/4RgTxCzK+YKufsCmAyYyTvWKVvuun
HhRNrg9ADqNjSj1sr7eDGm/VmCC338vICcxi5AcortZi4xzkWLfP8D2Qy3oO//AYwfqeuWLhBdwD
uP+lX8wN2vA1Lhm1nt27l0f7jav+LgpC9rT2wNwaULsiz+esNkrsk7TA0zgPLyDONIdtoeoh/adC
7JazUA99QEMYLmXCjziEWfiXJiA9uSPtTcZkVJrmh3VUN8Fvcpy98DpYF3LJE8WAQcVCK9PXBOFx
NXhd8b8bQb9ksbs/lWMYtsB9SlFlWQO6BWF6bmnA+AmAIq/3GaoOpfRKJNc68AW2WaN0IZPjjHi/
NjOjD8jj2b8p2oBWsc/unruO27bPS4tuwePzS2CRUMCrTxfKPLZUIP7iqBiaQ5nYSQdR0EOsz9H2
EfKX790/tFKKRNRJKGExgnaEF6UNToAgAO2SO/IiUkNJYi8YocEIpcokP0U+LUlFftQeFSCaiGvj
MToog6AbbulWeReScrCz0Y6gtSKU8W/bmmeypMp16WfQBxShqzbquaaXkSZ7JRiUufMX9xQR7v64
CS+0ivQoyzw+RaGULFKk/T/SycrfAaS6vRInEn05RKj0JkuXfrn+uL+PpfSyvt8JwiDqSmHFleDg
dyF4gecLWn1SllgjEU3jhnd/tbJodzGu21X9hwd/q+tNMmsm1gx+rnGXUH6HvD+lGGsQrvTjLtsU
3iA25mND/ipxramGlpFUMEap8VHqmVVDHZFY+KRdcjI/qGnS4mwgToAPTMT0TYI6OPlRYp0YpIwj
KkBGUGOI1tH565/jFDiumkr6G2PN5OvPKarc1aUY5jJE6TBXToAbD2cNLVq3m3FuqRvLa8jOhi9a
sHKW8i3f3Cv4f2+bSFvgDyc9y3jEaPbei3/mtHl3mO/KVTW1u0WWWCIGSBQm046qY1ZtOSk38TkU
bWDjYzspIAh0WK/y2uO2c2Ok39Q1JCWQdKqTrwKkJTDkqHzkwv9g+08we5DqAnn3GNq7ATpdGDiq
hgxLY8M8d1VQ/EcP5cJjpS2OxoQOgQX4TwxkSPHpFS4owX/EOOOQLQTda/wSdtgWpZN5XVh9+THn
smWShzGUyfGi4fzlTrAvIFsGmj5VX6dfgQfouMX3FyO3pgyKV6w/AiC7OhugpyORHPaWUFA85QJb
At+tHyMxi+4BdSCB8k/Zqa2ANoygDj86fDnxmL6KsUbRPiUaMKcu9lMpGDz1PBm/3Mbv5Gch2A10
Zhf4uwjaKNDfrB/Ntzvwn7/sI+Ys8plo2ygG2FBjS2ywF/OZPfW8Dg7aKGh/76w5fE97L0odNjzo
ebr3bnGW7kqDzG8L82xgS0WWHi+5QAkCPHUsIRNncd4EdpIdxScVXV+v1UwXeik9v+QncuytR9FO
GVhChRDQxDDI+8pQJSMen2ruKwf1eHckgK7q9EukaVTlJe+s+SwoozG49R1axInWs2jeOAgZ8a3u
mz8LSLf7qVoVnrcc96fenHOCgMgrglJv6I9kUaU0LV829VOZA0/5zeRYW6febLYMkX0rgFBijNAS
P3mqNYevdQBscyFattI+h+Jz9xx55rg5NYnydN3+P7rsDHVSuuYwmAdBAID7iqIhA7VYnNROFziF
lWu2SbkEfTcPP5FuN7xei9RctnsrjWNJ62Vj2yopgWo69GYxjkmoFN2iSBCjEpH3AqNKTYf+S14I
WzeQKZS8ZgSa0tpH9eRPhMUom4USPqWQpW61oKXphc8BlWrA/MknIi1b3CTacNc5U3Q0voAV7JOM
w05g+oykRgN/6/DjDzJqY4ZUMrelrFqW77Ge7oLqHtZC28f+TbHvLEvxrHWtX708X/aunScFggUm
Q/dREStGeeLKlOmVZRX63K0AtcbMI6qm5nUlAFcgHMXLfFIprwCRC7ia33/oNiTPHycelBWgwQGi
FDcLRkuElgK9GCr2lse/TK2+Ng4UeD3DhIX7iPuDFXVn+OO1M0VVjby3TKqKFqnD0exHc/W+a7Fq
lTnqjn9o3Bq6d4VdnHVNllbbVlxTw/wZCjtn59nxQTVFCzzXPyF67r5KxA4Mk2EMm+cZJ+7zJ9jR
dE5rKmMMM9eu45Lr1E7Q4XPrmsCVon2FJ1tV3sGiW4KP+fXLZaR/+CwC66bTten3bkCLpfkFwJ3q
SNng3JQwVcX3ZHxAF2gnjCRJ4mWWcaTVyaC4c17r67HYjViu026wKw3k7fQIKAhfLmrZ3V/ZnB67
ru9sZ5aZBknJIeXAwLm6Y8+yW3ptN3wcHhvyu78DDoKCzFhevDY5QngKttZplotzO8eIyfzwIaoL
L+YTnXOeWJ4TMoZaBiQf+SjmixG1u4wuA3G+zS4ELNn1FDf3TF5lAOPaeGiLXo/zFPMZzwbsPXqG
HZbqJp42OgF/wQMCGbSdp1Ddb+aWmLBy76z5C+4ZIFu3PvooZmTp0MLlKMEVjgpXhpXMg/hBuKdw
s5qmTCvZSX6FXD5hmU4yo4QzPimBKFFTZJqu9FXHoityeZyBS7plAekOv3ML/emoSNmYjag1qmCH
oyhXWpspSJWCHoSmFcK5GU6keikSQve1CxZeiEL2xcq/VB4I4+vc10fXdwYIcefw01YHLMTa6Uiv
BtsxbAWYHUXEEFBcBloQFH6S+0fG+UZGpvF9CQIOz7k6uSWaG6Yo+1PlW8c/+2FxVHJxxcTQmFup
qgkA8B7RZpeW3F9uqB/jAcG0CyPdJb3YXe4Psr4wal9vsOE7xn1YYGLtZhkpUiKEiUQ5iJMjXPwJ
cjsxLd7aWIhG2O/F2ujScLbg3U8gcyf3Z8Y3s4NaOy9tizArb1rB75fDICjj6xRb6kVAShgy0Tk0
VrXsruHg6q2vnvqEVpEzXg7AR5dtjigQ4k6IduQlEcTDP2E1L4oKCJ2veTj9pjnjFch9zfM/+uJA
gjP/yovY/L3eXKnGMUoLGQ62n0EWdnfQiVRduQex4SLIWlw2sBVxufUIph3ZkgaprAJZ4f9pXU4D
FAxKkfS1t1eSwshAAhZABMjjVzVdNdtfo5IZWUs0lo0rY0AcGia3QORKXMBL4eoADB1VAvsvbufQ
MVpb05UCaGskSEmKYMl8a16/+2HuXGjuBTf42vx0+2jrGWmkO7dG6u2vamz3IgZdcb0ZTECTthQ2
G10VVDHH3xgeyFdZP6nZFAEjdVQQ0ByLxXgn2sCZaFuGpYjINb0kxqpM6TtLqDWgRirpbWRzK25Y
d9MWQA0xW48UaUE+MzJkCB7xc61yOUm3kHBu9nuaArpr4OHDEKcTctTaPLIKtyA4mDZeRHukLmGC
jO2Golxtp7m1so0aDWvgI9MHcaLMJGS7ZkwqNeBfk0vXaWddNmZlrwTRJw6vhz8AxCuPFpRS/+c/
NWeHgkd/TCwqzFYMpxYcJETQ7AnirvIVEGx9kWUFFw2wBIRaPZ1tXICGS+HE7AjkePOzrKEB/isa
RVz26ugtROcQCiwIhuofIytH5cRl2/w67/WNDE+8hgPpazUfMb7x39Xi9o8ucKe3eHFVkwbIdzjA
/pAxEVWc04+XsvgHhA554zwbTSm4cw2xpnW4jmTw9R7rK97+tnokxQ3BQRg41lwvxPwmyEck47mE
Sm8n6slu7zKUaSVNUahmH9Dc+E9Q4NLjAYJouJyzS7mCtGQJh2ZiDzFrw9iTYhbRrx/I6ned+wDU
x8eTb9F70v0zxM2d05oK5CFnfY8/RfdRWr3Y2lWB+lyqvUudCwoO3raPwPbWL5rX44dOny9wKbbh
Ft9wbXovS3PMlpGJ4CvYf0jptDBgi/QQxgywuBI7fYNFo4UMygH6PXPuYYrLBJ3NGYusVkICvi3q
XynK3/zypUN4E5KrH4dOK60deQZGo+jx1S6VxIcZnS3ia52K6BC/rOfGu2AWOgrBfvzvfin77uI8
fAzuqkZW3sZVOhXPXnhq0GwuKMBhBPIDjTI5O8XMN63/1DBtJ5UXna6ACl29dKWL5lQObXRaii4+
Qi5G5Y2mXXqrZpwr/QlZ63wdPlW1nhJNDa8FSi2NuYtA4stSNREph+EsJ3aMsy/tfl38TmNE499k
rkYqOyzXjnb6pB19Je0ZZ2X9cl1A3VGPJkAoAvyk17wk9IvjdYpMm8afrBT58CqiqbVB5vqKVJLg
yGF4U90ZlOfEHwZ7IojDyBVCXp71YQAaBtjCabmF0zSptWSTm1maj8qasYTz4KiqaFNUVI+1RjTw
YxqOF/5SszTHNmZAg5WqfMxZ4v1kzurNTaD6b4ll9d/afqSRzgNW5nSSyErNZ3fP1hPMYuSgZext
cJyasFvWbxgdVKOHpGHfiB/udIJrAkFN1Tp+2bn5Hs/mQd29oeE4IECeehJFr5OsPHZszhB+N7K7
R50zdFfKwC96CYpI14M++u+/85Ik8BkUmcCEINNCAo+bOUHbg3T9Vy4DKpsBvvomDYlN3pbMAQV6
Cwt1zlUDhmigYpiv5opUHd3N/BRS05rsRlDSEBp0TzmX8Npv/UPSbQg6IQRW2q9xsAXQP6yYcYF9
8+jCZTPjPJOLdo+5RTPUE4i/hgCUsaZijthOzDdPiGPIHNnOUovUOXXlKum2/u6vSTwavhlnXhMJ
M9LJd1D+NSoxTzK5VuTkd9A4yUO3MtWZsE8/ehsmPzdFC7JQ1qQRvzqwYkn+QPVDbV1FjqdeigfU
6/WYkuZwKdxJfLq6I5Iy3DcevdaDs94HOGl+wljuWB6bReZnz14hDL6kHChHjdEgGnU12oFkmnZF
hcJb4skB24XsDxlfRgEFxDobme+kOfzFc0M3GZ/XKphSr3eE4eP7CeeEZWijo/aKKenIgDJNOmgT
VeYDkU/qHnTeY3aARsfsRN8M6FYS5XlQbyWCJFm2HXBYCD4HfxINcVGEPcM+MIEXGY67FV8tY10D
geZUxb3UMPCq9N3dfN7+3aBg1FiuMeUmcRRIAvf8BljrGkr3Kn9qfNQtJbydTlyW9nS74/5dSafi
y8PNwHtvrtAlOcwjnmHcU6LysF65YbOrekEOoxJOlryRVjD92tbz8t0RCzBS04qfMu4QzhZCJJH0
wSqFzyfkAGYsO9USew5oxdJIi5SjFNvawu7Rk3IX7y6jCC4vN4xvw44Sk9EoBamQ5jAgha2m+ntZ
/4ykZ+tctO6LPmcBaokCDSKB3zmwYhC5RWeHqQCmdUKKoxWPEC3SVAyV1a0EksFSrlSVWsuQJSQK
1M0GrjdiyUXbR7udP0Pu3eHQvkDmBfBBDHqWlkub/IxljxZyscrDaZGLyf//h+ZiOFKuIqMqSp+I
OCgYs3cLb7wnFW2mV1q++9r1xjyDELoG+VixN5urlkT65mie+Ef99CeWEMbRtd/OXfGhGGK0cQlI
2Lzr2gJ8olWFFS/15yMw8NCHbW/GDlG1pAZRU1V1p0+odzuM4k7+wedZEjhob8iBLkzAS5inaLqO
7oc3XO1cf+9ccI4oNYEKlCWbV15oygdvxw2OsBrIHM3U8ipBuMmL+Z2cwdgkrtAwk7vlAOJqJYkg
kIbYQ+v/jNSQxPDYNFzilo+zABFGAzBH5/vrPIhrKdQJTod8ndYxaQ48oE2AUdeEtcuf+uBF7Rsu
hQh1wP7GkhthKME9n/npi7hcOTftQYGqfFxiPvXDMp+xNshb/JjO2bxJrH9Fbqh8yh0NwPr9ZqnX
DfFzkT8CL9VfroddguMheQuMKra1VudWSVQ3CvRgWG6kMS4+D6et6Kg9+F0cJ7vzYp/WPFDOfA5M
4mBUU2VuhuP/QtUEv8FT4UB+G5gfyZEEc4ADJoS+1U31aND2/KQOu3wZ2CoCGwoFHmGkxrexY0rx
OizRqOLP9yKyp55akPIH1wL8yMk7h4pAnsJBGx/Vgg29LtApzW8jF2Sv8rXVFY4+AjAR0T2eawGr
kfquZqT/Dv6ZQV6OHGp4pUWVA0xWhG7pGW9o2BjXjcdIgHVSWRu1Q7hohf6jd7gY0xRg3VvqaUm8
2ttoNZ+rzTUFcYewtYaXp9BVquamcZdIW5hF+/M7YA/OI/Xmp7ZKVtE/jOZYadYfut9CUaf+DZr5
pelox0849NBkMN3u7Wp05763OQ5dTf90eDxmWOE3tjKgUnIMJt8zFKVbVI65HS/vEeFpNhdLoufz
Ttqt39YDozzadISHsrQkzrfYetHBevqDC84HIPJb5iuTEd6R4ipT9QJMdlWZ97Q45rI5xnt1cC/n
7baE/xxGkwaDkYzinDgbuDESsdUOH6dsX/SwAebRS2qp43kLIECRsSmLlHHYBJZ/GSva7psn4bhB
RQREJyCkxLhSCI02R7XPCzPi999TVQYpweZ6tCZzqr26GAWPg8zYLO7jF3+2s3JjdtxYlYz77GHg
2snIIVfsPxLB7ZVnpjOwf+O4DAO2980a+m2qSUriAPl3TBwJbs+fk82uZCNaytMG0WkZa1b3N+SC
pWPgM99MyaYmoGvd8n1xwJShWZCg2oeR1/iV0z6XW86QSFewep37580MOmM4gS4Qr6oOkrVgH9EC
0vIkGvTJW+jGkLmKHlVG15GqDexdML9OQcAtdWLB7PE8IInWTM9Dx2Zx4nlD+R45ctyb38v/uKTk
q6tXojLHX/W0+pQs0bgSCvoafXfddhW+HTKW7Rs1bgzC/fL9NziQ/Okp8UaKVWXG21BAmYbbDPRs
QWVBKRqtgEVs5yerxQEpUwq+/QUK3Xtc4ksoc5Dvf2DUOaAHp7uLb5rqJbPVdGRb0HinPa6CHJPD
o/WEM5F02+g7fxWEfI4KsUGLwkRVc8s/xGyjfVYeLnm02b+wHFAwax+VQhdyO2tTfxnpJQlXy2np
j+qfxjRSIg0k1VAVOdynSiz5PdSSztW5JSnFeRDdnHrNKldGdojZQ5Bueo4G7zH5n/YOKpdZDcBY
iaoIZ9fVWAu7mDbeSAeIFOEVTSLREHcwUBhsg123rvbUrWP7vy555D3glKoRNg0taFbpGhbBW8Gf
adwCQLPHyB2/GiG+8nbPXD8VkGYOEDveN7GfrF+Q8hmzck47r7qCFk2Bf492cM/m2i4u2toWuVxk
CQody+QnQChMu6jMG6j5caYn/KllZ89asi4YJZn4Owy1eecGJesaFFBvrxIoDEFTNYJv7cGM+hlU
Ooi5dR07yECs85iBF3sf4mmz782jlUfTLmeZCW0rSR//AiZvdLpxZAbHoWzvJX3XAFyoQ6L6U/69
j4TPNMHgPiYielbjx0cWf74WKySm8M7H0G/Ygizyp6ORY3xiUUynchstb8Afp7e71HVVr+lgw6Yq
wXDos7uO8CyxVeL+V94lxcX9XVbcibWJMefqPsTVLSZaorvSnpCp23ajEfuoUfQTp/MARFvEtQw5
Y7v0RnwApLRZvf4OYpahfxeD+YLJfGghdc84DMt3C618HRM0PJOtihXt8QBOwgk9JnRJYGR4tNwz
xsgSN7ui+X/F1MoJ78PophAx3uTyVIdOSIqBSsMnwkR3MQhksibpsBIyhi0Wq4TJina8/1dyFiE9
Rdi95oCOY8kvX+9X3Bb3QLOyR7YY/SJDhf8sTeDaCZWfwEiO/EFb7be9YjEU+c2Yj52cJ45bE3CW
CR33eW7AYQpRoujZHSLvw3uEmSVFryn1AZp2iRXFwBfPPuAaxvY9K/aRw9kpFvPOEHo3kXmIo0mR
XrTcEtl0emyp/fmnPUvFjLe8mVGYjt3nNT/X/sdDUOynQff8BptjOHvi6KNwI+e4BHDVmiio8Ezc
fyJ1dK46xLQxMVkXGWgM+y4QXJ1OV3C2HtHuehntHE12kd1w1tAZU+XfHj3j3yDHuJrp83edvodq
d2uk+8YT6NkerArEW03D13BBIi8ST49c8CWS0Myga7Et0sU1m5KQHGhtWTgiLlwe8amIVIBHd1E2
tC4hwr9QsKJ9tKJ/y+DzYj4J0ck01sA0s79M5tNQaAhHQVhCyryo0MWsE63wAv26XWJrtSY9DOnd
eDHURA9lRhwu/DfjEy5USYm/juY9wEACfZa9s2u96OBHtENCeO5IRbMCap41Xkf5mONZkJFXKSo2
xLqJxi8XPrdVnbtkJzYVeLHrrNtzrWM6luG5N+gKCiuVcPMSfVMMf0UUaxjD0Eoxz12co84ao6bm
pA+CYgdoBqBGPReBGPea6u6DudbtzB64JZjyXeoFTRoTAOvN6PJS/3RID7919AGzuuZQkprvt6Vt
pqYtl6r/YBYMaBAtFT48iefTCbtpGxIunMDGW6OZX4OFEwt2qWe/QKIKihlOHCO5LfA2rLrGl45n
nxE+yNqiMwpPbiXDD0nhffpkHcljPRCgwb7052kzNidRbSpmpVsrRfcVYWDC3D8EmTRVDBy+3k/z
rWkLRjC6XUNyLTrRdJMkAmps5qoET7wV5GQMzofp99yrWOo+WPEimAmxhb8hO4bvkH6CKZLQUSuL
vYlmvDAkYCJ1JoT0kt4q4c7ceh09ALufAKx6yspHB9kguLsPB6UaWmrHKIGOjXgv9QrITzAWE6e/
qg1pE100jQqhKU1V3j00bm+yFTkh+397mc7U5lUKBqpFiMm3yVdHJa+n8awTS/iUHnVCvK9Dovvo
swsejteyW5Q3Zv2sCtbFNfuM9EsDDkXsj2DqJFeW6n5zGPkQTSGYrvooWWy54sxqFxyU/NOkX5hJ
7cL/xMm8NpXTVMFbwr55co2YWUQHCzK9wOEaG7ZyXlp6UfALOqBdu65VwsPkvGxisieBb/qCS0nn
xubHD92nfQt77DQLi1rm5yNcSsz5+tgcxnCrUqXcMwPiKD3HpaTss7qLaxNrzHnmzSamfoQZGPIm
I+KbpdUcVXQumwOOZyGPKcfrCki0AF+4pkO4HZ0wRsyNn0aGMkYhfTYHuZLcw+Vz751pn6twIDIL
Tj3n9so3G+cXc20krv1M5oWbSWynzDlDvrF/kn1Jo0zjBv/CixenPvOTLYpgV8V8eXL2BdV7F44z
VnVI3CdiUAPg+ffh/IVR0Vr97pwxf/45gABUKuJlJEZhvqr8SzQWS3SuURGndlTIufBKb/nioyJ5
oZXhZIdXFGTxW1s5Z8kVzdDRMaqcngasKVtPGVJRJ2QLLa20KaiApya73gqa/afJBPNLwoIW8ynf
tFiFhjN0/T8qTH5YLI2vGfanvk9COLbvngpfUNTewithb1MRrNv/Zk08DmjQd73YfIaPb4cI3hfS
hHusf+kNjsrIOb+PFNaI03TdQ9y7/oV10OvNA0EOkYtJyVF+oC7HoCcoMLhcsmk0kZquA+F2ASCJ
7IdPhtEtIaiAPZeUcpyR5uSSBSg+SHU4WSbtPzbyGVusHLRvTc11QQ71G0wrxFnkbBrnV2lxZLqJ
k3RJkNk1Hvhlxiodv9McCBm5OxYIF9flC1k0cLSU4ncftKnwN3fUaLsphkMRBCFAZo9ApB832erW
2RJ8BuDdgE+otzUheewKJTieK0LupKte2QeUagTbFlkexIswINU0JI6TSjbeN0v7m8ZOs6j9iXHL
rFgCcwcgWGIIdr5OuyjLGXmIshgZyBcuyE5H2NG7OS32KpqmpB+MwNtUABzBxFvWsEu3iAGPV79i
oYIOt/vyT0knrctXine1dp9mgrwH+Tw0c0hEP4YQJhJlql45UpB2Taz+cEFcez7FAprhtfWzYimI
omvFzWahiQb17/WyFByXgT3ejxW3CjAxLnY05RoTbdTLKsUx/et1hvkLny1JvE8rKcpzKqd90Jl8
7kFSUQIqvSQMyrCVUEfzePmnZBeA5aHJOn6AF4R8o70Y15kId8oUJLTceCCID6j6h8cSroZAGFdE
LB+C/yWkX9VCzrmjoSjBW7LUwad39a1j3ukp0Wd4N0zK8+6QXDQ7xJ4q02H1VImXWEIBCBikx2pa
PnrI6zcbQnE6ip9zt1eYrB2f6qADe9NqZe2/U+wXRx2tHb9SbCmpuYeRYNu4hr0i8rrySBi4Drtb
jwc0bczEMwFsz/K7ySLf35B5XoEcgcfAIaztf0f8j3Cz8FbqK+Y+sB/82+xKSRK1yFIT8iZ1jmAl
mARHlQS8HnLfokcfphP0L8h1T0dvQ+0fN0CD8DiE8gyHwSMJB91YPfbkbvfqGKLdApeMV5aSxWM4
rbgcp8nH4Plu+et1YXCqtEB7DeYlz9IgADMadof5eTkqGTBRXfFujRo99MOkhT0Sd8GAmOZPE4rf
d8Dpw2nLhIlpJBFedf587XIWHzOpO9Xg5vnmbmsbyaVp5TbZtC2QmBgSBJPVXyYiQtL6dAewZ0p0
QzxTRmC2YfK1UT8yM0e6hXs8Pp6fWIaVhgC9xEKfj0cs6dCzK/Ns9xFCtS60MManhmpa4W/OkGq1
oFmQqS2PkaY+a+nTXNzzVIZf0t8KcmsHw5Up+GOM8lugRV7kz8wwDUD+jbNlR58WEWC+iDTv0NlD
WUeGJ88TmMp3vHAaxCVEFujv+b25NX4d3Ij7Z+xewaOCr2RtZi3A2WmeZPB46XZBWzcVuVptRAvX
2CUnYHVD0AugwoapG+mT8V3yKIGoBRhVEboM/lDvDqawGv0twttJ1OOt7hNQ/X8kj516QUKfmyVb
wI2K4Mk14KVqERBI2aFJEtuw+MSLUtlTq19N19kxhNAHPN0K+JSDxaCMXR06ROvzYaY71PddFhX3
/QePP6sVnwIwkxwSDNLuUug2Y/A5WTqUM0ahrnR2vnHpuyHaP9U8ys5HeMuP0x2jABycYaXdF/KE
iraFQLW85sCxSHPoMrFsYVaqyw2GvsG6enzUIAazVSMauFMtvkFUT1eI/cgDJJyb9uTtz6eO9yWG
C9cAWiAW4n0LM+EnGTzCBp84lSU3uSl8Ta9tGlsM7YiyrrDb6ck1sM/4YLU3BibgBNiGX+D+1fUT
dp5Iv8hf77Sn42gHXlVSpwJXVWsClS7DxUqHFn4QvcNv5emuXgjrytLoFxk/Am5anwNu6lvfc2o0
lzQFkVsjse00t6AKf7EP0zIuYc7ZZCSI0B8op/JcqlFjqGkLD37vLZP6FeAZKQ+yho6n/BYoGe7U
UsAUfhK35faQ1BWu3wRbGHwMUA1mfL2KCr97IgXu0vjr6wu4qHY4xVeDC3Mi7P9C86U4yU/cRFoP
D3O5jhPVG6L5Wnb/+yf6PWnRTZo73n9J7f38DVy0jPHdyhFs5ZXrpvdOfUKsGMkVi37gdSNWMOuk
06MCNeFjSmNDU3t9RTaVt0pmrv8GEz3nZZDFfs2hDyzDnNr5WcpnPvpAWoK0TTBIsYm/l5A/OElJ
g2eU3UcOAg4fa6gm2tRahUT2PTt3EL+vFlcO/32dX2BJSmhxOV73mcux9iYcfP5uRsbeGtVNsF/c
QVr+/RMivXJqmAhVmsCOnphKEb5MfARcJ4YQ3u0j7QL6sxwOqQ+c0c0cfXgLQwG2k1372M50VMc6
apLg4RwIi1NXkaruyGYPkgYnt2BqIqNFQUnlVftwimfzjapcEg3cPUr8DVXULE0uWAT7HT+JKFF3
cPHNrHhsgX5ojW2ZvuwL++sBnBapOoj0YL3302xDhKVYIczdYK4NONmzuFaUWXJOCVpVyFwVOktM
Pcdp1UkH1oixQjnujhzXzrPuL0axrz/dd8PFCfnzg8V8ppGTmqMtbxV66xlTDjqTcFRRNXy5m/gJ
bp5CzSqL5vKR1HcTd04voAqqoYTci4cS9tfNjR4xWI9GP2MUoBun5+R0oz5hbm+OS1C/qb3kTo/e
sUDiWtz+tw+i478Y55W0i5sTnWQTxvLms3XBPxCNJHKIMeeFuGBFfEI3fbYbzmeDrdGj3o4G/rbU
9HZeB0F42ASrH7YVOAOW+9GbtuwUevH/VDW0pXmM3DyY62dAsOeLgpkpMPliZ3ZTazgdB9Buy9Hk
MEpXn1YGI25trvabzJcfChUVHjmM3TVz0RG3PODGZzFRqh6JFKAZ/b7Oye+ePAxV7hy5XrcFea1e
xn8qL4Qye5fBTvBaz7h72KRBcdE6l01tTTs90EsgiKtc0f9iwd4ixNXLEMJGc1m7AnIPrjVZRJGi
EJPveN49Qso4qqR8CjzyM23VYvUSFu0rkems/wXi6VJ5KiseUUk6On7X5E768LP4fKFzjl8Sxht1
DI5tujiXet+QbruMvqwwc06Jz+EjyFoWBiE0GmVtmrX9OA3o2evymEXWIYN3K/LWxUzDWy3W0QUf
InNu7On8y1s/DxWOuBOEAhdkaE3bbFXdqlTuuXT/dIe+4a21odVzswGdAiEAi7WWVEWSimycyZZ8
t3gXtTZI7DWdpFFKvCn6SWBnZMFEuy1etekdsNEHrH4l7RzT0+ZkjMMM4f2wHS8x2LiMreXTAuZn
dDmo5SSf3NQwP/FjOwOlN3oekwoHt7YCtyX9NwW0Ec0t0n+A02wKTcFeQmoUloIia/O5H3k8r+im
+p/oRyIkPOLI2pMhI5f4RvlYjha18t5B72mM5iXbqCHX6No2sP/uk0Dupz9QsqaHBuhCvl+NVGcx
kLv3dlwZy6AsRVPNckPmPqNLFJIBHpT8fgS/pEuGs6j0WDFvEblxCzca2iUqEiTPVFfw0UvwzSey
ZsT2fp3pHnb+01TfYYXuDUUGqp+pT6gdRET7gnvCJ2l6BKA3kLL1cGG9dEWlVuJ9in6LynDn66Xi
VMMIx7lP3VKAHN8ikldnIfGhWkNu9w3PYcgRmRt8PlJdhzT73KDdszLoPx9+AaD8MXLT/JcNnf54
PUBu/NIQYCs0hjJ7MFg7407NNBlAq+7oCQBbIGnj/lqHL4neTSFHhiAymHAAjcoZp8lOqzU0kMV/
YyDoQrb4VzKCIhAQ+C13QiU1R7IDlFI5niPVlJ1TmXfk9VdhEzgg8YmglhOgKLO5xDfjfxVwfcJM
Hi39ChePfbfjq8Fi/HuHzqIvWYsYsKVzCmHlBOPCk1tCt+yGxLkYurUTuFuWMbpb8LnrkJvPxG1c
0eP0VLNL9oJEdvm7C4s3UNPM2PjLjXgEzj56HBcyqdCNkYbYt14SIPzQrmsOwVwCk6WSE7jg0zc/
lI8Vo6NYp+rMExUD6JKAIWFWdieS8Jb0yZ6anVa408jRxCWYAJBBfRPvw2QM7IUXxtcBgJgLw1Pg
Vn4kDpXfduqB1tz76NpyQeqBQkKczqbzpfJDnm51Tb7ttd9OrtHndnLioW6+9rP5KxvSVWkHsm/C
8ILnS2ElCqr9/KdPwesLOQqG42fytdfpGhP3ZOPKqUhUgw7o+f8eAzFyHI9i7argSRqZMbVMMN7I
RURKrmgcEsHXrwGnfe5qe/Es3XNIqtoVZePjRaLDvX2FPw+yKGXTkGQGQcqNMBV/qD+zjh+/REA8
+ChnRCL9QHqlwsgt1G+fKlTbYbkremU4ScWQgicmhOTlXreAPLC7RWhPjA2cer5Qq07Oo3rV1LGu
mZL/GftksA0oxEH3+2k6BHnZz4A6EfhrY1qLJx/2bAmLdH0fxKaaPkDmTH/yh/h9GfEaoTC0WPLk
gbnWpFzdO3U3YVdd7Di60Vt6TuQNFNI9EMGWp0/YJS8CT5FxlH2373GrydoyVSqJXaw2z6WKwHj/
/iOBWk0VML5ScNS9iziuVLjiOQslkFjFYHF8q/sGWy+pSOj6ejtNTeDJ0/O7UvtlsQGYHKIaAO+N
/7iqPq9t8U3jd5YluUME5nlwvhkB4rwYEg/C/yWQBlgEuGPMMB92dCGA3TWZ7JCpRcpnfq38cly4
GjkSJxcB66/2uZRPRtc9X30o6RItjphHRuSXmTYSucHeQraTREjO6JBuaZGJuefl5KSs4oriqKlp
O7E8ku032V70FaAVPlBVUxlb0Cg0meeqo3aL8zfVhDYUx+5ZozJ+uiSphl0RVfC0W+pwRUhOJxyj
21U+RwrqBlWT49JAWh5HxPsizpGFOla8OoE6nsDT1C3RxGF/KhyKjUphaivucwko6k+9/j8m1j7U
thYT3hh31LD5VenzhwiMwqSLk4gufXrkhieQRfbEVP3lJQDmfo5DGSY72ueGvgbCSQ02RxgYRwZU
E4elyzOHh5IkQrM+GRt+9g++UNQXaC+x6PR2gOuxRvGyzWVx/+dgSXop0pfkYpJMGHejeRYiXFcg
OhT6clyXWs/d3GY46Z1PZ7f3ZSgsiXuszgEYGX9wK7gRo5ZYG3qtTjVRw1zFu5YAuZL2ZhBSH0BI
NYIxadODsNy0c1IR4lVNXyFYxFgo6+vCJrZkQL50B00pj3ADN2o2iAk+syI506/ywvf2Cq4e57Y0
S9C4NHSeEbxpyQvh+dBzWE/qHUICiQYTHXrQevCm7cf2czLuMMFXQHBqeMcTb9/HatnzMwnfyKoF
K2djw6TZHedQnp7JJpBprNBJ/WI6d1DeWUVrrZiczPTHrf8B3BN6wEl+nBaTBQ4n+QA+7JtxiGF6
YIF7q1slTQV04jivgjaB3qjFPvMv0zYpdfrWiWnjwORExrcrCD/mYmmIfvVd84C+GyO2i1idBb82
GQ2BSy+zlGSLR3JXiadYCII86okHlg8F4qxrg3NC5PHGr2OL/pz/SwfR1gPT7aH8R+vRXKKvgYXH
zJySfnSi2h7uFAhOEbZwIltagSlLnkB9rCtKOnBsi+qZMCa4eQ9RBJJSSDOzOP6p1toYoyIDpdUk
ApfMPCQAOCb4iJz/EAcs4MrSOO9DTF3PtSIeBzF+DVkd14g7XmzyrG6a+cCMmq6sNZb63zaQKoHq
9oeTcDFrtTBN3OvdCD2RpCLqA+TeQ2Rv2/hOY9YCvnjCJqpWMWuDmfuxR/cnqlbQ/PbFMXYFD8r2
a+zRtv2ja7zoj7/ygR5dn9yrs2/6ol2e4KBwRxqlRLK/WircIQg9QbmGF8+b0QbpEbJV/jDicZ3N
JChUbMeJwItXGnYKU5ZfSlsfIAc0KYYJR1UjmHWK9LkyKEdZGfO+LumqeV/lm/LiL9NL6LxI7DOx
C8/UNmtrrM4bq1SjwIMPY+QcZ5gBuXt9R92W5DXo/hNFBPskAFytKWxs3ynUOCBkCwtpVQON7hjz
dhN5UPJuz5OhbcFH0JMpwsWIKZHlgMzjybTRm3gA9+EvVQttcUkIRlW5nXw9pIUzXeKEy77LVQD5
mc/X81zjrAtfRYUyXhlGWkyaw94fxMa5BxHsoUO+al+ZuOjIR2ohnlndscKiaUWjlAHQlT1QCyCI
o0dOVc9JzoRWyTB5K3wWL4btlU1IX+nVAmrXVMmylFIbUOzLOLLablzeJyP1VYyVLhfZ7z7qlI6m
MfSQR0Q+RdbRHHi74zu9DmnKGU4NZUxJsQs29XIMdOdY0Fs8Ut3dyuowgqA9LA+p79zpz4vMSW8E
apUVkfXQUi92TRqu3IAhaxQtJlLzoWMj9AdY2v8mzvkC2tTi8XEJrOQjF0zHFYPoYgw68gh+cquj
AXOFUSte8hepu+bca8Qp+Qh/U+br5x9NYfCibDNFdFwORsdsIhTy5xm1q5DHijKSmUZZpEJFzi9M
P4RS+TP45FmZC9ihJ6ZKzBgs6m3CgJJtXCVj6t4NLxy8C+AJJKzzgpsLf2tM7I9YTIrJhxL6UIc8
gKvR0Uju8RkaR5BF6DqCi45b/WbEdK3cv9lhEjo0MWcNz+xYzcoxUpnLjF2vcksOmoBReFHUYs3m
yh1u1xp7BzB9iVDBM2BPKficNKvaIU79PBKdSCnT5e+kCAukXtMOEeY1vrxxd+gHvigZyUhulkLO
eDTeZyPioGQf5Bifsxj0uBemYcCDoL9sWz2dUBEFaNxn3KwtmGGcmnWJz7uPX0eVcQ7Zg6D1zLBI
Hy9q4MnSCcBCxOwM8vj03qeaiDKvhxpapEkj8XryhO3IjphTC3jEkJOkDRQD8gYBERci+xdjh6TC
e4Uc/lKqZ3CD0AXVh/3T/87FzvT2eCeU3uUgvJIbLT9oS1tSnADHaw+IETsjhtQNL56igtnAsx7Y
R8uKubGwUPf0QL+Nf/EXPjzLSo96N6XBj5EZw8n6eA/sqcdotOtkUsIwYHCV89/gZKqHO9ktXXTh
SLOkY+R5PlLJsKXMAtUIApPMFyNdfcCrc4YDbf/5X2eTZUHCT4rN/K1/1U03+sXNTDe+35whmRWC
eSkTMtnP+P8jRfoYw+JFDcSbNf5Q3sICZtWPl9UPHHC22FyZZ7X/zrRAhPOc0eqDTnKJ3phTNQvq
+KOas8nEPOg7AJt+lZHyGGc+78vssbFuT/XpQT9uRWXl0AUf49te2lr3s8woDOixtI+SCF20uSZK
OINgD85wRiA+08wcpqivaGcnYmivHFJ1r5wfSHaFFNe2JlqMhYwyl22MEtgVY/wZEC1TG6put4QR
uPJl7EcQfgQ17NZb/BRU+gJ0990xFwCTIJf5RHQl7aBfbjsPG0ih5GrOwgeuJySMJRbqcpY4DiJl
Nr/Z5woP4fl7B4frsxesLrry+jRL98/qHTWv8Z6wt78XNmvVeg65d3I7PslXqUsdIIXdm4lvim0O
n1DhkX4tCIelYTd4GUIa42vwcFxv2FrF+tJdNEzJP9uqnsjTlY+7MuerkIhPmP/DiJY3Y1QEmzyt
kAnLr6zra9HpFx5mV9mw+X14O/EVLzb990vDIysPmozt9mLTDeQa4BnRMIG6KUy1/qmFjXfQFPn6
xN4UHkk783b3LosQJz4WA6Vk2j2DH5GWr4U6gLnOkw7xXh+is1ukBgU9i9iLVr0aFuGrBElETu8Q
D7BSRFMXngG/5UNnKH+39/qCkZNGIirKBZxROLrMuJ5YaO1NFDMkNco+K/SbMgVMpv971krxAcBi
XknRWNPlBTbAslHOLvRZMTlxzS9vSLMrALmyDmA7DFU6iEeTPvCsCQC/haqW0f6QCZfUvx3K4rQR
KIU9xqM5jr75aaYMbJfOZ7QrMZSuglH0tNIhpBj6U+BBXm4kt+fJLKHBLiYHcpLwdhshUYVJi8Ta
gbXDmFujWBwR0HtH8fXU8szLN2RfM2Va0RAp2X1eZ/BAXvVOxljRd9KAYzdgMi5uqe7iwVSuSyOm
4TVLgB+VhyoSqjCdznYqO3+FUPw6Lc7w42qrHe5jDP12q+PVM27K2y6WYcoQPFm7NTCTeNfu7D3X
f16F2ktcTHg8h9aLPYUyKV46o+GKR222GmDQDjCFv6lkQE62rKmUzWTmiP+lwaZyzAVwSPi8wP5v
fwdk3a5DJLJVhLLZph6qmQShg/Y1Zvq8HwcNvA4qQW6UE3DZXRXyGMeXNihM1NddylBd1jsVYneT
cEFLZL4W7WiUjeTL9J2wdk3akXINmT/3FT8DES7BVpkAdYnz8tSgbTB3oDejDKk+Ou6r34ILd8Bu
Utrw09kbFuDb7U9iS4dHoZ8Ru37bg4jv3fONZja1y0YVLVsGUKUAwFdWc1AOyX6Z51Ue8fYlLpSW
uQEA/R9oiK2lyEsUr8yjHVyZfNJR4ydeq26Yru66JAiFtLTN5yoIT+WHZ9omP7vF0nRZT2tYKIEQ
7w09UGE1CUGSZgMHeqSPiMoY7u2KXMnb3jkDbPBfWuBIh2iEBCgZRYz3Y8UToC9yjiJA7KK+E80o
1YXsbb6H2Cz81uSIzqq8/9jFCWLBqr/1d13u/w1+F0OHFb0rmCUV7Z1Q16KGgIgZ1QHY5yXlstg7
yejp1NJEnO2ZEKHTH//WEISxxwnlEvgLTVYeTFLe+YFdkl2w2fU5UeJLM+ZlKe+zkG/cdpM0xn7a
lxqK9t55J2cVaCi+re6n4dwhFviDpQI3dpR6UZeGmRxPwGwGrip3oc8ym60pvnFkaO3p67pyKneh
FtBL5vAUbesVRltzVtjl435dStOOVloYSaL8P4kA9BLTVsY2ea3CyxkpzsY3VQhQxxyxfTWyoCyn
SoFeOj00FXFG736e0YD7SR4jJPZmGfZ49cpWmhCcE1eEukJnmZcH+eVoSWx1I2G/iMO5wadA8jpG
OETPcVkqvqcOVh5Z199N2BJCoJTbg6Er6XADbFF9WZ6hMhZrvAEvn+2PLpc4pYZeoSqMir0K+goT
LshlZhhZIr4779sCpYAeW/1POtR4RP3aUz2YxSZP4D0q581oXw+p9uzly1FOu1mRNpM1vsTfI7+c
3tuw95Geyw09OTdBC7Ai7me9uswzsnqShF20hPiEHnEoohZT6awz1hDPAvLo1brr1fjmurmyr50m
UtdU3wzK2TAFZ449BQIhLaQSSckgo40Z+5dk4GosV1ARrhZIz4HRyPb4nyauJmwGxSpWP0XZwO/4
3TaXw9fZ7kBA9vYHANLjn6mhZBuQWGJdjBcAb1SAbfERxCIZ7qJwpwix0JU6I89xGPS0w2z7fN4Q
BI9ZNZ+Wfr92EYiOG/dOh94LX7u9616vb2lfA7bBNttQzb1AO/csNQyPQlIt/Xewo+ChF/dNOL6a
6yzlAH3uBDH028lhesHvidgs/h/H3nAEcHmKapVGhwIGtrRust6fk300etrhD2iEeIkeuU7ugFhS
oLYsTxtWk58JsCp+AaNaUU4L+0elpOsPa3AFlwuGsyuGna57dasvmOSBtYlNLQXlHSr5xgj/XkG+
kqUk5FtQ+2OOHhdp18/hTv3iRqFcSSNqDoQCMN2nl8C1CuVVgdL3gfFyUA/kzBYaciZ53hEQYIp8
soAHdfHDRSaooBDkjjoYd4ueEFAzmoD7RkVxeuPkU0DOtzVQzrFeutVIOUwnFo4eHP8Ze2p6kjLV
PgkBcpsoM0dWllC/k2DdeG7R8mchAKDxJfmIhXckywArFfnKOdUTbgMC7y/e1cWrLWX1QqO4jGmu
BeUSJF24MpE0Py59tkir71m41ba/G/+2JSgvk4rLiSp+C3BV5uVZpA4yDp7Kimu09rstYFVARzSd
J0D5CH7gKko2bsa62ulyypLH7r0+WfWmgTQ/DwVEaMviJm0xxmj6NRoXpktZcZgyQHK4SyYZ5Sfu
KkgeL2jsrB1EyZlGnv+ynGgXtyvp92gxNESds63m5w4P7WK8xlk+XJdby61aZysTFnJXS3WNIECj
hqUn94N0pm4ZaclO+qTp2f0e+okFlHdslzQPjY8e4Rnc0N8tB7wdoDTvJ2uDcH/94yGh0qnHNlBc
5b3cXJpJ23PFp8USaD/nvmM6hWweigwkB/HzqnBVey6i0rn70uqv6wOJ51EQJl1Kof4B1D8HJhGC
kbkzu8SGOowBe8PPqYf/9uCu6rYhjIUOQPTp7Lqb99fCotDsAu70CWjnI/7dW84Jbq17XbtZ1Aml
205Tcd74selxXVEWPNLIeaDZPYM/addFnBPTEaxjloPxrfJoCGuOX6389mNYNJ3oyk6vs0/iT/mb
jg7MqlE8TzV0QSvo5dR0WrYcDGDOTfcP+SC/rxoK7v7tcZ3b5i8+DSYWGehb2NXupS8td7MEyl4x
gtHQDWXL92dV19eiv4D96cvS95FwGkGqPX/sG7vYoHpbodEDaGl7NaOWPU0S5ClSw7bBSU8Yk5UW
fo7tu1H19NzhkIn0TwZilQ4pWdYEvrkUCDS3p3iHTlUtAVU89P7hRN4U/0JoZDZLfMAv1WcbZzOv
SrPjvvhvm+xX1A/aKenY4Ax2um3NolPRoQUGIkV/tcB3Z2+2/gQZ3hgGXkwplAEG2E4SjASlfiKc
cDKWxJMaaSmU/4SplwPbCn6UM4t1gVVOFbYJUz88tpisvydwls6X2BXD7bHHl0iyjnQy/S9q5pk/
UGp5rfolLcinmaucL/UbH3JwGYb6f0CHMQ2dn8IcVD/PDcDZTOrwIavyOXdRW/C8Ut4hCwwzLKH8
4+6kdQ2oUzYQB6sGzaYJJxyOqwY8EH4SRgMaTzMQ4hvn+eKQoZdG8wCR+As6iK2lt1pkDQHikGOs
3c8Yc0BSec6lwjvlj7RwhGAubi54GIcYDkKqD6HM9Sj46hqUAsWdEC0vaY86TX05eRBHxe+ob6ue
YBBS35TkBeQhQkQbR+g1QJlJ5jbc4v3lb5lYSMKmHYH13oVErdokg3F/htgxh9W68DHoyxeKX68Y
06b0m8h6A4rjm4GixKqStyiTRb17rqa6i62ekHp8YOksyaVJrXdQB5AZBKdMPH3cTgFDwlc1qK+e
sckHV+h9eRZumx7PyXXB5BGSKjrqxBGCUQO2m+GLLMXSggiPiyCUWeYVDm0+4tvy+2Vb460/JKkH
R2lTPfSWc2f3SMGpLdpbaMMJoNCGAqwC8rfbSMIVSeiBxpmuKHBgJ15JSfcIFvolFNp0gUEZPS9O
t3aRxwLcjywgB2m4WD9D2HNLDAFutk7kA67sPnONAFUKP2PV6bzD29w/Mst/NqmNIWA/2xi3fMN+
8YrPW2GzSITtqCA2c3aNSVSTJZ+i11QRyynqgO5mieRp777CJuyCqsUeejSL6B8+mrSeUgy4gqFP
XMe4cym8KVQ1JYSQom4Bfnrf+RiWJ8DuMAuiYt9Z3XGZLY3il2DH/Ql7FY8TXdqSgwgOKGrVSD1D
V/oDYsuShApbPjzTH6cpkq0kTcKzsPFem7diGkAsqujeqNVrfqxcCsR8LqX2ukYs3q0u511xkU17
Mt5aHtGL2TFNNrZ1Z8HiNIvPlHYoXd7nyV3YlLqIIbASdlBSweACIp6u9hkFHlPqDEXIN0EWTgcK
cTDPbbmhumNlYZgxy7LmtiHKcsrbDApw7XLZ2WpJab9BJQARTA2dexBl+MrclvJQ1l08JZ07Fqt4
NRNVb6mvTyX6QalprkU/27WPdFpGe0eO5cNSAza1rczm2K+iRkVVijncWWYdw8JzsUsWaMkctcKL
StB7a5b3lD68LxLAfMdjriKMZfGwUS1sM1qJ/k9VQGLUaSrwNRwSxaZkODjtIY2I5yzN0rY9hBzS
ta9pNc4NdauqKyRJUxKRGZjTLZOUcoFNWROxEERGWgO3CL2fxOUaqqH6UFzLAAU0/GxXOZ8K3d+h
nkL3DyMDAGrQbXBg/8pUpVLtqM75O2U6XE4pi4aQdumkZhiM+9WButIIxu1QRw5EOkcGZIUs2EB7
aRTkYjASkeyRt/oRrThDLt64/SAArEKhxV7sOlFOb2up266o8XCI4CfLgYJlhAMTL9jSWh82uFFG
5Ii5VNdz27s+ZhTuiIdzdhLU6KB2WT/iRTmTwgt1QxDswI7DmMPKK1fgCQBiXu2IJSr2JynIcWFf
BsQqvJ6a8wqMRb6X8Lqvi4NtmrurOdbviMYWSEg5L9ejEf8DVD8bWzIOIynE8sSEeW/UldPT1QoY
TZAdowYrOxdBjidiuk5XVbiv23R8MnL8l8eVU03D25G9WEUgI0R8XJ7fblBXsEyXM2WzATfNMSmu
ixnwWFjBaP0/U/GDmBI3IGW/Ilo0AZk+Lk7vkTi5kzB9R+/JzYpdhjfIH63w7OCGc1bmoteZkupR
PcD2FERRZ4OcIhLKeCdL+zgW+njSiG967TJujTGj/2KepiJHbxm1XJwV8rJ5GsjbaulnM9x47Xqh
PIUlmStpl3NGoCLiS6uzsi0K4E8Y8I/K8GSJrBLCnXLVMIBSxYqIjlHc+7IDrR61MP+gDfdWxxe0
P1LzXJilT4uQfaI0uZCOSRiuX6rE7ln45h1kAAEqlwLX4Q0WYhyhyVRCdbsJt00u+4Rs//06aWxE
ONBc+wPB1FkafI/u1wjJwpDYTRLBH1IpGP07qpv9jB2TUoAVLsEwe85HqEeoNIpcAXs2p8B4xGct
K08uujhFncWVQFURxxzfhcrO0+pU9STg4b1xATmc+bzES2ZcX+kESGHwtorOtEnI60uoCHniSGk8
moYdm+FtDkWdpJ6ZgC6ARPDzdz7OP8+wBpyDmQir/HksK+fMPFK9vIsYNLLTM5bStEfKK1yx3q5e
qdTBP2IoBi7lTk3T0p1EHq0qyLfc0aVjeNCZirXgvTN5rCdDZH/eMCNOE0RjxAlHPqRefuzJvDYc
SwQHpxo+/OvBt37Ud9pG0nMrKNt5jdHOjWuFoRMYJMvaNfg6Lnvl+fNOXp+1hZEoNzxMwEQPX9a7
ET2Ahi74vDTABTPmdGY1gzPuA6ByOVYGwmk4t/MHG/VHYeQP3GEX/B0J+GEp8EZks16wWuVbvnqn
Q1n4m+iEgR+X3D7eUTH6ZQYVIyoavWVzbkiL2scJrpIEbXv804cHQ7Ps1m3cRd0cV8dJyZSptnGO
0D0ZnaX4Es4CtC5uJiTNGK+Orq56jaSV60nWTJMlzYhl0nxhQs8pOa8rycwZgwKGNMY6MJxm0yv/
X0SXDXUTk/Glag92sw0NUMR+U8U5t1OQrfI4NtPwCBTa2Y7wbURfqU2GynYmmC3ncPweBX3slVk6
UR8ocqiZJ5jthcJbhfZ2AAvTbPN6PLj0+z7BexZPYmkl0bRr1q/3pk6WEf9YomjWM8OBtEiVJMvp
/8dTsnDQo1lzxt9TvU2Rkh1hA5nDlzzuYMz2fyFSd1nUck10DNcShzWTnCgfGV7nFy8ynqbQrbXj
HomDIk2afMcFJFYW97ivgTc/U37uGElGf6IDHSk4hF6GlyUl/tGKicBeLOr4nym0MAol0msEWyAc
hy92f0nN6eGGveMC1R+3ecAYNJTeIKfm4oglIFOLiExhCk0apClKdDx4tOPqc5ywbXKooT6kndw+
mi6sv0QJmcvJTz8fqAoJuiNnH1Ngc+jfZv9mmkjt0h4ySQ1ufJEUvLtk+D3VloUdt1ukWyw8+80d
S4RGDPVNlOs+IwocD8AYcdkS8aTyLXORVNl/0I/zK/8LXL8Y7pmu5nTdpVc7TAwZj5ZdrOP1J+Yv
TGOUKUPMoo0a1Tz0iOMN9l4l1YEAmXzs0Y/djS7B96Qd1/BlzA/irMPphILRiaUz8nqWnEWfjHFX
LJUxEOBXU0qYxJiGGTKQSvq/RKXGspn0icTH2B9OjnhyAbe6m52yrf6LsUImSTukvaot6V/eVvhg
pfgi6NtDJzY7tAShjdnS+ns4RO/PAGQ6wzTiAiD2A6ZsfBscP4waRTGliIMpttpvWRvvWl8vEdWG
PcRJsp+n5VIsMkHD9gDws6jjivRlfwyiIgI5aLstj7XPPF/7+kMRFnS6vADRGTGHyI04YJP5bCZ6
uW13K1/wk65ClCtJdrxIanPsdfOH5W5jPNDjjwSXM6nACICzMzXruQ6VOJGelBO4WwrZS/3fPY89
ZOr+bmVKPIDXsifdufsfGp/z2dZIZof3XXgKIXVLOnc8hJIAiWm+pf6iBMvQWQyqkpCQ5dkgdG9P
7aeQisvRx0Oya8DFAF6Mj3rmuE/caRXM65XBlXpZ+FtbS1XfhGw16w7TA4PWwO5+CvFvpMjELK85
SrDHt10LQaW6LtWdwMmfT+hFRygU1LjHsNEuk9OqF13NyLXP5gjpBYepzWWTn5PR7SghGyJTQxkh
riOX23I4xzHd8PmfqUSHdk4Vle5KSW7t1IAEBLe0R1IZs+Ubb56VTiM67wZNQh+6mqczpHXuqqJ5
DosoIsUpLUnh6tfoOpzr0qx0uUSqrPzbFQ6pwryuYIKcASmtV8fmhFCEDNeRseJ/R3sufat7Fr1f
OKqKpEnGVaD9fpaEODqsnRQmcIa6GQC3nAvcH4HIxd8FQZx9WquolEYZkTddvBOkILv2QGBQsFrK
M/EEo00yD2AOdjp2l0nnb9vf+jRMLgWigN8hzOYIcWYlMgZhiSWOVI8cPWbzuqihu/dqayORok+d
Nmi0CeXFna/7LiPMULBRyISC9DQSKHQeZ4MTgvagXRl7z02cUalMzyh7tKmh3EdGMcwvCZLqMfqI
K5AQ45MvRJNQF+aU8lIYMdeTSZbGdIt+JQyl4j8PmOjaAZtyjP0/CCG3vjZfKVE3TeIOwN0M3tjA
VImLydr0L9y1FZq3+Pe5Md+NAL21vw4NM7lFYTyYmVskeuoQ+99v0KulZnyGMGTL2blIvRlhMNTt
TqkQHz4Tw/jFHpN3i76z0hMkfBc2kbgYKUI3IG1BraQbFGtWZRT+xYCHqHHQGk4lMHrF86jcg0Cf
bfnQ4/W7pCg2KYUejdcm/C258jU4VeRjmTpUMFUszSwlI3yMfrTEmJ2DtcpGiNJbVqiV3JgQ/B/w
xj8Bvqxjc6XgOTYoXQyglmy/FFounJZMaJ/XAcEiELzhIj9u3mXRT6WAiovgvYeTRTlNvxwutFyu
4hBorSoS6ZIXDuVRkVy/u3Fx9XVx2ShaAi1h4RMdKX71WLsnQ0KIk5VU7U2TGn+BALGpR37J0ecy
8gJMvXQ3Be86ZmD2lB3OkSPsAOQ3SN4j4gs5X00EC2D4xnOstkADqbvmz5PrZG/HFTGEpd4awPz5
wJAiF0WNsdO+E80ARzUJ+xPMB0+y+MBOQM3oAr/leeTIKuTXiixiYQiZUljHkp6Wk9tb3/GcC3LO
ozDDqu6KzuaVUwjhUSEujiSbNRhj51W+n883CncAf79QmbWOKbCUtIIWFZ1cQhHyITuEERhN+RNx
FobHEu9sqGpVs5X6F99x/Ct1VJN3cI/2yVL4U9JmnZMzluIQOTDeRZ2uqmVDChTD1AcBqb8vYo9c
mHZWd9X3LfJC5aMjrNXTN7G+HYdun70SfeqfSXtGYQee7IauHkAaZ196qbQ/UxwwA768iO9ou+8q
I6JyeNXfKj+OT2gx6jTEFg/7SZuHnb1eSEJ9vo+Xn8vb1/c3FsrbfljPLJLVKS24rD9uvMK1S48h
MW2tH50Rt4F5SfUZIXUhebYjunDJxhvkxHFIkiLZ0gDO/eGCacP86VxaAGYgNHLSVq4nTcAKBpc/
U+aAGdGqhlP4D4eDZLVbkmsu2Kp0fpWAylCxnQLOGiy3yo2LO91159XTPl9hvKWzYwiH497QavXA
C8PevxHzmEyj0RCEiynQJCuTnuuhyEmmh76dDCI2nDX98mgFQA6NbkWcspxupmONbsQEMyKDObXv
0z77zqho/KHnBD3NmVzQT4P70prhd65HuNxEJ/fynzbLxYUNNjlHGWUYqBRrhJoqc3JtdydT5zG2
D3FdraoUaj5sqnLBQztHNnWDPKKfwT9MvttplZnjrMHXHA/qHoOheD/W4riL+BMfkr9YQ3V0Zrfu
fCAuSLkNix62O78BjXpApVcvOM20I53RuIIWNl0kl390vyi0ktyf34hh4S70CEp0FlfFWGjaccLO
CmaP9RyBJFBFISvVSc1YqgV4DzA5LG3isU4fnDXfewtJa8gjmF9D3J0s7entDV7i4zVKsNCyfn8k
spwV9/YBGKW58dQmcefxxi9j6geEbhf3+Nt9iUqW84lqxphuqRb5AkGBSG4tCiSeYiQMLCGYGrWA
kYdYqnqWV80CzUhaXW7tZLW7Ec3ZcaY+mmbZZeFGCkUw5An4Zg1Ty+ZdTsJ7cts36eHM+z5vAh9k
QrdjBWz833nJ3iNWvY8JCMFUmYDV08wI+IQHuLiNYzUb7q68MOJcBzPSscToF6d/pirOMOHMyxFM
x73RYC118+x5rWQJHkzrJ1raYL92dH9GcSgG+LQrXBXFE21BdzxZ+CRFWfuFgHAr4OJeaGfA7XHe
9qEGEIivVcrLfcC3I76oCtVCARTGdIQK2K2zE3r/8lzz1BlefupjrQjGk+bQoMWCIwG7mMW6eYrI
x98BlPt8BBfqeBKYM/ir3yMXmqLmZxgTox9hpsLnoZrBJZ27Ycf+r6eLeyKCZEu2dH8Y73/6DW2g
sEo6a62vFX3v0T510LEv4EW4MEOxKkH2Zwc/c0/gJaVEFL/ZTfr7B3GwjCR/Myuu0qiGts3hQffZ
v1ySg8vnIkEG1Q7J2bDExQ8CkPTNYacNgtxqz2C7wZWwCHwklYJdknmM9eR96sgeUUXE9tMLl2yn
n0310TaSFJg5eUhU5zdC5YYWRDUoIicAQU+0A/vJ2smkUM4M1HFqqsi7jFE1FhVH/C8//YCjQ9K7
1P1zk6pg3wrqhm2d8r0ZgrsSgG4PzpSkmTmUYlC8CiVTaZUS9dcT+P5dvNn7/RO41UqLVtFfgTnX
M0kPB4et+8dq31m5zFvidbjs9/CeU/Nr7A3y29TWX2bWToiwVINupnyD1zhqJZCF6F7x+3A4z4uB
qrUmBJ7HmvrcTfE40u6U2PKDSl3JNSgc53oQTNUmgENckNI8chrRzfSE3SnEr6C/wZZMzrj7qcp4
VrZCztQ4h71yqCwWSYHjoo0RvK/k5EKJ/8qUZkUQRZxHQfFp+0m99A5g+MwaJP3nXLA+AuONGBpa
wD0QDc2/Dr9b3QmWi9IlFmoyIFn1U+Lc1wZ2kCCKZEfDWjclLXHgeWbatd+Vf9tvY4wDYFEKU5Js
6SUt8yXtF0Ozjp9VVA5Ouaha+XHjW75KqO8PF2uJ0IWks4TsRB7ZxcjZKA16W+/4oS1klN+2vJV0
23hhnYE4utVkm88yTxeJ90chb7pz0ofuy5sw4AUwgRPkRzRuaDkOn8VYtXOXZwy6hZRtTH5N6nIy
Fev4sZ2aCQRksqrLNrLStpUpgr3kwQT8kc9gIrqYp+meVzIll7Or7gxj9Vxgys11mD9qom2YYwrI
U7Uek75t4HE4/lLAC0Ui2IG2oV6PVeMVGP4AtL225MYC65i99xXrBMzlxVeIy44eztV5ziRDXVZ9
xUzRBoc5L3NdX8gBxPz9OOEkZWxpN5iKa+XVM7EpCJcoUjnKyYrNCiNkyfC958h1O06jIHI9B/Q=
`protect end_protected
