--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
lYrygpN2r6+0f07cHiD+2pT9jHa8UxrTnhsBoowy7C/87YG+AHHRttfUYp5o1xkOn/r1salmAp+8
tfOQsV+NwDkXVC2VrCzoDL6eMIkX9OJ/P2PWEae3vb4Zr6m+iKv+MIyk6r5Qj39xb+pn+4Gcr39G
Hm6UJ0JTipcSWlJQ/UU/NU8rfooVocvGTamkbrUb7vFfJf7c3WmoN1hTqDGU9ci2NYVOyynOeYSq
Zb9SzzAu5G88b1Comip7QTKt4x4hzDTTSgCE+C3lTP+/WB4aEW/56LvUSbbLtLQ53BwrFcyfm+G4
oTklmJp7bmJCDVlj1eGYfhdakzSXjmmTELLhyw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="fs59I1Hr2PnTeNpuXWjCvM0WV9nahVs5tNApVOVEWaQ="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
MgYysmYEmxLEFPcoQslPhgdiOAtzuqen45kucOV7atBAL3j3wVd+DrouNk9b9eBBk8HH56xjNAYy
xvu4j/M5qMfmV4s/Bg/PZF6wvX66R7yi+XnYtc46c7br+H6eRZ4HNWH5NLvwOhOu7NOemzGw5US7
lV/adFtomQvOjJaTqMfMTng+cMs4KxQTaSOPeHk0lI3i1OZjG1LpIWtfx4g1zrbBDU11BFNcnA9Q
TxtsITQsQToipvpHm23iT84HaOXRIJRXtauE+v+EkFrI0bzjcJdWwy06Hr9YOw/ZAgZRGqIPhf3f
jU8BsX3DcDyCK/L2xFtNr0lsEEEOukxd+KUSzg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="DD+p9Ajk1a/86YYf7Ji9EPgnWm8BYE/0NUGPz2sS9ns="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3264)
`protect data_block
DBVmJ0/nXQlg1Q7gDWDjwDNVS+OdpPHVROLK4UrNNZxVD7GZVATVIcGBsfoaoayV2vkyQPNdPspA
vItX++cdO31bzqHK0ID4HciM7oIN+m7z5NhhCgUOXAwwi5SvsMIKCpt0xVdi2qTo/8czOTLFia1/
btQFjeC+7jN70GKVhgyCc2fqC5r6lfSiv2zGLhuOVR3DcFMHnBaTqkwv8fIqAPvkTw3QqTDkuBg3
LIB1UzqlW1c+Kke1S7Y/vzcKrgKKvYWQOtOMV6KjmPGqnuSvZKBwXHpchnSD4wIOTf0WrULlGVpl
1q40dglIaNUYc65saukQxFPdKjyABIfG/mcpJrLty3v/K5B1Y+ONvHa+dolNt7oB0nwpEq8n3mzl
NdzlZJipxyNIXyf6Ut1E2aRilvErMujfDlSoc3HPhc/iwYTPOWuOqoxRvfyI1LhLcjFTeJlB7Uo9
Dbe488dZWJPpC8zV01lbcIkzDZqfxuF8d5CRRZd4oV8CtJ+dUBg3JIpdZnL5VP+HUW1Bsde68NhO
Wl6F4qPE+GP08Vz+t0q2Arsb4v6Wd3jOEb+K0q+gEN+ntI1qPrspgh7u1JHkGu30ZD5nwvs4zxMf
H3d/r7Xfh59F87a0PMkU3eboM8IZk88BMQ6OP80Nvawc6VPyMUJWQAWO3h93YUtNiYNxQJgW2XPi
TNltOKndhXVemfS3wHjAbLnbVgL7C8f3fhV8pIaaLHvdUt7fELQs2f2RhFpa7TrxOataDRKqRxvb
NoXLupz4EKmgmnnSUlDM+3FRnSkGKjR2EobGS1WHZS71cZ+cV3kIJuT+cElQlsJno1kDx1kKGoaZ
bndFaH6mt+Z/Ngy5cGjHo36l93owDNUppLVzgmE9XcdglHfJUehWvhWoep7ie/xae272bAU9HcDh
L0rwjUSF/Lx47r+EPBbfxDleVhxXfZL8Ub9ed4QSf+o0AsH9l3o4iwTLW3b3k2P4LbIAo3mRYtMN
D3Xo2sEvy+k9fjSArhQS8O3rxsTNfNLQ+zDXCWB+0JHlqPybjeNmdFQ1Sr7V7bIum8Vb5dAa/wr0
7sXLjRPC1/qOd3cnkLUfcOtlRDF/KdbYwqaO0HYaOIdxkJIaZksUDDdyMC6Hp1+FktmRgDYGzPOo
vZL5++P1dkmDft+xqaqFHvUuVNLc+oOfQEUsV3EeoptCqFj2BbbD+KqwwHx97VFPS95NxrrXCa+z
fnafZWEVVs+no87JCYcdPhC1r+k7OL+nyKvK9aJaTig+tMNbftlog9BE735JkCYbdDMVOnIaOJLo
EDaUSjZy6+1HDCnDMp2fVucVMNE5QJpYeAWjGL4UIuBevxJCamI/RaiLjf8zCueZYzrkbOrj29sG
+6LW0G+9mVN7tHKG1nPqooXEPxh6HPzNS9i+LSadtx8wd08Uuw5tB1ykyAG0lXZRBNF0rmIEvTfS
l9Z2ugTQQvMiQ0FR1EFmExQosQIZigyV54r7Q46x3opt5p1a67qdTd5aaYK4AUV3hGzb2wfseFLg
lD9unWW+MtUwaLHxp1SE8c6lVnjmevVXHSD8JxEZY39Khj5NIi8T+VekcVBKk8gkwriw/zlohRLW
vgBsLiLDHApnXkWjr32q9izl2Ko2XXqH5BTP+tRv7jDipdSaAG+FHuaRvupVrlJhhE5igiQoJfbR
Pml8pmBtvgobZGrH5hOK/Fsj9FwX8E3AK6O9NUcVDFK3bn3h2MavH2NR3Jgxa4JNBsnemcMIcKw/
N1u5hNCV1gzQexMQx6pDvsXlZKkbJljKodyOjt5VBkJXCtPa3sfMwNad6n0z2HGQAP7SuLpGr+1L
H6TorkoO7lGkm/iDn+fD9OJbH55VY5zBQZY8jS18DwKJL0nYVLqQhfRmIWKDMW/sfFXuFERniCB5
LwhbBb7b0W/LQ/VaN97OoVt21ExAIxB1/ja+Us7PhEV043PeYcwW486Ln9PISd3qnur30L2xAF9G
0Str69USsePjeCHbisJdCwBkQqZmRgJwAZG1Rl2kYBCmYpzcW1EuXr6amIwOUZ+504P09qoCJgyS
6oMqdnAze+qk2PAU9MMPPN3hAXkVZ9EGh9LznKsv9Ma30/KoNCXWCRq3LkzFz8XYNdivK2gtU5eL
diElMSKYqVQo7f5U7YCU1E34vNR1zk2II79WzcFHzOqSC+7YBmEy69ZVkY0fTzNz6Ij1rYQmpHCP
mjFdkPTxTg7rFP3X8TOWAgoTm4+8ZRrA899+EsnvlHikR8/Dkz6dUJ5c8yoXh/sudXVyM9Conc42
UwxgwQ0vG05Jesx8z8mq4uU9emXFb5GAu2I8ljfee5X3pu56i5dxFxPZ20LVwN6Ve2AnUvLT/PwZ
JZF6QrO023PIqOgkVZuK6ti7u30LHXZQNlBY1PzJHqJr7GWBAV0qf1Wna5m+V09AIz8rkAIvO6Ty
P9a+CyCRSw8/yQVaWpUZQziFTsd0/Cp1Jhg3WGM8d7yJgQTX0Oq+21JhT/tdUifjOu7apb8l+4tR
LPfhGzhmAmcXPuDw7L/U9jE6J4a8OG8b5U0AaBB5E54IWvc8A/PMHgAnuzcBdCqVGUroxhX9ZMZG
SCfyql/cUwWpBF34XaYlj5Nr5R3fPv5Ezxwc09nsoSf2NCL6HkRJLn76aHrRY/ObCundqqFqwQxs
jYI35kleXx0LRos6mBGhVNaTrQ1Zb0FCydOOFLgj0dk1W7RnLk44P9QJGpEI+8yJmF7Dt5pCBKM+
fwQGW367FAQ4FWnZGYxY6hcgcAKVLHLadpiS1XQaBSwGY/7eCsD147V3RjMy/yJ3loKBalrTLqXm
mWj1UzOwbpe6p6PxD4/LrHdLVL/SKlJB9oRKZB53QiB53N+CkeKymWIJr/rAF+dR4qN12MjDiqKs
OqnyNDTOnf2ZT1SKNVj66IzDFbBm3Sz6N3qY3flYJao+dizFAIgAlZinJ/YR5bNk/Ux3NpvjDfqT
Oz5veep/YMxPrcGoIqV8gxGTjpf2/FC5AXENDt6MV1i5g0ueMFVTy1gFTdQVN+32XUn2dBbewUt0
QTQ+dI/v/wo6a0ebZLSmp3yf9c9kEC+cPzUZOD9QBYuivqkLAnDL+TVzKORHQY/xud6MRgI1kOow
hrnq4qU+jocA1dOIdonhSiTd0OYs+qBKfGUb6t+g/83VbPBtvlAnZ64ynPLtHy+htbJdHgBjT3ox
mWawTFBRPgMAewLsHnv5CLAIL8hq+KkKcYMqoGJmRRBH4Re0qW7l47kkQpCQ3jEDVjrAZSNPCEY2
cb4ZO4GgC32U9Zqcm4ICxG8mdEYZvu6cdvBvM/sObmPTV9PkrxHi6RkdqpXfcyBd224RkBIcCKkx
JDh/PB/J6DLks5LUNA9G4/bDm+dc0/VTkv4hiQicO3ZRgZt8jIwK6YUhYXf9/zRoFGOiAplUKk+m
juiyAIyu+5LIISGCx630nsuWGeqxQ+Qf172CUZ0OuRWh6+fVonhxBZ2EhWPn3r+HQzQmu0ZteaVr
F5kie/dXcdDhlS0bm6CxSFr6JlZrQog07DPGWU7MgSvIqfD0G+euUomPOVgjV8ZRFV83RAhZZ6o2
H9Vvvn9vTxYYi71SwW35hw+0DUDvhKwlLaWqT5F1otPRvG2i9Z55L7ssxwHTzG75NE/C6APpxS7P
NZ6CGAb4yyBN26jnM2aqx0WBBvnt26p0+5z5ETlNcwLBC6BfX9khnnWG70Z9Pb6bmJU7weXaCf1N
heFAQZ8xLvxRCkvD1bMFPwYdiCqe0Nvm+QFg/Oyahpv3Cu7+PR4nwaX4CJc0rf7I20dn+ny+Zk0b
9IG8uU2iGPnc5WwCX52dkue6Jf9BRlj7VH/WxCW+6ADkdtvYnOJ8SvvuVFHww5NnkzZ3oNFhb8GL
kqWpw/jePh0wC4yxBDC6+h9MR0mf2LSBeNilvwI/N+YQ58cmCbpW1+dJGjOYDiT6/RmlZwaSc3tc
ms71IACvFV3UwoPRXwd9BJOhrgXmbpqg5wEt/S5iqHv/XuwKsWprJkLPuApYIyVPfC4Fi4/X6jzK
8RComfzESOyyYppQYg8ZHZpa0D0ru0pVT4UJJPr7Q+IVyNljVFgPElkhA2E2CLwwP/D5pFTFU2q+
JUJ6C35a0HosCpMKnOLiaOnO/4VM6gk1CajLuGfqYWQmyZt3hiyeFgxWaQ6NFO5qkS2cdg6ilfJk
HonkAm2BwSdK1QavDDKGFGcw6aOwQa2Dtj9092JTdOpsIH0VyGYBeZupUtqIODwcmn5v8HfM9fJH
tdUsGAqbn6TemnlZL5SiBJEzZNSNUn2Fp3PJKVyf6L7S12gFMouPLa0+Ro6lYzGBQ8ebCPFHllMt
KVIFo0nWQ4+KSDDOyMeq
`protect end_protected
