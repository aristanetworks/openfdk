--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Z3IDADKqhF9j5jD9JGxiz5cc+3TER7zMdZX/7vE9NGkdAurj1rgJtj0gwD9G+MHxCMF8AztQOBRV
NEZNAQLw6vQzQZUkt5VPwtEnhxAypywRRdzMyMhT1Y+Ywnqn8d0X/iAbJf5FtjOPl2oS3UEHOORj
WJ9GsrBb3yh7aC8luK9HzJSTHzQ0l5v3Y52e2LjtYAAskA0S4jB1AJRMdy8bQs3o8tphv6COA97h
OVb65/U8PtfV4VzxYroKKbgRgyiafp6GDZP8qxCjGFUTlORduFQbghxo1A3FzvhhIdaWuGGkdvp1
MDo6gzGyP3GJEuioTFsDzDFZ77I6XvQPo1j3DQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="jLJewFyI587NsGrexG5niwQCD2l84Hn9t1uGN04+Rgs="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
eKTzW5V/224PdesfEms/omtx0KF/1qMdgO/kxJDwEReX1s4XgwbB5JSTmmk88VZJik3dVipoaonk
NB5MveLcN3Xm2LWch9DF9U4ItLXIrsInrKmk+GsCLqgdZCCWqc9UTfcjKs+E175ztlscFmhlCaHo
XWrGsSl9TJdrURqD1MGmHFkNxTOm9VxVr43y2CWyixNJ0gHd9Oa/2PKBzQjMG84OToa+JCv0l3FT
95Xdu2VWGa0yAa3rdmQnPjtbUCasOt5a8oLFDTteNZ2RPbJ/ScMm9Divqk8Rrh7seyU2ErrXUxm9
kkoYvxsJzS0g3z+enF/RfeVAkKMzWTew9dfW3w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="eNyKL0VuyAUJnKnkIjrXa7AEcvlLB7/+zs5I7erYGfM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6032)
`protect data_block
9eabcTxILzF8QdBVObUtpA578hXy2myLhGJU3zh1Xpblv1l3jogKoRBrubM3kdurPpBUP1ZZX8N6
HFLLCBAI/XrN7YxmKN+AksozgBZYgeOgxFJWcCz0ERuhZKUzSCsR82T5w0cgYvB1JHYkIruzo05X
PTwUgFCuMNkadLAhbEt8sIcCTsi6YEZtfFGa4Lc0EmLBqYYh6VDQM+dEteulahO2lwfoIqyzPWwS
3WTj0wy7I8Zv3YP0mftwyVCNG0EDcrHYgvSVCrPy8jUjtxGKPFam3Yc+8SvUZi8V7yJbCq8X5Jia
OjINBCiWmzZoIffHWmpbpCiHCAj8i4DxsLmZJxBPDrpl2HOMUuWKwLNTbEU81BkSu/tKx9YWO0yq
rvYaPAD5d7jT+2NBjWNR+7mTKvbw8IwdaHkuDIt1uP9xQaEeTP4N5khnOMByonnA/KGBnV6Qout/
0qn2Ik/3D9wld7XObtJiQ0ZLIn2yk1VVwcKhxUHe9Fc/Tx/xjTHAIBLrkaRguvkUeRdCKejxaPKo
OYMbx0yC9sn7F2BAi57hBBPgfSLiJ3A9eoALQd7weeRiyhyri8UJOQJG/RvR+QMfRAddZ5BoAJkt
KEA6tdH9erRvUpSP120hZ3k5qJFpcQAo7DcLJIvGV+1h8YlELiHjC8vRYE5knZVantanVlDeS6Wo
W0vNCnX6hpKvilEej54vwViGr6zwPOYVqFDowsifg01tzUNq5BpdCsjk2taWaZ8bgRHpDNvO/ooc
OuOH1KQNshUK9PkvQqTeZHZjdiR1dWWi+nRjWv7AdQQ9l90BzgvkWxK3hqM964AFq6Bhgq+Mh5hN
jwhrk9oTuZFhr3PHBhAiog/CMrW9g5yB/tiyjCIWRc818bZjxJjP2UT5t+J/oFCPui+QASCO3J9l
Ob1J7PqXVg6VbYZXNMgYzDQMeosLsqI8nMMnG4cTRVPm3quCe8bLw9y44cZW99IS0iWOXHILFOIn
YQK+YxS5SOVN5tSThboFGvw/53SZDCY5crZ0jJqdSrh5qpCvwggY6L4tOyMTmoT5oPcG5m2UQaED
mtnyzOqJwC6Hr3D6RNp1SKzHXse+Rh8VjUimiOvCW9A1Y7k2k5YDQpufaN8axyYlqwEoylo0fWL8
Zjhnq8BlbBVIn/et+1ORDxMe0rmoHz/AselHz3YEzzi/FIdmgG6TiXBJqUyaykoJu0UN1lI0o5g2
JFiuAsvlvEnyE4eRVFHjKR0Ia5BJcF722BD5kHOuOczfPqIspkv+YeGJVaCucPjFrsAw6PhxRe3o
0ddjuBW0hSsY4uLWf4rtYitmCq/QnMe0JAw9aC+1UFVQy3eidBee4CsQa1JgdeJAYUf3sNixHkgM
8BSr4/gGxinkKOxNnAeVYwFd94jU3gKeJ1Wu4J8pTWh0sl2Yg9n+yAUfWzx1dcejAM6BVH8voAOg
m/6n92aFjgB4w62r4DUJOJ8IQeaEewvmvA5D8IlbOG2j0NHopcGkMhCGMUPvYglciI77c09CleIE
C3kqL7Z5X90CmDnVw8eJHs697YWtzXpj2j5eom1QeQRM93BRK521s4dnc7UebCaQi+v97GoHGbId
J45zVTp4Uln7KGU/x0qAjR00CxA02zT55t0muVpKxQspKXsAWl+r/teCfq5z+cY1H6U5Sm3H7EbW
FP8rfpdCHu3OedhulQjZA0P5jLOrZjyvHjPMPuDl0UTPKLK1cEtYlSXtauMlJd/pipZgI93Pzx9y
fjx6dAL4NdOb1Aq6GHLrA+Hs3sZzoXFw42J0AXkBTnLF6yaQWa+fgy2EuMCHHpYv3MP3L5i+uz2u
7jqPlfEVflGfrIZ1cPZzSuAEVAnhpW3RR+0iJqntAoPHquLdYnq6EPo5t4tEBKu3oaJQzn+LaVBm
ugWyKsyc31ZUiWOwGGptRyOrZ/5mHT0RvheEL09qoqM2UNcgo7PnaMHfFfn5MmRc5xjsUvhQ5PtK
wDyMeJ1cnE3MkNuhHlL5b3XhGTVVUVP7orVWgRfRSQdiOEok7Ppg70s8twaj0DH4KTCsb5Ii8A7k
EuDc7ACu5Razflo2gV8j7ww/vgTh2FmnKS522heusD1lBmtNbdo+RRKH71sK3L9uNxzh1pYWWtGE
xi5Oi2jH18dSWBDqBzOFH+ipxqqqHyScP8n/zihhViaGdba31Afzhnxr8kKRimWFSjlThY0zONdN
Gdi0i9mbJBFBdumXPS3B+YorJb/SD4VkRpAaDjtX/+o1n70gpN939IfU0MAZPVUM2olw8r8yq3yI
EM7ZAFscHR+XeHyd93y1rFJLIUC5y9uXFdbgxz7xCGb+eP+lQrFoSAR1lKr/EO30MJfCq7ITJbdU
hFf6+r+AWw+QheNyULLf3SPfivi2dDWl8iM1Mv5oPvw0BJ/zXXmGklvPVOqor5gZSMwStqsHSBIh
hcMnfcTW6JVfk9CBEMN5S7C08tAXqmTRFq63Xf/E1SnwJCQMJA464HPTBGYl8B3+57kj/ojrk5Cq
w3HYdmzdSANP6fv3MTy374zAcJEHVjBEbTHpwkQnquj6QcX28/OG+Ro0FvxrY6VI6hmYcIDx8CJl
J2k0eFlhYe/y3jq+opSsiExFVJXr1OAZcRc9zS62X4KAeZzxr25uy4TeWsL9wwLiYAov8cMZ91z8
f6ZMVQSe8MVZWkaEUd7D90VesWlIKhDo09AHmcsplWodDCHYnGdS53nM60HiC2Kfj4MlYXrnhT/z
xl768P3p/bnN5FT3n3JRSmKt7ARY1VmTKhTb021laUfI2y8m1GxjN6eSO/aQ2J+SIeuZy0sHHS/z
JpjGvWmYhdPhzhfBtzBqJimv8CokCnUR8WWyb+cRDK/cqtwR4NBkXVVzMoD99rwrAYbaN2Yiyb4t
4UfwNkSs8Ve1CCX8Eima1nfBIQnxHwya/OAs23mQG1/NxzyYMKNGkQeLlsY5Ay14os2WO9q+Lhl4
CeBSIA6dagEUc+5hdgJJDorB1OEPA7hmdU9lcPIIV/pVU0yrxC9FrEHGT8UeTFdBjWDcXH9V0dMK
XG9iEPs7A/EtaMahqV3mAfT8r+xfTqayUFtnmTzsodzsiPGhyIm1hPYL7jON44HrAv0YMDUv7fov
nINcBnmx05y/l5WvyhZFaoRVorwyrVuF9ZFAItCn7S8goMvM6ehOnkhQZa/CyIU/mP/bTP+rlFx1
kB3k0EjgU1DxbaezRd63uxDAh/S6z6AvK0OhGbAB5f2K14LXSk/65i5SA4ObjR0zHC6IPFEwN1L0
BiTvi14f0CKJb/6MIWaT3qnfI9WllTf8Poy9R/fNIDB+f9lIdw1oZdkYG0QEOnL5QTkkASRwpySr
33GXsVHnIw1MDc8lbD5w4y/2FvILU2zqtHuSARE1/G2oRVF6DNkr7dpOsh3qAVJkZW3igVfBL6vQ
fWReKU4RQNMJXhArLFmdFLozGqqlv+piRjt2wdbIuip699RaKnwqfITc5p6yqZh42z6XJd69yINn
e4CFue9bJu61pGbydHrim4QkFCyt4+MGbju87wp5JDL9nZPcLrEbnpYe/esxJq02pil7ake/+Is1
35RVpxYnwBWkVFOSQYFJ+UCOFkgTRN/x8usVLEUF3AwGS1R0Tfql295+FOsLb2vvvYCyLPXO8Svi
5R7d5f/3DcoJ+lYAleM48NKLU/YebR5B3oJEU90KGGv/TbEP62aD6F97wndEgzXTfHsD/ZMtPr58
kq8koPiQvXXI0Gd60L2nF3WlqsWLND/ZXmCYkqg/V11AIM0jeOMONxvPEoDqWvm8luJ84bbrwxKf
oTHZx092inHhFvOHiLYt1mLU5qaQQgH+07XHd/ky6joJIYV+HpnFLxMeNFtKcP3wJ63LOXi5D0rq
B2FfSWHI+BnJOlQl+h1JIHfEmdXF0uXkqZIxV7YvXp3tb44kNOZuUq6JidXhyLUWBu5ORfK6P7AR
0PZ66Ozdq+HYWQPwFmrea7KCJfPoU22Z/ZwszMoRTIky4me2rH/kbrGl/AxkR8qnqirUlJ2VVD32
AqxOAEecae7EWNFoWtHQyr2yyQARw5zWDcLVOm5QpoaljsahZjg4GpEQXHwGgDciUU7M9Riuprfa
gH9VLLn6DC0Ak0fl9Z6MMBdbHhvWHg963dHsFSkzMfqL+PHnWn2am9Z/Kx7KJ6uv8bRHowTcunkZ
H5OO4uqxVCNE7s2nQZ14VlhzLiQ74GinKUPQXYvYyf4vsQaqypAjjdUM4mN7xo2UWSRzZq5OiLNq
2lHO6g04m0FIfM00Ssn75Zobe+lCVuhyuLAup/hfLnheeS0J5mlX8kBgDWcLNhk2hsTlim4FvqZs
R50FU/TJZu28cHaykuGCHgOvO7x5SxyocEMDmXqKYgxLSUMYHiX1BAgqvQiUHH1RYd+j8gwCp0oe
ArMxOuJAltBeIhzfSSMS37vd1GIRUw+rHudqAtzmP0AIOsPnPWbcho2/tenOfURn4QcN6/QpiF/b
9RR5OVgU/YBaRQ1yDGJG3qJu3sPRqUCnkjHw9Tke3FNoqkWlX/l2rpY9ukDdoBuaANyFGee9X7dm
BfFSYtFch+4emGWCWFiZA3fzkA6kNE8NLJWeS2p0xpVszFSXlGiGQfYANR3zzRDmZc9UziVs48XC
H8ziMhHkq61sv3QaQXOtO89YAsoH5ZcKM0wPlVNstD4/QVBFKdqRMyIGDP3d4TV0kN6gxMzMhbG0
ya7ktbY6fzurROxD3FpvIcXykW/mfgBSW1sbz3t2qExyuVfw4puyJPj1nTk/ajiluStVfxSP/TQE
OCb1ExwACT7y5DR+f4xE8HC7FF/XbYU3PvnjJ6i2F21wDHXshfcgQdqVfCmMj8fcNCiGTOKUapb1
Qh0faC3Uz32EKsN4VmKzUKkBe6OVI/KGwUMhkOavN9tIeJsJLw2ELLr/JUcDTlK6tRCErOCk2Mg7
KHxEh5unS8CXjw2wecvu+b1WK1adCJ/XYWG0LWPkKMaSVG4MKPuDSYDdB1qjpUyPYX+KxQ9f+jAL
73lnLUHJzpbOELaxBVXIQpSixP0DFimMcArgtPW+h3DLSRiXQS53quo9iqcN4IuFfRWzxcwyyg4l
LagQPnXPzk9tIA/qAMB6nsxLA+uGOLCSgNTnFd346RYdtXvS342AE7hBM63xGsHUlF2N4PzpVOm9
WmEh1xlC7sAzMBO1q0U402ahnewSRax/txdAikat7nN86Jb0TciAtrmDu9/9ZHcPGteWBOFbgy7G
oO3Iy9qtd0toFGuKnkvv6xsnCWQITsReWrtKIs2dOm6YZV5O/4A5BOMEhXI0YDQyH+bwStLqbTOq
BUi57i4qJs/vkMuS/BEwilsvb7EcJWV0gqfu631n0S8J428miKF2ASwM9BL/HMaseLAfr3H+WvrS
CdyszFieww2JxoE65ijedIEwiiUPFCMvYCMOaGdIIouaeM6WQi+7ks2QYsovMgiw9rHmGUG6Vsy/
7AY16rr0TCKOc8ykOtRFKH8XqU+XgdN6Gv9QvLVz0JKIVodLQcYHLu5OXcFe0C25J/vhtSlzjDI1
hdW6Z2vk6MrabWeeoEJniZu2eyEuUnnjtK7q0vcSniw+Pz2jtKfvWIhZSr0FJ1sU4GUM5mJGqHRe
ec3+yoJ8JAT86nHPIpIX/OlrauQKMzOZWwUijGgVvEcD+5mLlYQkht3uf7ScPBTIBltsqKXsHORZ
hiue2e+GH0KUtAACYaVdVJOiNJd2UWCVtCHnUWnGv55GBDusUcdnp+e6POEi96yAHFP6Y6ZuK4DX
rWwiutS5GrwZFdIRdVkrewbb5wzYO6E8/WC7xULS3SlMXX2aOdQvMOfZemN8wLUHFOjLbfGSD+HX
/jDYv0RhxXZc+TPwxCngwj62sozYxI7Gfep2Syh44bxwPQhVykJ8sxJLpH27Juqx31jywAmbfF2b
/aWD0zkydRTeX/y+gRi5ro60NAT9h8mr8QWqpymIeI3vTwZKkfxJrSPdneCv+QitAB6KViV+J9RO
wU++BeJrideZlKRldFWMK9UxrzrZqk/VGWdvm8m0gZh1OIDxTLTKhLToEeMHmovLgzUj8XUWH0vB
sStBsj1DuYn1c9g9xntvuubJMbVeZzct+nvBUPpxOaD4N3jFmwmZmAA7zM9Z+WZXhWwveWirOOTT
07qtvLvX6B+HWNsNHRsviSYWn3D0q/Bhdt0CaynZkTrzTXcHC9ou+eBTuMIelkR8cQ8cAM8LfYZR
TbJF10dp6fdiJ7sk5EgL4ov2izOxzSFSOJlsb8ezA2i18PeNXG1tYTAa6f4ZzsaAtDp8XQ67Wqdx
o7F+lqqlWpZsh0hlz42UxSS5VWFiphTZv8HunHcRFErDNBQgowixlO+fZRIJiTOfv/TdiyfsZzyU
yO/hRbWKVRFjH8g5fZSRf9fsPbCAgr3mj8fkzp0uIa9JIBaHdsogoHImxtGuNr3pDZyamtwUIR1v
YbvZATLNVbgu0riTu4Ewah9tEbwB57rXUxR497HUHYhSe+lvi5d/wvpUZu6ReCuyiexHbBLjzZ1M
qu9RQbZlrgpyIyvdo6PVBnaJ4DqY1HjWNPTt/my9M+1VcXcIo47WOYj7X97iD1oZayzZP3OawtHr
1QDxsy0nMHUBWt0krCMkULGT6P6VzkhkPSG2Ep9KKyAGthHeUqB2MVo4oe2c4Jf3XUG/T9A8QXqm
A1strXpf6sB9SpBEKxuhWZrI5DDAgkTXtH17dGtDlf3+HUCTizUZczdXRjjNM1S4kcphtOr1YKCL
BNxQLMgI7ES4yq92y/KI27WL1gzqE0Z8TEZn4N1mlLJgryTJn9w7zJpGxeeah6ePViqyC70bw6WT
D1gXF3qkr6cIyzKPIGRR69Sb34uF7SJIhYA5gnWmbMOtgJ60ir6qajeMEymSR5ZzGfFxQcBVEcaY
3iZJNKWVIF7kHXufdi7ormcAFx2+uXHzIy2RhMY+MFEz/NQf/xQcS5HsC6V7T48yXf11Zd/T4reZ
jnM7YKi7dfx7K07PXxy/FxebBtMvvh2+Wj0OMDchUpO137ds5XvSIQ86PMMLV6queRuLfJtyFtS7
vXgySnePRjeJWbJIbNZkYSe0szVvZJLdFyw4FZD9RYlBCB7fWqUSTHh5Yu0Eh97AU0QOqIx9y0eU
gfZnp/Qalbzk6IVAG85lvyRp7U6f4By6v0jX7DiHjR1g8v95+hU2raBLg2XiRxD5TYb/3RS7Vgaq
94T0qT1bHp7nfsiLAbKtkWQpIe6XWjFFZEtfjaYdJbk+vy6qh5hVE7OHVRObgkCTGRIvIDBXdqUD
vxsoUkAlvzkf3a22bX6YBMJX6DnF0xVhPBvs9W7xETET/WEVvpMl+MYNTMgQq1yTEP/W8olJNr0U
U3ojWlJLZXsednR6ghUUgoeDy2hPHSVZQkFi9J8/W43fd40S5l0ZhvNmjgoFkRZuyMGKHwBG84lh
cP9S/aQAfNCVxuNJQKBa6MuSx6BmPH6RdAqXg8VD0E6j9v+4NzQwVyUuHsZVTEKpMG1G1b9V6Z4M
D8pYUCsmqxdXGsVtKwgr1FHSvgs9znkU0fyLQIBX1XKaiVrsaaNduiWw+HiCU2FNXc32BTgmG1Hf
5lSRZvW7jAqTMXNM2vIBhVkJFIGp4u8b1sAMomRxWodkv+X/vo6OHRs9MJPi4R/xVirW1PupsbN2
U2L0I4zpLrcW3U0Fc5Vl1o3FRHygoEVcMVyWx0n5xnKt8it8DdGPQkKRbRtARgAi2q0hBk+fHITR
b0iq/VEW6K8LvLZMlTRnG2ClEGaDsvy+5PYQUe6gYxq2FdTX4CDidXq70IoEP5MxDmusEl4B8lyE
tiPVrSNYQDBG+Jcvz8OCisJJBT1nId03qsKDn+W8l6zloosrBtSUWs4YrxoUPOVaFVrHo92IdMjx
Ubtty2sNE1pTDTOpA8ZVRWvPXTwBZwXlNR/tULMHbfQPuOY7XVeoA2exGoaodIAChS2eb9PD4JST
TAG4tCtjpgpo1AzYNPP2fDMMEVM3/T51ho2gXbA6rVXP1kpgBnICArimwGkMcYc=
`protect end_protected
