--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
i00+5BPK/btINOqa5AvjUJRhLmM3GVmGtMoRvkhTO4H25uTcKiJ93XTP7H6zydMimpHXOCZkPqxY
UlN0lTK3rgDYiRPCmE2IZMruPR6FN808fe+m2l7eEoxndfJqA/OPw+4jt0/LAqgbz9YtktpBk39q
x6+XjJKB8tcqFfe+diF+heRbiA1Ufz7vzP4yI3os7Y0s4GfaRCM5V4yMhHecl5IB1FQ8BaIVDDQ0
lBUXdU1iIcPNkVqJNcq9HB2JXux4ZI8sfOHj7M3BxdRn35EkGtrhBuhXMchVNjw/AqYf9F6AfBgy
4MIEIP9766UkpNWHZamh2mbhXsMwdVBHhA3kwA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="ByAFKPDrRfiqdznNhPLDfKO999hjZFJ3FKFitah8FFc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
kuLxwi9iiMLSB3LLBtNYei2Bo5H9hEb123YUYwahSbOm4X0F622caJunYjxinJ1tG+IfJlzv7YVd
aZrEj8wMfnc+wkszEKmYtl+Q5Sd8qtzoMvQ51i1/r4/bbPFuKh6JOr0TNJIPYxFzv3vYwt4lUhju
FDiSLYNPcA7ogn77kYESAta//90i2KcZJU241oKkFgSelDaA6wAQU34ZUDkkLtV5OXL6dvW9frcM
Xyb5YRL3oG9CSL8D3XKeyoNEnAE+FiFiP2bA1DUvO3yxYpn7zRXkNkEIPtMeBVNAAMP6zvkbEoXA
swZbIRB2QwXErx5kgf8LeMHf5h9yIxA/mBbNVQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="++fxT74IdW+u41MwGy/OLMdDSt95GyGgNBJWnppQT7E="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2080)
`protect data_block
d05l8V2w4sqBHRA52GxZmbldd4zSswdLTOnbr4Oj3AzDUR/3kzyweL47co1l/MvKTF/V+/9Vq2h8
Q1L+uqiQGL7aN3m6PwUQVhpuCBpO1bQVANnqbC/eer2JeNaENpbR5j3uCzCaZs98S57j9n8pXpQN
VYzCl0aak0kksp0UCBUSpGF2+c0vvYEfxQGaZ/0Z4W9U8Zo9jGc65K8+gt7gDGkj1Wxs6V/f3aez
lpLMcOGwle75d/2zQGiA+G1/i+Br3PzjHgkAUu3cTSQY2MY3Mj289yuI5/bzH7VVRBdx01bclm25
hRFXDiVlSF4MS/xDenvQvoTmw8+uYSmxm7098UO5rLKB2tK/Uuer476G+Aa47/iNF4tzkV0g9DKa
D464pkEM9azexzwFymYXuInkRKZpbhN+9dgAOG5bEdTB821uVOKC0YChazb3xzo12X3ATDy23eQa
/ru2sxsZC6nQt4FoyrD+JP5D0wijpQU2M5MPTAMjBgekslW729+F6LtsUyUrwxfto756unMtp0rK
klKvzY6pXGeLOLa4o2Uun8fjy93h+auYafRzJqa7vBw5RVbrm/rTzMvtuMPz9ftNFp17219g9YgR
0jsM3t0FzMP1Dm5LiZrq/UAe9f1XT9XeI+BW4krSoneVgtDA7oaX7TlvzVfWbdy9pt1z+LNiPJ1a
ELFCWB4xy32awuDT4+Nqsf7Vuw18S+CpwmRtWYMZ+YypLFWNTIuC+onJU1mQqayoWJNnPtsnCs8o
sOMInXImy7w/znNrJsvm402RaCn+6Mam3HHhctJ4/qPr9WhvFNTvA2ntGeoo6SWCKt3T0PPf7QCR
EetHXjuinyATEwBeXc+gBWFtebgyDucV8SSb9ilXQ8iFuj2mtokjnBw4pAMnDMmLSB4SQjHHtXKS
1lnY9pjVDN9vUhldTy7V1JC6niZYx6SjifmHcSLo5LJRK8z73iGuQ2ZvKUtz1lh0VcvuXOwa4i5Q
X3mYq0lTK4we6n9Np3503TtA1xDmxM//to4lNlVbxPDPFeo7txCTERhFNvKoYv2gkBlAH2fProeM
/jnlfWTkuyt/r865+S9maz5O+TDzJxggI5JCA4erTIWFYzAJOonGtBlo3O2kRwCurd41J0k47ENW
o0Zg1H0t/rP/ttMvQRs2owa1n6TyBc3aAxBeZ93N7Z3+GCwXKc89zXd97MTE84q0YiNJGRq131+z
n0WvIj2I04oPoI57hxHXNcEFg1xQtrFzJygmSDlu39Zc2b7CpwBV8LDql1t7OuDSx/h8FFNY6kW6
H/YwoUxWzv9lPEpBvay6egpnxccCNKUnYHCp6zczbm1/PghTHc4+ZCXMca/WyDjTk96jopX0QOZE
5MZE+AP/b/+hRglDRioYaL2L4qBBBhwhaDEygMrLdm9NXWFaggnrf6EYHL1pm9fO9bUUTMVmbYHL
sx8j2fZ6oTbSrQ76bJWttFpOYty+M0Tx6fnwpJ7u5YhHVXDufCMR7YEshnV9FEcbrXCol5z43lM8
pICcU/y5ipR5ApBffIHylhcqvO16Rz/LSKYEswog+OFtVZKTrxx+zCa9PKKEMpeM/M3UeI85P7Dv
+/DWI96AcOg1WiPflhpJcR/EHHamwGFUtM3EjdBKKPr8lCmxSnK38EiNQdo05FOhZSegzgaLz/oB
GHQZ5tJDtJJ0uMJwKpD9OTYyqpSVa7v07W90LDmiWFUjkOChj2s94oOba1odHS1pjmCCsxaqPFAo
xS413ovIIOS4y4qN0FqDNoQUKEMFrO3V+1ei/0NiVILlcWhaQQGzgczoeGsFaKob5Mrrw8DsXbAH
irLrRcevsM6c3uiJkMJy2fIO4Xg1iNIcRecoZiLGUZBFmsvWXU7XLU/l/YKjWp8ry3vNhqD15TkD
i347m+T3LUWhRR/RsYy+it9c9e5EcUWAhWH+RYdFiFH4QS0oIeDX9Xr5D8D3P/5MjpHBCMEeQKxD
ROEE8V2c3ANP+cUKszJEUINaq6USWaINK8dEuEGOH3jAx/0WziqzHLcudxwf71T9LeDeS/dAGoId
slEvYy1j/lWkhw5i9V/ZGWG1tnOHPCrNbVSluGQ3CaQTjFuuKOQUSDgCRQlpAxWYA7ZKr9B/f247
E4sE88UgAqM05IR0pSf3w8lL3YkXcqkHhGTjB9hR+/kuTaICjEM3/VdjVsPmXxCLwDGQk/stEt5N
z+DUFiuPMhS7rertWBYPs5pPmMZ9eeVE+NYAaGtdtW01wDRXcKZMNBp7qT0JjHhra6MVPJn8WIAo
+mFEePCbjq8VZ4pmDZ9B/EqtiCzUyqgQmW1r/s1k9TywtLwkseEPcwZQknRDLEfzqtoR0LBBJY8O
pHpd7YPPbLJukusdPhT0j75RcI2KGSll/uve1xb8xoBq0Y2d2h9UZWCZYOEnNkhYVBYFnlfNETfo
kLfo8PIryhXPq00g2V1gPyzGaIXgCcnszsB2TYvjzWHr48dGpPab0WAj0uX/rdQFmoCXxfbDoqkG
mfi4M/9yvH86Ykz/RLJBAiuwsPAZVkllgNiXwr2iD4tm7kktFMk3R+AKWolgADtb53tLsVm8Nxgn
svTnrfCfm7bJF3E83H29LAC9sYhx273kyezjt+wPlOyyJ18RRVgM30LhJBB1jAWiC17TThTeziWN
I6+NfsK0luyi1jnaafj187BJn9Mh/Z/c0CVhvoiaCz0z2YeLBJkfoSubOXHPaysz3oyZ6Ii/z5s2
kgNf9ejNcsimGap/orDJOWew++ZgwXNZtsNdiA==
`protect end_protected
