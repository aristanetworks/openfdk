--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
lGRiPYFA9Ej5wcJAHCFuMveKHozgfIFCgKOouOiL6eJTxe6vZBrn0mUMTE5vpElfGsmW9LEyjWH2
CnCk2/oqF/+LBGKKTYFb1wWFi+rfRWlwTqkCtI5KUA7HcFkw2vxEeP7vUnGS8JBQUBFi2qMcfbZA
z3GIZY71vng/JzC1sFNKlNQ9a07g+wDrpKMWRcVU84si6d4B6jyQF5Els9/ufhY9la7JgSlLbPEt
SejkLbHe5g5gs2yrgdVcESaUrRF9OLtYKcYiz+/KorG+CTvNkudVHmTFT6N99ywS12UeX7NID5hN
MpcWSurGhwVuMW37rFLiN3GXfFPuB2BaBKXBzA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="mo3kywjp8yqQuqqNxm3QbTqSNNF9kPHreTZVr0All8M="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
qM31/rDXRY8Zr60lCSKXu5/PNX9nig78wsUyY168xhQ3bA7yX4j7IcDFoPQhjJ7+4yv0CK/GNeiQ
CasauOKb2/a5jzy4LFltRi+vlW9miDmkDSo/65DfgoECJV/e2ZqYg89iHJspV1xx3tZMetGgAw9j
DPBKt0kBoVkvsLWWJ/JwMQn6NcfWZQvonlerzfz2J1wVAygipjYERMCIPVAGBEf4SILE43if4tqk
6s+9QDFN6peW1wWMKkisNoxtcEjjnS7nvMT571Oj9YGUcCvMllRUM5a3GYBJ3lrC2DjsfcTc7saH
ZHwxlykqn9cXmq4c+J+ut4JlVAPwC/RJmBbjrw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Jn1Lb6xTrhvNnD27ZqEc6fu6/hcxjaVxQkoRcP3Mfvs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4208)
`protect data_block
eqeKs+nkhaX8HCq4/HupLGBH8PCzzo+r7LMfVQs/2uJOvFOKa9FcptEH9dfzx5ErwUCMYzrRApzB
71UrL274jDQjcEQ2gyNfmjKRIKYimFDI7UcosgNsUEITPoRy+USIvbYNIQAcnijCzKoyMk5/PCS9
ZAcfkj6jsSfR9morL8chmrdC4wKecOXCr0kwbk7SEjxWAEoPFRmfyss72XuQZdirG3tMChKXX6WC
K39m/4yhUaBtLuZ8AdpDflwEhg9gsUdCgi66j3QvLdeFo72riDzr7gJvaca5pCQNMqtmrwzhuKbh
YH5kiG97sk8QLA86rvoC3u1rVb2LS1fLvtfEvs8A5R0jFgq3lVbeolEfkhZOset+D7STKLlAFX/i
ybdCLxpaHNHkjzMiSRmQmg729SIB5h/jkkIaU14nF5s8xDSEsA3rqePq4XBswMgwY74HDnlsSc/+
HIRwDGlxVO8Dyz47tAgktPeB8lYeSQPmSa9sEcQoPDyeC15KL1vZaumMi6PyCs48DN9SOW1fvBbi
eBBdMFhZUBrKABbepR9o2gsBuVC43cPytGmNOgnn2bcSwG7M2C3hvYW/KJwkn9huMbj5BdVSQbTs
n2p+t50cIZQ9CqOMGQGwiDBplOrAsdgyaDZj9gLbKJTgGU9LDibnzw6s6Rv99c76wmiRnCz11GRx
zwFGEA+sKoe3OqmBsklELe59785ZDO05DSkWhqVg6WkUnlTv6lAl45RUUUMII55hmErXvpfBTjEp
xdVPTQpSQNe9MLRvT4n59imr52NwV5lkFmeTgXk5vaFCeduelBftilDXlH2e+bYtV6oZ5o1+nuEY
h9lwAdcJq+z8/VYYvx3zgNSI4axyKYKJlr3VVQYVPH05DKyzChW2+a/7wM7rNNgyy+4TRDr8w0Nu
Lc7xT76y4x3cPfTxhYwckNrpxv3BiecQvY/eAFxQWGkaCD/mo5rc7ewKkyaX4ZjMry91PskeX4v5
y1WIxx7UHKR2cSkxR8uDqiwuVcH8CbK6XJQkQRItywufKH9iYizJG2prb0kkaI/1lq5xkJcNrDWU
vetVp5nutylRCR0D6Kd0HCiezHKWMHqqKm5zD2+CQ/Ljnigvu8OMU7nWbHmOJkce1NPF0gWCOscQ
kyyae0IL4ZvCYiazMa6uodUI2EJ9HhoLVCG0uMgf1l4vtPppXc0oh5KlKKErHkw2Slr94wR/Ypva
y2BWLdiC7GH62dqE2Dur8mqhy6lysgTMmAGsAQhG3jUX222wQ4inaHhRl+4jS+GbwuCIt/U6n3Qb
Nksia0B5eZPu0XFC5oOW1u0+C2EBcw+7WnskdozIb5ZP9Aae7mnS77Ntykq8tqRZzGK/6ndwVTZB
YCncopUdPUrU01Yv0G8eJPQ0N394s+4SRfnIzoHjbM2EKmnnNbdz1otyOtfosHEPiK3yaLGeI057
0TZohuoKKzRGPxgd5Sf4SsAomx4Q5CEk2jEQmydU2NhHyux1GRCsLFyVRKcn6AEmQA116Y4/TX7L
pm5Dm1LiQvYYk2pJmGIcxpLPfeAfiVhglsOeINUqBugKSeXTRiaUxO5352YJqJ71Xj/UsibWABU7
S7ikbE62HWwN5o83kRBZpuqT4dtCF0wzX8tgZptverV7VFa4UlOVE4bjUedHclXsnS1mZdBXz+qY
DitPbKd5YkfgKHFS2JsibbCOsw6yDWgS5e5UN/+XnFF4hhLGxgzB/cDvFBVCLo/WfSAvTwUDdXib
K1Fsdj4+mUDLqMSFgB0nHnfS1gETrUFyO75yJJfZUq623wSN4utUnvAk+EqXVbhSzF1WvGc8QuOa
sWBQxgBEC1rA+GqosNbjZ4/5BF6jPNXLxLiW8fiKSy3/gMpF9FFi3gF6FhCxV8b5WLt65ECvsAQI
Br8cXn5+tv7LnFGMfWK67MOG7mgkG6DzAKngODBcWOzrBy42zqoJhK2WIb20VO/iuu5faID9ahfg
97EzAK7cMXCT5LnCIc66Z9O2rePZa2BuMd82tGOOGWTziIpTPNbTBbUdfo01IEkR0vB189p/6Gc9
Xqy5J+tVWHEk347+aszFuOHXyeycTSzUu4n6xOcfgONZnWRXG7Or4KOLUQsMW8MLDFbu3OdrhEU3
29+MocOQET8vCpjfjYggJE4cCUWCRXDSyDRAgmnFdz+Ev1Km9QH0L6FUrilYPCqFMlVcs1ntgPyT
n4UfolwtXePGvmtYgXZSxrTPwURSYR5XI02kRRKKWUgSoFMj7jYqCoCFAMQLrA1t857cBP4xzP1g
j5xmMNTydWXr00m8Q7wNvgbQL5rnx2JRvU4XgjU+2xF9mITURuKp3IjOUS4HRSHLyMsejI506Z84
AQCLrI4Bz95qJ1NbpIrX9GkJIVcun3L65LBIm6jqx52oxkJnbQfg0xpnOiD3V4iSfArmxvcVjxAT
fe4yLtcb2r5LRnyqT7qghR1iO5Q3lypMSNlxMkB8jatDWaZMIlVqKjay3sgTkUExSx+TadPsYQ7+
NRcKv9k2LiFgackqZPlTRo/Isus9tM7O8kS2FxX6g/cB2hFbtHFEdXSdqCa2CfAqusrnpFzgHOq5
LkkOqrwsdBCBK8TJGGHuRGL7vonf8GqQYgtoeiJVYAi9plAL/5x588rQkvfcZTlvpcMlTeHRJFxt
CTOINuX+C+1WEvZVB16cLCBAzGLhKS0eApVtljr50FyTwEAzXxPT9+JDFaZd8Qre/10xobR5Sx2y
R+jgu6wekJWc0NFW0pmATTsBJIW4LeXn5LTSuJdEInooWTm2pxImVm3Zf6XRjQs+qf2x2h+TAeWx
PTsnfqdovNy7D6LE6TNimHrPMPF+BcO8pGeW7lcPYwnbo1u9drZ7Tky24AAQAhn3w3zUn635zT1a
UvUtMunePuM1CQn4+5HLDdGh9kzvhILqDjS0zSJ0uxLJywaDeCMInMsF0U3ug3t5+wqSIsn9lYqU
V47MWiji/zENS7F4dibLKmGs8Kn8e1MoppEcAWe8ISV60AsmOTImGwbFkdQjuTd8Yqz/BjzSkYWU
1bXjOUJKmuIUeVwqc62TPCzdsd/P3ioEc9ITj0kmoG2BuFJ93nBOgPUc6Afu1C7JPxXRABPBJWpD
HLOfZqCfp0nAdonwpmm9Ek0kQCzxoH024USzR01GfMpXOiVSH7XYTOzRqkLTZTz9UGsw9+QUWUp5
flTY4ymcgqjtFxQB36yokqaCzJATZuKHWFs3bZ5q4z3X0XHnxoqRHURERWlDYIZ78MDg5FKdxfOe
lvlNaUchOgLfckyQuGKC8+rxN+seQ8GBB4e4rkeP809EImBuil2hRpNIjQ46RPygRtozoG9potUm
gWHDbS70Iym87xSn0h4JY8I41Qx22dFHvbY42mpW0zNVLhfpwF/Q+UO1F4rqSrXM74ELeX5+wPBB
shRw4akAiBOb64YJGA/Y79DysEsS/bw8ujPwVfHK4PDNoM1WHNGx6wvIDjmUAvWFj59ClPkIpiKE
WyBkAtyxhWWVi5GNgB2XK9ecDUTupLj8MxM8KHN2EVs3P6RRm7EyvNT6gDLZ7L4dfxqO8HNdmedr
rVJ3PaqHsqSMUuIVa7E+KQzD+S85Cku+3imi5jzlXHwIk6FYGOO39a1MzP9e4gLn6PgNfamy3ClJ
74IhJAaVVFF6uoe9KVGA5dM1dg1W9PmeKJ7dZucI4R+CJ8ane7sgfyW6qGKVmvZrqe8Cp1P/fMT+
QcA5CIuz2y4PEG7xB8ABG2szsiWu7lmwTwdr82rPuXO8tB32cqcdFbCvEQSTQngrY19owRLSzhua
qf5sFPLeBriYw9CQTlNJ6CP2fYz8D9v25fA7BabtqjxkdwFsJhQfiS6T1h5u72os1fFYj1L3F1un
YsaDgWXtvOPgIjCJ7GPL1b1ly1u2JDFaK57d4Dcx+7xR1POnYb8eQ51Quc9iFKurwhpNEDIl/8Rn
Wn76acYLeLaVDHiasvmeW7Xu7gkykF2vGIDaDv+dImWqDAY12kzZHO7fnXtzIdYEtXxNzoGwG9YJ
WFjafFJ2cAoNyBtliqGkdHMe+GVnI6AiI3D+SfuPU3qGZa7dFo/FNt96apsSWd7Q1UniNUS/m9cj
nFtoC7M0Oz9yBuula8ZW9dMZ7bblw1HzcOfyiVKnkt9ItWyyVNagq/XByze2ZrH3ITxIltpgpoiW
79uQ8W/idTYOMskxB8EhtDyBYO9R8Jc6MI0xX2GoQK6XwUT99cexv1czOVtPkdpmwIXx5efnnOjL
SYaYgMQJONSFcfDhyvtoF3FfKacvyibb180lDX30wgciUbcWOj7SD3tkvZKtEPLzkSdS8/X0Q1SM
Wgh0LviuWCW5WKdO1dK637yAadoMA/usJdxmj0YO+ujWTqHs5DBdWKOsEL0U/814oM0W4GFb1uJZ
TC8A3CImsvZFyuegRAWr173UvVPkSLx21D0AQY2KDOJ4zE2QsMWbfSLvtj4ZskMnb+flM3EhPW0A
uL1srNY5iJa3qNNLiVbjZW8H9BIsVKKJ1xY/UjAiA0JqrsoVIZ/sCavBhICPKUPZx9ne7AKrt0nN
qsO3UEvSwZ+U8/YqZ1DiBvt8SYA0wiSkb+a2oG6cI2AhaghhcgUrATPiSu38xqwc3faIePtka55O
qkzwhUmFf6sJEuKiO/RyeUFhMjmhKITgySxordqVdw5AfNafw5a2pxqd7bOMkM2aYPhr1Hp6cZTy
IgJhIVyxUFOohuDnTz6KKKiyO+mQCENAEtGVti/7i4E637Ob+GY2B7150a+9lEDOF1pxjxt6LKdK
vU5RtzCRit5pEPj5Flh565PYZ/dno/YFMFrWBnXCeA6Lx8gAiVHT2OT6ACZCO5j4pO8FMeiGUWDJ
95zyqlplTXNBTtMfxasbkVVnI+DRKs/+ZE/HlfK3Ow0eXtRDzf07XWnw1rrOIQvhOre3AeRtFOol
JATbfZpBBRdTY8xsZuczGQe3TPZ2QWz4QzWdecelwlwoKf/heykXWqwisrkIs1nlivqLyjwlBkyC
p5w3qdeFolaKvYclYQ+zL6xZ3vgrhOlPnDXaCQ9nnYYvwdzpS/+qHHEFc2Ww9OvsLUF+PWIegGff
R64lWkUCkwTc7qfQvyG/hY33RcdZTR83UYL2TkXRVo0ULYw758mQ1UpiWJjDJVQIk5xrVkb9bTG7
G/MwnRwNjsIFcT59Zrxj4VpMHmiBlcyWJxUOTABJHWw24nLTWzGY56XKTqS6f5rBKxDiFp53oUNm
ZRyCAFWSF7BXF8hcoFQPvLuBVNcv5hJrSUm3Ra0R4hR9uynVYIUKMzUvUPMFOaULqYGoDZElbsH2
17ftF+U5sQUnYSLtrsn08nc0eBiBEP+96TPt2xxNA+HW4C9EEO9QHG3e0CXLI1aNpmCFiLE3Yg8n
ZwSl3hAlJ2FJXKn3QDaNc/gucaEgogQ/D7rBz2GAA98+ueBDSU4qOYbwakrt9Iwzs4/7O3ZZUUhS
RXBH4XGy560VrzqYsMUTf8nyLxMjEa9k7YARMdOLqP4f0aYL81wIArFvON7Vlrypl6nJy28RWp/I
KkVysHCFCqgoRuidEP9ln3W4Uzg8TCIRK+iDSajMepMKs/DkHXD7nJkqcKtvSrk=
`protect end_protected
