--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
R4M7PaGE6kJDVbokS40T0kOVtNN4Xc64ocoOVu9ONZ6V0JdJB/BNQ9F7aeMHJBIUb2ROaSG8tzRZ
0aYf4tBYgCVnLNSsB+KH688i70y57rt8waLzWJjqKbVjWOLrJNeVwIazyyQY0nQ0DioaEbi8OT27
dcW882rDIM5ciMjyGR4b9d9LDuFqF6bdNAC1Ms/qAHL5OSh9HEjsP9nGnivlDoRwkkS+IYPuD0CB
xvbn3IlaCg/mSnBuaOcnx06GWDsm0LwuLIiRDIOG+Orff2k/VbpYD5GfeG4y2cjA12Ftjt5ulYyV
+r0K+rODcS2yhg9NK9Uvz+fxxtfuFfCXlmRi8Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="HEKLgg8SfnYKs3t4qOAP+HNosNoEj9217LcdKI2OuvM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
avLZ7mqWTprnwa/VGmfQozrCmWlBQQVvw8l1s2E7GfrgvfiLOQWkhU12PUlQqB9b/VfnN2jiLM8l
0Qax51EdWZ8WpSoSlfvwBDA5Ey0T4VMqlhfrgOdRsXs8WZ5aGz3H1irsjBbSD/puSd6wBY511osI
G27YuXbVuuUQ2e7xAlUmda396NqfTMJwplc3E+j2Uan2Bt1ySu7cRZ8Vhs140J3TWgrY9Xed3sIm
8nRmBBn9svw2TKFuT/QhqFcUA8h/GBG7W3sdlTgki6KGX4euybudPodLxwhkUy+NdcypmVRWtdyY
G3IubI/FRraKG8aXLzuyzYL9qxfVC9WHz3dhvw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="km430Is/Clnp37bvSlOxSXhfgfi9pqgsH/+1Z+Ppd64="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9440)
`protect data_block
utcP7wiD4tyRtIc7nmkn91iB0n4yfDJZJktXnEWILOcbFoBowKQ8KgT9qvNMieYhBExiokBj8Ima
DvIOnU52zHm9VmJWQLeQ3Epz2+ag0d1fS4V3kSTtAX059hfWBcMkYDQj6NjK0KGlCQKaSKZ+q6iB
rZYAcloGKZKEZNesB5qg+0gG6LatICAiZmmkp61KDWuNPFzAPqaEnZRlUGyq5gw3QdhsB7o79JhY
qltQsMJE82oi2theR869db5WPTuezQpUZaHLron9dNMQjQKyh6euogYrkpcbc1SU3xgUQKqHz/iB
VKwVmEDL167RHYamqUMVyxWRqt+3ppklKM4Gmymu3ZRDuunSpuTdSXTFLt41JfuHgkn9IE/zQlZI
BTz3qKyLvnbKxymKiX5CGKV+uB2dZwAZuPC/nXtQJZWAgCh8W0xMrxiUjIsCx1jY4b4OnoQ1x6tu
YjidddNgVz+ErU2Fp1h4GeVl25o9kscloduMDb9Q4JTK2/LpGAlrN569ckgXBue1SqG4yIe2xvXt
cC/q8ascfHeCkrTVQLvYiQO0byEDEgUZtW5agwPvqONYaPF9Torkki9R0UbTI2t3lhWvjOvOqO11
MVsq62cNeJLcKFggTXLzO9tB6O6ThxewNMh9bM8a0U4Et7ShUl8Zqsv7FlEqXIXnzJnBIJQ1RGZm
Puvlmyxo+WlrTOT/V5gNnnQyEpGXyn3NPVFvOMNRoStJCtT85ZlULtrEINHBLwGnbPdbhCJ7LXHi
J0cfbbYb8gEenlo99JwGTF1M1y9kP4kB5uhMNqFfRIJ0rlVRBEkCn1LOUd8dSWieXPPwUlHZWNvU
soaltnUwpS9gaVPw4p8ZDKVXQ9YKDV0K7J5GRUFKoFt7+tL1nrY9m5Lb7X2tj+zQ4JZ7MdjEel/P
vjPuEi0zJ9petpFzMeVRBoh1pWdospcBLFal6MQt2xKNvUTiBYTpXGgFxh7eLetjPvIK0afbHFoC
M6Z44/n6Lu3afYE6CRKQjtS2dNcpkbEHwtydXovSmN9vqKXk/b1R9kp7RVgFrrErFGHuL4xJQs4y
DuIlkGLN+WJ6rh7/gyqFa29GRw2fxawJ40usrxf0A8obNJec7Ajf7vBa9L4uPyrmPTYUinMcMEur
8mxU/N4Vc1nKHrwPXUO2W+++bygjSH/LxDY+MlhaD7y9tWzafeLLJ2dGEkMTcza3+mRfbxMdnuoP
h31rMgwPLwdlU5OF7ZHnb71nTrSUZKAzX/OhEHr8nJUgFGWHctXZ0W5wXyy0sHRKZfbgvSmSZWJw
yffnncOCOggbyNM5tOh203o1Fz2QrIDGPwavXfO6aTGLU/EVZHSm+a26J0aDfhihHW+vAMEMN8nB
8PHmTqVkWvbhQrcXdgwYQ8ShtbKzbMMrf8AwCABKznAT7RGme5YKgGYY98SbpMCZdEbYOIPcwjFd
EMOp2kE3ZR34kjTZoTcuiCNtIH64U9J6Zb+nM4zyHK5VNJ7IlBYRveDr1f4nROX8zzD0vt5kzFZj
w23BhSYy/i/bRQ7cOKO+vCqkD1KPDfh7BQEV6nyp88KV4R7eX3rjHol7ZmAVnHai2yHjy0NGpLgp
U1txgWCyWS4WHjzjl4LN10HM3y1yDlx9v2xO/zdo/wyJaSTHAzJ6W1LxJPoHsxsnI/c8aVcEGVQ1
1CQIjVTXZ4om9rwSLi9M6kkbDAZt1YtKHD1tNrVtDBQM8Lp8Ngl+2/kKOSZCyDmUXpR8mTwkRZSs
7OHmxLTmisoJP0d/vKd9eTYASTsUNZxEmxLlVG0NGmvbU7x7FMYUgNqCQMVIuZ1M3bBpntm2QTUG
x4fj016nyxq8onSDcjWseV+IULAQbgQpJ/Rm3kqfB7Fm9R7UBxw9T2GEFeRK/wrRBn+rfkYh879N
hWnbkGFXwLzhh6rv58/BRs+5fpA1Cq+HefqvAF9oJ4hKNWAizPnYgbBHyTE2kv2F9vmR0jzzjCi6
HjjnSKWPdWkfpnb9v+gkPFT4/AJRR1lrtMZX16lZjAgQhrpXgirkfyhnh439XkXAgqSuVpxsAVKF
+NJdlCkcYCB4CYcqyPNIurThZwqAT7Fl2z97ccvwlRTReU4xhNubnCCnYvAA5TMVzZynGECh8TDY
8KwW851flPXfSJoxkNZYgGoiVb0SDT9umje8E7PXdI/gXrtqs8DbNh/E4rNy6qArdF3RIPC58B67
zIcr6ddDwyw9YfXbq7S0hZdN/9sTseaId8ORmocUGxL/aw7QESlniIEDUyfQSuKQgGAcJKKCDDeM
MEilAjplGDwpL/9tU6ziZ3yPj0BmFByow+tIB499sSWyGK6kK+0AHSx3fT0CMjq3fjuD3SxS8Lbo
UbLV50SIkxmf2AP+n3Dl4P4Kn0zKZIqzXLnP0DWSKr/Ng9L3HHas5YF21cslvefoSJnky07+buus
gC0Ngz2LQmdUEz+ni21L0LW/hYYNTHOncwXTf37mSRLLRMKvTAPUyUAzj47qE5LcfmXwI97oEZZa
yCKb4/v2g4x/imZT+j6/LIemMjZtNxgHcjv7ILGi8MBkG8J7td5eI6oqq7KnIUQqnrkk7a0dm43v
e6qg8rnQ2wx2dAZzZKIhHJkwg1+oClc5bZN2S4bGuJz7/ycMRgc7aOUe7+xN7pzIvaPjdv3rf5JF
LZOoa1ZFosrzwD/Tuewcid4/NOiLEyCaqIeTiQhi3uWXPjEiwaRMh6GqFyzkdQJB7onrYfANLBmz
QDHGR2Mg0Mnnv3ywI058DzNvAQnP4t5l97/LDuw9vRGY1YjV/ChXGHMxtTMJkrERJtA1K09hQ1ex
p5JBusBNCQUWSL3xKKp/ipPJfWRBMXfwdHhpJub1pshd+qv2oehzvLtHqRfxfGT0lYTC4FOtU7td
p1HA5Okh+BLsv90COk0NlUrkBIMmSih7/JOvr2oH/+TY1ydeCFtsY7EiHzv+u2JPzcLyq2juZzDX
XSzFWcz0xKkJJc2ndqGGnFxG0/W860hfGntmqp6XD4VC+KOyOVE5fLL3Ev57oICKx4FivZi64oAm
LLjUGcIOe91uIrphBQHQxG6tAbKehqOpFQVcNUWk06b3lYbXBaimkUitjJbfPfSAZzR/WaThiRhG
SDKvoMi+zg47kGka3hUoQo0ogTGlowFYMol96D74oYcLcaC9a9PFEUok36gMuTEIbTZ4BA10Vg7M
1deQbKOsIMh7EQBGEW+/llRk0kuN2kPf7/uFccZVJNU2y5qvsbAFHODSDmHuqHkI7bkX/JrsVcNP
KigEj+fhgrMgZhJ9Jjuw11R533Ak0Fb3qbV7u2feytCC2noEDzSF5hNbA5N+dkFgJUYEjyxym03a
/nph2XuZ6eQ0EVOp1+nIynipZnlxeCBhoWEbGV5JrTZc2rmpNbTdHcWSBgdt/h2t9F015T1acYxs
XA42xLQJRxZoGMoRZtIPp3aIBnZDtG1zEV7ijRtVSfu8VBkFz6xDdGkc/OjClUookkEhC5kXsoDg
nD1X8wN7wugcskta3uJ9ZzbxFG5EY7YMOPHB63vIKOJoU34HUZxXTM3kFPVMP99IUDxfdMO6ebsh
anVYN7fOod5TW/vdlpw6CNkM0dewshvFYVz7nUIEwSnZVFkqEMs/tgPmO5ge9pDYg7knSnn7yyhd
COWXS3Y4/xt7dVgArciEXhxP69HUaRMy9jgmSKfDwqFH+q07R1+i2H5Gehpo4BcYSwC7S0eHQjUT
6MRjUZsvPwAg11cn1O6e4Bgef40kkDbW39D2k9WZnqH7lAU1jh7uZJGvCXS7qFS+oPVXanoAeeyx
ytuPq1cSSnxTveeqO/Y+069foalwwhi0jONQ3lnE2fon7T3Tp/+8Zx3fo8WY6aCNlasINrNHRhtK
+POz+PyX3DRYIHoJr5Em+xRtQLehKJ7+N3lAaA9SUoN+4Xr/5ldMuD2stAQcn8IlACiHq0DC0uBr
ZtPsbOUEZU2tURfGpONkWpWQ5Ol8mc46O8MKGJeu0Wn87nsP9rzwlQZsgPdoh1L5gtj8TU4mNoQF
i0hq8uhhAExbazVvjCJJulqCHBSRhx9A2/S03jUgA27DyGEN6Q6olbTtQJ24o/HscESnfkV9VXrg
WpjsDds+9Y2eTbMZyROOZ6kF1q1P6xDqSuK9ZzOyfHQYbGhtvgKjB1WJCWkXhfu6AawyMPTO3xD2
Ca49SzF7X0/0G2hWQUBZiX8unNYJt3iDU8bYAZIuXhe3mZwohGY3xEmFTQ+41N8IQptx4oWVKngM
FQ5TcD9Mf45hz3oQFuMqRX2AqCMzs5RDthkmVYQsEICudDS6qEpyc0bnhsZEOEUEeG7oQlt6MwvO
9PzDeKOYZDPVM75sqrWmKH2Cbn1Uox88UpSUMtkdjFW8DbqLGL/ZTqGf1JDOXI0p8I9o/DRPlqzW
GVn5BDjfnv2ev2mQGm5GvhaZcg0A/NeFb88jhuXdXNQ63x+HWee9Xf+2qGsvLf9d4484labA+GsX
afoB57KP8VTISUHco3OaHDKN4bRF54XZQSJFweJS83IfNgP/Am9FYaPC+PI/D6naNA9nYmMg1bhS
9cmFNj3529kgv0pp1eR59YYihO/lGsgAnILiQCGN0hL6tdKYwckQ4hDBVctwCFXpv2i6MGM1ap/n
chqht779rFx06YhbQQ2D9o+ZoTgVrCsRpWd0BcQRPVixoPdrK5yvnCXY/RCJLeu/8R7gDskj8LVJ
R3bt2J4D/ILeeGkDsPfh8tw3f5AR4t8Bu3jxwGKf7GNQ+aOkDowiKJk+ownWhOX7HP2iyQw2Jgoi
8LIblwJuUwPZUCzvSUI3r2hswKc0C5X6DRJ+2MAU1oMJwlOW+MHutpqpqf5tXOKnISY3/VavCoS4
eySWmVfvwk2X+vJ2glKNVqpPpPCofyjeqKf6nzOew+Ux3p0/b4sMqD/J/Aijc7G1XZl8P+1AOvVr
5Q924gcUjRqusNozYBCL7FUH2QQugpbamgcEX0+Zp7J2qh2fe10sA95TROZOXmgA+FTgFLd5xX5l
YJ262nC3jZtcc0E/HOkWYYHs0OpbQuNbeFCsb5JfyGic3XFEtjr+n+hyOIgxsOp64H72mxfvSNN4
46NBYB8OkrX6SOFzFJshBowOvlrN6fe+U677xbXAhD4Iy270E7j9PojSLfhE//xm1dBWslUoYLik
polsr+BR/fHslvDafcMLE004VEKVNq3BWBlDvZPyhsgiMmthK3MXOldhAmgpYvbNUTNNW/78dLuz
mXdyQieEuSMvCXEpUYOeseWnumr62F9MFlxN6PVG2A1KaKULYf2r04Yz/IO8UqfAifdF0a+FJcw1
jA077TgG9x/CwkQ9l8ejcSnL6k5lQzaZswzMnC1UquKNlp4/0AoTr8e2nv120wQjEfJaVOZPE+Vc
kOta6OuaXVPmfn7ZXK4scgbPz0dhKQyVLPjMtSh+iwzfzE4HtTLlb+qIrjkXhEwusMXyRZa9QQ+d
wZfPV908v4XMQywdLh0Jw2W4cpkHKM0tcnECinSNNVM9L4IGSAM+zuYRofFT8LrmGBPTmJcQR9Z7
r4elIbJ6sRRmO+VXDkQfeSlf72H1c74BbV/lOofZqDfSLE5DFNebNypZrnbop4uyEy15tg1fKAO8
Ju5kDt3EpdQGV5WMSlmM1g8nIzHhK1w635GRkFR02JqFygqySJdIRbcOFokm5anihPxsG9aMmODA
m6bz5N1xGyJa0ekDdNy0QHiOCCT9kD1vlSQalP1PzbGiNXq/cH/Obn954mHPGSmpG2AKpvusPUum
rmbL65EMZJmYV4w5YJ1QCFhZBYVSwb01HczLaAyK5WKe9LCugQZP85vA+72V0gcXiUSGz+IPkWfR
YY8avsDEC2uWN1TSy2K+nzATdSY9I8UCEmC9bNo2pgyuULCiLN2XU2SfEhg7uWxcIUgTov202T1I
JtGbS1k18W+BFSLkbIK4RAVgwFG08qrgqsGzk0/9l0MhuhYvfCM/2vVGQ9MK7GX1Yf8o5G+YpLql
K4DRu536kUE4xjDsQHz6hB+ZeI9ymzQ1W3pGMmKeM+S8uG2ZtBiLA+9FeZWiaWYdX+3M56dWX8VD
gq1xw6ymTw3Xo6sQ6/yURpoyc8w8eAvx68lGPZ+Tzfby7AzHA0AQ/YNHQskysMOK4cIZVZohZd33
glGoAg2siNHEnQ/W+UDI48JkODBY/fOmnaItUE+K1H+G2RzdTge2sgwkaxw0Qfg7CVd4MzGqTGjG
PIozVq8sjNV0sY4pnz3jQI5RQ4ZKz4zlFvV3FkFNGpKBx8vhsf2lqixG/kL1QJC2AESHDUGWRewX
p0LkvAa9f1P1BUGRW3mYQdVQ9d21TDZjJTGY+o2qb5J6IZegGcB9BHpXblJsuv5ietLmxL8fh6E/
e2pKK1eBYNkFUZLnIWOlLr+GYF/m1IWxNUWpvsE12SBBxIXj//E3owGWDiBP63rkmfJRXTMDl/qV
khZdr385kffhe7wv0NeIp4gbiAP178x2g1ztDuuhFzyHDCJFaPbaQ1aR/Psq5CdBmbcJrLxIELio
GcZElqtPqdPLmCX7QButSAa9MzJf8zjehB6zmQry9jmmC87lB+107MTIXpIe8NrYScsjnpb2Xz7+
NuBH0XHmmfMLQSF+5JGSFoV07LksSDlqjbpIbJLyUEnO7GtVbvICZWcXCw+7r10sGsjskLcFvoxZ
ZcpgWI4M8vzBofafQDX2BUeCRvVWmRPSjBJF/nZZT2ZMX4OBlM7p9EPr87H1GINfAEeIORmeqfVx
lRliBNnsfzh0CmZuwuwdscDfSAuejUdW9ZI8j2cNdIWER36qfPS/xDwtpf14zORQLD2iOuwWEZnt
C1vZfsRA59+DjSaMhoYD33TR2W0esLpHlXpkoIJH5DYaE6SV7JHONUHisdqAOmYGVjz4p/55Vzqu
QaP9hO+QjYRTf20gV2kJK+qqPp0A6zdZZL7Q7YqTTdOc20mhdVfD4oO6AYsIiyN0M4jROmHY1Xc6
xemtuUs6wMfkF6Ovvq+JGxkWJbcopjDiA7+m64FbtLYik9HSmNqtS40T+xyjPIJlC/oJaCcqemkl
Zmi6YtpZCp/mW87O5WbrKhdKVgXgcWRfdMEfYDf1u2EiomufgqKuwmBBjsHhFAiaZMgUzV04DooT
fgULlMcC6jIUZKcw1jQLIYrnSQ7Ne3RMtXqGMxdH1dpr0sE9E3ko01u2rPoZBc1aq3x+KBubovA5
CR8Oq1Mvv1mvk7d02eoprSTPXirAECz5/jwrxpfwHpbW4mImfQGYC1jD2FcR+hKmLlm8aCYrKeTc
1i5yYZL79iDRRe5l6cZVEl6OctIOS5hiMsCHD7M7J5UlYN0UoUnfb0fSnnxvQ0bdmsH89XxvqKyV
4wPdE9/OIE56ibbJ1pmm9HrjalSRwDEfhoX7J4bK4l80Pg5I+/nRXB34snKyoNtrnXV4rY0qWr6y
nmvshjr3E/jP1xe8ovFFWsXpWCeXM2gfTb2MJoV6z8zOl3yOr6359/a2qnryz/NY8BcH6MO8lhVT
518/Khtn9dUgMyUebR678NU4hC9TpDzSlERTmA24WH8DaZ5RXSpqQ4qBoO630+6Vv+wFioJJacih
6LO8fDR6dL6i8je6qGpIlLDpbp7XnPocc2v8WYx5Yf7nFJ+c9RfdR/H1slxRwr/sx0i9g2Ez+AUd
x6t24g962sP2QQxReC8korUh23kX3So3oYF8Gu0whPrkoU3Qy4w4pDXZzz1GRm4xKLLg8bbBD8I2
tYRyjlz0i+CLC4MgFZPOHs3kz4jbRbe0LlDr6InGc5YATKAvhJNhEdr6k4YLCrsACKTkL4UEwpXt
zpAV8ANDkyaeGBPADImvwp6wMnBglh86cIRPMAytqjbRPq5j1Rmk8RHuULLO6EHxZ56MVvgxWot4
7oDk4MfAJJGrM6nBSbApHRKGURObIZgLajcV2VJXCR7HBGzmUBjsGEfrMnqUCL+PB/vQeKXBtrUP
5c6rgJ5PaNLRxofcByQP+K/UQyo5Cp45WFgaw3zU9hYKOmrIEpuBLeVW1umbIaa1/X7I7oONsNy5
qGdZud3+YSxRoe2CHEa6E83ePHgX+CF0lNO1HZvPeI/LPVpXgYksQS4L7QV6kclT+z7TpryQsPXo
KIFUHF9d0yJ21Vg8bZq77Uw5Hl6CYnXr+YxGARf8/wivACwa01S75GS4hcgIpZVB0xl7N5VpNIss
iza1CTOeZqez/KM4b9pdSRoYJKYFEVY06tRXz4qfa4gaxrxC9XLiOGtlhEAoOCcYZSG+2EjVd1vI
+RjZD+7sGx86GmavZrZjSK7NOZmEyg0qwVFczz5l88MeE2h7VRxJnLXEAWpqorfaYHiE0krbrrw6
tiXoQc/TdhwhKmSUQ1fhSAUqyPNxTuzKpHja9u8yg3zfcDLhenu3utzQPrfPdl6m6prPjw9phvOF
vbF/YxPECYEs/o3vsUd6s0ApChpggF5q3rRqwLLmGFTi6c8AuYC1vq6+tsuBPCra2JFZQ5ZxYdaM
g02Vk3Em+9KH9Hkndn8eDmWJMyLqwjfe2ANVhuunvEf0OVL2Qb9VrEUtU2IH/uFSbzatTRLe7KKL
ORMkDEGOg2XP6qIX7TY9+NQXokbxtwJOXNKN+AsKv0LLZ+B5WVh/jSISawiMH1NhlmtF715CJLAG
D1oi3BjFFYn1uVZn2kNndMmp6siPZKGNqHuwuAJSp5x723rq5dRTWL83LKVxaDMwUzBwbVEqY5WB
EjjPM7Njznw7e+K12Syn/H9c0yrBrUH3jlSM4qp3MUnLyXk/q4Fhv5Yz+W9ivtQABaHpLLHmC9Kg
kJ2jL3jHvbW2G5F+Nc/FB2HYLoYdvnDbSJ9qYSuuh8iu6Xs80ivUgsr+D3rhuMNtrZisk7UoDvSL
mCmS6TYOzBI7aHJhiF4UMH7gQUKFiAk1XnaWbjX3penPffX7GUSvJJDq0Mn0s7+FP+2RY+/V/yvP
bQX8mHEGDtQNyQyYtZLjS/smQ5U4EC8uOTfMgJPfssHzuWA58rsHK0aqWG7aP0ydNeuVE3IbEm8r
nnNbgCtb1nJmBC7m+25Dk3OGzNanOH+E388DwIHA1b2Hb6aNHvOrOBrgAQqcxv5D+9B/dkSaPYRM
P48VpsOgzp+iMY1tLHnnHu9qS3I67330DTjyshmH85Z5F+F40+XbDhmHDIzTyjrf0cHXA1EoRfs8
OTKKcGm2xEwxtEj3U+40WWsVr0LeJJWT5Bqn6aFCYWACfzWaYdv0clLX79hHrZCSQ+rRrjWku9WL
gfWxSO8k2kK6Rm4TOYTUCF/QChZD/iCJ16NNScbErOGn9Qj497mTRCcqyIT/Zj1u6jx3NbcunTdb
Eu6/WDBIYtr4VUdFCQqbqPKX2Ri5u9MgMJGpO/oICGx2P0kOr4+RjOHrVvn2lXEW8E5/N2X/SzuJ
4usqdBSX6rNqtzBU7akpeVCnTD4/U290G+VTZcAXKKIjbhvqfiz/chZWCKsc3BsvIRih+Dqt4t2L
Cz/mCHk5wUV90Ll1/V0TEo7CE1k8Qn58f7UIZB5DtE5nMAxVBPMgpngcCWuVQvmvTqFSMe6pxS+Q
NhHKtUf9bZPT1MGBAw0phK+BTKPQ65SrURAI8Pe3R0H+N1IP87JHQ2kXR7/RnEVCz608mubek7Cw
FKAYa3iqdxctj7xoElstYOpi/7obxBiWx5sNoVWBTrvSrBvAT+thgFesy9G6FgNnQUUjC8JIjYS1
9mvVISTaETN+WMV/gvShuB/bxtKn1ntYp2qRbc4VrIARIT7RXFMzI7rigrgeJkms9HLMpWHU0yu6
oxENysiEwqkrJ0gGcAvotLkDFGl5wks1y7fIZx8HX2jHoDTXKvJ649h58dBqgGgu3vfnF9fzMhWC
fwwDcZKz91dC90Ih31MjPu+Kbdj1Ek22ny4GJWc946ozml/7NazTe3kl3y7EVuUm+loiUDljGS95
ThlK9pmDupsMfEfs0+E1+4K++YJDSuUdhp+1bDm8qcSOH/BJ+nUa2vprovHrUZvjCZfprRXx3ZTJ
O5iMf9uoN+IGnXlLd/Rp8hf2dgb/hAf0Xyxzg3nJyOTE9yN+9wBkdXh8Pp6Xu1AdDnmoJf1OMPri
PLY7cBxvvfC7GUqC8eLW2UaphPJphf/Epe/H3FRtDzHOmiSYrziycZQzsRQMXv1I2QSZ9x+qMQxJ
DYxpRIwzhLS462mJtNBorZGAzfMqM1tik3yDG82fF5+G90Xj5Xof8QOxK3xg3bR73M1rAcNKaXt+
Ivm80wFTIkiS6MMCWzasRkgIGamJIQsplRM/7PwftyQi+GJ6OmfIVp2lXo8w4/tQjIb8f/NAQp+8
x5fUaUrZ9SKDsEs4qz+EyC/OyjtAAE13Ox+P4MiV/W1LrBLII6dXPpjUcNDj6jMYNjRZhe3HUZRP
1QZZA2hDhN4/1kHGdjor2j+0e7QKS1HRyiYvGWLqSU+7cxwHKFbl5CJXTbiLAb/e12jgS2P5/D4j
xFrh0sLC5Hef/j/xYOz+Nv+CsRpB72Lp7PZqpZcKhaARijkq8mJ3YIQSH+bWPmwXadmDsqcy31Ps
6TTUp3CwT0p05hEEKfNu7OAAEc73ejCszDQw2IpUFIDpUO77NIhbkoYD0XKXonG0/NHi96pg2uu/
mV6K4qaUhE+fxW8WmGNOlKjmt9O2M5nU2fviLpAo+ps+PtSYrk894HdzwhoIm0LZBNsI7s3r9r5e
Khj5JU/tQA4MvXrt1wIp88curh4uG+APldL6w9vZOjR22mKsa3u0DeFy9mkMxmaho9KVemI5UWLJ
le1y1AqTPUIg0HlvVD8f/6Jgkwiyu/dEcXbxRq6kEliRcYiS763B7DFb6N1+10Fn7Zkn/eZhWor8
MP/+JgImp2C0fak2sbw2YdhDCptwVoRpc6E1uRXVdc4AB0ohX1S9MLcM1R4dDQZ1xfnOTQgqtFov
JXph343zv95wnIZnXfSHEiYnAAjns+IkTFuYuzskWqXT5ghY2EswyLgLLcnSKOS1KAIWV3qUV8nw
Fw+Z9IjwzNNRd3IC8fJBvBz2WG4Pp5YkjZzlt86e1vM4ps60KeMQ4iQ6GTf/3l+jLw9vVx7pZB5G
F6DiYqUNi3j2ijxZCBy9RD3nPJ4HgMerkMp7nbVb2858bfUBgP760rhf1YLkFl49jgDdWlaBRaSq
uAVGTqWP0n7yy3LQQ0WXDcv0JGltqtwy7rFiqpbwCKIO3gh7lwgDAqHeRFBFzpL+1JMxNM5b02tv
sMMPhij70CurwoAebZK2BmU40Mhm8hFlDsxOBLAmAdWoqls3gCTkmX2hfBneVbbhXa9BCopsK7JH
StKD2qguYg/c7PLy/pXwlfW/D6KB7Dma9xWkx7pkwnLByiUyhEvb8dcbc4xFiWlxbIPjpUYsL1+j
qSwcn7xd8P2+hJ2FVqLJuRO6E5pWD0EE7lRJhx2oU7H4PAGvjHntDpfS9CTkd5eOaYeV6rp7LrSw
dBVdqpuhK9w7DDetMq94vLa+cTdOJl09bWKKPTcMtb2CEIx5fp5kDY3SdYTeMjRL6moN0PEGsnBF
UPK7WfrIiemWxv+xrigIJ9i0prpGTvgOBZpdNIu3UHYuXTmTKSmNPRLzRvHTYXwSTZ0ZgskvUxfe
+VLov0BUCucdL0MlhM+H+eXyiV+ywmpQ112XTJ9f2htvTNcmqB+8EM+P2VVxX3Sapw6yCepVxcfU
sjgcg29hGEx0GhPJNM2+Uu3gUGdoruxQQ2xX+QkUkx1Woj3OHviQ846hw5+hDCzAtSDU+WQ0sqWR
bqYjp5P4PA0PoeftDThCGB95kHedJH38rygCnShgDxernZZ2RGdNTjieZd3/+uBkWw0DeI1hOl2I
szvimIBHEIcmHIp5Q1dHfLDoao9mpBbM+OizD8rt6eH1tq1c3kPRWzCGwBb/auCZSRkYYXvBoZIE
Xe7gks70ek8V1gFuimUZA+ldsLftViwaGoMyB3Y1uMHQzKID8SnzL1kafkDIxZtZSVb+h5EHA0vv
UPGsN/VPhA3ljwSilqhNq8Ohi+hRtVO2eMZLnTv+FnDz0Lsy3iznUSc8cC5nO1cIUNCwR5M77C8q
d3EB9QAchHSDu+o2+tKulbCXe1zjAXi9nX1iSUDCO9HbbYVbW9e1csenN3ytUnqSpk++KgTw5NZV
09TZSS0+3DKTVUV+zdI8wjPOK+iqN6ozEVfbiAiidu9+nfHj9DKoWJZRNQJoxaqfFtXezyDn+/3T
QLgOpJ4pdJKamVC+LSXXXwh5Qz0xlkVQFhZpmQpJ9cU7fGefmO00KQ7yvmwBThsfgm4MaBXD00cA
azoibs7iytavdjkRDWyAI6ndahsaOjkmbu+aN4vf0144JuKxnsGRYTZRcYR06hiRJkCXqfNoGMqc
eKYOreaLq9FzvvhXdHdVLLo0ZRgIyGOI90PiAx18tpxbou8r5dL3CLRqXtDwZvoHQr67aQOCRKsb
gNBLj8219unbBa3MCplw1H+NYWqG8AVYzCQkbyZgAEYs2rrbKKbV63VKa57Dw+hAxJKCBVdtcc9c
J07FjkLTocM4B6bMsgKmK8kQ/KwiEvrEB8lT1vRjd0MQq0Q=
`protect end_protected
