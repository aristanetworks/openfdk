--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
RGDFrFZkJkCHJlcRaWRybVBWKY5/IxZN8UUwqCd1U+7HPwYkAA0Gin8a3a54JHWlkL27A1bIxotG
H0Ayi+I9uxUJBnpADZ3JYs87SETSrKUNlZmk82wGDUCNTzKnJdW0TPyaEUeErkBpvFxpUa7oQ++s
+xzwnpPO37tcn8j8NqixJYTmsh0xNnWUNQZS3XzIIyDSyB7zpUOxTg7JIMWX9RyzX4QwQwv7ZNex
MEUyBJak7s+cbysrMF1gCL9PUQyIas/6KL4JZSWIRZDCuA0bQ9pmVe38c7ixvabWK5GuHjZcBFme
9mV2AfMLConEItrYMLm418nS0xa7bY3YEpufTQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="50zIFYxRhZ0B8LjrBMBcjBam93m/Ppfm2Rzw/zSN40M="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
r0KsAptAGanpfYw5e9BTGXtfPm/Qz+abLYbPuOT8L/tBBudfUJ1twLPgsT4qad0pA//NahY1nxZj
WvfWDGC4VSqK6CC0BsuNtyICZVacLHZbYvdC74NTUa743CJPkMPzq1zWlB+WvaoV1P4RqL5+plOc
LINBVVJOWqPVJR2Bh9Bk04+5WLEvTJ/M/cHWXMSZknyNaMc+QVYcFBeBtu4dnTbzMxQvHhXoeTXv
GjXoMa1OfwqVzM/mUKEKiFIggU4jYeOPFoYG82JTSveodS6YnjRMNXp2Ks+AcFsuTmzws8HNwOi3
TrRYxdiNy17dTkfDpK9PWTFk57Y31O9ds1mJ9g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="yxWF5r1hdznJwxAA6+tJMTbmZ7O4nVBXl4gE2H+zqC8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2464)
`protect data_block
BUzpWAB2DhPCKgHFupV+JNELIPYrG8uV7i64n+zXUzysq+hjDL65Lxk011WDUggJZuph+3fsO1b/
DTazfWl6ZNgatEGZ+Kq9qY7Fay9vUAAo/gn+Pdff/wcYXGIPAvJ4EHIP4Gpm4lKr0ga/8HCSCx2e
kQQykv9+yqcZRVHg6RKj057f0yBlIzWiGd14ZfQwL6RSmtCRB8uEzfrlp6nPF6yRGFX5PChRvOYu
NQWk/URwIwbpJjibtbhOYuAG4g88aJtLbwYYfi4QfD91uy/1lb3CO8Sfamjg0PUR4mt7LXcCJEYQ
ieCX40SMyT3sufLlxE59yTz6DoheKH45CqPjVN1uTuvPIWNbZxaVnTtj6+EPRzvDXEy5SphJuSgG
bRSivrLH1Hc/Rihd7sI+5qHC1wLsy0Y9aGyJQNwcgViWDMnbhc6DztEoL9zdeqsobODHd7bS9pcX
pKIxayVZ6agsshPUTQiQt1XU4e+kc4N3j33dkVRtzHIET7ejseQU1pMftJKdxSm7+Zrc07yHvNfP
K9He2GkYsCfMpXpGbHqkN3Ue6iuwbVnAMsxvy0EbPDKFHmDKNMZ2RnkgWCRW+wvHx1dRLHHjU3CW
Sb8E1XyYQJwpixHYLU7aeWJq5zLO6C1kqhBFqGlXLL6FmxrRRHkDvMTQG2CxQd2NlwowNe+6czAl
6xCcHCoa3BZ+Uh2H/f4qZNVT0jClEQr/exSxU7Ilb5ory02m2NBvom2Mfz+rHIwiKhVM8Dcq5gND
9u2SatMlLnU0KlQPHsrOTgTJ10CCWg7p43jCatJ2FlWftQM7M0VKVQ9mRlGhuRwyYu1zicZb5ytl
b+e3lfrAqhgTXxBNEZ2Kj4cc/SCxe/le9kR2vJ2OjIACz3QadUt5DWJyd8KSjOzmDBi90lFBNJwR
UyuhN3fc9CpOr6pTFANUi9jDt5oqzaKyOwQa6a7wwSdZ8zJkXXQFEToYHGXdki0aLJL1Op9HfEXN
joM+ojpP5zzEncmiZSTpIFofXLSHCR8x3wqrUZGhjYqZgzC9TsE255rxWRVfUQXsvr4A4AcdmjIA
L3y438QpzGPqPDeQyh1b4lze+Rt5j3xflrbP7h++4e9A8cXj7wYtRhF4iKig6HxJnXHOql4w4XEa
7Oi2nei/FZxUi7Qxfv7vHJQ/SLCgluxPmt//j6DojN9HV4+luAJiwukJ89q/nQHlz1JVf1kLuKKB
8TXn2q7al9/PylwH/UC0TkQAbzL9TUWKONpVph44kPZyAVF0s9JHKREoeNe2pedem7iPqWat96pb
lFy7ZpIntD+pNnOni8ZHPwhH1Go3Oh8Mlexu4Dqlh2A9SAprQ+VSo28Eo/2aU0K6zPkqDbU1+tMX
vB+npNZ53CSbIBTWGdxlBZFmtBYX27YSJXvSHABFY8P15jY/WNi/USJ7dYJbcy6ipTEjBtjG3h+x
r0F+84fmRN2wfeehXUJP08iouBNMzHIGMe8KBFnKmfE9w9zm3s9MGwjoHlVTjQMmlb5f59CEf/5h
O5j5FM/vwLPnx/auHA+/eo4X2aJxSE+VyMrV4r6Fx4F2glvyFDxkGedpb8Jqk5Q1gBXAs4DDULip
wq0ObrIm5uZvdllamf7q0ri10A7hX2AA8ulbQx0xNE240LFArffLFCLXpVG+KchTK+cCbOzWcUTe
7lEAMsJ2VOL3ea94a4Sj4MN/ZA/0ybn8LIbb/ko2pan15Ho17pR0YF2DD+k/dJBdVG00BDppU5xX
+Eaqb21je6Bi19s9tnehtxrOCpfD4Db7DLFSW6mA+aKx7Q64t0bfoanp+GQKD0Sj6EWnRSQHmXQx
mji5yGdPWrg1QccRhhMIt/VoxGIN6bdF5Pfginv90iH9/Ls0HQnvK/QJoCogRgjDwtXZVngvxIit
Bo0V2YnirOmvlNQeT9eFxz9n44dhXzRfjSVQZR9bILbMiiXiSc88JmeWQS37iY4Pf6b5yOO2iqrf
lrVgNaFXGqTClx+trXH+AjkgrPRA5lmRb4nlcAA+cW2zfiML9h2BK1sh1qQcrrlbYs0Qs22zZuxR
+G7fz4tSmNYEXDUuTPHzwJKaOM23vbjWR9SuPHcb/8JDca74Y6HPIEck2xjg6wHOW8Jale+YRoLK
LKku5P/6+1KAkkfGPtCOoGPjRtTPlWGu08cJvumN3N6AGRrs6KUxPrzbQNZ5n47rWPKkfEuaFtGk
n9c+MFpJl35Yw8ntHz/TRLzzXXbThrq/fPu02+OuWCfhSfryCbiQOiS4NV4kV1C6fg17cOm8uLuV
ezmKez1FdGQ5hQ9g9X3UbL/ICZ4gZKiXXqMhkkA4iNmGwF8Cjy9UkcUxa13iAYCo2QPkioY8I1PT
5M9DHvl7O0vanw1I7RjLFKpnv9H6Zh35LLBo4LAxjk46RZIyWI2YGVUfHoCb1k1jQPJa86NmQfeL
XShouJ260dwxWkBto5hxZMO3ZrhXi+w+OXtv9l3PL3MW/1gFIR1IkxoWt3K0R8wqK+sd7K38bBk0
ozxvxVyYdeOrw8j+mgMyh6Q3Un/jzKpSvrlo+VMDMDbzkR+BlPOqhkcxq/tPIXyPgi48Xqq4rFJg
uv14Mh82Vl40uJ0D0oRNY6g7GOpGzMAzVvoPT66tkHaU3LtVSK5oYSO4oO8+uxEb0W0l+YVkHjmt
vkoC/6ljHf4/4EWOrZQKE3gVKlNb0Itj79xUJA+YABEj0+fCosNIMHa3dXMLtYpask0Zz50DYWY0
Xkt4CJg+DLL3e8SK9ur1ul8WfwA6GtWkIZL9np+5hS3+D2mry1VMqSRCWV7EidMcG6kFC4sAuCvX
UvWvMZTri1y08isXNOct3C3I4yanRjkgWpFB3FeQNkXJ9CIHxzg3kpPdLour+TCLfGzKI/+cMO7Z
whvzdPrjrjBnVTFpWLyD5WBRidlTb+iSqlZDDpZJCk9EWD5EXX0VWy/lp1xAi1sV1OIzXr/RicO9
CWCX1d+YLyQLN7DwlBZvzGUdLi4aWqDI/UoFRW121kV3xE6u0ghWe5V8oDecLhmWYL66WD9V9S90
weIYMkTeZ7VD6oRZq8py2LQUfSt5vqZCTSqK2RRqjdAP7mcC4zpr0dDE5Jsl+W8icZY7wNsIS3CI
Y0SoAwX26DVYzi86eQf7I+uW3OBCYM/l/iwrAXUqIFhmk38hhb9ADurTaAwxq6LubuLA5bR7fFMJ
foBwa5LLiY242razZzKLmZWOIighQflDOTCNsYnbXbhqIZZKf/yHd4scKXYzz78zDdaj+YZ1UC/v
pNeDhJNUmNgY1KT40A==
`protect end_protected
