--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
VhtU4qXhNX8GsoxaeXVkoXGzqCNyEqV3wpdIrs8THdK+bdA5/9bitL+GEVeIbTwlH3m2xeKkIZup
fhLOKsatwgwc2F8QKenxQPmvzgEepdxGEPuw5+o1833EHD+slZMogf3ETtNYFchVcDDM91ALdKfn
OdWyc7aEdW2C5va77GOC5vKDxjcJXQImrOJ7PvTKjbsjzyil/FO2eUw+f0lbMv1qXUeJ+/bEavMY
ih85/Vx/S2xoFeNGozaXslli14tLlf2opz3icc6mv/t25n9r9nyHsC/TiGC/G5WnkXcHr88NcWHO
+YeHr4ji6O9FfurvO8VxBWW4POC+QxL8rIEKlQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Zm7KO6VcV1gLYu1dIWQApbkzrSXXyP+uzrokAleSlas="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
XbKMKkCEPHuGTvX8HsVuEexNplf+HcROS/u3SeBcQCYc32BQeqRMv0Ry9vyLjRKoXNiSDrq2IFHQ
6hCMyIVvBl2W+9Me8Yzx+EswNZUUDNYWwaNFUH/jaljhcPEa3bUGNeG8VH0CTelnGHXVDf/QlKNV
6ndLhjDtGQV5PQTw3dH/aiFxeXSR206UO9aBzx6p5yX6SxyGw5GyrjrxmPG4hbU+Bkdl9wJGsyqH
nqr7C2P4Wxuc5pXc6Kz0g4QdbrBn+A/mLlunxoe3q3GPDyUCkRlJGrDyc3GBiwpe2zOve8hZXSlm
hZxiNzhLu4D7s9zNblfJOWxmQz4Es6IA2MVw4A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="M6BuzCVmmXEP4FX6LjD4d4fZwDaHqy8AWHfwCGz4JYI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4128)
`protect data_block
dO48KXA35bhaEaRywMDtPS76LmWbDFIx6AOTo8HSnuhEwd/amVdJG3aunHOA39cSLFFAQrA9Sr3s
eIE5Y21DFzr+u/xSAneyy8SrmrI+IOlvnMEJTaB7sQtn7AFcf8U434i06GU2NqXgqceag4b4cCNq
XUrqeLzsYWn0bEpB4qJgp58R741VrnOfqe89eakH5hOJ8Ls4wwN4gNdE4ZR52oiqlPNe17l8Inau
GTHXJCagZM6cObS7S0L1MrrAmN3zydWy1V3WQJDw6AaLZX426TETw86GbMlOJNA0rNyu+A3k8oDa
2v+t+A8dFqzvI2eZObdnz1ani887OR5m8qhPXVd4MWPMMns5SUnweCdMBFCixISvyBdp6CkhKAYV
om51NptCRswyiNW2hYuQuU4SZoB8/pV2S4ftT85Rx4epc8IonxLMWT1wpNLQW4nvhhuH8xK6hb3d
u/IZOb6xdLDZ8PIVuaJ3fAYsjXGwn9cWbxZycDWfMI646tU0Mi0xn9DEqRJw0V3qaFRO7m8FakHg
iyLZ4YGJ8Lky55BT1u1FzvgG/JRdw/26uHg+addG4tKO4AbCEmTAGFP44GbbGkd61o/fD40WXNG5
kQVFM1h+elX9bHobFVuihANtmbDmLt9R+kJ7/hID6dpe06usyTBCEx7W1W4siZK3YQNnvNCuP8cb
hoWxFohrlpPz0x12d95Bj+RVCzNEcxKmTnBM7nRY78R34Cz9J7q7f5L6gdd8t/SFpU0cHqZYLXAz
pyDyWnl/Vo3BvMS9ld9xMmJR+SW3MBlCdry0XjBnIt2ZHNpev0r9DFTFozC0506yoIe/x1L9TBDo
Q1fnDAV+H3blizpU6yc460kCIcHGr5LBJVp86gEQWl8c4CmQU2EVyX1l+2zClZ3FsfqTZSjEZlRH
BqQaiASKxrNhcDbSZt4L2enYKndB7VsGXfFSoLy9t8NJOPsJJCr2OWKUbb7kkyEbBh2ZR+fjjA8W
gxC2ij9zOXGk8En6AUXMqlRae533Gi62DKyjcHjf4rrmKVIDcoWv4buKpk7vw3hInMKKCffIRTzU
34iHXkiXOgp80Qhf8i4uVvOd/dpeAf+Ql/bXZ9WE3ADsbALYpjZUuyk6WgBcsoZ9trGj1l4fGh6d
fig8sERTfquPSKFgPa0t2Op3qslPfHMRbWMkuen22hu233mtPiDuAtSZvvxBVAqGxQ+0DNbjDTSV
flB2PhmHXhzXdx/bsUJfSuZ5HiNvpSEWqvIGjgivC4dTIYQXUQI44/xxxzCmUknRxZ/TZ5Bw3o5W
cFRUHvlGGPcmgvdu6sCxL+dYQbClRGQjRCD/c/BfhgNg3WYl56RZVVhcX++I66X3vVwIalfRb49N
+5qXnszkrkDFvrGm1vgoUUbxpWhzs7KJFas+MB/4SzzUWlQvxw6q/k7Ts1eWaNWB3Qfp8agTJhtj
a+4DYesQsZ1UVPOiKKNqZmzY3J2bAzIssAbDlxPO5IijJwKcyWL22C6W723mLJkMnt8BuFCiCgzd
UtT6KwtvDRoWYy4FozNMAJRGeenDc9d3M7XVd1bHRUa1jH+YI6UH76z33vRTTScr9TNFoPH/sqHr
GOUr681nGdjWCRrcDIy8lUYJThxaawrkWzlLrw36K+qbdqr3U2nqLqTQgP2qeYvS9KBqWBNcQwsn
HdtR3h1D6WxG83vT8ibf24ZNEFVerE/n+c3IjwqRhzy52Wmhjncx8KsOW7mDWNof/jli0seWHTxv
j54u/VPKBzzNFt3eik/N8A9R6VW8SXj6EbnosVRZXckcAZ/97GLkbrY14oLWYPw8UNlZKCKHn2w4
i9Nj6DQ01DHBLmoBBjJPAWVhC/wScKmCPC/BEQhJWcc9Tqq05168h3d6plF3qUCcNV7O35OOy6qm
BarTZAyNiphO2Z+7CuczZhOTvqtV+/qCI+PZyckf2AoS/qgRG+E9rniVhcWQ0EiA+9zJ3Tqip3QP
0WS67R42Kcq+c5bmbLXfwts7Sndjc1xlz/Te4WU7Ez4cLRYrzkm7fgCywRQ0j++WMYYPSsdD/neb
/FcJ5+vLREK2i783e2pu/OhkWYVr+mmCX3mzcK2Dlp//D3VSY6HxN2XVBZK1Su9vtHweXk5so8qL
mImW0fnpuidueiLpUKv9wtesaXRm9dicBlx/RwQFjVHl7ADIzuwmO87h7IYPZwXZYeBxLZoQtN6X
n8dDYKyXyrayLUHBye5VnCPCMDvgAfhUkk5fE8Ni6TNoIQSi5UeAQzF16VauUBSKxSR4BTFXc7we
Bzl1KUp+6IMi1f5qtjeVHHAo7E0AWYQsfczGdXuWndegCSdluEtmbRDZ5UjAY8MnYwfA3yfwTY8N
TNlIebNOLCDc91rAfUEwKaabRhM3BsFIVF9GyIkW6CDmcRGJJuwmemJIv7WoVPBNr2Qwl7v2knqc
5ObsivznzOGVRZ3kV9vydqUSknyitZJtA068KyPTv7V7A9scODe9rPL+X6pT97fBbXaOejGZGPrc
BqK9INntYlICaFyjL0uy5TYBisqutP/5dsVZCl11zUBGbr0R0ih0YODdUl5Qq1mLup1I4HrtN5a0
epiqX2okeZdp1mFCKHWbJBkp94HZx5PJOnv5AA62lMXJTD03FbJvCLy7KGuYHkSOUeGop6zLDPil
8MHfEWDnvL2fPvVH7MiuwjlpdEy2mwbqNeIoNtmXNU7g4VrtrrL7zmY2xt3EyEn/P0bKQxLAls6h
+NhYWaLonsCWzr2YLnIiNnO+qSf/Ik8KayvhxewllZTyAkhm2AGfZr/V9JQYDln5PWno9oWFWGeG
cJmvpcDDeyiivYwGLOicgtYK9m15gV3kipBJAUVhNwQQk74LBTWdGdjky/Oj4LVkLbXQpBKihoj4
iahA8iqk74D1Z6sdStyBhHfrAeItk3Vx5i4safD+gi3Xeonssi4CTHz4mwcKJKq5j8rHHPe087T8
8U4VBl+DeK97maK7dCSZ79Z6sMgtN1yASJ+XBh9b3M2mhQ3xjSHUG3/ybR2hI5io8V7PatsKYjXw
U/vUrfFquoXFawQyfuFkEL515kj+qKGt7YH0RZC9MqcX+8L3EkiZZBq63HqKCuIMzQTdp50RZDmi
82Npl+OzRmS4b8MCrk1pOyBajyzBlaBHXIYEZFgJh+y6IV6SQgJgYeGeyF6tU1SQK9RiWnVVeKp1
b5MhnIl+2ZfSNYU/wUtO6goyP+15d1BD2g8m+4nCw0oGMBZ/nRhkR2OEVpgks7yqS+quVpnpXtTk
aUdmo/gy5bWq/nfHTJOdlU6EYtcr07xJhcDyi+uWLb85wLhQ4GKILrox0s7mHUkN4q346EmfBb3T
2a9zuUb7P/+SVQTI0tz9QuO9hOcbGSCkCBNrGS9Eyv4aNhF4kU6l2/EheHOe99fAAu28XdkQuHrG
YhFuUhN0E0MgPx2YpzxAN16rfuACu7uolNMntv2J2GQIo9OL96tzAVQgUmk4Ow+ra63gPYTUXqLF
QK/RiYpGaIgBO2eB50aiHvN/nkG6nlAN6t73RfrQTmG9L7B3SYJAhEHBa/fupltb6Ee1sU7KCJch
JT6vqzIzD8GCAwJOgWo5hMT8IcH7pKbbFWBbY7PE/MAYqrMz8uN7igJwpuN++w/bRwd+qQADcfbw
uu6nMXm5f6d5kCpl09k0RCisPKDxlWIoPJkLIxl2azmML0BvqbvgbiEPOt/PY5SV0JMp7TE3JqAT
9ErxNauX8R8d8MQ4IDFtZsJ8EVOQk1bEVPe5zoKbpSpoETrJyUl11vA3jJuhPDVW0ohrdPqHlE+u
WVevYrHVCXii+zDexRt0ccQXmt1gHHQy3gg4n9vcokPqEPbxAS0ciDYQDhMjaKPjvn1pOLI1qHwz
0lTqXErichhZ6+k16cISmZ75lmgeZz+tdZbOhZ8O9lbG42JY0pib2hd+5lFXNJnU12iiY+toViX6
tO2TMzqn9r80WvtUupvIlKZ6Vv3sn7geIyPFaBVHSW9g+JZxd8Vex7bwzin68uYJAuUCWoXr27yz
wT+EiuCOqCn75Xr+Knd2hLTBT1NEDItkfu0MIWj9EQawGT/ZS7EzqMXhymLu6v/nbUcYfNoZYCbX
YhxdvN6PaFlRLH00/MQ6F2tUez+8oYwCWrNCEmVElw6rzKhKOFi2g1qtxU/J/6BktKzkcCEr5u6q
o5fZdnd7HzNs+8iUVnTRgvdi2lXbGoMJDZcxVwJClrSasQbluTfNiTvOzropTQe/8VYzF5OW5HXh
jHR503+8M6kNweZMp8S9HR8v3Z3oKtHNx3wszws3cyzdwqpiba55UVRCJpfGBhSRAh4n6iX/9Er9
Q61d1ICsUmoVpWmVHVsH9goJnHWxyQ8/Uv8l+N5h6/qdOyuYH96VgzrXGIJJFeTAyn1J88Jhm2tC
ipDsxzfJcI8yP+KuPx7e8p4S68FVZoCVepbShhGpzi/68vF2vNRq2QWbqvRFKbQIcA+5aC6zDzdG
NfOBE/EccycO2baW6EYjx3okHSZwImGgFCK2MvEHYaHdhPAQOtVW+RQ0Q+GHxe2VunLGzUXqBvtK
aOuRnUAIEqgL6tiMkXEPFvtmGsb0mg2DWBz6R5xRQSoq5AxHe9c4E67Xq8QYf5kcIIOOL7iQjNwW
1EHuw7pNupk6RdYmAlzgJTXS2Eo1dEB68Pg5Hla3sdKU2OSeaEFHnatBoq6j2NgyeYzCHwy+9EIu
Z2xA6JeQUSPu36Wzb86aT9CTaEUlZbA4ZlDaXji65IK784seDsCI2rTNhRUcjS6xXoiJDaXOMty4
pqTmM8QGEA73jmtCxbphPeYeu1RK6iFfVuW6tVInvutL7qVlejO8N2TvzlusMBIOerOadAo44yXD
sRAPvAwC7kPvnjHQYVCRcTK6RvhQfMI6lomc7A4ELDHO0nHm5FtzYfCEuPrUrF2xOmCqHoTgJnKN
d319lDg4suo6gmHcif98AJT7NOvxzeGZg0CBCYkYpE6fnJvXWWA39A6P0tff6T2CpU8B5YVnR9+s
MZSkJUiwfd9Z1cg/kueBb6dFWV7MrLtwhCA2lbDzCS1gVkz3cYyC7Ykmp+LACuqMioF1xkVXq7hv
TLGghg27ZlVXVvSKWbl9XCziDKIta2kynUxvPJoKafBG7xnNTS8yY5mZYcu7uMbNFsdHu+s+D+Tl
zd0N1Ww62uNS9MsrSS2fJ2utBe0HOMrKCfCF0UPSC74YG30pnQhErA2DZXaPjcuzcVbiP1RTY1gD
H3ES2EkUC4cI9nO//NtmKNwUanf1DFczAWLNCBNQabGr+cHsPqluL4a9O1CORlYHTwQzA+eIkyb3
lFdug77p8j9huyDktb9Zy/3brTk1fBE5D3e8CRXx3SZe6IZBi1zt6x0CXmpHmXJuYmr8EyOyV5y2
mD73GPpCDpkLaDfMWorK2iP/KxpZPpqKHM1T0u91vfdXGmNd8/h1p6THHoG6/2TvX9ZCIQEmla5u
mTwvThADk644KwFDhFVV8Em0ysP2tZD/
`protect end_protected
