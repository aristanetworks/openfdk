--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
gGP8wcCFPyJj7aXICLMfxproQiuFY9DY267gCp3wSMclyjaJeXXZchgc6gUxD7mjHW7ERU4uIHM7
/lbLdg/E1xEvil2qKFt4KOHGb8Yzi+Tb/G9fEDkRduPt5qS8ZMc6Nkn79PX7JuzYdDjTeGd+to9x
vyNcEf4QxHvgru08G3f2n1ITYu7OhmP8jdYalLPeqoa2ZG6FUUYWfkV3ZcxQNgtoNohhojLX6Pli
CmEVVEBT3AdcVfObpieEe0XS6Ofs/QhylU1/yDuV45wMT751buMc5o0kBJlbOU+fPBYuNfo8SRDu
VYNXJUcIEV85aAhHXNcHwc/U7QCNEkfGWskNGA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Ii7tIwF4I/n9krTJryhkDho4JAK297v0yz5vdIFNMzw="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
kS22/WTeZ+Abix70EI1ekcQMucZNgFabKnJss2z1DOoCDrVjnfyWzJJXYU+DUWhIERCzhK92DgmI
W+rd2QtUMmLlK62tLrXkz/hZzEyZ2a5z5SNEVyEj11ZIvBtMCCQG3bYkDg6KnCJNNckQQ7c7zH79
YyOZPBmWoq3AM2NR57vTGFRnVQdNIH63WD3S4GFHZKqxhUdPLeX2CYqVrlEr2z2wwcVqd4/zWoC4
rKYcyYsexhUzLM92uWxNW0cOr16NyjGI1dqwglmVVnfXLNJ8338zVEXl54Ip8LYZoSqKqL77386W
CMNYQdWLl8GXcYHoodMWJt3LyUuRTyr56uX6zQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="ePLkeDdiUDIM641K/UCHE61PcGvm6DH7mx6x+s+Jm4A="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6048)
`protect data_block
7anlpmkxqsKqi/H0yQocKbC/k0mcAKkw4dry4fsiY962T+rX/7McUcM3aufd/fq9of3hpyzp9jh/
6JVEG6gTEBQmhFfHrxZy3Og0S9NcZqK1/5cypsUqOZgleMSimppdYdudE0DUzNJ8nVAh3x94R/m7
UB3QIrOfADsAGnpD9+gYj/oDyCjA7nh4oWty6RdCVXhkQNDVqtQjuWD3InCnlcPelB2QwhsX1npi
GbxWA7uvHTDbYs0ZypN6Y0mXU1LH38cHgGLSdWwYNtfNs9wTesPy37J93WBlartjUAO0YveY9+Sk
NxmYSNdMfIEWwevnDETqTub1IWSw2Mb3EiejQi8cDYg9EMHS4IvnodHtHdgknDUZGTyKP93ffNqP
ZiMUi75QBd2LzhI/jBE7dqELpYeo1Xr15KQhePS6zpcEGgM8c5+d60XjerWoRTQ2BIJNQJu2YoHC
fP6sO9f05Z8HtzPWs/28YUsZRV2kBWTtpIm5jnlX+We/JRVF4eKmkyAg1S75NenOml3YgsOboblM
9YqLwuXNKBHXRMCTMQKVEzM3qt/vSwKChSh1Z9h0itYvxjoHb29Y63bFhJrR9UZdgdv5pbrqGAZt
jYpYklgtgzpY829i6+G4vMM3mVGKIx5nQMSHdbnfxpV5vrQ6ZvFv+6ztRCWay+7TUo+89ylO3aon
HR/ibhFEY9HcZ6nQxlqJu0337JSYgwEqCbjZZUUCYju8/yNJeZCCNs3wTg/yehb3qCo1Qc16a3V3
4lJPgxcb2t31EJ1ejxNr9ZZrPKK4wUd59JgIamjSaHAxlPA9a1TiMEyw+m/VsMOj1AehCF8Q4jzc
NsvJ9SGf6UDJkTtnjKLl1qRozDuHYC3EQFnz9+LbJ7Q6Lqvek8eF8RaNwOpkSCyVlzNDb4lI5YHD
ylzq7D9dI9MOcHxTS9gtb0/MJLpklL1byaODgMvJ+UbMlBaRUUx5aDha7Ym2LZerovSPxN0nNDCh
2UAb418XpD7CKWXmai0o95iPsvp86oRfXDz1QWogBfVxSWmpnsCQY9SZYU2LfENrUEVjOMlW2IGy
vqDaxvqqq1k4fUSW87Il3kf0m8XWTHeDCXseAuADoYsu2tFiz+Y7/YutkQY107mH5ji4FqldyHxn
jsjnma47rj7L5sCvdkbYVtd8NNvyoALSg75jOn/fWtLKdYvkoIqHo0iTVIGcDBn4WTrTECbYy0FE
JQDGoxKi68Dmi+IQ4dk+EbB9+trlTGaVrlAFA2QSUi63YJfEjVuSqzNqor2ECvOJ9KAgjmCBiHjw
oMGITaTJXdjrRnUQ33std2YYOoNK5uBLAofUwucSswuD9weGDzZjxbzaQ4NdTzm0AECpoP0POyIZ
IvC+lCrAg6/VFQ4UEFgkI+ZhHrz8OAov6HLYtYM4ak/2c7JuRnyHvFSWuCU2KlexZto29VMMYaaT
nOGxrgqpcjbTvzvLdTsftePJzaefK9+ND6/V/pJRoqQJcqGsDDXcboVvVB6ozw7B+uOpfO8jNYm8
7Jq9TB3LiGalAZ5c7iGqEvU0U7PqQsuybUVGNwdl2VQQm6U4FMYXFQhdAH8XguKkcck7d7EwNHUq
KDn6w2TFHy0e+uQeLpTmz3vQy9NG/qkUow+HDnaYOcsZ8zmJXQXRqpS1Ly6I21hJZiwkxu/RLsfT
Zm1i3q/682+x4E0qVhLldCF0XwTUPt+oUuiCxrJUMkAeLPfLropOYdNbhAX21iSu8MsckltcO3kd
oDQndA846D2przyA8cI7Yz+VIJn2JjgDeyzJY//V2Qp+me45cPxceq3uS4jiwNXtIQKQngRGFV6n
PCJxTvcSEKfVlqG/YQU1X5HKfEkSgssyjNDxB/wrnFE8+k7CY8B6Fn4MGHuKMvuTCSEfTUBj6lsA
9Q7P8Pqr6AH3AkwVxuA7O9KizOqbDFe5CgVf6K7kX8do3TGeX5JSflFuDyOxXV1gJjCB0KN5+Apo
ZyupZ0vkZlpaflYjlqJM3LokskRrxcvFZmaXOIhbnEVHigXRmO4NdASdoFG4WTEaKm53ZhnaKfUH
BsWOYetd15J+axDG9UxJuj33XHSEjkxexQRaxLsqGIjZWopbt/ThZkK4IlEp7/sZRLM4LeM7bpl4
gBtO9/0g1wfrhTXF9og8cb7yTdVhPVz9UUnk7zs7+hcwGy3vGXW0ScgoFi6mnkY/7gFyAbU8pB5l
aHal/Q73GgMFuv/AwUv9n6k1RkeVpQw88cN6hs7OBABKgn22XDdUkZUCZ0N20YZMdipN+mOITe9I
ZDoaEYCPnVQTV7pc8CGfuBF9cKiSsQWHZUEfAPIDR0TPcjcw8xIpECni0y+TqqefETlXKreqq7yS
gqVYItAilSTHftHya0nha+psgu6tDeuoq4N91he3QnWv0+AsUVtzw5qDqupYeqVUmtFJqYOJ4fvC
tl9mgpJMqh1Nlc0NZSc+wqbU6hr+OgMt4bUmTM/IfaEAn5fDVPh/13QxCsru6yi32hE8OsVN85ll
cExYf6aTMvJEYkoL3bC2vceRm547Aiq5Gfr5nmShXVpqCOm15I9BbV1jSBlx8HWolNh2bslJOx00
yOidNyxTKpvBoTXOYcmLJSs8aaVwUC3h49B4+tuoL814Wl70Rnn+j9eXlj15gdfXhlk9yWd2ELNn
8Expwu2rnVUDoV3+9f/ztHe4tFnWeOioRe+o3yiMYrSJ52AWft+MHxDr+MqSsOhpWEFKRL/YQeo6
H+5KNvKMjEoKOK8SDDv3s9OmyJzw8QMbgxOlx9app9qYvTNNQ+kEuLAmb9beBqWPUG4YiI1vvLmo
6/67xmvSkM2JcQjHqsoskDCltOUCvPlNnbX9E8s769PBMJ0Tm3bSSHG+aJmJdmUb98jEpp2bo19v
fn4rE1brLlCA8v8h3Qx0baqGTG616voffR135rfJTiArVHYaGD3uWCU1DiJOs44gb684KDktNDmY
+58z/3CE8PwIb4kS1vqRB4M7lCrbZniAlSidu3CNq/ofKbNvwO+8/wQSvp7ObfqEWvSHEALnaC2T
bxN76HgKBoGoUn1PoWd68MhybLhXNQpEEaqTKifV3W1Sgb0u5uIsDsvcxR8hCra7E2j0vUzewPBC
ceakcR1NLmQBGXxT1FSP24Llr/HvNaceTnZiFeIhBKYt7mCLxfcSukfZlUSfIeqmIF2fz5ufm7Hk
zWCbg3vxzFKSanwy6aAuS/cg76ZMjGBySSAXdM/Z3dIT3qqANP6Enbdk7Rqq5jUMN7NMNO8XgCu+
AIqDoGJ2KU+X04GcyWxewu/ZL9XtAAGD7ZytprNGZ5FsBpjYEMuc0uieXd1t7Gl9Gtx+LWzQZjAB
prurwg18h0tLdZxJD3+Tg8JbiNIr7d+E5OJTXteeyY+fYGTzDJPQbcJWxlcXEyDcC9CmrhFZ0r6I
cvpyHPvYrOf/nJAfSg2cka1N5vqvojRCqImNxe5TF1LY8gkTt13pLTJKNXBpe6C1jf0KsM9vRO5A
bDpu/l/w0adv9dUzVJNoTxB6p2LCjtTVujKZfuAvg2qOG33V/mf9evzZJB/YQ1GCC/HO8t8dvXYf
HUX1Ks5zmo4jYTlMOrw7Bh7oZyZUAW16cKMHPDeqbNakZ3cA8U7R+nvaU2yaKPmDw7tQHDaHiWyK
2dSJ92kgFa+D2iNMWT/XWzXtQ8ER0ob6fufzakpnJ338jL/UC88OD9HzjDYCcipjdQQON+yTw4Ei
kr6UwbWMyvaR5YGpEQFfDfUQbmkRxTBUP95hXZ2bl2wZv6OU+XUzi3QU4yh7R5Cb7q5etqYIt0Rz
kFMZRhqtMSAba+Sh0VXWMIhJKj7KpIJdKhG6qVdoT3EaH/H/8gTiUvIErQT5S2o9Ndv7mhKgIrWC
Pp4nkKZFRy9tuluDUuSPFWfetyXYjg2IULA3dXyvHxjGON3Onhtpwi5HRm84RNP5TUdf7DzXyt2h
Gkk9+liVAxT2CgTfNcuF8lJLqLuczYoBIAjNj1e9EBr2RKBVz+keFHKFjULz+PidVlZ5PvHhj9cH
E7K1W2QsfZzQf+6KNt8/JnspRL8LxL2cPmxZDH9U8xW1oEqvhOacGM0e/b2GIrCfODeIocsrTnBm
Z9ABGZ3yWZjd7khtBr1w05rsn0IdNJ5FqPvXAOwIMycgfGT4lbvLOxQZDL0hr2el89REQF2B0D4/
jFdYm+fKapOLYZ/rbjC+wplFoFgp9HJu7eg8Qu8i3KqNziE4jBRw0Z7xfS9Gbab9A1HHbwJh2FhF
/k5uwRSt0hYdWKBEeU/6vuHGUZ3r0XqJKfmqQiOi4L+FZLum5PjwoB0i46AZLe0aIexi6U7Gq5qo
WTOuZeC+exnNvHKUQY5D+5DkIBfikHp/+1nfKBxptUKkK12L6oOKK2uLLg8KYZbbF4sGlSMgJ8Ee
xXVDXhVJjSXbhw1XT3SdlwaQB35dPriEgMyL9muAlB/zjerDF1B1fgtNBIusq3Vzicyw4A25Fcvc
8KGqtaofcxO9SbPzq+bcdFqz3+PbSIFE1GqAV+x7igBpexrlidAFBEzKxT3wgoZk/gGf4VsfJ/Qz
HsbFbkGKsJ3MVD+y/iLlMi8h58e74XyPG8jjaSpU1X0ACp9v8PNex9fVzguvsE8apQDO7xVoSUGm
4q65maPG9gRl99f0R/pTwt92u3OY3tdnDnUUjnIXJ0xtrD1DSvSZK6BEXb9oMDMKpp49y2KpS6GO
shI92ZNJZHliKmTzRXELTV0aq82WXnScqpAXqBTCgkA/UT5rCBE/i5lRBpdExkgn5M1beYpqMMq2
lMDvqJ1dzpo2jDnO3BN00DuKb7DHQBiOJWTAGjBFtYdAdAt2ijmTfwUr3k0in/hMfdmu5ll0iZDQ
F6lk0iqdT4mBitxwEp8yQrM9ufZJQVqT+mXfBDqkU2jjY2VF8A4JLUoKUdYZPf2sQjIfkOAjin7y
bnoNdC2r6XkiFGg+Xg+yahGqpd48Q2J4WB7JorEN9pKO9GyLBgfwaZre5YoXtwNKQ7ydRx968PpO
3jfmLh1yCjiqIs8XO/M9GjrHCgXM+3Pr/MW9STKVybRR9aLLPrreJ34CPXxj31Qsbz6P6Iwydrdl
RDiiDL44lSmaRPLdMcsapBD19vpEWvVaR7zfaBwZd9vDy+lyJYByGsFaxFtkxxepKvTHsBqoqshf
hgt4QSrvq6GyPJ0mCcA9eIMLyCuDSI7NcoWMnHFAH+rm+mA2h1j+H8yHOZKl+BMSrzqu61A4Rvr8
NydhHuqvYAZ68VhlWbiBtuWt8xgb404NkoTiQp/1ty7I5l/zr+nW0NEKimkyVsKcaygTU8up5NaU
f8SEFBmySAoW75vMTXS7wjw08DJvASMpz8Enid9HFBrDNzIsXCbi1U/7khJhIisbDLmQuAaHI4yT
IgunP4cL90OgBFNd747URm1MeyWCOnkFXOS7HAOu+fC7os+nlzpuEgNLZVeLywgUuA2R8TXDCQ0c
cTm5GDEw81vhVXVgvvVaVW/Eu/Pl0+nIcd3NHT7NrKIvESAj3rY2NL40yJmc5M6+hpxtMoyIZ09Y
eYqOUwbsbIuONNslioALL5gQfWyzoPCCNfTGhV+n4YDlV2xYERjvDYWeIOoJe/flVkM2W3lmcE5z
DeXeoFY/JJ2gt2GLBilLK9IS6ZZzGr3OL3km4Xu3tCYAoP/vLJKeahQ6eD08Sb4vwXcRsMHlk6yo
grKDVJIcpxcuNDf3wq4UsKa8iIq4ET44DOgN5ZawbCtuk7sZb73KzlZDqlwvVIKiXN2sNmTSpPD0
5qz39rdt+j10NSI7KLMgxjBR2xMMhdmN5l5aoXDVdnE5M1thRfAP4wb8TB1MmEcYCwxTf9c4YKm8
BccuO8afxlsXtw0TSiTCmx1a4o7cA6YGLftNG44oLmgoN2rTmQPyHwZ8rfvbV/RwXHrtIXq2Tcb1
VlebF/BIUyWHCMUVokZJVt54OPHZiXsliHzj/dKLNBG0wlhP5+dZloEpH0NmhJZr48ZKwZtUEole
gZVWm00fnedZ/bwXM/ohzyWzNB6WReX9fFWQm17yEwwuY8F5Zq9Gnb9CN2yRMzcqJHCyAPv9CIbd
mGYpExDbSR8BcYCmulCuy9A2Wv81Dde2vl15lh7sN6d086VOV4RzrRvJq0aaH26tagYp7bxZ/RTS
XZGIoNAjj8hT75+RoL/PmILI62b3B+fURtylwkXvxGqF9+FB4wV3hjQchkhBRHQCJ2zYH3e7m00M
9Q2oNibruNJbR5mV1ajFlAVkjPRLfAnM2+WKT41IfZovDAZYVZo/oSaKkUcPdvG0djKMu/CperfU
RhGUGn7gT2XsxsKkWcijvmguxhC5/QZh9udjwfAtraof2u/i/OiEc2InTxS2EZSesiKcKWQmHsCr
9CJ2tXqO1evMDb1wYcOL9ELju0U/tkg9vQhX5zO+jw7LQG/eJlTQnaDqF03s22TT5iGvf3Yq+vjc
3sAVUi5XxPKZ59gZa0UDba7cvpu6LC0zkzSCCUYahlFPF/JShBwPPTSMmfEUR43Qa2DGwHZzLjMd
7FiRAsIvgJ4x7TBI4bnXtKnPxfRFGmnlUGH6tCtheP7oPqjXGGv/cjGTkUN2VP5PpnliMn/cdDmr
cNfjriuEbpRxQkAUa+NT01JqRkJVcZ0OeKuffjGBUoxFplw0Gh4UwEhGEnEO8iCuKaNW4Wf6eRJp
XWM9bM/R86vtCSHm8Wn9ObKiys6yKUx2b3EKaTA2QwVZ5FKOwilOfUlnywb3Vvo5ucvcwAbE2pyF
++3cDXi8yXbiBolRmbzUHlK6KmJLTDyweUrOYrBPKxeM8b7cyPljZukqmVgul+lquMIf+aNbf0vG
HJxxuJYdMpXppLDngr+JMUKwHcIwK56JL7ucy7ZBJQDrzk2nObItEn5pAHLoJZqXWC5yvExOdJDW
nLK3RgpWeZ4XRoBLRnJNViDTrl2e2hbX3U+nocbUEwQdAXaYKcLdnoRSVx+i5QzNF7e8tLqjqNPq
u4cNAQ7ojblhWc+2rnk1OAu/xb+0Pd/8HkYwSV7OGiMIKriXje4ITwPS19FQUoNfAvPPK4L0kj5m
HJC5zr/cpDiWggr4IX+sU2eeODkUKgv41HbW9kZ08fq6rBXPCzqi0BewqfvRede3UemwTbcqFx4h
cG04XyuEgWdWtrGMKfkYxKYr032wtd5h6mIRRZUppj9MJw/qavdl3JIfE+Igs9T2+grabCEjl2dH
yQ+0vjSSdlOViPwd4PzxzvTaMH84ZaJwSg12X2256qZE1gNDfB7IIl+YiheIXDln8wHiXd20q2Bf
B/l7XD3C5IBm+Z8Bpk/WYItSfKIfP519n9nmnnXWgXK7L5PHpDG9AmCk8+1My783VFVeITg8ZMdI
kspwAunjtwgBvOy6N/suhv+Cc3U5l3pyFam/NR/ra237E7rGcvXIE35BZSyI8hKAuUq3d/xIvSkD
eqFHBp63bX+o+m+7KyBejnErwmOA6drEC/lWTKgM/Y6Jt53s3AJq5olsjZeCDHFLr2YNZToNmKtp
0UOXuNySUtxskq3y+ZHmpCNtWVjNxBQ+fUDiz7Jx4JAV9gpN8PHzO4om9AFaiV7AkiU3q8jkrFM2
REDwzU8i0bf2+YpqVRTVt00bgQ50lpig7L79OgADfNHTFncv6eXK9jTvNDy6WVP/uR/DGGmpWgh1
aiVK1CiecAWt66vy0/W7R4ifMUX1DFoafZpPwebqfJQaWpyx6i1gEcTjeKDxuvk9hAqMsSBP54Hd
LITNUiCoyAZvSSYEYWA0eIR82bnealgeCGkk+bJV+W5YWt80VOfSjaGXHRLLtshb0AtQu/6Lw5Lr
ByzOuj27E+QRm836lrf/tNLG/sPkNE6KNqhe3F781G0WK8NNZCqwNPtz23FOPkstkpFlN4hT3Uu5
3+C8hdPnV/K/qNTNTEelVnIK8h/acTrlxoAk5fsXycF0wv12Zntw8KUNxoO8AlupjvFZFFoFwk8x
hY3UGp4ElnNKGJFC6eKWWQsizNvUSsixjNbr7pmBAnDwJ9ZCJu+4x18uc8eCJV8SVo1PAVyu1ev0
whaXcsbf
`protect end_protected
