--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Xvv8QcwSUeTcxvj0JLRdfBPEBmbWAvvRVFvwAQfQu+5qg9Q4QRkonicHPQhAYNQ38H3QO34NXYNb
lLvjpyWBxrKl7R/LxgwkkU+QnGw38X2fVV14tSyFq349AC5hUF5/Z15SwMxOz5R6B1BSmJy6413G
slBU7Z0ZWTMHYuTv/U+A6+PvfVutMh51TyJBBkQGu84gqYjLRNa6vkbkgVsGAsyl13Yz/Nu2r5+k
DWTiz+XSKGKGSEWGaWxo4v/e+DX3zv8fWrJ6aB3q8hymnZrpVoyaSUX05EIt/0dvT729ey4oML6B
rj3tR9CDdNQA381hdeTyDxRbMukfHsMbTCfTmg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Beldm2aqCx8EPqCsceTpsG3pp5IzA6yd2otA86/BheA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
kacaXxx5g5I5HPe3lCadYQC6dbH5xbeZWUT1XXe72oRfy1qjkmLUR5PNASCZmFPRaCBQJO+3GSTK
9VT3nfQ6d4C14hnBcA5KMP0gOG99s3TZFGwFekYENek7yP82Ale9DpsE5GJ1RHiPCK4I/wVVZAW9
+2OCntHgs6LeOl9EdMopU37bFFSnqAlJGpOrAYqerPKicwNtob7MG/FNApI2Irk+qJvOfncM8Kvp
X5DIS6RlYuw/uW4Bk3Ub7XWARjgMxv7K/6KlK28PCl43oCzIhomvk466X5VweOnspHaoCEMIuVgX
RUsDo5QbI12FlvxusxxbiMjWPDRYEAaXGebu3w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="m8cm2Fhb2aAd8VFYU5ETBGwXoLj6S3ur5DEaikysZEw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10048)
`protect data_block
bGFuRQ6YATtnNw3JQkM2Y+i7b787DjX6Fuiyp6gxW6eyo6VBtHSjiZfWoVnOXb+yO0Vvu0/a68M3
gZ5fwHoFmJNa4baMsVfhmDGdlnx5/8/LpafLIZ+YJ2Eeys52lDlpXjRka+41RjZFsopZOecksmmf
E1ajD4ihTdjMYWwKwdDVLBOdJZIZeBiNTwKDUqDJw+cd0pJAQonBIqZ5lC1NTN2CEiMwbl/+GmRN
7Qg1Q+27epXCYBEVL/DW37hox+e41d/GmAEKmWfgf6Q2lWwhvIIGwWqsYSXAzf8ap/Stj276wFQJ
zR0M47Ar7UpaSj6Nod28H/RP48vPnySZpA6Stp5TGDQ4X0gb9YSVioF0C47u+8kUO+zdDEAVIpkV
YjTIXKNCeCvybAysyGuA49/87wpci4fPVZ0mRBoAK2QOmCdLSfAvmJtlFbWaGPsJSm1P5Wp4iGuU
8iXWzCeOhvR2KztlyVZEltMZh+x6hSfGldWip301UsSXuyhgo72+fAp29ZvijHHH9flpTrqOlxx2
YEwY0o6EWWDMY/uP4WqoXihFAl/3zdbPC+kVwtcAiZx1LR6mW3VeIe5p8vBBlQ73Ji3EvW8PIVBS
bQgM5G9Dd5BQFtX9Ew1pfVeA9wbHhsalMP+U1Eh/NH7fKBD4kfSIZcXt5dUn3WCoS9Rf5bULSs0w
br6lhdDZjM4cLNcb3C7IrcmLiwV8Fgk1bAulLks0p/WwKVZUrl4cFNykXUHHQ69UFjE7ji/q0SwZ
NgiFsQUuH2RZI6dKGXI4KMqcRBvntshvBFZa5ajnnuWR2ZnNlY+KvNzkfYzC4dwcNzwVi5R9Miq6
OQWv2kiIYEutpyHfrl5gFbxwvw2Q8SJiXXGgtlKpMDAB9Gb8YsXjZTKwK6B4bRn911O0h9iLLf30
+ijwsIjWd7x49W4636+wWj+DFfridUVZCDR9asJrjhDtlaYfve+ekq3AOdiCAzXCvkVj3rF1s6e0
UHTe6KRyX8uPRHqXyZ7AcZidVaQ1XPi70Tk+Lm4MSog8LyJWCe3OzLxztp4ZKxpIMv0ZzD6yKCe9
R0KRZotnU8qKdaXjQPntFyfxkqHN6ISXXH2go05eE9lcCXYM9G46y3ZGIT5sgZxc9SfnH9VXXwvY
PbA04lSuseH0TqpinbveDMZ7IuLP11V2RN5mf/KQZFoPdvRdpzpDTpwGnE5VJHZY54joByawFcJW
dpURg8XmSEzQmI7y4YkYJz99TD16otO8qzZKuUKNFMfyJCctkDzbKT+/KHjLfLiSKQwPY4iTmTFV
3Fgegr37Sk/2KftNlFkSdqMBJsEXcrCBPE+rtLI5nQpz7QG4fl5Do0xD7ULH3gfYDbzAYMr1hLpQ
gatB7dapi3dtRp8WHaqnEViHXe9DkMQcC9PFoVsbblN1Dz31foBjBVTjv16TUjOt3BvmN//swV1z
0kvohq1OT12HYVpy+jZjCKG7RJfB9vt6OQ0Mymbtma9pzBvYX3M8z5+K2c9NgXQLVe7ZEkUXJ2Wb
mXqS63NEPtfPUxbNTfAOyMBDadeplcz/DkRxhASAzMN68WAuwiGhR0I81sdiB3GXnGnAn/DrmcAc
gJEFuJdy5E/PrpfRyFC3gLGweRdgfvfcrC2ZxI/rloVIu7z7gYDFODKkzSx+oljBFx2/SXrkxVde
02ZAPXbhIsRuQt+AZkZZIauXKEFo61ztsRVuVtH5gxXRAYV9L80qZqeEeikCVdpP43akbT41q+z9
Lvc0QPxoJeGtUYrBx/+evmHFShT+iWYNGniOAoYxkok7VYOSmyvoz3IHXg4T5f1Q4Hlj59XwSGiq
STj18Eg1M4QOMMM8TzUd2O1Hlb/JoraoS2dKQ93HSls3WqbZpoizGrDf69q2nlOU5hxDOVW8DYK+
iyUe2RvAI8KRVtYdpQT6SOd1XOiukpxn8rKrOKxLODDuooBxGFKHwJ0G+/U8/ADqMQHFEJsVoQAP
X2qBJ0Ea9CSqgL+Q/FjOcqCB6WT6oHPnl3X7D97kFAokJJxGAixMGGi6cY7FQykOokDpiMkCMt7W
dQg3LEXZVLz6E/5JaecKwFfKkqKf2P3ajpSTJOwqOde3CoFT0sdo5TM5DPUKKNyZluwGflw5Ust3
uvJ/Of2HRHoL2dCYVCruWdfGN+Sc5eaOhi8p4loOnYAN6AyiETIP2TrStrEI3+XWsJjiYc+lL0iS
09ynQY421ujreMBBpCJ9dQQDVpGaL3PriF5lKeIKssajoih6JN11rxSCAKXpjuviLzYsR6FvSmNX
/AW5t+JHX6a9qRUCcTWw8yOF+Ryf8HaUnOwVOpF/rCM3RZjMRzDJvNBjhAEbTcfIoKYxczaaHOl+
w536L0+nS7Vhq5OwH7MIpGy38pEzwuOIwgnLhYB1gUdum+ATJqwoPYWTYen82RWuPehxpgUrY/0U
LtfWe4+SKSuH/AtN+N+wucrukzJlQ64RdRxWTwV0ZsI6BZG5LzqrRLLXVgZJGh1fVA6AXu9y2Tbc
vTVdgq6knUVvMJHEsxvwDd5sd9Xtxv2PCXn+ZSvrqsLlnS39EdMscbVQVoFv8Rabs35mdATGhhAt
oHtyMorjNpuOVlgE6UBgKUQNqukvQww9AHmt5VOuJyFex+2AiR6yny8NTTaGvd1y+wli/swkFr+u
UqJ7qCzXYLiLBjnbRFe7bs2aJHsf0j0X3x5F6DhVdBQeSorPbH+Px4XaWrQLBd3Njotz5uYb9nbd
EAObX52mOrAErnaaysPzZ8/LLRa/LSNO8zDinRfEhjdX6up6rWfVmBMfhgeC3VWbx+hludXCosoM
9y1ChupkFgt1avmafFsH7uIzyIIFHdApy3nIEkSdOKKohmG9SY5MUBl8pd/NUC6rYF0ohlRYzO3b
GG7JosFxP4wtXSkJF403M018HfGlPMCkOCnMpU9QZu9DdwOwAU7ves8pSmT7D4XNIO8f9b36N+w3
c2W7ngr2oZQtPlxNlmUyeG4jBOII6xhuB1CHfCkq2HAAFtyDF46QG4vcFdwXO6aZPDQr11LhJLlL
z3EX+gQ1eSs8xSnaEkFxSWzlJPOU/XAz+t3ZqJeB5vTVSfdw+WA3tanSBPJF19fLaGpPouO5hBB1
iOOEbvMHa+ufpeNxW5URYguHWXkYxBvDZbSyoxy7L485w4MNNiqW1v3doDqCd9ge7/lk/4PIv1bV
4PWMDfDPvNUAglSKW5w29Oel/gQjauH09gHiRQmJM5S9BATAfmRRpSYKPBq4V4NTPTePDJV0BkII
kRkFbsM2B+uOJMe+6boeM4wxlpRlJD82/vOlwI5c4GnRoTc66MlyzuiLVYz7UAG2V8wo+uFaIPy6
JpargcFDMqis9xhmLGw/MGSTl7e+Fp+unsZaIgkaa5El0GS+XPbGX+Ze0WzfL5GANjn8QXKD98sV
B3XHBQi1BqUeBTqsZRVKIPbuuvIF8KjRYkUTmooYIWi4iR9Hcin33LWw7twWaInJPqqadjon5LiO
9y1nAWCpKG5e78kIFFsvG3x59D2XogbfaPkUGQftoxPAVPSstQhSqQItmm3fv4yz55oJyDpciH7P
W1M64f1Mibr+MSeeuGFIv2tp1r6bl6VfsiaZCo2347KXf50ZU6M87ehW9FiNERMvj7FfRRSbpHmP
oULnXGSYURyX95wMjhKYDvPdBWaXwxI/68NFykX1utUH9Yp1tacwswRN9bQgerineSRHKiS5Vbr/
l428gyLLVZLwR9+qUHVMvmSRYxvomXdqC4mpsaMa7uKmc++0FAPQW/T3rNo1AsQoIqWo/JiNw4O8
f//twjLifS9QvMctwMcSHreUEUM3we9bS7OrlWoCkecd9nGWCK9LNw3aqe7z97IcpaeoH+uG6qmo
mCgpZjUzPSVhfzJ3Eb4fyrJbMs/SabPZ7hKmdrmMBl6JqRXwAwy+HXm3lV1/Yf2J9NKL/yp/VO0T
3wgtjxRzoiP1T/iOJDLeOA5n0LrWFUL8yH4v09A9lTcL/UK9unrk1ukhj7daTQ98c6lODDW96xd6
z/BG8zOAjeM5LiMXU9Anvmxhtqng/jtbJmHTNydh1q/IxPqzbOIhD+NOqBG0IvwK3w2EIV9PuN2S
uYRgCNn19jgmidpNDNIOCO3xQZ2VnA1wgs5P93CvIR9QUKc3UaRydFWCUL/6UpiMF/gh3nOXb1JV
0+EAHrvMXLAMkg8lpoCqzxEG1+SOdqAQm0z+XI/w8hbtg+6BpzRzJRc01zeZaJQqdwWg7p8bJGk/
kQ1IbGFdTJzARaaTArnJKYmnWKpTiN9hbpvfhqTbBGf/M6eoWUHUykx23NrtvntVe6ZgkBzgw84o
rUbdrJsdvjgEZkWAOVnHb5HFMKoWvFXoCiPdbWSnadgS3mKKYzsfXg+Ob8iRqLDExoceMqmV+Z8Q
ri9h2GO1gy1n7ZNRAAdPgZZdkNFpNaUtc0F1/Xyaowpsf2IlyFoOBRYSsh02Xgh71r3jltvwUTPL
Cn//KcZSn3263KAWnSmIeKuopjR0Nk7c0LKxazYfHcfp4ouAoME2RSisKK7bTN5oN0pRkltdoFMm
gA/lDEYemTdda+yK5UjKklsmpiJOsNHA4gDn1mN1+wsSLuTFtE/fFXQ3FvfWMmAKOLL0HLJqZLIW
jFe8CHwYCYKteJ+1vmTmEItqsjokJ7NkB5o1J0rTd26iFAX9NK6ps4WZ8Np+DuejarbuUBnIOQfi
ebgF1gRVLmpABWx67KI9ScMEozvV0ADWxL9naLoRz86cQKHeghuOt1Dz0YMwc6+C9YL5tTJpwRpK
9P0n511tdrIEKjF5NGt1q/Ica9o+YAkRHBRYat1V0B3CqTWBI+PYTfvPJhLM1ykvgSSNIcQOHMDB
3WvduwfACKlUfTgMMcuctrt16z+aMDnTqOlky0fgZY5jWr77kTt16eAMBpuLZ34GRVJdR2ZfT+ic
yXzgDYI9LGhtgda+9Ml7hO4qL6uPkW3sGsp+x+XfEyM1Ms+0oL/hEizN91wcn1DUJV2gCDoiklVC
Xf+JH/T1z+7G48xxQPyabNy9bTe0UwTFn1xWYCibXdsRM5q3Aj8pFfxZ92QsiqL35BBkEinkZ2bI
ZiEUZo1vrlRRGu7RtKRvwIo6hi/e4Q/PcxkHCP+KmBQ6tIuLnmEyOCBi1zXn16Utsq9x0lzsQe96
KxXFU6ZBW/BC2mFt4RzWghDw6svYS6zHmJ6GZxUA/qhGnO3D2XwSoaCV6fIbBfUtol/oHH8yqG3n
jxtq0zK5hQqP0QnruOfSO4TsvX3BJGZB4CgyD8ZYLK109OSmwQEnb3ztv+jodDQMgNme1zchSPlN
3t1eXtfJ/HuRIuC9iLaVgD0xEUiHe4ZdUogA87Rnfkxe+nr7lZNmyIgg8BF7udgv4tY8uLCl9tFC
kG/4TnTUdDVzdscLZlIgOdFr8zqQX9gOGVWZRq+gEdV1phLdyzvgo6d3gQ14eZh7suhhrG/RSsgl
KmAmz6CuK04OnhZ+13TkDo3gdNjQ8xrTOLn1YnyAhWmwh+jnaw01jeLXwBKuKmTi9ffVNoHRCKgX
Hr82kt2tLE2v+Lv90zAl0WWuWxjlyBAVzj8vlybBslb0N86ZNuLiER4ii51/7+UDFqzBgKlwRHx6
8Kx5QWMNK0gVXRB3rWliEtVW8/xCLEOWBxGgnKIdFnbR1hRDUAyuFvIwVWxr/8B0jZPU0DWHDLgY
MqVfRq+Z8ryeSBzgsq/oKQIwUG1tgtXo+9XMdxaLvoiUTi9sM3bcZazAkgawIhyh4hd6vnV81Y/X
4Fw/0WYXyIvOOFf206q4Nw7oT6tXR6v40AWZW9mEhAIm5B740/NdbhmZIXpk9L9DbJoINTi9Xgud
p86+y+TxNb76Xk/KXPp3nwarV7Iqgo4amtuE4bxbn8sprMiZmhAS3wnO/byx5T1+G3W2SjFb5qvH
O/bqv9VPhy33PyEv3gdqEj9v7UJgFIBVMa2X5xEu7WK8+E8wQE6iRilsF1OYaEkNmLGcA4n88zKR
QpnPV/hRxLy+TYMutYG6086a3HH2z2U4ApgtdnoMuRKoRRTmz/sZ1TO59+TncGr2nkaXcbpwrQBn
48UEc2IQI4fDfPDeTRIEiLzCys5On5jBQ1WfU7bxrCyzQfK+Ncw+s6AAOXNp4JGWl+oXFxgTrCfx
QmpdapAsNyl0pkSdmPMHb6Oe1e2dfBg21Vf/njslQPtQqcs4NfbMat1WkKaVQ+UsMufOyxrQQCmX
8mdJArQDFQcHBvruoQJelo95QJLdHW2T3icXEvV1qQAe/cn2Eb/W7FlzAkd6ES2HsqBsxNbE2KaW
ZBLLUUcpXSGXjsmWkcJWOCYM/HRpDReKt0Cz/i95CEdRPfcHpzM8Zc5TLTpzURxNWJo326LI74qr
GpHYd4SNJ+OrNYjccx4FkJ4J+yCpor3WyolmO09JER0Jr4h8f2RKHbzZlOwAAV7hDJD5I+JzP7TG
2w1UatJ3A6/M5WyxDItGCRPq6TcmSCF9rVxMX08uEMKjlOcEfIjmFYpww5DsNA0zzSifBLbges+8
8T16k39ZqSykClsJbMvDoiilNH46YGFXN+08w4Xh+mT2lsueeA+FIre7Y6jG3BtKQhmkd5oPob3F
4psjh4+4HuFZ65wRzYN6DOvR7zWeCVQnHSqnEWEpwRUPK2Dd0p3+blsawJI4b+WR93fFUEpdVnZC
d2wCLFWX2Z5xzQ5E7Jn5w1guXKYYWaWTb1ZFmFfXoa729+fX16AGPFrvRySuHzrmz6aNmp6tTUaQ
k9uytTf7Sfi66AtNAnqwK8HnnvX6g2jhjrjj25QASH9luH23+YawDxhCcwfA/JG0TFKjalQobYHj
i9P548kU26z5xaV65fufWQS3xaFw4Zn7TTiyrIDaExnXRdszpw669+eij36mv/LVYlzgWCo2nsVu
gi8V18KxXe6IsIZd2HAYFrvR5Gnn9wrv7bzN11WAgH80Vngl/IbFHJ/8TFeJuw3dIHfIA5q7Lhyn
PCcm1L05ftoz8Zo0+LmGeHG8fRneuZFC1JO5BLSlopmUgEwGLsEtupw4SG8MV5Hd9GcXFSUt3IYk
seYYFSrARuJuLg4mOOSmWHODs9oa92AUCWGRivHY1E2MsB3wpfhQt90qqVSlXcnzhXAMnlL5SaeZ
p3e3SIyx7RJjPTb3QB+4zMP+bksq122n5fjWLjXEyNnZRHZn2qetLvEXnSub6eKpkCorRAonuYYv
QWer46/a0c1F646jYA9MT4Gkr+jPIAqoizCJtmzUpqa5orH+qnshznP/0ye/N1G0XoaPBGeJBvGz
Dj7219RY5U2IM8DgiPNrqks93Sk8CmyyfXWdXFtEqKto85y6WFIbjR9+UopOQR5l4AqZUVPbnS8w
Xz12mWc7rKCjfUGSnASOD+GIMPPsaGiGujdkrH548GowJmj8mh2oTa9BSPJgGVW3f09ZXqJ1XgS9
YiGMluFt2T/kuzVINqKuhl9m4s2/Fpxnq76Uy9d+36ZAv5Zrmd9ILmUw4F6SSVMnok11tcIxmb2L
yCtPtVYiqPapk+UTrfCfYMdpda/TKEpYk6wX8JBp94czntXeRjoh0bS40CsCMpIsfrasRtbmzBmU
/mjXouFFoogOQTtzEsXWhp0p4Jfd8uqAcZI2x3ASuWZfE3mt1CgxnFCDqcSZOHC/sNIlgN86Yvxm
yGuSlLhbPE5ydEzbhuA2IbK3oWeItYEiV4nl+oXOwKz/DJewsFIYBsDcyzdr4RMrdFGgu23AARzZ
5L6KY0+hbbI6aOlh4oKNdwZGUJfulNIrS0HpmFNmqqb8TvKqltQesUSWns+lGaq2rYS3Q2O6CRVR
NtNEcW9snJ04ACEvq0oIRI8YWlaOvV1763/sU2sUMbKf4oLv1h1DcCsYCYraSCub+y/19x1np3yB
tZkWfeQl6OQkZP2hjTpRo9224745Lnpq6WH99OAzX+PIQA9XVF0Xcc0AbpT7S8l6AO21D1DqC7jU
XMbVXKvGbXBlnYlchKjacNP01Zsa8kcIc3a7Icy3Q5ySvBbJmYZtdbM331eL9oe8ijIsGu5n58GS
V1iiH60jumJKLdm7N8rPV8wk8rHWSClj1G9dw2kahWZsJ6L/DRGuTWYMz847t+fxlQsdNycWuM98
XuZuEZoTBuwifR7Dfd1jR2A1aAqpiyxWC98Xb36sNUG1sjuGqB7FS8n2OlJPJQeKRlkUSSoZmAC+
FErXoySCRhDdVB7HaijQ/5JP+norCC9c/iIxOQ2nCvtI8cGCE+cGbM3KDn7cY4G0G9O6eqZPWEjt
vAOMrkIVE8IUx7eKjAikUf8puhxZCAI06z7VNW0Rof57Mh97YEEUvB++chK4ZjTZnTDzOSQ8oPdB
sdWhiHYYR2oVhIs2rsEfGBatplTZDHrRjq8WVOSumeV1MivKj2lZKsVBcno7S7aBQHrzRTgjQhaO
onveQEVtrR1titOHLSrM2vfCTYxwuVM6eAqBfNvFvsyxFjx82+OrE0dRBXBQDrJc3hcd7T72AjD1
Bq9ngGU+CT0Nm4aHKmJPYZ/PyLW8KNJOsXQYzoZMJAxgQ7W/NQAtc8/1LHP1BFNhBkm0/SYMw//t
ijZhYsyUtT13E07ovvLE+qESaRNM2cXJnPhJL7qepRdJY86/Rn5h3Xk+zuPKMXEJjWTPJ/mi0vZO
At9/OFHF+g5KljZE9/Ji/TRxCIvVnscnK0aYxWwM8nRzumptyzlCdwVM4cQ+8hNwFZAc/iG3Z7nx
eVXAWzzU83TT60HMxv1PIVqN5z9vs8m4H3jF5klerFWes46USKFGVO2JzEWwfR/3DlSLy/A/9mnY
+10zalxlvgjZVxvxy1igeCiH/8m0DWNvoOVljeY/08BsHx/VFQCwNoeh2O3kuMokR2KBhQfDX4rI
0xkl/pq5Sk2uHyh6wZOXwigyITMo9pgrYYUpXYgwCIJaeY8R8r1krHY16PedJS8Zr/dzIFXdqXPQ
7FRJP1q9IqI/COCn0C8WKJmc+dkxN4J10Lu5EtXXuzG4xxgLIfktDCVHoFVSmsxVHkzZC52gnM14
JhUUTMTWfJnLn9UqIowSsmasr9R8qn/f8Iz6BvJvPEyC7bvfTKnVser47Rw+k7rSOLHKJzf1PoDg
m1A/RUAKRVziaZoqhRW1Ftz161omYw8xZ8+NlSZbLNzI6fS5pWMUJ7yRBjLxDNyW5Ip8b3cg/mAz
1A7pDYV3EEw+OkCHPfcxrX56S+2R9zhAmOC0C6hZPCF/vBTzBhmTVqH0IXI7ge+HeaFhEAFxw4Cd
jyU51XUhhbCwl4CmJRhhQVpmZ98cp+5XPdXXpySzNhgGbLQ9maajecnspZ3xK5ZSnBA2LNK1WWmI
uEgG6OHCyD8HZeDmhDIXZ7kVz+d5ZFRmAN6xeU5Kkv1hspnpZUDDDmGAypKckg5LETJl8IL8C3JO
UmECBluKF1LBqemUQNKuJE4aiOw3jqY/VP8S7iQ6N6sXbD2tNZhlXpXIlzzxGamnZNpgdWBlxOSZ
1XSHRK45T0d6teihoYqNAYXJonsgjOBT+U9WFySl63YVoeJKZyjcapwyvwMCzYReRpEKWwbFZDbR
Lw4hqj1EYCZ/CHu2tNTlgDjak0ZgUsCzpMIaFfk8XYjheRo4kLURidO9JlvYPNgno5b6ZNzf8iTc
v7daQzrb4GP2j4JD1FAHIDHWK6hScbUkAxse6+hyJggbnN/p6Tolc6HGvpnwvx1iA+Ob1ed66aMB
3KemNlLil6Y6ynTrMvGxQp20mHQU7ZymH2804RqPgqJAjeIzXAdT9jEXPhkHaIqOFXEFKprluWDN
tC1DQNDrjbVdSNcQ5srvyuN9L1GXmNY8heyZoZFQlcvMRn5o7D7L2LAe34R5QoBK4nuDMzm1T1EZ
CcNUQXcKJqeeTRHuHyAtpB5UgidPIrB2B3T/J9cBdcHNCEr5EdNVcVjv5yM+zXbB4oTbDpXdKa/S
BT+VrjF6RnMFEkyg3jQ273lAYVmouVI89E3HFhFCCOlFGTYO7OGY4Kjwg9/9oL5KasFjIEIE+yq4
xraVTVsCcGdQAB0QVkRwVrup73puW2UygMvefk/OzKKybrhPD2LfE808o53yUutTvyFNljFrBaxA
kuQR3m52drMqFF6YQHVNzFXAhjCTdKYQKflyFDvr8fxibGXialBKgHQCPK3qPcLFGrEHD0aZVoXD
pPolQZuHWLVHVAK0SNm204vlp8iaLeX4IqnKrdRWIpDYPSwUbY5HmtCw0HwI+B5nLlWdFHgpICfq
GL/N5CLL/ThKMZUWGoKllCid93SsTDIzar+0N8055IdRahftMiE5kRcvM8ggOdDqJ/t1DwC9a9lT
Fa6WluoJN2hqoekWrPIzW7ilwxc+OumpgXogmTHFZwyxPLJ4vEusysmPmo2nxrT0Ry3f1xbv/5Dg
7ZrRLDeZ5bTQqff53MyZW8IrwSBgns0xAqJqwGSVXbDzrdY3UqIE2mISQGVr+zgfnQHh/a/hQcHw
f7k07hIX5C7eZ1Pi1Ukd/QIG+LzqNPs4q0PLYRwYWiDmNFyCy5xqttUDDs3MLAyQdnnkDhZ4sBH9
gn4iMLRB/OjJAemGd9kyhl9CFMYhO/gG14yYY63NwA2dcTOqh2MEYpT4TclPZESnySBH+Rr35jrx
fwVsHWiq96bG0iJXp7JgYigUk3xG2jR9GKZwuMIfRG5h5tZaqBX/ymaiOA+sVOTbo6p3c0OUk4qG
RClr91OjriD4cEcw1mN1n+A8xCauQtBJshEc8YNE3/nzANu27RlmNtUSQe+/1jFsoAyXFu2/wWXZ
J/3kZ47wwug4nhkJ3CwzFtrtScKZ/MZ9hlOfQYTLq6KsB/X0klbvNSnT6J0fWNARniuFoGyaCl24
M9MHF4+6bTtkuvgXEBFpLkQRP9fPpRVI6bgrvRpKr9mCz0xQ9BOQC3GZJlLJjgpJlpSyWUGtMNH2
rC7sWG2g5HWm93BlUdF5j6ZPk4nwRqhCy8s/8T0OeEuxx8JJE6eTlv2vlnVFW+6Xhr9aYcVnBPHE
2F/9KMB1OSRXm5a1TxuyqgvYgSDOvvflUCkTfVSYmjQMutMkV1VjWJ6k1lzd9mK/+Jq4ot0T5VlU
312xjSTvDqDbjNWZZICmMzi43gMk2z3krVzqxLCWWGENwJcsqbV1oON4x1WXvK8oVfIbIqYbNXyE
K8apTsEzV7WfB03ZaRIV+mUx+nkJBwGFWIJmwkWsg6jPzCFEemto70Dzw5u43hPz5jBQRuXc3eRz
NSPVTtKpJJXrmAV+TLrhxStWIBjyDdWS+7LGwzlqYmw825K8/PHsF3L4ZLue5hqGXm/j9Mz1Wj+o
YcNri/tOFaXtcZiPg3C9/+kEjHSecsfNenT+CVnWm7X3wgKOSQ8CmethH4pBjfSZWvdCoL8NDuwm
q+RYN1Eev/D1z+KxggcAGdBELhk9olpFrVRgqeK4m5ZKczqhXtQ2nQuqQKzGV2sQ+Y4NdL5kugHO
nFU2JRqMGwhyw0ZJ8IDWtPifamP8P9X4N2EZ7mjrGfi/sr5gBpe1Fc4NtBWBopcxuzlkA8oBYZZZ
fHL6uexDaTv4g5iZANXz12SkvkLoLlBDsxZ7WrmnfpW30HxfLfBxIPf239+DmN1s7SHgOGqm+p/2
uGT+7kTYzHSb7lYR4tPBhFEzOt2mXGhLDjhwkv8PLmvwjMqHYHxESxnv3y5/smALtvrX2CAAb1pK
FE8xc5Ck0xQpdcVWo2zPibWxvBNLQYNDn+FXgQEj5XEsQyjkgGWqT7dU4yMecktb4lp1h4QiMIgg
4CsCncgD6c/+FajPdoiFS1CFzrnbHNSyZmx/C2Po9f4GlM4cxroZ5EX+/zvglZN2+kx8WAI3JHgF
f+rmus40+69VTOMBgSdM8IR27fjsN+Ij+uiSiuf6RiDvlyB1hPVBcnY21Wgk9zZrWl0vA0EAJWN1
9c3MS4JAFTIWkrSulIhqE3bfkFNtLoM49fJumhSinv9/OW1pYuivLlySz91ZTVPbL+zLTZu0hu6E
/2n98LYre8b+DcbnKf6ZX2dq74Aeywqe4d5wlqMlhBg7fw+TO4C0TkAI8QDeCYWf1SkEgYJzwN8e
OhAWHuRUt24LH/UmBwe/JP90XgkH4Pts2TKEr+Jtb9rkxbuCFNNUbpJTZCuQmBbwjolN7WeURXjS
9lMqJM80UyCcIuQGYnWhuMM9+K5nPDYx/BKHnJsMq+UBXmuKBfdQgoNqo2VwItCbsqli9c+VJdFF
a1YHa4Za/nRezc0hgeQEzDCgoPG87rCuH0QN8AyeOEaQNb1zy5795vyrlsKVIaUa3nyXdH7HjU9F
KHXKPblkthmpmBQcRAGd7vggBN2PH8MufId5Eih5k2rBxj+LlkvRwMBACAi3AoKqPIQLWRkRTA9u
kt6pf0qCXgS7y6lM+eTR3ihRfS8i9GUGNp8L7CUwxdTq8HlddSDlhEPvWSiSGCQwiUnFcRkswMaz
xPzYZXdqIx/q/wq/DeGI/HZi8P+Z4srtJMTfjLmf/Z96y8WBpHjaygdOHZ1JRklUeGtREk+APHCs
/dgNMble91OWce0bT+Onbn2oPo196KeJTyGU2rY9VwSSCfDzoi64D4p1TJpm9Mqj52e5N88R19o0
W/1ct8Otgp5dvzgkRX4TBlaXaf0Cl8ZYiTBCWvOVLL/AYbdHUZ/h3yMztNC7ddg4y0e6o/K0uj5Y
SIDf9fSJPGD1E/DiR20Lh0UAM2yIvnimCUM8kGexshx7XqHN0qcI/0a9/upVdtakjCSbUG1WLOt/
Gz6dM1KFn94d47Hio4k3Mn+ZFHhlb5SIc2gWc1d18KpxkWrmmbLl8FWEce4yYcMxMtUWlPPPBsx2
QWzAJdGx0SrJASRSmmXMlpxVAjhs09MaYKJm6TUSQ79pP84lb6H7J2B3QCkrtFN3Ies179KXpIGX
/Bq8b/UZz9dyK94GZZbT9FkrZJXWQ5gbP8i7oCsE5qJBFIPHM9dYSvdKkum/4iy7/YET7WyLkS2/
N38mmA8k9vAnHLUktf+XDTWM+pzInzv/2Y98wdjbNWfqBUxa9Q41lYiw02CAvs9qKHcc21kq2wOP
pL0jfsavy13BUnqV3AgpbbaM0Iasi2aQqmYoMnW49hOTJIjc3CyNhGw+x+GA8QzXu+wGr0vlXJ/B
3luQCuotapi2/Vj9XVS8lTw4l+4UfZdek8+VEvAxiTJ2ENVXPt5VQh6Cl5HtGsEFdJZ9D/wcxcLG
4B8DXn16Zv8HIPO2L6HUGANlcSCp2Gy0CPN1GWjz90hTVyxBQVH3JmcFdP81Q6KmZMHe2PRKP2EG
sS2JUTFyRQYHO7R7cZh4RmIg5TZyHhsdhgEsF9JfKSXi7XobEzAuDq47kiMwfM1RCMPwsSvAB3ix
oLalT905lDaXUgAxT+rbjQ==
`protect end_protected
