--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
gMomAn3JebljJgoDxv8vAJKHYZ/llbgKF52Krl3t/rQ7XJ9NQn+ezuh3H9MpXajPzFo7bv73zg+v
jKgEA8tDvOef9kJOK8tMWB0C1QmcFUbd8UhXfsgCFM4N2VdYkW0oTaUv/ofBkcUKf8rETs/q9dgh
jgN1Wc6n0JsPX/MhrusWoa58WvXQYdQU25HP/VGuEt0fF5N9QGsWJk312/pRWYhGYM2MfiQhc12u
IRMHOYkHPA+vFbynvHI1sIjpaipdPZxgSO3J82J6eCnOr0HGPbydbUbkPaq/6cGO+p+0C6gGGzRT
c+u/WkiXumEmy++m6ER0sc17Fn0PG3QsgTfG8g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="NUEBPNmahajnUBUQ/uP8zwaDoK15l9oNwosJjE6oo40="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
XJKUV7W9Sa/RNrc4BjYerfg/N4/JTGeEsAfjWX5htMkJA7jUeANRKzR+9YLGaJgrBIO4wjCyklOh
bJBEW/qaX9itTYxABy0BFDjc0scWO0DVOgZb0dmvGz34Gri1B3KcHliCF+T73Rg3HInwZQAQwnWZ
65n62jH35PN3nd/ifWvmnQlkbwmk9Z3iyYfVRJien4pzsZsxVJguin1lsBrYmi5JRqoT1k2rkv8O
sRArdv+WfQkhQlqqQofE8k/KEujwWi/9a3EGK59oYxkYQhovUJPFF15QIv1IJ0mnBx9nZeK8ZqOn
R9Y7XjpZm1MpVQQty5H0WH4DYK4vh5h7EAB3OA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="NLzIkmaf4FG5BdF2U/5HrqPnED2g5bMcgMcHFOzq/TM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4208)
`protect data_block
BZzIsjgJADs4JiSgkj8M9MdI4LSF+xBDTaxIVOnVEVNNPfQsu59ep5wpF1uCdpzv3BMqGdRDK6ve
sYon8uvgSTXWqnRFKZVcQpEarNhNVid84uH3ZZ8mrJpsck2G0BtqKwKLmH+P9Zt+FNe2gXWCJrUY
u3yVQOTR5Fj13XK/GdKSz4WLwkkzZ8yOEXLmkVoKORwL2709GE9Xtd7aMuJxmRARjHmVPKhNX6Zc
cdxlXXBxXHU7FXyIoyteGy0XAnNnItleSyk+gpclv+xzKzhcCalu46JKjYUPR71afBel7gLcLnhR
YuIrDblUgSnTMRfH5mtvJHl9EVo5YUnCIl3l3IESRzyks+GiDfidoXYfY1KaNUHi8Vd4GSbadNed
lR77YgcJVMM9tAzNxEiUxwcE1+1aV5zgZGxrR2uKc60UY29wh+SGumx/g+kUs6qvZ5ZRspa5Z30X
+atznc6hupuiK2n8acipvpmpjigF5HNZ3p2y0C3ny51S9Oto6pNAe9wsp0TTpOa1femQg71Cy/QR
Fu9ieq0edyOA4/PvKbgPmGUf2pIp+EmCU9pslDb3RIsG3VaWEqc37LMukk32ueciRVBBvzSGALr+
/gwjmpqA/CenQQVXnmikjbGsXzrrpBbHk4sZ8AUrzR0v0RIjF+Oj5mjNWbzH8oYACMRWtHRday4X
8yS4w0Jj42IwfVGgMwE2c11t7cNa0DTrdKcLtcfi+rzbbuogfy11WmGAhNjRcDqQW9hFvOli+DfI
TB6H9vaCuB6kij9IPyczsjUm8iKw98IRkIQ3dMUBdlx5g4ocOesfDkvpjh9ncgaDVgw2jFhO3pf7
YR6/hSDA+KlSUUvOZHl7jWbWBYVWshk6/de89MKdEAyqsZJdO0RCV2G2Iv7iyg8pMA0YaHdDDim1
GUC2pSH3XsbL+lPtlmd3hc8NiW5SMqrU0F6cTdrTu5P8MGaX9ZctCwaA9g0JpOLrM6/UX+5uRY0/
HlZrjxvMheQSaUAkAoQa9tpvygqtwdxq5ig686xGXe1NU6OvgnHwkm10bZ/JE3F5NH5JkokaG1D+
tt19L9SrpLO/o4IgGJsXc9HbWmUf5nJi2YHB2L/CZOx0ceIyP3nYlnSqdXDl7IdlymJ6mu4VQiIC
Ezrf3bDMqjtoSrcJXf+ENf4qAJWIDIiuFX8cwb48x7rGuw8uXfEe5/BkZNlLVlsUm5EBw2Je76TA
1BvJwKLnYrZQzJk6MskEAF/Ev5VJ18LR+RW1ECV7gVLiYCzXLzeTpskj6ND8z7ZNkaNlp/ElMBLF
jbjz9JSrWXnKOesdmnSSPF01DYSKr79I2BvDdOlwOjXV5aZEHJxDrz80BZXmEZeSrNImSOqUWTaF
mEpVssEEgra+0fi9UoqWnaXM800quH2V9X15plPsRU4yBGbNuaoIS/ZHsZTsuWq1rcGj60szZikw
SLaLU1Aqh1yzigT+8rprOMH1Y+bGuY2cPohwU/Ab1lFgvkzSQARE3jyhES+xPacol0aIiQVKxXGX
baXrssqvWG2Hxyp39FeOwJ3Dlc61z7BcErsQ0GJ3pN8jgbVof/aZnUUtxRx3Ay4gLaPPvgsCpYXA
BmW8IDuydFp6nQvf/gYZ9Ouk4RDrTbXxT59S4gDuticeNIOq3deAm5bG8aNTqD3ClxTEZkm+K33c
brXlaM50GCxbk5RASHxt+29qeW2JLIR+4NRbR49urgosg1rl7LYPA877u/tE0Ra3/Wu/UqEovI8f
D5Id70rLHG+NUe4/xQB5T58FT1QLCmRrzeAKq6SPVv/9sOBfQnIyYzGpLjGZXWZY2WwsqevAlI6M
xpb2ykc0Y4v4rZzjyeZaRr8WjTA942NK3BvxvQM7zZoLpYQ1Bo559FABR0gtNic3OgqcPmSN67Fb
SnWFf9h6qKeCs6vAWKwhpZHNeT6cpxpGTWdkeJTtVPcpe5xsD6ipNhxSw7s7nq+GVXhtYSQrbWj4
ClxNtvccKkfMxLjZtpPXMDuK7XOIKsIb4pXCUDhArkZWWp4zJYdedqSxU5/so8Riw3UM6NuoOfCi
XnOeNtLIJ0S/+pYGOsEwcUB7p1T5Bwkm31jk6m0mPbmEEzu7pk/dDkQKFYV/A5EBBq8clMnOgiaw
kB2TINMwM5GGkiZKpPPRbRQT5OlxCtONK7XshcPvyOuS/CyaRlvkeYjBWNJhkplrN5uCgn3P7Y/T
ZFmcvrtrJzZqyCMIPwRXUq6F3uEzxWFYQPUXYtUeHXwEcgdy600FV+q7LWsPXTlkPikwysYxVeuS
sVIIj+nYL3Axv2Aw3Nxw5VOPQU43QOOZZXt514NHXi7JfM5rzx6y9j1+fR5rXtwpmbYqZlRbSAxy
hUBXdptea/NjXJ+4QpV3uTpPOogd9GWKr/re6PTwGv6kWbmBBZNqDLEo+iUF+4JOoaS+IJOpB2Tx
nm1TO/nMGHcuM/99RgTJK9nBTH4PQEfeTZJ2Zh7SgciW/0iV8mcJk49avbCe7Dx5EoGpGOEoRrHA
7sl+yYY7UssF30P2fXZa7l9vBGm963/4NOXoxgnbfZuzSFtZ3EjC1t1TvEbGo5ehjIPxzCH8s4M3
5Bp5HSAD76Qrqt59GnE3zVWEGBIkmndDGfgfvkvwhT9jQo5AeEBpjkNzWD1CG3lMcju7zGICJ4Ri
b7tzYJ+b6KAC4S1hLIURsWWPJA6oEVXgOlZYfSAdYSsgmbDbo3yLIqgbrRDROVkyI/0WxbWpQ8da
opq9oQdIHAT1KuN40kBX5RVZqEzb7AAnBN58mT2iNerIrcPw/p7lXXIqFzaCgXw14JDA+7/QAHMD
mOiaf2Q8z2Zdijql6kKZ++82AAX85rSKoArOxfX9Mw6MNL+4K5MhxEeHoxCT+PERerFGrlFAMXp6
4KazU+QVbCN6hqJwgGOSFV73tgAxfmzQ7DQ2Dg/YcOrAzutojbkKstg6cLMSJjigbqMaNbBjKFhY
KSLeAFF6dIzHzeWVzQqAkQpXgQQVEQO6QuJ61t/rkOMQbJf3ivB+5f/lGDjvw8HbgWZQ5gTEljuu
bj+xQIQ1mTufCnSL6MlKRqxZuJzACcXtEAAbtTNr3P3MAHE3yhwA1XT9FG21vbiDdPiv+s49x6mX
Ci7KdCKXalBqH4E+t+Zwc5WBAU0x9uc8z6i6DBEOWE3AnrfvQkNBkwsXqdxwl0cHYRKvEuXZRHGM
0t7BMw4hV8OU0p1SDBVcu+6ON8oOCRpVe5XzhKaFEtKeIzn3A+kanPYJPUpmo0Sy25NKNnz2DJ7Y
suD0ytWnLuefD8PXzTRIZ8sMpnVYrWZo2F4q+J+kZZSNLf1rEF7ZPv94tMfCArtq1aSPCM5JXgam
esmkZojf30PI7wVO90EeeWPzOVVK+ktHWl8Df0AiTRiyR/kVYO2a/SV/MlYx54L/kASngPm7ipeX
YZuz6MJ9zEUbU+KzLJJRzV3sXMWAIlcd/7akbJJKI7YBRigs9ZMIwBU3U4LHfL6D8lWQgBpi5YaD
iY0lRE8gONx3tERSgLPMdvXNWHqLzBWt+TvnRu0Dx3AkcBo8VmwUirUwYqR2Gp95ivZ+0aaLzmPO
oiE8dK9GS+H7MmmAmDjJGKhP3h5pG/L/gXANL/7eVFIlGCGhN6FuqRkVE9+qo3lMAHgax1CneJfT
eoGW84thAzNZz2yV8hYu3WzZXE399BDvPybVpuXB8JX5V4PCKrJLHbimZ/wpVcF7OtLuoih9DQag
+1+l9Sz+SRoNKZWtgq7C15/Wdiv7aG+nJaqbxTRbiAClci0kFQ5q682iIC82pdk7nicgM4aS0w8i
Q6OBwV/O5zsCbjXHodaHfOqdWoEQtNv6zwiiKcm3g5fxl/AxKMdHLmbFngud07Fo7ag167HMPSus
Coe7Vhg4IwZ0lBoPul4N0+bgyuMka7baOA0e+Uk4tLx5fWrMT79Yk5VjipUd1qwXk7HcSvWABlyv
bMorUtl8O5PaMF6Fl3To8SNy0tPNHvImG03sjwGhA/vGpj1WBeStTgaMAYBQdCCELA18bWnaGZ0X
VqGe56htgpxhAGM1qi50CG56CP77fDu3VWDjgLGQtKeYXmju67u/hndyhjUz4kvLmVHUc6mpwLyz
FxvJEuQhKBHRNsgTnXFJEs715Zt/8ihoaJZTa/3le71HKyUwTkxUR05kDspzX4pxsgnukvdLqvDo
yLL0C16/PvINxq1D/jKr8JkmwHMbV/hTbvBV0GODoIDUnPZkZuDe52JCB4yih9l8nCyT6UnqEL1l
MM9NgeGpHZ9AWwKb1P/HV0+uwntcf4pu2pge023nJEh6ENEhtFmNaLfQhzlYJ5aTmw1yQicBBJKt
4oXF/g/BZgkAk1v6FF3ROX+2f/YkK4aj4An2Rqp0otAUE6QAMRvur9HX9msQzLey6QqdEEvhATFk
2X345l76G4o0G3XNks4uIvorFjhMejZDye0WYPXgvr7XG3k9fGWf/VrqquJmSzpBTDdah+1cN/2/
UzMrxu4dYrbpplcmVx9BEn4Cha8vro842l+w9ES9lohpPaNelEHxZAT/ReJStkpFaBwE5Z1dY/2f
VNSWANYEryydYre3U5ea6de8l8BRZUM2CbpI5A5r/14R0nG50sYn8+shlbD+0WM3OnFSgZ8s+eLi
+j6Mlp1jUY88W7N7th3O7X1O7Ngi6u8rF+JoRbmN1QHQkawXCs4WHwAneaaJtWkPL1ygz4UyawgM
4q0TZNenbFZ/Zr3L24o9gIheuxaU0/FhcT3WkqbhqnFmCBtISD2f9wz8sd6QgRlkK4bzxUsRUTk9
j15be/G/GVyfW+NzBioI2QRSwyWgXf1woipiUVW9rC/0qmLKtHNZ3Nn/YeOTKMjyUwG7Ekh4B51N
wyASXHBCIDSAwj+6EE/tuF16NsRNV50TakjMRpWPFcpSz81ZM8ytVZaqECbdaDkQQeVIYZUyni5t
G4ySBiirzOTZp6KBKwRosNa7hgk6F/uxOPxyDqgLPV8BZoBzDeI5OvDbtYg6S3z3+DdSZ2+EAvAS
zOXWbKMh6vdY/uTHpurqQ+OvWSZ2x5YvPiR6NHC54TBph2Bs1+mlP8tjZDFPMKboCC9/gbmzPK+u
QXj6EfX+mHuGeN3Ddhae2YEilL9Xnukg3NfjHDaQRx1OI8M2vX4LnHPCEHGnIaPgI0+cB15beH9U
bctVyuPJE7HeSL6x6CgFg+7Y8GcvQvUp+DatJToQ4IrfnWTBdmIVsu9ohrXxJCfuLld0dm60R9jz
F0B+67QqboSR+9s+uUdhvrzo3lOvg5OvehZv/J9KmuxWEc6k38IHJ4cPgSIT9b+sZXonfm2B5BGd
DEhLtckBhYrb42eiLvPYMB+0DTyLK7uNg6opmLSvxVNNqREstggLmx2ocmaI1rTu6IFFmySuQeLm
+JIVNyPAC/gCHpRqRXP6y7evE4Ew1yKJrn+WEUerG9RPjvNX5fK2Bkq7wCtG61yiLp30xU9yCuBY
bxgD51IvOQzvbOnrs2DAc5fsssvqb/s4hTjU/uGYK3s3MFT/mM+1mPftwnjWgfuSaKxyI935rcnL
n49QajjG5eIE4MJzDvFVRFiV/S1KphSpOln3DNRH7lJL4E09aJVvuwcX5QpIUC4=
`protect end_protected
