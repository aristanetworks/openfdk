--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
lguG5UpYS3EA7UN8sB983OAKgUivv0PoPTc868ZiPLW6lGpSU9SIwt4EwHtdmw7CyYdfHLuAE0xF
P3EePtMUiez1h8tlkyoOo+HqEd2RClYRUFDmZ6zIS2/bf5kxHzr0y4Wtck6m00CyOVHdrFEOf5hS
dJr13xZUsOBaHV1OcXm+57/EVMe/SPVztc3E+KnetFrrDEErH7wu94R5z99kkKQgr/tB0Prc4IH7
sxuw1GTFT3/K0z/orayfay2Lo0/yvF3UdYS9k0gMeXtenNozIeJKZSo29yWK0gM4Heb53PpSiyHG
R4vJfnejnifH1Sc7Eqhrqjt5Wc4ievLDg2IzTQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="/Ow/+hblc3ia6fCMmfj26SLQr1t8eoWf/w/nFWzasG4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
XLya5Xqa4ihqX/5zCleLU1FRlsh3vSrVIuE4TcuWr4cxBLrMXFC6sErEV0fqcv3S9a5yeR5h+uYv
lSD+XQHE1XCgJcrXN/N/O4U+MC/UZ3Ylhc97ETIxow6mcrcMW2iNX/Qtl+/t7vn60VIlCw2qPq/o
SLJvlWE4eHcflqUn0zcgwUkqM27tiiZkMg9tCc+95BVwM8fi9jrXdTS25JvzVDXEYob6E7F2fecv
y/VmGLS1n3/iK/nULlSNEJNp9qeMEKxBaFv1IpmrstNZoudI7TZR7xybypt0rtdXeCAGPJf1mvqv
DAqKCvy9Bb0Y0h7h52sMCld1cl3tAzXbCXe3uQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="HK/Vru/PZcf8fdXTM/rC+dP0m5dn0pHm61RRjBPblt8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3824)
`protect data_block
iplhbkyuSuJj2at7ZOZq9UbUTCtjDayOODCfMSFLNZOuU/7ARXAG1dJRM2yZEFQMCP4Yx5LMAAdT
WZK0OEOxIk9HZfNqdlMWOTqYt6apJfxJHJyzRW0bYtk/IPZHxIulh1lOGUNFfO/BL8qWaX7121K3
TMxDiMcjpYmndOgiG/o4fiIDYO6DHBkIcW1TRSKHyfQcqqSwJHgZOOpJdPFZM0TuY8lPDEak3P4t
V/pEn4DDVvO0Ui+jRjMjKvGxs56UmTmjx/yjlno9j+7MyjyO5U4pv2h1mGY40WUojzwn6tK6BBZy
GENB8wDVRtZLa4DkcBvdEptWGKDSaKlMbL6+bP5hQe9hdmJUluNJ61ickp+uJ+bo7PShSyOs/JZp
CuAK5YH/7QuzQJ+AGNEo+O4OgByiZt6IhIvtYe98fnA7+xHAtxX8g4eaKTV6FwixfC/LHBeRZqHd
KXItzlSFiF6gVRkl1SXZxQoPvBzyxBCAKUXYalGcLNmeAKCsSlJTvVwReXR83NGyCQr5OIIpm0HB
zZj/OdOAmUryslF+8pNxXOxxHZ0iHB/vHdz2OaXP/xEMTI2zJgcp0wbLSkZvLpwn2UtI1eXKyqVr
SN853WUDNm4YqjS/VHSnkPQih/Xk6XgsUeS9+LSflWavfn/NP2YAY1I/LHv2ggDCb6VcopFBciE7
WS35TmUk8RgomLx6eLXN+FyY//qdd+X6oJViRXHjHON79tqdaX4tD8E1W21/eV9y/FWmI0HFDWgt
xT2gK92ZVnDjkCvVyrI2P3dsNVwVmRdFBAgszKuYP1QB2W+OX8wDfFACWpbo+iLJjMTXlOdftLNm
00HeYoe/KmyCFg9aI43JwHGj4epBVcvqMileylwlw0HLG9pZG5JIZ0hDNRMhiqfu88xtupXP9zjj
mTLkk5At6X5rpbpiJIPbleg+opESCNJVavqmIWqqdfNQya2aHCQhqJmWDeVXfXHhOofQPwj9lrJH
7M4O9IZll+hSrSy0lOihnIKyf4Lr71UtSk55FU7YYlY31G57hEeUiJ6M5vJmAkuI6uN2fbUrg/YA
8Uv6WsT23Fa7qA5Kgm/a/xkQgROAh9JCv2gvCBYq+nbsHizz0xgCGbkBL4yXD+OBmDyoWLcTprGq
8FzpWLzbcuSJLB49eh/YCu25fYGwWHRIUfj2ZhMY4+a442Pticx6ROwwdlnzY0GNErO+iL5uinuD
K+1VhHykFPEzY4+uvFyp7zGBTGESirCDffmorWU5MYXXGkixE/wv26acaQVX14xQDRrDYUQtl0HA
6L0vzyt2ZPMPSq+TLPckdJLsWJyAHe4+a6ujhVd8shGLIFrW1xPrWHzPU6Mi8gU6ML700n6Mm/MN
CbYIazjv2Zw18/nUTHB/gYKjix6NikQ5evWMPppgNBTu60oUIc2nXTOsEsnEUHBSWPGFPqc+g1MI
zbYXVugq4bEjFdpG/WtpGTIJPXp3HEfcLMhwoNeB56AsoMZfWbbq63Mowu31lq88FYyutcgvfimn
xIaSlc2kY75XYqntLuup/t9S9iJqDMsNXbz//KV2ff/BuZnUvnnb7R8nNrUSE9Bkxl/fZysEImXD
bDzC3PiYTaIXfMECd5wV9c7RNSs+ku4mStwDLnB3/tDJx4ckbDkbUVTBilSSgFc+4BDPnlQ/mwTr
QRW6ajpE6bO5d8mEikJBxXWTPqWeinpv9trxR7rcSwVR+fTy+Iji1IxY1TgGyAWA8HK1tlBbwb6T
4itDPpUWi0ejk6ZiI5sc78M5Nr7NDvfutK/8wbbd5JpK6jiA4t/ynF3I0BJrnnfD4mYaNj2q8qAM
eO71A/a28Q7Ix9WXxp4/cYZ6PC8O5iM7cY8BHrkVOxXH7ivnD3e/PdnUT7ScgqNCgxYTKg8y9/rT
LC2v53BJoxUNGOXdkN79THMkpEg3ayq8o2d70g+OP8sFcgljBwVOtgd6yD9G0xd0lP2FxNYDNg3a
udAujmFINchrP0zi25Ku7iB0/FfQhta2Liud4SxglVWqioq7OdR9S+Vd1S0D1rIvOY2G2d5u35EQ
omCdeVzs3xIbKq3oh4Vfbqr7mTTpPKJ/ZFvKmVzkPWafa8qgBO+yV9D67yI+N57F7vVikQWdTcQR
xNVPrXn1r3tT9zCzi/e8Cx7GobwiLSZpktg8kDYWDgO2c4/Jo8jxlMqt9PEsOF5cwX3BXj+RpvjK
CfndiqaQGEbGvQdf3yycJNQZJvOfN2/npLQx1r1t/8ehgaTyYWDHTYOzTZULdIcCsPTFmr28z/DA
ueEfhQB4ZGZ4IyPftjAzZIQLuGn+zBOrdnfcKRM6XvYJIEUKI6wCHByz7ZZrlHMNfl0sA7lum6Ox
YQoYbyp71/WA3Y9ekPfqYucbxQgLYIps1OYPKzTvXXhOMKQj/WF9aMkKvEqnaP7Old/P3ytJBpt6
BPHQMQryIs87Xz9MiUsI7u5EFhOFv0G3w5WXULi0xSyEA92yHNXBx9DlT1/vBxIHQEmtDPi216tR
jvZdIXmRnvch7hejx7HF4jlROIZbtwu+JCJkOIzzLxQHKKCW6CBy7dv8ca5Duk9vx+UkA+losdHG
KkIb4M5TWpGmAl6skIHKV6uPj6UJ5uJxDQCns3lXByawxCZi13+H/4VA5aHjTe8DogJzJtF0GiHG
5fy3aofq1O+smC2V1fYxQYriSb3YL78py6EAwqSVhY0ne+glppwMeGesgIkWHLt8mcejjLMa6p2H
gfGrCcVdFircezpnSib7cubw/ioCnSgQquA6YUVtKr06O7e3gfje25cQ75Y1v5daGyv7UoK0nWHI
XuO3WHrhIUvU7r8mE7kwn4TEIXrwm1j6xe5/tiCPdq6EkZiP00iVt4u/GAsgdKJ1djnj9nq7hp4F
PwqJGDLxaOVGMcUYRlMFobeHq6EJuZtgtFG23Rn02AUtwVWFbMPIzJdpcWky/X46S+8+9UI/JHDG
pHpZfZKyCfPi3saMbSQVc6YGignhV1uL4a4tdBv++oZnkhp+xsHva/+IT7LVLF/ifcn/74hkXp7k
q7UitkUHZRq2bwkC2YKxbkC/WE0DpdZobgJxAr6UqwdKC/wopcLoBGvTlEDvqfPM7+MoicBvSs4B
mQGCZPCb4zYjdO21fMnpJKU6Eqc0UtqSqnpteZiUzLoC+HtKFiv+XKisBaHfEYCPmfiMMK8P30La
rUsX7uV6DC0+Rdf/1iGN+vxXFVKxyNv7hYraO5WwUzKJnNv5yo9ANHsxWDqf6teSv1KQXTf8Cmpl
EZ6V662lG8OnnaCKuVQ3eLjegUT+y7GdKnMbhim4AyqAKna4K+Q/h96SIzYHhPzkKzybrrmZSycB
uNdsofM3H3vyew1v9VTkO76OjWbHn8Q+yqz45/SCJPR1e+kPFOSMq/esSCBf8jhz54J06gfpagHx
adgtT9J9xXAd132ErhD3ZdbuHIQ4tEagt5Cy+SFbEg8/YXU4iJSUJbN0KDly/43RnzJDad6SRg5f
2dDNTJum1AmM3CBlcR2d5o4wGr4ZqKWuQH0BCSu5wZffBwKslSeimpzMvXYzqiNI3o5E1qj/Yyqw
HnCvbh7I6jKg/cexEEV4yP3at4YbcCciNTRilNIzAflHi1Z5+YWpNkjsziITZuLgUKzqUS3jim2u
OcSR+hpuFMi/G8dU1GqCt9kBPmTHD6WuJiHlTd/oaBoIRcugltU0B+DadElZqvLpPxTsbOrh7Zqk
Kq/Z94Q18tFBGCaBBwqkY4dh+kt0Y6usgfongM0f/Lwh8yN+pCcWLu5t1T+K+oF5Wc3OonfBCSgA
WWSdQ5PbVlVl6cazJfHTVNwWUfb2scKHKUgrGZIKs5WIqLqiHqlWN0AWmgBj5+UAT8zwxt5w98VB
7IJg2FPSIEcIFxmJBQJCt9KuidxVlLZB1VHRUSEF44PQgiz7pcBxvE9+nENssaJdhoF6zoNFA0L0
S6RaWiKO5IiYV0cyuj2/dkx+4h+COYpXTvcK2rtAoRcSPsoG94y1nFNBmrQ2aE9noLRq6RzAtVwv
+VbB6CdXUGPudAj0LfmjJej15zi+dFgMhnfEZMIcs60BtEQ78/8i+2YShXAdkiLfs1sl95DeAbFk
sw7uIQimYIXWsKS1YtyjoXa9iaaOsIlES+6tNlJTBRXWDjhzUbyIGIHASV7TPOZ+TLEEIqjPd3Ea
6OCTs/qo91hnph+ds6DO/Rgnt6BTAUt9qMz4gzRw0s5TMrgO49pFUkNd6H1/1a2mUzfY4Xz/LpS5
NZB87lk5WiA1Icj2PrpPEXUfwKXcNuF8M4pWrQ9jjBW68KLS5zr8fHNMveFKBEcnbGqJ1HBHnIzt
EV2PrU9WN27yolGOi3BgY2chuls6HBaTr1sXmIQthxeiB7NOniwMxGhI37hDLBApOhyqDa4BWznK
j/6mM96ic4Ulr6W+GeYHQPwKDmFtBM3Ffp1/DxFKnUwKiZ3BIMMBwF1hGXXzMNddmnEpFVCMrO3K
szbbyudMvW5vBZpByW+u2R/J/nZbJ+QfrldDa02Q7D3Gt/4trFEKdWEbQhdotIiGrq8KL/vQ8ovB
5y3l+zt37vNE7yBIIw0TQY6N1xHzpyVJ6dxZ84PXpuWg1mfZM8Sijgu85oiMRtvbbIbyM9JBQ3d6
iRDRZxpg3ZzPyziEhksjue4izDAYsNr9ZZBdnp+Da06I3T5rrA11js1Pu5bIS0mcl87ujUL9y0eY
xEztHt1QsJe4/VGiXm9NvsEV09dPtjhtObGL2BYCe4M+fSwpXMUvlcYU3DEeGINzlHaIvUl8Lb3P
DYi8nxUAof2mMqoUsLmoBt2LQom28MB9ISd1t5EEVxS4tuNIbxZD4QXIimtqMO8Dtje7oolT5hJm
IE8ZzjOnSX7dgBD+TFQkL4v2PNyAyU81/lfj3dsUJhpl5F4XuXrrRnOFn5XFPivBsGrKXjc9ZeCR
KYau+JMHwM8pjZduwuoFtQ83uJ1zsYDAPkZXnn6t7ODiNRcqZJPFZHQ0I4kQ4T3SvX6Nt9Z/HCLa
0Pzy6+NZ0Qa+hX2ONrYsEn0urqpc+vSfQyAcMjVDy/HkVZTODNuF5ha22ODkMEKCZrAMBOp+tkb1
cV3fgZk=
`protect end_protected
