--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Xy3ZBCadKTfC2i2NSxLmkQF2vyvVWVRDNXjQcBurixwq8Smw/bipmW3Z4jgd2yu1uM7jd7/zdsnp
m+ElcFoI2Gh5bzQp6nkCdp/JA9bX+PX5Rq0ANWieOspBMYvcq8K+Rw0ZXJSHO6zeHLV2UWaUnmUg
4eHxeCQIczigvSPA+Cjs1TxvLBCv74ok1YFV1zJWBQYTPj4ehiZZz64CigrA8LEsJQ/YqAw1sPvX
JRqt21cO6xXa0aqtLCOk+/JZ1EO+JNiKXiMvUPQXSgIrIBWw6ceaUmLhHtwRnUcaYtPupC7duc4B
mClBA6G8gIcFrl2tG5dsfrhbWxpT+L9k87BT4A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="o87AqlsMP1b7MmgpQwNCFp236El7iOgArbdjs4Pu8iM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
PX1NMb05auFdvWiN/hdE8DYYG8V78yfDllrpd2R8KLkij/yRFeGAVp27PkPXStapQ0UwH2PPjOMn
gizndLuSBp6t7/6T9+SVA43Gw2d6+r1d4nYzd64CS3ppnziQE/UU44d5N6s9LmDtDa2vKeXq9SpG
xCG05+xXaIX9s05YCFI/x5Zv5lsdVsoYvRxmz5ZNBfydbC5O/hxR9iBz9Wa43Iy41onHfi7xg4Sa
UeJyOA+Fh2128s3FfWqi2hM0jmAOK0Vu9QsP1fU2i6mcvUA74cFWhUrssxlQmrmS7vif3dJ7TucB
0Kf2UqS9S83mVbqukSFnHjHy9Gh8HCgNtgOJfg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="DyDsTL2OGxeeJc+R4WsPmRK+h+1woPcelAw+gZEb18g="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22064)
`protect data_block
md8eePcWWv3aJ+qPvybRei2stPenXXFz/CcZGC1wU+H+vH8nG0LvCzFkm5Qvay8PBXwipftNmX5p
aUu4I6vOkcZfIyypQ4dMp2rpR/29FTeislFafOB2x++KYr2D/FEMcjy6c4R6yCQp5iFaFzEEaV6z
rSy/JXUY9ZagM/ohj0X2CoQ2xlj5iFjsJ1a7Jb1sDVZ5gSGaUYf8DcjG15K4TnuZrCKYkqP42m2K
byvoynTM+lTS+T4CkBNy1LS94xvngFWldmZJdioEWV52KGONX9dN5/haLG0GTY655q8oagjJSygN
n135/J47yqh1VwVdMaf8SVy0u30vxoDp0caRh5n8K8lSRmNwtq95+QlkhHKIsIy3a+7fJoK2DmRo
AFc0atElumBsNV7pVo3cTwNrFTfMmTWMC+9coGZraVSmerCggLTsXruy9XiI7BE9it4qM1cLCQ/M
Z/5HUs4kwudagabqizfPti4qRsFDQc9gsXIt4QZ/ziZAbbQIy3orK2GqpjhvoselIwFgrLlaF/aE
sAuEL0Je/LsucFvv0dZbg27Z4ypEtNJRFHuo7JBexSHRtgD4sHtdM5eLwM76HHECnH6Flvlglbk3
H8UKZMeHV5YVbI5sYIun7c/qSuFxvbiQtQIhaGUqwg+tjTuaW8ZSF9eqQUlHdLCsHEYtPv2pPaBm
q8+qQ/RE1quw3u8p8i8+Jkq6x3sKLWFdILQ4GhxGzatlZZa6itLpqetH2/6cf34L4fuQTIIQh1bi
wwFnwk3cWY8mQAAyCu0FkVj8jWlNjePMhEsNvILcSz1tZmDchZjLSpUm4iiDo8yQvNDg69rBfTKK
UpyUSGktDELHZVWzML2IsWWuyA7F8kXvOZTIvGeLAgU+Bl2hsdJOy5LKTHnpEWW7GLmdast+phgb
Rejc19f1V/L0jjfL0So/4ZGO1A/ds6GTqowESTUzmABi6zIcOpdVj6Y17KTs3nSY6nQ8WdCI24B5
j0i2/uAlKj3ykwfEhp3R0MVvdBQJNqlGQGyEfAqSGg3KoEpSZdnh5IT3EF1lDbnxuDYoISXk4TdB
5VvSisnHGjaFPMmSoiiHciCPCXx0as11i2E21s5mhhu8lx39/XNtAVEV2+ftzlVkCtLwOv2Tuhte
d5E8qLhbLXms5/gopJ4AdX8oxJb8RMU2eTGJMJjwsgISYQ/5ffxbZk43bI4MnxFVaUbMSCwzzO3b
fhmp/Kf7Efa2lHxgTuTq5hIr1c9zubzEUAcTvUkI/1WBJdhsoOjXNBKBYLWVsSKeIhWM8iU55f2u
O5xbUhhEECstMaH6yN5kjsXLXmu29uzz2kpDh/PpTCI+0x9jkj7qQiZVLu1Ao1b1Rv+dVni4ea8X
N0YVKVpYnM3p/0nHgJS0M4EjymaErWa4vGaOJ8Y5bvumBWm9EQLQXv3lnFFAbq/zVyxHboGh+mbz
VLTALE9XBYOdHikgQgteFTNs+Q1qm/vY0xhRVzOOZFODjnuVZzLm7Y9Inabe4Svh6swDixyTiZld
mvii2zU2EAiP6g75c4GSqLVqouI/gcZzfHLN8JetA7PQgagAPPL8vLUgNYja0brHUKLiO1XvKLh9
GMkIEYuOpp/jbJHPjab49izJyzsb1lu0MDYQ1w0Uv5UY+Ut2uHvuNF1NMbgafS9Muov4dckAhEww
ISYARHXsqBC6PSxpe31KEsjR9zzvLx5Xp2l2nhPFEn815Fdn87cPL3mL6zOo7k2Exw36F68JWWAG
il8FlX9opPf3NT4fThlKLbgEQMn47B/jsBaBtzwqwIdpFwwQB5i7SHhctKPpkHItunZtEdAUcsEz
Mh9JTImELwEv1LVs16YDXSfJ1CuMyizo6yfYiM6g3fp3WRLuiZNtXAYnjf3Y9920qmZvI0596z6W
LZa+/pxrn1CNr1LICi/XL0E2pYO1QxLvG6atr4N/IAdM85c/72JVKCKiG4vmq8asXtgI5sPWFjsQ
kA7qmZvXzBbP0JeqrS+kwDB0hnkDBNGZQ4hKTC2TEGQGstgO36tsSqCFVNtUjHoZq8bWoUXslj0r
LWuf/w3WxKLycWeflDsnZJEKzOv9yZmmaHc9L77kvFuH9Gaj5MPQR8Gi6KykHHeKqdpgfV4wMUjv
KwdIBDRkn8GCKgcRmB9AwE+VpMg5uxjAtwh4/thD89EpdQTs8UgNOWqiqsiLpv007dtmkjlZHmtw
P67sTMcNPWnvTYpawZsZg5DsGH/IqfxoGYKxX/308KaTvAvMyoVA+sLOHnHnGX2AdajiZZ3TLA/c
pEKrsvL9srCGl82XLLQ3rL4lx0RhyK0Yv+Jk35u+Ub/lI0rLyQQ6U7J4U19emILrG2M0hMi8uOoj
kaEzSb/5C612hoeqlll6OBbj/K7QCOWIuP5ZzHs991uKuoEXs662t9OE5qoURclzT5faZhMwZpmk
oVMyncMoEIYkJz+vdxwEbj3g3OEI05YmkGzFRpCw62qZeJpDyXRvYi4wE1LyRkdrUmWB8qIDOJxV
qSIp+/KqmW4nMhzNsF8ubv/AwXvNhIN+LUGRzMgz1ltS99eap/LnTpNPY2nM2DmnX/VKbfPOl65R
4wJST0tnqdHlB/zNeRyme6gcUtfbu2+zzmvYgyoNmEl2pEJD/21joRZd2MnosuYoHQDFv5fYRmv6
aYbXXhZl5OIBUDwj9agUdyw9adMRE5M/Csd8Es78VBOJX4AKjWMt8myTd1iSLbiCh0eo0OGKsMC8
AeRS5i6Gzz00puw+jl3uZaHED9/J7XhDeIyrYr6P4vzBjWiAb+pkhD5sWE5ubES13wZEoFQ1EoLb
wmpnU/XQs7Tg77Hkm94YmEA/4BfpEjVhhbfZvZ2dfhAv1wm8ZaqeF4nhRZ8DgaPsGGJ48on6lwG0
0MycJMEF65zomj/p7SzcjYgDsciBndhKOHWys6Ezm1WXjn+X+q8Z6yqawXN6kP2slxrxdCo8mI3r
+xR/d3ui/ehVgZYVwqsc24omLvAEOPFEGBaRi64jwFvnnxH0K4i3ZorZCxVwiy9dLpeiy+F5ySTC
uw4U7zbv1FA+MCLpyz0FpD4YzoxOs8feegwmZS/gFmT7s/T4b4pAlzh+xcdjlQH4XHIRtYnzMNL+
iuRPKegC2jW4HzP2Hs/XxGvnuPAsmoCoJrc5yXvnVKtentb6xnLLNjmkvEyFlqv+m7nvXMhz83U3
ap6WJ8QK1JpAO5mXBQ9IL58PWO2suhq+iVBO8yO3/3iZ3EDXecIO2aZ4z+hCzf8pcL5g8HK3TBpu
yDebaIVUIl8GKzAMcL0WfTioaT6VkqsYca9Za3iofBcmhI31OThx5duv2XvLlgnLzYoDs2U5wIA7
sSNqH7ZfXuUzRtp6TnOtbo+FhbdSM9oQOI+Y+fxhnULBqbPK1FB+oX1AM85i9zx9lB2bRoGaq/B/
xBIEdHUSK640KHXmP7azoEwO4ny/mCvUXwyXYDsmCq6WcEthb/6Do3b+iZcUs2b5Wk3fpRBAhKQ2
HLpGBRr+9RHQ3W4XUOGvtCJVvGNTUJFznwufefEVKt9R832NuONAdRY8NGMdyJZtO3vOI56YQs3h
Cqi5cGx6PUP6RIt2AIXqIwQiiAoY/HaN/Wtd+aTDlWxuil41YTm5w9Bx8Vdno8cQY71D3MPjrphD
MaleAKo3A6fL2QD5H3s6YsCqfGCrLPCvOhfcK8ISF8PkycDwPxjRnGsPgo+vNJsKGWiUB+Mjnx+E
BfdQLmWgrUHGFFWQlDRYeApReWQhmAa6cEpompOeviL+eo3zOlinALHSa2718W4r1FKGpHUy8sDx
hTt8VXsMgJL7hWgDlgkWpFqAbYP9VX4VkZlME7ynmjcqgvpgnTxcWyECCRLRH+zxf5+co2v0FsSW
+cwl4sIt3/djPXLUdH1d6a1YQM0KeXgef5ja4bRWoxXuCB5HCyNuod6NIlo2oULuSJ6+763mUz/4
o2Fq1easGRrHxdq0I6eNUJktjDfwshMzs5JwKxswv5onft/VPmPYFw5g4QnWizZsvzPGC8YwmGBr
2wY0cjsZUSXBH8rh5ObPU3oCkfTY4BIdznCrGpUXrdIHtrpBLk15om+QO/HM36IwMUJOaTlZreRp
71KSwmSy10RVNR+SgGt31+ZX7HhkfqxU4FIgHKXtsgyrLmcBGWbBIYQigASejBPR1GvUQ0OnFt1L
mp73Q9QlvYbE6cxm2Inf5GOni8jNpT4Tx/wN8hAwIAG7PO563OGCFM82049mOuYmRcMAAyryNfTg
gA6ULtHwIzPh7AHGvSoSogedJuJD01fW5HCp/UTSqaHjtFsYfOpSGdlfwfTG+aWngcb1dOwaHVs5
WLN4RdP3WIictygWeQw6qeAKnremuDd2ZkLhrP8I/z5XM6x7WgeeM6uqC2LzbT1BCpA9YFNZ1lNT
Zdh/fg3i75wbxONCEhNnKH1ea5p75TvfRhYPOGrmKxqicOpZPcxsYcdC7V8ECPqWxyzT3uO3VhCZ
RYfYL2PR+qQx0PNr1lipnmwAY9eT2eSPfJVV6uRO4NhCwAVKxwbNToAfcM1LtYm4ByUnsrOmtdCQ
1NGKy34U8znJGFkmfOwJA5Oy4pAmsLqRlXfOyeG8MebDszOrY3ap0uN+vVE401IKc/fouL72BdsE
Xt6KuN4QYKJlWCjlTY1Svz+5Q1Zdp1nCSz01x/Mrg643OMHwUbZnuoKIQPxTvgc1AmNkGS8y31GY
z97WfBlZN/kAKI8tyNey+9JPWgNzXp8l8mwUp/V8UxyuwBRrTaVwN3BnLEGdDUla4Marswd/y2c0
k9TcTmauiU59FGLZI0vF7yTyX1cevoSfPuVaoR87zrgubZsoIfoqslCTRIcTx6gf5URYyB2mSPFb
wRBItM6iq7PLMQ6nR/3ViUhVxhplUFgmNkT7ekcqL3Dk+rWvTiQ0tTikw74++WLxwBS5MiiFOsD5
wL1kVXw67oxqlxVwY8xc6D8AhW/FeegYP15vwtIUKOe0rIjZgVlo5A3Aj/yWIpvqN8Zkww0Q/BV+
F5ePtBbrasfrJ6fXuW3mU3+LT3XiCla9a1pMYLTTd4feH/wPsoSNDnGkWKYTI6Jm4wlojTSP8XF0
kM4LCq1k/5p4U99qsdbDF6VuMAGHfVkE5xNF9c0gd7i+f9qGx1Y1on7+4OQvfsSRcW5AVIOmj+cm
hPdZylo8M79kFDO3R018PqiHrlNjCly2ZxsOug40e3a6j8mkZjBkAsIm2jnklwfi6gG/czBuM1WN
8jnbd7tim8mDsDVA+1kK9sZCiHOji9lt+r64bf1O6tKGJuWX3e0FxaxAwPRlUBPZSskXfq317Xgl
3RUGg0DbuZ1sq44iFC8H/MjIp4tAwO8ec4nSHRXCJiAwOeMu/o68veon19WFj8IHfYHy2ripOjVg
/ETEJWq+Yg2o6FzjsJhgb479eIo8upNnd15SKos7dFPfAMMaiVbOkzHmafbC1sE3kb6sADdXWTUx
y3DqwdONjZVU1MG5oJuzu+vSgBre98dzHVjCHe7udWR/hNfElbjOkvDSHrQrNeeR30x21l1y3ktN
25tVB1Q66PMqtmmn4TbXXGXlHc8d5KHNTOZNL5RBriF3S7V1Sn9ZricRe5+96wMqgBB8/2rKvbjq
nH9ERweCKXE+xGwUiNXLllZGuW7iMrcnNAz13zfz0XC/WTFnxezGwzUQovZiGznPrYEjKuDm0b9/
SU8FFjv+gaRyOX6WT1O1jC5MGwQvWIIVJyweRa/HNTGh5eSu0f196aXF49gWEBb/mYWFi0wTfOHd
5Vq2mpeSPW/TiD6V1MZkAftBKtfvmyepfOgByURKEIUML6AyaKlHkgPBPC7dI1jTepfJXCYiwQOh
ElbFA3QSCmxoFJQEeydEH0tEMFznaOMUF7yUVJ/zTXjrFYm7zsz1eV9TWqv+pY8Jv4vK1etKD7OT
osOquA8vIvOMamLFaK0GvvtDFWmX0RmCRTLUK1axBc+YvMdGUQM5KXtbuChwN0zWKIOKz2Q1t2K+
aECMfiy+nUSClffc7uVbSeHSlVzkzvL+n36tzSE8ElDVbcF8XM0EK2pMqm6SiXodJLhn8PUcWPNW
a3QeoaU2yscLpW/BSOgGCO0IqFR5J+khtchv2LdGEsSt1i1qfG8gqvkiJZ2ULQmKvEKJltupQxxh
oGzdzsR9q5fXrv/It2WvutUYEZy4fG/kiIcoYl5w55oz3XwnCj1v0lBZwMemOxNHeQSNfga6f7Um
C4NdDiz6bXGkAudgesgaIKTLDdgxgFT3HweSU5ucm7wQ3KhS4MdI3V5IHZnQFlXSS5JnB/Yqqjx2
UvS3qUF+fUunhvPFYFcOfkbHPfxuZgIPk5avURagXiM2Q3NpcQVAysF+fxTleCi+yqizqi4GrfrH
2l3F3Au/BBbZnVoxxTLH+NIv0JD4l2IZEnGbUys04WlyUS1L++oPENjIEaBDMk0qnypMHWPY7qCW
mKmLbPkjspuhIdwURekH6lwkFTjC329V4BoyoBtlqgaZGFVbQkl8gSR7EIxJzIDQgk1kXjThvt5O
dKW9qB/5yocH3Te03pCLZwsaJf+hK1HwgWwsIpKqCJPH0kR79PhBqnt47EnrFXtEf9wPFJhagSXZ
Dy3otDGjSvV3CLD0XL1e6eW+wv246cp8NXF5nQdDHzyS76xDWj6rekPgFGRRznSUd2sESFfK1ult
BG+MtUT6NPp01xPWBLVTyCZjm3e8n+jbUO+W0MwIcq+uyBv42eERJ3T8i4Vj+a1t+GmGDm8WnKNm
U2S8J3SdAiLqleGdc3nPoFV+YGKdbRQlL5KepUuTD2+/fHrMRuWImaJnwlxOCmVfqjdBzfgy55Lj
j1pnYVccjGNQCDB9kLj/AdxyVTXulrOsEIhJXuJYQlkVNDuXcVWnT6cmwo5PxB8MY4vPlBhH0YX+
k1BZKR9SRHUclrgfs6dbTtg/RIj9+FQTedvjbj63csOVvdFJfxbdyj4J5Y3BsRT9h2tVkga1mUcl
nG2q2jwGRy1tL5aZRP6HM+iuvDS/XeVrF3hX0AYzrEw92b8+Z/mQB83cbenTzkHg5k9+oPeQnFlv
LzpjOk4qCpe3LgSeoyfltIjiYZwLMOuGHP7MzjMYHvL7WkRQSiH1RKeapBlu0IHpManU41tnZeRK
6/Rqq78yL/4ydBRc78W9FJhfKJ64yJvxsiI1gKwwK3zuhj88E5M8GvRUACjzn7A7KqootKo0eM/7
02+UCYEsxjZPN9pPyLOBSaAeSE7q6ottvojt29JVVtxjjjeCc6Go13RsmraHOobLU3vlZHUjkeE7
MwIWU4+xnQ2EJ/PE6d7nDDQMx2lc+4vsdKURBwStMIo9HLdBbn6mZRRk0LKCHKeWUWm1e0hqMP2U
BySSfdMWuIipR/pUhIoxO2hrs4nuuAPkEaxChtjmCXylLG1NBuBENXaF7MKrrI6Yi1yBeyaWu5X6
MoQUc80YS8N+0ztq3Uy7c8zxyCtyIQbg/oimGqraIChGhmhLD5npIA051Hx7aAMIDzH0YWCH06xa
Kl9y5CbDg0oynAwrHyduJ3mo+tAT3Htc265JNPYeweWubMDigb07ey7lW9mgwx33fgcHEvVoh6qs
qxYFwr2fKSBLCjyZjRFuhL1cdWMFd0UsMHtL2Vmyi5N7I87Ye0QBfJa6tqotRsHo/FHCzDND3aPP
2401wuP6nL0rW9ejuTMR63CepMtwMAtGEAxQUoO6nSHXBiW1vz57Ctm1MUQzUEu91Ioo0t2jrW0Y
EKfE8QL8+xOrsbmYgbGQOz0NHW1hZRZMQiUCQ8zKaeVrh+Bj6aCZ4fQ6r4DDZ4Zj7DbBuzt3iE21
SyGdAqNNWznHxQk/we+NebLBI/bOFGra1Y/gkv23JZt/LI0WcTzYg/f4te5XJQRFgYTFF6cSPkTh
oZo4K1OP6RQ9P2+JFzezZAgKum3MLOgIGcBu4noKyvHCr23LZoYR/B5gj0vug88hL3AiBzlM6luG
0cD1HWTFNEW54DkiE63/rYIc3NJ3NTnIBkEYvNvwSb6B9r3r/BR+0vYdL9jKtVjgJHKyDVgdqC0J
slSQE0iRfenG/nld6o2p2GQefvPpSTwjvVuhMBDmrfXrtufNG3Te60r+gHK8Ml5ChA4vy68TFpvd
YsEWZ74Mfl31+uzPgf7Kl82+H0I7WwCEGvWSWdVNDdoZaLJQxy9p+13LCZju1MsZMEKKtfkM0BHO
Xc6B4dwfM8Ur4i0FPgJmgAFje0FUbc5hjPKq5qpf98vQmC3pLQjoDzqPTw6bTBOXfZZ0KmOso0gM
ipNfyNTF6IfIhi0h7ifYIdvBGPsTNDxk+AaaoaqzlOhmtodVzVXXPl7JhU9n1HAoh0bPKG6hNh9q
/GJ6VRE3BBiGghPTZd2FMfx/TegF98JV2RnIz8PqJjoMwVaPXx4u4c45DI7ZwcAIcATOEYG6gfBK
WXOT85Ch86pF2kTpMfGFKfPUOy9rUQ8DyBhibinfdcUtb8/Jut2g5Tvjt6ys8WC5E+Pe1KmORIOC
YVSx3vBQzd6QpZSAWmHNRiXZjR1WjQr7rDGK9OqvZmrR5+Fnf09cknSWB0GQi14noeQJQB5ofTEV
uETFphQp00Q1bUrLdtTWZ41EmyXplc/Y2CoWHXNtYZhG3VpLwW1J1jPx1iHUPKCxIK87wgzToy5t
VIoLCf7MVmy/dU1V69XIbqotDFTjnFkCwGJ4/wUAvhjibjsHun+i9e+TAIS+jipeAnqWK22sI1N1
Er4q6kRjFDAyZyzv99w9PtcoQ6sej6QA1j5Eh+YQ91MufKvzwjAGPDt/Gt1zyoBtSXS+Kgi0w2wi
EE/H+wSg/eXwhefApXoy7BbfCOzQQiAfM9n2/vtXGaqYQ82xu0cHLOeGnVfH76j0it/KoxjEQJ9+
4QKfqVWraUHN/TgZ0hDnOY+c+Ahh+REDlvqI9SOuFXCng/NRiFxM7+qYCw4vVWeuN6LAoV/K0g2q
1mtVjbWr7erbjMIGoH/EVhgZIq1E1tpuuPg2AcvywmeBMuQvtnDDKXZkhtgnQV+sr17tGC6HBCrm
yBffXMss0aRNYURmbAVw5wjOPLiFeNNp7rLfs9cGtl5cAihEaI1qw+p2zj6GfgxcLP/gLNhrUgDs
aa8kJAOq5eBsOeYr6s/DRkY70gV3eZNxuiOnjMTqEtSX90vqZ8K0ISNaqIRWx8Mpl3LxWZ38Kl5o
E/mkM8kEIhLX+k+iidfLHIk1azhDHFwWeZ8GTv32pGfXrcscGM6wW0AqzpUQd88fo2yTzyBr/3Lo
wnxZYicsXsYozCbfemXDoaQsju5lN/Q40eVgeMgORnJANhjLVc/gT2aMnY5z+CY6QvRDcZnzOM+3
VK+sEKhSRqbBB7nYnGlyqwlOMefHnC8X8F1eHODHSEgsx/x6kALH1BMt4AT9jJIJlb1MLJ/YGdNo
sx1n1wXn/TnzmQgPQBDKcKs0gz6sOlTn1k33omzyy5fuoVpgxnqpT4uY6HPO/64z8U4+psei9xZG
xTXtOdkFK9gUhR9cH1bfrjgoM3zEM6oUp11SG7GHC67sTiu5Sn2q3/piswhLtvSb0vXXvr8hhNjJ
EvbRM8ItJB0FXSFbDqGsrUoustNaSpiJHEJK9N+wVgIQMce8LiBGumT1LkZHYqTGCgcSg/VNtI9E
4gpJDgJmm22538LB19GFro4IdaCN31pI2RtZ6MLznYvO9aB4RTOkPqVO8tWNPpD9dCdypQtkvumo
z+cmuk605qmgO3rGB98Ng4BDTKJGqDMAYFiDQgqfKIPww0u93bl3pw77UQH0tYgNQWZoK2LGgYuh
xpTnTo2DjTewF9hfHDfuSR77kUjJGQKf0o087qknxJI5PTCYLEgp2jBOxTeRkZnXGdmFGcCo7PGb
SUeHDq5ikpWBVJrqb542Wr44Em7TkjUe0fD+kcivN/nCODec5LffW+SprMDYRfng0cUL+ViHYBDe
m/XG4+9T/8CxVoFxyjxHpB5wUfsunaNcdSzwZBcdy8PEpr7zQonUzPfKUewxGuBRqvV1Ati2RRkl
Y6R/wnV/XT4x0kSKTQtGwaBy1ypP8Ffixz7wjVNrn3I9TRF0LWfYFEwgcbEk9jOTyaRoXKBWXzKZ
SNj5oUqbOYFewt77OVXNO/urUH4L+zV7AkeMZ53nTUlFN2yb7v2cnabY9tDYUx5lEYnk8hXcA0D9
c2Ma+vI2kPC2CJRiFzgBwXpTu4bgwqr4x32YTvgAHHLpsc7/YTWS/wykCgL4l5UmC7uasj/fVG97
zsSbYA8AYu524pwu8Pv4RX7Kc8uAHTjiSIeawTvSZnqbBw9U4m7YpYAFHuIi4bvG6AVc88SMZvKP
ojmrV+cwjRlNfP2aOSGd6r+re4uNoY061IlIXuuKOo02oAX3mHCUKPJhc2tvKXnuBg8rjW8xX2BF
FgbzPEiMM7ZKF68CwgEPECG7YlPiJRO7hkH6B8+XsN2IBXe3Q3edTOQJIJJSTdVYudrBA3C2Ct6r
VQQHYDn5y21P+ycSwV8V2YfPhDdHRCKOpFz86p2yHgpbMweF2y/yDY6tMRIqDVxWbLupyGTu9JIf
hD7M9+vPEEBw6XoF0rOMZPb7TfXfPTR23tJgEjD2TCwmluR8AK8ZvbKzlAk2UAT/cvHl7mIjaaRW
yo3nrvk/fWh6FOJszK6EBnaxZkuH4doJKb43m35Wh3gib0PdT05qc1FaRNBuzakyY8h7P450kWuM
AauiT4pFhkQvUAXEx5r48rRfpimYzhPNKXz08rdUq4TaVHwJGpYmtIde9yywgzqUNg97o14nla8x
iBfonLFn+/hRnoJOA4EVAvxA81axhrbn7og/KQ/m38+SfMEEHppgpAQWyp7JVigbY0whAW5uqwje
BtqgJ85FWIFLHj1bfNZtIb3TE3YRAN47WGE4MdPZEHgLekACs5AAibYShJK4lRUO6G054goRCj/7
1AyI2PxSZG2s8F/tt0/Kr/PmygUThKZq5RpcuDq782xRw2zeKS6S343rzJ0f8PCXQYdkKVoGH3uh
WJKcZcAA42vd0Adq3sM31g3Eo6/OqbAneqm5J2VaCjmojRttWp7f7jFSFo5rmXdCEpjv9bPrLpzj
aIN4oQiWZGS9D2zjQgWvPU8Yvl99eQ4vQBSYbDFqpqgvfVLQz79Q3xbH+FE/y20mb+yeTCLWW+Uf
4oq5/X1yfInpBq4d4pIF9EKdv0BipUafEBgszBiwFLyoQ3Lki2UaJhwjCve2yoleoM8N6qDwthHw
e5qCnNDyYh6WcBqqZwBtrxmzO/H/KewE/9QUPj37TfawLbc1HOGlGYty1iO9xsIyLQHctmBXTJbe
vGvJrjyA3N9AtpTkFv91BrQd4Xx4R33+7VQPCzWn+ccMsgUotwpUV04BbG4slWfUjtjgGMFUBFgH
qTj5/CL45rO4+ILmify5SQ+uJILZTmgxX8l5R/TuEZ9PJPGdCnGvmckLaDlJ7xMjcXOJwmWYdTuI
JlVThT0XVoZQzJ04pQUDmQilxgSjsi9z4R+G1xgXVgBzh5s9rf0z5IshR/Ybc+bVNoq1i7QkiaOR
hBqy0jJytwpvUq81nJjffUDr2FJXhyqW/6VXlo/APdqjqO5HsYTF1ebEot1qdSOknJK2hh2+giyZ
Lge230r17cWvRNc7QJaYMGk4bGuu517dp8ghXDmXH8fZYK9UvUPQq00NuWKarZwwDHz2FHv1Kjv0
k1FVfBVSfTlXYKg+U4u0H9B4Z9bGtCs2R9T1yh7LZer8jHYQTj93yjq74L4OagsNmhNABux2ponA
1s9Ac7AefHLTlnlpxLA0Apzl7MgJHRNWaA1huMSsZfSQEfLuPup14oSQRCfkYivo5Fk7j6rvXjIG
UrcAPFizAhAy8MDz5CdVKivTLIDWPxEvlMHQO9IIijQF/u9cm9mjEQizlaPUzDeiPisvhdjvZes0
VaOsshgH8zLijR/+tXQjJ2QEmUkbVFI7/EvCKIIf7BPsZYi4eoFmOQmpC+24e7NesTWHR8wrsqzn
G3ttzfLObTFwge8GANBUrR/eQlIJWlpINYyhy4dt3WwJjTtFlUCzDUCw5XQVk8kDpSyd4OEXDs1F
/FzNRYVN0ZE1noMYVdboUn2M4hitFqbKOGhLxPDC8sEI9Rs6yEYW61GYWWnXjSIQ+R/ui8o+JAAo
Biwi+226TeJ10WKokLhO+ZT9DyVygEElntFjqf/e55moYDjtaEr8ob1WskBWPcuLJ5INvi2GIQUR
Ah0USXS+GX/QGe09RP5vwJL07ATZ8jrJKvKjSpPO1ApcNuGqvG8z2Ve4OYqCsWw/9Gb99bg3saOM
QvoAX0QFapxPHJf7QgF7FFhooq5SgzJ3FZsv4QUtRAm3Xgq0YDXENQnEr+eRSMVbEXjUato3KcI5
UHgT44NGH0h8JedjUNtNB7mte4ZFEaxKbBdyWAQHC8kUveaLYvifUNzgrR/O4xjUtwEzyk5zj5x5
x+SJ4dbEORuzP2aev1PtYm4wHnmQRsUI082I1hQI3iPNefJF5rEyqP9vOO1gicZfec5gOP1jOTLG
Ein/LZGL+krUgkdI45iTMX5Yn9XJnU2Gv6Mk0sXmkknnFlxDtO+hKFjzy6dB8pQTr+UEtzFyKcbj
EaKeAI5ovx+MFEADNtDbmFDb7JMj+eXThNrLzknBbHb36rPZi/m1m/hPAtqkfYLRVUKhjP5BA8ai
Q+PkoMfX89i6Xftl/D3gJXKAmgKshJlbfLjouizEBX5p/0xJHDMhhNlJ8EC7gZsqtFwdyEmFmbbr
4ntLhDnxtk5lggaqgGvJp31obLlZcyyVOYfhYhi9bL1qlQagBGQkxjyt5bUjakT9Zxycbq7vxi/2
DZnfwcr7/z5tLE+FW4IyB4ze5op/OI7Q1FEirhATfAcXTmGcsPhJCPH44wh3g6wyMyZVD6B7OwJI
WT/YatPPlJOK511Sv729laQGRatSMAcfNyf1O/VRNbRpspaLGkXSPySs8NrXtlVMB5o4bjVj1Z/M
qwd8DiGmWBNIngo2W/U7nOrrsGd+tuA165sarsx0YgQM93/DsxA9xbS4+MUH5pU+VuFGPGZYOwzY
FIIrNxso8Sl8Z7fZ9DVen75gUqtE09sCW52zxx3GVJqOXH+KAusOpC6s/O3Us2DH987M3SY9Bkjn
QrhMfodq6kChK5tqks9CG4TwP+tEdUnFoRhDkEot3YWv9eIuhOjveISdSNk0klYEV1swZQzX75ly
ypB55VGtewNuoVDA6dy7mgHnCKzKR1LqJpiz+yPHaC4rB21Aa/a08VgAlNsdD8sT5Cf0KPCuoHho
VF/H4XdrM5fF5ldgIu3ObRuxF/wMHQVb4Q5Sqb0REAl2tmnZjVVzQBuK0QNpxXiKir7YcoIMkVHe
m7Dfhkvq5g/6Wt7AgPvRkAfSfOKI/FmbLpw4Ezt+oWyp3WsR4dJMdYkxAfFLj0djyeRcvtUi5HzD
5N7vrevsFA9pKUABDqU9U2+bvjqUJrsghJQdogZgesxoIyviI4la3DK/PzynXF/2HeNVFpFQ0P65
V6rJB7FihP/v8O+av2mjC63FIpJ++wj31U/bnwXCs0GU/rK4gysvdb0MhwdmFVVVZuWFNZ4pCYi7
k4BfWo4UCN7sQV5sTUestxnsCWeow0iYfygaPWGe9ocNYqgj41o1WZt3KV6f5qYcbbMUdo4Dzrwr
1kewEq39b7p54ZcfafQcYal2Xo5DIJv75T9yMVT+ywghWAW69Rl1s4ew7jGSu18xVCIctSdMoKJ8
7Wp1GvVFP5WNCThCQGOA7Yp5HR8MCpr0ZRIrO7FVrJnPTpjKLynzsn/oVWHlYdwIdkjctzpe+F6O
IWZpSB+bvOZihPzlCmm9jUI/AqkWAQazAzPIN+Durp8wqumBqeLfhwMG14rhAFQ/PjXXoTwemREK
D+KR777zTsV3MTXZ1IE16C7gL17ugD2PX5bHkDb3yoeqh8EOrThi1NhJOgdIdLBeV28DKvkdvtjp
2k/k7uCROcYYxCxlnih+8NfouOokztF9vBTQ11dWGFxZGXRyo43FO82qi2xZQJVYVHBKngXfbAbL
bisf8A0l/wfJwYgocO3qSTicWv7Gi36EdG00e6VJmMTOX7KqvAgDXwYieLszIei3xWQi+eEaW+RV
mvmCyF41CE3aTH0FbNKHXTFFIBEpFSR7Ap0RRYyGnQFUlh6OckEDOzY4wljtsU7PffZMPY2ebUk0
cewitiHPMACG1x7qqMWtiN5CHXWzNMmZ3jiAXnsIFHAwZ6gZgPKR7KsdFjYSaMtf3b7VuZbmuFOR
zIIBLlXOhflEUoArV98QzhYx64OL0c3iTzRKge5OoQbBgiyI2m0DSXUOiQw0WMFfU7Q0DG/Qj+9O
B8zgMTKkVEwIGkRTJTyUNge19VqKxMymdUk4A/3KiEtDKCUM8ixmwR5ib+6foZF2Gn3cK2Q2B6bR
c8JZ3ezAP9s3JI8097rspCmLnzVjbKZHf29nLaKQ6aNrqTjPFbv0iU772XnwR5D5VB2DB6BLODRP
Xy34Cs3y78AhWrZX5lQgvwNn5JLCNsX3BYmiRHrLkULW6ucBXTN/3mgvsZJ5XzOaYat/YooN3HuW
sNWGwEyAXJUki+mpw20cnhJB1+k/wBdWQHCstkc3xyw1CUf9ZgkuuaLRWLbF+mg6HNmqeHAujTVK
3zm8+3J1vzKKX+A4WtAw5YCxJx3dQDqLOHE+IRbR/rKCcmY6TpsJKHVQS/RvAIk2XFCAD8JOtaQx
YqnHENF6aRAzRm01zT35azciCliXTaTVFFGfdlLVeEJ7d3p3ipSrwdF/LwD/ZxO7A6BpE7rBMyam
TTOYgQ2869YPnsv3TthAxic9fbPUg5aOscGX9/vJFJdj8ebhqBGEwH8MhIMS0wTgj+vsh63zGsQ+
zRU3Y+ixQ7nYwrTMm0PZidWvERDh5yAfB+VSkGkYnyZEt/m0X31C/FVs7v5qOZ8s1b9qTotWrHpQ
VCsVte1eSsoNRg6x4wbuDwpEVb0LwBYu48U4NMsmeG3Zqw/1ZhnTUXSAGVx+OrUJtZZP3mdrOufQ
Km5Koaec4JF8le/lf0MTbMJZxeHf7aZTlBpR1ySlP2uusEGXhey060VdTNEMVYuxkrg3lsaMm2X+
6FbXcoDQ6pH1yKMhdb83An+9KqS+uMHv63UXDebEFHu1OODVG5oA9GnnynumT9qycvEZ7jaVWRnY
Xz5sh3bCvJgWBmSlq1aquFZcgHMkt+L/3vebxBRCbI3+CR7k+6xgUuIgVXq5YCYb0Hipjun8luyi
1AXmZ0datV2gI1C+FSvgJEhenS2kiF9Zqx3XySYzAmMpLOb9noPeGBrkbxrioN3FiEv3Gk9nKwFX
2KzVmxSCwXgoO9610WaKtYw+a3td+sRi9K7TrDkI3q+ofZDEiE/n9xs8WkM4GJ6PTFHuOFzTqczw
7JmkeVDwM12Qb+bHIc2amj9QIMYX5LK0IqVetdr1dIVIcJNFJemregDnc2hxyaMVaR9FowXodReH
et27M2x2Iz1IFyPsr71mO1tUzNCTGQbopdau6lOtx5h4/IERKkHJ4o34MvztL9CgSwacr193uxkd
39VTPW8HHwZLEm5hetGWPaCYRiru9Di5J0zzgnpttlx7uGJ6un4i1NtrqiysSR0AfBIkHSomyFQf
1Cj6/HSLtDJv+hfCoveacAnYFRHuV3zkZTJeqNfVsxQVkJ14DtrWNrcVakwhq/yJVWv9edl2yoGG
J2LwnvkBkd2u9eAmM01EgDtKPQlYBQzzZh258GFjT4d5OC8AEHPU3JZFMsxuXi0Xj2rsxD6GJQEb
zH4iPJqtQj7Q/az0A3GYbnPKprFYJcexhjhmsqJRNLNU0Ma7uZL5iEbdA9+0sPS1+9ZrHL8Nr7kJ
EhxtJdn+mPzz3i7fFVa8sZVggmsAlM/i0w3vEZ37ZUguBf2aGIy3oiI17c/tDo7ZRSECkfggdww6
+9iArTO4HXoHXUx3tMsV1KEYH8M9BLVXsLIeyN11Z4BIFA+23dBduiVNrNUc/Ypilpd0Q2McVske
SlD3gI5vHn4t2kfpZ5pPJsOtGFm1Z2i3rzV4G9Ci2w6kqsa7mVu+DLMQVkZYxOo8rvoPNeYHQCNz
ybXHj/osdtvtmgKxSuLxFN9QBF+3mhguFGC88c8x8+SJ7IIdtbi+BV/CoCRGuexPd3oaEJm9Hl6h
04MD4X3FdnmKpyvuR4lwjBtbLDtCR4K8BHywZE/oQvKWYeMfdGbihWxTgEb+r3fQfxDmH+3NF6LD
b9E2WRMY5bOoMoCx714hXdc73PCCb/CLtNMEFcMVlTvrwz9Y7PWQ70wsy5VjB47aRcGWY1gNPjc4
QD2yjkcFKYjhRYMWSB7ujFz/l9Vgg3w4N81AYbTIQGChcDQJFVTfcjazz0ia2jgFmcIn9SByRoJP
kT9MlbZeVEGHXM2n32MigIQmO9hN61c9ln6BYpRyj+eMwcTqecBah8knoKr5rWq+WyyKn8adsZCO
AAoH0h6veLRukdwwZdP/v/9nps59KRxh0h0yJcRubZolws02S5981l08Rn4twvgk5T+JJl8Z27da
Zh/URpuZkGYYR6h73mERaslspZrBskcyEzblMJ1O4FaVD9YGmCr8+LPxvBMjTMyiqET3kTM/ugq7
M1+7UcGY2pmyPJbwTSyuilttFTsEuVkrc2H8FBKEbCs0GmLqYYZBqlNe/zdrNjJNKXTe4QzKpswy
w2TErLpwJ0WM8kDrop452q+cxC6chOn8+I0wsqEa5x3WjtvN+EygjyFGmk8vIlM9aMVrn4A4qJni
l1PD1RLdjiKOX0DU89+X7rypdss1WrnOMgtorDRhcGUX7Vom2QNvSc1snqz60avi7ks+KOdsHVst
Yz2439rnvqitut4qruTvBJCcS3mwgKEhbVgbOVzIM8r5wxMT8XmIzktr+UkXkD+QQ9RE/YwGQxxW
sCuWQG+yvWk6rLVe9rwT/AZRgpXJSAvQoAxWPS6NMOtfhQgnjjFYC/9VRHIGqafKMAHaK6ssOg4U
kG21lgFHVl/Jvow/JsirbRXzfsG25GBPYspV3Ql7lPmbYwEuE1lqwURaEMLdBUPLGAME/fvmqfI4
Cg/pyKLGSywKv8Ors9g9Ss1jFztxRp9bk2zG6C3luUn+uVayuocrd9CtmIISRGZh8pacSbc8spSq
Nb3zVahPWjVT2JvODpZUZdHB/VI5OzQnM65/nCNcuyflAaQC2CNN8AHdrntwO2Ybz1XPAMXJGFOg
wKvbNWR3yNc+9EK3F7cT0Uv+s3b31GlcaYUi5f+Cgt9xl1UdUE/bHByRatE8e+V4bEdPnytVCtjh
BjmXnv3j3eysNfM9pF2049YO0f7PLmVcxncrkMXe6pvpXmhTFjAvVHMKtDPuI1NaYUOC12OIjSGJ
3YRt9J4nQ82XKR6pv2+Xo2v9JfP8aRKyBz68cnZmvtqo1RfCEYAKHyKP9kwNQyqQfBGife0WMphp
VQvpceJ45ahNwencPkka+4hGw+73cu9xTSc8pkBB5qwpT0ca5OvmD4OlF+k0Ao3YxuzSKTXZ/DNn
xfFw4gffZ2peIk6J1V5ratrHkiWrXMAMUhCp8PLGVZKCF51QfN6TSz6o1lpSn5YZ9U8Vs4DxyrxI
3zkrj7Mezc5mODOYo3ePCjrHqdLT1N9lztmlvyjdMCHMptkve8j4l/5WZJnvrW0+cKpB8QNd5f/p
w9sG5jKwPVvTfDvGR9voNQ3TUQcr1nWnGXnDUjwKVo3xEHJTEZ9yJJfugA2l+bq/p3Yj1LGfpQEr
Ya7CHM5jLsOVbiH35ntcoEAViyn6cMd2VjcJdQkviKObbRfISE5ecPGkklwkmHCmLr559acFU1My
27/TILUQflG9iHWNGSxWs4N3kZXIQJZj5HkAb6X+e93pkcyaaW+LbBwW+kQ2xgCi932SgkW0Sros
TS9h7UDA5vKAdo3JjHL1mcuL/Bm4+yh/NyYfe8ajEsp1JdY98QuFLcn/iVN2Z+ggsPr4OvVEUXvG
oPp9qB4LD5E+EYgeBZl5vDbqGewJ9fPH8oMMEvBiom6TzKxW6EYdRe/vjRTmYypudEqJRWMhOMcz
/1N0J+1p8Es1ZyccbILbJPvg6TAfNW4ktCqTvn4aF6NS6p8RxnvKfnKzMa7ObOaLtJq1dcHXTqFY
8LIPEuxYPQ9Xitt5HWXOJCvPwG6hfy5Z28GbXhmSoZcOpG03rRqZEVVyQWawVhGv619d/4eHHBwN
3KTxHoAM/FWGQFl+XdqJ2COD6c4tlAWD6SMonpjGXIixb2oyGGVk4eh08fsgtO1MF6ucsebb5LA4
GOOpe9+4k5ltMm6NKh4DqM0EnjK8W7GF+WJsUYhad7pA4yC0yzA5qlqGNIEiSiXOxBA7fSfx2kLT
+3dHb4+aW/wAj6W3SKBwysvtVFumULTs+b4W/m3RvT9RjtrHTdDx2EL7ecMCIKxzpQl1aerOCEU2
XxWiBYOZ9DI6eY5QjDiIqgw1Ew8CM+J6vJMlU0Ec/fe/GBmBfXithACbSpHDtVIglDkmh1ptPDd3
NiQOMKiHrR4iJBs2u4YNhfAVTmZAl9egkY+cI5KFbvk3KfE9f3yk7nwP1xgLKaLMoh89IJPV0WSM
BzDG7TAu2K9JyK3KG5KGVOD3Tfh22YbUMIaqcevTyR7ghgeZj87xMfshBhO1CRmVPmjmxXXQD8+G
/po8N4ayjW/O3Nq3ZZVRvzC6Gl7R8xMB+eS3seIniKiN8lQDqRrZvcetZx/IaWFIgYSBGdHbteM4
tfhKgYzDahJ3/STKnzscuPUnxuDNIlMpUymKb+tg+Osa5o00TaZqiiJY+NvL69Tat4stWCNIHOBX
yYumsbuvF0KmtautLxYejPheibUQa7N3Tt20oHrb4jVzVd/XUulfa0z9H84FzFZP6AcYhtLDlHmR
zetlONbysYTm/vv4L1Xt6iKyJPoe68JkUrUjM3YeS6pZ0rp1lWR5omHFCw4VZvdAkF4FMo0pjsjt
hYVAqQfHpwOsog4fy4I9nz4fUWy6THFY5Cu3O97mrZ7+gQb6tbfoBBTgBO0g7SOT7A09X7xmv5cB
/V/3aa+wUp8WMVbJQOFc1ngFfUXhTSm//lnF0BWB8qaRw2RhPn5guERzBivwEos903zQUW9wQc9G
BXgBFwSM8eEAi2Vq9JlL/wIimlKFC6GjJJEF5BtDl2LBEwsVj+kKgSaE7xaUpfr6syuVgCSidYlY
zs4XRwQLiU1lHZGrCbW/sXJyrryoapGEbvb7NcZ/UCo/zIu0Nw0nlyDXnIATdTge+bR8NMpNTMn6
yxGqv1URstjtNEH21uU9ihANnF/IZp/a2OhomUcTLna/tIjuqy6TwVF9CJ4oZuji6IPwSq1Hu/og
0Y++KNNfjNdhJT9gLjIagOH+twPah++ahbjyjqtpK/Cd8uMpkne1j4dVOej82RuICKrSD/1/a29J
31te9A1hiNoCpEjlpxCXeePKxtL0nFbNEnfOcXOIWQtxjc/iAlD6Brtx6XYRCgrJaGt9Z/hYV/+0
haxzOAsEgab99401VGp0aGHCuOQfUaOAv6SYG3pDr41CmLfpck4DfIz+MOn51l5SiUPj8JZA5F7b
GwhDe+EqEdsea6BdOu4f0/xoObFDyv3n60jK7Q+G09Onz2oH9S+SZYbdADQlIzoJB/gjdKhzjnBt
gqjsI6ZetC7SrQvJ/9dCei8XDQernz4bvxcFIHoYI8a/lZb2mFvbtvgnnTmhqqNtNroVxo2Boj1F
7qD9AHNgZWy6EP8/1v5prTyepcufVtAVqW/Sd7SDIohFvILUGMkEKyaCwukqh6AKqtPlnZyo/OgF
ddWueLzx6D50J62Hwu7rL3dpsWn/W6WmAe+hJmTCLEUshA8e3A+KdR2lP0agu4SYdnW6y79pf2/D
YHtyZQ+honM+oKvsYw6cvKA6u8so2eAFAkuCCezi3kV2g22Ik1ZQ0oeDYZJXCCtWGW2UIRqe5+5A
H6cpopP5KFlKkWA6HKnpKj2z3hFG1DDn74Fs9v84jsOzSldHXJlqCvGoICJEQuhGaKo0CEPDNuGX
2r8uQuadIhGoNax6RGXRCnJ62wY1r5SbxyIAQ67jNzAaMurDvb+/241RiEqVh6GkT49xEUPa/4uU
bVWZV4KppX0K0DYW2StsuiH8jqiwjQL7N817uVKJRj7GelqZbIsVt0UwKdykeS/TTasc8kXc0bjO
rSacjG4svf82HC5CwjMJ7NshEIVDWRT5dn9aos454VyhXbVI4suCfjG/nKBmc/MlPpKh8btaj13c
maJ1rBCOkOimcn27wuhrT0vLeZO32gxKovi91g2PxDcZZVnkVFWskd6R7X5lh2dGPGC24M+LT7cA
UxP7DWT9GrThC7KZzzeUISKkO8v9etdYxsbrvBUDRRyH+iaj2bhJuyDbTlQ2h5ZfTIPlr9VDnW05
NKVy/LQaXAwGXEEwY+FVFAlBeO8ytsGgj6bl+smFo4A/30ctSWU1QSMcnTFRFgFhhUJ6ASM2FycD
2kUY5vwFz15QN7GcS+IfmRPSL2wiGxNqQzMX5lOuSZy7beyyFuCd860EYaoVOahtRrAivloisomH
cHJBqfT4lDgfeIX8ZQfAEe8yLOOTMxT5QuGp1LxPBEa5AA7muKi7hhjbMzG+3dqGaG1PunQLI1Ah
F9XtILGUHTliycwFYL4wpnLlV+TwhL5ueHz4ZHS0Y5wzsOYJJqJO4wWPE3tTyll4+jc0qRXIjKM7
m4giduJnwuJi7FNuuIOPNjYHMg9v/stTd6eHExycCcX+pn80JgDeNm5FAwf7n9rl5Cvq74JHZGpk
kby+fvf1NLrjNsYMMkoP/gh2/nDPwbBbKq7vrlugDgJRT/c+oEgPVWnrtpzyAYXFP3q/tZC6gbNa
Gthr6Hauuo7qCx3jjcXUN43VRr5h5PJg3FO73Uohwwv28PwPaKw6oINevCvnZS+Fb+M1/oAUTQb3
MRluCZPTiOSPSop6DJ3e0QZyx+E6bYbqezD9xlKf0fCa+kkLA7CBOO4uTbe6cRXR7SM97C02n6de
BKq4yUowZCNNbariUoHGxaLwuYHW6upRO4z0GMknxiklnqXBeVNPUMMLG548qVh1hjEkaXMG7QWt
HM+oKWTUmeXV3g8YIvnBd1FGRzFsfoUQ7QrBT526yVCEkIfovIRsp30PSGUtLzAJNIxlrgkjsXaC
P46xt9rHfKh0ozBARkJPgoMLpDem4PM0/+tZzVU6svyB1YIBEnul+KeFNh+fzexFt6bSQENdtALZ
pRPwbEXkEJS6b0fYzx+myCDRqZL72YPxqtVWkCZ7NOOyy3LKUSCMC7TP0Ns/KscvW9csYIiVwGcw
U/1NzN9+lDbDLNhqlPWZW3O/seLQLzyh6qgaecNzv1Oz3plLbI/a6ek7wnRIMlenc7pdJRluhHwT
W0oAYp/vuIS0k00swHmRtj6BeHnIl2N9dFoXMdC+qSyQ+t+26moEWApDSwlkvdZrMjibRVukFVt4
O/vSdQYynE4vLXaQRcI3x5FyEejhwnytjqAi+JOWe4dpfpmsuXxd/s038WApUh3GoSQHgdcoG0FD
saGtViY/cGJ2Rpgm766yCE4GHRnYHS1h/urnfbY206VWFRHUuG+jtcL0VgaoPdEZdN8RBoVs6emo
RzEswp83sC9EfTq7rBn2uPwWL9q0xdluQXf+mgOqPJvgmLMuKJPghm4HG8OkcdSWtiotFP5GCCAr
I25+IzvvOHdWScPcsQGliqbwzgG4tQ467q8XzB04/16WzarLnxgjXikM06PKY16U4V+ZH4bDG3Qh
jegxmlr7CMwgv5OaGu6gIroEmmFd/8JvaVyim4gh8pD378g6HwmhfvgBABrIijiXe+C/UjuJEZZo
8Vuhxv64uWgbCKKu77ZgNkj7HCKXZanc6MmixULM9OccB1dU5ym1kyNlZyORUe+J82FZ1AYmr9mP
uGwz+tCaXVxJXfa1TrAxQqjx7ZasTHUphEVJ8sArM+l0zDQW31AoJx1n3MYFhut1qLNioiD3IuIX
YvZcWRdbeW9Sy5+vy7fRMSoCXhut6Q8CcRLUbvGubI+/JC+3f9fX3mYxdo2WXdeJPaFoWh4R1Mrq
o9pAkm7VrKJ5eTp0KDQgjgzmlgMxWYznQmC90sYDMKNpp4Lzf/Gg4f3uWYKA6/ZrN7PFRJNx1u9f
csYbLgzcF8NHBxNMg4/Zy4K1Fe+QsRQJXAAo9zlj6LceyU1TpXcHiQ7S8lRZE9ckP1f22t+cjNx3
Zh+0c1runVI0LFQsDv1YgKi2K6Z0kJcBFJtGQgvCkg/4iHtOedweqRUHoUyPoBZcjRsh0AQyigMr
yivGYxbpNgn4UrmzqHKqzo0RYGqJKvU1sTjPOfjk7daFjeTk3VGSvd6xfRG4upkWoVMm/T7HHq2Z
MplljLFTpeG/7GDvLGwteLNVGZZN0QXDuCKaK85PlGQVNrMTiY64wDX2A5Y69o16PhMP+NT1mfoj
ROEg05PPLDMMdZAB5tCregtsa7p5bfZZcPqsqI2MmA/35HHCm72Qyszh56dn3NbsIrSUwnRRDjqc
6awgi0wanLbYkJJw++5YWs/45p/8yWbIuUhdIWtcrZh+IcyKxl66EnQpZcGlgo2RaRJGzdl2vWaX
82AFiINEaL5TlD/7lHkk9NPyzStZGTZgF6KvIA+Be5KaPssN7Xct34wSNu4vqQJQyDRbaUUNVMmd
m35ccnlCy9jFp9QnDl7vD35kAeNCOJGPKNEr250OHNke6ugX088ZVb6FwQAtpMqRwXyxFIms4rbs
EehPdFbE1S9Ne7Bk164Zv3ZIsEuyFkP2xuYbXjnQibhpC2byAwHO9cYH87MvAKCFOvGUOze8HvsW
pAsAdiAgGEfeHv+QIaR6aqHr2HG6sGJVoItzXFcokZw9AOShlCRMvjKG2RcvhqfHlw1Zd09m0Xs/
tO2wOsttrP9O+UiqEbYbvp7I4X5mXXVMUdFWh5YuhfIAMMnft1awlgUwSUGUVRfMNQoH9C6y8dfi
P69cOfQvjD39hz34yshyoyhc21RGdSMSKu2QGzbYjoiShhVbo4NuBheaPs55XQbF+p677S/sdUt3
Ki2Tq9ZzuiF1rM/EGfaDQbLuKO1q/exY6E7l4DAsNJVLkCEyT844RXTMqJOyBEnrNgjjdw89gY+2
QM6/9ZG35P6PDyEc+cdUAyr2SCJ4kfuuMJW1T1WHMn+Xk63QNZtUXT8KZLwUbr3l0K3qLBDK1ldL
9ZtInW3ATJ4daPS/L+gBDCIcbrzXsxe5pjIpzvJ4SY1PPp2YVBBcO+vdM/ph+gKGMdGrxFR1ZgyH
Thnp6TnzIrK2ylVhGHIOnZwzw4jk5ZaSB6woA2pJpQUv0wmOVyBAvExXSQ3JUPfXorQFRkAIXyAo
uTgTEfW0CmUh8dRHfk7oQ5KO5rQ131AkGwsLJ25armn2JkfSy0AtKIJR95HhjlFhSha80cMSuTOf
2AZzWsVJeASEhP/YI3ZSht2k03X5wYFUibOeWeD8n8SL16kf2if776OapGBJnTtqzdXak5Qyj2s0
v22qqwFYvq6KHYOpW/MxFU0h0UY+57j01j2I+JLhP3s3b40zJ+Dfu6wKhvZtpwm7F2n9EOtOiDA5
MGJ70IZ7WQ6VO8nsfApubhHDp84yNTpyzucga+bcVN7PqLqPK5wrq3Y71fot2uTYB00KYXrhc82I
BJ9bN9ueeQdbz5ChXtbrx1SD0UHmARabihEoHOF9BQXRgL2Bksbm4IdfnWfUQt893t6K5LGdicen
YRnZFXVdFhEL1NnFnAKcMrQFWC+DJElNp+0TWZpZpluJLBupUfmwXX6UTxlmpQf4FOOZM9jjRgom
iZ+pW4QWgQW18vpndGpdXsmWXoFvlvtsbm2liAYw0MPsLEIchZ8DeS9Ev4tNRQXFW8QJOt7kHl27
HpNp22bdWNkwnhX3ROsl++HNl4T8uhi/5Rnya+BqR2vEZyrUCZR9D1BTFnHNWPvhxD8NzkVjLpFD
gQ9fwXIP/7r68p8ELcCPHwWKq/LX4vSt5z1vHvBRPqRLfI81hv+L70qwLB4KTTp0W9hb+YCeOssY
AhkbYUz1HYGxCyJSmCnj0wMDzShyO5+wkn3Y5Fpzckr0E4BUFFr6329+QzePVwN11HdR1B8rHlJk
7BHGG+hbVw3oinRCsKz8586Gv1C7CECotYyrnkDjIw5upAFbtvD8+PhHg1fk5l31fGZBxx06pIJ3
IOTsNnpZkvIWnO71I58Qx1zZYB5Q96+39YX1X7TzJJuWyHWWYC/4SlcjE7NJcL/vS/oHYt/9ArnN
9PTqXSVdijFdEtQtpLCbeEClBqIluMBZwP414g+rbW2BsLBjVzEhIk3IbGbwazVdApqERP2Br9Vq
OaZp0GzipAfKXhj5hWboxliG4ZzQyhHabd8CEakzA9EhCO1OBXpQnw7Cjf1z2UeWEiCMcqZrc5YF
uTscgLPsfqfoCmZDlp8sZlL8+yQqs8tfcWNL6w2faiWLsyF6uJ+C4jOiKGHXK0nFpDRfQSaj8ZBH
fSoQs2x2Kb6PlWKhIj1WNrYXJQZjoBf6skmSm5hwqvRyS5AHxRddbzj+vonfWO3iOHITzSUX/350
h2mbnDi23Ht2eymE9yKwLdiiB0XeUIJf7I3nWDTAq5AG8tUSsIFwIe/Y8fwAHtjXaWX+sS55M20I
QysAPVDfF+Az516Vh9M5IrFOTnTWyDUh26DFOT/GxxR9jcl6BYII6czMr+BoNPL3lqFqY1GdpI+z
373grhOrJ5+u+IGq5BXr8eQCPrptDKAJchiJAqAp8W/L+iowZqV2Xf2f4s0bVu++gJKhn9PWObbx
+RvC8lVq2k/SeWfXzmV4rE0MKZWbIcRp/mVqVS9AXgnhOwoiwm4dd2fJg8qt4eeanHi4HTixHsMp
pxD5W6LMiy9PRlWnh63ilHTlnnW5M6+8fWni5f9Sx8XBifAeJE9vppBLFzbFPdoUPSIpdCxOd7M4
6n92+EETIUwT0tq9IkDIwK7UkI5y65lvE2ot+L6sISX6kKyRJnWBbiPnAbSJY5JlHAvrw3oAd+ZM
Elja14E2LxsLAj2lcKMdsmaKu27Fj1yp2IvMO+54lOnI+iH1UYXDSYdDu3eMAOBY7X/0cHY+hGZN
k3piFegzuhwgEJkYmZ5LLJqw/PjeyGgD3MH+6Bc8+Jwv66niHH01v7DyRSsmHqlOGU0LCthdpGIB
Atyi+K+4KOXzv/qEiZQm9cW6aEizjQSX80zOtz8x/dRZALbe9PE4znI/EsQBZ5ZhcBsE0vE7ZgKX
lipj3wydcP6EiyqtRIWy8MEL5P+E4IKE8jfoT/I+jJcS5GMbXTneVm71Ut1c+a+RVN8XcUOvYvzT
o8BMvcR2RCD5hYZT2xfEJSLv+CW4HZFoJx/dm943RdiVsgAm8OLqjUfvhCcZxWDJRDk/RXGOgS4J
/OLNz0jliprUVh8PuGbjRLazZkYISimfa5KtOFYdAujvZfrN2RvqZihSQKeYq53DhloGA3mOhT6/
JOJujIe6PhNdVdw6WIMW447ukE4C2GXkP4urureWHDrEwiw1alryLDD/1Ugu3wI5XlKUkYMpXS8G
bu3aSsHk6nUHLwOGtxnSpIoekqbGrNudzfdEksNNuytcVWHUuAuhM+BhOTlDrGRGqNPaMVmIwUK6
vor072D1TVJoEe3FqaQxqriqxgbb6qJc1vT3dW7nAwdZlq9fxvNj8J8MwkulbmkCThWNOd/6196l
yNxCXooF0F+wHxTsHe7Mt6feaxRJvphYkvul7MJ/DFum9/AjwigppjAfLjLIu1bPEq3LJt8/r91y
ONLzTAsRkGsDwx3TwfSwD0BqUVPoJ1sahP5PMxetgCU3IOgrFuP3P92GHbHZ3C/VX4+cv4Fxehog
Cgtlwv7OfwPHQ8zRXLXdhJ/isZ0Wx5NSgPDtgPM83+43NPLL4QsBl6hGm3t+ViSFZ5OxULekrsOm
Y7efapyg8WxejyoLkO07xVifWNkTr2i8NIbZo3fHQOUuPO9SWkWou0Q/oswRGJlDLGYta4PA/4Ot
EirUryu1LYTav2c0mGnUpQAHlchHBmNCDmtYid5RUGG77Bn3TkA4s8exy6vn4XSPDEW1NavyVLf3
NwAlvL65TKuLLC7PRCFptRr5ynbC7VLmYbV45QzlLVA0kDJ2KkKvNAF07+oF/2HW2yjweWFDoEzI
GEh5HGR7ji7rDZGLnz/GJdQhZnWpaqWTQoDaa4Yd7h3/2f2n/GLBLP6Jtm1hZPLOA48WsSXRqMlD
kWIrUC+PKmyTQOOajMpTwmX/FnLjOzEaZpWxRxbvbRqkqbvRX6Mtivn5eLIgsjt4ND84nmPZr4vd
jmwIU8M/RGpkETXKmjHYgzPJJOOEPxsdjvBaoRfEqnd9en/DSobKSe/WJtkCD4CDRUM89kEecyDB
we2ACK8iR7GVAzPPUgYzkcwkVJqnChQmMNd/UzBsIF0OISVHTrQzAtC30tKtlFzmlTjwT9xoPcGj
BZclxgWBgk36Fn8tzI5r5/pSzNGTO6R5sUNQTzrY1yKcC0tFnKvJid1GieI3hPidtt9wJYqQHSM0
YniO+eK+I2mt8br1f1ZNiv8SUu6qHvGyczZJ2fmFNR1UrA1O6Z1RtevFMu8AYG1YdgxIx+YtwB4k
cZMSrMr4tusupfHnt36BKF+XcOHWNBeYAizXtt/Y8tPjWgge7t/dJTqkuLG8Z1t98BpFSdfloQFk
HxvcyCZP6ZBzXHaBXqiDEMsIMrVtf1K/utofFCc1OMOH3Y4766dD46h+iAK0eG6Eu+/rf8EYDNOQ
YKrbI5eTw8Ku0JQ6au1X1vh7aUa/MwBHXK9FoUwLDotm7lM9z84LHKRbYTcaVXoGxE774s/S6OQX
CMAkaRFI89qGhXnGQgYfELRGxZajH9bFi9c0WupJCpWKv/bYZR7KO8DdA2HOJpijCMdipY1xZRNB
H0LlOyMhw3MuRpKOepM/z8ZAWRwZ2gf3uLZylHm4JsmLECMlAXxP3cw9IeT4BqqJ/Kdd3AXo1nTZ
RsDNFpteu9lbvcWdAyK5BWNH3umfekwGpIhcZuPSaaVukOWTuTJHtvs0fMOJw4GMAU5fOJ53M/y7
N/kdLIIkYaxa1DpIX7QU8mT5x3uCNHhFxcKv9WmhpeER0L5mKobytpyxMcbxg+rpD9PtreB9xLqZ
WyaMKX7alQMDpbDx7Sd9pIuLaZXI+r2X1pwisCv0Xb8x2u28SzlU4HzeZPUj2ufn0JI454gJP8A/
NCRtGXpST0Me/jNZHCxELPdAvRaEGuk+WEpVGi0W3wGTwf3tFla+CNj6KRZd6fbNiHn7GRP05sDR
pNWQkSXwpBs6KuYLL3nOTMu8tnMNnalSnIMlagH9PJHZJ/YZKmPzduJ5gs/sJBzcFEvjG57QbL4+
aly79F9SXpPhMtTOCo+/PcEpT+Q0yNcBx37gR5tYpip0qS/twCwaUGMlhwh0MOMaslwMsL96HcF9
pMq5qsyuWcSb60ROCuAZGoepHjA8YmApNgP4mOuVZJ8+oHtapWDhzEh3J+/3MNDpk0AhKGLwyHwV
pDRNQdlWckqpXBChmnB0DRqucWI4sh8V97LTk4HjNNfJcqRFDWf6lmA4SlR011HCyAqfske+OFAR
1iqKGGmwaVvWh65Ytm8NuY+gtaeQv/lGRtbeD3ZbJnEx8Y7pxJNBj8PYum9qDV6mz2M0T/p2065p
34pgcMqx1MOBBUXSzSDV/x6SHTGnu0l+SUTnA8j1sE3Ok+Pry8jYzMd7Cvp6IaMa1DudPbWWkREl
b4t3bKT+SkVskacyAZT0bp+0IEBNttvu5tzlz3WGmEpxOHaH2gP5WDqEzVDXDh1NvznoKtbcXC4M
1kdeFmZR7SDd8VbdI3sgxys93YmhMdBArMswFJ5wIEzscd9PIjFXFiZyXdm2rjSu9j9NZuPZtNyg
xrofgkY2D9YbFWYyZPgNOXkj7mwaVpPPJhzKSkN9YmLXOEyechABEeYLYXAFUFyCry/agltVtlqK
H32rhkK1L6I8nFrExYUjeGZbsPDS2cFAqecF4uyGQ43Y4OFOfzrCjwkCJ/7r9qkoc6LlefBSgGoY
82H/9brNq8eN1gBhtCvaI/EGsSZr9AzjnaR7CxmKffBtfTgCv0rBhBJEZhBTTjGxGWiq98NhGXQe
RLmuAJZ8aKauptMw0/lfFkwpHWWR6JwM1modqV7wkTaP9NQlVicArUWqLNMSaXF+I3cqMp3vARO4
+V0+UpkhctYvK1RFbBuSHdsATaFgYZPN1RAYw8NKqzNbx/KujTzFGVjUZgGMHmc9REnF5XXV6CZZ
JHc7tnp6BUEq1k9njM6nPWJAblRwese3bZOHyIukRsUFhC3xDpK1l7BqFovOQmhfXBVsuSkkUKTT
ytBkcmvTFm3WFLuMN6wTTsFtFK5mHSVRw+8b/iGU+93qLRn19jgYU3WLtNRnaEjf2BNsq9RyqPw1
myvdHZpDwbwJl/qfdmsWwrjKqX/MkTtla1ITEPkOQo7RpF/tJXW66SzbXgJ/0gj2tYE5sg1loR4C
90Cf8nykN3WrtNbIOW9p4e/R2J0kOmozKMW8wy5p3dX+u5lGDRYeOXh8PDhAdwzrBnsHLPcYVzR+
abtDwtrGptPOCR3Cty/8mfKG7FNLfrH9JVXB/q44PfB49ALNEQCMKoEqQAcMAHWmeo0V5JrViacU
f6FKhnmd4g2jQzc+mEzPadqEnjJ+xTq0XZF0FKLKQmeRGPpM9TxCM53YhdsjzE9/17sy4Fd9JemT
YLest9pdjXflqhk1VsILuxgpFchmu9OVEaMcVgQZEqGqYu9h1J0smuqmsRFkh63NGPvb93nJGIL+
9LMMkv+Piv9xK33aSp9PdcZhOHbE2xsLjPj+4wxNlgnvhulpNzBr7CTvAlfStaT3V1pG/cmuTYgq
Mv1nR0lyX8UkBntGxLMWmYq8rMSMblDnzhD7n1OX2PTh0sM6gTcEV4Ak7dN8CTIcNylggfQ4oyB3
RNFwxdysCW3V02PkeYF68VFwE6QVBYC/jHamrcY3iqle0UJke/VC5jaHfIYrvVaQ1UFFPmQa1ITD
QdziM3krJcaQZVG3g23GHD5jmwOmTztVf5zmVAAROVvuXkggwxT8Xg04UxLWV/vSG0LEeRym6wAf
khcHGo34XeI+uKI7KDadveaSmIDHHYL+yzigBa533GhSphrPBP9IPx7lQ2OMAgEV8hvNeYZsvyyT
gYRZHi58Xl6bh5ZC+pU+Fg17qZPv4wGiip1nVz/PWlOe2nlL+dOTDF2FRyrerfN0dfoBx1YSKEGX
Tep9usRlOOPCoj7sFdbGK7ef80p28XUOpA2sSNwIQ0cE7HAIBSPs8boc+WGZq5wx9TdMFgtRqwos
ggTNo80=
`protect end_protected
