--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
iu5eeTQDBHI6qec6ippdkJ5rwnXCqHe+BrmhLV6NM+atNkp/V/OhfFWZviPJJXSHL8KXRC1Ft+4D
0X2o+zJ++k2BX6V3n7+7SKpK40tNYmDLoij5L7trW8wRRH5bt8HaVLfkISK1uVjxlljsDiIvmpds
p+Holjvl19ZCGuR8ECwgRdCVynDMnvvgMvx048bd33U825v95Dm7G8tIdAloV6EfhypbZTZ2eF+g
yRAMqvOMXo4YLlzUOTJYVQyND/dholZifQIDuEwSIEW0laCnMvzgOWD1JaiivrsjL96XBKcpxlKl
VIolWJcEieTW1d6jCwUAedErb3zRp+I3fouTEg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="afWyvdBlPURjxTagKM6p+77nG4ibicupit5CPguKfVU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
VL9LCqN/Fq++CRK94AmJ8u0Xsk2DW42BUfZWYV1qXfzZHNB/v7u3am55RZR6HMqfE2dw8vGTe67/
SX+McmJTwwGpkZRfg7pxNkW3SPa+rpCfCHYKfMdegLuGMqXeLeCj3Wegz/EvKhl/RFE12fKhSY8X
U7fG4qTm8tqa5IP/j7jYrkEOUC9Nqmv9sLETyi92wTq0q/BV3BREpqX8igorLlMOgBFLPfUq68C0
ut52ZFVlsXmc2y7hQbzvCv8u3qLk5FfoJZ7IVMwBH3V77sucMTGSRYX/YuVp94keW5LmblK6/cX+
mA309ACsLFANJEVQL1EfMBYm7EqG4nseKdv/pw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="hj6QWzMOrniBBNeDiW687h2m8xvYQoV6chGlKNYLzvw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2608)
`protect data_block
uEq42W79icPJKZ3PXusj+tB0h/7Fl5lXmKnluKrsBcDpy3PLjEwy14AIYhzbNu++AjouCwiluSZI
oN19YqhMsxbAY34JmAL24QUmvKJCu5QQdsVGyJGDm8HIAOZ5Vh/xJLNAogNfcHKXPvzB/REujiPx
35AFHs4pMyA6fbAE0My0uy5QM6akAXTxwz6vsQxMlFsfQ7hc1hr1M2vQAppiTMbIPq+DMBTRE/Fd
tj2Bmhh92GyehOPSDKKTIoitcp1gpC195FwA/hVCvlGY7/mRiEWhQzshhS/N3G4Jn+lWmSeillrv
VsUeo71jAxHJI0vJHTJWCJBlxjTmlSpN/RWGUpQunnByYFAjSGOCLKduSkeKax6zqut3vchZ3Jyx
ekUmyAVbCh44aucQZXq7QGft8T4eJ9jrtYrDbVC1+StFkNmK02oR9x7Nu76szNfExxYPSH3vu6Ac
JN9cyatCeFr+W62GbxscK/azpSvsOhArjUsDPVDzNWAnyBzsLwGF9c27wOF2p0wCWr5PvG11PHCX
0ic8XDjemiH+Zss/vyYQQVpHrhNrOo7M0/tt187L8dfDqA804IOE129dver8ou3H+5lj5IIx8WbZ
crH8e0CCQnLzegANWG2TaQFDXvUaqlTyL0RVfwUoP2PlO9DI2KENws+iMfXkQEy0jBw6P5vVGAPT
XQVFcI5wKD5fCBS4P7mQ8fJtvgXDqn7rP37TyCtb13QQEnwApMboqgvatBD4dL/GzETJkvRI6NwA
nGsfYeT9iQ7qVsEYa5mwVLXbbYy0IJU8Hfo3xT06FJA19k8Wmh1AQ1kA3k9mQOABk3xXWCL6G8dj
ew6Ww4G00OI3f0IzZEEw0WXiqS0mQgCj4YeyKR0HqTy5YwvyVcCkwuPp9OQnkJMuP/oVM6Lz2oKk
YL7tNF8kWBK8Ly4EcaIWuxheSDBs2XkSIB4tq8GZFISDiiAP0lfe3L30E3IDXs41w/wxPOfXQZTz
7b4BOVs0YV5iD8cQC7060V08DOZ1Gtu04G3ofNiKwVBjyt7336WkJKxAC+1fVQnjVHtDZ3UTFiSQ
VKvDPPvCjS9KtOcgNTnvECyW/KmqeGugWvxGf+I/Exo6N7RNdMh2zwiZoT+Htuc1D0boXUFd4QAI
re69HyijC4DCX5BWpUQff8CeLDiSUzCnzbxXkFAmprpBvHiER2mWuz9Qu/llPLvOOwzOrIrOb5aR
ltNhV25uaZqIjBXNDIeONn1U71C3ybcmAeUgPrzovlCOceKCC28O2l3OQiZ+S4YsOVOS76mFSUXc
3Ful5h81VxS/ZwiLw2/W85VghuqtGPI15slpuAsNiLwrVqRPwqmVnxODy7OuPAxIZKSAMlTA2/RS
lv3TWOYXHx5BNJMn8WAi3+8dTwrWIX/sC4dgYWkF6dO538n2GYfMy59stcis07geQEla59fvbOYI
zTteeSZWoayriU+87RGCpoM0XBGTPyP5+hzOzLR4l7shVGvLJKvaxBR3NK7UTOgStYiY89loXYA6
bAr04VgY+wD2xL1oF01953IwNrICr9H37pb4RbCxYxS35kJa22x3ZbvnHqKr81Mfr1yQA8sYv9Y1
1RT8DOcbTpGkCFwLqOuCe1Z1ewI/NkYIHhgqlWxAgd/PfOOmSKSDzDPLNu7oaoUpiGMvzkighMr1
AKNG5Fx4dnslB+J/YdMoLxGepOucgkb9NR7TE/cPX7JYkeLSxqlgwzlnLvG9Es0qf+GaMkuTG9DL
rFIAanSQg0gmTNkUq2DXSyPsHpJe4j+Y3/jqWqcxGtHMOFGIhJYWZc7bMkw1Th+PXo+OkRw3uRoc
ssijN/lh66oNz9JpLMrmbeoX1hjXQQTD1djgBzvsoJ886aor8ONXvE0d3agiYBwY91fKh7xXtkPE
4pbppSotPcmxj/WWB0KogQhYX0PQ4GP1TiOdwIZUwxEJi0tK+WCBdT1uS+NraU+WTTJcBHGfnlYM
RiPekHZVj5VfrevSqxzr+GNuxrdnLR3e3ry/UOHnmXPKS7ikzICPHFu72TyY+d75sUSIMbW7jk8P
/f7Zo/qYaunrMUa54i6tnguK0Ng66VrajdLBfxNg5m9hF3jKVFDM98dV3k5l2g7KlhxUBPUP7D+V
9bqkGUGkrP7x4hVHbTym0d5EeVXEYnYJpP9uo8vOa96lp6fqOfeGxogHR/mM+pXXBRoKPjXzrfaR
9nVVnnvfYMx9p99VxA3zUbrS1qN8gV22lRCsxqBRWDQEaywQvGAPCcRIbOIzHGa8+xOVOzB0nnTx
50ISZELWtN0L7zI4LsbqAwWUt4Sdb8dCG2q4uRZH+obdVmv6SX9TFKwKnZVNC8obMMLrvANLc8vf
d9kslOrN51uZQeEORpFh/z+fZp5gnkcOWEEAgIfOoqRWupubaMGbQuca//IROTCQ1YOisTWBjxda
MqzoeQJcRsxkzObqSsJJp2BcNKEITNCKVmNL+wsizd26TvrMWwdomuphw0DhNBvaTFNrw0kZXIK4
83Mg9ocN5jBHWLhzLf4d+JyUwKlliC8UcT7gTj0zjErJNqloMJq4IILUAW3SsRxvyuzWIOKVqhRf
JwUSh+odpIBpJwaRlJubdvZ1aOUN0Rkm+byIG/ug6artFeiOQ+JMhXpjken0O87tiBY3PpxzrsBD
q5eGZQH1+2/OoNVcCCJ0IB/DA5UUGKzY9YdzY8uffYR4qOsodJ8CKRO/0eHsKN6sVRSu/psi8La4
Pw1pFiFAmsNpugoiy+TfIqJbdJbFvR7RNDjDLHSZJ/ldVnSPS7lQ9joBWCXQJMUetSTuLXSz67Hr
7gdOhgKyC8py++LplyNe5bfs6jzMNIOBH7xiuYfDPxsKmxGp5k8Zz/0tt/L+6X16HFhYNJZHc/ml
bWYSMY7y4uHhztJbosRoGIpGFFGBmAs7nXPVG17FBTMm9XBcwiQiMKTYMpBV9peD4pX2FGTTumvU
V0lfhOH4t0zluw6CO1Le6LHpU6xY6xLWNT01qicMdxp/ukOlse7mcSVJOoJ0W2+uFr8cXFC6sMHh
AsnEQuiA7rTFMwhT4hqJ49o2KetrDlfweTjhwEEKUFDXnMzwL6nn90UoQsJXFgtUTwWbJyGt1ixg
iZO6FSZ68A0+mPXxacziFpWm2M3Eu/obqsKCoOx5YDzfA5Ib332iSP/y7Xq5NaOXfXRXXkG/5gOj
uk9EuZYy64bumI/7Cpq2JX3ffXoJKFD2vCOsurHvg1HYOVHE1ryRMPQqDa8UlFcAbe2eSMpQL5mY
J2IYDnp1vVlleFg0k7ZiDcG1qgddFugLnvMXP1ArW9Ruh4p92ymSC4D/MhnMs4m3ESji8PZG5QXp
l06nEw64I6J++r1KPYoFuyZdt0GPr5noky2i3ja5P1gBvb2cA9RYvvetOZrP+N6t4XLhIHD5h7Pi
bgkTNTeG159AWuH96hYP1vpwj9bojst+Uz/YlSWY6jlqHv7Dyz/yB3mwTg==
`protect end_protected
