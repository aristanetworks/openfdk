--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
mBC1BwSv3oDwUZMNwkqinh4/W88sb/WWcCEL7mWIG5QCrHoe9eykgrKuM/1F0l0Sfpr7Dpyg0z1k
N7XhmRsGUyRMouv+cHsdQRrizHFmls/44D2nqHOxiXjnvDg3NLFjg8XT1JLUkAFTre9oWSJoT6wY
aDOpzjxsFdq4O2TlrF5O+pR0aKwwLFwyqDqpuIfbwp4FXgaS6ZoxUkmQV+tBmfcuVLZYhthVZaB8
6cILD3/WS3lrVuLLroWNmQaodTu5oGXay/D13W+FeKg3BvkMBvHJeJCl5N8hJiw5jYdQ72TxE+lQ
yT8X8NhBtB+Odrg+2seQoUgS+mqrsyqExQgZdg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="tMqrEY/l40ZykIzTA7G6f5J8gHKjNOfmdBId4sDDv7k="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
Pq5Y9ELPxfquT7DXO7YJ+Hxj/+hyGQ70eNVMkWuUGwXq4UNt98Nvg99XJhmgGYDeQBFGWRalo1DJ
K14irQug+nDdKkyybsKC5HsEuH3yDnUEXYNy6o0h7GWeFfqC+CR+X9EMSe2eRT/P55xK1zBC9nEh
V/Vhr41M+dVTUWCLCepX6u+3jlYStcCjUBjUdTV9mVVMbdeCTK4txjeOUpiS/FliljT9ufqC2yC8
1JdhfU0i4PqWUSMaoLRDoYtRvOaJQmljxrKWZv5TKfXxh3q/q1UrCHkquL715OjlAK1VHvh2m9xL
pZk5SiuVzT+fBcdgcdpkb6B4EBQ4kYP1gcUI2g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="kKl6rm/kmbi3MgcYxDOoBj5nCbYFZa54H5qKDccIc0k="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4208)
`protect data_block
YYFEdPRWVmAunV4haKnh/EayMh+eAIrq5l8E3Mltjf0osnpLFh25b5zIHBHRs3PjHpODGwu/d/p1
IlrrTMhvDs14Bc7j2ZInO3yLnNgVqLAHB68PCW0qntRrlhJ4Dyi828Nmzt5bEj6BLLCAfgeWQLTj
peNtI4CLqxgCJJIAtPcNUzsx+Knzkq9OdvPG50lLPfM+BZvfVYtzyRieb6L/p9YIYjHGTePDviSo
Tj8HkHYbq6kBPrIZa+AFjx0OoRMd4zCaCzmrjg9ZniP2zJBumokQ/cy+TrK8TToksKPqu7XzBlGg
3Ykg5EcOtEYA4+I+AhkOWwGUmHngRxbX+Q+7GQwTeyX8fLuhsEEq/YOzDbhYgmGGq7S+MxcFhPPA
MYfWdG0CF2bFQqo8esqgvyRxhH2EWuKeq3vCi8eGHzJrKhcfXAFUdDfv9TmL6v/xG7aZLclCF8K/
5gXcht+3mvHf2IRYoyKipjiPi9T3P+wsvpx69ZAOtO6XGsOrcxm1iGUh1opRtbZN1QvC0PtcVWX/
T/kb2RTlFah+UjG3GfiEDN7dOe/zGAfkHQIghm6nD53+V7bkMc/WFv+hSVPAA38Cq4eips1Y5Je0
O8YK45GaqBlvJmlZJX6a5FA/XJdNBHJD+6FRs/CasnJLh3p3mg/cuBT/3I2Di+hMHQvzGfPSxvGR
dnVVkbhjnMTX46mTQZ24N/0njcUHOqVJqOOqazsvTQd3R/cevC3p+rX6YwDVCh1Jq7Y7UWjR86Ha
VmGVi6yfdg84MR4GG6DI0lY5iFe+269I+FZWci/b6SkTNMkyOd28hg72skJMJf2BuQznwEvZ7fp2
Hrda02/TuZ7Ih0h0DZb7aUL4/lEO1iJBCg7bJ+3qyXO8pfuC7Kj6CBWg2UInDuqwoNNwI2MammMU
UeMJcTqcmtUtlmKlGk1y36jlfNBhm2+QxpWQTUK7r5VeRTICEm8jEJL9FPIzTXnC1hVdNaPzvxRK
RAIUcGCX04MzxThi9ehMUft4HvLZvcZYCEmrEpwt/3hIQVVc4CBwIZf4RdxbmlbHUqF9+MuSuYWp
qx6WSXRA4zaPpN/U9dhBSVT5paoXm3dmIJRHSGP7SnGH9anl+tyQ2UvDpauep/TnWF/2itPxGwf9
T+yb9RKdPzjyKJk1l4bcKjudDRH+JMEarSgAFEY+pclymLTLxnWJ7CjIxxMEFEagl5XkujOnjqUD
nCfDPkF8uPFH4P0mUoul5kN2BGm1mzM4fd27HazOW8r9H1Vjsb9IV9f2M1u+ixv441C3DiOwjzu1
Fw7BTyLaY8GfTl+FP6rHnvr8Pp99LsRwqpIanrwup8XiLanEDAAPrrUlyIRvRajBtzkx4RkUV1e6
besIBr0/8cFtgtec8AIsU15IN7WPBV6CEqQoNUBUyYatMDATGWxAs/C+VbqCdp2Ke2aZWTVVH8of
fXbljd1pY5FRFvdrPHuBnRu4qsFuUuEFE/7GtNy05N6mTqwcs03gH6C+gnAHNzYPyugCIFlEoetS
+smV4S3c99v7op24efrg4yD0vBpRZhoqGYfvZ0pDkBL422UPysZPw3fk+iXclEVlljPmUcOY9uh3
/SHD/FO/yoMM2KH8Jx9KpdTENC+KdJILgrRL9qUYa9hUoKr6sr0+hlEGoc+w7ms7NKvisLDNQ3A2
ekrM75XigoL30HiCc5UFYwodJqemn+eNJHO691ChvCwvWH/fmksNESzTlV1CUygn5wh4RmyD221o
MiEChudHlH5UMJKDpvaTmx8mpLgEDPLRwSd9gVVQh4dH8LPm9+txjpoMCQv0BGWQpiLY/jSlck36
TjEUI6VPvnR3QFzfya44+j1WZnrzwkG6fq1y9cxEYKTku9mYAk2N7OiFESJwJ9is7WE2kLlUOIOe
8hgWChVcv1O8BbD4nqCXmWTHNMP5U6ZtC1nlDZEFGxBKKt7sK0LTFSzI3xAj2h9rkkjknP8cJPIl
KBjv1JSe2c9sWTAJG4wKtwekGgVmLCO9U6utActbCzlnRg8EnbHD55GHNOVUZBGPVvePmhSqoE66
D5Bvuk37+NeyCHrCf3xIlCZ7WpyZlRZiBwO6hcd7832pP8zGrvvBWs5JVsej1g0WYAZTGBBPSYHL
LcHDJqM9m8tJH+Szsi1sIGx6iX1JcwQA0iJzI5nBgDhZsG10lolzewk3v4gjnmpx+BzO8yjc3pXO
0Ov5+66qIs02OPtdvxs7QUVrhT6MWb9huCYLAfk8rkRUfVhHsIDHoEQr7RFJgpzzlB3H0Fq2pPlB
Kj4i7AmKa3cRGvimaP2j/mTXRmG8YpQG599EalCnnROktgpk4CXmXiS7ETenKhy3xJKndktY5Tuh
1tjsMbNEV3bLdzufE9m6SfGQ45eIfjxoyv550hzowkByFwGcMAO4stiroJx0FWHxC+WiNN1wtXlI
u/yePdRaZzkZ+gu5r86Ec7X+QHTRvDraZNv25MFFRKr+2a1230GT8LOdO7MfzpeUNV57o/sXk6Nq
G/fDJKKTk9GDkZ8ysJDfmxif+MLPeqgCKSfXsE9AHjLw+lxiq7ZIAmShq5uWCDMtqP5eCTdTKP+T
Wxz9E5A25VWRlWsTB/y1OTGFQ+U89JEKjHSxbZ/rKpoE24Hy3Va1OQ0/CR9RAwJ0v4lDvcMXiOmm
cCoAhI4GjZcM6vXOc7VGkDANTl07qM+rvyPNxds188zIbX4gZn65mHbsI6LverqFiYv2OH4kEfc2
lfJIIyK3opJ76z1cwnhYQA7u3lH+/rXzzeFn/x5adgoxn0xbFM2QKUB8WZycvE5L6GRbGTfiq7Yd
wn1f9rV56MsdtDcX21CzGtyMI1TiD/xnxp1KRNhc0z23JJv1JgtmheQL8eBNm9f1F/qnhfh+EgVT
0ZYtPyVEH1PZCG2214StHaqScauChk7NsYl0Mi8uoW925+3zKaV0njw3PZyh0UWxe3ncKtfda1yW
6Uh+V2D3lh+FyW4eOC8ccoUY4ZtAGlPXTAOUCg7bVX9l8qEertCi2bk+XHd5h/v1sK4hYlVGU/pY
FfIEmthS4+4PDSC9Kk46iPDw732v6A5AETc9/Mop2inr9VfFtn+tt5itzCcXdQ5gzH6wBVvdWntw
CyRWvoJ+qDns7fMPEk7ndXYNGgnOLaS/4D9kCOHmhvSCSl9a3ktZPewoaZqvsth3yixgaJCxM5/B
Jq3wOQLlHYrO1nXBQTlL9Z/i4LYzCecwZvZ8L8Nx9EV36hLKRT7gFoTP03+/Pmfrt8BwkG4wgSPl
E3f76uCzyJvxNgm6VitPl0Qk97e1NiI/jZzJkXzxJeyD2D4vA/q+8Oyq0W6GIutB+ZawLj2w7JFg
bvoHAJT+vGtXpgg9qjM67y8FRnPa55uI0JbgZiADbs86CcrmSAx0svQjWnQxNsHtOQusILMpOTwN
NHJqybPEi9n+9NGC1pue5LC2xgrb2Bf/57naqk8BduFmxzzzyCPtLEbeCiRkDtpUkRSYXcNoyvty
SLKLdz+gy/Pj4DJq3YlKgEVCr22YOxmTp2qR5LNvPhvOlUSIty3ukZJICAQ62vVANXWgrTYKqzWl
x+/gh9Fb9FKuM2IwdEkAkebLf0KJhOACF83/FgyRC8jD5XRf7Wk37NAgRxK0SU8kl9kxVR1ygsE7
9xvObt+NuQP/lT9pyuxy/+2F8/wN68a8wwCZibva/E5/UnAW/c4zNEpNwA8c8tujMhgo8+x5xBnj
cvXChppLEY075gIAvDogslTNiFht7C6T5TediR7rJyq5aIvl5bl+BGzrAMj39fWJLxjLmFV8uO9s
NZzbCYBke3TpyJWHfQfFL3i2hjU+NPiPjuS81zg+GgL1UU0SHZ8xQcvVkME2RkuFacXOZd1GBDMk
dpuxejifKdFrF7GTlTcf4EYE7To5PWpJWaotiFoNFck1lJ8KYMxhzKpL4eauvyqn5q0GS5kcT/5T
zwT18hcD3pY2ZsOBC0Aq27dXSjyw0xesCBMVWuFvDMJdTqpfv7Rg3ZvnX7bzZUSw284smZ8ZHBls
hWjvPkUm6RfaoZb3QFvU6PnTOrz7d1avvtl4Hxm5ryYQ9+TFVKiR6hAGs3XdOyCv4ux+/4DYkKHS
b5QwUqWghdn0fJgtLKyGIYge6jCrgzPMRLURLg6K0Lr2+S/f+EKAY2UsaW1Q57bsV8mzAtwCjLnr
vXrLQynI3gy+MsJMrGo+JAMNhib33uqTm9EXGg/nkrhE8Cdg1Mr2WmuutMF1ClPYcf2daXXoJl4z
IJH36e9TLtmKYVSVx866HVPRIVF7LO6bXkV1HQ4OZRKByrOOn5q8UN1vWZcc0BVkgD7ViA5YacTy
sD43UXTtusPgtxfX2GsZ3OpXQVAU/BvE16CIXSCqfqmz0ijBgIdLkgRvhi2hKsxp2H7XVJYim4Fx
PrUdn0DE/ADwLCQIzgFcoDjf3k+GYgjEEAa9/IDXY3StKIF9TSGvqbn7//nzNsIrZ3VUAfrXR2xu
858lTS07HKk4KwlPEzIkRgXNZJqQL+Lx69Gpn2yC5RPBscA8tfTlapWvASMOaZN1uSh4agKPZQc1
7dUMk7T2r2fhxfla3eWgHxZCgrmbSXpAuVkQ4TX8laCqgaCNop1MHgOk05nbNEcfqUgVptu+eno4
v5paq6CR2b3rY4W8T59b37ZPWtznTw94ydSSzby6oXLOiM/3BgKVMoo9wMuZ1Fz3gkD7MunnD75M
+dszu1AB76mP62ezFd19v+7syDP6k0w7CEeEsKTg30F5evX8Zq5PT6c9P9H9io/V0mlykE/cEPLH
HVxMJGcSJUH2sTUm/mRCvVPw/3ERmOYDSygRSTJSzze9oH6ofh8uwj30c0LZEnff32vdEOaG4e+4
IYu/i1z++uX+T9qzfodRaAeyr5CSjp+rV//ymuHB4r8TJVoJR5lnhpxXQRDQnTlB4R4w4umtQF4x
GLaLZRlBzUIoOJfMDoVWl1W8EiJS7KgqpjGhC+LTpFyxiCxgh9L8m0S1H2NU6sdzuUGhhUX0R/AW
9Hk1vePUjyhTGW2YEzYmHMWtrFfMKGHATtIAV5pOkcGqAjAxONQx5sy9D/Ssm9LW5DDEJm6WCi2G
4p02kgPKuiAsez9VZgMVP5O9azEuDWrHPy7n7ocRewdb6pDJXxRcLluYK4RYwl6fvHicvzzwLjsQ
UkuJJ5pdN53uMojoD270w5nl4NO3zB6sPg0PPiwNET+OjbGtA0fd6VA21xIal7zaQTKJFWWFo56S
aKX12OhGD+lPOmjpiQ6uD3Q+/Re00wjBYgi5EOHfYKWlS9YeM0CL2CHCT7zmazbI9Kp3lUsp0RL4
TOylYuFoICO+pfiQLatpk0/4EMmWFezKhSqd5wR2R4xqA9jJtGCurBKOVhozh+S3cmqL9YbPBDkG
kyWMBopnfHFoh4bai7Bj/OSS2W6JonfIAfsZsf02rH4xruNZiKaXMaFm3E82fCkHmgIJ0jnsZ4pC
1Mg2Q7w+Rnk5XV3fGasIL+1xuOhjsBTrXiBuCoIabHEPIsU4/MbH91vREzZR4iPZ0Mc1CDosjE4P
xilVdPlAiO0m2O9s4/fzeWI0FoPi7B8Yi6ChJeKfr3N2oh/7ZLTXh69lxeVj+KQ=
`protect end_protected
