--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
I1iwTj8p19/iyV1Kj79i2k4YWYNpC7jgV5Mg4HOSLqDRqgurs4KC1S1WAz90ykG/sbsW/9POs8IJ
3e3d5Edp5iGXX+8NqiJgH+1o+KnVjccwIYeazIsnVozZt4nm9FsVWJLEb1T31uN9ALp70HYmBBw1
0/Hh8gNw7QJYFGA02ub2io9oL/FEs1jrxhv5igTpXKsXyCYmQLPSPiBGV6j32n8dmlz9g6+kQf2X
zfQwLSwHbdJdxsCwjOGpvHSzmAfaWu9cQtMW5a9rvp4OaWsKCs8vTDVJiuFS3PIUmoqxfIM623PL
J1+bsKWm7me111YDtoc9Zd14rfGCTaOxmdLdBg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="dTekUyjhHaE/kC+qG4ZmvrTlWh64+4wtQNmunULyooM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
iaxSJez/2z3oGFmh6WQ0a/YXJfcFQ/KPJxM2S0A4c9ffPy9gRtOd9hzgbC3jzI6ETqo+RvuxDZkS
cLrjoJX2dBne7+qw/53KRrWQQQZDZGAmeDIiCzHmKJ7FBCfRFdQCsUubAi77JgYQnUirYXQ076N9
TQ4ltlIcgDNLvJGWD1RqsJ7pCq0DzDf2PeF1BNGIoSXbz21VPJcBqcPjIAa1P64lOIMmTvNw3UtY
RueG5LnP6b2aank7qvr9C2CwsENmwG62nboguwLI3J3Fr3tB9fuSTMh6fO41E65fz7jv0tAgGTHx
dBpARHIWQfXC5wKQBBuAYq3wtHycvTGlELNmVg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="jrVuyBc//RFskTjnWlmKSXYXDKfVvkLQYiajajKWgJk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5040)
`protect data_block
zX2zNZyJlHQqgFcxwo4d/hAn1E75GpgdCOmb47VMbz+KtcyVCAAPTe/04nAgBqZp0gFIpcsXSsco
zCroCNECEoUFxPm1h3M35DzP82bHFDHcOA6AmhDPO7+q6/OO+nTO4Wxw3U9h2jzLEyud1nFBjN3L
oVq48tbG/AnX6bsOjQQ4dEWkneHM5TA7DsW8OUclL95MmugAgAp38xnAP6Fizew2dVPp+AnLnZDo
LjMNKpo+GeLNZaPbyy/49eDzBGim3IwP6NevSxUiEZjQFkwkCoTn19DJ7JlmwKbxaNS7HBPkxDRI
Pl+xDz6CZigTJ2DSUwTTqK44PHUCvAcgIRAEeezhcnz7Nx4gaACjp2VACVyndKnAYx6bv90W53JV
PpzANVnM2Bzx3DZH9yQ9aq+MrGnVtg6/b9FTfLDcAOf4YGGT8L93s49GJdRFauJw76yYM8pj64SS
mFW7acE4PkK/xD93+JSGbH5WxuTomDBbtcySsvbE7EeBvlM2CI61yliK5CZWOXXpx/Gy3WB4obvT
WRUzMRT+1mdxVOzwYUHGcMmR7+q6T/u4knRd/IqqDtulfv6JCIpnwCWw0uKuYK7tFL7tX1QrINud
Nu77Nb85TLfuI3lfgM8QkAt6q1cXBdYSDCsTz68za22V3x4FdNSNrJrKB0zAmprTQ2i+IHdciQqu
F/V9+UyiK6uvmapXIvfUzYdGO+cJRHzwvIDknJn5q8xY7rwmueE3OhobuVBXEp6ipzNxnfCupIm7
nag/fOJkyWEFJTCogC9GZDLq2SJ2eIbSJYWPdhSoEioDVqiT5mvbouqshMEhBryCG1VlEfQjhWhK
chkMSrJKvEOgVqNavsyNxsWHizqo6GsoCd2KzzMwGOJekQA66GTyEDP58ziM1feAct9u1XjZMVq5
CSZ2nU+aiUmuWdg+MZUKOjoBssxVUDiZ1rij7T9Sx3zWTnloAi+U81LlrBEteR1lLIIq4lyJMjME
Ay5ZDqLck3ecbkdx6Vkm4mU+duqoKS8hyMMc5jSj+xzYX54k7nmY8kUwTwdMzIMjs4eSJETdVp+c
IQuRALH79yGYsSUUZLlKd8lP3f68U2G+Qtp84fYj7JhyYoWYHVYfyeZRBY0s1SKU0GZ2zN4Lpiaq
w9NayZztGyttUwwynmag7SvcTUWa6bjggKI2L72Mqms3bvvziJ7D7nE7aPxrb97lGx48HXgHkW6t
x1ZOvmiVHCdLlVWid4hymw9WE8jwYWo4buXWOmkiZVxF9ceV2WM3P+2xqwRUm8RBXBwYwSHYupNX
IexQO2Izgdpsf9HcqfHwNaQn/HPxqJqkVkd5uCcnbYyyjTt/EU7k2wIcrWvmm0SSKANj7Lm2avjl
jiWRjF9KVXPjt2JdmvBBKfue9zjcpilCsr7PNv5djLP3UF7O+akbXf3DBs2Aepzh4+ysvypV3TVi
fME+h7W11dGCXmkr/ltrLObWYsTvD4pSjkqmApf5Tjl/U3KJDC60n0X/pSz6c5fC2Yc/OLuEvlkC
dIoM+yztB2JCOjRvAx0FwQT9v+8B0n8BTF9e4/xwt7O0mHFHM9BdIn5QDdA62CVuHezPEWS2mH9t
aDPF8Bv9nUdw0JuEEIGRXqwIALS1LDmYD1VJVY+26oKIP0HslBHvyfbZrI5aiU1fo3LUmTuuTFWM
kVPYYCvSrX0oTcJ27kD1eOlCcgvPJqeN9RUrneUmRNxSJr1P0j6+sRTuoOederbCXYYjPgrJQ2lP
EN+rNDkLvczDEOoLYGoplJTeQmULaRlsF7cnK1mBHb7nsgQKnYpAj2euM+k+5ebfAovhrl1uoI6d
CaO65PbAWd2GYWAR8wfJG55bEnwy+fzw/emPecf6fZbKdn5WuHE2DnE22uQ20tsr4rxXVLHFlO+J
LHGvvd5+W3fYLyuWd5tcpAEUbLJUs3L2KTpT/WRkLig6m6fnijYL8Nw5DChqNEukKBYhbRDSgPve
Xm/ky8/CYcpX4N7re22eCkcOZ0q6xfy0NmYoGM3es1KnaMVLLVjjPb/UHOaufFLE1anKnjyTD9o8
S/hFi4L5VR4/Y+SsPG2JY2QYLFm3V/CGrQSdn09vgkIHFagCOilGPCXXmZcECBAVZ8Vx1DlhKO2p
fNk8IjN8Cf/uV4ujPM59xoKV9hOs2+QK7gIjDfBws8yRff1ebH7aqs8tuKvw2NojeFuCwUZAfWj4
jATcp0Deof4oKa9khSulYZSk3s004/aMsjxaI8srn4gFD4uCSl2mp4Zam12k1kVBEKyqH0tr4CKM
oeZyFItAG/KosjVqsBvUthWrPCe1X4/mQG91HnDqg/sApt4nPyr5Ov4soNy2Du5rfYWVZfI8tICF
SgpSRE017yXJCfe5H90NWst4JVypb1CqndQk98UA/NpPr47AI5F4sgYMkpCP4zaOteDYOxUcTak1
WUqri14Nvp2M1Hj0A2jrnJZ93tUOcbRSZT+eaXgVrnGG5EXUelmmM07YApFwECwsCwFXVgSUz2J2
ZFd3FP95BICogOPW2btmp/KlpYlYcJ2Fa0im/tfv/4J6QQkDK2fgrf3USqhWW0CDnNHBpw9pdSE+
zKVPLQv7BCXj97L5buBap05bawu06PonC6BAPthWJYqvkIFx8ZrF4IB96+YeC5lryjAFy2mt4IE1
O4FPSILk3nW1o3dOSj9mshmTuSGs1K/TrEiB9rkKMLMa+lhIHGVx5TvMxyNUfk/CLPpv/EhtNl3q
kPCtgxf+cmgrOUeqpfB+NVBbf08EgaNyI+0Jam0LYkSmFdEEYhi+VsCL+4qZfLoFEXfeVTYkAjUQ
CYwIiVe+ZB4+kQ5JOHBfCEv55SWaFmzMlUHeA63uKtPk8HEfqHn34gUnaP/M+Labn+NykIbFM/1d
PwqkojBh+uU4frnF8krbnSb22ZO+mOc2oppFRjMbDUiJ/ngQ3vHeAgQdGh5EKFelAlTx9cnGBgI1
5DPGUCKnc3pdaxg6KcodS8Ck6SAPj/Wka5N9RuU3Y91C4IaX3mYQhbnitjpRA59o4ivs99ixVSfU
02cHiHvu3+3d8bAq9rIN9594SeXrNiHb3U4f9AKKbsmKA4RHYDSUv6Mt14JSCpNVS2C+CvQkOH4a
V9zIKW2A7Z74x81KYg3G5yUrOv45zpJUMByuiczQdThq55EdRnT55JfvQpV1pE5AJxeyODzaNOIP
IZsNRylKyKkkdIkSYgf/aVn49Bk1WZrm6HOEvOgwC/s2Ks+nIr5zOBRVWOjz8dAafMo8HGUyRSHD
KNLbWYDysKZw+v+YuS2roJxUFDtgmKbSPWbVSd/UJ8gLI7YVL3cv7ZBxgac1VMMwNi1Jd6jyxK+P
YMCCnLVr/Foay92zeKqc0Ax+14+Prn3kvkT6W1/eAdi9UvF1q+1PM6hunsOOa7xnDmzMAE8g9/nt
n2I6wLBPvOYjjubw5DZgslMqLDbuVea4Refo51Tu6SSiGKYC2ZMTzXH/y3xghnktS2QbbgnMbAGL
6Ju4ZzmcBKjWyx4A3U5V4+PGF2nCQVKYK5fXjSLWjHYpqpIGvE+tvXZeYQYueINKSexN3IxYDrSc
lXZsRfhPqW/yum6tFuvjObeS6sh6OOo08E4ylGdTC+SDBDsESNg7IW+YqpLUlcIKvtpBZHprfX6b
OdtU6YZKf9P4iQ9fvztQytVUSrd7GdsZE1dJhifqSkYYwFnGEOorRgiXbsjiGgrz1EHMN6f1TSlw
LacS/uNV5Zf37YZOOEXGZfxpr9HDLjbmUvqf/sytVdKs/q+uw4yZhdPGs/wP2oYvSi8fabM8Ik4J
lWvZg+6WMCaBOm2zAOyw34clozzA+C334W90pD4Qihq9E4qF0QEafIhS5XPPQ5gO5N3ZLwAEzelS
VOLMXpuDpMChT7EC9c1cLvXZY0mrGhml+YeztgVL2DmA92fE9mih35fjq1FatlfuC7uSljqRKKfx
pbOeGHGqVUys9JGJmAt1KtxMecHOvM81rb8F7tJlg6yiaOv8qC4FJj8jZweHbpLerswKW0JPeigO
ZWEagnm5RT4OeP+wEJk6VYyA0ONVWcdILvjQkNPGVmKkgb3CCPWVWaXCXQKTjJLlCz/98caRImYW
Gjwb2gPNiwpIu/kez7ZKL+DyJGIvTV/RDVWpCALbkKqTc2IM4tYjt0Jx7qiBOziI3kcc3Pta+NlU
VvpxjBg0Q2er+vsiFtczeC3VB3m5jqI+44dSi6yXi7BzXES/QTMteGBsp40QwUlwjrOltuE9lbx0
OOZQSLoJEqZ/GzHfvyWw/7LY+f415Vir4FK+tDwl1oeOQWZLcgpAqIgq2WXDf4JEDKyw2GJ1WR3W
RGB8TB5K6QVZ15GaR99hk/KVt9GdaB5tpzFONhULdtPBg3JgqUb/Rns6ALLrLzcTUQpMA/mK/Ur4
/Ra4jdr+BPoVR0yMzxxUQSs8Kt7uieIHjCHLfxDPUhXXBnisxF3B5JmvBK2lkUTImc0NDMc2quzM
EvP+1AmvMoOm5DEwHkdybIqr+OFxfJG63La2Vm8/1cIwIUwAgiaSIu1G/GDCHMngGv9fHaK/BZA0
/jv/DMnYFnKBDOtV7IYeVUx4QoMNNNkIW7mibaEm0CGlgcp1z11L6p0TBf/b2hKFbm4r7vril097
YRM0IQ3IJb2wO2MYBcQRZCZ+unqbP6a0mnLRApelXSJawuvVxk4jH/330y4HV+MNRFSiSOSNTu5U
nZxyFxRZ74bRF6Ec09isO47B2Q39NhNidJ9hn+UVwyv00Jrzzea/r7Dd1uOuNyftkIRNxzXDEPHh
izwweKq2KoqoHSJHlHljIaTD0Ka193qPmHkjBpyrKstONUUKIsaTN8A03GYxA2SwlSGUpp7WQba0
0AfQ0llWrJ2AgkCBEcUyHcMGxGksxhjje4WQFOwfcBSXAWjsto+Ip3Z+4g+11RdwpDKB9I0jxHDN
aX6+fX7k8ENjxbX7IUwxm0PilKfTwbTLafdT2MUO43k0OG3V581EbOCKu/39D4BFzpxbAtexulUJ
L1OmnLDM+1PEAiJ053d8JOMfOtyDiABh9tsn/OfsDIhpKysk3D9hMoUA9+YMoCti8Mm6iyBPscrA
MVawKGX3jYCKR1I5KGifrGNmwmV0/9OlcXHAZ5pV6md4MmqYLswA78bvgT4hb/hVWTeTz9rZBJ3A
NQxOAgyzHgnVOBqKA8ngBLlsgitjZ3Xmc7ddX5HbW7dz4imdloG50TO7/gMMmLbBVJKDaBKt/TKJ
nZfHk3z14FfJ50G9+mjwTcs90z1PdzOIUzBPVFJrtnw1ppO2n/ft5gq+n+up8Gq0OK39MLLWYIKx
l3ewjD3eEYSz5EtWM8fs4cINFT6l6r022Yq/sgCWHkYu4yOLPRekx1xwuHFkwIC7Lm8yAbw1wqU0
Hb1Ypsryp1WvP4QGP+oAPlaam7OS4anHmfvixYy0Moe7u/pYUcjsmy18Sf5q8nOuEqUOSAtkGMyA
FK34pqROm+ume0Oo+jZbomtbuu2sKXKR9WFfK0V7Nt2QnU9aSPlCCaiIWYgvA/ZogIWdvp5ar+57
Eldun/uyWV+n7+CIPnvnex0K7KsPBo3RZhCyiAIgIPUM4TVN8Edfj4Q0DB4mXhojeig7XKlkfSwB
oIgN6MbM9bbFT4saFYMJanHYqH3bJC689HRjlsUtXmKmL6CEkPA1awT5L2MugWyXzV1yqO60F47b
URoFqDBEpek3iqimHDrOKZMQGXlBARKsz/NdNm/ZWMknMiKOpXr7KuaaIlM4fyv6XZxxMyamSzD/
RVX5DjYIdmm2HIJ1FmW0HfE9RPax9VtfGhx4kELo0NVGi9o8bwy1zAspUC5J25ZJqkpvVeux/ayh
3dx5IvzW1oDOceF1xmmxU1JaCaKu4hpnIeW+Ywsggkfuu9wdYNwmMEh9/ApZwQJRZ+6I9UeWWUux
A2CkX33JFrA7SMRTL90rcdQhSSkKPzGTNPIIX53WECo/m1zdnSy4uOf0diBgZWeQerhtPn+DQXAq
K2B/psNyjJdmSsymu4MeehTIUrDQXKGT6vKDzz5ad5JBMP34Ne+jHPpKU9K2exBzeoC9DbdyqiRG
CSyrYpcVSn8XrQw2hQLr0FZtW2gLfrG8+SykinxI+2o07M39hOoMzqE5BsSUebf0ovGRKdX1+c4f
QlLUYHgn3zC7XXCpshHKZ3NFXXd7cQ1EZD+xUJgcDVOaLBbfmxNExr3BUv8Pv8xz0+PsZBRPmKTL
lGLd28G9uI+oCcliSYT8vo8e8tlGUOtb62mky85fHPaESWXZEzOaJlWj/Vh2Yw8go8CfgWpdVqTR
WlMqdNJp16K0ylQttclgzMqcwYDQj0lUqvF5JSiraYkGtdhV38/ewGqjQ86rFa7GliNTH4kohPxs
CVcTDTFY47M88gsFG8slC2hRoZHzI6k89kfhBo9f/8RLiI/E7iH3ioYX/k94Aud2nca/CdMq0a2W
eu0AQIN5amHfV6Lbz3+UvgnPWtkd0iUC1Y33RpOiYh9u2dNzxQ8SaOVk4YgcX4E1Ut5QeQdyhLjV
H5wE9i+35GmZDvxFu4Zj5f77/k+CIZjeh177AuXo68dudeeGD2u9V6/t0mcgYfoZHbfg2KWqWKqm
MNA7SbRzibUYij5UvTBtyOpdXAJyS4yTf7A6hMCLDp8RIX2tpKJ4KnhUxvRE8IqNfy2CBqDXpwRq
oAKDoAgV0W/6Zwu/EaAOrH7jTMhLbiUE
`protect end_protected
