--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
ccYv/KYKKCL6FqmlkwmRsAI/s93inHPF/QiXuZokT50E631ZUsHvX1nWz4aicYM3dncTAkJZbW3H
e65Osk3ajhIdMY1lnTR7y6xNsB2HdIH+h9bwesvVZs1T4GTpSUsdhRR7pc6mKL/nc5m0ANwwNHPq
CHP1BU3Q7Jy9PXgcxgOF6LgG95jTR+CSRANiiszueLbas8RKcG+4D/vfAtHzV3Xpr4GFfCwGW8gv
DQYJ/xoZTgXum+LepERlSndNKSxNEvPuexYUPFGbu+zDiny8U3jBNQOi8WnnVqENB/02OoIswpoA
ggmiyo5ARr8VOpwBtI2VQ1VXC7ZcKKFANEKF8g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="ui622MwrLPHV9rf7NYapNfxa8O5xWHqjByhrz3/PZ2k="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
hT2G6koSwTaMd/3T6SQjbRWnsN+rRa8jJZ0h9SKF1Re7wK2bJ7qcLK1ShcOQkA+84gGQsfk7Hy3T
7Dpj2itWlxJZPAQqK6ajyTPnZq2JmC8z2VUDUuOeZTj+nLpj1v6EmoSHrt+IR6mzbJZ+B/e789Zb
g/f5rCoMFpFxQXFyUAcSbAYLZHB3iNQLklSqUSHVL5szhrLISYtBeSDdxZk63cPgeAl3+vrS2i+w
mEqQL1XIkUUfF1QHHOJtyWBd0LXXCRyVuOZQXv3rjl1UgmVgTlDaZEoIW8PINRSun1NniRBzKDvR
Aw3XNrg4my2K5tn3DH/x3PyCWAlJmLZJ7SLXHQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="J4OotYS6RIv3YDtr0K7IgqyTSCxl2PPXICroOp5odBM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 29280)
`protect data_block
ww6L6FNmcphETDO1CxW+v+Y+fp6dDpecZrxp5wUzRBURW1AsFK7DYDFspr4v7+Cmyfq8/efhFsea
wJOb3mUxZvZcwFrPjNDBtToJMMWLkVSEgbSyMB6e/6TzJu5b6L4MMYqepbkJnnY/DqWzk4++kA2X
8hPA4YZq2nIo3b7kIt92LjfPDO89UNj/AAjvJGu8k8kii+g1KwpcQrPJh/P+CJbJX5H7qbNrc5Uz
YwjTgX64kSuCiqGtJi90Ka0iFhUJgodrDP46yKaYyEEjdHn9q81KhPI0Rs9HxS1ocuqGYvM0WIG0
zyUikmY0O4oNxz9QojraZ1hf8NeEXbYsZrZpFuOwnEowjOj6HkWj6Ny0NE12qzNOgJ3NNM3CMv4v
cNu/VxAKPWKFLExzRK/aAybO9N8kIAUgEiBMOc+vYPrfZ/jmf+BUkoTSFVgJ0SutJAKjdgvVzE96
zd4Wo+DfXGk0VqFfWXFsUGR6Yek5dyid1UCdfaMcZhi3rlhSbNMPbHJEwUQg7vr77J8IZ/fNGAeL
K/EleSrdS53VmjSZuLecX1+Gpi2m6nH/uyqJrzL9SkCkjZpwUW90Nuk+VnxlUMtiGCMrukdd4tIh
+Zs6YxOEJMJ2AcNrSFObNN1jaNORzQtE01UOGxVMZ8X68YuEYpeCHVNoOrG85pvQjgNH+QkCeHlT
KVetBXeJ/xyWM6QRcrIrKr/Zy3ZgjzaME2WC/tntoYlkPE2hsQ5xFHCEH4xt+rHNiTzxqTRQa8bm
LkwTnfVZ9hBc/tLqGh88S7wfALWRyTXJelmHXm+XMdngSYW6O2NMh7Qyjht4mfHRUKXYjmPYaz1d
Y0FgTUh4IkyGiq7tFf93+6MIU4rhLO11MY9GrR/jXUznJdoIU5yPOEVPmNeuEXIBhnHS0WLejtIg
frgvSP5ycjogiSj5NSvqCLbit7yhcyPXkrDzh8tRnv3pGuTRRLQ4AXRzASZ3CxLtlNP1PLtsL7sy
NoD0oIuCIcpUDB8hT4FtCmN4LeOmn8rvLdkT4rZkT2TqZb+XlOIKrWPTiNyPElPHTIjeP+0ePBfF
xMs2/NqPlmBJyUq7buyd9PkBtfznJfmAaB6SEFdGli9c0ktFISnLWP31OKFt6Exg3bMKqFv7Swgp
zVctvuOjIOlwKBphCrT9K9XmyIQwp+MuWQpw+UDT+pTGdWitf93kTIPdr4uQ6rk0xcnzI/waz6dJ
GMR6aD3sy9BVywvhxMlmPnBVyZABkD2PN2uwzngWIho0dtqkqI5iwqM/MAYYvsME4AW1oD9RqWe/
/bevCYVJAJ8kPDnCQG9pBDR9kL2GOZxs4sJZ0+YgTHNUBSigrQ4gxe1G5jBMgsbybXPtm92fDypV
zF9CrHrPYNjN9IG1fjrRWY9Sme83l8p3WVRtcKc0elgQjnWKYs722taq1nhpVams1k0abGlBk+aE
roXeEqLbnBC2/+EunDdhpqtOWsvYfF/8dgL33NKuVvQHvJI7qfqYltwic4vCrOOaWBe8HZnrYJ7V
tZcG+UEGewmCSbhTaRHsxj6Pr7ovTlzTY6SxmOHo0+/nra8wxHXlwa8E+UQakD2lZ74Ut1/fzYgK
KXgj0KITT9bwefxyla55gH1wyhchR/PtO1hQ9V5gCecPzvEgVrx730GxqECvAO/HNaM3pp26kElw
uvA/wY3eJqGq88TGJ1+zGiTWKtVNOfEL66c2eTvZRYN9el5d0CYlSRmBU6+KvTUWduEjb3wmrz3k
Ik3BBXrkthJ1akF+LM6I1Jtm74W7JkoGoBwPBTrVdGa+JiT83zvuZungx6xXUuOObnajIexWhJxk
yrjUNAbLaA3mQQKkvDKRedevxhQPd3D2oWZ2mw2EbSJsXWA6jwlduufl+uhYKQJopCzXj6KhDAEZ
Tg3vzVrbkVCig/UC/cjKOKUs2THRtPGi5CgO2Pe2VmUGcgt2MLtZV72MTMFGMiLWv7uRHtSqi65d
FuJsDRkzpvSqCzEbLpfHWQlTTxQDG6y+OBovTKJcmK6JMMO4AbVrGW0P21xjs2EIpMJnLhaNjdAR
qec166XO5M+POoxK65BBfDytGci2EnywjOs3g/8VIrXdaaHOzf1x+HibvIz0z7JT3tofPdVXkaTn
RQvxgqqCyi34hi4amfacLdZK8/BlgkOk/GU8+ATzwGA/c6iynKraLgXY0J4Klv1imJUbJoGW/MOv
D6vu8ty9SQvmPSnJPhDmTn15Ys9xzs9DMJnmkXPOGKL8pZs81Bevv7D4pXDDs4v1RVsMhjTHxVAs
l12vjlnIAJxrzMdw+Z/PzVml3W5r7tbg2ZABiM10cnzZF6WICQc8WidcKDBim5Pzsjd05sN3AdnX
PUY/djpdRtI84nz0l9dO4e8snWZaA5A+k8m0KxLRkJDsNM2V1XTAJ4V+Qe4EArB9K2JrSgc85y9J
99+HKJgR+rxmnypj0gfY8lJy0y1gUU1/kCOUH+1/Vi8qLg8t+5OB1ybkbhS+JVRuynVvU9l0y92L
CNiHxoDn2mRz7R7nQoB2XPAFQ5sjwhzkqJ+rVMcG8V175NcCBi4T3YUv58efyDrCWLzVPUGGcev0
vnA0QuUPMhTn2lSSCX5wrcWCDc1P9VZRRU91dQH+PEPS3CbWyCR+ZCnG4XQO4x/43LEox2oVZSKg
6fj6k+NZE8g7BXr472PZLrBo/CHVWBvjPonGfSuGNbH7TP3V+hGGW3JMI1FxKCkBHbNAxen031f/
wdFSQ8wXLmLuUL6KowN1dLSIVZvs3wZOIZZ724eanc9GJchYM47GILGVhDnr8V55yyt1h6d8wUb1
OXnw7B4qM2BCYGGk0S5ruSIKWvl8/u+Fp0qIz5lWZlsLyjfn0ALnT96sLvHg2I6ggfdXT0NPCIYV
1EJVuIxhMsjE1wAfZO+vGkFZsXIbZ86Aw+7eQ7vJZAzXYoy7bHt3CNPAUg55Ww62vHXtxZbf/8O3
EPAlFCcu6wFb1yMZ4eu+3SaU8amy7BAPoQ7PtZCwA8BI293OFolq5gffbXYIGP0c+O1TuTjqIUdx
Z7q5F+Rdf4QsgGzlVnctoHGGavmEEdmG5r9nsmKd7XWO+6zbL/mpxSOPpDS3OVq+6E2hBS5lLrbu
7WE8tORWBVCtGsTwIWTrNJzr2PSjzsonLNE8JvGd1dkCRmReyeTDAYvE1O5IzG2O1lm0OBJGgE0a
2N0S/XUQ+E0dIfZoW3XRXM3KFNoEQoo+SFqljdvdEfjFHsOgljQEeGjmuVVlwR0dX4KZufokRyda
NpaHzlYkPcBpBxHnavflJsbz6jueHLQ60QQM2+A+pcMTmCs7DROApSkAxU8y8u/gWREswXXawktU
bFtHN2m0yTfjSoRE9nwguTKoLaNz2lf42/GpknXb/pUzOkvoT1XSTAVamX7QWLKTLPsUmxbXoJqE
3oVg7DN3YW5Twh57B8HgnTy/goBad5srciAqGqYccw+qAwfxt+Wvho6Zq5dnnjL8KuDA99E082vD
XTcx7+voGJNoGmZ9b6WDZIoiZLM6XNJYoDkwQIieOh8jRqdZuyLK6eq5OGkp4utF4L+a2u/ciBeB
JZwSE3A/XOFLV8fkJcuRuGcp2HZ8ey21CLK36LfaIyBr7Yf7UEAAGBCwetxIzs0jp9+okz4VU0DC
IfI+An7xFCvffV5qA1ZSVSLvXxNCCHjWAUwudUazb8BwrIZi5wDtB9+RkQGsZYebeIdOV6+xPUt5
MYolcJTuRGd5+5dvYdU4xHdL4csbJq+5n5iqhs23D55NJNhSbDkXr5VZhs4LEm7QsYOcBgyGrQIq
BQ2PwlsxvbrJIHSF38FjNL1B9apYuagWG6bglxu/Wp8fI6s6rxrokaqs1REZZFPliS8hGwCuYTE7
zlHWd5sh8yBXMYbdE0ZkQwIY3Ue4Jp1qG/Sp6G8bYJwttnTRA8wtUTJFBdatDE/Pobv2zYq2Rj8K
IUJIV6Z3xsa3jABWJ1jvfPoHvkdJZ4OmAcHi5VkgstNBONuWeivv++ub6SN/pP/6enQfbE9XWnMB
P98phMYuChuTtl0cCAsnWYymzUpNVKvi12gcOJBmj3qhGYFr5unGWMxO1nLkyy8FYUamcjopFMCx
QZElfrLKlxZIDf4MfHUc23QUO5fldk27iNQbuY1O01nvgT9BTAl9PooCh6md6NW6dnzs6m9R5x0i
fdE1K9f3of7sWb194dDoYyCbzgBBCyzgFuGyJFzlZkBz/dvUp/aKW4i2QYF051o9KTgLUU22FtAq
WAxdIsYXvVy0aKTJyWv+nu2jpGhHo19YqeLZz9XDU2Jrhe2zrCSAcb4orpe6sbSpLi4i4obWFfxO
qQnP8xV59IQuV8T3neJN8oqJwQsVXxQo3Y2CceDnO5V4cwfuaoPAmcPejrUdcs88dElk4VNQ/dpr
5Rccen2i1cv/XmOx1ob+xLURoWPn8lKZ7r3bpgNtD5PGQxNysBd+VXTgsSgsyu4iBZkwG6PMo2Uc
/BkIw6cAjO3ZgAHlilNTs7XTIFrTgtaFXk068SwJtlywG+5TbWwHNiduFJN1HoicgwWKAwl+KBBM
uTpJgM5be7F8yxH7IGZlcGiscBOhZchPg4bz4OnrZf1vbOW3OaOh2XHNaNb4roPjtoxgc+UXrWSz
5c2x1teFZGdmogutDGjLe3dKwBUZk/Z7b8iuXkodfMEjpZH/1O2B/QvhLWsBEVNtv+W2R/9tTamR
v621kMtO4MoKTsdcBXzFNKmLKGeLI/VzTSw5Qz0ifw0bQ5NBzw0jYidW/IaAm/XkooYi8F9anp/v
MTdplHBYkIFMEf5WEKBNIZeovwwMiCm0FeZy1/+CTBkkGwrcau2jjIGg8SJZMOYHLrwXsRehvDQG
8CUWf2PIaWFHxJ1h0smWpKkoIxV2uW/dUJxL2AB3U+A7Qzsb4qupeIV60mNLIk0dEJZf2s4nnH9O
ZQXJQjNH84ARubqI0WrNF8ge8AOEqaLQpoBozuon8AYz/l/mGdQQAoeZcaATeld1OMKPuqsAjI+V
Tamc3PDhFex6/IroF6F7U2dO3rLfG65l9z1t4tN+P2Q0dCubd9bkJUcFqscVZouphK5vcxSS809T
eKmmkPK1Q0ouhvR9H3NuY1hX2KeACbZbwvVxNZVrvkorOSVeK12Z2qLpQinlw/aHSWIC+4nV5ofL
3d8CcC1f6jC1/OsSlP/Y2uy8VTK0VHFhfCE13Wea3iDBOU2knXD1QWAeCjmBOHDtG9hkLMm5a0ad
siogsA+oXnJ9Dtfh/MFHgnnzMIbBvw7h1ODi9Lm+eeOafVcetY6wPFaveNMuLp+4aT+HllN5QdDl
C8SKsv/LPN8BkfvMctUFTwru+Y1NdNXO+ASS3IVLe8mGmAJ7+J9kBSAQqagema6Cbm/mLm5PVrV0
7i75PhjYUBkv6EQ6LMWAB6Z77O+0WsSKgQFJR/ZbJ5LbEpSpPRzJe5Rk5usMf48hOgppkVQXkqrc
Ctpo3vuvbkPkeB50wOCOr/4ujAdp0z/W8a0+LkNge/mBHohzCTXd9G+esRqgcS9slYH+D47j06mC
qjHA63UFwt4vtrzprmWN3kS100PE7BuzMARLKwMFHzsHlF940YCv768GKLbInxSYj/snWVK0Vp4g
9QQveKaJDPSC3kjcnmqGyun8GbYxlzgqv+VhgWXlbFFlxhbDgb50mlE91IMt0hJyTo5TtqYYqbok
pFTIzWMvFsqPw4T/7trBZT34gYha/I6SBMu7bdsv9bCMeF4aIaDby7XnOgSo1jbRc4CfpCnUJFU5
HpkNFbtosTyQey40jzmsNkw7jJ1MZxNM+9CoBMJeJGUZuw7MmGKSdh8rDaarFl/spnbbhhR9pCuC
gck3EaltmKGnOCUu4sUk0IobG0QXXDDsiGmr1UuSyZFbxO96tuYUqRmOGPQ7ryweD0jZ/9FyUJNx
3aeWEWLbc7IsPgM23dvZtiH3uwh1UCrGZe+hgEGFaVmJG4NA7Yc/dYPRJYQincutqpm4+t54BjKs
FQ8Xlvwgpvcwv0chVPsgTCRrHywELkiGqbojsYHPwtLte55/4tjOl4qSr3V8rVaE5SWF0ycaX4ic
ACKyBZG3gkLRa0bVzkg/aiEHMfIqbbE6gE7JyfW/BB7yjlDgohqFlyV+FiURcVSQdfgDdeQ234bH
AkSO9cngAzBD3/nLKXhix3R9yAJRXGYZMQPEDY94LxnBa3xBklAWKhDi4lncPBb9/f0uwhiIEBik
Us4amI59SJPuSBefa6JrpnnY3RdxAD3XHLbZW8RKV/AeHvU9nSzeUEo4y4k4dbGL2yH8CKNi/sa2
MVM4VQo87c++KWvbuug/xwaoa66L/vTW+iXfawZP/vcb8eKx+VCeiz6qwAJBSA0hoilk05YM+qFB
jS/3byLlyqx0APxBw9s127p9CcJCs5r1Jj8RfhuYWi7f6DPPHoLjHHsLR17+jhkeRS7TH5Gw3AvU
wXt4FSfTGq6/Na2s+pgySPAlf8tkAC/zS9aa9KGcC5tpo3Vm5sy49KDXyfSuvNxRT7+hRs9VAump
F8snBKKGEyUhQkYOuKklYJXRLETNQWNK1uR6IUd0TiejGthNagPXRTWlf7CYY1nHAGZakh5SIUd8
xiB3SPHDhadJaFc1hMcbSZ/CTZXUkYuRyeK7ai0Wx3jjlO4VWc1Z7DHlok6ZiZJIAi/vzZHWTtcq
SVSirJT1bOrfZaU34K68/cbhtiL6IGNq2iuqe5VhvtiMY/ykQ46jLy0S15gdT3HKa5NuFnmDEwZX
kAbeXh9AdBfiHs+QIgUgVLDZIczpwkjyPc/jOgR7ZQ3+HOBikrbgtTk0PlOWu47ihFPRKyOPX1Mm
0W4hEu12Za6wFkpwwD0pqZ88kCQ5QZaXZWNeKYoA/gQAINhX5sW1Eju5l9v9LEXEE8/Ey00NDc+d
5daTuAS76bpvuAX3deC/6rJkDGsHSkgPJmfM0x3XKM+bSHS2Jhvq5WbUJys9GXkVjpUVCFg/8fPD
Aefyizfz+WSB9KHtzrTEbLCULDyXFKX9o7J39gkOcvNT/FLXeyz8UZO0LsLacEjWoJ0fNj49sTs/
8+ggg+/YWm26DMhJWiIDBKluCHiry2GFgOMbMPAJlDnmBmZxi2+KZsGQO2j8ONCY/NlSlRrzYOCY
3wOc3FlsIq+fAslQtXrQ1Gc6vdtsB9D2JGAeujLPUQ6NjxsqWPUEx7nU9kmoqU1gI3uxtUb46N9I
gGpN0zvCZoeD2wxq9ncwX6iwLz/bip4a+7gSlUV7CDmoRElUnkB6Wz6q8gycpfSZ++zOR+YguHgC
8xsNZfSnvfxzwN8FQtnjNTHU5cuO30PchbzQ4quJJ8IX9V4nrHP8PARU/3+3SQ0+KmywHyVC/weu
jU65ac5MErWHaKUfq2SLnBUjoiBcCnsTXS/uON72De80jYp4rf0Rh2ENzbTZGbEYybJGHvL1pGkb
GBeojsrBmLrfx6DaTGjKRe6AiMUQJSwt4tYVYVE6YkXVpsWAEiDErjfX947S8x6RoVlCqt/uC5nB
fTdOfj/A6jyXpJr7xTRALHKHdP9WcpEIiidN9KYe9hlURHRjTD9z0bVhEtwYIPpJrbqZwcs7C5GF
DL74Rsmj5MAy34Xc+DIc8JQ+YJwsvoxmNA30xpYNqZWImGxu1SdUkqlPeKKZDe+zoT2yAROHPDLh
7bkbT1SZijY7w3ENwaqX9H7b45mlOC6/BI6zMyEfqHCD/MM4+fLMsxlL9BgcUaCAIhf3eWmmDtN9
aY/m34K7c9M0kDYqW33Hto64jDiRE7RKt/4IZUNO5PQ5Odz5b+NqrR6IvEykySoF2yFeYyF5dwCz
UQEGZOkbDGW6UGUXvXPHCNfv1n2P18caYHuz7lv745fwIGbq5dUzIc12MNKOKshfeuZfuPP3p0x1
eehEnwj2IG/kCeFimu4VjxWEZwTGln2fp85dxWex2XuP3KF9a+X9i/ANjKJ/CEDmldk/eCUEJ4sj
5C6eNro6ulTBiBPywkOc6NDefyq6+wU3yWC87jzQqOhgTj5LdAiDS+8fJMdeJY2PNyiaiZwCY3J1
aQspuqfG6/Dh2OwbJPPpqDeyXOm2/iVvOqpV/P+aZKlQrskr3yONDkQ0ReNWTlXljpb/QwSZ+FJa
ruQt2zIy1YbSRTazidvYWqGkA4l6K/DMxVkTj+h7wKSBM2JrU31sV2ZM5KvwXAD3BRbVUJuf83fl
hHEYC7RaQFrbuJbsSJHljLRKdi2BX4p6SOizeZP1XtBTK9LdeREnImyFPLsSwsp+jRLEsfxsXB70
seY3eqopmtS25tlbM02b5bFsvWl7ipE+bhGjrAk1kWvJLkKwRbiqmQivETttU/rtBhqx7Tzwo7dH
mmthk8K8VmvaI4oo/WBUeJG6zrQRqfogUsIKm56UDOsbXAJWrqFKK/Uy6RKX7fDlVEOM6cnH1YQQ
OnHQbk/MhLm37N8f86cvhocuFomyNSur3rp20eOa70nOUY+wKlHGgjSC5nNhXW7DVsAi7HmRUwP6
4GKa0ggggD4AmVkcGBIYxFXrDpbVe4EAdmEMfw+hpM0mOCWXv6iLBXonzWN9c4fJ6yvDRaxYN3Sy
GSu5m0Ebffkjld3eH2gKZNrP3jpZuyx094GQ5HEYQ5S3m5hfr0X5KdZjUTgAdwjPsrP5+EG0z71D
HcyaLXIvxgfRIFMZwI8ANC/V3uvTRC4sery8PVS62i1p48IVAXUqNhAlPNFMA7UJBSEvAZOZAK+c
y1dL1I5oLySzMQN4KS9vy7PCwTEHGY5Lc2mAD+RSQZFMBcWNTisbbHpf1VtevsuF2SWVHkgAWGqJ
DBuhgQM2PGQgzKVZXgntZbBPrAdFgxl15R8Ls59+HC8qI+ms8jS0XpufIlqFH2j4Dl18r8FFt57S
ihZ5y9cVJyzQ0uSYdzEuD8NkKs2oac2xuIxoVfNo9cPadwp86/soQcfvuTLjifNdTY09gxjRMouS
KmpIgeXYxzrLknCWjuqEtJdUvkELmBWdGHQO+4O41654/QcWrVtBGS3TpBPqVoydNY0snwszsJF1
oNM/zW1lIry6uV7jR+3qWVWdzFr2OZOAf9t0vsGr4R3OXNUMBAT0Gt6+BcXkPmOEIpQ9HOvVRL8K
U0mU3VW5CzbPgTMCZ3ILWOfSCwdm/9mSIvlzI9AbAYyaoSI5imSV/yxfBqvPnacSpp6XtRzfoCTf
DSD1cWb4srmk6tohexKNZO18E2jyCTHWcwfYHVFeQY/5+yT9OTAHOSy56hqfuruWfLC98w7NChXT
cY0tcTBP0P8SO2PdRyJMHz5dN5hT7UYCdXHEjWNlVec8eWFAakFRtHAXyR2iXiTyVFPtI3kbz0xK
WCvccbAW6rU+CB1A4qjoYRIm14KdTNSa6Y3Fxf2TahKgufE0ECtDtv7WSrr0CuH9WzEBtnGT9wRj
3v8XrZnwQqq+UwPPD+sGmkVR/uI+FqYWNMkjWBdPV0JAz4ggV4OYKs4BlHFYi6aK3axuI29UX6xS
96HVu9Ci9lHzbC4a8gE5HMha+X7KNw/z9/vCJs9D58HEl7X42qZ1WmGXoGFu8ZB9BK5T5EzIDttt
GU/gyn3GrLisI39trSNp8fvkFNI3IK95IZ4gJtI+DS2TV/mYb6q2fUYtoXIZ4jHo3cSf68Z4QQpA
U4G3Je8+fOgm8TnAIhulJhr4Jj7o6/Kv0fJ2MlKWIZ5iYcbvRbgzFPWH6cdPlwMIgzfq+XDT/ShR
6fXPASCovRejar0OGoAdHY5U63pJ0a2/RqwpJjRGJhdhNPZ1pXWTfZJ1Xfn3B4H3Hu1QJRJwTByB
l/obhFGWwEl11kNNm4S8706tuWbdTtgZ0hIWNlUVTyugx3Xf87QyrIbCt8G9oY3Bj9Z6kzcIJyAJ
YO+wivu6xRdGsYOqV+edyhKVRP0+jQC0gZmddh7ptQv1SmARx8+4eEcalehCQZclwyOnhC2xbtto
X2icdP0yjpD8nFOANmeeWpTA5LDevt2it0e2pvR2HjQuy0qLe2Ehkskrr8k+IQ9k7ET9p8XrRo9f
nrQNllMr4xcScC7n/2spCySBK49v4J8bqc763mezdbONDLsx5vKruq8UyP/D3sSzph8U7AGJPi44
Pplg/Ve32+PgmLId2JrSIuSEEVx+UeTzMlWDWoVgtte43H691cckyibBA6QhaeI0ztRrhJ4shF8F
hNhC2yqk7F3j2ZPOl3YwoHBnX6sDSBH+tcz5lOj1Yk5WUI615DAX5dHY+mxklkdcQaNeflsZ/9PI
6q6w3FpNanUwy/S3/HqVxVBv5NcqsdR5rawoZzlLAgs4crvepZfW3LrHGRo2q+SAhv4P5tS65E9P
yTrCUUgHLMWZjdz/mwtbPZQJHPe7rP4wQvLRSb8WvRq2rNXDVesm3WzOlhg+yB54aS18OX1dvDCn
SEdNMFuMFE2JfwiGPruiAWmKDBeM3pYuxEZWa4vSLfQl9fYv5Fjp26s/Re+C8bG7F6MJIFds1CXk
kTWdVbyjlagVjCZEgeBp+JrwUiiIt1wvreI+ZF+5s/Kge3SJ4aWTOvaPCow9STLa7e8qSjw1vQLG
j8UvxcjBo3KpYKacSP/T1PN0mytuCew84aFeR8CWTNwBPkcFUHhK12R1op1spDaMowM1o3v8KWPs
yrhDY8KRg17pzHFKORkB9P4phIbTrPznyzFdQ7OoRVGLXeaHJCD/WbeYEY2lLIz3XLLmjs0hMoMz
p1v0ti7z1qnBC7ut05NeSO3W2cQgwKExI3YhhEM7l6gvHImIUo7fEcbXcJpl8fZnuBrgPMyuGQCh
mS1OVaxztDl8FEBj5ctB0Dq5VT+eRY+Ra1m94c8rIXOgbdpc404EwsHfAsvnhHYWalotfRUXLrEh
lcdoeO067adgJsLgjqXNX1xyAFifI+8TNKQ+WgcacQ3tMPhjHNkRCa9N7mOct3H4TocALwLW3v05
hh22v6UDShpv6Rj+Q0zbjTR6MeGqvfwY7KL/hmaCcyIull5LBw9Tl0oNh/Z5a2KUwL3a6O3eVmW/
e51QNY7OYejYYY5SbWKIwevZ3qAOamGTkzW2+FI6df3APtfu9DW0eaKGlRGUC2r6lbhzTMjCmpV6
ZTWRWPMk1rxU9KmkT2OlDGCd5eHK7/YBGySBstU6EVweD8YSX6yB3UCA6vbqjNHLEjLo9KpHw2Q2
VH/w7Ef36Qtx9VE15qkLnC3uBzNWp1UCeNYybzEBmQRo3LKCSPmk3G48tF8AS0lu6TN/kqP92YOU
3thrKMj0uY2vaXzbc8L8M22WPZaq2wD/04fgR8UQAUnhi+hik51HDXv+EDo8fzNp6aWUGxWR/HF1
8lE6hUbp2A03ACqCyXkWCckeePtSfMXDCImpsMR5O4qpqpJZyEdrGhwfY/axQnlD+wZGNUWt6fqZ
OPWGDADUxDZC9dKWAjNMNJVxiLRxh5r9S3XLHTBnpfTezqedYdNZdC2Q5xdioWsWGKbW3UuRKP2b
SKqwrlLzWmic7RGEVE+oAXkEAFIOk5MBhYtfM96nu/GKSbQXh4iePdYVhcvo/wOOE67DXUxj64p7
LUkFN/7j8BLoRVB8/rY4H57rp3kD6+MvXSNSCU3xkpBTKNn/ssbvr0SQ2gLGrWlJ8hB4xe9q8SC2
viFsbfWk4uX52+ioBR9CMy6VupHCHGTWooSNJcdEsgaTxasYQtRylpgv9u01DxPh4tyVNLfLtDKd
VHg0XHBNmwOZ/BQCBWC8NBv1NBIbmYfo1JTnBYw3Fe1BF06DpDEEw7kN5oxUdBNy6x1BrNE5GzWm
/xxxEzFg+o8zIR1zw9Rw6eEKzxjOkeZsnyplEWVsfwD5xyOn3jOwtYj46/IOCeNmmzV5i4MTji2F
hzia2RCxMqdHEvk05a/VDAXOxX5Ks/iZe47d2F195+MYSer0o/VRQUjuh74crBfP1GlK2PdPrGjc
VABNlvxuURE/+bamFaJq7Cd7uRiz9ZHNqsFbTOZPBW03Fq26vllattZZiLMZgvLxt/wNdyNKHKAe
WvjhumOJ3cj6aH4sidDaNHsiLUh6/jIVgrU3w4KWc0IuDgOkFyLFBd6tnUL5xPPMhEAfWwfvd3q4
nw6wjUZ+T5btFNjyj2uhmj1DOFGlRLddlR5ZtQvOIY6YJtFgMEDommDGSDoOvMwvRvUqA0WT6Zr2
j9vFznyt8vWF4seCNZhLQzHdiQUU2mayde6Huvwon0sDMGo9ztjwSB56bSmCQVh1iHfTHIW3nguN
Va3Tx4oiGzPYs4YEJJUYY4NoRXMclNdb5Wi/DUqYOfAWZFTeV/009NI3/1IbfYbFtoqrYeZWliYh
NgI0zGm/Joq0nAniTsR6fXJIhB8MNAmzhFXAu/Gj/zUqBrXZZlFHkTPrWXObHjo7W2HJKt+OBTVY
+02Wa872qIasJEe7vpy5yVScz+Scu6akEuJjVpfd71+XsNG4Na+HwXDD+nBW7feZxNXQ4kycnoNd
2R92IxLM6Yaf8oux6tez3D2v9a4nZzLGEZjEmWqBvWMdzba95eCFm54YF45DQEK/iQCKj5Jj2Is6
N7gC43wZu/zGhL8pQZdL+IVovV28hbHPAWl++bYqHksmVIagLa2kcvOlfLMruvo8TzbrbCu7UO9s
IfNpjGKhTpnx7P2ryQsOsyQBP4g4gUi6RyyKWfyM0dPDMXCI9m3It9nDoSVYJGNkXBn6klec1Rry
tlvBKKC9uvKA2yV7mpzKx1+gK/Pek2xdHJgT4G/TFAevs9atRymF6YHbOT0gne22Z9q85zFykZ5b
JYsPJymUclbET2fqMfcVECmBL8nylRdRqUFKMmiAkwSPBYq0NJWLV/I3emBLjWYp+kr8WiGsJt1Y
+4qxKBUIs+Xzib4WeWs5yGsv9WbgGp90GHiQqsKbtjmSJUgqMYPBaw+KIpxN/KydSA5FvebgA303
V28xBsSOgXeOb0OmYh/3R1Xh5RUmOFUetOiKGkcFu0Y21X9uutJ+D6m6Hlph1+RT9RPo/InqF+sV
NYzVsSPEkkZdEplaxUDEv2G3YaU6b/yMklXapMGKgw1d2378FtRcybrrQtX378rXS4Dd/tIPsp7x
MNcOQYnJvZz+w800AslDPyoyEr512J2841aF1+dw0sd3lyTzAIL6H968NuXMGnTsf3cj+Fkmeh9N
+zJ5R0S8zeUgms++QmG32AZYLyOZ0J94kTYr67sDh3c64X7hwGmJb4+z8R8S9GMjSR7Cd8CggDVR
15zp+w91VMwA40DIwgm1ynhJz3GI8lMlBEpaU7bcl56puz/bOkzYk515VHb3cY5uLePrG6g/tcsm
LPE+tbjiFMeyx0a5d85qz1DhQ0hiAndKkiJZyOyPojanuAYSXq1lLG3XFvpZmHAvw5qCa73fRf6S
0zMp4MZDb3pPBkwApQKpFuh00KB+SVhAuFmYh0SPf4l+mxJzHb9tu4DHuAgQFmPVk3KdsSYIRbGs
CtPRAYdp1fk7KO2ioVMlc6h+NUu3x64q5XT5c/jc4mla4qQxgx92qHMvAZ71y4cdj8Ot2r8US5u9
IpKADb9WSBr/SRDIi4maS41eCltZqqFoHfwh4Ufv7W9mO8LdAt21fbBQrqW3LL7ar2nYAjlHP+5H
95C9yVTJUyH5zCIj7SXQ9RrWHhh9HAPbuEutqkbOhQxBy88I7nev4Oh+Y+L0q4mECuGu/Mirtpeq
pU0wb58/nHE6lcqCgj/N6Lrw90aM7NCNOVhO0+D4Q6QJyuFLKLfU7ykf+VT/NhQWsmx/2s7R8PkK
vRf9y06u7KOWXrADFRQQhQOZLP7DkfzOhdWwr/A3XFzILLwidKoBv8vrNTaZ1kIoP+NaQIH3t4LN
yiqtmOX5K0BRaaoiaXAJJ3izGuSVMQEATGpAsMJjdZI95Vf7bjNof8zHfl0bxAPsCQ3/uPDJMsGM
2TXW9TX1gf4Z2YDv930+GX+4HFe+0rL0jaQYBb1Lcwqd9vv7gmhBGh/f4m1zHiH2KOyz445qQyN8
ImRwSrbi4GUy5jntV9lgPMcX2jlKG5T1CwXXub9TOOMtMA03WcqFX7qkX8MfI9E4AlyyBK67ud1K
JGSKr7rzkIneGFNQlD4j+4jf+6oHB7jMQNZTNB77PJ6vZTkIS4PxTXUszuwZCGFx6bWNuHykce08
sZJ4NgRQ6JiAZXq98YLiu2ECgmTcP4exucIHhJzD8zptrY+P1+85McYCSG4TFg0bIhAw6FX0MYEh
X6VqaGZj/08XweHoxgsRkfx8/Y0+Ue2QIMRdGo9uFn+5pvSmBrIBmy+fZ0vDhZJrahsWngw4/CNp
WM67i0nZoKVlWJBTtbrkyQ/RlTXQ1bNn1enT1H4VGXjCENHjjxVhDC2WBZZWkSuvTIKhmY74lGbp
VptXEU+MKRmiRsxcTLhDx/2TDRCZeJWsEoL2w0dIO4CBWFUhHpCvej8BcprLJ2/62PBYxW5Ug39l
7d05KNtrPoVWk9pkhKDGvlVf7niglDg1ParbbOUrY3ZahFNfH1cGlg7vAcnhzJG2DH8F0wGMxaJe
IvEXAGgQ90LAn8nAukbMGQEdgRVMMDC7v8Nh1GhH9gbr42i6fljYJv4Tvbg/5FUcSTCKAxCW/ATD
J1Xa3M6Rx55OB0iWxaCOWy9GNCgEkaUzvXCkFPOVpDfnrhEmPQ1PpomFxV1iUa5dxIEbmqW8QxME
z3AxO0NY5gWhNgj+7VQQZqhaOYz4YG/1R3tqQjMB15OERHkWnyZVZ/E6S2ldgl2UTzIFvSm3UUkj
QyGAr0xuNcq39efbeZ1IEgbYV9b3KUdG571mduXUww6QsYFx33zOFcnJAomJSSvYwcSa2LAug2Q2
Bkl2UWu3yWVACbW2LKnesn2Lyw3b/u8Sb7loELpqFer0zqrj3zFM/oWM7Brfh35F14jHlvNi2aRK
OKhzSnCR2If/nTn+Gn04COYFeYBWMiHWwlzQQWHOX3Lm2EgCFw/mU1H3BUFPBgKcYVbk393GNxdX
vd04V4o3TACGKg6Kwe0eHQMt4ckt87n1OZejChWZBvDAk446XybTgYIhVlhnzvmcyYDdoNjBOULy
HKuNUfITaMMaKJXjpbXlZ229LwUiZ2jiHcheF3+/LTiVs3lruEGjj3HL7LY0BPW8qWjLR+S31hc5
B1pQ0lSk/y29CXcJtuOpL1btmvy027o9LibMbpL5GmzdvL3l3kNCMw7l7t0QAlfCyNMU3ZVRe0gI
lnhRcqwUgm7yoyW6y+KQHVhoy3E8YfP6Eajstdt5IYbDBZ3BQK/u0iwVrA6FkTQv2s4M5eKjpe+5
f22hAKnFH8uwb+gKSt320TX+HgiJwxtO2k3mJ17eJZm2Sj4UwbTb7O2AvqYawULgT0OkUH9eDf24
8v7qJDZoY6gx3W8WvabpvNCD2ZT6mDPWVxZjeniMdjYwPR6O/2SXfzvizvLd0Ww4kRhoNbS+IE8Y
1GPYVNdtyTIzF/hKZRPI+1vK3vwYs0KRERmcU5M23nJFBioTLXTO4je5tdFJqNDzQ+7du+YsrmSG
uBOhvSQ8qIQaDMCYIIqICPdBwfJ8a4Gpje4JpRQbNxwhjtFhwtI0B1W1FDCfyp4iyYyeFy3xq9EG
gcqiOSv/m9wjAifabZEHZZoBuNXX9X9ClBcFhD3wK6nrOZX+vqEAFYSn30OtAQ2TrdmHh/3UgjJS
yVG6glMSYJ00KfjAYNwU7AaHbpJxCDboo48ixXaN0D8rYTA3W6nCfOWjpuI7KhdaHQL5hCtoCBT5
vGTMlGoEZoMOXgYWr5vp2ptXzSy2xKBp52yR9ypg5VS6wDYvy7jtopMGUsx7wUUXsgTdB2Ldk8Hj
a/ozR4MUJLmfatyyKmfg0zIwdB8ZFlqEHXBkkrEQ8DU/FtnQ7nJx5xBe81oOIlQmvMKeunjAtqRK
ERrEywjmMb3KgDerjW4OHNzMz3wFF6Mbxdt0NLc/8BuNxao6GJZWjRmUkMOYSp9DDarWhKmrIaez
x9cAYrzv71/xg9Vh41a5r3VrAyXoGakjhZBmc1m2wezsx4nGZO7/Hqc9iCfIxJ1kb6aJja+ZwnKF
AYFf4tBlCW1GSQa/5RePtr3/MkH2kOAK097dhpSwrYIAK6//UqmGwll5FzWugK80Q+5iCv42VgJh
x2nkos1NrSnT8xQCAgLOtCkZlk2Qe+zRVG5gMwAQZIsRN296CjXDUcGRrcALlMlWeQnettdGdTCp
gh5dpnkEjOaB6pfX4l0qj70idtNuGVGTqW0hbHqLNJTIUWCYW4SW2gF9AbGHhbdoEtipIUHewx5E
7LGcNvK9pI5fzD8COE0Tawh5SApOgUsgUdrQKorD73cXmeSYRZcHZ3W1FIU2nX+bmtX2rm+vzg3I
eCzeGP7+ZR5HqdqbyIe20M7jxgeyVFdFAqT8VSktJ6oj/52h56saMvc4t+hDzYNODAOtp0Mp0eK+
4KLIvfyu51YLkwoIq6cdFOo+m0TiTVswxXXrGCtaiUrn07466g7jJv0NT7CKk4D7fsk3IHbL0Cpn
xWfa6drkh1GdBaVgrlRBj9cAlEt/HVQeswQEmtVBcJzLhLiRBKHKBCnEhokihTcu8VBYFgWMcjaX
Kl0LMGfVcsOknzMMKi1hoNI7UIVU9qaajF5I21tBXvpvcLyOeK9hITFE19R6aTbM/AEYqNe1iipv
Wa1q3/m9znMKRSKn1+xzGrlybJJMkFOfCpstv6/WeXuLvmuGpZFQ+utgXadxviFj/fESeCQ93nmG
FBsqSWH7QTdrN5+hqbMk0grRDjTAsb/h9ubaJkt1l8BPvpeOAQu/rNkyN4T7ZkOc/Lk5ULxKNe5I
1RdYRMN3Ly2JWMls17F2Knj1eJmthLHMKjhno1bOU2YSulPsxLUDAXcf+6ucsIqGujO3YlAby9/7
btqzZ/Xyg567i0TcOkprwj6MaIfT7sCITeCU6LwTuV2dUI+zRtViqBYbYz6nuhcEozLAsEG/CaK0
rGhNoWQrYs50xUc7vLHecTUW0K4u8rtNY91DIzi/d0wz37OEeM5WJ86rgTRk1dvuy/IqOaXA1OwL
cnqko7SyoL8ScQb1XZ0X25ZVL1Eg3yVCaWTxBjs/1VjRd91n61Ik5iFAljClMXkKkYYsRf+nuIw1
O4PNsrGlp5hLsK74sTwtQqlbErpS9jBR8eqM3TchrEdfOBJuosZQSfUj8wa6InYp9ufMk9uWEyhk
gGB67W5L0vMtspufvIDAJY52euM0ewa3+y4kudrjYflp2UwdmtlO05fcmAjMUOqH2Zc5za99mmXZ
pT6B8Rd+OBPPy1RIIvxuIwnDq7/VcZ5ApA6Mx6mPdTn/lYztnpOM3Ab3+N+mWwCsdURu5i+TLFAt
oeHVMIQKZ4NmQvuK9746r4z8dncP1+ZkydJVPk+a0zyrrKQOVtkeTjseQGiiZNq3YviM16AA7ZYa
EdkoniRb8FvuRRcsLvBXKsY7PkxPauGDugpnVRBgSHnEFdfmuy65wEbwob3cSYnbP/jjTSKEk6iE
YuVW0CtAaxjvA1+Is1/Z2dmoMMXM1sgYisX6dVHWi85CLrC19HyGdTxZ7yWy7ebqcyOJ7z4NcePi
/sFMoo/CG5xhA9Lct8mKW+pN3gMeyKpbGv5Qdpt/OmVly8B9vqxJlOMgxvNEZyncOmqJ4bE7s6Yw
zt6InocMMxhTYksXAW2ix5feb2dg/ChoqLl8uc66PIjqpHojMcCzIeiQB/YcUButyWAT94yhLvdL
J8BtTzljeJIMjuyUpYcQ+fiavLpFXA7/ta6/dJ166Ap71zNTbGUIgKeGl9rbEGjuYLDCdAmVS4Dh
dOQGLMyrzeZaaqsfFykJZmdBbnG4GNIaW0jhmRnYzurUur7eA44Xlt+wCtrHdm7G2Yvbol/fcIAU
BrAfvAuov2FXxxlIN9ZJ5eDf8l6mIFPF0mVpdYVJOHRm+V+7SK+URzCeGsLcW4AevUv7qe1nE5iJ
vfxDr0rK8c/b7ezGgDLu+EEKHl2m3Vanm3HuIjUdpEl/ogh2j5W9/g+W0FuhKf7GA9OR+BL6ngri
wB7kpakzTaiSi/0sd5JeuPnn6hlAJ6KRquL90e+6/kZ+ngRfFdq5QmIB/Kzl0Q2EMj2a6jtdX6el
CH3QxVoN0fdPHoF+ofSg8yyGXUBLM4yVD2vJQoXT0tlgoJKQH1PFNRkR0XVvqdSdUFFyusQH9Unr
vOxKsdOleV05ds9Ix4DqG2+lq6v6OtahM+e/4QprQw/x8C2sx3tP3PSZnxOpYUBA776mEZhotDot
LIgpUJFZnx3yzhvwTUUTLRv45pV4a86mo4yS6JzIdsZ5GaJNE8vmI5ARb6ySdJehubu3zIw2PfsY
nWyYXJqQ+72AYXoi8tymPNPNHjJOpUS7uZJyrWh0OlWkF9tXjT8rHkR/DL7dLXP9JyzwWDmBQPtx
NSpfDjr/cpugwylISN/Gq4Fl9lK73ueVN1HXLqn4Nd2ZETmwMJ9IYsaEuJ+IpUUzS2lZEDsSSned
Qrt/Emx25tA1t5DfI1LIgqXxclqfoW+ES4PrjTBPnkHPk/nL++i/JLaCb+mjVyDN9K4DOgjaNkLN
G7hBjG8eVeGv2amCTF3GeAAX3gaK7nwF13jfUHISGsJ+EdpXVDZqEaH+vuOO6EUu3VrpsSVRc7mr
GzVO5Wpksd7O+vSmNXlAsH9JwPAd3tYe690MwuLlxDQaYe2krmUVyILjriW+xFqLAZoLEHqTFI8n
zC2K31KPMY1Ry1GhjHwPyUAcof0zQ4nKNQCX/OVOh0lWqdk+UXJ3OyNGvrug+SzHl0C7XmxRPzeY
wDCToMLNLzymhZgrEFwUW64mEyjLuIatUvPt5qsOzJ2ie0AbBYdRTtEBvh54ow9P1hfZgKNEWDNy
uk07loy3OXjXWp3WFoNuZJH4cwORmU4m8BUfUdWMmIzCxjyuGL3tFWeQfzVJ649FstIH9/1/Zqaw
fFiWqvRGkAgp7j3sSAGGiOhYPDaYJ+K7lzw8ez7BclCA/6KzBZtbk01I/Hmy5ARLKgvR6Z5XwHHO
xhL326zDmX+ae8p/YaRfu2KHVC5cnHZ1niMH/xs/WXZ7eISmFjBjx0m6EHWvVP76MH+Gym2LTs02
SNUbkuZIdoO/Yp6Pw176tZ4PIa1TmpQdb+a8IyOBhLjZ9ddteOKBKtu/EiTZZ+5mxicF+r2S1c6e
MkRKC/pJGGOVWITa1rSJ5Hvnx5o68KK1tsS+zhe8fVMYwn0SVqM0mR3HUGGf8s73UwTyWSF70qSs
glgwmXzn1Q5dJzyCAEY7vHBGumwipw/F+rVvCE+OUpaZJtL95Y8iik9oF8q7outhroaVlPCbajxN
fk0TwWkpfM+sOz4RSvTvu81RQWBpFqN94noy9jlk2ABuzK3Rn+ViVauvEbCG4InpQaJ/z8/8DCeU
Qrh3oUQ5v2oFOOYY+YBMmvJKY0IRyRnD5wrd/d7rDbW8BDcuOKJM0XUymKjfZ91vO4rrY7u8P1Il
S6csTjyfq0eoo0Va4N91kiJfFc2cgiyAySv4iT8pUHJVLuPUM/j31oKuAa67LmaF+W36n0c+d1l8
I/vrhmAHRhITj/2tPcV9D9VhdXDL6qiOI2DKJouTxNYphzYXAk2OYQL0ar7oJW6EU1oAfu+HxM0v
kzFHGdVfXX9U1aUM6g0dKRC+fhgXDL3PDakXb+FpRrw34kPGT3RvtPBChm0+34F8sxN/z/oMEw7o
NUKmrf23G642O0xeGQvQSrQpSomSYq1YFdzNQQT8gDXfEj8ySRb0/2DLWqo3mMwwPtPLiB0XcMlK
FGbyDB+t31Y1t5wEcruVJy9PF6az/bVzt/284TXXx+A2+bzpthV8bG+TVbizSS8UOoARUyjEEAv4
yVaPo/mBIyWXQbJUXq8PE3br1l8YTW+1Pptbtq52QvQ2Q+7AbUoSaTgdCgEm5Q+2TicQMY/Su0pb
758fmPC3fR57VFnkB2JgDhE9bp4Gx+EVJVmttn2iLnezZQvSQXFgP2AbnUEoSvdmudeEcFN8eWF6
iQlvn5/cUCX/wrmoRwN3Mj01+dM5wnUhvipZ2VOa2JcXgM6fWHVmd9P1IANgCqW4nSYuO+jPA4/A
HYu1peE+Rxvhx1MagDsSbNd2j6QsJ8ExLAVQPxZ3/wyHuwRqcj/JYkLq+i3mjJeBHnN8BdkcIV40
Eq0xcU2vuArPKkiTEfun/0U2nJ3mmYtW/rGg0bBWnBDKjC0U3tjCK62KmD8VvgUa4aJwYmxw7igc
V+BNNu93tZC9hJ7kM8kHW8cARjxcWr3LfR3BkmmrIedt5QoXUYjBa/mxxjgZnHCvqfhU3FgXS7n0
MORqUcoOHptn/QUDAVEu+/bao4SqqqcYazZ3owWQaIO0705zTxZbFs81ys7kPwp1fjJ5CmNc1Mub
EFsPOCjGOdlAWSw4XtqZ1HgJ4JI+JC72p48Zd3SMYYub0vWCAtMhSKtlDv6Q4fbf/KJlhgOyRRLk
Y5nvTr6a1hWlmC88eEWvFj/FhrD5ixVN0a2368pMFCGRx4F9gfEsYjEpkSerH4+PkDNAQw1BWdsR
l4Ifu9nE0QF2VvKXfo4ePRnpPgngXA+NDvTfVEYs0rTsC2TzCWeN5Zg+JMhLKWchyBou6eQE9jXZ
QyMM5C+IkVcI5xLhDfbX9A8VZeyRi8PYZovvJaNksnTZXrjEMEea7SD5u0gLCjgQNvL44ICcvQdf
n6xSHr4iALcew5DXKJIdnSgFHwsJM06y1KPGeLzr+KDv4L93TpK2wcbZ9EtGBek33jOvofQOmiQI
kDXqR59W5N7alZFZ89Yt1z4t0LQvKZlyy60lj9J8x7FLJ4nPheKWPgl9lCoRE8PzqHjeVC1m9Hhy
hKJVBB4kOQasM/OkW4ruEP/t7Ej1m9TqUqZKIqba1X7p1YearIrxnXk6FfnP6G8F2g/AwNYCCu4R
Eq8RgX9jE1izw4lOClSuz1qIuf/WSJPnSHVM/j+tp/kTBNnPqxd5DZXquxjW0tK7KDT7cxuHYXRd
rdYH/j5aanBqrk+XVxsBYPc+2d/uea1nIbkT62d/oZ0ZFw3O7EKsx1M1Jjfsn36+g34dkYgEaKhm
aRTMgimZ7Valiq4aX6YGsSD1HBOkaHzHSOhl+FnmZruccKgN7YF7+3fIdgyrfeyagFb0tvHW0Y3+
QsK1A11uHLJC9iZUZtPe2NRthz8bJE3TIA1Nt3FVypM0B3NiZgkKBbqn4wXjhFz9mbkEvBEWSDZW
klceib+rRjDbFUT7aY0LxuGjJMmmgYKmJ1c9wto4aJwIyfeogRxD1NMgLO8oiC+o4xDU3I0wax1K
7iqTOdeh90moid5rVrDfZe/BRgZKuoiVwqLP44wCoA2YqrFCSQThCXfLxc3isjLh8YBpW0KmsnM6
K9H5gpluMf7IanFmDiRTC282mhbK5UaeLmlsrx+h0PJtJ6DsWHPqPW2+YUxg6JDCZ63HWk1YwDxX
ff0ENhxJ8295NkfiqB5hC+SxLzvScgIdy5BOPSn1EGaSoSL93R+rgukKH2HF1JetApJJhlfu1JzX
ksqW7EK2Tt4LF3gaHRFHslh6BiDJCMpItW9rMqt8e8QG5+TFFdFiF3PAuWxQyBiUZNFOdbERq3wC
4ki9JTZ3jXEkAcchaTroYetnvBjT2t5DUn8LDuw6rS5xmnujvIHEzGA9c3JxcvJGzoNk4XGCSTlj
SHS17T8zBStmxnbJoJO3EnckP4iCqdMMXMFHtpsNMk9x5qkaEBA/My+5A0ROKWs7reXKPqCUHcXi
s0S7F8vef95GWZ77vRl0M5KRTRngwilMV9H2YmnOc8vicem4tHbWO2auyaA/4zeP66+ZoDIpyydd
HbUs3CPj2VKSzZ3Kz8Fg0VhqNat5Cu7tmzDtsjvd2dp0xa5A1ACmENyajctSOnKhTpW7vFEhaDin
v6zsMxTzyYF3DZK088YLYPt4CF+LnyNYQ8CQCjLo4rFIGVf/xXa7aDCKAmU7zJ0H3hEIhTJKMfs6
bcdjdLWzhQuuIk/PxOrizIrV7p0akuGBp1+79iDqTUo1Mq9/+9PCDOEzX5KiJA6XgWxpX+C1nb6c
GXvyzuv2MguPVOtgoWGjP+IVyXHQiNpsWfNGR3ekZCz6WJMbxLDAmmTHTvMH3IpqZoUIw+ylqvGI
9CfsNzz5HdyQx3IDHQTPxiBG0QnzGnvR3R/T1sOeVk55TCFKgLREJGhYrNWurcDgiIA88H1tvwiE
4WISIomEZmmBxyXhqyUNYkDMhDc/5O6gZI9XCq4M9V6hclYcDBpVAG2MEaAUd77bRT9lAUkYDYya
HyeQzyZ185PdbqvtD7dD7inUS3zsVZ8JYy0OahSjl2FVOP8esBZcY86zL0/QU4Ir84p14JI1EN3E
Oe7j7ETtEoWS2SxeF2OGNFnE/Sdg8FfUMBrKheVAS1odSlsvxatztEDG3hfFmlfunVtBXtf2yX2b
AgqqYlIGFSahZfr/tUn6NA6Wg1ZFiDeE1ymmvOlwEWUFaXeiWLENSpqOvq0BmTfZ8jsmMLk5u8z5
ATHwF0E6gm180CHnBHf4NW5e5RGDI29iwlVDjivMJ4jVXWZATfdfnRh14qHl+2HgnwP3Fgh+Unp7
sxrC0TJHdyGlsO1DKK/gJg6xyNoIkxtv763/bi2GbQ8YXrbd6aYssSiHwInPs8ysoglFifikl8tc
tSWqvGAe04nRG+xyxAuEPflprlZWknzKIFTw7rpAoS3YA2XpKSHKZa1PdlU9OurVKS58mmzemrsa
dLkPvL39ITrJZh+PS4bKPhE2MDpddJyPkPEQWO1UA9tWpEFo1ReuyLKofrsyHBPOoruswM6qbvdD
2fgNr8TnJNHCfrCJJ05g3z/2NeKWA8usqPnz9TF7ncSPrNCdE/zvgcX2mHgHyuXV9OqP9fQqP5+k
N44psnOkvyTVSPbNhtv4jr658p2CIoKgVymvCKmCZkta+WEbarYOryYCRLe08ULscynN6OkqYLzq
5AsYnrd7pH9R9WEmyG/EAsF2bfgUDE3WBvXK7k28tVimmcsxgGFFVhwZiX7HqCcRvZWhLFPc0rHt
bTdCUDcoG9F8pHv9SHKCMCd5xG8gyyTYY1MMbN7zI8R3tf+L1u2rmabj/g7vq2xh5gF16Au3vF5K
KB1i4yT3aLNujeUiqR9qkiP4PMmBqv+P5ED1qrLEog+FwpWMFb1l+BxNSIbUHCWvKRINzRquSpbY
uMYm6/S04+NwoEg52QvNZ/PF/em2RS+u5xch/01gmn6FcbcP1cLMF7aKTZgtLTELiv43RCOl6TsF
hBDVAujkk2IVbqOjocLJfjPOdRC/9S8dglGfi6Fn2rrecIsxQxEmht1T8d9NzQX9UH/L89y7gSz8
8j+iPfC5+Cy/kB5Dhn5WAmZVLnP76/6+7KV8K8A7W9rHLbpCbZS/LhO3i5xfk4notqfMoe8QS+ec
Ib8yitr81M2qd0dL1cBPhcjD1679mKUFxwtxRtkianc9j8UCU0bXjyrkLkYovByrcJJZJ2bScDty
VPkCSqSsaUXISzlUE2HF/Kx2adwYYuWNw2wp95CmSGi4jtK6ddOpHTgprvUmsQUKXyoZKbNbJHV0
ZWNEZaPRmKn0aH++hEv0Jr+80D+SDiPqcECU0Z95kffNmrjsWUOhLXf7aPnlX1Avrs+rVqW24WQk
QJ+9warg/3NB4X+uZ4cPWx5fgv0XXWGXLg0fec0K7u25dd6erCv65LXHeVyuzFlENODIDzSbAkzE
5tM9UneS3Hytpbxw7B6nteu5sMldfl9T5wxs9WAMsb0mUOnoaQEY9+ENbnQtNXN71PGe7HTEknfW
wB+Lr2TnrJw60bPET5TrOxToTWNZzLy+ttHv7lqy4jEv1LHGFnXm0uRGGwl7gghCmWNGwVkWCguA
+09Y8c/XtsRXP8wJjCTpKumfQnNACB3bqBmTidxVQJKOGfvdm/8WOSVlTKxTcVNDjNr+C4rpn8G6
FJCPNywJgp9ze0Y1V4Y6tnd2ZqskCb63BapJlW9io2AQIJniTuVcnm2s8SUrgmk40FJtgUg9/6VX
O61CwTZ6O580pHTRJXMG9XOaLeJK1w33hfZTdf+x5eKoeaq6sKamDVGhIhtARikN8FJeMIRrrSgD
gUhx5CSo5ISnpSZTsOCsZ9NhBM5BX1fCDUqldImwVMnOkJ/4Gn1mWZQu7SJYQQe1ItugUCVn0VTv
wHxk5RzqGiir8D3wYXrv9jvx03pThrcRHi1ctgWXPqjHX77eS/LMhjAhaMeNmlmvdB8pzdf+O11b
yUh6+ypDk4CxJe9mW23QZbY1B+GBdnYOH8ULrs5xsSJb5y0kgZRGTSInIoEFkpaamshHhojqaUbV
nyLA3yqmiL6vKPwp06E3Ts862R/+LbrF1mjh60COmAB3nXCV7t+y2HpMhaQcmIwAYL74CuTm4+rz
0x02Ab7DcCr/J/vEkr8qRsQxjSkNTAGKuhkeXBdkkGo7nlxePOfrOgMVAQepO09s21a0zc61rfj3
OQXcpsY/j7tcABuXUxawo7UdpD1Z2i5LQgRdWnQ9UY/6FcTyTeeUX3bxYjCw2UyYxx7WAmtbj+fx
3z1hVILgPkwIczHFlrS4WU8C63ASA5Vq0j23tPj5jkeN4St8SPunnRVgspDFiYBruZSUtGwdw5Ku
phQH3XWqCMyO19qhA6Kj2Ak7oESNQYdTZkgpIh3tbZFTTOj2hmiDq/f+yVlJJx5c7doYTLWwX30J
kEKjE0xafg9fj+3eE77VlK9w+KTQHDPAJcnKIulf9mJiT5zuu12wPGRPNE9gAckHTMoNTH+OSKPT
TZWcceVvuXvOJT1i4ffjqILuBkhFDuTRwnbmyFihG8PtF3lZPAzZkCt975wQ3bnYaOy+C1YH2LW6
sBeMWXEzzwmgSGE6cJpBoh+L/oKlZkXho4ZK5iHTokM74akCm2Gi/v7xboG29BcFO0Gk70LmZtKw
Quu9ab9ad/61YzqAy3Bjg9QCpJ6YHlKNVWU2kzGk22M0Tzwcb7l4Ug2g4w0cQ2iUd9vEiOu3k5bo
bRIcDLYRdlJM0/LQ6Acsau8yq33BKmNU6u10sV63H0lficclUt0HB3/tXfum3+xvpnNGnIFiJQXh
hQv2pnwAPXhQVYs+2Zi4g3kO0PA+b+0lwUPFjBSIo7fF8vyV1BA8eoS3h6uFf63avkz5haoE7Ag1
iN/gERYtNT5yeWM2OB4Hk9paIYgqGeR12f2X2vY0UvG7PTh6b01eiYSeoMbjzG92z+LWL3rCtfJ0
UifoH0yDxgi0QheMujXQEbly38O9I7/s50YoxIucrKwXMU0aR9be/kgsf1lBWHAUERbzG5al5PKA
6a6L66l11Ih6E0FqjkwJ8fbAxVbM0Hu/eNKqhAuELBRDfBVUm0BE3UFwUpykaR2ktAIfTD42nB9X
5wJVEwqLmHX/pEc5D8QYw450nH1cOc6HAhRxDOX5yFzydKuwQX7KZb0EwD6WZFDNotnR+i3F9aSp
yprVpy/FeasJe5wb7DEdHl17OgVaJTIlfe0D6jTdO1P3hzz3dcvu1C8t8rTq9uWP5J9Uit0lq3l6
dPClc7iKJSMhVnEbR91+B+uLYD9jUawOgGm+4Nr9VhobxuThhF+2JY18Yx3JQ7qt0Vj4EdBT55bn
8mZWu4w3/Ual8SEK7hG3G9TM51/PzV4i7tNCKi6uNEDvlcdZDGQEGd4J2hVNAM+andRP5bp3Qq00
AmicytfViuLJfL95OBR2t/f5RjTxdCIeBOcddjF6eCiLBdRorPDxTy0dvqmQipqsD6Or7n0sTlSN
JpRU7cfSUTqhM4erHMwyx033dJDrJ4ycnZrwKR1dHYeyGRUIVmYnVEH0CsZ/AOr+9wZyDEXkWEMp
uelSSuc15nOtsqnkbznX95YXKeqmNZo9zYzPHOrCfGJSNEah7zqBJM1+cY4h/dBGzgSXSDpL5Nj/
7SDTxinfZo87i0xX5ecMtKBwzAJ3j8yEokNDLvdccyaXQ01SA7pSuCAd653xZPIRFfoB0LF5Sf8o
laoIgSFakP1GRIYJ5ZJ8rKAAFDWfF5r5F4bxUueirga0Wzokk4O6wXeZu6sfttbak32WyEP6XZPE
Ti+6f4Ngd9CxOigB1+xDFI9rHbzVJpJXfcf3gbhmfUd5BfLuGqBQNIlJAK+zhQ1bjfqjPlhxh5sJ
nSq+Jc0ak/elznRb8RBWTxwUyy9Aeq+H7awRt5yIgjoqhGnCkyfmz4zDn1k8m+cAeLlavrJIC7EG
gLRhkIzY3Jiwk9T3mU4Xj8WfqHHw7M1BkfVIQ7DqKy2py93qHdlK7SeinMRSezjhWD9X4PRuQ48N
NOAuy5zSUNlrNuh+OxyCFxJ3iCdO5dyXJIwAzaywfV653uPG2amD35ZyVJUM1PL4FBeqVoX8Kq1O
ndxQFZRTtsD6Fc4HEjtxutP+7JdcANjQhlPfKlJVqQm33qzJBmd+/yURySm6yMajP/fj/BqLrn/z
hgdD3KtSXpUd99oYXfUX4/5QALsydqKq4EqdonRqQndCTMz/oFRUYutlAvYcH8nYYw3y52dpVJGY
bBHvBTdT5d6qQ7iJhZlVlz8J6sYewrcOiMtXg/zC8bgcHhyQjItdbYD2OjhIkV6ZQkn+ItTJfaW9
Vc/QDINXqv2qqdre+JKQ/NZGZRe33+yFEzUmSgplv6eBC3JPMVfPhM+GGL6D42W4x6usOD3fTvXX
vJEqw5KfAoIT9WjZ3D2Xteu1Qg+uJ5BGCDYres+yKRFqiy75H2iPB+7zSV9DBll4MKedqUCMlJ1W
JOHMONsFt+u9c9KDgey+l0g/9yZeacMfTh4hq7FadehgA6h+SoVguiw1/ODAmxLodOvJHNIdIKyL
BtPnKS0IfRaTqU0GYspjKKuLLjDbPLdnLf1z710CU7g6v65hqozh95ioFzyQRtkdDdgrnv503q64
UloMAh4s+I9Qm81nu28r+taHJAjAwnA6izMDTohXdW+Q1efVa4kpZQ4mt/vMOvstfgar2+3w+r+B
ypHd6A8uZUuE/mhZevadtlL4lQQWqygKYQsNz5vHPToOlY//99THk7KnPzin8RwSZSvaZutC0kFa
+ds6A/pBu+Xof3B4zyTohCgGTKlsFqz68dei3YP+CsjCFXOr+jJvIwslcyjbfha/yHMkF++3W7Pd
I96JWxwYbVgnofQ0O/l3sEqUxRumjRrkN+6kNNzvkDgv9jWH74Num9F/AE7e0BAaxlBDAJleGIrQ
ziLD6EbzolSuvSb1eNNn8+LVlTtehktv1hJEKpEMncrphRdEDpzxbTtJL7ODwQZ9UwwCGCZJFPhc
DUU3LNdtj0WntinS5A71aFnDUd7xXlbWUGv7GKrFMWBhtU4mh0ET0DysYmQTD2FS6lAMDrfllF3T
kRkcocDpA/4h+EdjP1FVR3CHkTfyiHP6F88wa5DYNX0kU7+pfxc8W3uCHM/qHU8UmfKT68L6i/wu
qOy5jwhDYsPS9p9HYwVPUkk2bueO8RGu75hL9g3X2+fe5YT4FkuWH8oGiHW0/D/zM9VMYgSGkErz
zV+8tJ2MlI8V4NhjDptbI/WuPKL554lIf11gnTE/t++lAlYuXZH8Qf4BN9uf6v1LmWIBRwBTlLrc
NuLKvhDbmdEUDhhzVFO3Gr3V+L+ErEyGXyS9qkNVe5xaqk9HRC4wYTALrO4ar24rFm/uxYMDJ9H8
6nP6IzdVenXV1HjvEoEAwhXkeFzs1bxH0V/b0maR/FYdw7TRB8BLHcvl5GVPGTVeaR6BY0BvaeDO
zTWftdIehG0cwTjuf4JNBnGPMv0L/lvVuvQhZSsJADudqDQI6Q4ya+2u48r3trarookG0ElRjUxt
net45vfhaT2OxmZzzua9D2vcc0qd/ljRddEVNyEw8rcSZLUSxDy5opOfuId2QtubQJvM9Rpt1Lj3
0cSzpXVOWu3oDKhym9rQhl9P6odMbhqVwUAiwLr1iYukHAgpImMv9pw60ebOD8urRaEqyHdScvh3
7nmxQM52IT/YwOLm8YAzTS8i26/FkidfRthdu5ncdiEXlZ0tOAUd5lEcehzVbUda9fjQi6/VQA0n
ZCOaaJ2Ll2hsHBIGqJsrJmu0HWjbsZrkq4JIk4B6lG5yAkrqxFGPYyjS+dpkVKAdsgD2x1p5Mv9y
qnPWfRJs2Kk5EjlpY8oZ6H2G/U1jQV5EYG/pcwYjtF0nXnqa4l6fvmPZO9W27PP2q4QJgDv2sjkM
C0gew1JPtxrVYHY0oCW/BezhHXMo8qP1zeYFu/tJ/p8xRB0oEryvNjW/JD656xE07Gz8W35xvlV1
YuQZbyf4E4jcAQucpsxVDMjNkl35b6pJRJz+fhrsuvg/Ug8C1xZ3IQ4ZHvHscxCh7w0sPLXd7GhX
Xhkt6keHWVKR8/1u9kBIosgl6cHUqHuSvPbrE0u/uUelK3bPy9tnlz4l6hCwDJzFKAWKnPgHg0Gt
nwaZaFmgCMJYN9Q3va3QgUn0Sweo6FMk4spLfBeGN/Q1u7Uwj9GaGMJUuyNOpk/3HuC/o83T2Bo0
5kYtPb01kcnvc9Cz93I47bJ7RyvnIY79FUq938G3WbuAU7A9jkitkxj6Sz93arMVBQSTsoIynB8n
0zsqWorpMvORbxmc5Vu6oLFprBm6nH0DlXqnJB/vQnvHjsfyAyifbOKVWeHQItjspH+UMmR0ulsY
+CcpsJaO9eUwNDzf7VPXDmpDL/Td/k2lKNjepB/zHcdMqe/dKLBut8XzfCei+MsbAuSH0h36q4rC
PpWEvgDUohmHlevQAeQTxHw0ZRiJAi2k+2fIMNyP4SzAjgyRY9biyeVvREf8a29jknnsi6yl8bRB
aaNUWYEGqhvNaE9ewEwtPqX+azmooVBVNmwwSM8PkI7+V35ETq25pfFpFO6RGaoJ4A4kCkmDQQ2i
noyiUJUMjAQcpLDmxqLXL6HkRA6YC0T+3bbrGj75oLmTYOUDJ1GjDXnESbViaETxS3wpUqTaJNyJ
1H28r4pa0UEQQVDr3pBS+PtgwKnsR85+9N1HW3U2hWjD4D/Qdnuffh3pDDi1CVx7AlplTexdmkvU
dkJfuXqltNM2wZ+R73ukQpK61Oj4IfDWEebMiJ8ZMlbwxHdoy2nhTcw+YAKfmCdlBT+mx+3iSdin
bx6dv+P1RNA/Tuzun1mtRLb7sKuGoWWCGQaSl3MTDp0G3DMLRC0WEeo2aaJLPMBW4BasK+49YvAU
iCzy2iFt3VP5eARNYVPW5R9sn+nK0Pp4CjMRcA5o53KtX6HkhKTtvLTzUfZKW2B10MJkZ57/lVWh
NYh/HdUclsYJ9yiaAu4Yh45uroSlyO++FlmOhuXSNxghlX4MXY6xleHW9tMEtDRb81k2RUmCaz6d
Ya4495taJKEKzJzf2lm9Cfrc4CVnuD6MzwX0w1Rf+ai/L610FznQtTsZ6QDhlKkoqF1uTh425rbl
tNYy85iLVtbmWP2pzuwN3G78qipZpPQqBtZ+xohTvhLhA6YjsC8uc2+zZq4KC1zZxIfol3hLDbRW
6u9nV+5cJZUNW14R+AsLt6XRdNmBwjYOHjqpsCHux1f6383UcAp1u3kRgAeaPpApz7Gqt1UeW/2S
VeShVhVWGbuf51OfkwA+odQE/zFF1BrhRD4EKjKH/ykzTYbvl17+mdwtYFE0AP4chg07P4xykHax
qvnR8x7CaWcqXncx04+5vZ6rYP1+Olhqa+YXYjhLNHOwjtwRGWgf3KAlYHiJpWnKxfRxvo9oftH3
O5n0fFPltWIOLoQvM8x5zBSoJNw2E332yQa4TN+CZtAPfppf3eLp3Xcua+9xzD9NRwj3M4GdgHgq
sCl5/oOPG5GyQP3w4d6NQG/BAnAVK2tCWEBAyui8OwjGEguDiT+A9TgMKfXRYVFEULZjK6yUEo4V
CULr4VFmRiRr7LQmh2NMYJy4LAk06r7qtGt4/OdwQOqy9ysNb9HHvXWjXumnSWuGowrJAnV9zMVD
tc11GUHYi8Q/S0t0vwOZi8v8yfDTnW2XyascJ/bOXuXf3noCxdpev/kDYviem1/pNV/TQohD+CgF
hDbmBslz3CMq+07E5XBKZl5U5pkgARf6hOacZDWV+X3p4Je8Z911Km8EZJF66BFN+tcAMu8U4uCN
21EYV9D+TbfxRQDXJtzjFG7oVX3aGOgdvTvXOPtqvsyOK/xsAOR91b6I6E+oPBTFY4nM1neXqqIk
MEIVKwwFfo80VeOrI1JCyF7LxRYX65cikDZxoE2tNRLPw6eZZMgra88jTq98Ai5PKPVcV/CRDuUL
SRewaULW9O5IK5pLWB/Gysd0CNl7mH8rrmtiE4pGMRIvlSMrLM1oyuXKUZWXu8Ia/VveA1jlUKj7
QB0cJgwRWEH/fXDLIHI6noeJ3ymRYYjyokcNBWDEWtxY5ct7TlS4Nwzl4gJvnrTatg1sP3oDtAAC
qQZmuCCWtvfoYZRVQRMcdXyAwYBCVIUhrOrJZoL7aDuKh5QrRPNzpPzxwtZHW4IPJtxuUNj9C1rz
0P2sx4A9xoYpdKlXb4w6VyIJsX3+aQhdhk4n9/pwFZsQhqc9cRmp8BEWBwWvd9UCpgUUoqNnr5f1
QvCSS5fgkCw9P3fGTqrXChAoq5I+idPIYw1qEkzlvJEwnH6vSEqlbfgfF+fPTW9TJhX2JXpE4qps
ac3QHw3Emn4QE/eVdPZl6dfT7fRS6IWX6mQ+RjRSTlosN2bE5VBl4Ml38rp6lmJoYQB/7/ScHCWp
i7/QIwykWhcR9mnZvOIH/Ewhy5A2KdbRseAcea+vNrQZeoVsZIGtHNn/kcew8+0WKRDZrhFbPejc
JR75wZS9HtrEzXldXOGPrF4GeLQSqa0PnYokuXjI4uQFYOWI9jvXbvMdIWQAvlEvnsMOPGGPrux3
hXxicygh+/EM7ZaMoadmo5ymOspweMjXJMgAYpbhbbyF2BER/yhUncRWmkUuQWwh3C0E2qGPyV4G
6Ivoo56qAhw+CdAcnFpxkpbR0rJTs2J/7+aQWEZgYH0XSJapLpLkf4/wMO07yDmfEv0n+Q9MexH4
QZF8encY7HvdwIFHpnH2UD47xoEfuvuVYRnu5kgCD0xgMrxetnPLONtiD5TJZ3I8joAgZoGeuCt0
mSDwF55WnEjetdh+mvcI9Htsar7n59YOrTDI713hCGrDUVbOvgbPj6MCCMnXgchKsec0gRF5wyDh
VsMAb0sEo4SH1LD1BQOdDuE+l5s3JXs8CVLTxznar0HJiSgIuZw9UHVL1ax5nXRVj7yf5I84kadQ
zItDqXKSVUtsrigk5IBYjQJjR/J3v+5nS+5UPtFk7RKonXi5JhAcm3VUP95OJlfE3H0IK+g8RNeQ
hXWq4MbbCsyNTS5j1u/j/6NEQI8U/20vLVdrM4NMZE2zHAo1lzH6kQ0mV7OxQ/S0QJzzLH/RTll/
a5czVt/xT4W8xgs7vACg49wQpocKnz8aLwgih4Ai4n0Dlrojxd9/Ifeg258qga/nl2F6i8swdibd
q8zLNKZx3KltbwX4l6hFOWV42T0JfA94zXIJU2NFv7A3h+TE+quMYEN+3E+63qCDoZTdDZ/Hc5tQ
QW9PmPbxKq+7rs3YV0yrMqcEKt1kH6azGRs0ipZOvE/ElYcltP4McdRDX/kL+6JkXHC2P4clCo5c
wnuSMmdGb9zuFWDB5LgwfcyGHN2kRxP1K2IdhVHhXM0zdXCYjjbOtjTFA4Uh066CZ6tT7hbYXblW
R9hZDD9O1ebUyl7Ht36u73k33tdBj3RCdKC8JKTCqmqCOZKJZNE+8HV0EY1WNxHPJ9WJE5udT/Xk
aZx6sdIAELjPLVGZUpEfIrQs1CVN32qk64ifYvDFP41ex+7rMfiAWq9CRQy/qUDdxl7I5avr6TEU
z2MM2aEagfvXrc/GzU/HkebwNfDBXgsXcin5q9qsR8RV+KrUwSKmEyVF/un4ehtqVnx3lfrh0BtI
QjRGoIH7LSKZKb3uewDo9Y2lpX92YhMyyFPSKZR+AEqjsSP2/XFaf9S3/aQfVoPS+rFI242Uhlot
Nrls/Ux5+iBve4LELZJ28/EJ5Dzkj422HKp+VLrCXW3V7qY8MxeYiBlSY+vlV/g2gzClBTaI+YwZ
YNwQ5Yc1Ef0j6g7Tpo2QhwqKBQgzqmiewuz46TzWJD6jpYFrV5v2xltjYAaVL5UJ767zMgmPfL8r
l9FYHWktdIWaHlf84fx8tAsxE4zv3hqL6MnsVYVcVk+m249G3253s0g49UFhYhkXwn8N5zq2+z5C
yE0vPQVTMMmGXJjkLPppPyqnt34W6XrawJLtRRk1RTqgnw590UK71GY5vLziiWGZ5Jo/tfNjdAC6
t7R7bYuKL1zRJRG9ifmVZSBY6qQas1Gpphq7NbFP9l3aWCOEgDYAhCNwzNJWpTW9XYqq4jqGL7nk
Y8KWBzC/0m9l1Nj/af1QHNV9Ayi9gU9N/vBI1r6rORxDTrlL4UFQ5VeGOAMfTjQPVgaXekYV87Cf
12hk+xk6QdjJocWIgjy/ANZPx92cg3QW/yYRCBUQqfke3ukTcpD357ez55XD8S39kUfwjy1zBQtp
J+d7sTGVIKzkUulgf6THF4h6H4nMgrcEq+8jTaC7sDJz6DFgAogD3fxzYOP1p65g2lWN36BM0Oo0
z3QronFCrJn2ZesrtMPRTlfc+pfWe0qLAXMtryeVSpIkqfzqsRD00JFZ/n4eZr5pogd+VVBjB+l8
sIepKNC5TQH+qF9v7F8UfAnkAlYL4cfkGaIqRnc2rlTNp6u+/mxxg+QYKa8G+Mt9bJOfe6z7cXGZ
xXWdkiPsJ0cl8SOh1I4RV8qXZKRfydXXfZKUYNs1QBcveJuN4cr2KPGZsTMgdiSD66w2KqWQoZue
1rxjJBTKtA49RCJn+7HDnwn0okFONLHsqxYIwe61kq0l2FZotdbxWV2zyse+o8+kYrvyHi5C7Ebg
L8OXyaBUp1YawXXN4OmfaztRJFokkTunIxxXXim9mp9jd5MeQYcgmwgR2Pyk67St/hpTdwic5TMA
lWFBDztI2B9EVJwPxY6b5V1idvGS+6A54TqSwOHnbkWsJcIyhQgPXYC8RP796OP1KHKbmxkMa8Ln
frZUC7slpJ/VOWYXgkoZ3pQljAewqCt2+catWCw2bnaNHbbmjl+rCF4sayqVAfUWyzrHxyfHkLsI
Ohixwik+fzPFoKWD0WMh5lp+DMfAEfMuGNX3AOXiB3r4WYgjhNyZ7uIakRARLWIXGWmQcM3kscBF
mUsiHaSYgLvbyPL2TxOnWC481u2l39VQSC1HVIezuOUA48P7dSDnS+LYtiSTCs3Zrr9zqm2zPhbQ
jdUp8ankXTws+BklztaVqhuk6z06E10nggQkIR3z/oOSr5NtEa3Nt+zF19e5woGjcSFqvTVy//fj
T4jdAXrvRnTHZBE5sVMSDv2oE2LT5wHikFE2BrNJVwFc4yTbRvhRzXnjpi/oF7ZdaMrA5AUhp43J
Hd/hOCnHuNoy8ZqrR0WIln64X4PJoQu2ytPFFaSvzTq6XQqRy/EG/XxvwmH0cdhMg5aHEJU1VMXx
IYAbVt6IZO/DjGjRjrkVrQ4VFvAeLxjcRXwAy8ZOGrG27MpNhHBJiR4OqgntiPSq5aMRBSzRMmtD
ekciNVwhkacuqmh0EhXS+XR60omw8MAsm14u7eggHeCe04eVKLq6++1QKRT927qogsBhwbUAl8Tj
lT+/Q3PGuBmKOi3KWwMIIWGREzFPiSG7uuvk6885Xg9inuy06lBvYw8pWWbb1VIxi7XOBOIMhoyX
8ZthYP2SJVNYEaJ3JbS7iAQs/vcPL58wXP7xGG/FQLMbDTvvHWpTjcU4Rfo9BNS5mrKpSocvpxrO
izxKp0E9nrZp7STyunzjRUvb3DGvGg+ssZdGTd/8spt3xv89qICJAyj/jqSPZXW38/H6BVOPdf47
vtu91WL0sVLbXUX2C5OTW+l6139F9JxL4gELtvvCxkNtZZ3uqmTmpSjiQfuCgpirtb124KlkxAyk
6WahHKDVxcBCQ4Md8XYPhyKkf/DTiuiNHAKNrilCJmpFbbJ7eaxahZWdT300SGX+pPdk0jA99JMe
ffLU8JAmCzvdyOZJTykgmUrcL3jO/aAY6vLpPMtvAs/lKGWObx29A0sevkdKZHtU5o0WlUvZYKek
5K0P1KolmTnjQrtSUVFo0i3CNjPXBWRsMZD04OsSxNRGDe0FUf7GzWC5ccvFXkSq3hAheQENFJ2g
jg2Uwmh6JN+/ybBJCKTHfR4zDsNhgkyBYtM4t4XrbAuADs294QhzLD417uHyudW1yq+1c/5gn2fo
XtbiacdJ1VN3zWTzxNCIo9XMBVGDh7umCIV8mbHMrPfGWiy8N3kR8NxXAyukuBWEixJKuaEzACRp
ma3QzfYn4ilInxkLH4icn/zr2FZxKBGANfTTu1HtA1+UcejYM8gTIl/HOMHcykS7+GnJJJ2g9PSx
CxVL2QWNeR+atF3k83HeeYTFV8OniGSBrZh7Q+z25yPOHiOPBXwAi5d7h2sbVjEGyFzctwtyHFn2
XJAmzDxq1WgEuTOeE7rVXGXrtL+1XfslB+/GQCcrONcsD9sQBYMVpIIucJYIM82urO2KOVqTrk/z
hOvku1fg7OpUApKW2mxo6Pubslj9xviJv6YWcFrvX00Xnz3pfeC3FgOI6O6gDo1e4iJMOdDP8MVV
ltDFReDE6LUpaYCrZ2H6i5auUvFqdzIOsl1MrQplG75Fo39s3G/i/w5Yb8ZJPlsMxuiylzdFNAN+
EJ24QDjhgXm3MrERQqzQo//1KHRSHwWiE/PGf57rNBMSCv1S0AHd2Lc4BIO1I4rfw/dI+0OsVlpC
lIVWxCkoIrnYngBFc+iGXBipxRiRz8zlihlkvreYuAFtzp0Po+1E4DcukAqEF1nV76OnC10/l25Q
fHL2w0/8nKJTNMgMxbCx4pXEHhB7v4sJHWDU9UO5Gpf8+iS0bdn3obm8tAKhITgM+ZWtAYOhYhHc
nubCwoK7XZ8A9a0KnyBtX75AAgAu1QtaDv3le3Kv964PP4YDKF5vllE65VhwZFOizPRf1CBjT5me
cKgf4Ev2yuukrEmxB5uSSqO9CCbCiw8f27S4Idm5AWfjY3qfl5C/6XVQ50TvJUATjnLeyk6j1fdi
WyU3CeLP2Cl6b8auZC1adQ5MW/bbtDx2lucxD5X4/zoJo2mQRkVDLcSopUOYjhTOgbu1SA3ncvMS
hTOX7cbsGbTglRHRMY9FbT2rzbZoZtpZVjvnkGPPmrMsqpQgSZGqvOt/pyTMYul1yv+6hb/RLsvc
2kui4mhB7MZYCI7wVrYHsOpIag932vIF9gwo1wSfQZ334pMP2iBoaF82t0gZro2Ag38ahZ7w9RG6
J+Y2a8iVGVXZCyYwEmAIefGY89u9mi26aT8Hv7kE5pxQs4el/DHSCNb5GfuA3KEsKhQfQIknM4fi
PNWn1wCvDPYm5p2pO+M5HwUQ7jrE4Nl5Gdtzy/sXBJ1gIKT7aJhiG00hJnHiSMbz7OWzY8OU/jcD
Wm+jB4n0ZImviCAgUUNPPvF52qdKrDFfK52Ww8MOOzV+5oOyiNUyXZCN2zjHWfExQoX3ssABBvjK
zeVkYDGN7e5ONFezEsk530zplt32+2gp46Ms4kPmbTKOuo/ZomLXemNAm3KjCfKaRTCukyxm+hr0
BXyWexMqRIAIYGigtYd4uoLT/KnczORvodqXwMonbuNsVe6dEzIA1e4K74dQ0tFaqV7YeNK1xTUg
+iuUeyAIRKgYYhpDCs1g1Bogh78bGThwnU5EP7gPZde8mIcWC4JcBYbXWiChGlYerd/Fqc1/qJ9+
sPjJISsyvz2/NOyS9+zdQRbYYRucaVBsO010uxE0mMKzAg+NPcc7aiQCL9fStu7rqyBPMeefARpm
TM+IJhRNEea5oYFABku8OETt79Ed/NIXLTmFlPrqW50LNsVAXxo59afj6LpX+7hqKFu8cTw7MifA
3KIO9sDmSJxr0fREiADwVHinVY0WuTiE19mubCBF6runI+djH3d6zdHf+jqeicJdGFs1RbsUPVCJ
bpa+717SgwDWopTVhzvho0zVXV3rnuNzijdhykuxZ6RR4Puxkahg/QprbjDjUmW44hpTDcc78smI
3DWTEl5UxKH55jVzrHVq6ZF2fceNTo1Jf7CdBbJhBzZJlxIPBS50GOLPmShlwTjBf96rFW50AoGf
LYno0qdx03fWI30NAQ+yhSyj9a3Q6JYGQwFBmhOgmgbl0t1nTEI4V3YACS1scZh/iBD4APuQY/2G
qANjIG/uCp3iRtHBV2jhNvhiMK1ed3oF+A9X+ZFfL5wiKQPryavcXRRpViW2RjOewAMOMPBE6X1p
eVN3FLHDk7iVVDUKfHikOKBXOSzGtOUOd2cSELDs+ZvZ79a+gNwEjbrDUQpRbpCg0r8QsOEjB66X
WvrTonqDQ3pCLb+BvBjOIzrm6Muc6plCLpFqr8zge1MGwjutdyDrNTuRXPRMtAzxJsHnuDni2m0a
NZq5O76rPhLYQ4CuYSMEzl7K0QjWqouIqNgYZaD8thmfqEiYCmW2mi/Vo+yO+b50/iUwf8vF3r8+
VTV0EHqG0iTE/hKLwMnlXtT9FITSqf1haR6iPS4NQZ0sSz/IVdFQirjhQ2ix2Uy96csniXFMXZSe
JlyYbuTXF06g/5wZNIrPAsSZhk7C4MZqpUHObU9yI3CL5d8FtEDQ1lZMDzrccvWY8pygEDUfYc4S
1uhSBYfNJqDiO1PQ5f5A0EqLA9ps1SMQXJPqTCmOy9bMJ3V2yW3ayEo+MBfV/ICaGxGHssH4CIeU
qeM5iASfE3zm2TPkLlGsBFKzwmpNESn6RQxV6NUM653uN1f/T4V6VW5rWmjLKBLyzfIkkVj1bUeY
btDJZ41SGprGxM7+S2FwyxOgU8aDWlKE7WrAGbDoJWr8eDLxjrewSDjQoBLMWJHmIG4HrsAp12Vj
P8uWVnFCSjoX6oP+VHw+qr52xcrNAjq0pu3u00+YSq+8//GjncVd1j+KpmuE5x7jvQlJuuMc0KrS
Az3zxfnurLmD5gfvGTn4DBvHOvAk7EB8uNOI+LbNsNG0cEeRGjnJmPLOrm2orqyW4GBQHH/c49m8
zzHcQOoFwPh13gWWXtquzP6qCy+OLn8XJ2ElO8poqJV1xZWPCLXJKYde5n60V/2QgBLm+nt8w7wT
36TxoeumGgRpRww0pwD/tzE7ziR7BL+0Dnv5n7BDfSWP/pz6ijmkqFbgXBAekU/alBPrIrf9Lxzg
OReQjR0ylFBUUP79x3FsmYXILcl4vrvX5cOPCMFMsbYNIBwYpPET23i68zG6eAD+r6C1gJBRzY1g
O5QBAX3oIeEE09Pp2DoHenOz359LfflKoWmr/PcR3unJhFJtBN0Cavf3YTHqQwIQUsyLOs76ZsAy
5M/EdxSgF+OzpKrpnCSlhSV2XgvM9yocNm+9JskKNMNK9i/AIElhMeuYArQ28En0qAXgMyKegy47
F4azVUZ/9qWzTqtUoF0TcOhlSR3ckwZKNbgsP4ulsBVfOo8LZBDL8LYBGzwrFMtgSa05PT5MeGvA
5ETQ8wT/PmmUuTztOrjH2XRDaxo7/PmKonkuqTHNg9ObqUflB8t+DwYDzzfLpHhCUKgGJxPzqGzT
wrcHr3aVP+fAwrR71+h4D6bi+pG8rN3S63Jcfs9h9tEdCdj5VZj0wJq7U6thA7k9L6jOBz6U0bIK
ad86KTtabPLDt8ZJwYBPYu3NS2Kq3NOy1HAF60SPvIFgzBlh0+vNbbxjNkyXivbhVFN6NQz7phHJ
Pvc6DhFFK91xJ0SxoqWxGAWK8o3bDIoeBruuzCtUFDlXpgQmUJ06m5ObTCyfTHcZZF8eHJHteRYD
9O0ylMtVa4F48wbQZE2imRDvjg9/r8NWNLwcHLRH2d1CXC8l1fojd0+0/yPUWJlmo+pb+E1zUHDP
fRVg2vtvv7JB0zYwLBmaf4an26m07l2t4Fd03ez6b4eqJOjl9pwbNq//4c4ex6/zfNY+qhN7/R5v
NtBRszOBH+84p2vrAM0dg9RD0q5LYb7CncIlKvKsEMv+MMAAiglApsT1rKxojrrQ6kA36LaVwJBF
000Lrjif6qwleDzps2OfYN5JB5vkF9C4VO8PdgZR1AMxfRIyuHMXQlDCGsM/PPSVN6itZ7LqKxGh
C9DCv4eRNF7xo5tv3jpOTljOkQfaCA0R36sx+qUqA5BXXt3Jfs+l/9sstH2MalG86SPiIF6XH30p
oiMnbsCrD5OIG8iHM4Gc5y+t0p21V2YauADQtnNvE44GSv5xoJRCCbghTKVNrGH9Cj47nBlqv+QZ
eKqW+F3ILSi17yzeA1a4JdMqrHqUfVo6R5hXlvTqnoBS25tnALS0iwwKdH0MSvyHIPHUKlF1m8P8
NnkWVMH482Mt8i8fhNPFww+UgM93fEjINqKTfCUe7IpldjSuLr8jWIKnk6GTsr9BpTH0WC4kE6PT
EVj3hj388nXxYchzt/KWR5Clq11Av8RvqODx3TJpbn6vX4M//zvKaNQ1GVxdy2s80/JuA6Wx+Wle
FDqThazE/EM8Oc1Xf21svhsDXsu51TAfl0oKR2Rl+0X6gDi54azG2jn2nKYk26E9uj6WSKPXhOLh
eGPkoKdAvwi+K6r2/H1evQVHS4h0J9RrLeuxn7fOJ/+vHJynP9uDheNes5gzWOBAlz4mKESYKPaI
B2TCheo42MjDu0F7vE6heE64eiGbkkrvqVQXKZr+6YadEQOBAQ8iHWz/jgjfq1Vn4xnUpZ4fOTOD
IoNnDwEWKOKk0xDxcDwksWqovqYILbd59/yjHIURqCRgFrKRsbJ9j2rKfqShV8zfkIH8e1GXad1O
ACIc00wRrB/qrvJMisyuKcgenecENFgPMa6eVk5FIz2DM5u5vpP1I5EU70JebYGBPJwjC+2odK0c
7m8t0Zg0MYkhYo6n7DqLy+bWhsiaRSi3iK53gcpPuKQKYOMOOBEOuf9IA5jdwKROo3dX3sgU5Ien
T7P/vzhUnoRIp8nnp+Db4ol/TXJHuGujzp3t771KM+mPicki2bQO
`protect end_protected
