--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
m1QSX0NvSKFsBX4ViNaneG83+/Hfawd+AEvP2ODOKagocUQDekiBt5pgTbf5H6hu8+HKKMuG63iM
lUuVgW0C+efNP3RM3PnR9Ll8sq2yrOHTpuT4WNUCRDIPYtMtnJghr2IpvbsQYhrSiSUwXraaOzKH
HnZT2IaF+wN2Uutq5mouXodyVeXdqUkCb+2wsuWZcKYQgiwOD+DrtnmRS3sqpw04QTdBXlprsgid
RezP1LLCgd0N+drRjD0eA0A5Yie6DX8G5RzG5XBWObVexCqqbrKkfNnz6rIAqvj1fn46Hp0MQLuB
jgf2lumGaolzIPzYne5KkoSk/hzFOUBOA4b9KQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="fAYu3SJMQgoge17S3k3+n/F1Ybx+nEPoDBqN9kJesJU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
EGhHm1GeRM9TtdlmJRLTt5zigl+3CeHzuVnaz9Fhz1rV0CECFzlXSJHgdcXhHvMuNzSLWXGsJ7J5
qhI4WqgZn88Zt8xgdpCAunsXnrUsIo+1TMOnuH06XAhF6MEdpzktB9jJIgHyfA9FlbZE6YPd5fHb
MLEDP14hm6kvr0OlqEfyafg6YljnFWkBKtnjjrqOg93eJvWxvCQBBdbaDdVKw1vT6uM5iFLMSy4p
PxBRYPM/SEe0lkbAurMH2mFfZ52uptqe6j+0pEmQ6FP0Z84fGn9G/5ksdrNbn5w0iutJ46MkVyzP
eGUd9Xv9E6bxlQgAfdz8wMavFxjcEck0uQZaNA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="ctGyJ76cOt6CBDm0OPjc+xsQDOMui6cTQnfQokt3JPM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 61728)
`protect data_block
2xDwsOIql4BFbJ/fpHPwGi8Uq+ELZJobjv0EGdPUVzdwPybwtASZcb0rTy7/0hXEtXwavpoAzzum
L31tRihNoOz/hCXy8kl12FVWxqrLEmgLU8oThRfXSTBHCmgEu34Y1Clnhh+UNoYmZDnQ7FTSn/lz
+m4VuH8YsudOm5/khNMeMZNauBwV1PfUGW67rEGKK7q3nWGbMtFMyF9qxio1jSTlio10Q/rB6O58
kQNGlb2iKeSVEXnjb8Jlc/g/amutkWWzo/EvEG+OHjuh/hXvK8xn41pSQCTOr6teXk0jvCUTB0NU
zWgJyDhQVOG63r1A3zICm9o+FiD2vKSJ6EZE/sge8DjQy/Kk1yNW0paTxc7QOQUuU43edQ7Zkb/J
FYldh1g5ls7jiZZGG+jZqMlDfgJRUwMNP2KSBKvcuGPsYfMzNDwAhc7kM8cwyRPHTrKJPD6Zngcw
sVmXZyIUvkSJGKIDAtFqgexuWrWv7N3HJFbhYdoI1PJwVzUhyujLrYzYkxy5w+gt3SJIXYxFShiG
pJ9cLgIyTzn8iaOAb9q6EgVyOQNP7h8UuDHP3G+jT2wKjh71HQE1P6yLjfUWQfnx6SDbR+3BEwNJ
fNi9AckEysVJkdGVal/F6w0DKoox/3uPeXZLR+eaJsI5oQBNejTTcwqBsIM8YZMTRwcp+3ZkCVvH
SV8FeOkp0kVLYtDQZR2HpZQxbyOzHqardkmS3mtujfUChZMhI61U8OrfFqLiQn5nrgNeSQ0mNH7t
MnYWHj83V3jRU2EvgW4g1KM6ZUwoicqgXB1GapxMpYAk/OEM+CwTWf95NAo6IPiAg+sXSusLYkuE
Vg9s+jeMd/3fkz/AYa5yTW36c/PeuadJ4ROBqunjnVyDKy62lZtpIs3YN2/t3XmFbS4PdHaXHyfR
4h2HWImZXK7FEqRuyQ7SyB9y/4jik66jkFhabF2xELLSvus/LfVqdaPRgcIkymgrZeR5xdWfeyTG
K/9awqWnIW9rp2AtniR8INfKJhmG3XCOpS3R388diW65wIDsTNwBjk044V7ROeDaT0kA7URD+e8y
aXQT5b5jzkqmJGJ2Me1kzqS6WtPuCnrq+JwwEjnrlmaCvecO461SgKou3xEQqoo38LPFUWihN/te
UpWH/ToTyd1fLx6rmeXfvwGOm6P7KOM/jTMHRts+OY/x6ektQo1wU8WQMdZVrvtGHqfZoj75b1En
ddp4RCWNoh4fF7IoPS68EibwpNG/yn3e8f2SBBR3hmfjOrnEKyB5/n45IgNl8Bp5Zie3HfWvi8Mu
sq8kHJsvS5dO5d+gEV+HNa/H0yklvlnQxRjKS7TNp1fKtoOzpaCRQ+H8Q+zbUsKZdYenFDItCANj
hRQjzAz0vZ5XPYKwqPHU0Z90iiCidzGTfSA6C3wwz+hZqGL2nAOifMNvCoyEacv1nwyqtJuNMDZj
3cnTpK0qPP0q0fUr78fakQE1MAEWCM/UKIWQamy5Wb3WWIy7X2VJ03ADeCMEz66TbsYhkrPG+EnM
F9KDdIgEz7nEVQQKhnV7ykjGmtvc+Ehp+ZI9mG9cgT0yv00DDDO6CIrv937X8FKrFQu4MJ51S9pP
UOz0AgMdAm4deQx5wM3SfdNF7SX8o1C9/SEppptINleAsUFNUtgEpWlZf498Hv4qfG0Rt2wI1zdd
HeSw5sUAhlMiyi//o8xh/zFhN1knCoo79V9G2QpYhqq06ycampZX7IeEKAN2kbhSf89cwjHEL3HG
NhL1SguEWiuR658wrcHxZ3S2qdtHkPXvNixk6qTIYGCfqxR4nAYZYhCI1yqmL08g3RRE4obhz88N
uDHPkQCC7S/vv3BR4dyu6mNJrcKHpx2QPrYg2y8dl8R7eyF8eoCOpuU1s9bxn+Rp7Tx/4+Pyph3U
na6k2H064DMV3sNQPA9qHRL/740hScfV1QKIHrsgyYreCyamvdWkjAo4xXJJThwRNkt4ayC4aJQw
JXxC4eIONHTZhVx0apY+XqKCWxGcH8dFAekNHSiVC3M5t8bO0h5Z4u9G92Sj3xiK4ISYE0eA5oF2
JZdZalCXaC3ZuZgbLywk1w34qnqOAneZkCbycuwhmnm5yLg2nkxmaIOc41YhhktL4f5lPa5CZRvt
qUEC7pawXRHLmHKnNHZxQVlToQinaVi8Ld6DMd+jbTZPKdPXHstUL7rFVgl6W41r7L2HXJG2gQLi
+YyVzKcLIaYH4uXufdvZJ6bmw1OBnwb/jBwLawM5iWddYbIPCWOU9pRHq/ehbYunkZE6pklqRQxb
oAUQAAlmqgR0t6nOKmyuJaJp9cXMRngnrmDIPcM2V50c+OqGbXV93UILl/b9wQdvzdgmOoNwkcwr
4B6Qr3V45hLvYSKDWGVe15DR2ATLgBnzUU0DJOhamU751zjC2ZA5cC3DDDuRlaCl48QEtgVNPS8G
uA78B2CeEV+BafFY2Az/oJUiWi2NUzVToPB4xzNCq/tOvnChPqRyxscS9HnkM4l/ip6mlzBSNh2Z
VPViMhEwaMWRn5neIwcl33Kz90JzxqJeqbl4CoxM53ZL3eWuVEZXkrnx75V7nxBAl5Q9M2yg6I1o
fBNUhDJd9jmWZIH+zqAYbFNqgbk/6bnzeSDiTq/I86ypiddvM7ytdshteKPmP7G2cGaXs1kN/ADx
MxEh1PtotS9XM4UdRINv9IPXLKR2ru7FyfEagcPDMWtal9OUCxR2oGAtspiXCLIQ6mvNJPQYyA4Y
Vn8boPWt0Ws9kHH/LXkYStxPzJj5WPdd3AGZMYrQD6SOaRA7yn6xiLV0uH3blj8ZpCWDTjlxSHr6
9UH8kUaAl7yJR9ZDKuOWCeOloFIwwhX8mzZih/uIvrCK0O9FRSTiI+9M9Lk9Lx/SSHN/20AwZva4
ynpMvPEezy1g+mXRXqCgLwzdVXbssIz3qw6kh/3YmptkMvrCBgh1bu/zMXTnHwkRX59VDSd+I34j
wZJOBLp3eeoSpE+GaVy/3HhF27ws7t8gdGBpHVa+9x/swaV25vbxf5g97oAPeSTTpV5jrhHmvnt2
CuwG9evVYA3YAcG1fpYUUroqQpd/Tl1GvrU0XEEENloCwL+hr8iQpJAIzBXUTCjRWQIls9SsjkfG
ie11OtTeWuZ7pU1qVcV3GS5cvW7tkaNw3ru1S/IjYpM74AAlFYz924Sph54wV7eggYcH41NFPeoT
V1WFTnT40Qoszr5dmUkbhlWjP85aFJ9fHJyQBeKbYTLva71u7SffkxI2UXqVEsmJduyMQphRuzPJ
lkh0p5aDUXjA3w1pHD6G9GPZgUoqfqyn1rBb4nGvob/6/ltThYZ09QknJDV2rORDQZ0hu6fNIZ6R
0Ao+pplagVMTpK0mSMf6snju+QMaylX7ggMY40wPARne5zqCk5bJJVxlQgt2U8oo5tziT9F8P4bI
Zs0OU5Zk/WqYUTijGtRyG2eBFxJbbwAMx5f2eRZyEjyn+4HSduxKTaF3ELOIYsBmyiZZb+ZOJPvw
CdizfJe9U4ufgI2AjDH+T36NU+o4VDXFtJ4KQKoHU+xu54suVZ2ZT1mF27fYwW1eWKXu1e1U9S/5
uB5E8HGzvkc6i74c6nXWVnzM26lsilzb40yOP2RCuIYaKsRjAzjE2koPZYSMTcwDRYdd7hbl5tNY
uhUeYgU4WGapBhU/4N3qZlEIufeb/v2sEWTABeCvTAy+PrbOUjdB1w0xyb/2vUOku927CLBdw+46
ZwoVQpiBIsVwFTt1U+A9g/qBFCZeicclZUcn9jkjF0GeATghRfCoz7Wh3qM6YgNdAS+fPGReluEK
K3kWl9APFuZqEM1J3zP2Eq1IJQMoFIuO4j3nruPKZr4j9+K8FfFv1MF4ks1ZU/RR8wMNEuAEDetJ
xrtu4j6bHVC8xWzLvZz2tkR+a4by/E8fEqMhfpQa+sTemwVxv1Q7FViSl0JYqDYzz0SYprrH80TS
2v5yiUjjm9U9yOTZnY3eH3I9xGjrwDznFu63w9BB1fZMWYMGlUmubbDtMYd4ZNtoM/EOjd4n2kDA
eAF5N8tymOEDrGhDtYzULUPifBsfwZY658jubcIGMV1B18TOL7MnozZ6/M5tK/hutZKCWPDqIcAv
uia3gFvL93egzOk1xzd5AbFZ9SYeF6MrAGBqM2ibl3LXUXL0Kjf4qWyAzP7K7G/4YI9zcEa0dXdA
iBkKzJOwLhUZZ9WRGmTWVe3l10AXMGzlyXNP1GNNl/s8kXpmNZm7k7D0r0oE14Cv59fdXzMA1Sk9
qQv86cTBlrh7KYALvD+OEvG1wi2rPNj2b2kY/2qqy/NNNmk/HCF1E1zyfZnEcmHrz16xtA5HZCiA
n3co8FLcrZw/6ECeJOEsiXn1qEJE/Icz/SrbzMcWKDz789ppfeaLCQwYkJy1qV0oFtK5YkUcuaz2
tRi7VPNHYtDh0Uiopu+oHBfk3uafp/wPHQVGlm6Eyo6Nl0ywQkmTLG4AmNmDxx9m2J2iibWyxiQD
tPYlbeMpbUFBymo2K28fHhyRdBUUoaPjL9TVpfE2KGazzp7M1yO9E+1MsX7DKtYLnXF9vte95rKF
XdJnK/StspstR6Z8z2cxDa8bVYWJEGs3i33eB7pYNoSfKJrCJiHu05hUjLB/X6+2Yi4k5BD6OJJT
3ySU0ocG7I8Lnv/Po0TrXqsMQjw1uoVEFujErib9S3mu2D4B/yCo5D3yJQQ/CR68is8zc00DT5tn
NvkoXqBu5MB6/am4fkJtRwl/jxA0FcvdJWFX3QQ1JmBUfQfMdQCZYkWtpZDn5U2eImY5aRcvUx1M
zbfd60GtQ5kWCeGW+rTTzObtjiMCqjy4Sz9kLARDoY6tAiEEcJQOtgp2dkku0rOYE6L5B/ftGz68
lAdqotjot1O/Cf9xOgxXqKmRzGoH43abqLt4umsDtEWLKilIBTsy91rpujx0p6i40KqB2ULV3SlT
IXKEhRFDKQNatGe/WCnIZY9eBb30G2VvGrrVHUteGMdtQB5fcqzHEErot08U0PBbvwk7lEFJgNJ+
QZWZb66p1itLhYoQIbAm4mWCdeEB83+HYK9KsxD96bn5g4i2OJSRT1HZVhYwu3BGudtBXgLe0tgo
jsBxK8IM+GGy5PQm6qrWMrLM0oBDF/29VNPTXr9OXJO4NWQH+KE2bEGz4xbVhCxb/7uohJEZDf9p
iYlwEnH+XvGB9UExdv9Wr4M3pNShqBwG8T80O/00LHd9yjl1fY4QwFKVY57jxjQ6DK3EyVpJem9f
3hKFtF9m4G/naTYtX48bNZrq2ErVWcvSGndPI30lbLaQxgVZpCrluptWHBrU3sElf5sQ91hWL4eE
LhqAVcjdcPICj2XNFjDdsL+/6zrztHn15tUwO3Zf3Vae2JIC1/CafwB1NFnPUoQzE8t6TVxIWqTl
OKGXcgypk7hPMr+NORbFMclgpxHX0BsFWCYq4/MmWgbeF0tk3H/h2sesTTjP+92uAq+e1I1ArORJ
IKsf+xFcFSWOoCF/MZxGWPdOPDoikDMxqgURNrld8FJ3QesUmZDApdgsA+b+z4GVsrY7o1IvTWzq
Z9lBnEw9vHKac5DqhVddvw5LvNPDGLhfa3SZ3sjKBchqg6LSwPZwnF6VMT8Ma61g2anaZ7pR2eFV
HHoqKPDCYq3cMcBauhb/Vmdg+VpgwB4r+VTen+qrHYa25TPN3S2S7cCoN3ClrpGRJ1huF7gg+iX9
b5kpF1iXkdNITvFLXd3zI/YGOdzRgK9oTb19C2FBeKbg9fJ1r9d7XyVDgUnnCfZSMM9IT8MXsXVV
kFKphuDGV4//R2MbeU0cCNaxl658S3mJcLV7wXCH7wuKWiFKKu2pvDMOuV45V5KWO1/7UPm9SKPs
BHQ6ONfUthkDT5iGMMpaAOEo2BdmTC/em8cYpMFj9DWa5P00a4U9I9ZRH/pLJUauREoRa+iXhZKL
caTWJQQMUamhJIaKXyaMBd8RKQph3WjmV2GYY05lsNsaGIY163bSaxr5sxxI1/1NgZdMbrxcFhpi
n0zDnr8kU/ZkdWyczrnpoBn61e5EFb2MbhuaGCVRwIrBv1tn/CFZbtev1HzET+jAfy3phIwVwch4
w/SSgYHQNGVhxeTSXBQgBvI5KI1Qzv/MvziUvJ646GrCbEFpCoDQ0ZvRqobyMgaElBIOq4BGCi0R
S2k4kDtBbdbCRnSwYl8y66NR4NzYYGsaP90l+RvMAxKbAf5OaJDfP8N/U5NsdgzHNLvPm+UDZlYO
DVNA2+eagt+lsVG9mXYEl8odliIygfkxj3kbifb37UPFp9smD2CPNr63kAOEnSEJqA/h1f5ae+Tr
yqa5xRPKWlox8tWlPf/Uv2N6hbYDqI6ynvnZAkuGQsOaYxQ+9786y6eLLwipzIcj9iXeju1kmOKq
+zcboq2vKJnoW//0ivRpYI4qHMLGUz8Hh1H8Gs80Hpb927OfPxEPpLCFykgbBGWUshBWCHPSeCEr
2+koFxOU+ysv8ArzqX0KWv9XOyzdkJFAX0r/Un32lRCf3H1oo/Qdwc3XSJZfwiXLJZiyQ9d1kNQa
51UKlNvPubMDvrFcLjp72HVRlQO5itA/aKHjtJkLQA/GrUkUlCIb4Gn2p2QzSukZfo4tAzXscsIk
YVX2z5rFDcFj0fcf0wWzEKKJEn5CIASJ8GaH4VtTYPaf5jdFjxq1084inRYtsy3B/CsBLtfFcNwT
O85h9OZ4XGT8RrE4A/EeDuf23yV/3SqROK6tC72YD1JdqQpuZOnqOAr2Lwy36mZHGiWp5RPpNbr+
DEyIqWA8m1704F6vawUq0en9zeNFcBEDUaDy11Vm634U9TVDv7JxZyxFZyxZQx7cLgSgobGXpuXh
9lhe+LsquxXP8C3OR4Tf+JCBSq0MUXHZxkkzJbGiCn8H1NbwRFt6uK2rFNIvtzi5qcwW0RVRApdk
aV25QKqXzdmrCo4SvPuZCm6V0x2Qn370CT0iyVFoO31vIMXbIidcWMPlsYW+oogKWylJT6jj3Uif
Zbq4oc4UdzASMZ7cJ4e08Mpc2O1WXRWlwi+3IlB5x1Gv4RxJso8d4/Sexpx7zyIdxx3e6QvkOTy0
0yIVLxUZfa0fRk30P4mI2w4Q5UqtlINms6VIur6SNgpuQXZMnhdP165bENFwCjt7pWSVO0DbU14x
QJoOkmjXn3QOeTCDXkoYNFwssshCJM2oOrbm6KQqjsjBgFNItpnGOHgUuxqNtqf1bCODNMnFcSqO
y59i255fbedXoIOqZ6Bal7hoHRQwevmjXjAJBywoxeNmDs5VmPPg44Bf+49NM7ydufG7s8DnHWJU
2wtTPUYOdxMOvizTJwAE1/UVnYYE6b4+I8c06NlhuPDCZtOL5rRiTNpmxzN6ZTeZ6njooBpxKe5p
4pA8OK8x4Ioua9f2P/ptpi3bCpk3VDqKud8UL0CkjdIW8BRRIkrssy/JNurUfOcX5XBw2UNd6L4Z
cDu9XJhVyWYnM8Dz+s9W+2WPbuNxBntDE/7REaogTQsu1nHkevHvuYDymHb97b04LlWafFDllteU
ooboRVf4kyzXejyv/hDlG0WWyfSraY4I8N0ldjWFMlC0/VutGhjxD3zqmwcs5RVVzBHvOkYcm5xv
z5VMz2wOI3mlGEEbTswadnvnT9bQmiCYibf7w6Xjg+ck9yzzkWFqdpF2rtcCGcaRIEKydKXJiPGa
oSSUdAzPM65YQuk/tk9maIXAKoOiS2Spkwxd7B6ehK6fFMUI3G/7DuWz0DfgWKwbkQ3xKyMUX9tv
+9x2g41JNX0jodm1Jxk6csrB674cOKOHPX4SZNgymW35dCX4F+XY7usOJGBQWZZonj8qXa49N7pi
6IxJ3JEKddjUBsUFDMxjYJPDWfgnF5J4L8otPfQhEUI6fnCV6PWbiy+5pX1CZeEFfGiI0vIdqSMg
ypaU3Oy57v8fTNymTIeMww5PumhyRh0u0fuGYN3+0QKH/AcDl1UpchmeLukCTUICHxtfbSGc/Jr8
TmKwG5WsctH6OItA9K6AYQbmrQD3+iHevsp18hu5rgJ9gjCs8LkxIwxE9kvApNzP7/ANi8FxNdk0
DVmSZ6JSC8NvrvN87HKuG3sM9jsvZE2xx2mGaq4rCgAmpARDU6l6z2pOhSLW/geApu6C3I5v36uf
DRJmZVqG2ZTisdCzFtPMbo4fi4iROUPojnbh7BTJ3gartDcPPGnxiNf1Wx50uTNjb/q1fzq+1YTX
BPBp+0kIGP97uk6+e753Z+LZeGwf+PNjMdeMMcVUGVtWtO+9Z7rwMABWpzQG8hF3W4OsdEO1fkj9
Id+RZKDfsBaixkss3PP7x5QV1ZCdvUvGmhF0Ie4ploPJsoSsilhSt+0KpQ1TGQl4mFDRn8g1C9jL
qHHzur3FWEdQ8ftGfcD/ymbTF76qRJMArzZCupusG32vzKZ8II5hC9IhP63VL3Avirip8P+Jmj68
IMSNK1ZfY3wvI7A7FLg8KRcE/kni6lwbJOfu9MC8i2W0eewxPrkv9UtIXPCAF+RmJ3Jjd46AENLl
u7rsQ16DugRnO5g2jL/vMvyZUr2cL0Xwf2VipYVk16fppCa1ZwkNs20u9aoS35t9x3Mv7e0Nueqi
VU+094Q3PiGYYimhjG64cDK0bdGk3QHs/erkqtZdMeUew2e3xxz4hYuXUREFPIcMeglgFrHx4Zyu
RClri28MFqWDpBuuh6umJ4qkze+ZUr/XhVyr6wBwXLVooTUv2cE68TEyc0tn9UCVxgxaeJa8jBaj
y1zNLjhBHvNMvS+ku+dK52DSFQwSre+K7DW+yL7cb7rjkGJSy/N/QD3sh4WeTdVGYABc61esxKJV
TO5C+3GTO+p27aUt2p1RrCbYAYnpe+KLXkwpmzpkR8qg2JJwqyPXKUyzQWuxT7fxmTcvRDHb0mw9
w6NqdW+BG4GP2uxJFPm389pN9Bby30KKiyUoh8ZQVt7w9HjjsMdaa9u12N3e/vK8CzeQgnkF+VoA
xRINElk9Ke2Wm+heCCK1zN/QyQWWF9UovKMMzfHMzZjpOt+X5A39QMBSe3GQAOPzo3futKQ43S1Z
7Lxw4DpxrdQ5Z30U1SyJyfFIRXcQZ296oRUxkJEgN10kH3lhd6j3bBnXQDV+hRj4N4Vrafx//k08
mZ0+L1eSepUVgnnILZs6/uC3Y8Eow7euys35V0BwT/0+HJZGOb99eyd/phZsQ/V3huQvwX1lSfMI
G71GrIy5GSCuhzlLYrhA6IiXSNqDnU7gTV4i5478EqixMQ0I+pcGasKWpFz8hGvXsy1kzIoK1E63
smlDpBIDV1iq0cYbWIJ3IlVCTJHsqUMGB0HdVBGuMeTkE4MDc17DuST2IEYuR2uF7QUq6QOuqmnM
uQaw9fLqoD4rnKz6aTH4xK5TjZn4/Fi1RYpFMqBkMCk1tvH+lGW8We6AWCa/Sz7fIMUklipZ/ZD3
ikd507RIZ8/5TN11Lg47zvlJtlr3ZFZvJcjefYfzibbhuk8EVeyDsqr/B+VGlAlngcfADbK5cDhz
KOeWcWjnUkWiBc68UjNVpizkBiEwEgEJjMD7JRDa7IxMyXpZJPFkvEWBkOce7SpuNCGapfUBEDFD
3iMEjDqHkF9JOuKQAeC/zfQwFEWVCRDUFrl7UF43XGIdFblAPyBHU1GXpIMsdJUgk1yO4z9Pj7Zh
ulD89/I9wozFDXJGcOkt+jpMb4eoMXy6+THffjpa4b1CwMNdtJbtgM8bgna5qu3XfGASCH75OrfU
7RMW+zJLyT9ilfPtqFp2UxTEaOusSIswSDNyM/PI/7c72uAzTtcXRbpZwXd6SV4S5vSZzFor05ED
9rJGWnxIkAe/B9J4pqJr5/W0J5EiJ9VR24W0ewSr7nMvoaVZ8wQZhFGk4Dmg5sT+q0eqlpxG/Ob+
z955aw1bm70LH28zQoPnTx45JlQdM1C2AtvKMw+NNqaQxC4TEWFx6TQLn3cHwqvkDG0XO3ZQgETQ
U1FauHxGuS2zy+4CHBnFKdNgEiJe1Fsu70+Dhn8OqPRMe4WLj1EkAIG2S4teCJxUBd5U+UQ8ikrl
ylUhm29MDfafmnKi2ZjupaHjhym9XW4QGAsd5Dq95Hvy+qEkvpdV5iwTpSm9vjOF+tJyfheIZBHf
GNK0vkKlwCu24Q8//nulWkBoz8bQI3iKK0PmZFMVkmP6KCGKXfO+h6C2RGgG67y8+TObrPoZMugy
siiD3EirpOfG8gv+J8p3SEomcJ94qrBjRqNsie6GT+Tcel2wbk0G6kOjk/r+q5MwI1/QvgSfDWOQ
iRrKmZZIOfaSu9hIz3C9i3ohndNeo49rjs22wOBgck7CyvcP0UjAIYg9HN+O9kSiHdPQnnc1ulWU
a6RB3zdNBMmeT4DOaZeRbKNFs0UlfvwXW9AwtG71RY+9VI3Q+nApu0hf7oOkQN1fUdUU38zwrioI
jdgaebuEGAx6UvK/B4SQF7kClVYX0SGWv1dbWsDaMGeoONyq0oN9Fj+2tJGyYgOPaYMLuisiCdQf
xSy8oGdsjJt6dvarYSpGY5OkHW3S5waH4Xdxx0hX6blpMVZ5gfulkawR61knxK5SJ9XH1/jzyw+q
P3noyIJvoQpbzIKZUgNZGlZGcvPcIzc4KcniYXly+riip7y/xcfGCIvCCYWCOJrVk0PwcJE8uoW6
iOuO6+mZLaR0Hjrfr2x6AAzfyyHgX4/2h6GcrOdKZ8OY1VqLH4wbvjNtH+9jFMtPEDV7EyZ3YN90
zM8gMzLaIl95Xwh6bgxc4i4yEBBANX1gkEyX1LdBKH08Kwa5lpacHwVnJ+C3CPiPCv1Sn5XxXBOh
8ZZm8+dz3k9jb61QyIX4OgF+DO67lp2POlNoboJNhC4Su+C5tInZQIVhAsgeevGhV0a8NmSFmuDS
g6lVf+9sWdhCGIBHf90zCdkZnJyY5jznRaHSBNYhcZmFPjlGuTYYWdq7h/IQRwB692Fp2ScZQhyq
71mWsDg1a3s3cPnp96733yKG84JeIGsmFo7pySvAcwMmSRQuorbW/Ik5pxNvLXH7Y1G9M4qt5o7O
7hupjhRiQGiajK2kYYUTSf1xfu9G28jK88xkQOJGKOppkiulMhP2m9KYpRd13vzjGTyVDy2ajkYH
Y4UWY0dezuo/M+IbFyaGlh4tfsLOSe48l3b75pc2m+NoKx3qLCufYcMtAEHUrKcThng285GPyLk8
SAQpyCUu9lrYCenzhjYrm5WZQy4f0pRWSZizcmOdsdaDb6t0JpKP8k0hktaR7+5AUUNu85uQk5B2
RRyEXpn+80aTMjW2h2DERkj3lvMtIPQtaPDyX7ZTMADfF4emYkDcOi1tyClb5rXcRQj34SDtQ4oB
P+5FPEPWbyqThjpg9e/Ia/NTjP/foUXv0z7pIVJbs86ZOMVxVNVTchZv3dt5s6aCBJNexRBwMX2s
qOXLWZP1bBAfHa/8BTJ5BCKE5Phymdn6WSOr63db3kQP1MEJhAqV5qHPTEWRpTYEfnjtofRa1AB0
plW+6IGCGUvy9VHbXX93CxD6AnxpK4z6GWtY/plag/tvEFT+hJpmnR1AleM0tcG5e4EYRqUOwC2i
oHT7nWoHaKH5taP5l/cKmow5E/sp4a9XLjlB43K6v2w+Uu7XNIcJNa/TaAdILaMhJH4XIM9Uj7RR
xyZHvT7nRJkY/172Ua8pnrMbYOVTw7QkMGJKp0XKIjEWbPtb5ZqvE4+epFmZPgCCl23PYKPALEU2
aAhnuIZMEsTXRXTUWDGhpGOr/JsrKfwmeIS652nMpl1H+U8DIs8SwloaoPaJvQWibEYJK6GCglJt
9uq2/l+xu3sNlEYYysvJ6L4Q6gw35yeTTD+ucKSb+1mYg+cBWcB72rckKkS9P6ovkNJIZT8Y93jG
ezkEnozoc9ZCo91sWPX+8NDtzFgftJuQgCUEJ3yl5ZDTfUWDiDQzAOr+Q8PhHMVG13Sj/xoudvnV
PaT2bnNbfmCRlGxHHWjooSjL5+NPAXunoEEDHRGMJ7UMWcJPagvR4/UPIrS7l8D1TDtjPLux+sI8
hOLoO2Z9Veq91b9qvlXSD2zP0j8kbpM7Sj8VfAufdP0lpAWGoboA3wrAXMEJqWyWaOtHz3gavR+V
ZQwYWTYbcstKGB563yHATAM5KYuvF76IGZA2qLqlATlL/h6Or5FsUtB7fCxJVTdUh0O/mCjQG3z1
qRF2kJcmsJ+mp7d3YsARACu3435oHFDxz753Dq98i1hJ7soR11YpiX0c0YfgjB0z5Mps1GhFdU9J
s+ZrDmImcj8/9+j1vJDTTmRVKpjtSyjZCCce4qXn60hvujbSG6gr8utBKEmwYaHYsqdvZHbowHxU
2nIjIFKcybJpsBgW9lhX43+NTJrpoU9bVpJbnK3UElSZVhBT9vNR322L46YTqx/lgPPLhtfx5AgO
PbD9R5FEjehcEIH5HZeZmdBacxkaYpnXVXW3hmxmwj8K3ip7eZCnTPgUi9yo4kLAeiHMfcuXGK0f
MkP58+d3pEgawhApsXjoKGz87IZuVDyB4oZ4kn+eQWizC3J18YQ52aBHUSbx4cKOwkr/8w2GADMz
Zm7yXRUEOhAY8/tN1XbtAPlfxvDFtNLBy6L6BoPGoTvpYJSufTtBqyqp9CWJXxw2mtTauc6A7K1T
1FN/LuC0r+ZGozmMPucJRIwtYnPqrFReji+PEa/6nioOVWIVOItive9ZZvfTqzHkagD1BpqdeAiw
D2xQ3CO40UBYydVINT0wAg0Dhzj3A8TpgJgiMVlvKyoiWpMIwgdAwdrX20ZIRHDklqkWYSPKhQrY
Q8jmU+hqYdtRPZJW/XeX6jflp+3UGojKFVT9GAqj+ImqVNEzlzKiSfOi8jig1o2AF1/TXVGnQVW4
NeW6niSOFl2jFmMNb96L6QK3b2EUFnuxlhlk7eW71z9nP5v57fl2Ifg8cS6R4+j/MCvUncWJig7R
2C4+8xxvo5FIFHAv+UpzGlPsKxv1lNuBbvJwcTW6Sg381ZOY1OG63/lhdTSZdGhg6xF/JTUz3lsK
lu53uxN7Fh4srfdAUIDCyKfvSGVLbVD7OoX8MCTFpRH4ynQrLyUSoclkyVym7qJveNR5V7zs4RA7
znHnjK/NRyZsgr2SldnvGHljtN3hMsMjKJIvluwbgSyydf3ukvYvZiqvBamJwI0d/BBcz6vTZTtW
66XDgjXk9Ea26fgrNTQCPOoyEHJ8aXFJ4ecVsfe9T/IvDCt/la8ys7xDzWra1D3+fdodBS7ZQDf1
WnV55bNrkyuzFWDODLVa8a3IeV1t94q8l3OGhbnJt3U1TQjVRDUFZYORKH7kPo/vm6A2tua+d33j
KKQKOK+33+Ec7pD77tXELMFS+QZjE2m9rR9s6WtTIpfEKhfKWswkrpj22LjX5wuLU/bc53lKj+aY
Vaa3V78EsAx+n7NwWTbXS9DDOIwOki8Xh2c3IN5yhEjszpHlTfN6Kjw9HoipqZJdG9yLVCcYCntq
zh0tPi5GMM0wmCKDKPPlf8o1HUmu4BPAfiKs70QPY99xfZFcQLWGDTE7IusGwg9Yx4oOvXaUwPrI
TJjej0YQn5NtOTrNDOeT6Ct2d3g1e2RI/aXuPzR7SKFOAvSgCdIYUEiVjTHpRbKr7ySsTdAc4Qrk
PeX80vJKHNZLjraqJFOEhOroz3ZIXJwaPbzjYoMX2463QFGBGP7CutdPF1n7kdGnQUeAdtcYEnmx
6dktA3dq6QoTrpUStJOyGiniXsWbzobdSNA83tcvc+pMY4XL1SCNc/iFNWB7ZjGUud2vfvGMEBoY
Wtf12p9TfrFt6+O1eCXH5QL8SH02ujjIOTZE+Slx677MXFxdmaUoKZGvFIYwXHYOkFdP2IbKcI4y
GURsXPxPmnna4cv0YGh7xNptg+CURlTONk2KQrbmStM1wMQDpUTi9LqGKLzaarMlWm1X8Rfo70fv
mgfOqbKRqIIqgGU+Hspy3fhoJkS7QqGq9bYONJit6VsvOBjyMdTBZRJ2BnHdpD3622IsiRsuRtoJ
ckHLHAfuEIMLhYVZ1++YIWOx6Dol6Z8R/IIYbKXYtAmTUWcLILKEW6A8B29QKeTzqInKIZHedYex
1Qz5qIBUxxcFsdc5V4ZzF1H5tZhUcHPFtxWl8NbgfLBkr4NFpX48qna4n0RCYXyK5A5ffo/ivCyM
nOLGQsSmO2JHTAnNjBlsYnqmw/oq6xdcjP6mFzsONKQBHkgcx0egXJTRtPsmedTVUBLG4cEVQPoW
Hg8r9FJ3F4UnHIaijJtswY+ZGb3w8eMUjmGsYKrGmKzJA7b2VKdf3lRBRMn3nntfdR+8BtpM0K+d
6YAKrURWwdRszkecDN9MZrV3TUoK9KhXG1PsEfhj+GLVTgQtU1Mur7rQDWdk10lS9lu4GFKhG3Mq
xI8h0JPeGTxmgTdCJ9jUlRZN2raffhBuwvYhXEuEmODH8se0Ut1CPPxqcwwxCzrI1HC4KIJl+/xb
mEuNWBCZcA1Fwx8oCTuyvNRfe0Hm5YbmrRrOwnrfA0aR3TY2GvnzacYRXapgQB0Ige8r1eIOVgjT
clr3lkWbAI2D2WfMgPeL+7QMq1rMYFyJ4QiMCCHJXBQ8LohRJOXdljTKuj0g9e2/gKItBZ5bug0B
WVBUQa/DdxC8vjsm2WnBK/qDwQe9bca3JIvQl3Vicnz5iCO9byJVkcmO+YfVX5Ib/fQKALHNkWGQ
u5Qx5LmyyCRNK8DJSQqVQJRAWQMVKwqVpH5/elEBgE/3rj6/9ERTW3oV3evihJBv/UKwbiCJkR1M
FFI2RATiPfR3OLuowvq4QrfWqx2MCFTnpLP9yvaANfpVz0Z3B9YnqzW+uEGXk+8aJhtOVJNwjcL0
MLWH7myp+8MIBncmOovHyMk7+Hnb8ODaxyyGetfU4VnqTxDbfPER/TkPlqgZRY3xQEMue5ikl188
lPhEEijKRhSJu/D9Ci8QWIBjpmOQDQROtwEtnd99xuMgLejCHoQIDTM+R+lbNNO9k6s6MMONXO3X
vrucDTdJISLRFe2ZSK0U4tDBkqPDiwG9omPrKYJT3fZt+jr5sTRgugXF6RFmZRKn2tseWY0ZWxzs
Txxn6LMTgAuOcWnAbMca4y86DuMdjDzG1/wZylvyN+rRsoys8APwDGFfT7I9EmEdfSeIktEqU6mg
scXM2yWA2stlDuJ0bgCQWtBugVCOYuTbQoyvWkHNF8ymEd2v8LVHoX5Ywa4ThNN+Af3AEAD5PPO4
UQ7FWchDve9xaK8+ILfxeUBZ5xWukrL2rnu0hWPyoVv0Alv0wiG2bkF4kKTzikdNTZG7DVYM8wOb
67TDIBpQ1qJo76PkCujpIUcGhH2IE6NYqerVjOXTIfFla7Krq6MpBTE2s4DIqKrzlHvG4vtdLZcp
yDZhKo4lBgZZFbn36fPyHjHP505JZ6SGAXXD7j3q89keY0nfe2VOxGgkSQ+2k7EWTWScq7Eo8nUh
61PG+NPfbC9gCvX/jWdMGOV83RhOCWxcmzHWwmfZvW640Zt35RhoI/VdCOYdZcxdL+WbwkyOuSOC
g+/RME1wtZGVTSckxmXFraJHoeXgNVr2L4+rVAZAbqRduVRdrYJBLwdzDY2sloacbGDAWmfM7Ix8
/szu5SGcFuzhS3SflpwdRiZOJomtkBm/RaiGdF13oSjI2qGOs5IsUSg+NdAww6Xb2oxKAEs/qBFm
bonKpq8X7ntNJSGTKmT0/+c3a/5aNa4IRnOCshm2GoeIzBOY6Lk3xvRO1a/GTs8qsbpY7vuKjYV7
tO/Kdp3dcEXQY7+HNkLYmQaCNXiDwI6jIWTbE9/+7K5a2aG9aDxlPwf/HVIHeG2Kb+rV0gnPmTO7
Fc8cPgDx5OebwdESSne95LLuQM0D0XvoP0fkgpA5//KxYi0DEfPfGz9mObulKmCVMxoVAT6HOsV2
20/MNfdjWdfgZ6PhdeVKWovi9DoZQRVAI7QTL8A9K+ZGZELxDSBpNaOjm8c4ujEPRLVzWBqSM3tF
558rtWxLP80MAr/E5Ly+RwGG/tvhw1pWeXjO6uhvX7rNO9QHVs51aV2FUuIUZ5bs27cZfRKV7xHn
xwFn8ClnAhKEv8Ajm+PaQprmkWP9sKCZiqbDNLq/N9Cs0ACj7tWySJ1QT+CAvuzq6clPPUqJooVB
iDxp4dMGQPx/IKVihu1307ckXmNFqLrUHD8VEbtyGM549hB4p2zC5xjw0jv+t8u7pW006QExYV4H
Iln3ii3RwsdbScEY5EX4czii7se/dETV5azunEW9uWVGSGUfGlRBFLTFqJqMF18s5WaSoyEpZB+S
fi0ymaEy06LdH0J8cj/wj4UGBkpvosndfTYodrGXWLutrK4TdA/M+wcAWqS044xdcIAg1UAm3Dz+
5W9OK5l4J0CJPaiHWkBm8xw0U7rL1L1E/w5GOuet5769rez0GlhhcVw0QSzk/fBmXvCEBE31aSqa
GYdactpamSjFpJ3dIQFIu7oZJhGbXujJHx4VnE2WEosPebSacCz9nanixVkXUe67z5C4w8BNdez5
9EIhjfaCyCmbKI1/9ZbrQzRgcGIXC/krGGItsqBWbJIUAyNIf3sM6qgzpj55oDLzZ3jCYp5+hwgM
Lagzf7MoNHmqYyPcOwBNBKS8PYI/sHKVdvG4TnrivesdLXYtGqrbWGTi4JB7KX4tlyQKFM5GsAcC
oz+VyLMAhp5J4ettwJhfIo7owmBEtq1HTpexAd0qwWmdA0yuUiM0nl0I8Y22jtDsY1HLGVIuWp7u
WqFl7YFnbQVZ1JuIRFq6BdXr6aSLqn/mdIqeEQF3neVCrC4BxFybGbP8XflnngvSfJJ37j6EJDQV
YWhKT7Dx31bWI3L1b98LUW7twYdMWIfCImUmtJcaFaXYDl81ljDdr23ZyYF48lCKCdRvzlvUWgUW
jHVerpNo3gWiMYMNkAGb7VhOq/4Y2j2TYMxHlA1lc0+MBNAjAUTDyZghXhsCTp+eDqSmifkhib2x
3h/cOhHFr34eijCeBmuxBucILvLuSsRi8bMXO1OYBu9HfmAqHbSiO1VsMKD/MvH+e3wMiBbUZXt3
iMxeCoih9Wb0KpMX6RRr4VWoQwlU7mwb2EkT2OLt9KlQOydCFXK+2Dh96CmYu89QUzGcG+d520cv
wIV48prHLnDkRwSDBLt0T1Uc2YNHQmsKWz+27ixwe3RvngjoJxAGHl2slTxEoMSiw/W1AhJQl8XE
i6kuApXN51XD+b3c99dtTaMf8CaEsneM2Ww1+dfLqip/LBgCJmqWA5x3FIl7dZYIJR29Kdp5Kv8P
GJpdTJYdXU/x1jwt6w09zHrZf6+aUCJrZM2GYTSptdiTUH8yLczSN/MO27CGWEqeMYTPi+XQxJmx
s53RIMbjtJOVTrZnxsycKrEvgHo6kqACfbDzJ9A+zkLhjIwFVjZR4hhVB1G0Vv9LKySr0jDj0cyg
Otwp8tuhaZuWnRDz6IyRpWdHGMUCESQjnY6dKWfXA80Qfio72m5toIraqRey7kv1qGq/C3k77Mi0
CWzfx4uOjaqY4eugASoom98YmuOgNDuxdyP0XxMCLeEn6BH0hiHQOVftwsGyG0z8nHPFt4t+JJ3T
24jYfu7a/Bt9FSO02VZ35+yKCmC5adUe9nQdeMkXdMNwdNj4uRGgpfJ83Jk/2fF/lT9Gk7/5SrrR
HRHNeXDSOwUggEgMqXzycrI+ISHBRZdC1VS98q/sHbbOG7Vthu3eOMV4tnNWO+1+nqwMCVA8limW
JHlEOUvi8wOV7o2ELfh5gzotqOL6EgKIwUWzV3GrN+mhSOaIs/XfEP7hlgEoAwDQdxhGHvhQaPE6
HZ06nhjbGEXgv3YdOunOThn5H9ZAfxT7mucSLr04HsUv73b+EUqCO1+HUX6r7ckn70yt8zcGZMEz
DRNtzZtoabm2YrsVmrcU+cMMlVryFTLQJGi6fnUiq52+Pz4Vjk2biOHdGyOlYelINvuGbraaV0Bp
WddP/Tvzjbvbu5LlUJI5LrsvlK1UIbys0RmQtSIEF682Eak3n1u6pc2x5qQCZNJUVV8cf9Ba7PRD
DbyhteIe+MzAAcLkE8caQ1JLvUe+EVf51fjGOP+I2vG34UPkBRJ182tgDDCtRCOsVx+gh3n4i0Dv
H9pkihz2SGVS/SeBKV5AW19NkxiIfn4ra4B5AtJ17nHnN/k578ip2KXgGkyzd1iITuGhXxtuNauU
r8cWXixqCcakQrPJqIACNdQi0h1UNkTAH++fVxUnpmASyMd3S5gXWHwrrnOoD7efJO/ftXcUPIGN
T2bZ6SZ7okknEVK/zGVsA2tdr015CN1c6tUZEBxf8XB9Jyq8V3HoTCidqqr22j+KTKHxLRG4MNag
tR+GzDpg54l1+ApgYiDvX1eiOhWfesuJkgtw2Rvu1QvZoGBb9xPYcFsd1rRbSF++f0oIYlOWBQyN
qJAUtwrKSN8YoSjvQOmB1IbWk+UK1QihSK8hueDaaFxANZDxU4keT1XyDceFzehkkNMiCLFybN/v
AXNvnui4XYqSSFLMZBDOqatockszgRIYZLjBZug+13U3CyLwHelFcyHCLyD+EaG12POHQoVG9AoX
JNAZXS6JaGv3GEwPtLFESA9BC1bWN1Of9GJMBWJHIGD053RHvN9r6AXxbwzTlIDa8RikAYTTCGRm
rVbeqRHGb8+WUVwxImVqeLnQVkIAOYv9kpU+8xs0auEYU4fCjCNwvmZ1hhf+wz/dmF6bYvgzl+Hq
Qw0sFXwmYNaLBkavUWhI5KdXF/KnDm1FwRznRSjkweMFzsMErQ1J/XF3K6qV0MFQgeCsF5zHpCl2
PMreNjxETVDYlAA83tfFLWl/9nL1AGZdcks5Y8xCnmDk3vYyoe6DTF3bPpYx+yYYM8ceIv140kOT
BRXsuGUfy+XRBmho58oibT4eBTKfEHYbE10lAURcWYcoUh92eeL3moOxqQHpvmqIpwkfBMmMdHsU
4xcK3U+LMJF5ekDaSrpqnE+JyOshmqEgVCa6YdLoOsYxLJTme4iHpWNUuejHLqAGeF5uhwvhV2uT
JGkTCYwExZgE3AOZzDHHJ3B/bvelUMJT749/Pzql4PMp08M0zHQe2uEC4t1LegY4WV6N5oSTP4y4
4mkTLtdh9lSizbLKCsKFtn8eSgw88kAL0+H+W1s9c3OznJrj9+aSCmT6O5/96uD3PmgjAhnaZ3uZ
K3LSTbgYFNqViw7TGm2OLwwWoN8dLU+VG5UwYbyU2bDsbtTico1Y6RkidzrEbQXNzPCXP65391o/
ooWb9D+ObvmEoGDIfa4StCy8OOuQBbXUeYx4E3wAp0l3uRLSLmJH8I/uNHDtcpImfeoMg3UeYG4p
51TXvQQbAk32Lx9p5RDZ8MHsKDI6oDezRL5ID4AukBaOdyEupSlk/Z0t1vdL/mYARBTe3AQ8+yYV
YLqRuvyVoK7lYri3qHM88Dsuzq7X56FaaXHHeU7ohKl4Ce6pe/2mBJ7xvanksWzIJSy/lSKr5+oy
KOqadr33tNRAtKC1twaPqGur+KqfPNrLlyrAW6MlC7SWXAjPsRVPs/L7qndYhaMvH5Cv72ePsE5k
B7M+GqwnqNcohmHYtOIYF9QXvUws2ixBaaBjALKDFKoTAosuFVWrsI1iRnyEqRinXzIR7Bams5TK
qgN5/8ZXzUfxlVYJV75LiNY2iME4vUSYA/JafcavrZT8Pkw5mwfzl9rTnBxXB4OhoRDasPXxNmJF
k04OqhZ5cpSBH7OTrABfOLoCPwZEr37j04bLhcG39WleAELej7XWBDSALpco6nyvP+Ftg21nGnE6
g8Jn4jz58QWsLPa0n5lYDYPApdQ1vHG/vWbK7nXwVpw/qrRgWN7I4kZTHMbtQibTllzzyR3FR4fF
Kkh6ogRCXIGUURL9sUjNZRB7KNSTjGWvQsQ8hoZrWHACpYgeBe8CIf1D23KA6poF7FoNXYV8gnl1
SLEgejdThHDeqNsjLzlu61fG33hEQOMJex0tc+f2HFDniZ7FRlz5IEAFf4ESSpnJ6td39sJnzC1R
n6rkB0dvUExorabiUNdSeQEkcmQi3ChtkWro24B5JlTJw4/OwrhlA++PZh1ayO8eLqyvnNzs8IJL
fnM07955nK0mlE6Y+W0A/2VoOMoLYsbp40/loGmAlVs39NoIAtRL8H19w9T/P9YIdo180Jk9Y4yi
pzhWhRnJ4oq4+JcEoqdPZ0lHTYZjb9fx0o0DfKGW/2Kb7nw9TBdq70As01ATv6ZQiCWbRmUmmFgK
MLIRESDNJTUW4r8jXVTJzCMDEEmjoeXm/2pBR1dO8icSHLhYOheA01KCjVkM14vpUXDBO8RecHVX
+cvtnOi4SFn9TNSxgYFBjT1+jDeJIQtRBdOH9cwHYgSxFKlINZDSUZGmC/H6oLvTJ/c+Dyw5GxSc
Z2BHUD/oAbfHh0wJeK88gJobFLFZCEwnHr7LjIBc59Cg8FVED7DVN/kdrLPkPC6pz2Kem9ZFPcfM
cEcWXV+sAuH3BX1xZRTGb3mxq8RY7AjI8JKBuzX2xtbCvAwCXek6eBVdGEyhDsRX5ovplDRghr37
AHLoI4mYEVnS+sSAN9EnkD/5Fz68Wztq7weQAn90vi6/LbjA5kNfGK0f7r6QAYPe3fz4s7vVCBDp
bWb725YHAdMyu/dq+zniAcqnNuCaD8gdE9sW4H2TOrFXl2QadcyTArn1wNoPErRIVxaEu8mJPGC3
R3mDstXiROZZ7KIwbDXG0IKZxS9bYTc7mJBpQN0lu/LtdmETAXe8yQ8RO1DxI8H08czns3e85bMO
YkncL5z9Ke6dE7GeaIlJ2OpPvM37SfqetRAPwSQQ3shL5xWFerSr7O3e396oDrVCe7Wyz6ETMso/
PeK6zcYLTp+DEHeZ+s/wuxODQeYza4GyI693mBBmLMuhenQylxvB0NXf23jJgqzfSez0eQBNMoSh
MmW7U2E79tvAI7Y5mcX5mjxtCRDy2PoAKEBcwsi8q1In9QzxdsNOVfqxOUZ2/PMjx09SCBy4bE87
6Bk66JgtzFFGhSOx0tXfdYVVMg7MbZwcdIFSPEcKpbM/f+jkka6cIDbyWEO5D9RR9QxfXCdFFa4w
lIdd4PKBcV9/2J9ONKnl/6THnvXrN6xeu2NYYtT/rOt8rg8xU26WTuI7rw75Lmb/ZUj6Fe3Cq2K1
46c3XhC3iNjqqswBSQK54vyseJzt/5oTNkYirF4Z44foDys5u/peDLOlCPMtJvPgMuxRhZ/Yb5eQ
upGVfGCNL21yjD7dUzBas6rCHhHUidXEzZnKwy4v7Bp8/ZagpzOPlOPnZTncfDV4HOy4IORO637M
XInILN8KADEouSoG5Ja//+CLYcvktX+144k+EC1yBKcUvjOnOAsqjoojYwmN1zdMO2eSBE+ZcWKw
iP4NdM8rMy8nvfgZFWQ+HGHM9DYupz40+f5VnTKw/FiNDZtb+GjW/3w05v8Tk5vAoCHsz6k/oLI1
wKCAiKfKNBvCurkGgqapjSRtWrGw1xDtSab67JcGgyz4HT9IoCB4B9wI9ojL+JFINll90qd2iMZp
Wv3/CUDNAwQWBcr+gs2iQKxIMuU60eN7QhlpgOcC/0iPFvcSJsuW5cYrXHLHugYrPQxa9ByO7UJ1
Hp3yapW7C8PCKa3CPgn72s93M0UjZjT61zsAt+H2J7RXmL99i7xszW134ptDXwsZkWh/90fpUt0P
5lt4zYtXY7DertPZEU+CIMwhn7Dr7/coKsgnr/sk7x5UhH3KCjkTSvCB3sdd7bW+jcvuk/gxg+AH
lxrZCGl3M5A3kFNnyjH/wpxYGbjxFLmiOuhq3oeJTb2JuSRA3KFNb/z0nyCY8Wvy4GKo7Y88vi9u
7uf36y6PH96mOyUCvfVzFU21IfR9aEdqAlZgD7Sal+9zNy8NHkxytL82J3TsWOpkzl7R7j8psYaL
K82DaUvDdOGQ/T2UDUAWTbPfAnBF7uxWKHBWjN8pKiLtKKyUrkEtz0dvszcyFns9OePO/6ScfnbM
Dp56ifhJ5f3aHVFfqKfSHzOY6AMQYYgZqKeGwL0kbaw11V3zzz72NZEkJdjGDgqsrnN41UHvLB4p
uL6o9YOXojkDKI+XkYpVz/HXip1c9+aJ1CTLDX6S7RCgdo+AHPVAEDfYnhPGfT8BcAAhDPvW/Q7i
eui6sFEKp76UhfluAOi7Lk3uP/jlIDeFNk7ZJEUEoiEdMm+PZhfpI2ciIEcgZBp4GAU7flTmIXlr
gYiBGL6Zuc+IXHmFvxubZ7ac9vZGnmAdhi0mKhkbzlrqE1VaiyDhy61hR75njS7e2rP90qN90+TH
7/Wz7L4CFSaMUPcOK1T4HUrxwC8LfpxrqqGyW/gTHnKxO45O8/vxdd/mw0b8kSrxr5wM/MIELBfw
3lFvfw0OkDDsMzABWD5mAtGWv9cUZwFonkODoldp52kztddvUW+Se+RC0s+Io3/mV+0bpC7jJYSF
5EwjGwMp3qI9kwBmy1qrniFP8ifX4zJxibiWAnGq/JVeONoLON3T9EKKeo8icNerL+Dm3W1ZXDVT
kbsgWKijA6YhtaKrGOvimsKM0Sxsu4cDESCuyu16maN/QBmCDKy/4s84N/FuOsmmxq0cMZ9x1XOY
OHvk06zCxln33EG9qFzrzKitz5zwxg7NHEnZJjJVW8obDqSogWa/D4Lnl+xgi2rASrjaUR+QZy/B
EKJ9mnSSlWFTXZdebbwnHTv7L4/QEvv9s15XKKajP5YXwTAjklS7BCLFqjwwzc6O9QYwJ1R+tRp9
icgakWZGmlq6kSmMXvoIXol6H710sudZsA8P6JuE/bKsW5wM+97TQkbEe3flytBDJfNFWVSBZoS0
Chv2pT24igEPaBwqPq1K86oh8RQZYWPU8oYQ6jvxjHU1RB/O6QqTPpK0xHqH914P5nWWpr/bCGAn
OvXHpzwS+zdQbEavTPGcuxE6DER9cwWvFvJWnHz+awIMDNW/uQiy/PK2DFAn7yNKkRBQhWutDVGK
Ead6egjEa4db9gxlhdOC/i8Rz70bqBGXeNxmxc2yCtmMyuYLJMH1aIuG9D2L6moqBpm158X0fAZi
RfGx4Uk7yA+TAF+QqrfnM8B6HrEA9YMOP5zepdrRQAZQNN2QHJpPi6/pZee+/n0hwTrp8jk++Z32
KiJW5+EcJLpquVh0cihdzAWZcy5AdNDr0n9Ojj6WcRmgGpNiLeIJnKi0ZzFSppbrEXrxFAnmOigV
js5IvYM4llRqJIR7ZC9aMcbJ4INQctvy8OZEHNLxenb5xCe+uJ3VeiSIxTa5oxL+VYleKsn3p18I
TUe1GFVAau2vaT7EJ3V+8qA+J9qaHjdVEaVKG9aTCRwb2eagBVInCOX44yWdub6Cu04LoswxnBML
qg/QNa4if4CyVVtwuBMBybf9/7jgXEs1er3J+xBNTdcr7wsTj5TI6FSURPUSealnFOetF6oom/eU
6uQpMYcZYGZVBDCvTBjSPkoKisAD0eobYf94xyXtrajzftT4Ha8fuYH18Nw1/v0X5b3f/SlyGLzT
GQx6VoxySzls1mGJMSsCxi0mITd5mu5uV6WIEHVRkzir872c/ml46UxtcX5s+wnySi8YayYpG6ZW
3xIeulpgmIo2nSeEXM9OXbicPJxC0xAvsFOeWR0AUofXFwMht2uLm9l5fulGEtqm1AC+wO/Erzro
CPxXDigFg6/GPmFb/BChHAeayXUtumai4kGJi7fCirTb/TVgvAGIHfqsgb6Wgva9nrTJx+96FvOx
Kh3y0/t/5I9KuZs1HfHN8qEnG1XNA/kvHHOVqAsra5vSqiPjbO8e28Mx+ZD6twzmr0KB6Fm8Lt8B
b9AAqeXyx8W0qh5Uy7Fd/fRHMfQXA9QWEUZLd0tPOcJYwqTM1xiRLZ4OgC9J6yAa+9a63wkHCY5z
cijhaquwxKoKnN7dlgnN3TUwa46QAAVVa6avjEMp2gCsV8FM1of1/+g44PMuU+/wzz2TXZOsPAZ4
/rTOXj+d3lFIyNL5apd7yg88PBF+b5/8G7Xgz8Idwkt5EgmUIz1+EbybNlHPWNeekMe0xTHUCdMC
H0dSkdajlAGxx9b47/n3XChxLMA1shCHb+9LUo3VRQyLjqY+1x86j2oBeIQfQBDLWZZOFEXJxbCo
UyGo4du6roTm6DA/aPeBmnC85/RHlgOC/mwmahAtvT1x2BQm2IHfF8P9Nbk2R5Rkb8JUH7tVmvYh
h+pu00LVR56ZNc3AHxCDVknp0pHTzYgz4lLhTsVAt8FyU7x3qCGhqJpDec00V9bYG1R9kXucH6wZ
3im8PfMkHyvwYB+zqDDDP863JtLIhPr/D1OsfMSjJZFYUV4GmvOgAnhY0bVwnqAYsAsuLeYpEXWM
f9Di+9dnXgKRrVst0Qp0hYknQesAVNN4vSESbYW4s18ZNf9ddKtq1ZWOntdsBEtXDZPBC3Elqa52
WPbQeaLF53ZQRCbQyx9wa19I5HLoXiQAeFvudJwCtaqSU0+1hfPFJkiNrZ8UJo0VQYYRvVRUAFkT
qeJj2ozQIAbzvIlEmrGZj2WSUVHXrkBmHTnznlyKo+rLrVM7M8KMv1KAcg8nCxNJRoM5YK8Y4FYf
hgX565U2/k4CjejwzlhZUyTzHW9scfNklwaH7/XiJdJ4T+sBFu7/GuyFSWtqLKeUqVlh7vbZgcYT
ncNorzX+Dgq87hOHTkrkap/ftUWnC25jLAprTdwVLTzjNjGaie9hpuLFbfb1M9g+z5rnWkOebBuN
defgCM3eak1oHWvCfMdnELVF8cNZTlvE/ZV8Ub+dC6igy9Pn+eRiSYAZ951JCl2vNGJVIik3Rpc5
rjT3S7tlR7dH9qhxOiXojBcVqT74MYomQJU1SVaIOICBWhZo4dj4JM5v9wd9ycupJ/HTw5eSdWOT
yWSfBp/tybCDA0Nos9l4eQGGb+Dmj4RkF+r61SstCTN7JeBHTLsovIyVQblXXnhtE1RDHK0AWyNM
3+EcimVt+nLrlZsV6mLkNWUclgLrxzPUhQ3zkRknmWu55CXb8N6GYy6dEXJbvzV96hTXCT79+tO7
jv8PxtpmMIOA7azN85uis+watpnEjzWaXvIBBTUEMm89Hwb1t47jOA8IDIKyF3GgAcFTQvhNWSns
tsTfIqNXUenQwlaJuJ+WR68rkifYlDZwJOUpliA6KiOvA9rOr2Mhwia2UVmd/2K/0hJnbnNUnET/
VPnopCX5I5+bx7AQXzd2H8ZinxVeUsXXi2/SAzxvjNfKLmQU7bqqDm2EsP6zpmuvP4+jlAx6A5Ey
j0ETJTaRxHNuDn6luNzNPMN8B/h+D7lEC98MKPm8U018EEXYMXbnjPWCQwJLI7ToXkI/L6O/kdtT
wkArC26MgbOcbn4zm28E6oYzJCiFGfgwPhX7fdntpn8yTJtB1LxBJCjfKvGaWMIDXAfItbCG6ysL
z7TQ+zjJLdtfRobxyiqxkKYuiIoYwdggWcQG6DXGxQrkB9Z059cfBJ0/aV/AZCMLIzUfxORlkULl
0hL/WrNziFs3OBCYRoYHnfVekrWM4MjH5ew1ePf0WPdAtnYxJwiKQasz0c6tGb8X2RDVkCeeY65B
0XL8PeE1fbOSHWTTa90GmDunF62VI0CL6JhosvSb6Jwoq6ThlJ4AszXbc4Q/F3da5MVq4QX40nOq
/2MkluZL2gktrls5J/ZWpx5kSkPjX9Mrgkp83xQtOt1QHHBV3mCdxl1qe0bXZ45X8nbsLKSgWCzQ
3vnitLgeX9sfpHKOBY8WI9FWSaWRJe6VPNBVKPaMk2NteGYcxCGRxFR4QkRDjZV0FocJZLm1IibQ
CXDtCNyiFHP/PjX/WJBZlTW2c3FV3NGkbFfCdGEZQ3L8L9jxJ5qfBMfVuH7ckjtb3OZlVcAPcQk2
b4UFWATDDXRGjz+9cs+EXrsdqEMb1/II6+XyeLD06YcCINBMNxmTD9oM/AT87aiLixICTMrRa4oc
YRQQlzQaZquHOu9R5EjK5xsC2pDGFmUPV7ibd4HD9HrPw/cs7lScqj/vGODHFkbVw5QtJInxXUam
3x5R7xYMiz3pibpgh4biw9rWia4siNOtR5fPMRW6OqU/ff2hR/ZVFvJM/vqYlAFThyCFGOxKf9ub
phuOyUM+RVF42mMNEm9jX6PyyoircHc3KOPG6oRhhoQRj82j36s4UmKGNrSLStip57SkWrHYtrhK
u7C1wUwfHdgJrmtg5xBEmhfm97jP2tvXep8KG4hMC1B3i6kbf4T4zr551WEfC9YthddHGczCKzKi
MigeJsfCSgXOxHyGlH72ezdGoOdfJsY75AWau+jHdMxFMydJ0171XVTjHcwBYCWsY1UdKwOF+m7O
Fnw7XXKjpY5IU3Yd+b+mXEo+2Jk+BjPIhUPHDSB/LHMIbmLoklzkHv3ivh6dTzxYLWWBATwmyxto
kc7go5Tge2/LJZZ/JPBkl2QdWfXSFp9YZMexN7B8IUYESsOGQZPgzclM2ISpPqNT2F+uRyQOVFW2
WqqdYWLb8sxVswhFt2hZZJZ4rD8m9l2kMkPDiPihrfopoWF+SDKYA44pd686W7DysERb4umGEAJr
l/FSO9fUGpIDN7R4a313EKNtrH9t6lIpWiRsLEFaRNLgEr8ZFJ/cLZr8NS6MTowNAyD3RaL/n+wB
uyJhEr7QIovDM7VlwKijcgEd0pZIVHMHHso9d3u1Mn8ykv0CGDcAnxcixaCkGlsG7AEEmbXw3JEN
MJbwZzTafAOtVAnt52xIi0JHDchsb8a7QZkq2tfn0U0xsNp0P4GxS3IKjsrq6Klt71tANP2IVZs5
CfMEuv1JmjGppENrhAAio8f+GeRLWJOfFnkGp2f8nyO685ZVmA5hFDs1Hz4ZSEyPUAVVlC/SngF7
+dScr5HAcdM/JksP9rrnT07EZqq5veQZuq5VhqwLcnoM1gbgnfs1a6NIB2vTrPdHINheqgKGPx76
QjxTvGyibEhiq4PEjwl58tPT8wFSMP+XtZoDSPhS7g9pkZ4SXfXh2trmSehtJUowLYWwSUiY2oXr
InvL4Ek6h6ngyh/GkKXVP3Q6sRLpxDlyu/nJ2P4zSNPM4CXVXiUWB7+Dd8aa4ghDI+vutTv3nwzY
fFYVWksUsUa2k22YzALCLws2kbZ3/14BeVQKHWjTQcby+7A6iSv1skwqBN4xNlT7GIEHvIZSuIgi
NmehD5BpErSfejEdgedMjyFpuzSh+iBFVOLaRt47fExmbVD3pHq5BZlu1LXsIBdcxTkakhYiqnz5
NsxZ8jNpgSvwVDLT8AuhD77nn/ijHZKErjimBdHQIfyUymso4+RRN6V9Y5pWUPsNSx7ziEcncXwg
2l6j0BFXjX/RMd6abtIWzf1nEIjEHEd+RhVtdYlPlCn7hkgIsSDqdtazLfo8wwF4sKyNEjLYJM+q
mLlp2k0vi5xfaxxdmtHuBgsgAUGlB0Yty/16QNwJRuwFh8JFJoeJe6rhl4j8YtLTxsoBdx3eMUbz
WO9WH2/4j9Acq6RVQDJOaz5JdiH6ZDmAqzQ35pecJ3bDTTA9L8zlTqSqnvYkmyqjBRDQaISzxEsk
TkDrtiN8TcetUDPuR2AHvCbdWRDA8RldzknDaYSK7ICpjWiN3eexjatt0vfhImv1C4D2Vt6JLVeP
Uxz9K0hUCAWE6kv4mE8y3vlP+AO84zOO2mHdMRf4Em6fuqkl5k6oV8qMA5utiBLRsp9Q0dLxUctf
b3j77EMWelvctfhWA5vQqRvb9Gk47pGlsB/Y7MPqSxQEryr8hU1jO9KijKzP4h3oJIKLqTzPpi1x
Sjp0/dsaQwfS8W/CIWPlHFbXHgyKsu6SL3rd1fXWXuzKlzdf/cDKPkClVA01klGE8nRHr/l9TDhd
vNw54onLkezXv54lKLRFKR3DMVfOWYj7Fa91gWFPmxJ5EPWhTN73fGNwrCmHoZ9IsaDBz1DXGgIo
OVn2sgLE1EUL+Aglxus8IzpBMfXkXm9dKKhGLsS6djDjK/AkrqQCuXyIOBUrgMVmGILVVG1iwfje
f+UD+yfQon8kAJfoGpQ/Ap1Ya06BdN6P7EL1NGJUZXmQWmxkfbPM7lvPqvD9xUT/y+H0BXGsbkAi
Ol1l7SqemOz8pOgwfnOGfJn0rvR/nA2IU6GmGt1QioPVHg8gLTi3w0ZjlC2kundgy9Y3AGCfGA4z
cDuNwZeEgjPTPLFAOE5ZlECSQvB2pLClSfm9Idp02nRfd2WmwZhnXthfwGviVMwFoq/LMR5ay6iO
iR5fvNEY56Cv+OOZntlecrFCuwUIuffa9UX5Yx7fBIPwlkcrDSZNtUNom/XcBC8Wq7NUIOuOrZkF
H1t92Ol8oPkb7WyiS3m13lIZW7/5XkpeDZpvnS35VVsD1BKbyjZE5oel4Od8eOW/DR7wvF/2U55c
E08yQzBdtuVmkzsnPFxq1MP1N7AY+xVB8kNPlaeYJZDzj8so3Fg63Ztzz9uXGkOPcyp2cvZdJlQQ
ww5EdrMkhh4Ce20wCl5isRcvqrgdFwvKaLe6OxH09SBBR/oq5DZFzYwFpI1m9LbBzV+I1A3nhqm1
ct/XMsX/Zom1FDFh4aV5LGsa9Tl3DVkJWCnpvotVPnt0HR3PDBbRl77ZLfPverde1cAEEET6GiPU
58ve8gxDMoWjojOsY+QnFre70FZ76jMy0eYwQlAzfsBkN/K5YP/2oRWxFFTReaDjbzo0CwEi1CfF
qI2IRL49/Xn5g0FLqhWT17hpfU2X1BHjv0lHuljCWTivPsE0dxNERTqBTmijCSRfKqG3EwPn/eVa
2We3373N06igUQITqqyitp9fvqtFGTfoYvPskOMTDglv3ZQEDL4pbwTotPmoBSR0bc3ehXvJuDWF
BnuRMUHc5XhI5V413fKX/H0U3XRKMvI7vIm65/0i01juNFKLG14l7dMvNnICBmn50X8oRs17Dl/s
Q1NWw51kdPNGF5gpnruwS6OQGxdeis1a4lFq85FYKaotCPeET85ljlOX6gRO8+uzohGCvspv3fXh
ssvn0Mu4CVW4R+I7qO4yzXqpORwaaZplV/aMalrN8s8gaxKWot1f4ewGlwXJLvIV6otDwPuhqm1U
0gCUeib5P6Yt1GVeacGBzQGrA2TUPaDJT9y9bsqBj3aspCRLRdsKAga0mueXKe3Msk86Ae3KZZBy
dMbn8uaUvqUcMuTaz3K+/fBjec8L9wtQLpeq+Rl57mmE/bxr4jxMJ4uAOv+nmt2c/mxyvc/DhkQ3
JpnL4hQkmvquiD+xW9H9r3miSOW+XJlV4vsYBdRz8vcRhJwsNwyag+jipaZ1xp494zdpLi5XnaWg
YWYGzFWX+4t8Yv0rY1nE5zfi3j2gRoKygo4RdH8g74J1+x1xtF2u9DvAdftg31cbHOQH+ixxy2es
MA2SyOZXPIIl0WG22E07eqnXXoMlQe8ifrr6tigV7Q8rmjhbZv9dys5W22OWnuzUFFLgYwqMW6Fh
SakHc1VpbpNFYhCSPM/mqfGNzDPiSu1U2GaQmmRALyiaxAHU3iINj5jvDdANrWyOid1DUVvgwEaJ
etLeznP7bhaRHYizFqmg9RxAEKIF20THIYfdo5Rt5hsponncNtK8U2YkGPWpXUX/lyfMEIoLl/nE
g+51J9tVeu83XRTrTxXoQ0WdnWPjKZculvWU87dT/zAgeI5TQt7b5QWp6nngU/MQ/WDkKz2DnVw2
WiwGfgDn86uphUM7Lu8Y1JchugrHxlUL/LV/+c8FEy6pBxDAAJNqOvkJVcoQ0iNjW5ogoiSobI6A
OLUnOoIUzJxhfcfL2aV4T3iZemuGbi5KYyxLUZ/bR13xcg1UvyRGePqc1waJlenBl1S0hl5r/u1X
125PvQUDEslV7TT+R7+a0k30yK5B6e959+cLww1Plsg9dRG/zCuv/yfIkbAJOjtTVKjix8AVbwIy
cgXTfiTgy+IA04rIiMQZY1P+pcNk8ITQk0GExU32QwkxShvm6hqU1lsQRNhQMbX/mQm2YHQuIAxN
TTETmw0v/JzFvQ/QGV9+8hg+BCO3gJF0JjBiBUgkcttNYksB/8yWrU8kkOYllQmJGZz8nfvu2UlC
UY/Ww3PgPNeVvpf+D3yFZq2SzcZaeQpZt2q34WpMEb89055sF8JfytJ0QWKoWbMQpbsFeBca/Wsc
ossDlME9j5SKnvr9Ta2WS80+oEV9f25/EqlKpDe3xqu0z038ql/A3cvg1LoRw2II/t/h6snw4N1+
kExeTvl27o//BPXxktWIb8a9GY9JJNnM/Bxto3VciNP2MTjc1YPLoKb8zc1woKalSCxLX1oH5iqC
3wtf+84yRd/id1z4Jh6wKlgPzpBHbHZYI0QWWOHno2pgqfrxdS9UJeBUFvOxEWGPDAHESSVQF+ym
3S81AtkdY4Y6XfflsylH91NBGsHZyCe5fgwG4FHwO6RWzRAKyxHHCs8H3ESSLrRJbNNY+PQxbI4B
hMZ1M7dxrEt2w5P/U4jUQI7ENdT0uP3RUj0fNKFmhvaBHqCAhS4LFLoSWfYlI3nDCu4r30MtSTsj
wjq11GFUSCzzqe3AI73AnfDQXEay2bD0xA/zDK9zoz/+6y9oC4FmTZlSCVMBiI9brK4xfp9Li59l
h2J1m0XonGIX+Qnf6vIHk44ktIZbh9IB1Z9mS7EyvdLyfdir69wo2vyGxhACGIw0dDLKLg5o6hKX
DHjC3ttoyn8NtBx56cGysr2LW2ySptCTFJAdKwZXH8ga1n9lLov01frOHNiE85DA9Uoq0i7598wI
mEk2OksJ02e+cb1hvQ8FWbj5yJFbRvE6790Y51QZ3WtBaKlzNtN030AeDO9F45GO1yrQmYkWlwTx
gM5Zi9bQN9qvCQKOz93F7u9PRpkz14tijPeCWp+KNjXTKBhSRWKxa6jg1HZMcKOMtJsOFB+VjAk7
rX2UhlWl95p5vzjYnkPsqBkeERVSy8mVdoAdbOyznOxn2uO4MZtJtJVn9LyoSpVgwD9UGmQfd33o
pssGb9IqO8OOPgz6o1Ys3m3p4ug2+TPRRJhZYjEKi4dXZotts5y/vN51+7RAbUuF+zNvfuV4Lif+
c5eKbJTE3KhmJA0e907jav3C5sFtLbv3FHckuKSUsLDa0RMOGT7kx3limOJd9/Fpy9mj33iXlI7h
n43e/W9KfCp0mlSfTZPpE0hlZMn024iLTGJHfDCyOpRuCgc2yFTnxScNedtSeA6fwJtuz4W2rTOT
CHkyDOLvTEyRLNKfM83nOcFFlisGbamOo9tVVVqjSVPfS3/LQ37zzxCGWr82MPwEOjCM69BQqRGD
aCACjV69T2hleyvbgGx6bzQxdpeiLNE/pp3BR0PNgU8RJOXd4ksJ7Yn/tX5ydTaGLFchX4Ymos89
vcKXoY6aCDYEDlv3O/o0nuorv402NhygKBWNl+8kSUVxOjrgIpHcOsq48Mj9PztD8X0QSGIfE3kj
7PgheRMxu9NWcu/6oHKtOtiAv9lhbTWYiX4EeucVaBW0X+y/tXTy6o98pAN37PV0VbFhJUwy1gQR
mNPSek3cyPjMb2EZq3xaSy5oft/4IwGlNDqDanZb5HJ7Jh1gN9dbKaoWq5NctaNWdE4WQjI09ip0
LqTtbR7p69Kx/EqqYJFBrONgkHaA5pCPMgNvnrdX2WdFmnqUmQadNWy1RUoZh8v4MFqD6+MLdL2T
tdCGypRhp9ntLKffo30kFYrsAiaAjVTcBPKGnWdJLi4ULePg1ibeng8X5B3q/L9z/G28cJTOExWl
/tyF6/VuyaBjHfiWX3apkUIGxO9Du3AboQQk8gaIqCdAVWPe0ewwjSZYEtMFot9nFfIApUneN+j3
VQ2pBxXh48UFSS2it7RBJoOSnSG9KGCyoKga80kc/wyjK2oi+cFjg0UsPTWh4WrfyQYIz3Bd2/Ud
W8phx2kmfm4qPjBzZOQgUyvCeN2fWcuU6W2iLD0/cv8nCdWZJ7VD7ZbsE/O32Crp3SSsh+/SntqR
UfuPrBlySNm+V47NiMcsDT8BOTmoMMp+69uh1BrUmsdyvuHmlUDgQipCkieMNjRwRmaqj5SMegB3
Mec895FOeI2cXvb5gGt+JHGJDyN7SQ17UtIkNRPvQxwfn73SngDvhYQKrgMGnrwm2h/loabdnH8X
KMBLycJckllZbamrJ+3fv8899Si1d5ry2/UzyZ/lwOXDR+mUKQ3wfZiOT9JgekSUS2TkBt9s1zUA
2xSBJHiSczZxxuXXl/upu4+d3So/Y/nXsUWH/PMvx5/xU2CV/HCjQ5QBLSVI8V/+ExpOR5ccHiR8
VrpZDInReGsC4mCJ9upygwNaRApmhgwLekczY+KNoxpLP8PkSoQZ35kklvPZ/dsfoD85THp2ayS2
mjhL2b8nxyriRRkuNt45nZAjMFJXkN4j7XbFh3i/Zp+BISB686JCp6bxrGFtKPSDn+nsMIwQH+MO
jt3BaYS4iBKGPOtIfkqt9JjG+JMM2sxlps+dQff1vqBvijVQ42y+WFGifvf278Koksj76HBXlrSi
d7GTn3EwYZbTMc5c6/F6XHYo6ZSnQ4ANFQFdR3BmRbOFagNFJzJts9w6JiSaTG7PALB7QKRcVtTp
Fv/0us3jIQ8FAi2YtKhHcPY2cdUhUBDZVxwsPC1BRZy8D4OoXrRuR8jaNKJ+VHI+pQShZP+8GWKZ
y49AyhJVrReB74xR1RHwPvNtSVeUYaeKCsgCeDDuvnwVGclap51Zj4mr4H8zNU5Z0qru7J7s5dfX
UAzwnq61t8XvSpEvdbXjUDFL2YwzefkJub59HtS4DgtV5p0hLejq0FxCnCgiqGFgUSS42uJVLYQR
kKiEquf3c7yjCMz1sILbgdS3oM4KudJSfju1hPGZBoOkBaWqNP9szhBebsYmeeuP6Wn7GI2Bgduz
mFSdOUdq5Illp56j23V3zyGDa4xCt3BRubsl+0K+WrwxH+PR4iwOdtXt+3RJ5qSU0FYLq2F6ND+m
qjf0z5HHyGQfEb/gc7w/iI1CwEyL0bUICxbGRmWkE5hxZzGhF2vow7YS6o7VLDIFZGXW/w3pKS0X
5VyDIYhI9CS7crQ1G5cSk4AtYAqWvJSbCcmXEnUyVc2edmQJYNJonNQWt/QN4zY9/rWTfVHmD/rD
0HFKmLfEfJvx2xMY/LmsXqtGbhg3yVov0M4z/LIE98Asyot/H1wo9ngT62LJ63PKTu8rl1lnr8CO
kUtb0tL7ZcuV8QDk7jeVrkNSX4xvYddBZvLUROJEgLd4SVmGtGtAOeGtPIDH14y6OSwUGaJYuwtN
f6MANBEu5wmGgMKCbuwHP73chAKaYtfBbjqoFWAInP7eCy4ryWF0TvwBV3E2uWOYh5u2bQbdX+0T
eDyEJdP72m1jIQMSm//Bb0wXTqBE3kTB12KqOtJ51rl3ADsUS+m6b5KVgKFOwI3FLDGKsAp6UDuy
gmN2U3zlA4HG9O3+l8Yecdtfxtbwasd340/47KH0UdtH40KsU7DvfUeNaOp3lTesmpTz7eomBmnB
XHoNMjHL+J+NiEB5D41pvEmcTXu5YHccvJcfEMuNfw+Z+TUwNNZXP07/HlG8hfZ5GzTAr8ipJnGT
/Lik5o+Rh2zMQTM3O7hSo21i+2Q19ZOVO8oQjyT7AbAWMVULJlZTKABACtav04HIkJomzklEH0O2
qN0U4rchw969ZKcOOO+uWGCNtvGdJUqsRmv+5VGDQlSSPU11Q8gTP95rMucdIRGaaAwto+vXvicd
nrNHKFL0Uwvdw2ea6BnhInFX8z5mR8hnaR0XMLOjL0GLAS+LTPrrboCJ6A7tW/8z1Xv1SiR5EVCu
MGTPLPt8nubLiKXP+V5bUtU+LI1N651W3QgK5Nqoc2g/QujKwrlNZNJKOeQO7rq+lQtprdDl0Vrs
wI+3JuZ0VCbKe/hhYi9G3Z5yGeYcMaJxQyBLN4GucardEnlweB260LjjJL3ZzpG/9Gsxvl5e0OV5
U+XOHeXd04oEcuSx/eX8npTfwXqXOJmKeG/O94GPu2CPSBTlejm/Kcd83XfvvuRjINCakZtarfaW
3DcWepRDj6eU3APUdPhNn0hemM+us9iht9Qio7Go4CVMI17cz71cjWC+YGhF8lYPPO624TIWHG1n
1NeOe2HDC9aovWXT1M26kO+1KHYJTtSZ8yunwsmeA+1hyATEpfUs0HlaJcqWrniG3+tGIYTLSXoc
l7BWZ3tscEcOQ64ZSeo4duPpiG5BPaTW0IBuwtWxYg4cS0SqAHeDpt3u/k9Mnq1FgmY8r1xqhFdi
Zb6kQE2HRbOii6sJQD9fZp4Q8IiyFVkOeH3phYUuTJlREJtBcAEPlvwOE/i09BFwoVSrRpgw/x2A
AhBN3jQ+REYPuVrROPrLlH2jTSWx+J+K+vkfBZwgJg4HX6lKTQw7gfLH/2zVMSqZ97B44jcccRQl
l3iG5PET0LGpTmgyONWDeSWxZypTH7kXeMqv0ySf4vH3AqIbzq+TOv6asyAvE13vSyyl1s4NR+kU
KDwr1uyaBmk7YFHocBxAZmbxOej2IO4Y/7LdX8qCNyQuoQIaEo1g/7VZbPlNxaAOSnJKRk4bLn8X
xtwXqQ+VUQLzj6EsiJPTEg2I+KheRAJM8yqIHObjGPt1mAegPvjsCIm3QRD2RYJ4fSsdtFB3ggDE
T/Jz0gjexsc8kx9CD59dOR9HqYKBGLwTBfRYBemStN/6JjBusvuTjam3SyDf/kcfy64GVVah6d+M
1kkG7MqV3WPZeMQeH4cP0+Y3ZRjskwVNz4Nb4XCLM41TRovQLUm896rTIb5hNeeto7eHX0Ewqy49
TnxwUWbWW864uES+nBZ+fnVOIOKTQPuf8TL0M+Cfdd2022rPQuRaWi7f9TUpaNo6DtYsB+Xmnx/g
oxsqK7SDAa0DOT6xmin74k0nX1JJGyQMPM5TQ7dGKGHuviWpA7C8Zrn9W63uk98sueV58P1CgETl
ZnvViOuaBiq10cLj1EGdyedv3HNuSEPeVZe6U7xWNYAgn8h5WEdp6njHU3rbbJI9fr+p2UtZYsDb
V8gkFiOf6YPjHDEJ67F2frcO7eCUSf1ZuJCH4cAzOKSBFo09EOJ977urD1hvU1mUeqitqdcNOCeT
Z73hhIw7M9XU+kvpC7ZeKRcSzmsQVl/uTsh4tTJxSu492ZqF93N73doqtbuMlmyC0iTAStWJKLzy
JpPS0Zl0tgEydK5hby2v057ScSkI/rTichgIe3lCxWPAAZyXI2m/9r5uWBWI7tsGvJKo+eLiRyXs
3WcQlxatAH39/4EU1jg4UV6jxQT03tjU96G84TSGlVSKUFCZ1UNF64UWp56VlEwR2Kk5dNEWQtFe
Zhatx1ZKhe/deBZ8TjHn0rrSKi6JwMwJ2fRgRKOsupRC+PE/NJlx9ZFFTKFelxmewdni5OF/5dML
gjeLImAB6ZoTSkw9cdAqxOEhEbm1QIBN7/81VaGAycUEcOmsnnqafgo19k28CTGj1sHS/+H0jQA2
41fIAlnfAQ5f42e4F8RNdl+AXLfkTW/O44EuJAvVg3YgAFFzleZCCpaNDs50pLDocSx6az3fAKdk
852TDCla3udWaTHwLc7GC5nKJqVJg+4BG3+VT18kPN6AynWWORsnjYEiXCBlOe860wx6poKbBPS1
Lss/rduKicTC678CUUTdTyInO2B6GEaTCcDUmIy24zGuddPz0OMrhlMtHmYt5tZ9Mk8jv4X5Du1v
2pSexwUB0Cp01q9oT+ewo5xW2OLNJI/FeV3+t/7EduFXwJdjgcuvDOlT2A/beW1+DoQft8SxyWeW
TMvD+2Mm6w2on3XML/uLAoFqLSMqQ9XVsPVau1r841AoIH+SZDe1HhP0JFTTvun+3nIOh+fX8AxE
fwJ0vGjkj77Et+5ExiZ+O4uYsUQ1pXt4yLfp8cAXxKLrghx8KAkoOjBU6FtYuaz2uhEKw+jZm6il
Nb2Far5ClUC/cHuuXC9PD6qF2Wvpxj24cdZ1bvTL5lF0MO3e+5g2Gbs8IBSbjQH25R99DzJQ/fRk
Vr7lBzn86tD/XEIvAJSHgHnhx1tjksLCwKy5zpNy5kt3cFhPkzOLJ2JSLu13Z5LM6/3r8zFV2cRx
jwPFSX3RR+gZ7GpwpMi0dk0h28ltD8t7VRoapXYBrYMgn3WxBMtBBHpIsefhGhow1/sPE+1Qvh/d
bfL01hTpNmiE9JRiIGS87IbuQOVpaG0wPM9ltnQB7suU+2QFxhnwvlbjNw5sGeX9Sr6Llh0aBcmr
rhI8tvmgQycs+pQFIIoNY9jeAJc5uouersc/bROlWkxW9DH33hPbpNZyVrMFGACgodSw2FUSek7/
UVVjmt+FfK1dI/et1ARihmB/FA1lBbFLdpR0rC9ZM4JLNqh43Yr6fj4VXrrke710qAsJawG5qdlU
qS+kj6KmlKb/vPF08Mn51uZt6U8yL6iYv8RQJGYj/Cq9c0WJyncPqG1hd+Cu1EGs31rdQpFCxcST
Vubieodwu2YORt8C1c0SehiIPqgr6okGYbRMbvT7LfRf44W6D4+33FlXD4flvft3h9eD6u3s4Zfk
D4j1M+RbPUX0OOkxEx6MUQI1HD7ey1nDWHPZNWopueM2nE0P/hYd6bYSiQtwiAnnE7yG4yBnZTuH
JCZxomvqGcxzHOrtAfkp9b2nFtb0DUMF8VjoqFisLx3/ioKzg2nVPr7aVf/v3AvDSqyDCPlr8gKl
jdyGKoFgcxIT3EVcru9acopwroSacs8l7xJScmoYDkbXLYsvvWbiRD1Y7zSGs/xPaodHkhS1pywZ
NVuz7cYtFOzZIsRkcfXSUj8AiGAzpWWrn8jbzThg+L0MuAAK8oK5G0o+GKbPPd3MRup0713/puqI
uMrD9PVutSQUt7EQ1M5af8RNGAz95SudfwzMpq1rw9g/qdayifJZeiZ8OnQGL807jOT+4eK4y9bX
QO2oUkabd4MWl/FeTaYiUxAvw9GVHKWXw6m9rXeV/LHolrqRZxbc9naUfova4QH5C3dwqlJiiu5x
3HdGlztzg4HFMfAYb3tixa4ay5uODUsbwz0OqUxdJC4eO4C3TzbKdT/HalEnp/76tV6TE5a2lVvq
L4ciHmYHnAOBV/ZIYYV72tDkiRLYIzn2ZLTlE0skP7vP/SDPL/nKtD2HjaM9KrGDAcYQAVLhktY8
u1XGooAt3sBU93GcZLR5nU3qkfNa5fZkp7BaITMz9pU+lNz/21pBLGEE0lrJL0HpWIsT7iKU1nr0
V6L5XeCpyYE+sILe6B00bv4P3slWPZ3c88DQ8GOqxJmaicNwQ/5iVAhtp4bD+oEPWK34nEcFfzsD
NOKPQqX7Iy57vTkpEcn5pDmsMvLDTX8On136W9gvFjHCF1kU6S3pvnquHpZQWRBWGL8Br6Q6KBfX
VKVd3wBiGwCcZSR9H1XdzS8RuHGrkgJsupbWOiZ54JFApeRx80Z+jtab7lipdjcUE6uZMFASbcqq
Sl6kS0bpF/qxTbns8nzFs8u76npIA++Ux6i1O0fViOxfa12iTVIErQBxVbhXRKymt8D2fTzL0MIo
6a6dHnxfpJ+oRU9chmQOcio4dgAAh8C9Ra4Na3WY49oPDnhocYbkPVx4IJiLnXEdOMUBYJANLjve
JkPla76jA4LQ21aztlopexwVFIMOnwk6wy2AD3FSf7O+4wiHaF9wimDv2jIMypIPDD8hW8E4BVrP
Tneo1qYDrTUzduEOub37tJ8WUBOykgW31YDYAhqFTe1+iw/Ud4JOqTmRUObR8pt2571KBTkqN7xs
eoyaPbYvxrEDhxhWAi2kNcS4MIC+5EVTDB2nEDmty3aw3/gXoSZWl1uYoarhPY23C/4GuaqB4FVw
ZHgJglOeV52DCHq83Wx5ZK1IkVExM/Q/vFYKo4w2Igzx7Dkgxb4VW+jmfqlo2CdGfsW6mUR9vwBh
S21Jo7InZDRwJRDEzBu2/dIeJPss2qsRpq1MPn7AzKFFBpQhPrgnrLB2oZpmrOFQQw5D3tfxhGaC
HpCreAxYkFluJrDitgon7CrMNl0VoOZDB8J7XGThyZMLGtOJWtWPyxVwS9DaeGs+46zJKV0TNR3Y
I7WRNZIffHvpw+M6aNA+I1TZ7/EdCaPeSIh3rCTmqikZAX0mgVrOvQNGp+qOT9Or1QNGh2JbNyWZ
9TW6xFZCcwxD7FLUguS0yFCquXHMlTd6LoxlQ9FKf6JUxYiMReJyx0Hbm84lfXbSiuUeYaPvYYeb
Lfcq45d+JSkyvqIIE9WyDacuxPUFxTBjyBqcixq8Ps9Kn+TClgyUIiGrMquYZefd6rJ2cu/L1SHc
dS+R2rHJwBIPP2Qqq5PJxDzYvtrrX/zuTuEXCdoCHfYdnSA9q8ig8YC7DHXyWn3jnFj4rpNSgVO2
QGFyjNKXiEe9dh8T+j0sRYEq/oGP5ERosgMfI5fx3WXadQ+df2O/Tgj2K+AoC5bQAzyPPDB9PcKe
maQ0zYjemwecam9/BvQI/0+WN44I2LxgQXPu9mpQ0La3fyerQU3303KhFB/59YQhvlj0/kk8FF+g
RCUArjabEvt/RUC4X6FE1PPQrdtrDCgQs6Qqd4dgpRn1viEgO/WrlyCcT+/z7gGkmSpTR+X9Upvp
Hrir9G9KHa6GMhM41a1GmJVhOfhVV2FiqSQZlX/20SyVscPs2awlP0bK2c/8rVVlPgYYBVEW3HZ2
Psa2W3R78zr0Xvdm2RJPplJMx4RpQDS6f2os6usfXObtXjozvKK2HMWdZ97S2zAv2VIpjCExg6SP
c6Qv8MG6cgMBroOeoWEzrqViVTo852AxH5iE1Por+GuziI7jzGeIjzW/QbM4e6b0+FJ3tve6W7Zk
zSfkIvc26cEjipy+hn3DJOE4dDnT69M8fnzuQUsu06dsqYsEuX0Uckpw7Zn2DqdjlqNVsxKehXOO
pW6v2+8wVfF590tBIlN/ZqbzsIOso/ukSUeSRubz4seMAjVAgdSKcGMZPYoZDDBTlFCMO+emOJEL
rZPwr//QrApzCIZq3PzDWEjQ5UjBCB3SIQ55V3uzzCDxm8M4gLq2NvC3qcMSm9NwTpDA8X0prV5w
EERg/Hij3NgvSkb1yWOBG2IvUiRor7W46PUJ23w/of/CjAqPVgJd/3Z/9C68GPwMsmvnoxfqaCVJ
NGw/qfEwznyQiVqLqX2G0aKXx0R09qNWRLj4JVlwEImWra2ea2VLQ/b8fvc0LmjfFfFqe2BRv3pt
UbfU9YLb5Km9udNJPqdL+FI20prKlz0VazrzWDEa53qe0CXg9UKCWyPGcGdB2vpTTl+NEV+jSAKV
hZn9zkfxzUxJ06xk/0JTNljFCqBrjlDuGEKuNPN7lAudgOmiiLOdTEqMIr8ZI0ipSGcEgMfpgSOr
2811S9O245Kp2dtD4fS9sKtLFtL2YdtQqPiub+L/Zae/r0wPHnRIK7w3QcIRMsG8rsvvXDyJDllT
Jd7kiwpxD7B6GyQ5LuSPhoGgS8cIDEttmOIoHM9ebz2kgKjWOAGeBglqEB+xt/RSwR5CFFq/zz1s
1Cz79X5cSaXk75siBteoBSntOOWEeKFniM4wKaZBD1bxfDO2VkIt3UjjKjHDTL6LyzEqw9NqtvTF
VmsBTxqIF8Iep81mR2KYjIxD/eb4nQzlIXESf5tc1SBUw8WiZ3aUcsKjvpnw+TZInB0qYYjdStSm
DMqC+CiYNjykZUThGrFRcraL28vSMm5BOusBbJxTOw8eEjTh1W61/uc/Fu/BfhldTsxMWRwMTMVk
oQ+ElWDYCCTOJrolL+IvS4LslFJFw4aRz0d2SqFQl+NrIMpmN/FBDvDgVzQQm5XaLCaDeEQaRfuv
ogvMHH6D2/g3FmeRXE9D4FeuJK4xotrrYN/+jr2jWBoWKLToPx5A7OgT/qJ2YxDDQCEzt/qGzx6t
LMtkahtbzmQX5T+nJJUH63a/K24b5ua3/fdGJfk9Xn2Qb6SWi3h9ozhp5RtfnqyOZCtlX5VLxZMc
AA3RiCpx1IeqoAVqkOg3LS5fZDRcIf4iCN/thop7x071uHZk/hsIJhKl10er1gUh00obW+o8WB/y
A+fvmUse186JvAKoT+OdZQGZshKscYpTDfHlh1hgANjqFB0YdPf73TMdR+rJSION/4sIrXaU3kud
ELC0lKtypRPjQ9G8LUovVIxc7EkrGccMyAru+8wwgYeafcROsYbULvHIKB6Bb+S4Hoh7vyOaV7pR
5AvkL0IHaq+dbkPfKxCLqEM+qocYR5zlHGwH4sW8SxWSg25PgpxpwMruEQMBimapzDQX222l7ZVt
Qj7KaSB0UInwCsAgEarqA3Cj0GsP/aCFNIxqLgQHYorN5NPtq1R0Kk8umBcNPEwdiQT2+bmXo6mK
4OWEtwE/u0q7QEI7ecYYPa5bzcTfncU6vLCQyhJILQLcdsPzOs9r4T/pY32ObTzAV9SN85+1Koxb
DVB1gWA3IqdFo+Vg+GZ7MEqB1WEQv6EGzlF+mmsS4iTQOq+lnTPdRk7sEOZiQL3IxbdE9psqe+FE
iam4gF1YUAhQboBz1oKHiaomXVUCt0SQCF0CEuRyTZJlrt4q6DdfZNLcH/6+m7g6iWXNJKzgFJp7
DLMjBoaTNq90Fp3pzk+e0UlCq1g9khQ2YWEL4rk/dkZB7MjbpFBp2bUWKTZYRgDy2nV6+8xX1CqL
17bt0d2ipJRc/0zou8Tq5E+BFE4C5xcIMLp6Jy+iWilpeY6DqTup50dDSU3LqMKxXtYVzyeKOoV1
jvilvoHCswKrjoyUxb1qyeWalmH1k86o123KertPhxzE/iclUmSOT/aaBiLgqHyFDNA/OXGe1lbs
aEXKEuzxRY2f3H2gkCw2RUvrvSkTDFzvxfKUikh3/3nvNH2aa9e4jV0JohVP/AQ5m51ckLHp704M
h1l1uDEtkt4w4tfOKNJFI0Qi0kyxZ98UBsgSl/H3yH4lb5swrYJ05tT3DjazSc42oY13pgfGFS+e
cZHNsjIQ947IzPvhIYZ2ruURRgjDV1MgEYb6t8cz8Czqqh8AF2NxBZXdW5cJLP2r37kzGIZra5I+
mSpOuZA0/Hs+C6ZsDlbwdsVVSbBhRSqDJUkdGmKeCWxAilUeG74cA2hZOKet/eKWLYbChYTidgQk
/JSd9pBe9Wu+kcQlvug045bmzqj04m4zcUV5mkuDc75DYgwva/YyA6L7QWsmLOTGurJPOWabudi1
x/WsqRSdc2zhDp+AqHo1q4VHGMiRMHlQtohAMZCReRyMTJFxhh/EcFfY3dVNqmTl7QR8LxSyxFag
8j9MQTU5Gpv0trc9Y9Wv1FBhO5pVf3yLcg/e3/Ci5isVt5gomK9wSG02r5Ebvty5nDpx9LT11Zgp
5utI2wMNo4xCdo0IjNfjh7tkbswokjqhjSC9QDR3BV5cTcouOJsHoblsw6StSOMCF1EYodREV8e3
vQG4vQeUI6QOwnPXi+dPPLu1CY6oBa5kK0ghEoIDs4cSI93rknwhepi2gHz/CTNFWv+KrA742Wxs
TI9h/uHRCtb/cU//zF+uX+S1WiXIOFIiHxhW7Hy85uCMTmIlrZ23wQl9KUHgsmdYpdrJVgfC/bL3
3e9huVE3KcvxSwEbawhl3Ov4FAZfTRn3wDPPsB7O82fVfq/avquiRSFOKNARAxl70iRILWb6H0AQ
ot9MjRcnwHyoI7Fs/8wynaPmlFFFlwko1je2Ed5kJA3DXo3rYH+HZKvfow/0OHT6lsNXQepc+uYe
CPWUtNd/J+NTO+t9o9R97PEe61K8AT0wTIVxGLOfFbX4CSvjEcnjZRXH5hXfuAdc95isbmJUBs8O
zVhRgS+rrfRz0Od3LufGOA0TGYCcv9aqnZsBq16djwX4AQO+v6Q4KaiAVM+n3xoQMrduc93CfE6T
chzUuLwLc4jwgBV5MMt6TFK8ANgXrzotmgl8FpTaJFck1vy0YkA3Sj4F6XFa0cI16Xv2V98o8ltn
jPLO4+w6OqG06BG17omeaSgr+DHDR99frnJdv/kmZoPwyH+XProApsmDWcYCoHgNdJUBVWPLWuOn
PZR/b8KP+uVpRRtPGj4hKAn1YYd9LbyyJDtvz+/MUdw6Bp3fNUHWPBo/CNQn8UzgSgY1v4EJ9ee/
6U8DJu4cPqlkGIq6zQuM7LGMnuN2+UNk4DvkDRp0Egp3K/HEK+LBcw5phOSwpVcH+RczcVNRaWqF
rQeC0BR+oZyEFbMi/+SPI0tK8TPoxJEKke3ik8VkkjCTAvGV7mcju75zoILDGYlmUvGLECovKR69
QcNqxXQNmkykwKuSCg2vKDS4775nxVOi86DpkpO9veZ2b5IHFlix4JP9dIbJIVSH/55ms89aAs1c
9rTPZQd/GT727V3p+Ul/UgeQYNhH+WOx1HxXU9FvrRoA7chV+lTOAFWOh4aTReNJjZsJfX8PzYNX
GGNlku0kPXcsas9nCEIqZP6ZxflQgisQXvKDrW4iByXYhxAYS4WQ52rSNvy692vaLkIpEoICtYX0
WHF5raVKNRu57IWPH3sXsxsFkrQ+k0VpTyge3ZPWQQ+nx3/FP4yTCoyJSJR+YdGUEVCZD/t1b6le
dhEdl//9ohOCKct98g73PzJiPF65IgCe46dKpEJDQrr3yOWrVzWZcnziWdNsan3fLn1BCmrXPBAC
EOm92zD+KWrugcUQLJGLDy781ScpHn2gxW+qvEvN+qWjNwf69HpmX5v/L6vRNi+quEIuFo1UzDo6
hmaYnF7D6+qnIt4L4RJGAsa6iwzn+3OI80IYXOoAcB4MotJ9qRy74YeErJgm1rMC7kcxJ321x6Fq
FdJsihDQ1/Cxj9vCjd/ouUFcW7pg/+B212Ei1HNLK1+Ht9bRTuVaYRvWIMLUd+oaULtHitRTMkVH
9ZFm4bkkdWHoK3elaMjNlFe6dT1I5TwABDzB+mu5InInBj9pU25ZUPqHSL2Ze2Bt6xJhLeaWgjMq
7v9gKpW917fFGGuExcWa4e0G4R3itcvlnpAKVHfkHXNYYW/A1mREF2L87CUbC6MJmmwAX7/RADc9
jwCjvAJMWdWzsukztSvQruVbV33ypg9ElzAMJq9V1I5TG32eqTmfPsmvjnn0iU5OEq8L8ELSHW+9
wuTT9ukR3sI1PK1xPv8CC/xJZS6Fhf2L1oTne2ofxD2kb4xJrC8wXObUv+9BcPuBK8mGJXmcLJaa
JkGQFLS3pe+AzG5AZK21KRuHvivot3S+fF0WXjeu9lBYR+S7bm018E2w35YGoVqCqo59KDhrCUi5
ucWC+paPbxeJOZLv1MJbgGlaeiEXhnCyV0bG+LiwrTeIhPfMoy29/eRaaRj/fnYeh7OV9BTcljOr
/l1PmlEjcmXEuFWucFO4J83+SfRX2HVfjOW0B5F/iV1LacknGhXW1fel6lVCKjc0nIpsTWDZ44tX
jXmknnUYEG8PCpb3FeH2i05txMXdqWJp71waVJ/vHnXJpkmTwNQg1b8Rau9XXmZQuJqNQG2U5xwu
xoLwr8/RMzj2pa5wAsXCvpRXHH9RfZCFVUjSGA0tHQdwSnwoW83NmO7IBF9OKqu7WUUMOKPgDZdx
NKm/faoag23nJmYFH2ufTuDmaIOFUoI9EZ0JQc0xyI1yQrAydWoeXTf2g5fdwDi+dcsG3H6HNL8f
+RX/SXb6tNK5ov3rrKEprraPAMvvzWM4XnBxw42wViqi3pZso8QevAqMotH/qGAzp6izp6Rrlxc1
xmCM5B7tHINj6oU4Qmohr6qMv62sFilGmI3+Ol8W2FVkWQr9F+rZ+fmqtELpaU+JvqjzKLS23UIY
AL8U/1ufJRDqaaeAplkxe0FhMFxVb4YcdT2sVtKpYG3CEY/9WWgP8CXgBYNdfNoADawFMH+9vcjh
kV0Kuntz6LJHdCeI6wpSIoV7ti20t5aG81rE/hy2oScwK0uN2G2/DPN+zcgi+OmaAtn5FhzTGck0
cDH6eFxzptWXocX4dFPCtpn3HH7A0C28eIcq27DMLCuILqoXBHESiHZv4gNfXtDBFyHrHBD7aU5c
XNQkq1y32s8t3nxCJ3gNcmt4Stis39JzajA+w2NvS6jdggijf5RpBUZdQBJ5vS8TI1+jj6L2zuB5
1yHut460yuNCEnGwNbcQYeZO2rkDpDnffiulaICt5uPrHUJMyhQffY7PZCmZhrUAHN5CRukWIT2G
iPzwILBjHYS0B3+GTUeHL04gbHxtjB3wlqSvgedq++HWGmNueR/uP23dlOC0R4BZcA0udImcerVF
Ef/yDPFMqjupxFd3/OfjUyYdK8GHoVuni1+JDxCAsQT1/xjv1RldQZNN6ha2WKNnAf/MxHMc3Hyo
XROUDwkS6JteNze7LkJNUtAHu6AE0yztR7Psr0eepN7YKEtkMn4FM8ceWYaVIuuYv8qQMMfu+6uY
6nfMgiVp6ScyUBGboI8I7H3gEcVvxW4/UCZHCroAv3RHd0CjO7uPvf890P/7QIMRTEM8R7i/HRvo
uAkiaKqOfQ6CT+sdUXM+4NhIUZAULLQ9txq5ItWlK0LllotTm5KgafDyIZVB0s13+xKMYlss92MV
LqsidPTo2xpBKsWQt1PryapEAMJiqv3ntwhu5EtPGaJSOl/VtPgVNH0M2TEjyvdrEJ7OasLWRma5
wHLlC+39mgMFkGJYyqWSw5AkKJ0HYPlwY4Qwi1jSkMqd7LyoySH8QkCvu7PO7Y9u2shwzYbrtoDM
Rx/MdrXJbp2tg0gwMtdJCBSW4l//RsglR+Z6XYhhh8pbtjGFZgFlcCn6t4aR5S4qWZOsqGYwczhB
CB4XVIISVgbvTD6UHNDJC30b+Nl8vibG23+Sk6RiWFVciPicilHHRIUQGeyhaWvSE5ldpY0K2nJU
S716IQ1MzmTM3Bmag/77gv7+2nP1aTpNp/h4REVSBnuIgkfSfpuAiAmqzup6FPbS/bH+IxBTMSum
4HgNidSP/X7dntnxiHvD84gWmAaEwTieaJ6BWLR2Sa9L7tu3965YRx05dMDpIyLl2kZ7BUvp7UG1
7fZ24cWH575rzLgF8AxX7vX5zsCILd1u74cY9q+HsJns9KugQyr1JqpoK7H0b2Q358mrI261DFBE
2hz8B4f5/ZZ1JZX4kN5XotckfkiiHbiL5z1m6kLBPjSMN1+4aHzym9XOJvWLxq+7wjCLCaSnbj/W
skIQoNo8i7Txuv0ZrdqNcOTyZZcCIkJ6ZwqCsHQinmNiHQv1WKLy1guD5BelGBoAYrdE6OjmwUxf
DA7HVqBRWDz/Xkfav5GHDsugb1LYdqqFxCmhIO8Nt3++w64/YGOx1pcgz+ZEwihwNo476ff0Q5Kc
A04IacVzC0qKgLsk7ffcXQAR+b4VdAbVpvb4fIZxE28Da6xkKOWt2kQcWl43XayHm8GIy0Sh6gyg
Kz8R2xHJtpB0L8T/X81Svi0lR/jnKGVQ9Cg62++faeJroa/oakqcPRSgFG+vZiyr9/EQDr4c/kOl
FWU8DRFSIaDYCMbvVyZhylj+skmYikOEKcYABKYjx6T5H3l5bNZ61eIMr2qjju5be9I5R8dFerT3
/tgchmHM7osH3D6MWSAnT8uVgIcPocT4a/hGMrtlOGYLDSXHCnVd9yviwHI6Qoscg5c1mYsaOuQ2
WzwhdG6cfzEJU52ojIWe3+9XU15NpFmLItdSRatz5uAsuoNbFAJhaRcZaGRSjXbQTw/YC7Q3dwGH
R/ibc1JkYWnF4G3DrDAAsW3P52Mpigo9A4x3vJ+5xYV1KXPewQKnEsLNkSPYNoZPRoCinXJk7SMP
YoKOG8Wcr/o5subytt/vJsvsAQXMjVzqlRLFbNG+Xhp1sNJo6C4SVVCijI00/3C7Zs7akHswxdfl
ppOjlwdjKx7r377dbvRLxRwvYgpMFbMZfgpUz+TI6nfJe9arleA6R012CZ1mGtSByrdwzJMQHsOc
uGgQOPw4OxxHUjQqXKwBaFZSp90QXyfpCojht8SQW+djN4+mj1WwD+bTXpln505ZzlLQ4rjtVJ2j
Tj1VgSxjPK5R+OsVHnLFEwXZ+TiAm6PeuFF0J/PIu8Oe3RQBOqRAZZcodf5ujT3Z4wyG49xtv+Tc
gLyA+ZSZqWbvoxT06vL1bX6liuIIvYFvoQGsJnerAiQeiiPHnpF2qmZLk8uRyA5xjuS5o1WOOwFC
ykuK+ek/DDADAO5OPei3XzSUMF6V81tsSwRUE30vhXj2h3zWhZtk1dEYdG9zLObkQfyWi6x84cI3
eK7FntMRyFgpUfgjRASQLMaDVa4YXikTrDtTPsfUkCrdkrVDuyaX1qKRAWIIJNONvUu7B9VHvP/S
RbacfC1HL4v/5OADi2dECjooLSlnPqsukQgrJmNmH0cSlIRNAbzh4kuC/i3fH2Ne73vucuTFtR/p
AJLH2BaDcuUEYWu7wV7x2niEdpqWADHORJ+iJ3bCEaXSbs3MqOSaj8BbNoTYd5QwKVeSuLqt1tcV
ebr8NfFyzxzo/Fvolt+2XthRsEqJleU3ZlrjEPJdIAsWTo55t8Rg1K+g/GbfetnesIoJVdDoXgj/
2o1/sBGVK/C9hszNRpmvOW2mPC4ANP+ZGUm2Dolrf6/MsDoHC7jTgk4N1ZR+eAnlB0qu0OKc7to1
m9lVxbmYXLvSYZ+qAAkMus9WAO+xrB1h2TR/UzmnD7mtxaMxr0yHiVdybFjWSRGpeFRdzguAb+ZI
esfBlrjiSJ/kWxLTpUzBCoTZdOWX8cUqcrWNwJiV4IE0t05tBMxSPHhxn+cmWkg/LSCUZcJFFikG
uDw/s2yqzOVcpAJboN84w7/NN5nMxrPn7PkNupkzEDujZKyyyHNGCBa7AtZylN/sNMX43JbdgerO
WfZoLnmEeOQKPAUaFgiAQkSACiN8mFwQDy9Io2cfmhU9oH3XhOh22UTOkeJU54ErrDvutDgA0Cdj
HCm54R81v/XWneqLroDs4UpHbkqmMa87mmASxI7EJi1MTenJEqGwM3sEp73RmW6UtV6LQf07m7oW
gFKLS8Hr7L3bg+Njqu1GbvwHqUTB9UkjQ0Kk68CqumEBUL+AL8sUUZUiAnLpPCNN2tgpMPDgg9ju
ZCh14CQiBBMthXyUbzcZJz3cAXwEm4ZiDEQHYRsp/vsZG8kgoU1NZ1ZjnVuq36XA4U1IoxOBQelg
GpHKwkvg2qdYK+nz59qpihHvN4ExaU17kofXDiRoojk3d1/YBjS934chjXl+1o/KkKw/Rbr2Iu5x
D3+5+yXAW0vOCfQXaCqgR6uOh7JJF+SWfHClczvMQnQAMqRcLqZpY4Ak62vL4c1ouYjLHgeZzDg1
QM05fLBS0Hi0bmHF1wykCvlRmdzy3EO/HVUe+hM7HaY4xLmgofCNX9KoWj3C/3Wnrho5pcJuNUGp
sq3Y4PvrVhFFc0A/NJ1n8Cv2C5UsDA0AeLFhV5hehmejc/kak1J0tX3xqu5fOVyIOCQj5t72p+HS
8ClIUt1KmRgjVZtQE+FF6JGMsbz6EI4//2F33xH7ig+Rk+rVJtoefcRDbtKxV/XqKLkbvM3uqO8l
Vb+iqXalkqa+H8gfy38byfDlEqLVEbU+YfLU/2Izm4VAkloxx7bvr+khFcvLxyJ7OWe4yMQspbUu
3xL5PHBE2mSYqPUdwX5sTZBCplbj+YHKlKrnu6tgEixQHQM0bwt1agl92GV00kySEEC8h9BWr/Ij
dDYjJZ2pNdBIS1ipVZa0Hnj71aG8g7z7Z3vgkyQJrVLxybcAZaO6ok34PLUASIXnrWqzbwYQ5gOB
WohKczFZAHjP6AAL7HkgEn4D4FKYjPtBtjLXFGf2iMRYw0SgS18Kcl+s/GYIVBvxNe7EZAUonVgf
l4rkV6GL7Skasdfilpbg3B68NNIOnxAdvE2mW4TgRAUj6oVx4ZEp4nwhT9KZI1+DzRJI9mxWd2pT
xkePuPEoLVsU1dxL7BLSReA2Jx6SBJdcvuwMDAGfHbm3ujT7bZuc4FfdlGjin/UVoPgq3UzVi37b
i3GNd4zwx08SX4eQkLK82nFYg4x+Mqv9ViYW5dMmST1+7zQhl+W2zyFT3dUUmXT0VHjHZG2xh5Tz
VtTeInyZVVN+lonIaPRzTDMJ7suB15x6M3at5y5WZx3AEnTAho1GMwVTXAh7ehmfPvV5LLuNJguY
1Fq50JP78H8pL+0MZTD3l0sLCQG6EJwV7aT6KKClveAhPJkp7jKjoHVT1FOLh0mIa6RtrjLrr1pj
ME+J5vdInT4+5rKGBbnsQ5X3k7KffFR9AiQ+/64P05puJ4w23lGyhUpjH+6x4VLPAc8WHyBHAU8T
XzcqTH31IsevQlDxmWg0mhOn6Z2EU97rI7q6yzHBQ5bwfa/V20b0S+WNgZYciM9rskVsk9Oy9Y6r
bu3FpCujihk7FTpJf8kDRKTuXOcl7Y4zDUfIpWVOkHdpSnRiu2GFY0mZi9IUEO9S6R01et1TRLDN
VnFPvQAxquC2tukXEUTxduUXF4DVOFlIuqfV+dCBHA/VOMKnGZCUMBTPp3d13y7rOP8V7kWyBjnC
sSk1XThVCjtOamlimhGfjLxk5IZNKLWikNgbodi7IOTfeDJTm17uSerW/F1sCxPsoUDQmEw//pYt
8/dCWVuCNc0AXAkBw/jQnms2n6mlbCcIpwYSUz+K0TQeYWhvVmbXgaX9zrLkRCZ8eNSROgwZ6aPA
m8N6bq5BIkOmf+jBhG+xHADokRxtNBJFdL9JCWM8nQSQ6T7ZqqZzAZco2fCiCnl7V9QZ25lcQapS
Ubwn85OE2uhHxuBWyiSL10xQCweUzEFDEl5aeilR0xuF4wikq8w9q4D9qelq4CHM21YeazMM3W/w
a/8VVgk5VB0JAcJHLmiLWmIq42T7yIRFtrz2D3RxL94GNTCPsh3MKFjxjctHZgeFhj40oCeWSP9N
ELezfBGuDtECfDfid965DW+wss3E1CVnRIVqKYm3Qpa3WUx6dCBp3d/zLtBE56Oxg+RodhksEdg/
JAvQigAf3Wgl3pap2FnFKmNrlgH3efLBFtykZXDrg2uYm+rDpIpxUxQ/6RRoNmwucvQ74b/+2EoN
bZpYaO1hDJuHEea0RLRLRntP0LTRe71h2fAcGLV6FQ2qrvw5ArzMmQoKQbwb07qrqfQpWcvdlfXs
vChFMC/8BjTC9twaC5LpbOJq17Jd/L1d7IQ91ZDL9nMo/50MLd9IDaeEWmUgK3lMcRB/8y7K1kF9
yVoL52EvoT1NjX8XKIBy/BT/P2alzkIuibjhIugseZUqU4A5HRcwvnMMP+ypJzstaoJ5EtDV5CKd
bPoJWGEwGyiaJazdr+dNxoNdLBny7IOYR3OLRgIy8KGN4PpPEcZ1vuXc6vmCGUdL0du9HuupsG1Q
mQMLVI5kGYVyISNJCLA21PUIqfyC+lE260JmKmMGYPINyMHCdYCHTzhUaZZq9RgLWVS49bTWMxUr
kQlwa/zlTs3H/c5Y9alz6nFwASPBL0oc3Z+9DoSIOXx9kNWRQC9lnHdJlHl9Hejhhp5DzU/AzND0
V11D1ZY48ViQEDWoZG8Z7vDq+8PraHKYgFAWh33g+xLeExdBtYy/LGRUo6PBnmmqTL5DBq6Z+iRf
jtOouXKQBv7KFBIhzFWE6OnyX+EjnQ7MGGRifR+F2LFpK+sNU4ppwpweMBsfLwJcrzO2oc83Y1gF
ZsJU30UYi4/PTsrDryUbzFnZ0Apx5FG6GV2Mrj4Q9DZKXnnIPIVcXEa19nr/kLa7Bmj73lbWYEVE
v6qRLeoCHz8EXvktS5oU/eXGc6q4nvcMaewvuNZIgSllFie0/r0HrPbwYfrDWOIArjHxFoCp5mJi
AwPDaY+tPVCGaheY8cGb32nPSjzhix3gI92qhhaFdsTZ35Wv61MihbveOAUi37NucpovQ+mWRbTE
JjZ1PBt1SB18oLPK+e/vTXENw0jzy7yR0nawRhTgKqCMEmNHdemlgfUjkcbtbOT7wW2WJANQB3fF
YcSpk7AMNyCJCx69/O7TbE/d/vbA0lV08LHk3G9uhODVR8s55OuboEyig1Rat2RvxfsZvhNrSiAu
4FTE7uyjEuHJEViF5LVv2mCCIIN2SsPTCHSCU7hjuvHhuf1C3dLBHEWNROG1T57wQ4j8Zspz7g0a
WcAT8AIUM5aiUOYEpwmJRIs3cuNy0R+dhD6VOzNG6fSoWZY5DEcnOslHcXqX6cjAv9zUGN2MBroC
YajoaPWCYVfLn1heWHZCOeKCM2ckJ/88bMlMkcgQOjTaW2HvwMBpmZTgIaXThbzqD4CT9WEDwZju
waUaXxJlcSFN/u/zkl64eveQEVd6Hq6X7rBOvpnebrh2EMDXueqqQ0JlYaZyRyKwzYAjHxGyriaB
PIpaljOlqLUs2UMAjsSWLqz7dASzr3AStX0aEORNARnq1BjG6wJfn5opUlkQQW8pNit6uGsbByOL
xxaCoAMEAT4t3hrz/ZLdWczQU1OPkUIjnwvtO5LqgZTGU82YnY2+1FdgtCCVfRBMO2tFogErX2Aq
PPz6J0kXyFcuOF9h8F4vDbTJsNmSvRojGkqvT0BvTbjGEjaR6ktkdKT2QnpmIp0zyIxkF6L+PoiJ
P6Tkzv4fUkUeuTeDlHXHib020+xynN42PdVwi6zWBSRzYxzAXAEy+y/psFUuN4mHH8nSffQUpevD
JR6LiJKEiAXxToD0JO94o1kvLSgFIQmXlRpRm0jXatfWAU1rQqq4n+nh1frqfSN8wYm7oxHkXo7i
dpmSX65BLYn1+NPRC5gleiH2guEo3xOSatp+xjzn6958FABS+nmYmel4RenN1i6R1/pswae1gj9R
NPHRT8kZo9hVsO2l6k6xwk5NueCPac5KSr+PSxx7J/BMH1+oEqC3jsd4gQ3AzFV+cyBemF69ZJv9
lqMB3zLLwHCxTaOwSyp//l0DOV9Uh8j+bX/k67ATVwBx19JyEOvJ9pAXkypzpQLPizBDOPdK7D4L
kyTbeFkmwjdvhOxMVmhqPXG5xf8i8dSRZHxdz8676ynUMtbBaqk/RPFXINfgnxATuAHi78JNGZ+J
5x/rRLPLQNgI3h6MDfYQzwC5Puf7IITzN0jV5AnC9GNoze+kZgwi0O6zt4THTQLbMAAPH3IGJKZa
Mp4WxO92I2hrX0bA6oz92sK9ZK9kLycEZ2s4PTGgRTKtpwENepW7+ixwIGTmUuU/Kd4SVu0reBge
SS4W8t5COgnQhdYwxT0ibkLgluEgOGfkim2KBvwJm9wCd1mi7hUkV11lqT86xzxDoU3bDBjVnw8y
AWvWfcOdSx67ihTlEdLZjK1UN9boZm6TXvybTg0aDLJDSdfdXYGiX/1ch4x4n/UCxEnC9r2ALkzL
3/LhmSkE6TG275NYCiOaMzM4HqHOnUUetFFQO1VRxtuwHZaBLN0oqlzMNkO6HmjtdxdrltcozFOd
CSN+2qr0VwUspZaho23D445lbJvtpeVSYsmaBkdLFGyz5MRvg1VtpJkAV27Uyjqce9xuhpqzo7Pa
mSacDzSOx0nGFUr4LwneQh3AQ9+Chu+q3DZLhZZUO7nxomq58p1N/8jyHh1PiGSGKBVqPCZBtcdg
KAqJpeIkfMJMx+isHZRs+m01H/Ha8jmjLl7BeV7bAD6WtlrbhhvdoWJp+xeqMzgoaKzgcSAvGMd9
ZnIzsDquPNTDvrDXSj2MyNtpNWglokwI0jsnaugtbeBCjtgEXqXbBSiRzhQdb6G5OlJ1/jEziYH0
6Utq+QxdNcnCC8R1oVykHPHOVxddoYWvpqfHNKK+Nk43ZgRo5fId1HR+01m9XRiNBA790Hijl2Bg
xtbw8+TvaJvqXJxku9eHzw3pmnix/GpjQTqvexqyH9CSRE41wAYnq1SbgtRafSfDqk4DP+ydxxIz
l91eDtNJ0NYBFkiYASxv+mMCSKe7Z9kONrl4FpOvuLPYGMpDMxf+6PjKDguFXsOXvytQl0VWDB2C
B/I5zmogK1r9FEyMym90ldr70CgMQ28FLACMAVUWtspAM2EIFNT7Iai7/ePM4vne2iUsAS6Y1Edw
gw5VblMZuGrOjmjX6xDIc5KVqGtC5KDh+D6DKV7MAzbYO9gxO7e4QgI94spyJoumPCvYxuMl3rv7
kfu0KxmmeigZ1NMfHQM/X5cm5uEZMLHUbBj2iebuUpdnSp+7e/DEDalu7pY263f4xgB3/cCQCI2B
zXEkjDEedKsxCcb+KFQ3gFGR/Lk6iO2Zv3v0AAP/OuhNde+mCcvXpVy2lUu5vFXyfXd4Le/deHMo
fMq+vf1CnV6pRcLpBNwJEudyz5jo06yaqnxwR9oBexKBgn1kFpdy4Kuz+bCMaDdVMRaf7Z20JYHE
7hZTJtyz4YqbWHvRLhrbhgK8gfbdHMrdwyehzLU+uFfda+AOZL8BsteCymzJM6IMpCALBtNde43w
ntm1CPVhzjaoHsnGqXXnaI4Mg68hM8T95H0+e6ldE0hOrihuEMIBM6vklFx8+Z69QtJTo5owMwTF
yuFE3VuhXjGsW0+KBw08bX9ggfy2Hhw11FsClnuGK3jZnOCX8sXDGUKswE376EVFkMxRyaCU9biH
CJ9oJmzfWkI5Aiqa2v8oY57FD5Jj/Qop/latKhSkYR6HZz3LfTq3Doe+xtfJSrlE5QCEioZLKJ8Z
kI61AyYFpHYOeYDm/coF4HTYa+hlm35phtt/ii4fP481X3AcqLM9X2GhaR1FH1kWQC5b/4cQqbJ2
rcQENWWcaN93PmzgdSVpILFjO9PSVyycN9Bd2+gc8EYHI0GM3FUgxAxoykH9XYDbxcZ8GVubqklo
4Hq000Orja2f7DZFCL4fdQ3t459jydXhtHdf+1rTX74rBkc4N9j3P48GGbR4vlTxbDboBlav9Y8y
eeaTGVwLdfeEl3AESyBJUc5M7pjHA0CWWX8t6RPyP9dj/qReRS2ZEmvd675qSIhS7TGEwqK4jEXR
3e2ThGzMdVe9HgtnfX5tBDhrkY+1RL8gOmXHgJas7/6xAHPETjCcY9dBw54UpJdgOY9bKt33Ma9g
OZ+wiQ9pvl882ji3dDJijgE7FskfK6UtKYryBngLvbYlYEZ3yPysayNynFigGbzBrmWxumwjSJzj
u9R/vRAL+mV7Ue2FQxUKy4wIJQslWPXDxtHCayEl04Dx71pNAwfGtEhwq2tDHcpyiaABNXUgvn1j
jHvk6KvHI4M1s8wOBKWw0yliQuk/tP+4PaEjXqqeAFoOVhVuoO+9Dadg3RKi2XOwetGx29IqKBIC
6etQ9vT11KteN1u/Mu1FGzXoraIDDpWWkc9UAL/TXInTNmCIIR2yivNnnABP7jWXB4iz66MtarkX
kwRcwS0vzPKl9hFO9/k6zegfty6wq8T0NsKT1lX5MwogYuTIIPtwevhY1GHVUhKwzgoua8WIwMr6
QSeQ2dDKyVe7L7SgcFqXa2EY7uIT0W3bgsG4PQMcD/27ZIHI3IAdREZGd9GSpXWnCl1nerqhwKKa
8ctQ2eb0jcS3C8iuyW8v4C5eLjimUrjipj4KurjXS2I62qo5qpLo/xM9TjyHbfZV9CIfiU8jJB2+
5jHKyMjJhVq39F/0r5icHbTU3MMJPZ9x1hZuihB+rqCWm/4usZrnwVdiyKYALFmOLxZRjNZMC3sU
CfEMo53eifOf0g/NwbycKQje0vMmfHbl0i/t64KxETVujvvvnBvqwJT9zmREOba0utj2Fa43j3Kh
Hf9SIH4TsKBKy1xOOeiNcVgwjeax3ItnCi4nLZtF9G8PKP7Ml0E8HxumgLsb010sggr4Nv18gn8I
7vb8jhE8ecDFdk/6pc3shJVSAJsm+jIEqCUXlvHakNGa83+zRBVVa4lvKRYjFyucGM3zq3wTHrzT
VSWrajG3OMRJuH5cAbrBNWD7DRqVu7mYVIqBOZBFNcnftwzaVvK19JTh9TKSgkE4CjHA3dCNLLve
NE6K4Dj0q8mOb4UoZ2RE5bNAkHZgqQ6wYPFgnXqaNylQsFXAb6luGRgSWY+Nuos9ZyFL46bCKJFx
clvfAroYVqYMsUY4Y0YmxDdIroERNbRmRuZceuFGzx6u1C9kX0ysUFfgWiTWqfPBbSyuI6Sv6Aea
NMF79f6VQDArCjTs598FJmquXpfyddAjBQbPpg92SHBepHudG77athmKGi3U/rwcE0JVcaAM7V0c
Pf0SqobFbSOqzM0R1gMnxxS2lYwOUeHKYETFu7YtX67xXq6uj+snynCw61VCZvdrX1z8gwM+lrsR
SFhzyT71on/Ycv1SIijKEUsZbVj4TeDSmDVTzv93fJB/SNBiMpsjoHW1KVyzN5upKFJqzhI9XrjB
5rTRjaD02zb7Gh9Anq4kYExYadO+85Qfa7BBwVDWdGmLyqykXm32W9AmuXF1NYV0ws5RxfotAKIf
e/vzLZCJpWouJCJ6f1QXUavEX6vX5/a2JIesbfU4mEfXiAKYbR8+8kp+MGEUnpJaAiuausYjKtWG
zMk9RI3a5barcsr3SV3JyyRiRzv0YAzMmCZvieaDfLfvcHvqLvzS5sCzR/Y1G+FDslymSXwJscKw
SN2lIhdc4jcKWT5hkEGGE79wrIC8ZPbtEx/ncV0NW996c94gdRTa+eYjYlQyDiUwNWFogbkQbS79
hFlt24T74DCcgju6yKO4V4XCCg0tjQb6G29Gl9hjWR9K5EZSEeBppRbLVqOecz1fevyr2BgHi+0l
h6HjC4jj2dA80OmnmEwYgy6I6xH386GUpjlnsfeo0Lczp17lI9B/wmazbdPevnRNh1lQ+etIZL54
IgRuBvI0K4opwVqGwQlOFfyW/zRi/o1QWzEPhGFy8fHN2TZpQ/MwkDX7iyyy3fmcDSlBeKsHq0Ra
JlqZENxNUrPP7EfGruTZd2iUn20jHNNCSA71j/UeLK2OImmKXAvh6SXItdQ6WgNiqnHGWODbv+BP
fWvkSTqA13g4TiZmYK8waYkDcxIaYCFVmkhwUUZQzEVzQfPKiRejtoSxiDLwFZpD8ObMcDHCNoNK
q5d+czN0a3xYKiymogFhpneYZ1h6uO5lAyFt1l4gRvVGf1lbR78dy5Jt+UYnD55tBdhWEqXcXpIt
MTipWPd5ZaBm1ExhtrQx7Ge597NNMfXIEOi4u3OC1V6IKOykHyurYbFm+WtRrmAygMQ7E4royw/h
1nwfnsb2lo75ss7jLGye/jjF7iY6Xn8bUJLV62Tw+j6ug47z3JWuv4bVMihORhFkX64IWWDqz4Jj
pmXvJl8ZO1FDyCE0ZrrMx/pNHIn/uY3/MP5ezg5BwV4gkvpylAC9yQ8fegi2RcLdFqajjuIw/wxn
jxXDENvlVJSCWlf3WC0PRfUsrezwhkU8zKlGp28wyHqIjrrWane5VELn6rnvvVeLSu9PETZm1f7t
ElrQWHu/PHqLxVL1FnFDNvr82+UFHu3m6ElRjZBBs9R0y4IZIEPGs0ZrZUy/veymGFDACxN18GE3
tFWR3RaS7sl0M0p6DzWkjVGZ3ssxMlSmM7Cgq3W2AXEM6ZowCeF5woTHBUU6M0GPvhaDQSGYfizR
YMBnXEjhcDQbAO48mMmEqai7pI/CZydEKyih1reN/Cp5BTlPo4oImoyiXUxu+BO0uIWDIVjC/vlu
q0AdYRtA4JRHM8l8evnmXbYrxY1oYrkdP/mOvOcYztDFb64JJIdjciN3PpRMOm7aDnlbVToDWc1/
wIaJ+b/lPwyKv3V4tzG9P9Z/O1Fv//wAI7Gi9/ACyQn0H2DMuLaxfQadVPUu3HImK/nog/eJF1FL
Iw09rSqLx176bpGqxT7LNX64y77HkHbE0fyzgYIpS8uhlVLaw4GtDR+wcIHDsNQrRW0S/yKYlmEX
jJ5k2XM7h1wFh0vGCQC1NVBqNbXSh52LYWQ/8s133q5Cu9YOU3QzC5l+MMadI9cYEIApRPMcYBIj
ON2YflZ/hquna9wQ5DASBVy+Wol2dr7wKqW/cbBVT4svWC0GS3kXPdmklPz8oFQ9k1gV8igV9yoz
NAHvl0GVyHQWmZ8u4nOaSZtvq3ZARRb5xpgwPMiQWJL5NzmtXneePEBFd/N3/CbKCB/zoTJoGCB1
dfbEyg0utt4hMbRxTswdzW8SHBCoLIJGM8wbk2kwAVRgrv1ClUn05yOJ8/7lwQwZDVwvkgMC0Xyv
1lUh7CfmOWZjfndZemJei3FJWJwgPPS+uHN0doXHIfW6tfCLz6n3AEcAoPzT09dowS5okSHdCDWu
Gezp8Ja139BSS1MklnJS7D3NXfU5ioiOQHHn6CYmpvige1AH88LQ5bjacWZkxmg+j6dQBBHrHflz
RhZ8ldmSy0MvxVcJGP8uxqavYbnUo82IzHQzDYaK13H84/fQUZry1GwtVrzXhA5VTAb6ebNfFy0D
7wFE8vagp9XS6h9rQ/zlAtkIgjNQp5gGU5K+WdO7MDHGDEsasuHmW8stxbUv63qinpCsR6hWmJy7
4KlLvKVFVGBeceY6Lt3kVEm0KVpYLu5sptX+J8z/JV/zgyXYK/bOJMwcGj7QOAKLXumwaG+rNNA/
bKhaCszY0fmblWqOsUDRPatPDxIQqk0ewOtvaOwdL8S2bxmBQM1q+OdxNFg72+bZIpy2mQymWevd
xtEduIIilX7mTqDnafHanXzkYNwovOZmZScVGqYLEg+LSjzpVldamQajmYkIRv4gVKwko/M0q8gQ
lYeC1XDi8aijzyN4waBucbrxAhelhRo3YcvyHd5/cFiMn7Z+cx3WXhRaPiawOD+vaY76N/cayshq
oc93wB6s9KLSgpG69Ae6TVUHZjHdScuSgBhf35pbm5gbMFMs0/VXQovv7IBiR0frl7ys/xkGo4Bx
rs2KwChg33dVo5tpd1r1ZZNSu5NZE4tXgyXGPzfRg3Xj/2rpU+5ndqzEQQ90dxClhM4gFTnIAHnE
kd7brPfjfrA7EazdRrMlsS57K7B3sKK/vkLqLANHrl2Yyyv8kMeOzIB2JMe1pcIujQImv4vK6oiE
1BdoWtdB61qKQNOZ6pSHKAsawTcUIw5/LhbpNfWEY+BQ42S6KytgRa+WmMU7e8SjkqSh0eBN/mn4
UsJjQCmLzNXfOB77648+tiKvIabOupnx6sPZwNK6j59bWY+/7CI3HlR0MApxbLmgZvtakGO+aiyK
LxfofouZcG3KJiX5F++1rJ0bMv9+n1u1+HHer3dg/CBt2LxrqijLsTf5Ion39RizI5oahyg6YVWh
LUOkJVN7RPcpw8qmR7ltx8oW+AuskE02Ujtw2XyAET3P/xSrrix+AY0ZVeHrNCs/jvXUeRnBebHZ
fpEC2rziMKRct3HTrp6jTGUN3T4017Jyfd1sVR4f1QBRA915YGHDax8eRyaI7iWe6DDkwPjjq0nD
ZS+QMf0mM7/IZhFoAzLRGMCCOruGIa1zMOD7ALMXdJCVUYRHtWPweociSlvzm7E3Q8Ty03WTwslf
FOKnms74956QZqzs5QASlmwIESn/sZZVbChBmRokLVJ3xMkZkQifCAT2fAibOdlc3J0ZvGQdAp2V
nEV+wCCe9RqBeqEXy1XbMfJBsJJ7IlKjB+nUmK/RwtBpQy1PK2SYlzTr2cl0Z2rPN3mKhI+21h9n
e1+oS8rTzR3CDAOcfgE7EYqNvodDIdnbnLEd4wGxnRupozboeQyxIITh7q0K8R1rp1CN4LERDmA1
fY9xcF6VJxzbaUai66kbV1WTBpOrquFA7a1o8kAVYX3jEyALxKqMwUmLTDJdlypE95nCuK+eDcf8
Yh2G7AbXXys+qxPe3YBpUcjbjtuBUjBRN3c2kfFmw7nZR927gzBm3dzO1hm/2Way+8PY0UQa27nG
Fvm1b/VrPez0GfPt9wrNCNFCYCcGWwnr0ZlkWtK9yCYh3+NVLcD42CucrD8dAWBK7uFvzGfnmOa5
X+71cNG/ObOdvlWbvHlwytD6YUGTCSr53vwxlYNcq6EGiqRZKvXrhQlaE5qFUASEdXZAsjeI3W8G
kuI5WW/xhXBFDNQx4i1Otki9Ak7c4yoxLb33RXADY+iyQvhLSwLIOFwIuMUmau/pQ+Sl3h8EfjFb
pW+ihf+Rkw86D2QR7hQDUxIUH1ZaqUllm9c87dsTPZmGmyJnw4twricfn1lAZ7mrn7S4jP5BXHCS
0reYy5ELBPvy62TGt4yfK6UMqgOTV8k3pRylEDvBHCpFSUFJ0+6UI7s/47Moirc9bjL3+IW3SPLV
Lyny2EPKTwui5Rxr+C4dC3kNO/YvHuShT30MkoBtO/RvzMwF+VcT5UVTisjeHd+8TB8kB5i03WRm
5jSDtAAB6YLUHjeOtaEpjmBJRbhbbhtLOf9na6/GJyzflidposK4KzcOnzsN7xvqAWImSJ7Y6eTd
d89EGQjlQog8LZ72Ug8l444GR2oPhwagSWuZy9HL3MYWqeGwfPlGh5ug7tTQyepo0FbI//LucBcl
Mpz926v0nePNbVFG6QsOLGja7zf/47AlqARC/RSfnOyi0Q6Kt30IIOZKtPFeMDlfHjL5siZL0i9E
odr8lhLjoOX7yGsyphkrXZiaY5OA/jeYjDhPTdjzCBvkSy1VtKACcGxkSjj0IcuZ68P1NTfU1xBV
qj43Wa9xUSVD3GLMmgpjdnyKzQvMHYM3zG1RhjZo6SlFlGCaqQ1cHFY+m3PUJJSVwbFBRRA0W4Qm
cPmmp8RpSp1CLZ6yv9G/WxzusgjdUmejPpirz7l1esrw8oNfy6Vjv/TJIA/rg1YxhKuCvNeAzft3
bzD3Tnt/KdIRN/X4hhwT4UaDvrNy+vbEFZRuN2fdoaF52UFQ4drmt1mvNonvzjaHfYMQS292Xl/0
M4YyiR8LhIhXpediQTVYTEF691xc+oEeXoVOZV1eAQSf16nCWqTYrT0Rm2JNMoH3eEaLX7HAGT37
wasl4i1jN/52/x7LadLV332qcLny9kzefLdYoE6hscEELZPMm/wkgjSU5k3uy2ADJDdIg9tQiUVB
T9hFRgU5mMDprEK7wVn1bTCrmS/eFCrMUmVXr/QRj9odzm8zJ3RBUFMoIYdeOf6xFlc9IkjlTWVs
xldS++OdZ7ZfV3ZOArPMI/OwUWAzN2AcxM58RlIGYeIoI9+8TUTwRsqkF5+I3PhqKeT0LgNFOYh4
tiZE8Kmoe7ycqElH7hWkTWCdNM5TjNlaMplmc5TLdT3YKABd8QWxghx6MIfxz65mhgep36OSlotr
txgYQLydSCU+l9o/XjrcsYh7W+0FFjl3cmCjVt5qdxjG1VituWX1F+AD5WSAI57WGP640BZPpOA6
x/uS2O+3pUns/7YaU+KIpdYVHNZsIDCtJKm6B4CqQcZEVWAQKZt60s+p5wvQCQob1UAxAF4gYyKk
mCmR1M5qQjyR+fmLnRqJHvt+3H/C1cLu+das+9ksQibdXM9m0lBLCGFdBkQDESs72L+79B31n8hY
WHBP3KIzwPelJckM6+oYui78NRMiTu41ZknULW4XTZ2j9wQ2O9MQLwoLr1K1fHOGF2/rYPq4QpFW
G9OxmkSNJyV6RdCtIVJJQQwL9uRKvmlhUXstE3PDvH/8axbnnvzcNZpHf8tuMYHsvu50E/slEkjj
q1dpdOeOIGWsjUhJo+l3rSgtu/RD2Gx36PyzCXU3x9QPM5z6MJz8FQ0/UabDx1GQYhSvK/FqSpUX
ndXUD963E7ImA68x/6lGZ8rZ/cnxPHLnAQXSZZfUV2LCC7YOdQXgvXjhbbwAXaJJHU20dMb+R1/j
nC7TdDVQ+RuA93Jbcehk5eM5KRd5CyoOTRP9Ks70dTPCYM/shrA4IThCMsCi0AHG83HBCV3IjJDy
BBj0UowXIxKdDGZyrqUuX4F0oRv1Jgh9T03xIvGrzp4EQIdcG5drKfuREDsqe1WP0bgZH1ygsAUV
mk4Rrk12j4fdH25ccQZhYWbgzOY0P/Q/J5I8Z2gVQQy4lbARUBpKH6dvSgFHebhxtit1H3nJBqos
W3qDW3zxH7Ui/boxksGNoV61+D4or+zUjnDapxw5KxgmUcSfd9GhqVBHTg/u+fJ2sZDz2MiCS6rl
l0hZHlWKLndf1C0l5d1U82GWh1g9V2C9DSSqU07zCsmgSorGhqt8X2uaWxALtEiQUjink2KSiDb3
6IZ3XE3OSrwCA2ywYyfKx8arVKV75oHrUuYnTyHtIg5hVDzl7UI7smPqv4nPEJ+LnPX7+CQt4Ibs
ryP+GqCGmJl52ikSY0wTALGIFvFCxPaOshq3Mm89T7dlBaJZCqdTONSJ1bXkuW99l0mKzp7Ss4Hg
mZeVBsomEQDkK0bLVpnCCKbZNKG/pDSsanl2ZtrI6qvEc15bsz+KJ/wwG5+hkZkV1DaTzJZCWrqY
AoH5q7kxk6rOhpityyvmj8Z23FYeMT6xR1tiLg/flLZF+14yecOLLcqKfqoqeVBC8r38pikioXEZ
LvNgwizC43n6+zZkvP3aAv7dGzDngFbs0wYlMsC9HCRjDm0zp6AQGKBmmxr6fRngvPiA9Qilw22P
HbGyVSCBjcx5pEWmtN7mIUTwLl3YEqFOZzwXNDgckg1Xdsm8nBDTEthCL5Y03/4K0LOXPyTNFmC2
jvIi8ghcUMhn/nbyPQss/GzJbM57uEd8sErv54W6EY3+7eFROkneTEH2jMCMQd+CAR/K6o6jdNIc
ZaHNMLvKfpbt7W1a39eg/J69qzZOxOTXJBb+exndLB7HZ9sqxNt32W7nBE53UElvQv9HkTgREMU+
xhLz81aQnmV0nfAwGGNKOF/nrgPYhM7A8/RnBk6ZKLR6XZE5bnpE3453cOR12WlONQiOHXxVEdlJ
LhlKECPiBNbtUUmA11BT4/3sG5StHxC7hjl5pR2pPwQT8NK5bI5oBvV1YyJB+ePZC0pMQRJeGQ65
RAxACP538xc05YYlo3/29kLibgPXGgyQg7f37KArS2SMrVGVxayg73dd4xKHMYGjDBnsA5ZCm7su
Pvg0HDyydEF/CjK9OkLdL74Wj6t+aMCbNp1QdKwxhY72LGMwOXK+WeG8CZkHVYJwz2yGHJKXYjqS
MlkD2P8OfbSWlSXr5jWZ/pA/LeiO/iMQQ3a0B0KIC8/0zkZch2N6f1MpnPWHzHqHO7QCZJhZwWQj
2Dd0lVMtl+WBORxbi1Vq2hBx5TdwFmYPOmM75CmC3PU9T9IIsvXeLx0CIlBv/IO1tcVjNJPNAmTq
28V79Bgm90FKJtecAHAZgQfwb1DvNLv7SX3zg4bMt5C4W6iml5HjU/vMabiq2a5oV1a5yT1mThb6
+27sqwd4fDMnlEY7dpDgGIos1JSRyXZqiwzt6WxAIAP7cEGAkeBi9rj2BDZ/AqhLPq1gwdfAH/Vn
4oijG2gyNiMtJAHd6/Ki0KE+q6eW01bvF//PQraqqlSfcU19/MI6k3UEgkbj2GXjTmvvcbm7s1Pi
InDJR/CFFnPk9zgvF5RXfJ0TeDpvoQfhsG/MLZjgrT2Hu3K6Kyilng5m/K5EXkK6acX3XJ0elsMP
qjLE8mE+NMhdVveC2VSKXTVbT2kQpZKlOx+/CPGZ52GFyKtotLgFCG2faRyMjcsxXGs41AqOMEAf
bqRn8lSDZq48ivCgAfYsPMWC8wwneJ5ZgoqlLZd4ru7nYcJaITVTDPZ34WrPp6Op951TS1+381tO
A/02Hi4re0NZSw00j6PBpLC7X4f0QUSfEG6yRNeMjhmLHPZUovET5eQ082aqE5o4WMQRN368cKT8
JHp5i2PVLf8SoKxne2c7lIOGotj3RRDzcvXxBPLvCW00GzfhgeRmervbXQ/fRwBnb678Gl54Dn3v
13TROL2G7dFrYjVGFkYMMHb71MlIi2p6FgGPuih2GPX2coS4rGhHBhrI9TNA0y3K5mXMr2r5+eDc
6HfLZ2aF+GdV2SyhS9pXuE1DfpwtCW7e7BcjfLvgT7X1unheJI8il0EEKVttkTAJjfgidO95JQX0
Gzs1LOWnC6y4q26jmToP/rDexF6RUMfsIPLkTfypQtAgEJ6HzxfGCUJRFIISkkBuePc/NDx5Is1d
yESPcciMBjC+mCTvkyUKKdxKu+hthzkk1aT5DF3fxssq5jZy/zv+ypDd+0+peUIFrD6NoHsjgUeE
MTPN5xXadADFSBTZFRTXBpE8pEehO26GLObn2K7lwv2vVwLoUXP5lpY2id02OBTkZHs79l6AR576
dH8vVJppNKdA0XLKOJ1+4vjEOY/Tf91DeIvvWWQfUibh+te0mp4fBJgJ3SiK+R9vZpJAj028qfeD
YFYcg+XimUWgJLCUbkFiU/S7wu9VSCHtnCWSZ+hRwtG1SC5yzpMkycAfIzRvRoBTf/TdZRlDbNMt
bxkFyca4yi1GNWKbDHD9cTCXd2HM2e3sGXa+BWsfi82aYm+06xanPyNQmyBTQeqSkzHSDj3zrKrC
rH11jOrzxjVGByrjOKbVSJ/jRRwhEDN9QnkcOolg8HqjutVbO3heJBVAqHwKlLygF4HIpM7cPec0
/vT8TKBgz7XmficWPTq3PLhyU5a1DPA3vL/M/i+Y4wBcT+kdmhggEYqPaBX1qUfeyuU15VqM4AuV
Uy6QMqMJbwR4DcLYCtuwEkIHoWR0Byz3n3OEE5rsvdRDfEuDypwH0ZcSZzffBMcN40x6AEs7q5wW
bJgTetgjynS36DM6oX2ovCssACt0LRHM66+jw+jfU5cdwXupRziVfjNuMNVY5okgF6Tp3/QGtGyQ
fNNbaDHw8VjqED8Bv46UUIUiixhsJX6+jo7h3473QA/T5Rv5IVuVHYDKEgPeWG4gQufjR39kplNh
l8Hv1j4bf6o0SfvnL/XL33CxuFffPHpjSiylhVERxZQObg1NlzOCppt/UbSjV1NniT0JnLv3fAI8
a9IA/CsdT9LtIiBPym6sqesnbjWwkxcxGZ+gKejKqxd3ORS5Dq16dlCAS/n2AVaF1iuKEOoTTiS4
a7bH28OI+VplrrAoUNwaGMYesY0hBO+yO7oMDJY3aaCAyzfdDxiMfJtNOf2LDmLX6H7jc97mNZTb
aNTeOYzSY2S0VrMSn8u4hquGjiR1IrHrq6s63fj/RrI++W1cH8i3S4VynAyLXmQjFnwQ5Zbdwt29
sCA5YNWkriNI/Ku/N4vYJ51fPTgtWYDSKHZwEaV/Hfsr/W34BApkNpjL3oBUCkzmYjmF+WrJ7wze
P51U5Jyc825thT4kWQSAKcW1bjVAs8kdusdStzqTtmWgpgvk2mLuucEgsK6R+A+Y/zv8d5lGcvuT
cm2SqJ2ZmR8nP0SDV/KKpFtfVbb3Th331TR6jGePy6WHzGI9u3ebq1Dia7OmgkXlYY7WV/Oxr24L
qRiTmwZhWSb6MbEPmBb6lN7k/iQc4bNEJXCRo5gocfFOjPGZiZF/yYXe7/LjkVtJYfhg9Gw716gw
jxyv0A/KZQZ8CSSt1RcvYIvvRE9trtSA92Lt9W97mqjWwH1c1FZJ3z3pW2HEXDfyO/htX4IGKLUi
JMNfmB9xq/KP8+b1A9rooCLyMPlVBDgSbV8evrMLituGYDBEfFcwl9xxawet8W3UezPcEZXgomwq
BkiEtRpp5e1Stlmys37tA1M2+Z03qWa0yivd5uDyGgBc3qQF/HocL862B9qk4n7pi3GtiKM/8SNl
5RRmifdW5hG92+uLMFpTVsVL6Jhu7oLEuBtTgjhfPgKemJALq0ignBCNTsJIpKuWMFvyefia2dFy
LpHGBXeeL6rI1tiy4cETXQBspqxAAqgr2bhb6KRe244HtA29fxSRSsIRhseK0teUOMcYPbjzTRK4
sGm8/QvvylAisdbXmDGq92eEcGHiNKC5pIBihmXFU/kAQkpmCSsbgnjAcdyuElCEsjgAIOcpKow9
a5vyrO9/rUrc+KsaIdTpy8EuIFPYEOjf0fjYLkcsfiilHM/x3vcXCWt1HlvnkVtrIhbeQ4YiboLj
pjoNf1+GZiaRtXzA/CTTNcT8aBo/L4rjR1eHYAUt3OpHJTJJD5N0ydgG6piGTzs4k4VE0bItQhiJ
F4HkuuwOxR9OiEE+g+M75ho4uaMEVa2nnyRpbiTuZ1MFrxW//T7Gsi97JiYj9jZ4lprSBWXONRYm
d/NQzwwVPICTRze4qtOMccWPwFd5P4eyb8gQ0S6AQUpLqfNXFEi2CpMnUCSNA+hkMyQQmpYFYz5j
2sjffA6mg83RVBt7GSlbxc16mTW2xvOMwQMyDkJ/803XiEY6FKXdyZ+f2qABNpbMlRfUvjsLciGi
5PbF51Fke1FWunG0MeYNKOA74rBfD+cgU88jRQ562llFy9fiwWzGTjsgHRpD7MBW0cF9CYAOLYzo
V7E2lgebQ/6krV0ZgV7jMKBFNcy6SAOxil0Vsx7BU/M7Py4tMFuadeddGJvViE84VnbhqVkdyNkp
1yNVUCZbYpC8h8NhSWVvksmLZDqXZ262uuwJAfKyT7OPmkjsRU92lLUvjVXrm3QJYs4soz8CFIHY
VOjkMVVyNaYZ0syjZeo1euzCHxoFRd0S0qCY8goyZebMHGa0OCmY7HTX4wABqKKBnNdTvgQnUo2+
28XVi6VLF+Vlk4JwetNfeUDAMyQFBxdlsKZ2He5RDiYa0L0nXPFNtH83hBf5/i5HQPH7+PxwSv84
NGDI9naAWgAoO0Itlp/kbNfLdhKPZ2kiOWKArPGyVMhO8czqO8ILUbUFISSmSS+lp/+IqTE2ciFZ
TK5a37H5wPYJ08UEgLa4O5pMYHVFbYezCyk3CXy8ITV2XPaTzI9XTzyMNOvU/33K8sEqTUqodGGo
UT4470L6g+WKUUOCLPonbGFCRNQKgBRZIuYS8hGi6X0NSAIgftBhGbOKWX3qGs9bBmVcPlUPmLob
Wh4D8SyGYi9jqSBIMF3ZYMnaK87+cP5I3K/v03EoWq9MC27128ZDKS+qLeGTDOTkFOiBrWhnqc09
WBv2M5TTN4TLb4q87xWBqmDiIujP+ikoR9dUcCqBKXUOaTETLyaIHfM6TCW0JKxUTXQUO5MLXTkZ
yYmiMsaZ0RBD4Ji9qBvKTsvXmdKC7nVda00DaOzx1W9bwOmY9i4NLoVuC/YhxaggmaAeIqra0gYo
rOJ44uZr3TsDOQU2ZMV3YsQ+9KVM4BynrbYQaBPrLoLXmimr4tiY4DwVIj3otLb9gPCdBJ9Q2TdA
3YSTs7MbibMTwxfdKINR0xe6A/xCHkqTfj9pyFH2pUK3z4tAmDqTAB0Ne9MwTMzmnoslOL4ScZYM
LIYy2cGUyGgi+iZHYCT33tkmpkXV4GGoj9P4t/CtsymzBcbqu38OeqICa2KQ5m+JQIHO4eDhlpb9
NC+obLyxcooIusPN2pKwfkdaG0RkKxdnqYoWovoAXDHvy3vwUTs7y/B4A3vfZfXgFkQEpNBIqGXO
a/lmbPsOLpOuN7MtN3vOsdusA7JBZ1spfxJBkRXbSEkeUwNqqwBOWg82xb2me2Ul/nI0FFfIPMAh
hxm/4wlRI1XLd3WGvTfU62tLuXr9i8W5vIUp0v5WYMOhOpjdqoG+wWWKxBJmwCuEg44+xkMMTzFR
rIyM0sn54uYjJYfF3odfEu4QD3ubqVjrQRteHofSQMW9gyJ83LiaiA3iydhtBVp4YvXFekKRhNG6
Hua76Kym4Vo0442/WLarVx6ZyYelV/9UJ5Y6+JUXk9DbFfltyXeUj/tcgeYnoKZ60bD5QyFf2sRX
kfDR64pkT3UF39Ru+T8Dkkf40BevOjf8ow03kXssTPFdg1tDB+8jJkWeeIEd/i4TskeSRC1uEoqp
cECydYHlHUNoIK4/InDPZaIGka3KDeHh3+eyVpwYENzMsec94eF5W5dl1O9rKEcXJKg0V74iZn/V
KQHGiqA1tS4p8OEch3Z58726COa3mdwJAE9dG7bs3aQZYbqqOSZG9miqC+ujT6Oaz946oxuj2lSi
qrXROEdgPs5KtAoXE0ZbzUaDeDisd6DKPAziFTmYXtqo7aDZ7Q/68aKFBd1gRcc4M6Q7gLNLjgwD
PY9Ccz4l159cm5cE6YsEyZUNVtd1ekQjMcFMX1mKbZb7zXhrb2UWpGZWETCCFfQUBu7QCC9ofYE/
pVDBYfr9oOKzZFkUscWcg1us4lVncKyk+At4hag8DkRC5X0Lfry6kRSD+C0b30Fj9FHh6ehVAQkX
gYsRmrqG0lvNyDKsBrpmGFDvc4Z6UtYm+mjXqbtYdPzKSOyXCBDr3JuLpkl1eHu9kxihMdNnouJ/
AUuAZTIDX1wsaskPYs47uFdUJuKbXZ2OYJ/ryNU/CxN0w+AAHL+yut207a6rRjzjJWtZYgubXyp7
hbV1m1JVdh+iaUwS6jEHw2NGS3pngiXWUKvgGNhEtC8Nn9LmSdNo6wcu2sqC7IBzvLZp8/RN0uHO
qu7xGUjq4wFIYwRmqhLkOPn6gd5h4bPa2KeuC4MXec9U88cRryodSwLnYwIvrFqSaTopUaSCEkCE
2MEV0hhsBjpnwX5xIxtEx1KTCb50qri7u01+vjFM3wwlQ1rkHEszJchBTo8hW7xBQVLtIELNH9Kk
QiUp51Blbg5fNIPt9a3ut6Z8U+h9BspJNODnZ6XocbVfAnOdCCCxuZo8hzPGuTOsXdjW4qbboY6g
njgVp9yXM8oTamc4X6ybdUQGS+H86C+dUVOhQFqQG8cWjyMN166IC5LDL2lFqWj7i45TSawtCuUA
S1OwKE3vkU/B8UUjyTisZ+GsE857Cke1jQlW1U6fN9g1No/1aCOZRL1hYaMzfIcF64xR6s7d+2m6
3slhIIM5yaFaz0XegKmfgL1iLBKbMnvNi8XdvnRwtsMN/jAxub3/L12TbG2mOYCTk5LgjXrsGKhB
/LGpM5gEFky5CUlrCF+xaCDyZbeDYiNaeLvHu5G0hb1bxZvaAbeIdykQwIh8cz9XYvCjB6m/ux0z
Kvs+0n/M66Uvr57AAxWGma+Mj45eeyDMvKHvLJ2PHpmEI9Q+lLDeCa204IwlPs8eGJRKr7SLrQG0
oP/u7jx2gXrslMDit0p9DG1GaGrak4nixg4pDtugUNaD1I+LyES4dgqBl6KGoiaDB4gaVLpid0r7
kwAtKPh666CcNrToBpXb3Bf/TRWBP2aqOPv/n2mPmtvK/ChfSLHV+90QThXPiUY4Q6xPnm0l+PmS
ambZJB2nwECn5FGqmogg6LWVMJ7KvQ82croGMYfKgCZcDL3pXLFQGebMSTdelBZGXady+uvHrfZB
YQPp4j8zwmhrJh/F2C8HSCXRqWzhHbZsG0HI9HfE6yHBTW2nSw/k13lNGS3iJ2JKH1CCnWYgEa6/
GEM34weUXwFnjbtr4/MPKYF/GZbX/L6AChsdmfHZXRgjXGKZZ6jYtuHNdvwd05519WDSXqbbv2Pg
6zP1V8Qv3jr287jh+7EL6LpCM1idorNne9CwmPhN2HH9WczmGzv2A6KlgsQwZRLLTEoVFl5aYvXL
cuKC8kXvRU34ShUyeGcvsBBQvGc7Gl5X1TIBIB+FKbOMylWg35Darujf92kMPPa2zF6cU1m/jvcD
dEIFcfKO99TA8w/2OBWWlPRMIFVHR3FHZ1svAJsVu3sppT6ETxp1iJ4TRufaMBIhoT7HyARRPr0r
ODPMEaMBwizrGHCBbZs4x4f4haUJKKpjki0jlXkHv5HLkNNugFm7BwhJHFZ/IyGG3npdavUPW0HY
uwvQzRTz1xpZONaE10TRoRgwdyvi/uOo0RaQEyMQBG8RdrTeBCKO8bvzB8da0VeLy0cGh3yruOy2
JDCu6i10t1GWH/w7SJ7/n6Ny9WFQ8SlZjzxVSVdwkif7UM7M/sT5yVr09tXyQZjDcmTGOrbPkkBj
+y7QBdeek5POb0BxqCgpWqKp7b0ICpIyFUNIMFqIFizSjIi5RLeS4ZjLpja3nta2vLcjdj0FgKxr
foQTLsidXR9YMpXa6c+av/PQWt9Y8SQIPi3bFtkssYr1FoTeGFMytg709sNpM7xsgWHSIws0UAYa
N96veGZK0wD56XCxvV3cEfYV8iVqHaTenuVLvTDnClL9P3rrcBSZ3WjTRFIPmdH9zdyRyry8r+4z
fbI6TgzGJZJFnzcPvHDWgFjpB5UrAcziwlT4wHylJNWU/ByYnmjOw5LNNiDMiHpwF6opKfhcbvSS
XYraQR1yIomp+fANh92asWP9nuSCKxqWworSoLAMRBVYDm98E/qYGp0LJUyxgWj9dCVP0wWQ6Sfl
umfpRmDSA+4hvg495R1gJRhFhbpuYW66WmJS3YnbRoQhnlIDIJF1d1s/Srz6amgSUlIcipjBdDZf
aq0lF9f+3Pi+6U2StxJpgUinehb0coCkfOFlZWRQM2AoYhAP9pLul2O8AuuOOHnGM3rXOI1C6N4j
fCFwXDKKKQaSJgEtCU2Gu3BmFr4s1ByOu8PLGGjEuq8I+UkbLKmLxlmo0XwkDbqMa7f05/+8BhR5
7WgG//RWxPbp1trCTU1BR9dK1iA1osqkR568vMa8fcI8NxSJmyWqvrPuaFn0eUjX6FWh9umHtnqK
/Kjd3B62fVfdDx2IPwe2GgHqT0zoB5j0wuJdbmmLQpux161JjX4v/PW+e2zJN+9I9Yflwp4A90L5
i0blSPOrLepn8Ow5ySS2j7G285xysHqHwgkeDNdVjOc4fHNE5LFXba0W5T9Kwj1NSXN9kerTR9Kw
OAJ42UQ+XwgYP+3/9K8XzIp9wjCF05cbLkBadRJRGakcVv2ONPYZFdefzOat1YeUqsHPtZFQdzh7
3UZXenuHVOTq024YhexH1gt2YFtRXLa4EHr/P0i04OZ/qviWD0OjlDrm8jH9bsq2aXYga0FB8V5Y
oU9ekbKm2ivB/F1bG2SkJGVww8cIs86mS8Hw0s8M9LxpwuSHXbRR5gWgvQmM3Bl5SMX6QK1iicqr
00+Z+NqQBD8eYvdkmtJPRajloltBRXuB2cOoClqFL6YakxZFrfXBeGaLLjNGUSmDcb1iIU/wR+9q
iAzp6S7qR5PB/+dEYgPPSeJYv/P9VRef9okD0U+QUrc1QJzP4dHB+clRJngB7Wj3ebT6M4BoZoiR
T4HdhVWTmvlkor+yR+azJQS28lzeNY+MLHAKKwpwfMJOV/RLaPAsAtus2CWkajBauKdCoVWSwOrE
qchhBLVx9PhG8ZAZpae/89jk/aZCeteU4R6azTOujwj/8J8KjPhZqpo8Ho6lg/R5jLmhMfZM1IhS
MazkMi52rGbUUr2ipqbEKsu6faxIbhIvQVmT3JnqX9lNURsdh8cB/mDWdHKnvtrMHq3zC6/cv7ax
6qqbFNuKh2mKWe47mewI2RUm0NKuxfKkuh0Y1KHCr8v2zug73BxyZseETPOh/gEVGkz0C+7xj7pM
AdBSu7ukVvGVgLHQN+BkUkH19g3zVy+TpmptM5RtahmOIAhFTRu6S6lJ20K5ZYtT99qoIUXzFaFy
SWqjaAd0XnppyVnWJG9VykqYchsBSUPrhjYhTqWd7HqSqWWM4/FmuM1iKdKwytz6vzYZgycMOikP
IBs2lCZIWWnzSezi6u18PQoA22eDCRElE4YpnMInpo2ziG/k03QYV2w3As80pcBPEg+HzvWh31L0
IcwEBVZi0HW03yh/d0J3RLXnba7nUkvM/C8StCATFa4Tj9dYlgIo4q3V5fiFzGDaqNsFXan7qQPk
ip/uPVL2bx4rDObF6Yn46n/HxmxazYf5by47qGlcYDWxOkpAvSGLi+P7aGx74TJL2NneqBUa5EbM
JI7GocEAF2fGmtuQqoUlmHwHcbjM53i3MdEfwzJ7f/+nlO9MntTl000a7YqgrMbwplv0SaUDsHQS
ls6U+GzSRq/Pl0i45Ro6ldiZexg0G0/7zXuXfU31VGDL63jl91mhIgZtpx3sY/733V0yxsuKf2LB
EWZV7rVVwUmVUfIPMei2efxR1N/FyRk0Nbf12HdsvnlY7xZQ9EnY1YJfle3rZxuAu0BA2jCaL2oB
w2BOd9YOhDZFFygx/1iKc8Csqp7xFVdAqt5ROz9mJjaeqitRIAIE3sdD/DZP6WcjS4LwYkIkG0fK
VOtXk4k2SHHL1Na88KvVvOhSVium1BtZrcQ/efSR6Pp74eUbsRckrQVJlGagcNcZAUej1zd5xyls
flm2CBbzsZucXhp9DHWYHaYVlcyN0gHEVZkAE0Ak+nCKo8U4ZDcNjNOlEONiRcn0dPv+wff0a1lK
k5DkvXxbgtFMr1kJ8uVbzD8D//54UwsOeDIWp5SveKOhnPnnCRJikfBSugbvZwrpcRw6XmtmXwe6
R9Y+LAl1MyN0ORuXeWj0Wb6+0ADr0JsjIPs9Hr3lhI+THN3wBoYTH6JhBeq/3H08+JlpIb0gfuyY
K3QDrrxdjFPXr66ZgD6Xa0cNr3c5L9Lf7I9dGQjh7OuZq1k/vLG9j2nP2ZIJ7qiWCOWianLtPCTp
jGtyyhK82t+WVwQzjyll8Rli0xNuLfUFEOAejvTzeTIRS1qSxvRZ7xC1oamhbTrzo6ZvPtpM2Omc
KtpS8U11m3TgR1ssQo0/IzGt6dTjj57gHcEP+NzxEuHycHGuqCy+c+bt88Wms8kQDQEA0RguN/u/
q/ceFgQGf3HF7ucZd6alqExwY1lIBSS2tb3cIFns27aOd7Q8r2tdLIIYLeF5ZaT26ZKcDFEJRdcj
WymIEeKE3/RWX+GfdMNU0cTr1wcg+lBYh5GYLAQHN9MFrjm9p8mY3rPu8qgEo39qX65vXKecsiGd
ARe9jiVba6Fjvk6lSwdgtygT2dy3Se0dOxsIHHWfhJQIWDTPELJiPbHWzrKVqnOCKh5VVwoB8ZAy
ZMG1wUPCKOIwPCUqn9DzX+bNlWhGmHvtWoUI+YDYmCGEfqokF5Oxfg2BnzIEnLbuLcSC0YVJDvsx
KcG1eXAlk59wlFiCi4aNPo+aub63yj9W/aZVRpI4RVkK9fSYW2u7sLdeXjLXsdGBHPxLucvPbYMM
tTN2rbxl3g/5Tj/8ifVaRW8zmTMbCCHCEgLP5xz1fzzZLcucKYoi28Rali7Un3P7ejSxEBUQBjqQ
dncMUQz5H2Gz6rh8iAAe6rCtZyimRZZc4o5Npu0pcudQraT4W99EgNinqK1zwAwRzD63ssM/a+lW
D0Q87e9XO8dIEo50YQSduJ8eET2UCAXNEYWywG2yLD6IudJGPcHqTg4aBxZTeAiA+SGcygW4vSew
2am3NbojkW6jETe7Ynpd8CZNR2RgiDBQy9nC/aV8JQnxzSAD1gw1bCtdhnNAYRDUQAKcsAcTakMd
Wpl8P6ImvxXoVeZtuKM1FPvop0uBtq49ya1MzIzx7mFfNS4WVEU0PrZQZgrukyKj5D2b/JnhmQ6n
zqIX850Isci6iEZQ4GZ9210DgLuJXyc0d/pZMS7P7Lc0a7HrjTYUd3G9LOvmjpxdwLfPxUQsO9jc
6dRF/6ST8UQ3CWGWfRqaZbjS+9CPHkcAPtthiXk/a1BM44Trg4clKPQK74v+yTT85Zcngvxf1QJc
9nfLuqTz24cxlGUxoKL8sfqIRPFI/f4tgBFTRm4ob+P0RSTlCAHhv0n7ByCG1FLOh7odo4YQyKH7
+QjEFJOGZ5oegeq+YKH5rsl/ejlNfHwxIeby2Ii1KmCIGkACsK8eK47Hi28Cg4FG0ZYyLVKbpGP5
/z2AzZ8GN09sBN2xKhsaShVNbEu4Md+IlHQoaihWTp8dXDi3WfgfmubHVbhnynRYiY4usbaZcV7a
zLKH4dMowSnkpN9Y2lPWfHmTV0w7tHwF7prOOfHFTcb+us3R9bm8gLk5moZgNT+kwRPR6z3W5uBO
+JjhdcYWzRLP3n6SQDxi3gsl12BNey1p6LmfuSCWZffJmBO11U4vbLor0YxplftXDP6f48T2FzYu
SXyXvsmQTcoh2hMUxfwbW2Fpxsi1YYRQnzqj+IujYMb0saED0XcQYcwORiaQWULASvfaPCDa+JGr
+BRcU+U42iZsuxrw1eAL2XFPb1RkqGGPN43N/Tr88RK4KwdUJWi9bsUDa86ukHv43ZWn6zYe1N7S
tDChuiVx6ZYEHa0rChICJm4+qPhCF+qCK/QrhqEhEOSU+aP4KnSthZPaecW6AIIKg+xvHscm0a42
jdHeeWeap55l9O8UZcTD6vLA4SDGhhwgZPs1hBi0LK6bzJ4TtZwwVUEKdFl+m6ef8wfyFaUVkXhl
OdGw4rYDXSAZ7SgbPlEaWFYX6d4LpdMI16kp+EX+ocaAb/rrGvPB0F8+cumBBp/MGTkBlaRIZIRf
j2EzwIoP68wGf0tQMCkihXTCIgH9US5G1FQfRhL15cY+qDMrRPqMZ8yT9/FeSQcvso/5wc9JvcLt
QUtnAQt1gflGMy9W3XyffpMJjLycabb5VpgXXN9x7OQEbzxJHpLfyw/LOxgBPfPJ4foEk9Y6vwX6
HS1aO9hFZaG+83r8GCUf4W5t/A1jM6OX52RLHTDmBO6tSNMrbupoQofXT9DqOLF4wDec2iTPJvwO
+dTp32mI69e37MzqPSnTySGefErmapTd5cg+KX2eWT8a0KdOes4W0zFMHNDcHYhn04mdtUdcFCwg
pgeqJL5/IFJ7O9TXxQrURWjQRPHvf0rmo+VPYQBZPS0r/PBzzkc5Jy/VOwHdkjFRBHrJE9Pv5g3d
G+HfCywNTPIO9vP+ISJAOdQCi/fZdw3ZbzS4II/C+rWQWtFKgskRtMBUV20OfjPQ048WHJJvS7sq
XZP9L63MOKBu5JKZu+ZIKq0NfNmkHWanv7x75JNIhaSMsMfxw+QWBkhZwRBybQaq71c/VGhyqIZO
AxNBQES7fUbzFudJik3xRH2WhPD/7QG1Z3rQHWt7gh7ugHTzflEptuvBVzufVT2/50dgO2GXQDkv
Rv59ntB9JxexRC0/2R7ZPRBz9fRZVdC2G6OBGJWnVxF7NJ/gVul0SEZCN5zEEJ9bxZG3a5amF+pf
KCRjqM5+odOxX1cXQtDOed+in2FdeDIe9BX4AGG1IOSFqj6O3lW8AytDIhBsikAVlRwvXPuiW/PC
rktCpxp10nZFjyJvRKxKHSCLki+HqvAWxVrl6lCBtulnDVG7i7X93VN+MPfSAWKDUmLSbggy5PWc
gWkpK7bHSIP6fvQo5uLpvpi3f+5Uiz6PCSFCVQLAAVuGhB1yxQolMAnJ71XkCmrr/11sbs24Fy0A
SO0duaV0aFt6jt5qfSemz/nQ1F2IJHPd20ghAU1HXTZZ1gyNO6MOwJlCgEvQYJhXPj10Kq0NOk/E
4zWI00L3Wx/ujXqTXXAZ3bW2QA74D0vD2pKb1N7ZpbaCNcNdhjAPlsZ5rKwocZf3879tqzPgrWz3
fHPLbjfZc8PWuf9XOUZnXE1uluhVt60i45rIFZv4jalGOv85nWp7MfvhEu4C+DuR04mG8aoNCoBp
zk0YOpKHYsKBL9L9NIhse5uQj40JFLsOIbH8KuO4CRFh2+LeWn4vcN6LL61ymKSJhBlp2BSahOUr
6muOXydSqZm1RxeCIS6sxP9i1ecYmOe1t8Mer5soQFwYRU+dbAtQNWsPryarodPDxZZcEYhHuaU/
0TqueIFkc8lGSnGjYUan+jxu5hTqn4lSpVv4AlCiqSeOw90Amck6XN0n9XXl9vPIi2GyO0DfEiM/
jdAXusZN0x2bq3AlkXqximnAxAA/HM4SBDKBUDzPHKlXtPGuSHO7XB0sZDhWhwz3cn6dL9TQCrnc
u0WxyMBdlPyhyEIqxiH1awX6Fg1zZwULu4rcvNpdOmtPWCMdL+2AVHs1yONRclIKalZbviV7827R
emXmVHT8ttiyzY1TFe+blZmDoGZrXLrFwR+NuiMuhs4mOMrxwP3ks5tBg8wZwm3yI2SShmNHzkpy
jUm/ZoCuGMnwvyoUoRdXSTuzmj2VFaVXoE6uMMWtOaVvh2aW9aS1GXB75N6wba1JvOhgeLD/qg/e
DWnL8Iw3cMXvBydtJ706CiJoFOTtU83to6vrl5yZvcNJpll9isZxE8mTHqh7uQXESxbim93ZzSDC
9eK1ItQ0hBJa75HZT4rFaTbN29rT7Hn9u69eleskZ0PUuv4/0T9lSHd9ND4NdSRdJ5TZsGpssPs/
qcd1qZb9ukZEKwLY1TtO3C+xnYssi4+6DfokSwsRm3MFjVHrYTdYuEq2ZaRqpsIymrz7xIKFXP3z
o/7npSn8b6G59n4qXEFGfLUE9bkdrhxfEj5nYQh5cQXgaIV8kFr2sEIOIKxDQOh6lvySej4/JJ/+
PyufZ5hkhyNkj8yeHc8CQjYWlBatXRkmXc5SKp2YUwq09I7nasI8X68BILpX/WO3q2xxmW7e4gPw
8Jlt0RvqlWXljH1npQBrZlHBN9gxXO+bTdeq18YWa0p3DIer99DdLBV/061xykuwt50gMQkdqieW
r8KWhVn+lFdnd+2QbvHhDjcZpqjFL/PEbyM4ELRFdqsGQ4UznKMpSalPcYF8iGxRy0ZjfDEXYpmV
chCt68ub/ci8+f/CaDKNmkPxTnurh0yfzEe0Y81NmTA/QfwKOosC2UYjt/p7zi186RGzGNFp6Wwa
KPQRgQC3mvEeAFJ3HbxIYNzC21qRlI6yQcDvNZ3abgDlZP/mGyahWJN2vwC19v8GiYKoWk/bC1Da
fQgiffwqYYSSi3aE+4YzisgMGNWC6hEb2mA28Ax0d07wksU5mjK3vHFNK0giq+rlTtMhrzVQTd2q
DYXvADFLVBGteULN7AhDHASZpaFWhgWADe96ttjoEN3C+MevEz4ae3SXf/Y06ShzzA2bsXwkZCZP
7eZ4NNM8dr2Id/uIwgcIGvWgcGYnUvYT2KJBE5ucNguUwjnCygY26wk3YWUzBiNODC3Rm5sD3DeK
CUYMtWH9aMYtEvS62iTUu9+CYtyPuXFnyP3wonPtCRDFqSWlAvwTPIa+1zvHfYhmFsMpnfkTa7/c
9dyAeg2X1ivp3XRwHIsUe/x5358wRWAWtC7lC+2fEGr2PGgse8gNbPyflqcqGoKmpcEfjXrN9yc8
R3TmXGzuWMYNlJXCDDEz4e4QDXSVGEewvfSLkKFkfE7lQrYBVjUmBR4lfrvhNBufRn90H9XacFOv
VI8GZUESA0W47pp+C2uqo8GfAnPG+2pcTkePS+wac73bTDiLYs8ZrrKizy+2a7746pz1Y8Yu5UFb
FBtYhb2WwxnsZ0D93qPuv14yOt/Vzza7ZBomEJJgQp7jtGMl3ocPHN1V2pS75exbvDP38mEBoC17
rYpFqZOwDJs/GaXaLcaf9O1N4H5/hU8GB+ztdl6FR26Jg0hfvQe3Ei/shfwOuU9KFenzOk6Iiw6B
HWhdcjHn34dWWo2CbeaF/PoSlOPw+ObFcGQSj8T+yo4R46BaBMik7vgqkOumfzh1YnQ3cG9JgLQ5
xKLVhh+P63l4K0ExoffKeEGw8gNP2BI6uzpfhZg90uCRPm7gQ1xccllJRyWzL0CcaUms8dS+Nell
/o7b0Ie8+w5Xn654JVcFazNN1nruXb+NosKJTXT8eAqvPLhqWdiTXHlBzYBfPIGejDyIsEnpRKBj
iAwMVl1zek1UneBPqiRzbN4901uvYrEX7EB/hSiENPjDJ7lwm2WV2NOmtRTs8FNA6iNHfO+WHJOv
83ybPFfullh9rSac1Fzhpk4veOIY9unXz/jol54OhT9yiDQMeVXKCnlc1Rv+kJB7oPYNdPN5W8B8
o0l644bMFtCs82/4wXrRICSnb+vTR3ronagobPt5P62nC5gI9KO0cLC/2fmNTHtQzeRZDfGGPg/+
x3Jro0l3+N+hqu3GmbmKH7jBwYP2MxgioNRp4AXeuFFrth38OkFiG1wEXrW4v+lK4/0MH2veo5q7
ar7Jy6o/9sCFashkH6dNpcE03+vHb6+bKhYxTtWpCA2SxmPCAjYxM8VbE3zmsTjqQX+oS/xnBnVG
lnfzFHmsYILhwP3enAecWz0cv4pO4ojD0D+4KcCH5PCQHAH1Fkge2gOJWFHTrhQYBrdoZFhzmYfb
2IWcs+nC1FSSkKyeu2dZGjJucX2Iela1qO+SO1Se9kuWaNtqmVCALsjqDKJu5Qgl9vDwMJcVbVtP
RV2bOjvYjVrN+c9R4hg0OebeIIOntku+7/tALDNvfkodm62iIWfbMHu8OAMagG0EgwlTKyEzLtK6
AqV6NczfCbOeEWiTIRg6M9gdTxIK9+zv6ER9t5Da8HpwObgNqk6YN9Gr5ZqaXm7xbh6XjerP1CjO
Tv7ArWjSWKIcSrP8F5rNxTp+0IWQNFGnHNSaLbsFcSZZZUqhYwG0sX98z79l9KrWQXAYJEPL7wxh
2TYvdbkG0fWDqogC2AWMV9piklJrOegyT88Kzd91eZNXMPVB9W/ds4FqlKtXmkhYk4pGYgeZ06t6
ksKwNedYrOln/3KRqE3X68U8U0Y3OkmGO4OSse7VV3k5cjBYkgz/qrBVkxE9JolQcxiaQ+Io+T9D
OKIIA/2OLOG5zCsRUHT2dRn3CU0R+OV0fINWD82A/rsHR0EH4shKNVDCW4iVMqthQUTE0p31sAa9
REbtAkmbtmZJPB8FkiUX3KxxrSHI3qwCF+oHy5O4IVyzAJD4jjjvt5bWg2RT7IZF+bqxkimWbFMV
P0VGTHa6n/Ft+VXtF5kKbqlTkPgV12uZjRFJOrWmdB8tsm03tOQfUZk2TPqmq76z2Pe1EB2JOcrz
gQuBhUBzBylUXM5qRDpVc5Q6Ae9DHL6eoI/Kes4lCCEcpuPtrTugMFICi34scX/7WzNe2f5T5T3L
ZEDX0/5wKeeEb9sfdXMMzjCh3KSvR3VC5PiCkq0YEpB+trItILgexdl1R1xueYKn1jHHl8rOiOjn
CHgJlXASXqXPysutVHtO8EdQZNnAnOsi7yxQAvu5RjJwivaQA7g/076Z2gjaxQmxJeIAFAk2LzCl
7yJSGd9NQzXO/Z88sjO2E50AaE92f8HwcOnYWqzl3ZAaTK3Ef/VXSLdKoQKi55DFMUMfUpWsI8uO
OvX8Kr8h8KV+AnJ9ZLAsTxhodYsaLUs1lxsFa9MvgNVVrxemo2DihaQ2D7s8eDAWdTq+N1mE9mAJ
MJL39wxXJ3wo3xutxS9jGFzniHrqC3LgDh4tGZviBXBztN+462u4FQa/RNRzGPTF0x3SdnxG6zKF
WKftIy+wLxfJBXuWytgVXBxfb22HsXRx+kYbWS/LmA6UYls6JRN7lvmZH6HDMHyB55erjjwLtClB
GYJoWdqesVV5bYnH8Yhyovmxzx1/sJwsYZQGcqqOYi8S8iqjJULFMqA2W8lhBJe8nBWC6tKMcA7P
1LOq73UxIv6+d3kEohoEtDIzWZ762mZ+MRUUSHNhQoZ80Gk3x85HP6cM5yEZwJ5YTlkoppPAH0Rd
TPVnIIi4d26F33DRM5PVN7F8udh2Gv+4vdIYfiFwOO5+zv+mZyrH5dMOnTxfa7tznCUSIy/2u7kD
R4QY1isePQKK8wwQSa6UdSASYPUDllGLc2BNRVzu5EqI4+Sxyyk9j+WIl+8zoh8U3x7Itbki38mK
N17uUeYmT5z6IvE+VJUL0c4c4qK36K+PkqXbXKwKnsHsAKGAHV98QxEFMkZUlDFWvlCc1fZaIC6J
BfIdfZNUPKJEXISNisgqqYXqzBT1aoPURgOg7xh22Xqu7GfgrTdugprR7PiLKumag1+0fIkkgeqC
SWvclaySzWfcq14R2RZbc4xaFCB4FzQ9RPDlX60vfAPTxeejOVe7lvjHkQjNXRvaXcPJXuVWnwvj
yZJd0/u0QSlVNnACZTiQg88AovEZTS7kO9U90v/IZBIRdvzCnu7RhzXEVe5Var+laiyUU5KXSjxL
9QMoqm73ktw36VkUHwfxsvpoGIjGxcW6+lj3fkbZfU6RtoIbo6W+YM/xAU8dscOw1lkayIX0rdqT
EU/lOmecR5EPZuOCYQe6S5qgxNtmSRWOFV03EAOzIRdTjHDriW40svqSick7abud/op/K0IDUKzq
b/YBF1K7/gI1mLBlBkNEKSfG8Sa7BGyjyj1p0wEzFUaeqgK2zfCq3BMlGSZNt+Omj4aTnK9dOcOz
K/JIta/oPFBxWyyZdvTJVfskCmyfieFF4+LDoBaLeAIfFCrYME2zSGaw7BfwmJYKeZp0bzM014Ol
V6jJh1nbQxYPTxsFZ0uncqV3nvEbFrBbyFOi8NYjwWsJYQqN254qbjallHR9iRbY5viNCXvFlm69
gIBgFYVm6TB4kGgTK/7EVhqvUrqRacdZYpZZ/0JbBW5OYLRq4y79EboHBkPv7MOafbQM9AJVH78V
BPPIT2LvuaE99p4CvvvNGfr31WxVAgTDhSXIdhEP6I/ZUbjwWg4AUdd7KgqJDPg2iutEMI3YDa+n
D2AnjxxNJjjwXwQG3DQnD+dztin/NIQcZeZ3NxmkXNIv3iEpa6BBWzkJCWUVF+Sd/Vdt0KgoJrM7
Np2O1bsZ72f93qZ8y5gBfjJIzAwJrDG1hVvEQ7KqwtMyF/d2aJAv6JEXXtJwsvIbyQbqnPt0vg0r
DjqPh9n4XmfvQuq3ZcnBm2GtfS2EvHogmNwqtLIr3zKepRVliNZnAAFGAuaSXGtoRK8NYh74yijg
BA28O3+7NBvEgEGhEp6Dc197M5Og6ecilYqnkJpK0chUmsRQiQQgRH6XBUr92btkrcK1R1ZGFxm5
lOYV+EL+lx/+kOVrgXd89y9m22SHEoAVPz3olhKE+6YILy+xfqAxUIwFhM1z8BQb7sNlWgQOH7x1
8wEki/tzRKKp2VUmgP0jSEmeMYEh0xeVLiOvEZSgAXF5aFOq5vHCQRhl3FbVWNUmtNk+U3+cp7Ux
Oz+48QIwHxu7oHSog+HmCATJ3W0Yfpu0YUUmPUxfSzdppUNlpH1GOV44FOsqd6Wm5DCGEgQ6kLPU
JpadNwdESxej4tptddmbNp5N4lC540dgdLkK9/n5aCkJznBlGJaVxP+HIHwmbJ0+N6Ys4VianLnC
4kcwucv8tiEe9+OzrUYk0aCje2MogQ4iSY9fouWv1a7MqsggTNhslygpW2/buL2z3p6sTHbEyYw3
iEyaxhd5CWRYVLxVc93L5GwegfnFn9Es0f95iHlnLItzHaD17wEdUtR9eBZI1o28hZH4t2HlZPb/
MmZRhnL0tMal0l4iMOocwQtXD27EnSs/Z+Mv7m2irQ1SesmtzUOZktujEmts04gv3LqCSB2Gbq3p
iD+T+Ll9+2G7hv188F6lFq96UYagTnbjxTx1/xiuYZBjPzVNiYPs5uAwx+6YwqD4cvYSue41cA0K
CNmGuWZsQt8hqE4NalLl+FK77b0s32W6yhpFESzGrzSakrW/20dae/nbOIP1k3Go8Djy4Ca3rBOW
37OfC94X/N+0ijabEjtWSyil4wv1igj4Gn/ANrRuSmNQ77nIUmuzGWwl8EcF/avpqOQhCDQdfMW1
/VCARq/fVobWEPbGHyfmAoumdGGqP/Z+Tt76Lz+7y10F2ZfFR8VYHMBe8zTJFuWIetvq5qU7EPf0
6w8RydeuL/+VMS0w4YA1uvKecY0iBI+v6RNOnBvCh/O7qt+BtEEScm6IgECxlZwBoyx0jSCJVa4A
tdnifhAHfxqvmgxAgYVFkgqqTs81iGxv3Mr2N+yMMgcmU/9GWSg6MyjuVufmy4uWpSuP6mvyE8Oe
HPNWzvCu7sK//DXXcdCV3oVdOrLJS9QyLUquaryFytUwJBeml9B8furfETNonS2D94A5f2Rf5891
5QMWonSQqmINtX7lwryBJKCYJ/x9A0rVlZqn/ALrsYT/t3Y/Z0VT6oqKCVTxC966pM3piYZlcc+i
49slVUgSKaYIgNYEQd7CElhBB2RH7Jn+ZiUG4pnNlg8t48mx31v+8XARoAWy3Eypi3zGugE/vJ7p
NIfM/jquLgywC6urVMFrvU0Qt6rylL24MHDEBqUnIgfK3GrjvvLyVf8Sg367hmOOLWtnvqtNgn+9
Bbj8N6oXDbfKD8+HKxRyKVeZ2O0e+rSP67CCtmkoanJLji8QgB04qoD+hU3P6gwdd2RUAWM4EW7W
7HyZO8QQNHUVttanAcBBPe2ixQ+BnuXlzpQHhSiFXdSP0denD78Tw10yNNq11CKoOu0JzAK3+CpO
M0A0r0aNqLyTtr2QfpTywU2LxR0O3ZY18YfLzTFiVmGazXJIHQ4eTgG9kKSjeyXRIVRvluhog8cO
Pe4HrAl/xng7Ymr/xTSfBt2staycY0QYug/7mp+gZwCCdD5xyXYsyUVCAOkERATSc0isTXfOl76E
uNu+tzRu37QQW/4iB+JC7DHlW1Fpa/XHrOehkxGhuWjCFmRYqVQVqX2xGUbH8K43i4RCTCNm2CJJ
T1iGdp20edTFYk8lEwnNS6M59ZTWvaTZUc1Db1z6whoGWBKU185ajIxy2il8c6geVP8d5QrgK0Dc
pLLDHrUtuhxPOWNrIAHsUm3zbCzPf0YzoSThs4WuDAQuDOb6Ae58P6MDjouUmXGsYK1s21EqhnHP
YlHpuTNYow2dmV2Lw8RTZ+TNHTkabTGFt0zx1Y0yzr817RA5uiBRs3iqPiJ2a/FF+PR6Cwkjt0MA
lpWXEwg5P6/OtOoK9F/Ck/10Dpib+scuep1m3zYJAr1DSXT9/3AMi/61+MiYqTKFgs3gjGbz5cJN
MUhXA6UOYCn0UFOXqFGWd27MK3L/VcziCfo1Fa489OYhe3lofq/PItqItlKlDLKA+uIWms/9F+K2
CYZ/o4QRsI5xQeqJwD/gkwsr6cNnRyQhr+EqVaqZcyoBqO8Sn23BRxYvVLCwZNEWmC5lqmIQMgRn
cxl1450LW7V0+y/H4Fy95mGx1BsY4AYFe7K9S+Z1uOz4M1gdnnA6Mn58z+mq5f78Ueo0mnJGsDx3
HvH1K+m+To9+CPknXAJYeRIOj8JHwtnhMHFeJbTM3s5NdB8+4sfIWtvhDwTF7Mt33NvLDsy8af0U
mILHCVRWonxR52NijKgjqFosD10iQEb+wjbdZ5Dl+4gwSEl7rSzMFgs8xRCGYwCO+VYGxz2bUVJJ
bjdNB3nKS2t50Kz37cPa68IfFsItZKA7sHoObL3BJ1qS/zVWedGiomR0Z+pTSKAc5so7qGU64DKQ
8+3LjZ0Lsy610H6CduoXx7hWHG3REmsoeonma6Taqf8ye5ToHHeiZ/jHhQaRA8DtLlUZ4CA+3JSN
FGpLDnJYKSgWOdTMRC6k5WYYOtx9YxmN6HMDa+lIcx4xgTNTH5F6SmecfUcADUM/YIzu9aahYSXE
HAkIQAInUOzv4N7CCIX6IVOh7H0EPV+IGcPn3MYLYknQHrYPnm/H6W4IbzUPtnfzedgDSfYZUqLu
RulDkVB9hhyhV+CgGbXzRVUSpO9ewec3/mjtI7eDFzXd75GeDgDlUEgozYyuRUsJwZ8KyXJFxU9t
hWgZS1mcmbGcytO9H3nQbSSjY8GeMOXkP4x43cDIeXf5bYVCHQ9wM47YQQG8t2o17sKePBjbV2Wl
4pRlP6x9GfdMLSkPBIdmIaFZTSmHBQ4JFu5kQg+Xg+RcMUGlG/EDKYp9RZ30B/4Yp+Jlihm9f55h
au/JmZo04eGr1fM9iNk0PA3GpcYCGs1MMpDcpCUvpfnq/Bi4u3SgV9g6ojnAnUc/3fFjEFo02sTM
tsP5ZtxGb8enh/qm6+3Sz6UMg6UmgL4Pa22eoo57x9M6JOfhiWNksAwz4kPwIzCMMkHZKRZLymwc
4pbQ18fPZtjuLsFjfn2EqzIxOcDoRtTYvbXyH+RwMsSf53rHmX4p1eX9kLecM4nhMgbqyjuoMdME
2fjX3QH0gfPnxLx0QjeNE5ZwR+LTxwPtiGsGU4+H62rgjNkbhIVzAHI5I2329M6bdCvfq8VASNtU
MkxIyJ0c7ZtWz4+EP9I1p82ySh2QWxtvxwFxxZM2bJ7Lk9We2YP/fF07TCsOHn47Vvae9GLY2Mh3
GpZzsL+7JTWDH/QVH1rvYCz3khfDG1TSHNtzr6GVtC/jW0/CiJSsDtWnCwrZN8RXyxF4X6kSY34B
x3yDLiBaiLQzBu/j7BDnOzlH/VRWN7WpVn4NkXVKq7nAfgf2nGCXugcKO8PiC3upktrMuefkzO/U
7HmJEcqsu3Eq6An9EmDS0c0ZCR4NDI5bMEMO18UIcfI8ac7xTWmDC2j1gOkvf+aOZUYjNcKmg6NC
g+s6WAIxi970RyeJaFPOdG/NJv1qrfbo818Nj8B6996UQInn6H/dOjAtptLL3w+YpU1sHKZQAtSr
qpRDJkmfnAJCmRnfu8jRFqYn2lMfjZLiPyk7l07VYzKIu177y/vRuwz4KIQVSWmxD/ae+R039U0I
BuQTO1xW3gBq8Lbc6kZsm1Dgwu++kaluZlbV8QtcTP/KcLS1DyUsquo1hsZpmU+zP5Na22WSkTWU
FBltJd+DSjsTbdc2y8mpD1mA8EtlAdxfTK0F0MfjSCok+AOAArLOObYm1YxH6NX+xiq+evnyBQDZ
eSuQKuKullws6WCBrVZFzWleKK8NzQBRisbS5skVBby0mdLjl2CjOu4AD3z/a9R+/KZDSFhp
`protect end_protected
