--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
ktM7BYSUNDIoCP4iXzZ+jJlwxH2eO/Odaux98RPbBkLuwzEY8utVHL7X7MEhlTFo3rs9659X0TbF
uNpHboHjbb9WUzozH9vw88zt//GEOu6/8duDFuNLbLl8q3zkKK0YFy4FjnZL+gPSm/kPfkbVBlQA
AlTKhDnkw34qTYhIlfK86Xgmn0+Gv7ryHb0XI/Fdrgdi4FMAM0PdJ/BdlEvnZJLiSIl/vHS+BMpk
7EisCqpsq6s8Btu/7+5mjv5s2ACZMN/VDTUgEDLOWRqKyh1REsWcJ02SJuBax9jndnhqNogJzVUp
/TnSI1G44sFpTSisSXlzHQKB/djiSUj+INVpJw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="5FwyDk4YiMxbWs0FC37QPDrsJ4t6LDbt/dQk/Rb6jgo="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
WvRhFN0d0Hx2zgLFoLeo4yTnlCyWKGAwt/LQFTNyfIIreqMiAWcSNVMnqvpp4FdVwfvcvlRCRv+f
KZq9SZ0NAOgmPPTt2kvGt7z/gMSxyoz4GwVbMvTCI0lkLMUzISqNVTOwh+tX0HJFTnxWsf7oAxQ3
ReyvzQRX81uVZJtWmbqMaSTpeBZNrMcBbaZimL+d8mRb4SuME3/LpyC/CTNKWPhxpWnySNw8xN5j
ShYZJ+KvyIF6pRqm5XI1/ML/aWJBr554Lk4CYlci56vpYIThkKe7fO3Ow4/ORw7ID38IwzAvxvhQ
VRFUTSH2bJ2H4OZszj3nqlfbTiSG6qDxyqtZ8A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="zk7a6Mk25ZjhLmQcy1NHDZoFPppPqH5hwpEZj0TNiQk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13888)
`protect data_block
n78JOQ5U92sfVeLdAMITwTBoQf5tDlI66aslTQPJRXKqAKkQr/hmoPFpR9kFuO6Om2KrCuP7OjKT
2q6IoQaICZH3j4jzyk4jYzxAuc+iXDcLVHNwPuBQAXQTha/Mlr6csWGm8+5nqWBC7vK4ShUAaHj8
u6+yF7vyORnPeoBVhxuowJJYTA/i/x0G3FfWiXnm60wm5xdHUoBLIJujI5dK4HaZs2YFPw1t9A+6
mfLiYwHl3uTFJedpy5aIfmuqGgVJVRI9MaTFKdMeNpW/3EcqWdi/RvcKy8ordc+zoWx72xuo8H+S
HhC1wkciL1khDumN/N1sghP8iXJzB6V63A72NMsIm6FSS1CNpJWjAXEaUSZLA22+5k06HEflVctA
MVQNd6p102754UZ6iTJtL3xK2ave8q3X3mFPUR9LzTkRjlgtfFe5kcGjLc4NDbUD0VpVPScjmkd4
yl9/ZyBMcJ0OIRhJp7/JYWMf9qlMHqrFFQUga9oMM5Ri+2XT09UaPBte+lWx0VB+PGMnDzrSHVp5
QH7geTMpm07qwrbqZcmVf1ILfo0gFJAXffD4SIVGZO+eIizNsYstr2CHc57AImNOFZJm4RV9ro8m
lygzdg5Urx31o6mwrzbKo9S+f5mKU9um+ELNJ70aPLwY0MfXL4ZBKEz3c3hnYn+4shnyFXkhFTho
KA2ts0QHsrPfcl+ZPb4HGd3scCVUbw+Fpch9xV7Kf+GhZnBFSaZI9FzzQFS9XuvPZIOjHK9F5ndm
UNDv2NCOf4QwEfB6rrASndE1BeoerTNJvcBjjiJDoOz536yx6bPAD3wyro09/MurX07yBH6EGb6u
aIoMNYCQQpOAeaydsYfh0ZqZ/Lot1kag9yKjJH3Un4wl8EjY1GAE7FgbYwTv4EzYIeSCyMCgI1UO
QcWCaYqHCk66GiYORnflfsOzuC3DZHAbDMLBHYarGQh4dUPvyKEWhWf0sGE3X//5fQsoJeSDEcSo
30FkdrCpnPXyVxkjU7hlmxYxpUOr2FfH/MVFbH1xNWqZA+LjC/lXVseb3QYGUS4UQTVtUW2V9GKi
qWtn7KkRpwzD+291FHJWDKax6/q7IwcqJglJXPOHN/xM0InwHbY9B5d8Z2RrB8l5ZxxzbfvZ6Gl+
3WSDS3Re+zlS2jAcH0aRnrsTgOVrCO2+wO9NJUIH3u7hmjrlyNMc0FZGSAreE4hpDNo6Qo+4UiyS
A+BuZfCDqjsSTYHINHF1jXZL9Zns7dwb86sSb0ntHvVwhLOojGKQx4UeK0KwfRnk53un+mdtGS1o
whp5VjEnDwMeD0rEP3fEQl5Xsz+LMmwM15W4FFwDTn9YmRkgpw8WUYN7cVUVMwm3D1bDW+zooYaW
saY3HYIAJ0jtf82AVr0++D3mao4WEgC8u7qir8XTtTQoP3r5HQrRHcauL/W1alKj4bbjfCmys0w6
HstIhDqmKkBrgehywgKT9Mn51CTuiXA5zYiHaaNoCFAyqj8YH63Nc+3RE7iFnVKixvo2p63StF3q
As8z8bOraSNdzQfCd4uHGSEoIG/z/YDoVBH8dCQtGugsdzwMX6XDxNqSTgaKMKzP6UNbLCNg5qxw
XOuRs9xCsN1JWRNLwZ/OQiSX8x43DrC93nBQL3B3sR3hhBofLeX1FmECZ7gG+kGhSPPS8F5CWsii
ldN41TZ/41Pp13msaqHXprxYuz9Ty6Wl9wK6xcwGHQ3ziyWbOykNjrEWFSccYMsyMFLr0oFSi4od
PbIOjCBJtWO3A/xBRwtI9HPPhgjP1VYx5LUabGIiu8D1lKrpy0mBBKacu/gWlbWUFilbJsRoLmeq
Zfyei5fo0vtpZ16C+q7D8Dn8QdL4PyCUzQe+g9w17DBiWKzCVpFViZBozeG+Y5llHwJvr/+v3i8k
08F6UDM1gEUOCMGFkuvA+CexH+kNXrTAclQEWV2y+bFVRpvvBO3nbeN5Om2lghe8uY2zNTIsflTF
HimLMT0ZgErTaLsyV7772YLza+CRgpiAxdBxsrxi00H5Zy5NGFhGtaLO+o4SgZ2SpAk93fW6udyc
OQEb2XO4zJ+Iz7773raAaygsjiuNysNdi3ywlkRspNzEVofQnVuim9gijH994BXCkIO30w7fSVlT
P/unQkEw5/H5x0bcJQsbiDPfPqmAkoUEqEoYCIkJTSNIPwyhIlubs0VqhBHtejMSmlrMGI/BDlRz
EIhCsVaqI3Vb2qitAQsgrbJNDb517DDMFtgRM7wFMmrk8XXKtT0eLCWzFIQpREntx5x2qq4GtYmx
AuwUS7h6DZmMvWpRplKiOBYgQbI6lqI/2RZzecB+5NHrMCqfC0OKhpuJHXHNal4zMrz3rARUr8uH
Mr4LMt4SAYezrHHKowCBX9ilnZxKSwnpSiHD0qoR56TS4AzMTiRziOYF7XiUBRXt1P89q0BFQTGL
TguXxGQg5k6V4i2NuBFeu/hINhq+UAKj2vwOu1KTQFRogJPtB7IQd2SVrHridvG1HV/Kq4Lr0klf
k/4gUDq17nrwlwvj9zGE1/ioe0EounwKsHxtAvbCJjg8rF/Mey6b+gHvzbPGU/TWM4OShcWwyGRy
A37UjxNgCPa/oHOZ+YMqY5wvZAWahGu6FKiXwWu2SW+kMKL4z4eq+XOoqvwH7iJKo8MtKtGBUo5d
9Tjx/JU1RoRc4arC4NcORUHM6QHbLnt3CiypjqUfreScUyiNAILUr1/+KaP/f9H1NrXZkH4Vx8hl
EDFtPyAvQloxDj83rIbDCcVjkza7ermyhV9ZYNP5+/J1VDIp3DsEapRXj2iXJyny2Y9OuxCx0CyQ
ZrB5Zo8UPPcpZzXOuqJeKKgB3pAoIGKklRaP5dgIaCEWpWl0SMS0xb7tVKS+vOnBrRBOMqLJFHUl
nuxv608QT9DijeFynJyHCJiBPVr+P7yEYrfKHSAMnThXI8VRoFGppzcWW4oKvWz3EDfCidpHaKkl
MwCeJtgw75+sYV2dNe3H4OEWWmS7rPxli0NU+JM7QjoL/CDOIwJLBsgTK3qjtjzMlY6v2hzdP+Di
X3i+MTC+Y5Mr273El+J3T3LKxWl/aS9yUjPyfTzhSIV53eh+ApUfKxiT8Kz+mWCVtr9RtRyOAcHm
kwsvhyzeKWfj7JNzy8GKBhEDxC5rd9fcsyHQx0cC3dYpOn2dcCEcW+f72FPWUXRymxQVt5u4npPw
C5NEoq5Ds+zEUEveQYRO/dI+ynmKeCHEiCqvWykUsLOPSrq/LBlxfMr3oH1Aibium29kfc/PVZ1T
WcaWPeR9vmybkWuTnH0hdRsGgwRnqk33dYpBp2Okmmb0kqbkMiC2FDmQ+i4qCr5ePBWyt1b6W11t
3OFVMHoKNdJGIdmMBYC/95YL6mJNf3ZlQbPsC7n5It8QPZ6FYldJ8OsY7Rq76nERS15EwnjDTjpb
DSuJhpR298WyQG6la862JAIYx+6L/IvNoOpnJCWL7xKeeTxizv2o4qnNfswmcgARZF7B4fPHdNxI
MqLcSuqXEE5t6Q0XKy3RuhVpd3RYKHPzJsaszmsmW3z9Jh/cTKeWI0v3Q3dxRMmmYm+L8casw/Yq
T4/0oB1nawk/xpLFzLSJ0EeL0apLRM3LZA029dt1ef+6urAajvWX06ZvI4CsCD4+5JHfXYTa/EBW
HWUgGVWWbrjCcjYnCWevz6fLHxNMoHX6BhrWA1sORFbypsMBI2BYsVIk6gjHtA+tQCQR5SUttlvb
x7gdaaahkPL36cXF+l7KGKzBW0GgaTG38l88cn+U6hUPZdgXUAxdpStS7JlPH6ml9QkZ231Qy9Et
Np5NbwNnp6GGFP//z7NhU4nk7VmzuS7oOW2wsVTVVPo0oFxEB156tSvw3/erQz5c5FIMn6A314aZ
vdVTBUB0QwZGQINALPv+aeLbh0hPZR1ZszjlRUZRtjtZkOveBitF3IkAioxSqqeoEnGUFxrHIwOM
s+UieVS/Oe1omjQzBC787foLIe7q3wnWUUx8T5BAtWvR37OHoFVKU6VBLCU2ZGB7HmLFw4PMqZYj
trFJSebZ3K3yqtUDhSR8a0Lai1+AT7+s3gMwQUTabMqWstICoTx8huiHFXlXYQk5UZdK7dSyyCdN
GwoEhiF+5r8Kv90IoXGFMnFNaOJeS35GrwXaLpwBUa1yN6dfnigZLf9OS6pEMkAhFx6jKVQvd9Uf
6LJTC7OG8ZLYYOQ29xZMVpjeo7AvTIYD7B+O9B3YREBcki+xIN9AjCZapJKwcOVb9I4/itEWQM+J
3KA0RLpGEtbyxqvIG7j168UEA/mQI/wsafl/AJhHucwk3+F8SkkEoDsAiBQ9XC8jvfJUfkP06bk+
LsW/KAfg0ZahqBN6wxWE/lxJTNygN5OkOnviYUbccNd41bV8Ha/s4TbsAo0YxDIkwTyDV8jMqx+L
qV2KU2agkmNZtG9lyEz2+936DF5GJ+EkrFB3vd6sAb6B9YFMOzBMzecySebpGH3lWKalNwxubVQj
KnnlV36X+vvPA5LXqwgbsQRVaiIFubI3lLkHvUDqKfGmz8DK172O8/tD7b5aOnupaA8ZdTp062Ia
4xzf6QPUUB4fpkFjtoVprqAQYINiaSQ+QLO7E9UBbqJtAm8VFqB8Ad6eBS4a01T/N3OQHEczeTsY
YTbYt/QtaoGL9NZkosb7wVzh8iWzXKqEdFCp2Vq1Bk1uZ1AXEtRrrIuTpLiZ9pWLx5SD2fG7cOwe
r0S6MGfKKJQLM6SxQt9hRqQW1s8aJJGcrJj8EKJzeocJ0z7b9JtcOoXXcEuKqfOYsW8CL5H9/ix+
I/deB6pu5iJaYUoaO/ka2EXi1M4++kMa/HF1rH//A8e4rHRV6XePaFVJbdAIkDWO4CgNsSO58lRl
79GYtoWBBfESVEvfgWHSMKJSPaaNYyZv5bP2juJiJp1rhXRtJlBey7Vc2hfln+/cCKe0NyI8f7hS
Xl0UbZMvPgOXt9f6JUM4zAhsc8zw66bDcLNZMl0hzYuTJMYzz4BOmc1aIDVnZ6azba4Nw8OMY93A
bHLfkqEpZa2RnMjU2xEDqdTN/LlWZmitC1vSkBi4+6me0Xew5hjwMeoZwdoSKjJd2awjhte5Thof
7vGUzlgcxQg5V7l6DizqJoEu9tq6om587qLFF6g3y2YwJBSCH+yML1BpHQuK9Wb7Npl4vQP1UlEX
USPq81iR5L4z03O1CoaN+jU6jZB0facvHn2+vemWAxI1ZJLFlvxDeskd3MK+VfPkgViiPHD5m5AP
mmZJlj2URSHsm1ZNxj1ipw0GWbMKOoeDreu2MeBGTlJMP2oL5cPqVSzoADMcLxTfnlTiCSu29qd/
g/yS8opESlVIQ5tNw9zqnKGRtvBv9h9D3c9uwwKhgNExgNudcY+4Dw8T6Mb7E4jkHpL51Zpr1cEY
XbVbCeU7L6EcfrqRBOAOPUp6duNhy6ZnG5s0Xm5euu7yXGP7DVSfQjAjSzFHGhXOMOJOgfge7K6G
6OV796/IMZGav9ioSATZbqgm8YjUVhU/poTJiSVMieuDO5UDXidAjG7bAZon+Iz78maltNDyk9q1
OyPNHJSBqQ3Ibz5S+Mg742MH6mLwO/LuV3leCg3zv7yxbeEc51ygW9yd4UXSXBelXIRtQt/Hhy90
c2RtB3AUaQZIBeiqOQL1H7zVojBLQvbbWXNov1iEHBRwHaa8n5WIoZ+YIIunkLA0832lhOmF+bJ9
NQVwe8Ot784mVqI1eK77tySGSBqeRdT28dBmYNoUEvFyN0AasOW1+ZmydPakAWJ8cGqMhiWOB949
FV8oSiO9ajAC+yA8Q+TObNuVE4Hkauor1J+wu+dlIHBVdZBVnAtaXlMyMmYW/nlSSMVhDouCh3VA
2bR/mubNMEs9FpqD6UX3TBG5YoZ+4nwkVM1lNEgNjqyZ3rwfDrtAO92hfIqwCQoG8tUy0Sdzn12Q
0U9WOziiY69UOgUcGTPJUFUuEpmueoNZWraCXvhI8YhwGCbF4+on+K+VhtrnkpNPaKQNOZTlWYuz
yGazMaBn8QxmQRfc3STtbhov5z6/LMaGvczGtV4wBcaJEeK9CTQMIK9AJSBizaulJkoHlahTiha/
hPMlQ/7sfqQwt2m6MdfQvwWXE1IrLEW7AblFj0UYXeMxUxCVQzH210DrluJP37bGcI3bP25YKr1r
imZlKWAfi0tN1txqh9VwUdOM7l7oeFTBplKPD1s3TyLTb3eOW0AwtcARbFnsvAOIYjl1N6fJgedd
az1CjLu85ArOZ7QL5+a6m6vhXrfeC+yttoDRbzS1NjIT+iLT4FcEuro+O/v/Lru/V+Kn2Ol4CTfw
Zs8AqoKKzxf8Yv/3VR+q0iW3pi16iytosCYIXtrnuK+wNJF6AI88vmaTQ1jGgGnKH4uRBfQdIWOb
JpT2l1A7UslQ4G8lz02XGB3Yp41YJ7em0Eon1y9cF2MtELBtjWcQfEzAZcN5fkZUNlikqsiheAuV
Do0InMArXumZKyF79Xv/BpZ4PEUhLuc3Dr/K7Fe5QtXIioQr4Z/Yt1/boyJ+3bnp/FyEtlbM3Nz6
weqgfU+PJoVfXnd9FsK1iNx1dUiI/5db8IOgk7MHsCuFX8SkYPGw1B/IPtmYuW7I9ZWZtXR2fOns
Rp7aHrTjr0XPDO37/SfaBaML6AvY0rF2T7rSvYzwCIE9DfiVoHETSKWTBnkO2xZrpzhD8rEOnDYc
hVLEoXgqK6EBUaSIslNEBG2QfMYufQ7XvqUsG0tybayl4ibBPOu2ik86Gm37nxCxgCRiXfLBM7Wi
KkDdHudgSFl4aTtHHAD0GMIrnZmZFp72y/ahaorItJTbwkVwlMKtTlUi94V0jABUOqQWJvVszLCV
vrmyKkmCoSc0E/EIKOCYGugDk0RWbVZ6skhtnSsb0PxL3ZwOP4JVjsCp9Lm3izhrNofT4qRVK/b1
AzpJiC9sw4Od/SurVsGSQGM/eap0KM/uCPW6Ks7b93riq1Bk3Yy2NERvpabBWPsM1JaTmdT/l7tn
oEHu2y/sY4tXN2HUbzwBZhXL8mGZ8Qw0OYFGg3pdsGh4OLaCVOwOYghAjQELZRNvqW+cRtPgQjuf
8R1q0AO1BqePWFxNeMclOMnFDt7CKxKM2HlmsXUgY9uInWdxdXKTuiZ9sHua33zzDeWFphUQk/ma
JNdlZMCnJO+G5TjqCJbT8g5bfVxQmTH6w0C9TXiugQjiN7h10wxI3Sk6UuT0wu94Yp7X7j2il8cy
55QaIsBfpY5QOcDH9iXxYKzF2PAEPHMHpHSTwRJHq46mFjEzx2SiyYfaRPw7RT0NdXj0hEFDMo/P
U3cpDZ/t8Z98hGU13Td9HGDlyDMv70PxMGq7mX93UDrsG5QWtUB3YVGAnaPF3UwugQC0L01imFom
hzE/7Vu4ex/fAf/ETwFeiSanvV+FH7Raxtzyv0DY4lWmcNvLfg+hQaJ1+hcq6Kze6AomAfWL6oW6
ZXIOM9uMjLBr5rpkkBD2Q5ToCDouJ+L6q/+U3yDt10w6EqJIFwDfgBBCMkBeVghKlVXyDpzSG1Dp
Wj1Dh4UVUkKy3eV+4JC2yFCI4TfWty6VvgEmyrc07JmeympxRYVkZydKIx00ezjoUWJEtK21rZe5
KzNDg482Pne3Bc4vRt7r+OW7LfBZrgWmcU2o2nKahSutFQXfFYEfFdj8OQN/kxHnYZeqQqXWXsLP
fEXOoQsn3VC6N5K149COkoUJNmxywgOF4/ePRaaveApk9xqAsMz9SiIZG6NhNZZtD/7UHybmeoLm
U4kCqgFizle9oWpL2AWIOVYvXuf9g00dleyAWPq0tDulWEDaNfjPEXTVHtKHo0Jsgu2Po1NXk2G4
8ujYqDyEtrV/v4bZ2m9tipIAm+D6lWRqUw0PPZ1YpZefEKeE5q+E17vmMgSkOn41XwZAszDAkBna
9zz+TsH/fKOQtMLw2DAkXGs2JJUWzEj1ITAvwO92k65Ve2ewc/Lda0FVKUEH31dCqQbcFyBn2rms
HmR227HPJPCQRfnH8Ydscy9tSRW3xmz6sWJceEduSjVD4MQEs2isx/y3T5SLWoAiqV1/o2nMbcFI
rOqtxsJmngs/jQ8hEtn5RSSHdkgbzfiUa2sphjiVA4ARcR5k9/sLa+RJVfOzgMGeRT4wEe72t+jY
hZaZYDJK0v+m3W1LLd78I/rZB/x/1OkziDEfbofl5uHA/CxO/HVrzrE6dF6ADW2gTgiT5Qf83xKa
X8yTVV3wh6oIghky5vdAfRFDPl17lEZvw1d1G+b2reuRWExKq9UmAJCi2mm9aYN+NCSkJQcTiCh/
yEETq83Tdi48nhtZ1L+Zu44M6bhU/vTt6trmQp/Lw23xe+IpUTefI1Nghn2PzTBRH1MhexRnFq2w
jpljHnsmGLZT3rcUX7fO+qrnw2oYebyL2Ukf5sdVvVBz4PPcL0q17LZ/iHUv2JvFqlr+4X69Bfbd
zOLDsspTEZN8uRhFhCuLHgyv5ft6gzKm0Je0O4U5Nl9ZV+upGO8bIOK+mE2xBG6WDMEW+ALq82/h
T+h/oZAwPJ6iph1hhhaDisZKYKwj9wy6Hc6NzeC0zZ0vznpZleGzBjlAUclB4KlEEUb4J2sZhV0k
9tUVXPa0/aUCWOGzm+1+CK1zd2da1lHjerXCRa6fEGyf0cBVNoWvW/WgdY1SRRLLy+3dnkKt0O/w
LwuwrcJvEWC4IG53n6qS1Di8vADQlYMnV2PujT6S6RwZs9AKSGKIFcOyco6SRsVqR3suLCELxV1W
2gaOUxKIU+4xCWDvXeuDhU79Y2F9OONSpjNYb/3qRMSwiMdkqaVq6IGiqpxoLooY33JjYIv3uo91
itZ3a6I57YQDOV/oF/hwxoPfMTqGoZoz0YxX3vg5U+nh3U5yeHQxJBkppJBsz7ORrJxW39foXay6
SDF1nrFUR9feU+Z+PNOCwPePkCtFsTnOidRbN5WfN+lo1ZQ822O/XZEM2bPQvQfkoLQetB03dI5S
4tVImCTCEYthSZl9fqIhZpDRipwJ5CdFDFeVdZXROdyI4Ev1y9R4JbxGVlXVfeyT+PRySw5Y7TCf
bTWV+ZiRBjxkzewZjf3x0vQgR7lr2W2c5sv3ZC+tVEaH3JUSYzp463uY+5gR0UQiyQHdllfHk3q5
rWlCHmnEcL2HpI1lUDkFIUkgxU2fynR4nWMsEebn9hmzrT6lz2vvlSZBsO/zXnM491J7O/2gRAQ3
YLVoxi79B/I4Tzy/fmOWWQOeESX1S2M40692LLI/HabzlwlqykvFFCxH2DDjbXlI8gbEg73d7hTK
0pE0AamrpDYZiN9oPEwFC4ecPjfd2BCwgLak8C26T4w9I8wyEwSG845mHwCBCBXTw3jz88gG99om
4hCOFTcLllJRFa7Ua9ubR1Rf+gfJ6QRc1PiJRiPGSaLA2VvLK5I4AiLGj7d98FP7IKS2TtR6PmK9
zLGX5oLTwIWVNCsNU4Iq/yWTwi6GViLpGj35vSZ+OWYiBt+fu9ZpHR4T/eFgjutJsa3JxgACIpEY
tJ9GteOjKPafZoH6MTKpniRRqHv891VXEG4XRgZfF0AHVVTkQ49VINPx5KLY8AgPSkvFH8gWQkF3
hfFzF0CGJhBMKF2ReEXSIcgZr4LI2kdfH6Ic/r0iepPdXXqu2GTVHOlDDLPvkvUuU2WjUM9ZkYLh
pYlmIjqCA6mDfq7Xm1DSxr72QkkdxMzSV9a0e2VHtVon72u39pR8XGMMv1+kfRRTzfL5kyrPGkTw
5Nw8evPsH6j59kEMTiTIEZ7tFiEMf6SuHsHDK4uVFehLREji+wl1Rtl+sEMITUr1dYBpcSS7Bs8Z
6lgGap1zK0VUrfHelUQS/PuYj1a8H+n5nkpfoFpSHRand81fuv2S8foQ/I7pWOY2+S144S1wMT1C
7fpYVI5yurtS0qoqE8kVW8V9jyF4+RVbAFXUxbeRT2J8WtlBlMgg1l3MWXBHJDZH+1PfbC0DAjb1
GADvNQ8BcqIXzNxlqwuimUIiLNnPVxZ5++XhDnRTaUTTj+0hR6lUZMwqZ2Y6TZqXBo/a8w3psqG6
8NUP6HwQ968wRHEdAbYj4DqRfZI8O1lZfveIPSsilXJvqjroyEB3Jn/b5Is1bQcWvLu98gHVr6na
IQWYAR+9344aWvdKrPEwgz8IRlyNB5ePiLeHgJjdPYDiHygWXJ0ftrTpfBzvtv2/692OKIPtIzeq
73cJe1LWL4glpypAcoai9y4ew2aoCMxbfc7+bBExqRBaXJpQE5VFeuEseTnLCWw46fRXnSuW8L4u
CJzBTC7zqlkRxZ31hCk/2hEBsGWhtnL+AZACqPCr68OlUp+iZhxBD8RnPskAqn8bGNkDFnqGkGaW
AXF92Y5tVN40/Thy55aPcq2t1Z0IWsDIAMGV0q9t84C+dO6Q93Fz1UCuYVgxz2u8tCoPgyF4oN3m
QZijuB5n3bcrn69nKqyDm6h8DnJibrQa3iIpsOxQ0oSmsQB2qVmpN8foY8bSyozawtRxouwlk96t
ZEu0xHNF2BsxRCO71BUcJ5nEAk5CPSsziSETriBHPenMsBv1vEYUYXrhKt4gABZrgNA/I6SnvBML
6d7yagb5rHBB0ogFxnmXpxMzLdiJMA7He13LugNxoZQuplOn4ph12e9dUleDVk9ytBpeNv51NZt1
vkhEuqmZ0Tbc6uWPYsJJflE5NDH4PtcvXggW848+vNrb1Z7h8s5nxwPTZ0Vl+18fMgeyzOOC1t4p
FWNw10AfpjBpAUiIIGFwjfOkf67rgq8QWRo1vYDhBjdytG11ECMiTOnTfXRFhe2LMHe0VDfUU9VW
DDdMCYijihjoELCM4V67aGUIgfDsWVvOZFU8H7dmak/l9h2fa2mD5+2ebPQfTwGVBsKFp2/lFzAD
AjR376xDJO2kCOtbFgkohyJmnmR2o/Ezg1Dqi6gOd20qek2Eiltsh07Pgs0/Fn5Lx7pYjRa5BGg6
M4mTLEcEANljLvmPTBuOZecWwjY/+keSqn/iAKskerRMtdVGGddZqHHN0ufQc9ecEd3M8RA8n1L5
N5SGNnh5z8zd4BFmSrXvbVzDjuH2iVN2axTjdX2lyofPKPJRWCLupHuVWHkIjz+hzq1fUSL8zyYL
FRYn9CyOR3lQvbRjix90htXbS9Gk0EX4n8AlsDsyeGdU15hw/zfwslVueW2U01dA7G0k+bXr27ao
TyK1EtjqHC3OWGVUlvNT4JPstXCa7RgU10MYpE3d+sz5EHmIwqMUAirs04m3D9d6VgzV4k0JU7GA
Y/O6pkQ5bagDLkgtGnCJ7enyo521mBAICERnvlfhQF43Tw7wKdGi/7kjv7iLB6IcJ/+kNmiFiMLI
ad73jbwNAzywi9fJmf+wrGzYqgaIM8Q/U5UtWx0bQ5CJUJOCXWHPNk0yMuXMHUBYn7uIYpCYfM0P
nZYbkq9zZ64CCDNoN+N+95q44SEVP+IoM5DEOWal1RF0T5kGy41Ho/+0LcgJVM9NYVUnJ81DhDYt
Qt4wrbhE6dogfwxrFOppdEMHbHzvfAMW6vszZ2L6M3Uh6h8ApYSw+Xu32UwK9ryzvHnXFpxvb+V7
rMjX5IOkedMeamVAZSRM3ENq0+FroHG5XT+Inkx7VKG3bJ4zwgfFu4vuKRlDrjmVyAmw5VGgf7JW
1Yb9Qmdp+K3gOXR1BLAHBrVcIxi9+wrJxcct3i1gPZeVsN2DuuxrnGjpM13nrWo5BujzrSTmRw32
Mn5vS2tcmO+vK7LzqrJhp/nNt3lLo+/9wiFoFVYTU6sy06U5MyBGaTbOa1h9OUpSeJ04brvqaIsN
5HCFwawjIo0UyObaKrXJ/5acqGNaD9MdnagX74v4vLkAEo155tlH6s+DhTfUWVUZ/M+yyO2GGzvJ
ff6ZzFZIpCXiSvKvqYcpwjJTvTTNpwtUpcL+wGFfqvO2k5P3u3XwEUPG+qxqSUP2CYBTcEADVrQq
F13OPtIqSfiyjE3dZ7OhaBm6jpyeqNVfH4uh+urYhMnVn1Tm+FJ6yO7/hSmYmVQem6nmYkw12+RL
LIQIxxC4ASC9VMevf0Jc9auAiw5Uk9zkOwpHmB1wRHiSFQUuPL/N+bVTE5t5oZ7fcyNG/JuY0VrN
fVHuANnyQ9umOa7EEC141ekP9pouuuTtBoCdEw705X+i8XTcpvxdKNBp8pLPG9X0ZE8UnLke9+Tw
er9hcowX5gePMHopQ8a6dW4TDdVQ30y59+jbFIW9lDux3pXmABtWV8gEZMGrjgwoQ4ElTv4VUznr
x8ORHSMIfD2YN/X88GlQ2Ey8AU1ET4gDMghVprNp6l1Dc47TesWevobs+Ean7gbPpg+EEf1AJ/lU
eYv7X18RrKvhmbDPSsQ4V951cbadR9mzikOxt0JRVwDh8D38UTfnFBQK9UsKoQMNHbyVbmSetWG3
2dUFuD67kcdglL03uDjY54dhpbOUKky03cUJKB3QzkbmVVqYQH0+jxrhD+6+1s5z/XqQR5SFhpHN
JpMJsX5Ty9efubmoZQipy3PB0DxkvyLLEhE+Wp8852ZRsA6QgU0xfZCqjl4V0owzc5LHTj/izUu1
3qDtt5XK5b3BxQqO/agGGdPKmgvDVkY0ifhvkAM/W1qU3qWDl7SbZ63TaVYqJ4Ik3GC/5VVoAPiC
2H6w83OcJaT4LsUX/yUYv3SIajz8yXI0LM0FIHcg89tJSLyELDWgVN6Pet7eK/AF96IIYYcpgXl2
pcl5lC7Z81aAIdtehsPexssndhD1fyouYsoOvhNRIfZUaU9XnWKU4N28aaFbkgiPe/l+BW3leqDo
CvnZvtqXYKVxzSKEBW/w6zSO5WBgCV3yRYtUQ589OLKQGrQqvfwkdpV7CMEDUw8U2P2gsftrPbXk
dVsJcBIIuBkDQQ6ZFpJjJtgT9c94GzJlGQEw4EVB6YgpF774Zfl/b/YkqGJ2vjUHc0I85hyuGa7V
wx8Pc4TFw1Zgj+butI9auwjy7LZHPYm4EGlaMOpOcwFMv43IrFzj5rw5so87ENOVCqTHqHUb4sZ/
cj2HcuCNjshyxNTqYM8hjc1jGICnwF3J2a91WBhS527z2GgN3RcXkncLDqUjP8kaO6ysPEMy0l1a
jHm8OAZC5Fgpb1F+CVgVRAwIybaMIa7fPSUeXZzoPujMY7LZAJyi3mQCOrkTiHDpGuhIwgj04JmC
EWQiElx4uBesE9wIemaQeUt9WObu2wlgDtmF7OsLXGfQVYwolvj7aYnl6X7gSNxdWlpThhfaVoob
SGzrCHv+WooVKnVKr06GhMlHJ42c5pfdOj9/cE2HdvZLEFh3Uc10XoNLuHpm8jwntFzX5oQRsaKf
CJswd7XbM12KqJDwvykqXEcNGfGmGK4I3PLrCy/oCcptIIuahUYIi2Z0vMZuRJW5rmliCccAy20h
Ac71lojfwDT9UblJtGC/1ImHpW0sJdkmb41GaKqZ8s4SMQDJmSXrZLXfKadmdOpGLIdmtMH4ZEB7
VEtsKpt/z66Z9gHSLapeMijpu3KWvuy96EsNxiD+BMMIWnROWkFGq1sPz5Euh66b++RZj0A0Ujal
W5MTGn2TN9eLnw3+B0IBZA3h19H/eB3sQ4vbdwm52y6juGL3SwBTiNBR4R1aJNNilEzgT9bH80dH
7QdZyG1p6BmSefr1fw29qfdTV6JQkHBim9JxClQxCjMPeJlJLwE/vAOlF/KQgBLAFME3E3ihFOrB
n6I9p/Xv5z+vRKCx2PnN7P1Brsagtni5YPbqHiUzjfyzo1QRhE4FVAFN6U4NgTjtIb7he5TVswgI
3nWWVdhbIYtlUy9FXokPS++TTP8uPIr1Cs3XHPpiMVFqg8VGeGfpwVDKmZnQCFVbdxnWq7CANdGK
cC29W5YWj1j5hDJIfqEkvDVl6rg11nZHnWTE0kvex7Pjg1foOHofbHoXmyad6+ORm//YvysowxOq
Fs/t7oBIy0XqPAcLjJJ0yteEhAUGul1ltgD4taIvGT3oLlCetTF78cxIzYl5/02X49IVoZkoR00H
Sh1/qtC5r16BmyQ+ZG/bnz/tm88MWyylQZIXxECrv8H5hE+kH78KBv5oFdXoqW9c+5LPPH69dYKh
Hfa1MvgtM9VjsbVjbg51z6+Dk+g2gbVgfKfxJKa3R84mrQHS6jwbidrnYFE44UPl+YU8OAxhhVgA
U8+E2JAEXoONL+e+XRGfBuaYL9B4/QObFwftg+HVWqYxxaAl46WN3KRVdzQqu70fBuYgrO4fmWGQ
/TWLip/WaV4UVEaqfLh+1oJyG0zhAx1zBs3rctUnsGJLNiHSQ7D41Nh3c6McQR7FeJ2epw3YsiMW
sjpWkN6OWxRgTWjfjAVcyCfs+56fVc5bfjEQbmzo2d24sOoQtRUW9JAbiXSfqb/XnTWf4ZzZ82qz
/1MMNWN3X7u5r3dox+UGHvihpvrkvBc0OZ0Id05xeY6Ib8KuXds/1j+KU28IjD0HdTejIO98xED9
XPdXPdV4ql0sA2U5cRaT8iW+3e0ZDP6pxP8k0uIPQQHnlucHgsXfMyK7w+AG2RhuwnJG6MnoBjJR
Dt6Uo+hvqBVgVVf8hR70hVjn4NvW2ROJDExaxxGfqoLNXulgrhXkF8lSFqXGV6r1Ow/lI1RuZ/Ey
aFfXPXqiO0sv8WjuDOPDY7XGI4h+KMPeM2EF5T2kM6lZgAu390jYHzmEurxX/T+gWBY78cu8x2P4
s1Z4VW9RgQUvz0EImWDP1xjYst/V/XMgy8ftglEMJg/9WuT8MBqV9cvjm9guM+PHBRFhHh6jjeQR
1oOw5m12tSCPh8tc641SESVNueNhs2QTucxX99UDeaTTTilIjwkV5U7xXODCvM/EveWojexcPJ4E
a69gfmAGodjZv0DeOeVPiGge8eGCS60C3VZiNq0LOddhMeTNm44zU55MW2QVHvGcJHkzWOE+s3MU
RR4LspgcQau07Rn8dUCFBz5C5ZcaNhUykfMpT+g+UVOu+sfkI2md7xWAhp52Q4gyleeH31SduT3U
z0SFlKL5Et0pc6Lg9hDvNxbQB+Gm1PZ4eY19gmBUwbStdgG8udKsfG3cRD4OJR6v6mIkgNiesAED
eY2xTRtJc+gil1+YVTaBYQcLZmNpc9LWwBpYJtqrK1C8kgJ+OBs3UJMBuwleubsvR7BQNbwKkqyu
tO3OaKraO8uEFIbM7RvLo6fYME3FbWPomPL+lpMqVxDRcvG0bm6XRLTdqAIfIQZ42LJagcG+ep6v
kpp68lTYGFBoICXQHfzLO85veT1M6SF7T4cZnZZUn5nthEhvUtrkA+SolzcHg1KvmYoGw3eb5CzV
9MNvOpnSzE8456UgYbMZZbenJtWDYS2ec/uZS28tb+ICIEkbjmubrBfzjsHty2WyVvEkwEGQ1ypr
vhW1RXHAK5jSmcnhXanSwn8SkRrbpwNAfkWBeiN3Las5JSV+XbGu0buMpmW+1CriUumLCX8PmEzy
n5wLF6nxIzX50YxsbOCU5C//+GazN/Wrk8G+/230QwlnzZQgRsSU2CB0aqhW1FJ1+QW6yR8oWvPe
k4A5Dv8FpZ3mVP/btgxQ7n2BYNa5I4Agt8EHVYzoKvZtx0NWUCR1OG5AKNY+CRRKaU1SRiRENyz2
ATEAL73tBD6YMeatgA05zj+KeWzV0a05vQU0hvLlM9OK5Hwa8E59jk1rY4MP++ABGgbmSyJPVEGg
GWXdMBu9hGWE96VNJu5fq6xCHPS82VQKYWKQMfEyt5421sc/PdFi8otyrTOsY/Cz/2ydUGSoumpP
tIHJg0ZsxxGapsU88wVgwhm9CsViAf/tPkWvZrcyEL1HGwM+Q2h+Dkd4YbIz/lRgcrrX+J/TcdVS
oUQ2QaXpsB6R6bE9QkbcBC9nZXB9S2HsFnpKQWNRC/VwXdXCmMAbCuvdyxAWNRJXg/k3xXxGgaGw
1DPi3sVRf3yyCDxBgDGtkKst8vqh2od24A96d1FrGjSbDASbPRU7evhdbM6tKoDtxgwc3nnzOoQV
kk4OydBK6OE4yi0Xyq6cryPFx1h5a3BTe/qrbNJkGiFNnuqSY2RyvNkI856na9e19LWHON8GfExc
X+4kyd7iWsYllS/3bKPOCbrhPKrKy1yJJkZHcpsN11g9gUXtHLzGAvpnk9ODGW5kGcP6296cqICg
lDhtsDIr3/mR5DX5e7yLEMJ0AYWgWHFapcEEbV8xo9dg4EKjVVgvo8p4wV4LUEhiU38/6sggvl53
77ns1cBijrDS9cFYJVF/EWxff0Rag6lbDhbJpmzFV9jpcE/QpbSJ4CjLmBIdw03esgd4r8qa1a8r
ZP0oWNBVZ8T9T9eUSoUqum37VMigEOTsJazCs9f6w4CRVur3NfD8cx0d2IKwgvH6hoNXR0u0vYkc
Paaxm5cdJxMa2tpe6a2REXjlHHpNYx1UZsVVywyx30jB6ss23WIjlVctIXP+FO49RfqAAfttV+JP
qmgozCf76qaODjFejTq2qv2+OtqQjKVxAOveJJ74sOfp0i7ilXjSuebO+h3/B4Z7F644d5e6zOHz
SnIGTGD6/IAn+K6zk3J5dzezbypO53xW/prwk1tUBqNgKra1mZswnZUyJtW2SbJ3SglVd2dU0+Kf
ufX5CgEhQyHn7yXQUQuaP1u4ASfddATHG83fxF58JEyLs5lbM6obwX3fcQZnwsPKQFQUWC8CFjwd
x7F+0zWNp4pAtOEcbA7oA2OL0bTgs90iJeju+6CayVB+bAABXkc8uxdxFjrSYLczMYr/hF3vS3Dj
bE2kRLbOGYKDlr2ZHXrBMfUjm6K0QgFFh+T5gVIMAjHGxAXfMpzjeKEK/dYceCBi6qBGonPV6Xx+
tUcRvFt9wq+wUlYp5OHGi68+vsVqscqWOGGJ6rGYMeDnZ+6pM/SIZE0DCoBUzw/PKE/vK6dc73CA
AVit6giWbwAe5Aj/FE1PU6KHWNxEKkfd66Kh7ek9tIPSpMbKGLsaV+lwQ6bk1GPe3qUyMayaxcMF
SEjS8mGWsU+dc8qvL3ZjZ2z2Sqx4oqVAT7mKjidQzI/r+G4p3YaQgMXKRk0DtE4lUgmudxJEkZ4c
owzJA4HW0VLD2/FFICLTBMbGdnyjMjnPp/kpgYdgWMn9pQeki9QfrVZhJls3v08NvFAox4yxzML/
NNJDKLXqUPd5+YDBOGCXJef08v2QjXsl8TgweTyZF1fW6NWeKadzVUJQePj4zZ5jaHxC19+YEVd+
UxpLIRCNjAhl8L8IMyBm+Syvhg6phbFJDUhxqK7roBfjodfVf+uUdWXwr4siCmjHjPbOK4gObaXv
A+Dr/WzyyODl7hUxmleYx5GS+VmwQ05Cfs5D4+cvgoXOiRHL8faMRPNPigcqcnWnHYdPR7MJN3Yv
K0T5sDk7dtKL9A/wQgcTr4wTQLaymIhNk/gwpCn9XLcZwXN3Gna5IX5AnrK05sDir0VVrc/oB5Ft
N2ihX9uur3IhKBEEqLeoDGkywF3UfkYRYKRCzHnjcu6XKsOVqVnS50Mkeejz++tyM+eMz5IJFYsF
o3nFL3+qCWHfhGNFep3YM30YoXdZIt5Dwc+/W3GJ7l7xd7j8m6XEY/W6zrHVP2LYH41msOgIPSVF
TFENmVrdTtslieRMyIjnXj2UUuh5F/N0012nBXNvaZsUVzvUnezrpfadxWXzD7jx96PA7Ej9Cxwf
MWZmpDXje5kcA0rvnUO6RIx6ad8lv9vEbmaLC5TeZ2IPwForxrZl+BOpqC3+mkFBoh6rf6F/odhE
r0cIwwtAixf23VQoEo+nC+W2Q5I+/M5s72Lhe0JQZfPmj9miM79u4+oj7VTXeS6xUUO/SdNBYgh4
lWXd5zKqYuxBRjDCD6Iu19vbCgyj2RBp4ZX8omS7EUbkA/UhwAMneJTynOWzY0+HPvg8G1BB5mDY
30sNFJrR6iM/+6GmswggJZZhcDZ2PVpa08bMncIoVVojJxgRUsKmYaFaf+m0uDQYbTNpYq4vjcCh
8b2iQxRHnbIbA1z6z4KNyFxojd3H57UQthIBTJjwfHM528FvWUrHhSiAJsAb35TOfdq8fxspgPwV
L3WXNXGtiF7XgUW/5mx/+k5XyGdR+DQ7HxEN5sjG2583edOAa/b4rULn83djg3AB3RHiUYfA6qTI
ZVk5TI360Kd4LQINbYXpkb6QwPB22IWgUInWek+HG/pLOpJvdRcD2u4dKfKJf8LPQ/1ZNpBm2Xl3
q6ynyk6syFgoUx6nAQ2KAtVW8nl5ccmQEU+HGlU0jPnA558QxFpejXSxu/NhvcCQ9IAObmkNTveC
l7TDJDKnKMdIxJj7MfrRZjtily566E1ebKVcXELTDS2FlZzbgQPUXDwdiePELTHCkas2JLs4stKM
k++b2N/dMyIT4YsvK35xo8JUcouxO/eO3NOqJz4RQbXEE3OjcDqrYaZBCnE+lWAIkm3GtoE/lbxb
sCEfhVAjIBgg1hCk0JO0ON95Vz+Um61di+s7WWjoz6MCSIjq600hrcOXhigN03fU4918pkDNNanx
4EMFyR9ZuidlDTbfrV+HJaOBo5DK/UXzkxhnzMUPAt5Mbf0zyw==
`protect end_protected
