--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
V+rcMYzWydrxYXeQqU9bTJM7wB4KsCLY1R6jGLE9O1IQSMAUUNapByLseCRwERERprUch+hEMvXj
K1FiVAZyNFI+NHhCpygmf9221w97+cGL7eNI1PW24MmG3CAN3wcXkWLtIV0gm8dfAOZeEqhEhTqr
IM4f5N2eiG99p9UiMJGcfN3dc/2OqH8egiCiU63Mm7gPIPnAnHjiRPvStGv9BO3PUZjBlHMXM+KV
UWnzqyvpRWNN+LWbLQE/VRXfAtWkEsfsKPoN+OB++KOoMzJdQc0sO3t4Ea6KQ/H65qAMPgkQBgMy
24FJRcOL9pxeQNwK42XsvMz7oJUnkOKLOg431g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="1dwXWFIdA+eD73XYrA9m6b6VAQ0RDCCNsLfNMQHjSVc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
JUFTgLLiSIF5p8XT9N2mwFtUd0LF4wG2RGLIWgxRvFIUNs0FEnUdO1TxrUf0CuHoUX88taRaM1i8
jDHD7ZwIGM1nCfNakDOxNs5zdqiIE+Bf8eEH3j1OL2Lzfh2PYil3a0wNN1aBFrTa3S72G+tdSifv
npuRXycXYVRyib6odPG/VpXhhSLpM943QmBwQApD66AMhr7VhSfqZnuehS8HGyzUqYmm3HYKCQGu
dVh7JmkRUC1apNY/tvHY625pNDkcuHXMmK1vagfgZvIE2SgB/KxgcaEbElcJSFf1111+k3M0xYka
SYBJqx2aWWeK8kKltjtyFi26vpNDXqj7sfj8FA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="IL1Xh+UbypupmhP17Wx/6mpDrO+YtO+42QKS/QlcuYs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 36560)
`protect data_block
2ay5W/k1nMBXayWxHG35w7y6PMH4LmdLKfd2akIHa3KpXdZ7bGC/9qBPkv4mJ8WnlxFAfdR9vAGY
QRuQkuHhG0wl5DXe0t63c15Xcoi74dOB0fLYro55Pkk8+Re2X6Mq9emRbyK56zznpevMlitk13y7
uCm6br33KGWKY680kXlt07Gjw2xn7RoxJCaX35dIN2abf/HC8NmwvlXuZVzo69i+3bFRtBreLXtc
H4+GtvIxLVu6/PVSuV7fsQ2aOaZvQKXccoOYI0s2PdfbiWZEkA63BoL+GD6nakxZgWnWfQmkt8qh
oh5e/LjGHFih5vYmIlyXke0hFIBjk1e1jGCQSruBKPWAtif3x3zW+Qyj/srS6jx0irqvMAq9zvoL
QGfSkO/4ephX0a3l1ogERubUyNWc0ifCblxWF0R55oNSSG5A/BSeJRUQ7A6BQwp0hov27Prezc2t
E0ooJ9YdjKRdSXaiMEJBY5B+ZpTVIJSDolXC9AYsadE8bpVQ2c5YTBptGXY5GiCp1UPSj6AhJ68X
dWjF1BJdxzQRXcJ7EZNyDgEuIjVrkDGw/FuxX3dftQgz0Wf6je6f9lmxlhD7siDJO+2uCTGNL3Wk
hWZjC2k4vpAE7K03XHD1MccJnl4BYcC8I3XykaolF4AMap2ihO/ikYSN5ofKIuv+ZlG37dfbyh6h
WcDrQ/bZKUfKVPgCdAhgpPiXz/QO6o1arwmG2haweKj1N/GjLAN0J7XVKXNneUzOJTe7yrKVK+g8
oxtD5XNfOUsF8FDSr9oPmXlaEfHSAb0sIvWRSQ93/+l4eJzoyXXLhIkfw24UHAApEfPY+VaSrPKS
EKRHDmsuVumcBqUpJVT6ccDd7eKjtaiCzkVVkOEjBtnOXAhsRZLUXv3mX82P6zyfVR9MK9UPKmeO
+6y9exs48ZEiL7XdPy8EvI+k6pyrWfsZ8Rd+nSHYEmiNq8x4bUnv9X3sNnYpVz5pUNFIr6A/Hf5q
wNViyYQkM+zESfAKRlCZqfiyMuvp/41XrihC4DJpVJgof3EHkG09oAfO54fNzLCjJE4+omnAQwqp
+1B06Oz8Q0788VdXudZEEYgwgwTtYPo+FwgnL15aIuOokk2pMats43VD60+ufmQIU3owNl+TsZZA
m459005efJgLETRgvvAc/cWCRE4l8zpwh600WmGaJrYDAMzxOMONokZm/795cNK07zDDm12ZsUs+
cqbMLV6CBVgDiVWTPKFNHjpcLlTegy6nLoruuDkP6wa9nlpPK2Cws+/N6cJ4qeil+b8/BKg75Exx
7JsQLeDaP7UgV6XrfGDV+x1GxvXf2UEV9zQjH6Ih5T2Qrl+aGaKFbwgpK9m4V3LStygDFqg1B2Vi
v1h5NdbtfqO5k6ThrNb3yCEpaQ64CnMmnGdlSSUbHSxoaJWls7TIIneiWevrOdMpIf2Zx+wBPCTi
hnfeTK6m6xWIsvs0z+f5THXoA725nHBQmncSz0xx10cWBpfv6X/wS5PGIZwcUV3xv/4eQQ030Lb/
OtZ+8bDhelzNuzw80t+C0Df/olgoV2VaeR0d7/qF1nS9RcAijG282O4iqsD+7YchBDY/E7gEfowq
HURtIXWRLhlidCRSitZ+NXHeFr2zdabOnZ1fKbocctQgN4KvVohsEVKRFV50PGNEILJ8eVl4mKGU
Wel/HyvCYd8U9Pu4U6Aobg4T73fqbJuJWDJ5wVpfNCDsXFOows1KreV4T/pOPdhnEWlsChwfbSH7
8P3FSR8h6HlpuKa7Ad696tZCBnpik2p48HotTp8zMdiQr4KObx49k1Rtr2aTsNKzZavcIvMmp4W/
Qh7RCsbQ1+cCjo92NEilhEHliz8TIaYaqhkS4ZcIzJdDrALpVdvTvXdb4t6qmJ2R5VbzBASbHHPv
Djr7xy40WajL8kA48CxgEqF0UUO5/wr84I3OoMfixouRt1UbFnfZ5iIUbCxWYcwqoNSaKs6S+Lkh
IazZtR6m+4ftOoJWRpq53/uQtgTt0W2haWX/ocAUEZU6d5OtmOHyoxH6GO1rr6uS7T0KIQKGpcln
HD3iADW3ZhEdzrZhUwPd+GJmsOKwp8PKPKeQIE5/DpVdMVby/aCuQCf3mXbcJ5xtfdh6IkFDji91
Aqjd8nN6ZXXC2pgVCw0zhvf5ZNQRCYP6pljX3GDY7y8qm9d4f+bJJyquT1lN0RgsiTO1vukrdoD6
4ntvvgrx7lvC7mvQf91HjrpS3PqmFf78GexUZiSo/hL6sXXOOuKvDGZnZl+ugJsdrKM91o2GTJzf
u2lTdN3hQXyhtC6FiNv5QCIyJ0HvlODR91jpuEyM7s/8fFVHZ9tHB2PX+niUHGEUeXaa9WIQZ8sJ
O9qiVN1QfdO0ngu2ioH+ikYGmpXbzNuRlPK48RldA4M/zpDV9NTi6iwrktpCi4qcaWKWfayjt8Zv
qD3NMgApQQjGrzH9C7Xds+GpLTkS/1Q5jG4eWpyHDhv/Cu7fEitxYZAu6bH0VBOei8BDrCpycWAI
hPzt9TAa92mMhhOKkpPBusYXiyiCGtcqazngU9+IR+QKWm1YvX8GhqDCduorbKm5LB3EWa1bTjHY
owO7mjwe+tl9qe2CvrdodvSkQTdIdKU2TIh0gN0UZsDUQ/OcfTEcN/ZLr5nY8+ERcs9J6Dqu2669
PR2XVlcUut4LQE8//TlUEyxq+wfJEBHNPiPacCmCA/ABl/08pczn0dUAbqj7snSowZHp6oEHWY1q
A09zkxpzYwUx0lstP9aZu9Alsloy+CTmg/U9IfS4FYWG5m/03tr4WsQQz95bBtN7D6KXVimTWdjC
N2U5Ww2JSh31SrrPFFx89U8fh9vcyn/l/4l4IpECw0NXkhyagIZZ1cd6ODsR02mryLDbYEdVGYIk
zkQZcnBCivGsoMafrNpRQ5HCh7xataWxH9Wayk+b3gt30uU5BY6piHH8d7Xv+ue2lGhYdUJCgZbc
UHRtj466fsquMRcHiXCzohB9ieh8SUoyD5NNccXkFVCSrqo44P1tc0wMOZyP0hrU6C27DgwuRmut
LJjGmVleRm0I7J2LoJrVwkwIS0JPS7PBvsr3o/kwZHjl10Snbgiip5YQx8SvEdCBRc/JtEPNeV1w
p44zwWoRib2BQuIKoSQhkJQXQ4aCsSA4nGspxwXYjHsONtmoRlDty+pfC9cQps8zW/w5+Cz3x5rC
jju7/D3fjPgLP4cXNiApJHYDFN9MZJyRP8NjtEgXLJsiEz568vPMkkhdYMT5TEzI/0gcaleZx6g5
hi1vOXqxTaK6GJeZLDieb7uEW0gk6FIMPBpGc+FSA4dgejpEx2phGyMxZ9bIZJhArvxI8JgkFjmq
KCN9a0p5DOSdF7ECkEfC6PHNHUSHBE355wK6MXbGIzekvYfFJL4Q97NSUhygZbB8t10caesAQKQI
PjFTXCvE1I23P9SrQJuHWs8VzTV6DzObDupLXm92H96wP9hp6FnDiGkTgzAJqRxwv4duY1CxE6WL
KmE8WziaKRIQPr0BGpbVINr8tox8t0SXZ8sINJE1yMJ1zs2avjisu9hnSpJVxOS2eFMPBwXAb7ge
p9KBTjNzQYQVRdstvLJNXbZixrFoQnzYf3nTGgmUO7Y7iTvcq77r0bUkTkGN1WgJgld3xqyVjeBQ
++9KGxmCNvw6b5umZjWdDOF5ylkiG4A6Qh6QUN50WJLawOlIgJtCkUpEHTpR+McR8u/fsxv1T61n
/S8ruIv5X1Wi/FeqY0KLe7fhkXDvJdgqEGp+XuPw1A69d0ao+ePADOIVcjOQFoIa0Imm+Q26qoSd
ZeFEBjKmsTCzmFMO80+p8eJ8VtZW/3AEvCRxIW0F8Q4BiVO6J0YdRE44pUx4VUuo1S/ZZ31btxui
ZGOOqewvtoi0C/NXcqh4o0h6As9sxyrDp+rj9z48ciXwAee7enJPYu+x4/uHgAu8HFKtcYOXLUoT
y0/Tk+ERAcQryWhylXz33lBDTxpZ5Jrbf/pU2UXjGSiLr/w6tK/vKTREjvwb86puntxYlHbPZNqI
oSq/AtfTzsSM9Hk4fNLbr+x1YT/RPzFbnjQrw0wyVy1w7R0dkDLU/HSAlPVL7rS/l+8t0lTbodsE
ftbOEHb0j2E8cmEmi+Vau101w/o6mnxmWbyZ6EeGGPaX8WhA9+8dSdwQ9O7XY7lUZuj/Ee6PBDCq
u6kwE6qvu6N25poJNswM2piPUxnKTpLx1OEwsxd9uBvcYA048/1vxvBw0G/lMF0AmCvimrM7Of9x
0gz85QPENjifb7rKGGYpWrnx2SBNMEFIpsbez45ecyvOEofjiNL98yU5yAIawCN42zbfVLYriY6r
zGvupCmdvjIJKKN8xPl/nLCj43i69CYnhdHAy5x1bedjh0VUV5FQU8iTqauWJ1eWG5WFfbFheVGJ
WrlRIgSWB8Cxk/HmN6LBlUr415Z5Lourn/PWCrh0uKjGXMes3bf83cso4hQF2wcMY6vw04djyajP
lU6cNU/k97MeXy9IW6OJKtdiR8nCdBkk266yJ5her8VUhxQawUHRw3NDlm+7WIS0yQjIi0PClHtO
IMhbPP4WBLpIBBYPbifxuhMUxeoTQ4EzXkwZAeZRgCktfVzhQ3M3+MzfK46EOdHGuAd9/3s+5Fej
iox3cL0oF1Ys2Lejq24Ve8VqZCVDCHK8L+FjV2koT3vaPfYtndcBTaF4uuNKxU7tleDbfVveqpUM
7LQPgLXmOWk20LnWmNEmtoaRasS0Qz8WUxqrUvgzJFLY2JrYv/rjOlGmGzJW95vEhQJ7fmm/OXrY
5rcH5WTPSJ0pKo7b4Eu+EnbTqD/n8MD8TA0rk8O4DrlHRr1tzGczCHh8uEudL9cZRW3tGgqy4Nwu
G4ueyzjRi3NibJE8Q+bzDUKrUDwVXcS2QW8J5hdNvxoKliP2h15rFXxXyqaU/aHr8SiJs4Sg9947
AupFB2MovsMfxev0Kp6DWiWDdQCpfNX0B3cJxJNyY4aI9Ebvtm6GbLYBQOkD16Fp5uKAUjv1jSj3
Rt6DxJRgYfJxFCRgOEv73tgNa7u0FSdRuVPYFOPi1AQ84i6k2di7rr7jum2DwqLMEjy7fMP9/b63
i763hx8f5/kyhV6X/Mcazqw+0WXvHyUCQuKzpxFbJSiyy9wcn/eTff49Yr0Iygn6GwQJxwQpdQJv
mdKJ+R6LcdZzNlJ2TX0qh7uVsYOE8zXiP46g3/3KHRs1EfpcyjJaGcCAAqCWTbkkLGnipyGX4Am5
+TJPCKpTMhs7Wp8NEIvu4FB0y0eH/3zVLygZYiifnoX4NURqfXgu3Y8JeV9rah78EgkwTW/B9Mrs
vjBkWas0Wmqz7blD1QDFxgUd8F2cQsvb40I9ijocAZdvUj/2/WecvsFprxDbtsdTDhppCRK7aklI
rpNIhki1Fm18rgwNKo5IdcO9lF1QGvD2gVb4RVmi9FRiNbRrPeoAcjrt5TmSRNwEDkAggEyu9NpD
/gA9VtXTd0lJ38DA9mfbK1vyzfc9b0/xcJAXZbDtE1dE+QAlskTrdZQVJFC2U/D3WRKEHCnyZTdo
I9Cl28ECxxkkC5Www3674MGmTFToC/ZvNAOl6euVwGfw47uDU0vNl21r7tQiA9mXOVSQOnqUrtVP
O689rKMoHi+Oo4YYEFaHLAmHO+u8TrA5UiHr1CdN+w5qOLp9AQaJVGaVWP8pZbT3KRcWAe/YhCrL
fV6uy62vuWomcjwCPp3lvjogJY1/qmz5xnCJMtaOz2QXh3fW5a6eZid4yFjyM0H7XgbOqKMRcQk1
rSaqVByM0B+DFDnaxaU6q01scyyHJZBsy2q1qalF8R6AkOuEpfAvfcEaQjwm61ICTZMxC7zFnYja
rNteD0x7fmNiSm5c2DCR2wcQuNFLuaxVRW+0PwvTqyGOLcoC0xob1Q2y8bLMYJPGF/Sn9iHZNoBP
1TtkwQ1DoBPUdiCxwBVapIK+bDdB2j9lzIjsKj/1llXsVxJVdJ56vXRPQneVkgkVw/5kAjFb4UMe
OQy7LrPru18Xh5jjshF2d1EqD0+N30qNybeS2IBNnJDvcAJ1FnAv3LG78P3YdZHUCAAU/HNrWc4v
Ysiu6Yw2F6WG2Io2W1hkCgXwHcMmN5IDcxCqQ3gX2694IijY9+kSO8NohFp3BG9lI/ixwOUjyiJk
1jkvprEKZhV2K6pODGjLQNfJGfcwrzxgs8+HzYAXsH+UAdTMVaXLCBGMls3lN8KDhegYQWGs45zB
l+Fgmjibseox6Rt/7jWq5+qavHNcQQJ1jfFdK12wujPWQcEXDc01GIbvZUyr8t2yyNE/aZNUuLhm
wmiP0XpMf6zC6Gh/R5Z7FaGEU34y85f8ckRHUyGNmKe94wuZwZ85V5aTKU47+ZFBjHpuObZ+NYCq
hYOXC4biCNvcNGHjTQMHOpx2ds0N48pfJ0zKvGAzyCpswVg0zCpzftali2ZEO0iBRENb2ZerAtRH
iG97suyAcquAejg+FFrpunbqIFjlpChZmP+5I9xgLxH0UNe12HNKXBBaOxe5jSAYrpe4ZW1zMrX5
ybT1U6xxSj9Y9Hfb+i50l04CfaZUqGH2lHsxMi/sPPHu27an9QkdpcwMJ4yBeysw3lzvunZL6wxV
8Z764CQqkTRnHazQtyaMBoBtpBsqglN/sd2CKwn9W7zdaZozK43CYUivI8mMUQE5w6Rh7BUxJ3uj
igFy23JQDQc8qDrk/Kp/nF8hKWRUs3tNwA4jlft6UnL9H4lmCfE6XFhXKUBt2RJS9q+ABHpZhnnl
yth0zZ7AatfKN7pg0doBQ8thrSoZ8osNngh7/8jiFr49Txqux2LZ5C7l3W8kvoGoVe+BBCaWWWdU
mgrN40ONR52Pm8evNDddYx62dmbiTgtnfn4HDg7Aq4SvhLDlNEllrrj0SXkJlVSPwSJoIHP6nbUW
JZnszwb7BZEHkHnh+u9vuWKImcA6Izryd2QmMrJqsE9wbNqur+qdsfy3N9MkEUayv93TSiJqeqyk
qVHb8O7EgH6kZIywLUblTZw+Dya8oPBlBKPuQQB5nyPRHBi+D6ujzhqgEwp0oXBxALeyMNKdW0Ut
MbihsTRa/0JWu/vSV4vq9oBL0bLMgg048PfcVHB975bbwdhAfPulN0E/VngYGz/I6U2ZB7S1u+nS
4J29PGUC6/lZADVAKExTmiLYpnmcHbMlVJCB6klkI4oCuimUx8sS5vGq3AejhKcvtWiMHv8w7Iku
yVTeVoeOvBYeTj/85+VcwlLyYpf7+/4z6JmRtmU2CHtp/ZsBugT5v39pw1dSOD4klUFdxmieqOPp
0NMlRQEgY2vz5LI6RT4rvjd9pI1zjtW3mmfksVif9ix/hYP6Beva9wo0D53zpYGNqX7QbIUOhjzs
HY61wvQosjgV2fZMcan1zrSpCzKjDyD0KdroaiGQw3YzuZ2SfCqbIzVcPEAQ+jc8Nj7WQdjQAMst
b0+DVPAaf1sb2qbhTnjKBHGMx7KJkuwiwdKqFRPV+J09vmwxM4Tt9T7RrRAa/yi76Cw1enFPaWFX
xNpbyYnAp1GYl4f9kedwfp6jpsSRguFcP11UNnltxiDrQ0MW9icjVl5duimxu5CxpEFAvtOwVGpT
vIDfu4R6CaqrXiz0yrAz3MmhhIQdOjNNsj+Uf/CMxeH0Q4sxsiuNrGYLYtR9PtP1dvGO/Q14o9kp
bL863zm0j3HfcEkjA3PzuEMVAqb5Qy8SdeF+pFC2IzrcvFBEWasdS6zgAPtUr+VE3oenNdHGdput
OOOV3t3pp3O8sXcTaLQIn4sPoSChCoKMF94rSH6Gm09Xwot4MBXA1e9oPclYICzYkxLfX9pmx9Fv
nHFoJTOTLNjrcbDdnHyGGwVG3K4k1Gl+oUeBTk+TGSo4uGu+An7MLvQWFQVkFINPYH5729s/DN0e
v5Z3MC93GcANakW7ud2H2FeHIVSBMiiSPDNG9P1DbeV/hHha5JJ0EZhWGd3Jj8VMNRxq0hMu0JLk
iGjr5qSombebfWtCc0gXQ9gsH2O7YDfxTvjW15lDNLcwcQaaUOMiV6pV57+PhBpjRdaoqbM5njNf
VBK4N177I2ZjEaMB+SBMPYgOkCChQAMGmIoyEOgAUSlQ1DN+8T48ef/2QI/oP0wQ2CFkTSNomhsm
ceo56NHav+X1P8Cu+F16Q76QaPyYjFWiC4WItIULH03cYGnG0Uk8M1wqL8xRaIYvZrPTSxag+qia
Rq9GasHRa9h2uEyo74dUzk7PkvSYtZUZksRkDMdLnqHef04JpUC/wpYu8Oe8DISBGrSgV1QZEMaZ
p1mPkGOYk1mhbslQ6bJHBDvFwjdno0kTR4vBI8nC7UzrBkRh5HA9t+GTdKqEeKxy4S5uztGj0eCm
jK4DhFBEo20TolfqlWXxzoM6/m8VTsFz7rsB82PwY7pBWPlrBTEHLn5WIO4W5hudWeMwm3pF09gN
05btWBYq5CfD6gdUmkKpljkPh9fhTUzhWTQ6LYYgssyARbcGCVOj+NOh2GsKx5RzR8R086ShP2Ox
dIXPvzLDdaO27LIS2pp1kKnkk96GQjbAXkMI5IJIbGq8U8Mh/V60i69WquSIeL4WUtrFZAkDF/gh
454E+5uwbJraslohAPr0OQ+UOjnAR3/xYbA+k43zgbnS5pzgst6m/Azl85F9tPN0XIlLkxbCq73L
aHPVhOqw9eR5mJByX+0XMczRuTFuEw4Vl1TTMl0JZW25KXYBuB8kMIfVjFSh2db95u1ZRyYpAW3s
wQkJw2dyKrhDUJFhrCGXOY7QLR6gm0qlrpKupBT5kSn+iqUg/g4Pi46LooJxWP61RsiWXAtDkJri
kRHktyKlmKxqpmWSb6lre8i26DoWA68A2tHnzvQsnh46G8USsOSmFWouzFksYzfZTUKjfzMjBQ1w
5fRyN2XPTdoVjm92sZpGeowXLibw7IUc5LBH+K39DSEV5csSqkhQo5xiPrj1D12HiEfuhaota2tt
IHLPsntdoVBK8+tQIDAzGAaiKUMRSLx0kfZRVUpNJOyyac2JN1hdP+PzvBjLbvVxUz/xMKlfs9bk
gLAaoaPe+vTvzVi0mBLo1oDlsaj0LCisTxzC3fN0sQkrMzlrYJ9osiI2EpV6agOy7mf/9NkeLU8q
E5Ltab4wv4Ih95y9BArLJO/6izjuKh4vNkHrse/J1dTEeJaC9SKmwGa1Z0KIXMV/xY3SVzgbUb7E
kglIUdYln0afIuF2cKsEzZmyLYJgX5JvD3pg3llrTyC9QgpBSOiv7nkohRClR41sOZeu1Me6RGVn
EANmm1ydAa97jzKuba8Z10NvQAENOj5uvrwS9WriUMkbZzJLKw9VjheCFz6MesUorXt87/idks6q
CMQZPq72MNYjVCXseTQQg6btHYxvXFkg/BBpZh3b/E3g+okN96xTV/kxzrb0Pi9mvnnsEMrQ9s2M
0QO7qHd19yJLXFHF8mHFAnXjuAbjBHs8DEsDUTIhqkx9T+2/1gf6mOsYRFZoMRSB+5jdDifU++fv
h8/Dk6m0pvJ3AFXEvfOv9KszvEfFypYosudoQnPx4MmXphdz2kTo/B7t5o6/OzJwoWxAJcgJm3iA
rpf0GJMis6ez5F4mVzETO/NmAKtuuDuYO2CU3bmI54cn66aRAZiO7u6lrVMmBLITdvACiWaF7OCQ
jvxDg6vxDcWgYgssatolLjg8V+6YR4WJSfQijH/NnPcYueKlbt0sVZRRyhJTjisjxHIkUfA299g0
XyaNY9P8ZqXuuL3PFdVeh4FXXIFVsa4cE/Qn0mqpyWhHDuYzelSiaUeCL0ZksuwQ1CtiQ9uQhjrJ
AbjnaHjxXbK0x7YsTOaQaj3wewMfbZ0Yb25kYdX4N/ZuQS1TPV3mgMQbR8xS9J6MApiVAX+qa4MB
kuqUI8AfW8Dq3YdXPXZeCelyCE8749BhAoUrhOzLn2BW3JMJt5M1SaJqdzw9u4+l2pvoMSjG0fmY
KxcYu7vcaHRk2iAFUt+7Tw9urM5ZuS/UNhyT62EpyweVTm8JXFtxcO2Hcwr2tAxPFtVBfZkp/Gzj
5odLBCeCWsik3kdr6avw2cBIuXzKTVeDlv9baKJWm9oMg5LJzJWgQkemK0PTie9ZmT1RVlWUXopi
r+O2KmFm1nAEadxMZ3iJHb2ti4Fm3kvYlPxDkGgHOi1+jBIJfGfSoM/lxGdcHBEI8Y/PzGCPvw51
VqawxhyL6gbnSi1J2WvPu6Sx7mxTGpMTKHtn7O4joDGZ81/82zg+8p8XZNs3xANBEq+gEbn7/B/n
xMH9gJiZhr7LaQo77FeDOKPo4+NAsGiG/n6S8Q4phGTiCAoS092kMaU33m9ME0Zxu7LY2/2ezHQD
AvIUorzLclDsJIwhMdWusNJYMjZZgljChdn39NC37LCx/qjwnGamvG+BCfZvRSAPl6dkNiqHgTrk
GGzmvVpwkYM1RTVP/U/YoGtymC5GUEGDG+yInSdt7OLA9774FLdbfB/DXoPQLfufFxFy1livb82O
LXfBuYwZnuKcHKI36KThe8SUV+/YgKsXX0EvuptiNKcexBuxWrUIrJQJpnQI8FLHu9Sy2lgvv4io
Rg85Y+NfB5QyQSC+Jrm1UkhT7CcotXfgiK68z3fvIDf3JWs/87mtUH2B7f4TAHsiU2YpR+r6ZLXv
gR9JGS5+cpjkhsGCA9wo8NiZ98mL03JWL8r/iaHi6sJXN39wM2g0tnJa3+j3GwfNIGd7Hk1ILCWl
mkkQyzBFGTHG/dUFHlbAsi4gus96O/QCdNfmiF4KD683QQL398V3Nxae1Sc0MVbQCLxgS+PSGTgc
uQZasYWkDNp21oTZJhwzdagx32I6aV7RyyidXjZ+4jxaKODTwMhOCcFnYx5++3dLX72VUwSsMGVY
GaqK1QjVuwS2sUfHTxJ0NZMFXMq1IBtIVIobTWd40AaTqhYbmVDKZHNuMEv0Eh09S4oeM1dyx5tl
F9UaBxC/oRoi/1Ic8n82yoZ6AKEBfmMz0CL8hDk3ItFo60KvnYsDqy/icbpJcZVK/+fBHEIKk45S
H0/Yc45xVdp3XTsZfES1x9x6jZ9/D9o1FS+ap9f2yud75rl0ZSmOyGdtOCTpEDVg5fTgXbkRSX/0
VM/mTGuEPN0hXAg7if7yguFyge39jXe98wKR2uYiSBWVabGz+PKvJDCdksXlcYU7Wdaw408VJ0IZ
C2gwlZes9AcRAeEiUYcat2HIe+rBLFjRoRJl22zeokcyz1KrX/ziQnYPubmhHOoDDKVDZoSmhIpR
sFQwKSfJeblHGwcJgLK61tBNdJ5ijhSE1Z59HdtA+wxZ/kuOhJmqnsqjvOKElTC87E2uXQoTfbo8
/lMVg7xQPyyO6tJaEej7cNRaawtfCF2kpWiCpAwk1GGxQYU9SqWrKEiC/8oQpZVLOSUWTqrSIi6y
+kzpePMsIkyJQKNoKNB+q9mfnfwu8MgKHEChG/+8EBYWOKmyuTWqtRy698DA43znuAGI5JZxNPjA
DP31F1hqrrPZA/ISA0wUfau/I5H/kNbxfoui2VfMM7rgRWGbLGXjRnu8GrIr23hDvfCocOJSf/l4
CNOkJFi++r06nH7EAGKQAs62EdXOB3yoiaUOTA5c7fgMdYUF6dBz3jPLTyOL7IKciUnHtb93aqhV
7rjROQHFSxzRwby53rc62GYyscvBXj6MuDOa7dnD41aKH8DuD85BggXIUAbwSRC/kBDzRIPYNXN4
ttCIhHFdSZYk1CB7WusrXWwyMQxyrAGiSSEgEXtIAtcEw/R7BRIrMI7LKGNNYwpJ34GdlbcvrQjM
MsuYu2bor834HxYBLqzGFKR3BtxdaUzXRMTBd55wB0oBT/7P9MqIyMKa7IWrsYxwUvX9CT0PwtZ6
u0uoaA9nsYzXzXN/K7Uel43k4GEVI4D8NV3hK+MaeTEX6h5BTi2MW8/LpiX48+Fb5/81Vr26Mx9H
QIpvVYqp5vtkZ3yRE1kFNTvYKBhafsr/BbbUYHwv+YHkJVqHCjHiU4WkPZujiQgRgaJx81ghK13r
JQetSKPGx9EbOXLQdkq9FmeAHHvMUCWjsV0lNLqmiTVWxqfWtrsrWmefp63qr7yn6YT7KSBACiTi
ESHHCu8vKQaqrMbR/T3I6F6LOrSmCBPHy+fRrk8t8tSiUOeWoBLoORwC6CetnxDQTSseuqkgxgTd
WSOVSqHVK74p8uNedHT0lK7+GAJh2O8cLSlzctsyZfaiZXw7fLJzp50lHuOBPr3C9uXgK0qXxhEZ
DpaQaEF5qqxnTMvG2+qKlfRk5hyapPPu9/yml33ENz0/BlvRFashHUrwChBy154j9ACoIix0BuHC
VpIM3BsNoOay+DnH3X6b5vh9sTCLIQBqf2EjGHZ4LJgu85hRD7/vYYsy7e9kmUFuQWsXhQQIszi1
IOoa1NdnK1f/7LSdAm5PlKuyzZ1Ja+km6lGILBGiHcxrBhtSUYYGsWBM9/U0yUO1bHRM9TWSBqy9
7IFfwH6FmVKemkDO3XBcpV2yvjxA791gosaUAKH7b74chugl/aSLwKrbjxuw2NkZ3i8kXP134oci
ME5dsI1ra7BM5evts4fT86x1sNgxegSaBwsU5HRfm2SgD9QKw2a9FnVeVQJj9hFZYTa2dXHc7fEo
kw/w2qr2g4g3CAk01sKMeReFcb/4Jkiz3X9yNDqpthxE8GBi3HSk/AYJo6U5MznsYdcaGRVdyZZd
ZmVr4yNnArL1RiZfBrtq5ym6vfD8qTn8iK7qWi/DMh9r+l5+yzxjYamp1LtcpS65OhFyqayv/jI0
RgtP5y2iRbQsL5BRJcgUWOEDkgvzs2oHlNpHR1DCqXFee177JH9qFclJtIDRqVdxneJiSvXi1oMj
uUIUqmXS/VO7/jC2ShffiFAeNdztuk9V12cc9XeW0h2wTjbLfXAZatzwHVVv08j9529Fqz/YwNNk
lje/TshZazGgGbN4a9InazWmSeENQYYexrE1zjUvz2VBtpTPTDFFRQ7vzUbSfq213DHdTEJsPoOr
a0MyfpGgyQXgcbSy6HVJBQAQdDY06FIFKv3iSsPCr6D3lF8dRmwyynSM+rlaRnjR2R1MK9z5HNjL
jwwpnWvFvwc/r0EOZF6UGykU0ctK3sL/DyUCVWgsNKli9jI+d7MwfwbYTEfVJfQcDTVm0z24gcFz
IezlwibBiZmiOuI4qF9sBX6SDe1cWW4EiYvhLIlBDOH5Weg1/6iW8OIYDo7fDqoVKRtkrCQLqCBp
9wPiwJCYt3okEfL2Rhc1jYWxsyG3HMWVka1BJ1Y6XEqrpc/xEa1/OTaiSWgQSl7A/p50mKPgxKgD
xkNI7dWACDG0dFb1SYkrNtvu6Oe9W+FxdF6cigSFibxwJi+6W2LAsYzWR90gqHvzRPgHXhu57ndr
RT++z9WmReEhdB/kkMPrFb3TdWm993llUluMftfRSgLxiGTo7msCS3y9t1LPYFq9N3JbdKtq/joY
D6cBTZ0xXSWTIUY8s57oP9Ify5ny0ZB+KMwwRGjo6lhfNrIKILRs/xERjBzdmWO2P5IOnrkmkGEz
yFW9V4vsN02sY7MjV3rgHZWR8iCUHaqL0IqOpyg4M7st9c9z4SrePdIcRUblDPixz7ASFluGlHHn
Uz/vHkJ9sDQWrKo9SsvjKf9aVy11sPZ6uPvzGycdgK0miJglPO4m0pE0pZkPndiqhPSVbtoyikAW
3SQy34hpf7LcPl0WVtsOqgowmlWvnrGb9QzMtGUvkULYvwrTjo5tIRaE3jSZcavY88KHvtbZ27+H
ejh1ASR/8dbM75gnmSD2NmM6SyQNT/mMapsjuX5sCKWysnZ/H8Ym0Af0gV768J5NrfwPaTVESPE3
hox0OGhcFFvSCVepl6M86iFTVOVjb4tyXZlPWpT6Kh9mFw44YcFs8A1bj+NJGR4vVy+utVAn+9jp
HSTBCbBAO0Nd++l7h2ECl4YQxj6rIGq908qTfXqblV2wOU1p/RUEk9ifXfU8atggtX9iTPGxuQle
2BqGs6PhxxDbo/2eaMSj5rPIQZAX/ZHo8oVUe0RK/tDNt0hTAk5XZuciwH3axrVAMM8F3/JgBvmh
ee+6eOclWSoyXNJ7BDY4KXaShOgZESrotHlSVvvyX3PzdDfRh03f4UYTN/C5ezjbS6oGPW4aKsrc
MgfOiFgtzorq0PIDSg9znqONeYGp1Qp8WuNNQSOi9FhiUvmNvqqZSzxMAgn5zerBelqM/zMeybsL
LRWSS3xgK8SeTIXZvygRD/FX3ao+TMTdr9QLHwhkjRM1czpKt8FFxQ4VaSzoutMOaMXDreI+XU+3
qRMMMBa+AxnxF8R3JzGxDQJFhTURnbh6bV8wvcT4biL8SK6jMNGVPyBspw9Dq8yIp0n1cyUoAf5a
r76ny5d9jDvdcG5uFPQP02yNKzZfBQ5GtObAC3moTZCIWEMshgJEOEKmmZtxI0OFtlLCbwLPjlSA
YfakZfV2Cd/ouaZOF45RDFHhYq4ngei7oYIlDcuPY6zILQLimtTMkmxuo7TEjt6kcAB8H+Uui49T
guT5wwsQe7vglM5s2Ut8XtZS+ddVsVgM4bROVxZy7Cz3zy+NbPauOZg2OUCTWZC9VdJ80mJcXDvw
xxMJlY62E2QA4kJEzHp2HtXnz6KGl+7dIAK4d9NCAApdSVkD5UyNYtOm6k8bHxBeBeeBFxe0Gzad
rUbHQ5eDLfXsirUmRThh/QmoU8IB53MsB51jbVmJJJ87j02qa036+LUbBHZei1wWD/fiLjcXW+b+
eeLoXltlPbf0r7h9fW0VAvYMTnOCNbBS3uN2Jhss9hP35l3DZ+yMTAGnoVE4AVLH18rSkgAPfDzO
vHpB/+iqHjZRaBqOcyFGEdhB8KFK9lSicCoiPT0L1c5u02jjPn2Za42AstXnsU8jl4FXxEPcQlYg
al3KB4kEiyQ4zLl7bwb5FStX5Bn9gF7pBqY74ON0q9nPWuG4Or162i3buFTadaXW2eOrjN6j4bEc
t77W/+M4DPnPHHJ80nay7R0J7OrtfN8QQPhwNaMsdMN/FDxxttSDC7ppEVKJRH/r7iPtXpzpCzZn
fnvV5GRKq0+EMhu+9KZR10tV/tZmlc3P7ullvnB9Wq4sT+lUckJzCP43vqLUHMP8jtS4lbpe4GrN
IqSM6+k/l/lG26NXkMxPYsFvjXD5aTVderAhsZkMazhlvAvT2p5eTZuEsmLC9g5MSzs2gP4MfREY
cTMbUQEm6PF5uVM39xibGPJ2sB4z/VYYAJtrZo9vSJdLXVxOexgyKpOnffftkD+pNKdj/vKT86sE
K9vsUiigFkd7pf3ZUD2g9j/aqtKl+eiij8WNzy7UaxL1+XDN87uUPPWYv3ZJY2BYczQLIRo/Tej5
2jRlFOy6lmBGZtjDZSwcG0s+qkrtLcvuMEN8lof34zyOej3eCRRN54eAL8jilaTBIHv944/B9Qff
8cIi/jAFA3r7P3vTG8xL4xgx2nvfZqT+FVidWuaXJJVXsZy24mZJQd5jA9p56pKft8w6oo86nl2S
ajVPS97Osgpm3vhAyHlIcAe9MjDBmMi+iefnPmCO2piIgm4gCj96c+XexDiRetTLiM2k8tKoWXQl
Rs3wtvdvWPbeODQEluKVpOlPHOKbyglVF/Mip/N3gtEo1iPsRTnPEDfoFX1pU4AtvKEg8PhmNByb
kPHOT7M8k2Qpf6MwK3Abc1YwzGBw4/rnx+NxHa+6f3sQVrpo5s3St0Z4UsEUWiiri4YNFd9DrzMr
pVvLHeAIBeDem+UD7MS58Qgbc+zw4FLoYFyYoSUjZZRfsuhr/tXfjNo9SSRCIfUmJ5qAcBn2jndj
2vFlVGuXjwPGUPj8IjUizgWQnxW9fUzzoT86FabT7CqR2eL1nc9i7RXF4aeBLlG8Dqf0j04nlHUx
ROPRhxJD7j+vC7SDsCMe1PU+fwfNmIcOanqMhxUMYg5Iny4Am3/AruvwCToFcJ9pWqR/2EwIiGAH
QzEAU5bs/A2MalstYJUhdIG/0Nz04Yc9+Xvnjcudv31fJtYHi0K988iZwIiIWywYtwHkKha6BXjU
ftq7IC2ieuWMNMokegk5Frqez2EqPHcZ00S1RAQZLTgS9tliH+GPP4FIy+YLd81/G4xCj7h2pZV9
h7MCGFJE9wHwzr6O0qURGMeYFwdqbPm1r58e/Nov7VKLUihoRC78LSvdbGZ7s0Il/mXMNRFUvCKu
USgjc9s0kqZMcyAEdbbjNRg+GTjI+0HgETtE4DSVhXHeXnhWJgp8mlgmKWEQm7qytWltJFGwVp5T
x1wZv8k1tWI/cjIpZxsq8IT18ICkCDiBqmmXE4lZtGu8Ch4dFvfXdwIUsbDuIvDtrcJMAYRuxjcX
QIdukw/bOB5vDPHQaEFijV/tufxbL8y2c5ZTCH1pTeZZZsBNlbHmBxQjZsjLIdiki1kCXhlLNzta
jJWVgCrJhChYZO8+qNPSjsmWdF2quekFzebTmQM0IKSZvzotZ+S3ZwlM061Vl9qyTZMHuajw3Qw9
wa8YUgpQk0FmUHiKMyv3qATJb3NQc5ULqSmSJU3ALf1/Dm2rivIDP3C1swtG1arm50ohehPdVH/d
LLbfKIA6moI7vbG9atY8Aea7fmRF5Vme0Yo02Kn94Uz9RCMx5bd//dLHIZZzDD9z0AMCg6tHQkWj
JfPKfjruxqXhqhtAJNk1a9ne31U5swizlCRbwFHH3CfSOIHgUyezSH6X5VDdsf39NlaO+pkzZZmg
1sx0W7v+NOqts3M3VZeaSdI9yYblM1bEHtZMlJBAGjv/JW1fN14poi8oLaVz/ZzeVrAPHIO0M9tw
PnwZl/WE+LYrKUYNl9U7FcJ90lMak2LpeaOiuIH5DXKHXqP1ZghgGMMAlftcN3iQ7fk5jsSC2ZME
NltC6wSTr/Gww0P1EkFgAUziVvYBSSowLQ8NsOcer83gyoywAtzYfn/MRkYXtvrVPGUSgM+SJh1s
Btno/DiaDw+zBalHam98iMEE1jebEvbDZv+QZuPRHIHaZ3DN4qAgDyYX79LY3ZKxgovnwDVvKJpT
4wbV2PImg5LsVm2ScwaaNzweXGd23BA5XXeOAjD6sDDuUbqZprYzWDDfqLjcrx0lD2vcdAjejOX8
7IVTfyXhcBduCLdRCDElgspszHwawD3azdWoxdmgQoMuqrTqOj2rk2Yx259gRxFkmop/f9ZmOSqJ
g+YX6C+CqukTGofDHfp+vRtxv2jzq9hzWrG94GR3tWrFO5KDtzF/jN2hIPB/Wc6lgtNbJWIUuqi3
KaCkxdCFUeaKrDaQQYhsdVs6hYkLEnJ/5QlayFXYj8vkPlpraAWYeax1p9TC+LjmuE3ms8vdWkck
MK3CUhBhjzufYdqH7wXfhc4RdQ+FhvXXOEs/j9VYiIr4fxSY00K4l/Drtt9n5+o+0+9ERUpywKy/
/mDFrAr5XYYBYPpfqV4CrIsX2VN2CmacoxOwpFP9BbdOphjpvb+kjsrEAddWZmMA6cu60adfdYIc
NP/ylEtZLNotI6KvLv1xZaMk7NX9WaCNSEWuJvAxKk1cJ8dfQdugEzRgYQp5w7Y0LdDXfK573h2f
3dFXzIjwHQztUGm394H+pJUKwIZ7voRkR4pdNC5rbfg1TS5EKRqdgGK4pez2DFTB6IPYxBP/NBxp
lhgKZUbzesrxkzbCBNAIpWhwjImc2eCaI3YD/BMnlErnRpYXrUfnE1AVb917K+uZwtTHfRyxoWu1
x5/mIx9MZuqwtPQj5JeNB++LT4bKOukFB15QDgOTkq79dh7puQ5G0AAP3XW9CvcLM27SSSPHIInW
jPB4rpQYOI/Rt2wVnziSKGlN1IqtB80Srl2eYyxknBU0v9kX9b83dOSDWfky+KyUQoAOEUZaG2AI
VavY0w2iIN44nx/IAoDEE1xS+MRKbZgUOsK2sRY3yxoBwDyXlvaxbruxfrkSIwv2LIRP1ciG8IOZ
Rsqtc34YpRI6qsD+Py+Jo91QROuxLoHSTCaRbE2zn3Q7Cbb2PJgvqAs/zr/y5WfaJjyhlqLUfuIf
1bLUFGsxWYFfSBlkYMZF1Qqgk1khCeTcESxeYwtpl+bPw1xyxl/kPotMbZg66QIFEECl/8+2Iw96
pDQtrkDHdA4IcQSSS5rOT9TMrTmv0ZPRKMbScDztSLWSmRAxcfKZ7SlAq1Zp8VZPycIWnaelv62L
dZkfV7QYRhiWtFq/XCoAMp7Q7Qol1hnzCwuQK7NxlumgvIAnG2l+ABzPee+OxVaXi/6hX2Nmnpq8
TcCso22IRtn3/dWS8Zs0skfo2DwLe56rQpcLcL4/A4IKv6N04IS/2nkZ33CjtoE+41Z+o4KpX9bN
DALaDNDGJ7ehaesP1wzO+ORhfenX4x0KL6Hy6ASlbnF2X/ixrnqdfllSqxcH13BbgPo4K0PssYm4
jAiZi3Rf6F4d2A6j2VEMhv15SHSRAgmYybPeBal0zlpp8lkbWNOsN7XgsnqHPrZwd88f3zJuSb0a
ji1qEz3EIw1wn2yoQdgOl7Du8RXgRK5+5X/BwKI2po+Qv6EuEeLUun99BhdSpGX924RnYUX26ZFn
J78f6EY+no3uxg9KqGRw7ir5A8HE5wBleCcWJry/ST10aT1+2ZQbE/+iJ+3j8apm7JAajVolQwns
KN1HP3ShE4IFdFBDkauYAaF4KY0YunqNjXk3pC5H/wlqRKjI6aqrI/cgj3q2FP5gs1OTwxgvpqjX
LQbQqTv+fuaNQpQDxAhQwDZIjKzuyDsFaLTPfODqNMHaDEZhjv7bx81HSwW99mW9FYqpSIYfrQXA
bMCCuMn13eDL2gWuAkclux3fl3sGygpsYP+qHtJDe0ianzeIeW3puKjsWMrNhnqE7r5JscLrT+ki
4CLvMkIkaZhWOfLTyWvTllDMZebg6lg4DfrRlE2i+ULppgm6ES+39QIyB/2jN/wngk+Pn9ZiLRgQ
p/FZGPDTICX+dldPN0P0drQ/Q1SJgub8D2mDGwkfMrqwIlwELJveyygz6gvXIEoyqIT7QMZsdgYA
po2uFchUAebvrSdq+tUoyxDDMUBV2yuKIANofoBBIzAZl+eMUuvCYaZI6K0eehIjhRC8SPDqXEGU
7+Ht8NNv+/nyF3AsvhQY+dxpuquNDf0X0pbku+CKDigSq9zG+mDmA4N7uTMjFt/p1YC4jdNIavuS
nsoP+RK+TR2avqOpLtdEYh7HHY5p3ASKycgwUOUfGPBnN9dJAbFUkScSqxDvnB6cASQnrKZ3vXTb
n6jizPIeCFWOERySJ7VKtFGGzsjbUEq8WqfGMOks9WJDdY0boV2VBtrR3cynzGDqZVnsOdfSbjcZ
9VwhnC9zSWEfS/7DM2lCmJxFD+WnGAfsNGZRHClR7Z5+vrpZFf3vsAWMBxUchdkGqVCsvZcqfm/r
+akUCth1gIF0Qrpl4TO0dtwL2hwd8MHiJY/qeH0uPoQ8UGbgbQvyOBzDUw2UHfIjYykuUy2mz7RC
i4DbzFK+G0g3wnxpwxrK/VQyUx99R7kVM2Ri615grgG2UfBKQzJPaFlKLsTEYLZUcQQ/ekYS0tP0
82k+ZETkCO/nw689iOvzw1rXrmUQVoJ8KZf3lr1/nc97GISIQf/ArxhD5u8w4rCyTtjNOghWXfeE
S2Xcg6ttZrlx31cHuwf8tfdFx9J7DG0rnI6lMN82/rxGK2XjucPqV2q+YWTsoxFLBj3BRvWtvT9E
LBxGMz88TW620h2Ar6e1aaQCQLVk20ZqMvMpCJAH9hdokY+6SO8rVS2FLgL/0thX4T3nQnuD9e12
94eJe2GybT4aWaGGhGlZqgNg6pcSJAyCMUqzGGSWiwoQFZJWzyEEzn6hk+RUMpUHNY2BdOzd/ADt
XC+NGoX3HQTQiwm61g0Kh2pq0o8+VQlJcruW+M2WfvBqPxD8enP3xmxmAEKFmsAoWh6lprvhBU4H
ufRoelAWQrrqKUjxE0KDgBIZouVxz4gQM8VRZWQFXdAlEkJmwoRWqT/1wakNoQC0XHNDGfbfljny
Esjh0dN0MSKJujoFHHzF08uvvg1JWCiz8/pbqzXTFzWQwxIl7IsJt6r2iOHNhR4sGTOSCCssMHzK
iS2ev2cNATpFhDhtDyWgkNubrPeieNOQFWqiCiUdRut1jd7rQaJcpqUN1JwRHZr9bBvkMrKaEcl3
PGTV0oSQdXKKd5zp117IPq08gPJtjqc58Dv5EnJD4PA7Gen0LyeephOpG9w0bU1togCK8Vw7oV/X
uXJEk/uNXuJ+eYIdJAx8t1N9mX+gyvn7t1UW0saIxQzii2BXljeCIo3ewpNoS0BmkjuxzPMxRsK/
2MAXyMJCPDum0DfYQzWh1wXIfKmxxnCvznmHoX7AFhzx2tmOL886NrRrIB/fnllTi7S7ZBodCQuh
6viO2uZLeqOiiGxpHKiK3IcJSqb+YVb8G0yY3FphNbAstwuRjP1AI+Bk01mx4TVW4L8bzNEH4nKU
k52vS4gADc6NnBXbk8Op55nkMNGbxTFf0/kzan7fOu1aji8EymSt/VfLhIUmM2zTFXkUd3al1SbL
OWpISInawxKLcFsITI4DTn6jaqSHvPmjWrKGMl8FGEfr0lcGajljLwjucuBE5aori2btTcWweJLX
TX1asC5KDF61gmVN8pKKf6GeN2irQdOJwn5SpMCIQaxAAgHLwNQufrlgkWtt5uHILTCkDrG6SAPk
4j/37Do/s2ADNQvz0glF8xZvRcu8jUhH723fnL/oE5cMGh+U2IQOnsl4zw4kciCfO2ZOpbnXMNn9
yfJa+g8Crd+plQoAcJKaO5ilxNT/FeqA0Q+L0nDTyhjDR/28gH/FxLii6E+Ch0huxkfD2TnNooe7
DAszd4lIQ03wTVpmY313ByrWmwZ0l0IHNJ1nwHc7GuLm6twi4G2qTraRS66wzqVsvw5wwa1zMtd0
fUz0l+m9M7bup389Ac2g0fi8nY4yh1pxXi/a6XtpLBfDMQeQiA37raNdPNwHJEUMaNInOi2XOEJx
Agrvf+hQTv1Mm5vYUF1vz3r0DqjHL+6X5akPIiFmNX1EC0IOjlODh642JHyMbcNHXeA7IOa/vtc7
3aGq2suZHsfWnkYhMSIIfgcMdl/56fgfKhDoHKJgOYcnjb0OpvC4tBuk7flfVFNs15Xy4rQ/iSIa
oFqz3u/JqmwGMf3J/9L6ND+bHbbANpZCPuJWxNgYQJhh+JojPpXZOJ8fpp0UBn23U+BgmE6ZOYVw
WO837uXBteTkcG16StlP93HXHfeb8yncRoS4eYfXmz2VmfVe7Je3I24UiHoYLz2sNglEx19vnn/J
LZDCq6/yu+3SvIX8G3hHlyrBCQViQInwLlMp5KJ5GXmy62WlwOATJvRSQOwrv0DZ5g3vF4QMKHTx
leZatdnbPQoTul4csejxpBZOAe0bEQObYli0mHFjQDOIbv49Yvhr93F8DlNJW1IumZdtwcmEnaJj
G9loahnxYdjvP8V1NFJOWP4cLE28WUzdzt6sCz4s39IEA34PYmleikIwCpSXJN4gt+8ebYXX79gC
IPFNfMChfXtcYDJF5HVi+taWACzPaLZNDE8xDFEP1gq+MmKtbHVjpqc3dfn1iWPOZHBpd6R/5t4v
ziyKgDmDeI3enSJdJPpkqI24fZ03U2rhAsz9qYmTi19lVq3QLb5RzYqTRRHazAgNvDyAMiNAt8Jo
EG52M/96TxQcVMjgL/gWdgQBX6eCg6m3YJSqoDWBEAW5ngSLCN6chhvuHzllTe2TVFAa1i9btyY4
Qs19oBW/vBQR/WujkDBpvvoRHPGgTVUEaY2fjJk+YcIx9/NZthuwDyaIrfYT/heiQWP+d52l5mvX
QbZ+ErzkDIsS7dbIfgbwdqbYX3EC/ppfewwMRP6wCcNBmoE5deorqCtPdYKQ8NM/+bEEDRtkrUsG
xicJva/2vDCrZ/k3Ib1hwOjzNltwAJcyBRWwmCRltcQ7bPQnueo7nEHPBIqXb6Gs56aiETMMhOk3
kdBdhfmIq4ZdRPA6teU6Ol7KseXwaEKGN2AT9N22xaWmhqRKW4a00GL08/i9896zDg1UinjVG3Mx
vhgmkPzQdUt+aeWhGwghN2uFE6K33fwH1lgCBeIr5blDO4w1uZfFicgoNkua/XAfMFat14LGivrw
BcKTGHJS8j9BDW1lNI6HOUTwkM00zFtcnla/VKS1NA90YlvebSCWAGs/oQin/AJ1sS3YmKzPnTxZ
Ln7q++0lbY3W9L18kvO9Vju+hySQ7OZ6bNiLulO5UwzoZT6YanFyGDw5QNkgrcAMOc79tBqbAwUv
qDGhsnQu4J+81S6BuLNySd/sBwZ8hCgz6yzbX7zF5/BCF56KBPvZFQyiSAhjmPD6F6/cd4DsNtXz
J/tTDrfE//2O6LDimLaqbnSj9ZXoSqwvpDPbKYl7ZXdiETO7DVdUouLnGrl2QGC+BVi60LsSlofm
XOToTAojXnT5YCa/PSVg/s2x9J6kPf1IJWpNYjqB0XszFrhCOXRH7sfyY6lVXgA8a86CrV2ZVhcd
1i8F/SiRo4vpiRhDi5PCimvKdGcIq7SSVKC4vXh6pBs3L0iOlCgUXT59LG567xuJjQKixtb4dwQv
b/MYUTMpbDfxkOcIWhRW0tgj6Hh6HN1loUc5yigRxwkrgo73wWkDaSrN5R6izuOrN+kRWbtgT3qN
qPjwnQXl4Aur1hespiV7078fRDkQcg/2y6qPmdP3eVkdfEpzkJdJb3mKRz0RfYrQj308HSr2gIRH
FMz2HCo/wGUukDYlOjcDXyvfp6bhpC7QtlPNyjWj1UtP0J/fZi+2RNR9l4w+WRW83WUzPlVB3J2S
IWGwHWGs7zx+u/H71ce2761w36QnXnAu0bGLpYBuNRSSsmkKoO2VNGiGS2Jso2HHJ8MU6dN7/Kxl
J2MNphAcH89dwQsHnSc+SJHUQ5nLPZMnMaTvQ4pObfk6RIp+01tBnfv9qfTQKNVxNImC/o1VLtE4
8t6eRRFm+1Y1PHqpYR42nAbln8LWfoqkDTGnUphcX33KTgLCzjsrd+aSZt8gVwxD3C9K3ylSVcUm
CuN6cX7RA13BRYSTBoTKfD+E9Na0Q0r/vbk7lX9certwnwwUjXitr81LFPgTpW1ZBFlAuvXVLsBc
gbI805RrtChCxekm79L3Q7Ubux00MatEOVu142t0PnJjOvLo9o98MbttiKLm20JjYCja6EKzGApX
VMylP3a8wnYIOj0XOvmYZ+76Eig/v3OSaTEJrDbNmh6Dyk+Ea7xT121TI0NfKuv6LOb4T2gAEy2D
m7zA7FkIzf2ppp/8BwFK3rDj+nzk+0/KE7yP67j2AcLGUDvLRFfUM5esC2V36tbtngkQEaXhD1wu
qex24+s1gxDiDkJkpQh9TFR6mJcXlC6756DifFAl1Z1oExbrFoWAasa52UvibORdZqB53JrRs+Fy
XMIWqnc1jqraU6DY96sYwBwD3y7rWeoEUy/rTkEvEFMForc9aBN4/G2aG65bvUq8jVtdxuYa6sp1
0vp9uyhqnGGzZPDbjjsPTFTuFCMCCiGuqCOiSd0YWgMvhiCDx07TvWR5tqtRotUQ/TysvalM/CKR
62Ode1SjxjiSwvYlGdR7qC/zq1wxfEk3Vap8guUGG6DmBDDW/B18Smr0izBYoYObbrgCucXnmtrD
Zz6Uz8WXUkJuvchdgV3Dy3teyaCFhsDR58q+2zfHl5BwM2+qYfp8A/Y+DlIoTlWYl2m3x6xQ5s4W
yi8NsHjFMVAOtv1PRmCUrkwYbMd9cKoQkzWPPNVXEm0pLJKEi2AqCEChtAXR7afUttLkh66OEPdB
IVCPi18Sl+syW42uo219e2EF/V0WYY+2ndj4+KVw/O1FwNNUUjBkzo85xEaE28vAl8nSNRLh9wT8
wyYuaeGKONpvc9jhUtF1Ho5R7AIP+MonhBbzW7/J1utY16i3UMioaHxYeFzEkDgtYpMaPO8kzezS
UGd1s/XsP8LpZkNXsF5P4ezesgHnwp2ERNNA0rYKVnR6kzKHS7QcVEfCiXBm2ZXuqgTQgr1CTwBk
1DiD057NatlDKIIR+KzG6tUdQXwDLxGPNaNB0BOKmyvLc93Mam9tPOVN2R55Om0bNG1pn/To0THj
WbtMy/yGQMYSEbaiq1vXs3F2cLR+ReNiUDhS0nl3uQAyZOAXfJz1ZUG9VjF92w1qCRJT9zWvZtAz
vFQtvwmzN/hP46zkKpm2+FoJn0WK6UAjmXd7Q2lozkeKj6vX884v83f66K78sVi2BsImXzbXXXR1
jZUD1Gvy5dyknJ5IwvXHeKSHvt1QFQuMT2L+yTd6TZL4Cl06RteVekFrtA0G0Uhdt+AXAFTqUE9a
/48MWTCRk67J9gQdkbE1W85wqoqep73TBUsn8oYMgQxOuX67lWh1MQ/RwcXv5SW0tZG5mMomUr7G
UqMAVXymA5FPu6qd1YjVejdYl9bNy/ZxDeSKfCpDfA5bB4ATTQjA6GFosJVjGmI37EVHzXKNxu7l
xSfialInm5cvGdqe4Lc7FPEgJ3ag9pJfwH8nTT38LULYeOIi4iYsoV1PJ7LKRZBd2TK6v1Sn3qML
ko+WdHRcsHzQa5LnoFv6iNDlmJRtqKyB5tiS9B9x9koLud2J9VMoIX8c/FfoVu51d1nT+u+AEknP
I3T2rphqJtgH1c0BbZxbQYnxSQrKnGZhDR9WH3c5tKHdg6ETHKR6Anb0Wv2e2BhUydOBDdo6UTXj
wrvOfQ3dboNolscZYCq/6P4sEGAhTttryl6bQhZ08zyJrF1CB9p/qfHvLfwHXKyOqoplAnrSVKlc
4+lO8n23w5R04XKdnjU0wsC9md5r9vb+olJeJERyXvzzSs32EDTx72hQI8YYxAFp+rgPzTiqH+ll
8GTebBcQ9J+wqTzv9c4tEiKS1OipGcW8/g/OhWPOH3kvXmkPNFcQeck8y4IQHzdHXbWQJJk36sFH
FYFVa73dwqq9ekqTZoRzF23qXeNbzMYl2QE5JjsRs8FVZUwH376okd0g/xRkBwEv2UslVOHG7htS
e2NCalBfCYSMhdIkbx14U2+nrF4MvLrSMOzQ3gZD8lyFYQkl1kfXD3iXpHgvcnwMkCS7ZZyHAfYu
6t/uzMT5UF8Whn9raCJmswprToWJFqqlLPGuChiNQ3zvgyW3C+6RDJWukfgOG5Cq8m7VMnk4Q/gc
4Oz3rb+2FBhaxDV6hnjfqfiYMPr0DOvI2aGFiW+ZTaXMYGAPRac4OSRbUj/5ORPHe6pdcCW2T0mp
eZh1Ew81awtSGQitpeo4YQTIyEnZyYQ9lZKN3N/sF8aHmfjmtKJcTTj1eoR3XI4sn8cBQBB3Cxx/
OYYW8RYpcK2oNkB8NqAYAfctqVlCyneGXUGu7Qy2fJ/aItxQvYWe5ZwXbe7SopRr9k+O9KcuCsii
CYng5UjOPaRWCc2RnZ8JyTEc+0J7YMJBrFlps7PpBx1fEETj4JZqlLTZ4eEBGFswxd44NlzT7MyC
EQ973SLtcHgIGU+L8CDmn+0ehaKTo1F1EexPdQgSGKZ5T4LJClk/9IIY9GI1dexPU/NeJYQDTC2i
MwiNAuuFFI0pqVSaOYah10naL2NDEJzidBs46LHA2DLc/ThhKVdDoyABcklsdQVITAJtovS9cFfq
vNDo2LU/5Z2El3ES1/SCziN0GdPG2Kl98XFhhXHWN4kbn49q7GPqw2jJ0uShUeA26xEah2vF2MDy
IzefZtiwdiYNhIshMLU+03mS1ztOERf3vnIzIpjEsbLi/aUYWCmWvi62Nvjj4ybYcrPdB4paYXqY
RWF+kXbEyIXns7A1R7j5F86UYv511vu20o+zFaIYN+b2lNtXcb1TunMewb6ZIi3dXpTvOEm9AECU
YySN2k6h6sQPNSd3tvP1Fj7x957FOdObk7EdDcj9OnloBDdIs6t0zhp1Wgeo5+jKaFxaNcdbXFxm
dof44lJ1pXExxy3/ppuRs+kbaVkRiaZx1TA7Uhn55L2oxiQPckVXsqQ6up7EiFxxX+Vbb26sYj3l
MaMlLGHfSayAPhMjrfY/XoSu86Qtx7ldYVSNKspWpoN7/mep49HqqK+VrmOz15w8gHHJeZVEW01l
5pTDnPdZV/eWZXhNdTV3//y3IjaJVC03eadqaKBkjijenJbl4Hw+iGpGODqC6D1sHGyWUQ4GdP3A
aXjKUlcbbtiWWykkHVsvt/APAuxg6tRYMd4W0XVU18B6hAcklhBlqkiTnitqWM8NpSxhkDEvaQej
P2M4PqDAMonmgAzIJR0F5f/zPOtcJUNpMzBRThShFbHWyX2m8Thqb1uDKnB3NVRL+jwQZWvCLcnP
mjdQ1U7x5PPo6cfq/jvztVKg1rEW2FiqDWBJFtY6gYCJ5Xhoypn8ZtfaNU55HrBvks2JncDIqDic
SPzO1hG9fp6kbQOckcjT7lQnIoamos54mfH56hBUs8qE9+X8Gl1ABOd04Mk6bt9zYFsgIJesHOXx
H2fAARtW2SleA8SPWjcHj+hnjNJBrH1HDkLAnMp+/TalCz5opfPkJNl0S2zq9OkGu6igS+PxscPl
TaS3/VLIDdKj0oeBFA2jrOyAWZq1I1YuE2hcYlYZwgME8meoC3duoXTRBgjExtSlFr+lE7zR/aiF
+HqALolOc3bQZiVHBdXkCrUcX93dYTUFpUYCyKMDzD80rT+sz9trc9kRejqDH25poyA6uuna3KaQ
bCvKrnEZ/4Pnp5Lu3tol2zhFrzNVPOcRtqK96n2N4WOn0OOM88p94uOJt1xkqEFyOmbWIY61m2GL
JxoaBQg+aMMvYn7iUTHlmI8vTTvTnJcBvgOXfPGWIjyT1S2M7a1SX0/IdQU4m6SgFNlffTwh8Fio
QbrR94UF8PbC52WncgvCL1mfGswUNj8ArqoLzpnb4WKbyV/d/ro/TAK63MCBD3dhza4c27O+7kVI
1qqslwsnqHO7pFpLLzJRphUzdggeNXd8tzsUN+7f7R9qwDkkHAQU97waJAEhZ8X7+FiRa+KFJIAR
bbCuct7N/+zNzwPdzzXr+O1szz6yd2wXccwur2JmXIYO+TNcgiK6rYB8t0RNzp1tCIo7910uyvGG
Rx0fXXSuvIKR6W4bOfN+l2/6cYiqeYtO+nK/7hBqCEu/Q639fiJc5WSxMrm5rT7FO10wj8w5nL4i
h1LD2mFuVu0W81QdzrulR3JKYqFkfPwDK0J2eMlqcXbvB2byQCmqmfJyCo+YQtja4/0BlcFsaWH9
OE/HQMuMaql/dFQHiAh5pdmbEGYbvbHGB91V+rcgIbm+cO4mEw4SLEzHEQMF14acippAdQ8xR4F5
1ywdxRuZpU4aTAdcEzwyyMDo1OVdrWQKmFhk/G4hRHAt2OjDTRxZ959D37SYGyPXXue0UGHQYJ+w
4/XhwGEDkc+Ly2VxsIQfwT7gswF7M6CdbC5hk9dUkBXQxTkjAQIHlNk36QmcWUGc4A+P7WasC2A+
4CTNgjK9sHsTeLftfTnQyepfp++7aAwgIUcomvTnR46Xjg6Id3ficdl8+witM+Eda2ADdbSujw84
qsHFXBBlsfwpxC4M9Dt47MXZiFT3VT75t+u8KPklSpGoYKLabL2Zq2pQtEJpDYBQp3+AFot2CYPn
8kXnEqZDPEsORQ93Gqdoj3MHEzjaSvbJoZFiWTIg1HhzPuG7nlRj8eoU9S3QADtP6h2f+0MsRgfg
xAsnFgSDMF+bzW8bdY1biEIHqaaua0gp8u2CeDkAgfJyoEbqBNEI20Nt3OujHOWCKMFiAR7GcYsg
EKaYJFvzeUD3sAmTu/DE/WkOSpHrc8BspJiNQRhy0nbAtvKKv8TqjYzUc4UuTxWvGnzl6XjD8ycB
reIQNd3juqbgyR6cVZeio7wphSh70a3dEGCOhtS5yfYr8N1Sr8Me1hFBuzJrkDO60Or1uuJyQj3C
7HCD5PS0lnawrG9HK6EF6YbA+ZwyDkwvQ0PudLTfx19IeHwbmJN2GrYJjUau9xKe7lEMKBENWIsW
1gSUHPGarRH4VZhftvTaMdInyvFm+htoqOe595YePP/lGe3B4hItRqw9yw8/zJadjumgHYgynufl
iDNxVxWyd7Lo4kiSsPig9/yN+3/Du8EhfaQxM4YOMBij86gV0HuTDpikvcgCSTnZ8n4KCUnHYTVJ
ZAQQgsDRJDVro1mfnB74nZptKqhwXXGFtfFRwGreR1LYCtGjxFQPSFZMO7rsBzvH6BlKMzmQxhd3
JP53bkFfuQXqUsVxxlZtOOSZ/UqzCYCiE4FLfyaHgYDZ1HYluafbeYonFGM0kPI/dg+7HXibIEE3
I97n3BZPAJTgQl/910TdNSdmZ/PEz1Uy7d+WTLyIDtuwLZzhjT+HLQnOJVWUhGeQyngiRWYdCSUA
Vumdp6+MX2dzvnj2PhgYjlMECBUgResTzD2+bgA1TqKKmgTqyvBVpH/Q4JVovvT2uJ4vb1BfqN+K
fs4p0kuR6lCkApXpo56D58EDDlvtMQmGCiIhY53snYL9X7RDMxNUFSYCK186IANcZEEVs3LsgAmJ
iNIzgzFalBLioYRuezkZg2VFcaMfbSo67wnqUHpnCL3pi3rVKx8tVsV5yxmQ0azUw3zbQn9eyQ+W
PifNOg6ScKvGWdfpviu+WM6cG6/TILrhGG8FezDrj/FofT1cl0tuyLZXrm3+6+im9WpjQXzKI4Q2
07jMwwKYiok136vvKCnFo5ongdbNZZKe0GJtSVqlYOHrhu5/D2rA/PHO8+soeAs000+okt476sMG
UxsGHSsgUa1w7T5T7kcAfOJTR103rQqkPHsWElmTBdXfvd0HXm/yHbA0WValx+3BvyP2LnSxGeQD
ffT596p4mpBgW/dbxNgCWqe0X/6WWR9vx9OfZZxikqkGlTUuCoEntKjM2+DtCvPwSLyDK+NXGJuU
nPUoYzz3JCC2DOEh3CX0QbPxVI+AqTEdfiQPN+s1V14GYsca/H82LFRLcO6h8IRkk8fp4cp37zQM
HuXWpnz2HQgPQA/0D82i/QUVvtCgczW0KqbVUM8Av5zA14x5ju/v2n7oPLvMrN9fYkRDJsGKa2HL
9dwVrb2hUwYMIpkYi9BjV41fsWoQIV5SlTge2g2/wdan3nbPnwMr3KC58r4NKAKgxXNQQcZ44Lmv
nwHxtjOIRRn8BlR0DKQgFbpTdt5A7dsNjK2KIVdel2Jd9KnFVDTyeWsr3P6UPfuWXViPo5tyvYJ1
mCrnCV/z6mh10qKUwrS0r4og/AorA9bM1opA3WJ0UUo53ap2hyO9TbClwpYBsWgks8vwanByoZCw
1fkMed61RBEX68RBZne5Gy83U6zIpYiDEOwuPUToxmzHsvG+js1KkStiS80kILopuo6bcWJZz3uF
qee+3SRsxRnv0bnRFNT8KwOoUnUVNSMc/j4zZqsi9TDx4mOHNpyYVc5s19MBQsJ2I/CDPvBYsnjL
Kw/YxUYJza4Bzf1KgcRIsgYoE6YWx47KqEFz/HXmm9r8D4ZuzthiRbPAd71hGxJ+VL9pWuIVajRC
DNfzDkdSUxYlX1YpnSolAHVmQdBUPY3ztZrw25FL09NymOSi8PXaBjo8gvkOARjSdZxunUKzBHm6
+y0sjMVSVaH63L95mxhljl9KtSulcRwPxAxm6Q5WCNheHujIPMc5MLrCYeGw5iE9Nd4lutvA8Ei9
AlvJzFKagAwmjJ7mIhsj0oOEnmnjeHY+emF2Ckv/jfP9Go1rGw8puDL9EyaTts+giSy3d7ghDHaH
DUyLsSdI51C8wERnRxK5ftj7+XEAGjHTIkNjxEJPAtA1TyNHrvPeG4dJwpZ7k1RoyV2BPuI1DVab
zrAI/JojvUVaFjitMxhkNk6PqGrdnfxR5LwCz7S1kU3JKsrHddapmUXXA640PAKuIDYzXrqhJ41/
KJ5dgI/ijvOOVXbRxJv0veH5PlzXX6XewCc3os5cyGsejQNAxQYeCTcJRbNpkW+cR7egFiUEiT2O
lKFkll0MlbtpPoNS2sditLtidBH/308fjIJLKB3o58PSb/QWcc870eErfUfpsJqrWqnnBy4358G/
P0zeSP2fDi2dxtm7bEGRaeiI0fVjpgiL0XtAH8UNpbEFPxR0sPWD/Fh3Mw6+Z9f+j6D7kqt1Ax4u
5AbItZ0L+vqleCjauNjRcEwA7t6lAHDoae5Ef1chyEY7BqI7UAzCLMFTSNfG2zuREjlgp6C7LjUg
IVFYTu1r2FnfoL5CIkU01Aqd667L8S5QkYnmfrZq37mtRWH1/Gx5d5lsdKe4SYlpQinAXxxsO1F9
zPYXVEMUxkRh3UejEjwhqXxQOPdWm7AyxBXmnTH8iDpqTFMajXbDKRd3Fb5FgqpNUgo99rZ3GM8p
aW70FQn0X1rgfGE6x4C6ttpztJIoo81WqmK4I/nd1SbND/igCifmyIomwGQIGePZP6mQADdTW56P
I5CHOh65avzEaDZSIC4us3e0crsmiMBac31W08xSo7P0JNkmCpP9wy1rLAKLEDxuuRXMRkj8L6aD
+UTdKuOjeiB+Nx/o0+ODSTJ2t184TGVm/Uo+VuF2pk30V+12z4pzHvCLGcQHX8PJVwbGx1V6AHsl
ipyzJrItuIlMu6ZOSHwF5+4i0DEN5ddLAAR0LYoJ/hYZ5naCPzJXho3ca2S9Xmc6GrMiCzrD05sq
pHdwryV9Tk6FMc5rs814q72e14k4PJoo+/ReaJHIRUiHFUhXEK/aQR2MManJXu+voi+eeAp9ffQF
SeIZLLB7G5hby6ZQ5E/nV9Ti7TfcrJO5csvtQKBfWwrOG/OJcYplXr7yrwcLSZJ180IkVsca4JWB
DVoC4FIKNgwjjzVulkI7HHDVGx4D0enxotJXpgilxLvOdQWq/3tnnzyVMrOY10WyIFVaGrVJ+DcN
a+fw5sWgnjoTTSpk/nzyko3eG/jqDQz+HekhVKr6cbeTFUI64P4RNDyNeG+EXKNVrUwXjlrhVGtb
uyZWJ24RM4E/NYA4JBxByGxTE2yg114zgHosU5bP/eiyJiZrLiiTTyz9UH9Idm0dEZiSQrgNkWZ9
oN+aFfZokS4IKpN9caxRvsBCZXKc//IwWUAlKm9Da3WvoZ92cBRaqpURsLitcghwU54IKmKAxh6m
1q8kzHprSP9vuEdYoEKK52nrwNvWspUrgrMOyvespH+91Phq2wBYEYY1CQOHno2VbcYePKHX8ksg
D/uLeljf7Yi8UPgtdstRq1WOsOSHtjRSiTXc6W6HYwjVZaeE35YkiqPlKnreinKHt3VANX5PcPRo
g8hF5gT0XiSzpma+S3Sgl8+NXbwjI138RDErIGw9NoItdsGUwS/rtRidiqzkFp+M2apAYLKdFgmf
TIB9pjD9XGYkHxKn+nc/1Rp8OEMzgIU5w7ClXMm5JQjQWtZGS2bTet4989tkA1EomOhuelMFHVKu
01QkJq80w/IyJRuO/1UgiC7FAk3wyzr15KGgp9IFpcH3wxJOu9uKMd+NIf0hwOEi19Ln6JspsAmE
0e2UA3ho16CLrN3qov8u8BKx8Az4N+MtaD/eldEHIqNVWIOIwqpH3if4Z83gBYHuwHeHtvXCblw6
J8UivNSHnJiCrblKx9HbRxl7lMsbqvOLuaSDvMeL4476LPTuBxOb2qjEjFkRs9SNRvqcagNmbISc
4TqEJcq2vSbg0L0eU0g9U/nkSiw6bcAFl1HHYzrWFmLk+BjcdJzjYJeu7WhrUHbTk5RfNm+kyKYO
IutATICrWvK7A0WPZRplooe82f6JF8H1bANwhpsneygd/Nj90QNGVLys7C3hxYTfcuhpPEY0868E
0aCDIRXHU4TE0aOFHVrbA3bNty0uaykCYilwzCAgTpmu/8yXLE8kOOS6WY4AbhtapU8QSIYHrNhR
PG7+VJGcQS8Om643ERxle4ygtLOM5LRTkoVma5gqhgDy2eQ6IUXu3KKIUUdOFljv3XjQyjKTlgm3
s9o4IDiEJrwBHJuDBm3oDp4D8amrjPB0tHh3Vv/PNaBjMLdKTlM/lyJqlkDK6GzxuuHm7dfr48AI
rxsuNu4iLNeq7uIWpwzksJYa32Dyv2W2oefoXR07c8CbJfLksJY9xQcsfFYjWe0XsOBGM04ilGFI
u9ctc8XVk+wlPA7oIcJA01R8EHq+FBIKGEG43w4f6RByxXClWvFr7i1EabfNKG/bJbpPU8UayPKz
vMIAX9tJgzzYdPBBgIzGp8fZ0aYT1Ue4HtdASjW2UmrffwxerS1iXmOk7NmfA+8vnn0ZsZwqao/c
gnMbWqDlls1YKI/D1/OI4kkyMlFF3o4z1FtxQq8VqlM+Rd9Zsu0u9WXfQ/VfLERlpPbsUwV8yCt1
KlZm6gsf7roJejIofahH2C3t29iAVr9PpnvGA6ZPdv3msLFx+ThNYLzFYBSqew6rLoxnlIp1rAEb
Y84XtbcFCJIvZq5W1KdW/y55XUQQYn1bRiHNNc/HwuqGNrHuVpH9/kzIGVS0sQnbH07laAIBl8gQ
X1WymupeOk4BAom1Yp4kyOrkWh0H5cTZZEfrXfmIIL2T0S28+IZb5QIqM6TXuBSoFPKPX4BS7MkD
yj34koa3k/pNMbueSXzvLPdr+/UjZ4EfItHCkaWSTXFJKn8Ry9S+40DbQdHh7VvTba5YMuu5OZN5
vnN+lVVIw6IcBhlqIKOwIBntxlnHiERYpsHP58HLNIo25aZx5IYhiOOgOE+Dtfqex5E8T+fDnMfe
gE5Q7c8IHDtLMGp3gZXQHNcCfJP02nv750bMMsBE+0X1zndsZMyHeX0+F4WM44q6y0Av1/2fPLCS
yMLqdl1a3XXjwCdalkzuW3HOLS6z6Zc7rVNekpZZ9hfFWzuH9BMey0k2ytVxnXN5w7RIbSrp6BXq
fSJ8WiD1D9bmHWzdqJnDL1eu31iL061zMljMaIZS9igQSxebEZ5W7tBUVERTUZVAUoNzAg3DLW13
kp/2jzQPoKLUODw1jcPWk7xrUPyRR1iwYyXdAWYwpWMsaQlwzf2Lv9EmLRLiPQ7GEyLXZdjkNL5L
cQ2lgyWmUr1GieK6YvhYPP/Oq0D7ZeDfueISh40U8/kJXCJSgTq11MajwkHJOL2b9guDCh+iy7KW
+ucEXX74LI2MCW3A5JYy8eSJ/vomRRM8wEYQVabUqllDv0Apag4N6R4Fzt/LiS4pnRRgRwTb+f2k
1oEKEJTNkBR87Um+SFrvKohYFqoCB/XIO5bXyFkOmC/suRSWIwS1GK4tD5dgM3ZYZd8Fv88njxty
fzR2dQ9LsbfJlDibBlY3DmpqFjs8HA4sCN8Cq9ZTHqC1E1UPe9qvj6leszv4PPAqK7I4M9IxAk8k
dyLxtxJYOUWEIH1AKYSVG9PFsEoiW+Vl0trUaClKefFosVVXMq10hR409O2BTHiscxZ616YTfgfQ
cq1RRB5nNU3wkFQmMkvdejp3GQIdD2wU04Czvahds5RYH3i63eCHGmUGZajbAnAOe89+m3jYxskx
9gv/8Pi9r4ZjxLBf7QH3asLYtsBYT4VQklr39fTqYaFYyA1I4dLxHCfpZ/SqPCKRKgiSe8VNUQjC
6tzrdhseS0vVoR0JtdIxur+6J7P3YL0912sPRx+GaxICwRRazna8APrTNtL+f2pcEYJyYl8BhaQi
fR+x9RwUW+O8dxpVAKpaeFEoW2i9lCBIg4Uwj79h9bW4lWSMclH4ZymvYaNKO5ss5Xe+J2hW8uYS
8JkzDX8vdN5Bcj8wKPXAFSkS74tZrxymvqHoAH0xyMJJC6WIk/Xvw7LE23t6rppAcocY2Yk9iHyi
8hYGjdoc0yFYWc8XdvoCjn5GCtcIPy7mBrla8g21e3AhdWNior+MuqvzTxyGBTIfhdaZ6V1CZhYF
Q5Z9yB1d5Guz9iCFc6wgdeclKG/aW7SqUPAYpxMi4qUQ1a9vNRgE3ODaaNEA1N3NtU4/ftClE1+2
jftlQXOU2qBiBy5T3Fo3HjClOCk8mKZsHnRycAbeJQCStjk77SxswK+XkyGctl3AjEPeofxGf9K/
GTlxwsKEjcIpRG4Q23YDkNhkpP6dCGOwIQkQzw+JDm7ko1Ts2I95hpLkyZEmQ2dkyk6NuoT+4trY
RCrXnjwJ7/AR7ESfGriN0sCR56h7j7ShL0VSPyqda5K+l8zx0egZ+Sl/4+iZ0erfJC90WKeogctG
o5+/+c6wa8uUknDTEAJ8pVgkFqKhpBtXt5inx4hCvklfghxBX4FGJ62upN0PxU6PgHfzx0aUd4ep
iZ949pdS50x+kwyi+yKAxcOD0ZUt/ttetvdJrla4lGQPR2LfuXielx0W1hAvt/IcZ4wc4x1Mx13h
KHGkpXrd4ADnnW4DY6FUjz6dvUib5Cs+O27BPTJbZylqKiYmmoPY8A1Upksqq/JmAHdsW6GnS/r9
u32MNY/q4U81gHmwSEdp1ubLUwzM+7UNzuBMQ5tAetFGWEllpa3dVs0oPq3/9P3wR5NnLTPN2HJv
ChgiH/Z9IhU992zzQpcydJJ7zJ0+4iNNMeHdEIfBMuadLIZrYCHVAjwwnKhAExK4zlZsX3ZC44xf
WqST18+Pilmm3w7UA69Qjq4gd9VJecZRsr2qE0gaJfLgq9t3kFwwYJt/CgO0bhy5BK7MYaW7x6S6
UPFTFz5J6JmM23WJ7ZNTRk3ojh7GN/9rPU9TMZaVeGVcCGTZSXuj/KP6RbtZRb/xxEYs7rwM2QEI
w20xGtpMxLH3nDFo+wxAPsdu5a2irSBr2ErW+ycGfxZeRAvWBQvxNOvnAreX19X9yRUhpIHVzVCn
wZsmaa4lz0kzfawskDNfiDfnxoTLp7DdiRFlE599Ds27oz1qTnZnFpUXaxq+MKbFneroPrt8lB8E
/t3d5227D43VnSimHJgRbYVKjzrlLt4sZ0vyKLoEaNaCBt50Yci6YIIdhMDOYp5JfrvMdcc3Lwkh
5W1YFqI4W1KTGsRTLwcdKoME7VICPiIwlWD7ZgK2xwwhy7tffNXsAYLLG/1o9xZSz3RvLn+IED9s
OjfF+ddZWXy66kETwXoUlHRSGHnz88BkvaHsvU5UnXQbGg78ORBJZ/Lhr4XVI150o7POBncUYM28
qMxG1AvCjvitPuSsLCYBRcFZrFxZaRetH3c2beHYCRDUQrxvT6HreUMZZMrVuE+6ed5YDCD0ZoeC
Bt663Wi4iS7eZnCaEd3/8z8x+w9UqooUJWoe/W51IE1PFwLduGPdPpRdEPAT/ZN1L5XeLJ3ALiLH
ujynNYj3w078BXmtTOv4K9rni/3xnW6u+FhUAeXeSQoz7ueOxj6ovJt8PiaNMqsiNXFYMxyWLaGH
w4HXmQ9KszRnk4G52CPGB5tDyZ5OKEhjBnBJAR65tcV2co0crHKUGc10v9MJpCrbbYlaKR8iYOjn
cjB9dBuNRKwWA5BxBb31hYAJEZBMpDIrC8Ekkur0+KEis8rGsLJhJo8LbzFyCjMakRNb517D2oyJ
krobG0VVGlEaun2FiJZLS8w/uqHwyQEoOczqjeLv752RH7QKprb4E/ReuxCH8/7lb2u1UiUK5HkB
bnLdqEg5o7ir8BLdT1I7gaouyM+33Or+3HXqtYIYlnh7k0TUr1DdvOTyMcq9+WdoR/SQHM+8jgD1
kcqQpHuvIvh+TfIZEwWGfo6MawghAQ2wELLrCLHrV+TMn8MageEB55NSK/FUxkuHnvHH4FTDq2Qy
aY88owLRvk/YmIn03NMDEZ5WfuI+tM3gKuUwiROzxvSXMWNhh11zOKEU4djRE5jU8B3MccUoZseF
ICdBn2aw2rLh7xLsVfHxd3F7SMsl3Jzfd19DG3jYw/r7fUDFUqJmaMXGtJJN1O26+iZb+a91cXE4
thFVd2wFn4l5S+8x54+7G4AHtcng1N0sHdd/zoMo62auu7Fr2Lu2p8NrjDXE8frlVwQiYQFMempH
+R4irnzTP49bSHikKx7VoTUFHCcaoprl8Cycgbv/tFfkOxMJ0HZ40XZfk/OhLfVA7vYvc57rRRd4
BcHDFpZs1c446x96HMYCnV1G7cnuHFgao0TVL2utA1WZVwteB9B6VXHSYmLnWH55uW82uv+6VjxO
G97k5ISly92Ft1NYcjWkIircSBTYIXNvoKM4B4eb8ykXRR+T96X06SzJCAOQc1xhqS/ZC0L4fMyB
I5pRa1E7UJg58e32Dr7YhKPem7Emeuayc3/PvISPEqpN2HRRxGx1vmpbJoKCvc/43IV/wXyVUII1
i9VFaJOWE4D1V3dovrTtOzNPjM3MZRCo/OG3161uWTuXmwa3GtIu7jLDd10kQXHn8H+UoLTcrO3Y
GTV8ogoD/p5hGUD1xaj2f3cETjKMcMCBOle6Ytxu8QdH9qqlDpLQl0gwNU/9LAEEm7yB4D/P/SrI
YIzglCtQkqTtsnr6s0IrhMh59EQRCFAxUQIoOKz3p21vBX34WNgwZlHVlWJpGvXdo2H9Ko26vxvV
46eYUetVDpM71hukNJtixu0eFfa9Vo+rjf5BzYNXWJYimG/V/2HNxwR6Bybb+iah4r9GGU+pKIR2
tWMkbE8LXwulKSR0wdXQzvudtGwt4EZmYn/91kc1Ngmi1XzplIJCQUHv7hkomnh8VnOkZSGd+l6j
GqV64Sgw19/IIl4RxTeIIh0n2busRtBT4g3yqjdmdW83TUR7INTlWgrdThYXQDc8VJlLSsktXoIu
AOxbvaRON7K98WbdBzR4EpwOtrci6LKSx1sJcq0NWGTtMlsK6ItuW5AkQAcymlYRZDVDvjRTOL95
A+xArgFPVwxO1Tnc+EiQVhq6aDw7YhvTkC7BSfzw90UBwFPg9uNxx9weLCBDAaTzzjG6+OzmDFc/
clZcj3Gy0UoDRI5EJobQh/q8V+81fI0Lr8k/SU6JeTlly+nHr1xpXAlm4SvKsrq13d755Lj6ZB4K
xsT1aTi1iWiGyJqs22lCnIoiQNcG3XXBtjRqmbAwddjTjN4qZpccZkDrzymGZb7ak08+hv2kthHi
SX7LMWp6pmLV5d/CZ+0kv3Xa7lbgMyaJdfAJ5wta0XQJEeJP8IGlIkNjwoFU4dEeYxUMkwKXA/Mo
/orJ9M+TzLZk+9/papyIVIsGJ/+4pPmtpzT3qjELSdI+K+G45LCg70JXm2hW1i2XiWWy4+NXvcf7
pMJIKEr2R54G4kjrr48gQqCHd9jbMH8ALLlbWn7xvEgxnG1/E/ASoloRWJMHw3HrAl5fH469PZNt
Mx1inxRBUAcraMu6cPvT4APfluAMuwWTve8B783XioWDqCKre/aTTonohbuRpWulRRi2biWC9qUP
YPPgv89+C2OmjikG1zDlk1gaMDFNcaj9UOmbFWs5UTqAT4l8iJnlb28P2kyu59lLi2U1LtO5L+OS
iFlf9TQXpqC/0mVmMcZGnthY/0Zl9t118RH5S4DVPuZUorIYDxU+b4bSiiHzEnFt71axVO29Yf6o
wxalXbXfsLhnH/XQgwQmAplpHGHErFUBe1hbXW43SxgHszKUndpIW52yEhorfDwrBYBfr36LiY2M
gir+9qQ6/egpsGWqd+6sXgjmrZRRCDT1fmQFlCdeJ1uVmrI8ja0ItcgLCS5rzU2/2w/FKSsl7T4o
NyEcRMTBSeH5GsjfpZQfkvx40jyKzg7QF2xdIN7/f4kuep9QI+rAhGbGzoe+gc/dxbKeJEoWx+Y/
3yt0G0VucsIXCnKcbx7a9rrnr1Jso30UfujLeEqL7yG3yWrNVgTuAZju/lep7fCjxsHENP5mEgjS
dUSr4/YWRK0Kb722UaZoZkxrLH6ovlm0ipOlHF314/Fdq7Cw8XDRnjrzfFvLoL49fE14pOfLnONK
5TIxD+yMQWQ8a/+BqsiBionNh/RAKzxnGQRHXiWhV/t/X8vJPwgY1PdEvwj22ZFoMUirRNkBBltc
Y6QNgcxQA0pYBfbEOYsn7ydeXYqnkrqeKFKgwjCKoUZmlCSz0AwkpacE7LkBG2xCfegQoLXUJ4ot
25JnFdxpGQ+moQ1b+kuDy+ZKw98HNGQuxI1TIAJskTr7FA7wO578V/sLrZSdKEGNr7fJub2cWJa0
9dbuno9Q0CtZs5R8d8yVQjLFJ05qND9015t4d3JyGLfPVC5FIEH45be4J8hov0xKLIfDNTOUuQMM
iBNIH/4Nt+FVwbgPRW3HhI85bPcawoJH5MyO8f9LEGCWlSeuVpjwRGev+8QZN4iqaETK4UIb/V4E
90HsE4BSBO644akN8ZBMymtKVjuF7lA2y0Ru7pvEndWqVRE3meddBEIhL3Z9fiUe/NXhRGc8FIUr
JtuIejtCEuPw/8nutRWLMvu4l22QH0qO8FCzjuArzj90J9SkHi9CwVg73WtLzbw7OCkjrpJEz1ZX
Hyw3EDKytpqUi4tqOTNpDOH+aLPxorijLpW89TC2ML+/TngfjTzEuWr1uvqFrLbjSiLFAJNbTitB
KHnGKDqQwqw2LLL9dpglPq5sX+MyVhXruhFSaMAQFjy7TCSe/0OAY3EVTms8BJ9Uknqbk+ySdPll
gyzAgRMN+c/MBFyskcfsWFgMyq9oY7boMgIRAzpKGIHapfoFCzMM3cBGGSYEYcT6FiNiowS91GQZ
fsyo/06ki1BSU69+2MuIRk2sdkJi7BepYp7X3tE7XSMND0h8i2gKJ2EM2ldMslwXDwKgC7xrErQT
dQ4fhaCNbH5USAHQCzVHi0z9yGBl6cxComn3aMlufqgZw3yUI4xLr+4a5JsehBt8nICNxPY2E3bB
EB5YLjih8K5iGV76RDomlDrKZWkOzxVTpOVOI6EZBeWfM8fDjuRUP0qm8XeaPDbc0Lp4owg8zOqo
VN7/uIAxOr9dXPF72lsuQqdEBiyGsMP+FpwJYUqcsT2l5O34YM+b7CW6tSyon5kHHc0PNocDjUXR
PPv33r17jOOSAO1zgFZPEaK5qjZrj3+bMTBDyUp9/QeWVQp2wJDRgn4S+RSudLjDvhTOWe5YihJ1
xHoEHeK5ulFDRezlFKIYf2rXEMz1+sSYA2F1ICqWYj61/lLCyFYBsODcdk5Dhe+5TTeufgobzGr+
K7wwrSf6mTLlbXVpTt9CHvY897VCtdhmRO/E1jAk5vy3mTmUuuyUEHBrlEMmpI8XsO7BEdDi2G9s
maoqtmP3W6NIKIHPHEBqARhOKjjKBXhleFINixhuL27mS2lQofQvmTtw0Oa/vLIjZ3hD+u4PL4xW
zQtHTgZ9M+0L7ynOYzFjIhT+3F8W525o3zdjWg7fZBor0e3rF5GLWtD4ZjwIckF7jl8GmxV31uhE
822eIVi7/IInAtILE7dZfpwRdVETDrxTvUNGmrzIrvXIlCX2cA2pJPMxYz1S1hyp3I1LO5thODg0
RiVTkMOLINu+ZOtIGSpkrEoJtgwLVclcCl2XX8bgzM1IdHjUyMTRa0BwUKP5Bq9v/qpYd11QDeTc
NeDPJAdc8h1R1CLNadojxjsuAUpVGlhRGNEibmq3837uUiqYYS6lFjM6iFnGtGEoDtZLu/+8TFMh
e+0+WRa2ylLoBrTlHgWlXcZb6aE9rfeX155eFiOHYJdzNJu6icfUPDIxAHGilnAFdOk/Bn/w7+3o
OsHflJhHgAxh+W9WAOrYvnP/5FqKmrLaiLXCnMgBd9Mad+0HHPk6qlCFJeADvmuXN9tqNx0+UaKQ
v9z0wlNZ4je9O/CM4ZNeORuEwM6wYvD2PCa5ksP7gkOQekEMOnVQiF4dTC33G+4gS8b7h/1S+LrT
lQr3eNGKlyth1ZA+a8fEMg3dthGdAk89/IeEznNaBTTwlsnseMZxTon7AwYzGrKH7MHHnjpUhW4E
fjffXBcvxKrcQ7AArQi9lroh2WRw4Gi4SLKrfwvl/rWWXRZrigzaxG3wT88+wHqYxxb2pG+kdjhQ
A1gvilVapXWavF9vHDv6iG1My01rKoajEKAeRD5rx+6vgw/vgKMQKICX5cXq6eWzfHJSkTSDf08K
CuFN9a3/YsqxIwk6Ji8hC+GbKl8OeDIbo7WB/tlSVKWgyIoINTEk5HCPfLnHkcGpFFqbbSfmhUpV
W1FXQHyi3/1MI5JNVr3pICUkvey48bnNLbiPQZ+kf5e0/FmORsGMjfctZnaRydjeYT5P+vPO+wf2
MGAQ/fLOdAlMiB0pzmvrQWk7z0seWZ2rNDzWbJKxbGtWpNShshW7225/6kUSlVxNu8XBo/OxOsFo
DHdY6R7pOXHSILAKte3X1dakRs4Q0cx3MIwEha9N3JhCOrPRtWAxu/+ux2pbmeLM5tNsVR5EQI0b
oFHgNSkt2UyQlJJokSrtqAFY1DNLgWNvetqCY+LrjQM42J0lD5vexvBvpTGTQe6JcjoJk8/sc6MJ
QWWhjgcFq7n5HIRjMRuMghEUNtcCcXheL5LSF4RTkEVHRPo04CGL/5BVPb1YFTxKVWpw5fC8lsjv
1fq59ShBODWRxhDhurIwPcDbXcRydb6Nw/qPLdK2T2X668zy933HIDQeir78YoeRhLPNDDuyzVIL
cAzms6DMSpk9ZQy8AkYUsGS4gHUyOD0XtvdT/6gQpgvH/rfnw7oZUY75KR0dB2ts8FtTyNGgFj4v
A3V39hDHFnULp9++2pYNbf2G1d9bBhGTVnU7y+5LHHoDXB24sMiYXS5gzQTcDl+THttXuOhHd6Mb
LxWubytsh00U5OuP7qGYTeACW4i/mB7/qCYvJo8vOnq/iuuZJfJTuY2skx8zq1/we25PzCQlRP24
W63xkYmIpu5cYV3Hp2lcjj4kEB14qaHhVQyb0+eMHDTpSzUl++oegni4/EmLO3dZuMKdn+a9GGzh
P2fT2bz6nbUL75/+HlKTioYANJ3hPZZcifXhR+LT6Qae7wgDpt+nv2UIcPCbe4WPTCJNKOzdZH9d
Sxsu0lbg5wYCMsXu5I5Wpv+C89tS2no9ER0a6fQJfplG7rcOzKZbDyOqPyTtwBOLAxEjIfPI8c0m
cModrMo9ZHkcYk1iutvtt+1ewlNy+5+HzTnynae+V4Fq589C9GJxu+i+wh936LcjVjf7YPOYz2YJ
p21YZNQfzssmkj9wcEkBfxDlI8IihWIQ02G7Ct2Boydsu4/9O/s9RXAdk3iQTgLB7kdNKLT7kHMu
NYfm8/xURvJPlKj/vmlqORTI11vwrmKY/tJxaiWCO13LhVhhwMbBSwOXxszop0k3nErCdQ90zOAG
OSQQawPJQg5jQfBx/Dgmbal95Nj/uu3JY6/HWZslM9nFnaAfxvSuVSXOoiFCQZGG1rkO2pJ+7Tl4
KDM+Df7u76XeNRwgapb7SOG8/BPOxHXkqV72qeTAj20qH1sSsAr6yU5SKtsH4d4Stu3TsSYOwp6J
IIiXT5YaJHwGPrTDsRQ5sqDMfsSx7uiREkDmLh3oJ6m2rPtQny+aHCG7K3oqj5w2rSCRehmCF4vg
rwzfsMiOxQG18tFM4uh2TogWyNDuCY6c0WcVtdAffSU+ElJRZsBvcZMXKfbnS6tT6wjT1VLesAGi
mBuGZtEoulLeb8LEHNnd3uEUWcKnk88j/9AKQOOBC63i7+vC8j5oH8g9qIVJWklAHIkFxz192w7J
eic5RuCoWf3RbYy/YVJ4gZbeLFsI36UNxn7LqFMP1I9pTuu2fmpEn8xtvuBmv2ykZIqNo9DIuofV
sUUSUahP4xLFhqbieWS8vP6c6dfNEw1zJJiDKYekWI/C5QHvfvTopZKRVwnMrcNm+clOlMQsFYGJ
g+TRW6H3wnQyHPCMcu7oDt/MB0U2kd2Veyf8+gKtkqQxXzajro0AkpsbTlOdBd2fpiJI17Ropskx
DUjtoFTFrSj1rPYnDB/drv9WL4bYpvCvbEpyUaKJTtclTvasSqM8CQ9IQ3UKXH5FPTLnjgPAE8Rh
/fYdRjOwu2/dwThS3SXyQVl2RTVREgtCGa8kwmFdK9HSH21adyZ74xyEWsBE6rNazSw2qtJMm4/c
KhQDOAUuVGlOKQs2WYcHkOQ+mF8NrXnexuXeHGfRSLYILJMZVK9avlJdeLPU1M3vmSZ1tO4VOOu/
dGIsQoFH3U4XnEY4C+yYJtfTSBjwUIPe6l2ell1lzdpQFn0e/H9oXxIE0MffOBtwQ+M4BU4OCtzI
ToQGU6cqLwrlkEK0BfY2SWKVcBLnGZjufWGphAlTr/sljaAEuDu7zC6XEkp0UC24dJWOlnAeG4y8
EN6NqiarvboT2fblkBWbfPK6YrIdfaCdVIvTtk+V9ZtGQUx4h4p+HJw2iEVufQWCa4th6xTA/cEF
uicGsTnyYFXKvbsl4OKY7EjYxIl7b6/85uObB7d00NTOZFubdUVKRxdPLRIYYvSVP1008Y3rTDCl
pFdvtokXo6NbfJxa+mR6p12nY0G507zdRSypm3glxR7ktAzZ07WU5JWQHtWBuusHfbqazxKBmd+Q
IjfcQLkQ7F+8w2U+tK2X8lAjI00EehEFwWq8kAymHqXzfGONUbISOGifmSw3yAXdeX85v0aD0E27
V9P/OJ952zEyiTMmS+5H0Cpexw4rHAX6G3iWpzTyjat5ccKOqd2eEtar/AuRt/K3sLTeWUtdvYaD
DYvi4Nw+/5eAy3vOZnJ1OtMFPAd3+R0XtOOkz8maj3xnq4UXCe1y5i3og18eoyoEnYFM/9FqDdFh
zvj8mWPMF9NEXcqGoAFOc7SFB+Aacske3vj76DxGqSBVIC4TA+NQia7iCF0Mq1KH85kywV+cbb2i
zF27Kymuw08f0ZHv8vzd8H0mLuufZng8k17z2UA3aRhv5f2iiYwdbjWWKVka2wX64/dHKxdzpH3u
LWhVv57mGL12P8JO1/AJfYQgEWC5OPmfvGGYbRCp2dPnSdM5QMVQ4mhbmYPvB8x4YiL3fdMl0CZq
X5wTqyZS1Ol0cP1OlbOZjmN0v7NB9zIJ3q7xAwsNivJNBFC3lC8sbXpb87S3eluLwLy2pO7Toy3a
L26dFuxNdnZhYjHI2vqiu73Z7fjpqOXTNZq9ZO+tNe/zUz87MyynnyVANdkB8WCa3WePrXMzPZKC
CgjJmzaVg0RehvIftGkC8JTugPwibnKrRUsfddQxDk09iEWx3x+IKnCn63Yj1phe5EwSmkoUNpYl
QuENft7RyRGbDydwVF/KZvHE9DaglQHM2vPgK1ZnMH5XSGBTueuPYIMiIt5yB1kT9X3wu11CV5LX
dwocT5ThWtfVNadylusYGtsmgKkREFxz1AmGk3oCvlOU8PhMvIzsK/AkjlGBDVGcbBIamUcN6zs5
sSpe01drXJZVSBlcei0qCn43XjbeEVRp9D/ZQGug0w06LHRI479ez7Liqd2UFi/SDXNV/HnKh766
0LNYpXC5weUxb7ZTYa9NseprkLNOFdSraR1RLaeSg2uwSg3zqliABd5EUZRzNiITVL96N3zRr5Cd
m6L6QYqXLVZJyI3glmqWRTP4Pjr+lqt9rBMrH7PazgTIVPIL5kdETJvaZQcldNinbf6a3ZEh4H1K
N7yye8xHNTXdTrLi0iIaApaV0zd2z39wyjV6oivaXVT2suaRh0z6WZpgD7z+mn8NJY41DcrIoJ51
5MPA6lqFMXW0Uw17qx6yDVsn/jxfJ5XyaM4MH1E08+goeNgZInsUb94AxRQjBjdDhf5IHQYs8Y1+
pGPiyuX9l4N5R/mxWkC4+NvohPN3cZVeO5ZZyRK+en6RP24GhWZOrFD9GeY5z610/QHe9o6zzf4E
b8tdidp2sLB8Uoan+gdQe8yFER/VcVQhywTnmDvS5TmziK414kVxra7Ukvp9vmqnXIbk5r4eJcS2
raGB5vudY6aoJ8W+ouxkwnqYUPhkd0u7YuzAbwdIwKV9YHHC/AmS3o8W8AfHhKMgHsRxXnJs/n3C
wfuFmn2fs6EOlRUCi1RY+/CB/92sCuFu9P0BPqsUfO7EtI4e1YuGWoO8VCL1zfWOb3hSck7JNDEp
fXdjUmjjJaNo7qh9kM/DLOP4rOMVxa+2nW2UuZs7/XOWktwU+sbMupawyCCSKnVPINzcth30MSKZ
EIsF2SpqoPFDBnhLAF/bRxA2lS7tfcn4JB3VL3FlkXl61Zba1IkG6w6VmLAWrxbUllicjFWnmhtl
uSTETGCMtJiU7HpzgHB8hEXTi8vi5uXdZ2QaUFcQdGIsN6f++BU0kSdgbZCzNULFSc6Z3GPq4hAg
WD+EAc0liCoEnnb2WNmWGFmIUj5+PqKqYTr7kgglTq9kSQxwVhynAYIpdjPtfB4noLoPnA0F11Sv
WA3G0SMTlKkwZM329rNTVDAusZ/B/ufwAFElYpNJ2j6DR+sUgI4mXou/ENZ7CMTypw/NwvG2yFHT
9DOP4UnsXpQGwqCAo2CWMfi72aWhyFajLTRwZNAmrbyhFS5Ns3LXX2LLrkTbX859wsz/kg9ERBVC
bInXLK6j+MHqHJQ6ioR22wT7eV+ao14V9HWkianeeSnmdZsVpQZ36Snm31L4RBxC2PgXXftvg+u/
OjIY0HlNp2aTFgPDklI19eptCMTar4FDgoSUWeBTchGI7kHcp/X2RaEsaOFJPB20R1hrrCtrBvB1
S8WD7yR4kfO/ZjB4mJZni4qtBrdR0jDCU6sCzQfgak/NjVf+Cyb0Cc33quXFFzc2u+iA9AMdZSf4
mje3CwOzlqrm3AtkzPsjNJbsDGsHDWp6mFPdDDR8vX3YrtAAuviiYrKrsA7M9gQWWrnt9jR1hgA5
MkNd3r/FhRg5QviKxaBNvcS4gbboPHiNgc3u4u087TAHEgT5aL3EMHy0f20bZON/9SN7pMWBQ9Yf
oh9yzy2w8J8iTf57b2B9Gjz7O86I4VLAO/UQT192kxN6c2YjZMWEdj6feUMeX7ejLbZw5CWwY6CD
UhNuQHjLbsdeMjEX6K2+qH3hO/iNbN2/JPf+RGiv/ti8Fzwf+aS75RgiMDry3VYdYJHzps9lMc4x
JDnLpgAWh1vb7uFPnOP8+z7HKbuC6XHUiM2zcsITb/pdeG2bT1nbqJnDuX/fJbH/Azih7IhjODqg
XjgGrSFWGIAJNSMR3s+V0pJ5wcCWtvGSC0s8KbIKyRBkxdSj2/QI5eoz0JsZgfCqh/2QZ4o6ZWJ3
Jp5ubHhEvXB5fhpl8t8VemxJYRUqPoPeKfrXi8IrIQjZ9+Ltf/W5JJmIOn9VFedmDb6Ii4AVVPiz
uAbZO3ofv5d8Oy6yR6gY6SJc+njcIImXAtTOg+kTwOZR6MvHaAy477VTMBEW8NO81rvDLsPH/0ns
s3EoIkb+3H89QdWmzWFR/fl8kndmz8MkeSGJXMZrQ6gsIi0VSqNOH7udxXpUXLfAUwp7pWYoMzXJ
wFiuZ4zovMUY4YmCr32YQi6pGTA0852n1EZpvlmYcto1BihEV7fui1gaj1Z3hg4n0/jOuSnPwP5g
kOCwhpA1kkjWDznu4VSJ+rfpnwP6nMswbCavcngtWyxw1MHF6adte8GFqYTPIVirgOD9l3Yv6gY3
wjFSPvTxTxmZ8sgfb+5qaN1yD7Es0XUyJs2/nLVEk2WaymuXrplFkMx+cuPJrh35R0j6tnl/Je02
LxEcvEi4Om/PcVUu2/UuUIPJQytYtOWz9pduUtHNKAQ+fKa/SEl6eRUhlrgSab3DVXyiFUt5VpAs
+4tt5AxRZBChbbyKyDDtBzCRb0EdU+x97LuPDg0ZQ6eoIb5H+wfLek4MsVn4q1dDVDDucRnVw/z2
yu5RiWOyyuG8Rx9tzGEamVp3rbwpxlZQ21S+fk5Ycxf3J/EDTqTJGkpBt67yJb63XRPD5LoXvD66
AkO7PCVAbgAvtAsgItIgtoo2z7NVkygGZN3LDf7kTQ633UUH2MQbDFgOYCtxm5DbalcetOYqurAh
GbkfzQz+fb76d1drw6LCBFNQS12+mw+DBKGe6jF5DJFN+BS1FxnyQ8sP7NbV+Yi9nP8Je46lcxCl
ydBq9F+zZsMs4f+B1d/3aUXJmIQ1Agl42svMH/5hnQe5ylT0p+xqVpuI+Tfj5d4HvgtZP5mp2AYO
K9l2hdw+5JmXHGCoCfo9uLHXPY5EB2yJ9RNvDwn8aF2ZjUWKPo6pR9WvuZvCMAiRYDQwAAxt2Crh
k+9saFFVSrDmwwQC5B279nd/qeIs3KNHxtvg6Zm4cGNovntWHrzDiNd54Lez01xD0BtC/8Snpc+e
KHGBH83j0EEXsmwSRpvaxBPMrtrd0zybSgksWJc5YTsHCgMjuefDJdZevxY9eQIqYSN+pgEZJTPO
qxElIeQH1V//Msy16ASb8UYeQWrC8SDeozyAHx9Ly5Po3yUT2es8GfWrXOZLJhO4Lb52BGkx790i
QP8m0vEmriAF80masI8m/OoSTX/KLkLNC/hAF3sKKg//4hdPhUxS3FptJVz3Vn0KUVHVtWey5J2d
jVXhTZ1ggPSP8V+cWN/j0R14K1sUVURr+6WpNfgw2gv7CWxthm5+j4mNR4ZGvldjVYEFDGIZF8HK
AoUNsRdgzbkwfwUZRIWEiAr2rzehCqVgKtyobWXC5jn0k3IX+8yqoEFYrSPltZHJfGAQBKJosjUb
TXad5E9p9McE77Y///oq/j2SZ01YqapY5Pu3/J0GW61ZyEKLrAWtfNp4sSLuk7TCwvgdHRRPJM4p
zx+an/0Z6yolv5rY4/H/zWvpWEeRoo+f+q8dTNvZ9mSHpdbUJDylkaQV06qMFjBwcNECrNhtfwCp
u+XAChZuTDhZL1C4BeUmZV6UCN3J6V3dceS+MDuKuhG6mBZgunlgJPxRevo62HL9oYdBC2PN5Nol
tTQXEVCpPBo892Nv+2gDVb+qrJoL/Jzl58wd8ibqSw22LjRSyFynjRbmdsIJx6lZYTI03UbTzmPw
3Q/gRyu+PXUPUcyJRlU2sivK/dOEONUJrJBX7gBb7iw9+N8PS4VJ7RyoHh4o+C8deReaEx98YUto
6S+PHfAY3UtxsSXPeluckgmO/yp3uoQuBC38woLbY1fs3Zx0Tbhus1dshznrdV0U21x1Zv+CdVVz
l6SSDtcHePeO+SAC6lKp7YYyvqboGRih592zUqB0BJwvLeyTi1dfRXat4nui9n+ZaXeW2+5hAmNW
bANISemWBkc4YiQatS7qfd1Vy6Q6IdEaX5xPKLuFGV+r5ahtt1QUsW3/JNkuE3FDtaWlRZE/bF09
ihjLEqSO21wrgCI3q4x1jxaxtfZSnLx2qbZ5WyBdbrQ5UH7J0K6neb6AMbzHBn9bW0ZiKEbkTp/2
BhBVL2waD9CJLJ0obEu1dhvqyWvd+z+6HA6NnribOPab8ZlO7tRGrf6LwPtk8OS6X+j1PzjjV5RB
cMUAPbWCIILD3e6e1gx/N7cERIkMRaE7556DxjfVFisye+U1lNi8M71ZKwcJpSxVNlDsnp5TKlnR
TRJvYHyLE6LxLe3ftCXv334STzvtSAljxXniXntEj/j40EBVAoW0UHG9MTlaS9ZAOt/05Styj1Mx
kr+JWNFe8MWLKtuh+pk09dUF+IjrhtsZsAGHlS55pCLHVO5kktxrGswDiWhghRtm7B/RM2ay3Ves
MdGVZhxB8y4GvSC4EC1nQUIoXJVxjLv1+tg24anVgYTEgcx5swdU94eN6W41fO+i0q3nc/VRkhIy
WY/swMUbYNnAHBhrAbeLofc0peqxX/Kh+I/zVqRicIRLa/WQtUaNlgv2TMCpd/E7S8VdNRoW9SCi
+bpMgjbmMBCG5iJAON+SACwxNIPHZUA1m4mfUPHNZ9E9W3ALwAmfxZcymNdNxs/jgcTcUz1RRIfj
0n0uK+ledWzqGlaoXnTwxXHSBBqBmAJ6V9x2T4npqqDOm2T9vKpmq5ZAZm9n+MxchiIj24Be28Xh
bs3kKMF5l1R6uL6bpyJYVKf9BTFYi4MKtjWeudFo232+MSsSjG/Ah+kHf+N4MxHCdFDp92SCb4e2
GbhkETsXhuHzxWH4+mbjihH9KksJdFeoWW+IM6PVaHqHOiZkSPNpnhXShl202uAgk/RG1v8BKLr5
wCWsDSZrqbU3I/7zcsUxT71FX5CrntmnXkNCTPoqYwdHqBx3Luir+AsJus14EnBeqTKPLGVFjPez
7ZEKwgyLmWKs71kn4GE55To2mHsZQO5GVs7u6bKtFBzl/Gu3B4iWMoMxybwdmOZLLKmj+Ay/cWA6
/IuMs36rzY0Q8jv6bSog1oRdbJG9PyEmtT1Eny4/Z4G/yDu/roNDwlSn5Sd8Xrjz9k9+bQ0Tmch1
yzjxvc7ak78EulfAMEdSuQFtHaSzRh/V+iuHvWLqvFs53jhv4xrkV6i05+nhnxef2riHbHQf1WhB
+pEnYGFltDm9xA5QomRbf6sFSRb8LMnMhTMdB7B6GFrmtJn2CZepEZlQ5Fz+x2Crt7qA9xFMis6V
WU1AJmhr1hV5oUxcwiJt+9xuSVViUcfyGHw5gTuNB5Nm29K0M2+l8PhGC9FrkHiSi+p26BqvN2zL
yth5rhkNAe/ju98UNigatqkOYVkxNlNFWNuN+/FgkRscOA9IFtH7l0MwAxYdjcI1BJWUOOdIWzf5
jph8uuY24KeQmbLp1yJXONNbWIN+brY6/MbnoQ16E2sdb82oZ/h8JUJDoqAMQrd5uDcoAFUiXHjU
gvFsyUEqZMo2NnmRCbOkfkqhQVTDyc+ODaM1pHkm0met/GF3Cs8bVZ7a1piAoqEwXnFi8lEQGj8k
Mp/KqiepokyedBhIjbirmMDp3vQoSr4f6gBs8HqAPb1VCG5SDKmATM+Ej5psjSNMnWCjQ7PnTFCZ
kH1gN5HurqKAVffExZ+8F6zuGFX8FXsdsAStBaO3kSwyRFX1BoIsK+WgqolCbW2CFqtbVutn0gz5
xPQcZ3JBPqJJCc0+iQgvzBbTrt95jRU=
`protect end_protected
