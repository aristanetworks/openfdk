--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
gquRCGTHrvPON47E6kBP6O41DCX7aKj9PnkqlGTxBr0UBamUXY7S0xTpKpIQGmiaOKWHx7GZeC4K
nIa/xcIJdJPj/Jb6dV7NOFQtkXVf1/x/WIqPKa+qMJgN0aFFREC7ezBgASey/Y4E3NdLaev/vQSo
386A2IF6o0gXESThONfaktVpRiC8n4oJ3K4RTV1YIGHL54FLk/U7lz6oMo7ugCBY6N2mOmYzJ7GE
XRmqG45H89IqxgFyXKnlWXg2p/u9v+vrY/FHcZEcOsD4yfF01L41oxlyE+bwktw7aJdaGgMufk0B
mVjAmRcianebfv9lVpt8I7SxCqfFLS5vW27gLw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="AQuV4asYM2+KFugLdrFSZ4tb8r/n/qhGsSKnTgbAKc4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
qY4jflry0886jBvkf7rZFpTLHPVec3s1A3ymq8xEHGbkFytw0+HKz97XMe9bPHD8TKeGoGUdquMB
zJJYEN7QU7QNY5ua64/6egHvvO5UI/HO/7bH8qdBTMMcRW4b4pQP/Sk9J0YLB/miD19CSveuIMnY
Dh6WZD5LL4h6qbkhjL8pQHZ1hMAKsMzykP4J8cMSeWeevBBaY87gzq66jsHpXkjhtq9M5LdyV2GD
JPecvGYDkpJQbdW2eWu2TJ1/VlmVHK5Rt/qAiL0ETolh0RMUMuISGoAPX+tq1l08R4alaNGT4uYg
Lk8oxJFcBsO3mw6IjmFEFKvL7D/DaJKxnQkbkw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="puyg4MBGdaFiENpEMQg2IleljpoeWjhpMct6Rrm8I4g="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13888)
`protect data_block
lsPki/my474JFZr4P5xvcJwX+GsQzHSbiPDAXENCKbYdtKA+Zp6PL3J0NWXHx688gsqrzfRkT20P
0ZV//+H0j1miQvzJ6RE0nIRyyyWBbdQKghFSneiShw3r5EdYMnYZ79CDR7QIADLAVxSQRzbFHCY4
wkgNVAFBSWv4GN+PBDYtICPfWBTc/CSUqtDrE805aTohjeU9k66lYFOPwRSJnmziD8q1E794AHAB
rKCtY/pVLUcX3DQk3Jkc31CIDz8ESu2Vc1WTEKUzvRtWV9IaMW7fHuiSfFbR1bTqmL2m3vAOVn9r
R+Vn1KfZgs0t54+kyq3Q71+N/eQFB7DKQGFbaek+E9hFPUlkrJGUvGOkCRGeD9yLw35iCOnOdcpv
KC34lHENkZgmogQphb8ckKmpiIRoFVEqYbRtOJHEL6JWys18zUj9xoXDDjvvNcYMFuyDsSQapegd
Xs+rRFEfD7HwEuEez+ERi8XbQrZNdSPCw7pqF917wy5bvMs/hEOv7lRTJraBg6U0XhzP+NyWwFYM
WpGkEd+Wxr66zaHOJZt3s3UWH7t6oni9uuUjUzgrOXcfvvjfqa+ssHD95llGUr3dzmY9fQuJCk1i
Jq7bA0nNMLu9q5yzDyanqdjMnEJx5aaigYZKs5ztmE9t411ULnSXqcdIAQEKfKA8Fb0yEuwYu+EP
U8aw+luw1Gaaf7hrDH2iWzIuj1e1bYSD0LSkZ2DsuxnrrWKPYzbnPlPzc0VOXPWFQKFzDKY9rJmk
uOTzpsytNvJnXxLDdVpVMqtojc1Lv/IzPNzaxQUa8gsNMa9d67gmYHmA0awz5HRCNF1AR9xs7DRb
gr9lRhifWHS7X07//08SWt/gQnEaU2Uwp9rVvjdcALQQELRvflOnsgX2ygohRO/sEBd/Du8ev/dc
einIiOefCw4oodJ8VrFXI1ir7TqKWewUNMgzHvF2jPbY2y9J2d9FbULIjpmHok1B9zBCKzjhj/jP
SwJxHye0VjmkdlZQ4Gvlqtk2IhNEmxe12y1Q2D13sLq12lHvuk7Y90L9J9KTSlNj2Yh2iwWeoARC
ekpEg01VNvCT5reLZj7dWXxjVNZOujnmfbUICdoDI3JSJKVy93cHsY0bU03TdmJTRmPJBL9AwLrs
Ucfpmo+nseQGN5veEEkt2GU9ElsUOkVP+l1ZQ6ogSNYsqlc2HElg+AskNXZjf2xBsdP2eA7zR0+k
QqmLFAI4zC7khQ9rgRefdQvWl+wpSLMD7pywMW8bu8rOxVIxu88BOcxfHLQwPsJIyRpW3qH/lb8a
4DwqJQ3OeKw8pcAdhMScMC0+Mui5UQXbs5z2SyWU4WocyaqKpqTATHiZ6V5PavZ2YnxV7A/zGO2N
F3BEKeP3Ey1cdK0ZfPYpTS8AwEgx0H+vAPMukIgmIIeVxagt/4f6/cN8+Wq4peg898rUxUPVzPNQ
y2FBPHSRicF4DgC4xfsFFkWSAcGGr0dDDRcZ1hKRtHfaJ97Khdju8EvvrRu5XRrZ8vqNtFJ35tV/
mOEgjbvbYNgA7oiObB7r/ta12U1FTAF1QUjmZM9BoHgl0vPSvucCUl634EOMiquUsNFjoCWLnc1c
FQm6gbGBSG0fR0gM9u+xRmGKkh9At+2L2b2+8etUP3n79+jXHaZa4KRFUhSJhChFXRuPe5++tEum
Z2Qk9DlZPdlxfKqGZ/tfYGGYfpWeaBvXeMzwHHFtAlD8QQAMQNzxXXxI5v0KuDTCr7fCjNcGn3Op
GswCZb+ajPSv/cVIL38xjXlctijlKrpoNL3VCIEC8tQHW/dPhYXivirlUOnjq8ivsFGU/Qke3cKS
TqKFtVYHS7QpvqD5v/TlZ85IiOWa3hEimw5AF4Mz2839oCoTx9oPfEkrj7DneRp7EGCZsYvMkyZV
WWVnysy+KWlh30Lx13zg2T2A00ABpTqBPnzomwpuJLeSlwSlZ7mLoWclWXahZJFfrEUogtgP1k12
VS02hfiqyNh8DqqnVX/6E5/OEOiZNbtj5aFe+8zZo5FEgDdDKsgoMwtCEGN1idrLW913E9Xwi4Sy
gJlX9u3V5l0rC9u7FPTwKWY/0Hp8HD4s1kKAOWeGHgQSf3HiZ3Max0EjEYXpZMKmzAKtZwjvmsyz
1CWxP40wAkiDwdhZy6E/LfECNB4LLWaqYQRHHSpKWKyUx4O7HO1PQVAb4n7mnmpjoz9J1c+wnmAN
DicqyUE0R28CjCBxKvmTcHNGSap2i9/Hrk8muyHOetXznScDVyvbgabwU3OMAeCbLvMt/yELUeuI
pHG4C6o9ZOjlJ8m9pgrR1L4gwKnCT29iqFnxcwdLKmvELI9QMNJlsOkDcvg6IJusClGJum1claZm
ttCZc/EvQTo9J1zmBxw6nShQlrEMMqMQSNAgns+SPrdDDucfJBsBRkWE2kF3Z26nUb7uj2/m++Hx
NFou7zgluZQ60jKeX6hk6Ia4Avy5RPM/ZG6QbVyyzGChvVWPB/zyRvbyKNPPF6MrBKqT7hTZP5n/
DEQeM5AGjGux6NXU4Nh4NcDfgGBseU2rZFcq1f3GIfkidfJyhI9wptOygaVlJTBelKYFmBJBfuei
WppCMbXqp/iOdp/zXIIRSvNPdBAHiWmGbe0WqW7EXB14/jhTgbM7n29c4ldiufnCZGYXAWMpGJqN
c+n6eyzN+fEpijSAxZooru/7Fd9Xh2HlQgL4hSysYrzY2jUzpMq94ApEo/BYKUrEoU0e7csCrtS4
qxwTo9b9ESSnS4Cy0+cnFZuXAjnnY28jybzSn+wNbK6wZIcZS/D6bC0wnkapG4EZ7U5TVMETdf6D
tPdkarPEeozYERuF+lhUypG/AwIgIyQFOnKqMd+B9IG6R0hxuAZMzJ7mkRPI07ltDaN5jHRwsMCx
TSzLn4X5g4W4FAAEvj19RrXZFpKaAw2nI+iaWtODXfo7zQAGayGy+WbK+/j5YgWaD5s0nxqEo9yb
TF2KcvYgK2etU/dnh+JI8+kkDsX6a6YomNph9t1moqcUvYorb4FKGP5oWQIB53mygMYjDHgBFQKN
nKTCuB841WoxbgyuaigpNBtipB6xRGz9Q77RzUHeSgLg68hXuHR8pNH7NPUXCvFCfYBjqjyu+EcZ
D23RbWW00iu6hnB9dwQhXk/hBYRaIS4yJyKTt5OtzGoZZHS/QB9nLEGlY5P5CE95UcZ39SP6jm5i
xBgfz04+4b1caYQluloIg4UXV0Sn8KrdnkYAFYSYBccWW0w7KLj7QBo9kpd09/qRI126muAWBvLd
gQglSGm65wT+8BxzxqRfjEdc1gI9amF43rQ68uele2OHHfH6oWzfVpcNnlPlyjim5yWj7WIohB1L
tpEbpzm1Lfi3U913dKJZj9BxQn51pnMiCg2JHVMA2MFXszgaiBk1GzxUXJCKEmuT5OHiV16d++9A
jJ+qyf7AaVZtvgMCEK0PDnOwHzGsVPq7j5yRKYJI1QAPL4QeT+c2T2uTlQ/npf++m5qTy9KKP5f4
sVqpKl1MGRSXTc3vyGsaSItxy5PiMmQ6jlgd0QW8Rczbxsxq/In1ShqPD6jF2txhQMmR6YPnlg6l
i+Rr5RLWW00l41jF4jf4W9Ja/TPfjRxL3MS593X/EnNiVqIkOmwBRtNMTR9ZjSpaCCRPFdc0LcaL
2GpZ5MHlwvsk7GYDxfWrkdqGmnMZxg7qC46plRc323SfH9GwfIvfEDQsyO+iWvXbvgYxGMnkHAuL
sWn+Um8RZ4bfySpnqqJLc4O0nQ3TUgqjDaXcu1KfedbhzV5dbDNmS6ia390WLfqLKRL5bcZVflJb
Wfoe5yxfvIcKcpcseyeoybE0faAak0r74tJVuzmXeFDDE6DrrnNUCvnqmf4M/QAzXNUHrKYe3CHP
BGila8oJJHBtFE50smmlJTZWJcFinIptL/u58os0d4ilLFOKDjrnsI9Je3DLHdabR/mLhftt9iWg
CnaJyiwo5sk1dBnRUB3P0xH834n//+Yb470B1y68XqRQ+d+uUo0k2xy6DIBew9tYTudtKr5RY2Xh
3EUZmdNHWQb2iCiIGFZQ4ar4XPlm/AAcNjkDR8Sc7yQ6I7RcgLlsgIPmj4k5dfzPVcMYstjPhY+M
tTDxGmzUOSfkRvJ3WduRkQACnFvrLJyvoTcLCaT6/Qex6ChC4s8N70DugOTW01EiTaDdDH7Jcplc
Xq3NStINDFaDvlb1qolHZq6mijnZN0G7piLZM60uJpz1x5GUCBD+Ews9w0Pkj1WNv7U68nW/hTF1
DirHhbHMuYEVLSjjddk4BZm2F4Xg3Kea1WrjTX6UjZQ8N5m4NNoMXwwEc2NEZd3QZtau8YhRzQ9+
CyxAgApwrYU8UnuaE14CcBaWTT5MyvYMj1fuHYWWSAIXJsCwJJF1ghyiVgAZpK0iOLjOzYNC4Njt
YS/sZf9Bsh5Iq2c3BTTi0HNihTNWt406vr8TIwqKKVAdkY+4loAqKoNKGKDVxG4PlEbILVcLbFV6
jrvJN73/33AqtRqo7uhPVSGAz2fY18bCxsNpAuEksQFUJWPcAz8veZCBft15FpdpCF28qa3uGffD
M30Ot4s66gw7PK+/0G6PYHdwyX1yF/8LmwSwy9OYOLJZyGph6oErR8nWqZZqbgAlMN5bYvGB5zBW
dbLCOw+eMt0iUNEYrfSoIupUrx77xwElnokLsib9mJnVhm7+HWcTzj8cFgF+ydrMkoJAaVGcQlPj
rsFPvxmmYI8RUHyGLL/o7DPa2QrOJcKo3DwmVzMqWmPOYpbK4jV0sES1vQHQYfuikJ9u8dNBAc5Y
Rp2a12oPk5PhCDeL++EzWWoG5/Msoh+shEN2zCRFfh/z/aQ7+uK/KXN3D1o3byDirPWK0mNtURyj
NW0lYklz69TT960srRBHHx1C4Yhm8ct4ojuqyDuD8yN7vez6jtsiF3Of7gbfUMpL/LxCi3p7RAif
8/4kShwDzw1Pid7hgrpxpm1FnK1aZ3WUnXxqO4Y4R+oC09VcWsL1A4DDfnWOAcp4JAk6hMM41Zss
Z0Jrw0ouz00VXmW/8o1I7udahOStUO2X8SLPfe/PMFig5koxW6+yHslcNXCFS3qaJIaW1KKRAMS4
Vh0HZoVJDRlLpWTLgGFKk7JM8D1HYLu/0UA0Y2Me2fqpDpVPchUFNN85ywEvFhVREdJI78jPI3IP
BVxLjf7CVS/+kwdeAm1s/bqyImv7Z+BuFCMcd63wMk6vo6+i3L0zlmQVTQuVdiCtbkO+XfTlTk2+
r868dcEi1v23t9aKoP2/ueOv5bwrNNoSsIzlShqF+bVQpTTaDU3Vxx47Bis8yCCEW/G4nFzxi7Zu
jPO+iPsNSw7cFnsCu5owHpj+WpUDnfX77hqBsyPXfSEmtE98e8Fekmj6a7knfBdtHc4Gb3ekk53K
+veQehJEiPRWaZWI4eL09wmFZ+vuZ6w/CWiztpkus2nPj3TVbBorXx/NMi78cl8/gUXa/Qiv8aEo
6IxgZSgRbFuk0CiKW+RECqMABY+SPXAGU6U2/1IuNGZs3XpA4QiPqjgS53Fc+UYRt9FG/lbu9C8I
yzh9bCeUoUvntlSYG2L/pc249DnMwHZZp1t8wxZkXW9nZxQJpQhP3uBoG966P1SvtgpvImn2NlNQ
VC9iF/FafDEmKkGnsGSe2Mkd6bY6tyAhHJSE7868KLnaiUwNuvyKwAiHOpkmAz58qvs9uDkJ+0xe
YH1saUOGO5u4Cg9QK38CRLEPxiBDtZ/X36Cdg8dz+bBvM6e6ShgfQYv9ums5qGPjs0aCMxcUEZwm
Iol3jnvEsuF4uFJeJrxm/PXpwaFZ2Wxl6SpDezuhM6Qa9RZbgwBvHf9zf7ZU5icrfT0z4kpBfkVg
dUZinEPQ/pxS+HjU2mMM1z/xKPkdMhoYueVoC2LVecr9Ht4bnq0X1tFe7mAmVUUPjivynOsnMwng
jmB6CiZMB7bDcKxvh4sNW4VPtwr/A5sgogdRZwcEdlyXV8Pxxq0uq7Ex8AjQHOx68uj3CFrHKoKk
Bb1RWX4yZbGGZJg3/rLQA7u3OL738a6cbeIBw0/3SVwVz0ICK7ySh8pQ2RXlfhEauL4CJb4aMN7q
zC2j1v0NwL7K+s54uaaikecf4X8IWihSVvTpfVJND6F+tJZ79jBm/eSdd2uUC3Kzyi0580SOXUvM
r9TdRjSX672PJNgFt00FdjwcIFOCO2l1Xf96k6PCAXIXVjhHqX6EXRzz1QrW1FUIz3OsDySOHJCC
KhAM7MRF5Gww4sctUyKTTf0IhDODVcuXTaRnVI4d4ntsb6uB2YDQYu9yAMZPI71vJgtLeoP1VuXy
nYe9O48vGCDLmv8h4irF2RATuPmGRWRbObOrcjje8UwnIQiT2AzF4b8B8IFw9WGJVxVnjm9RKBvL
uuNZj611qNALGTR1dGAlysT1KHlrXxqtD+5FrTBa1CLbChVh1X9viN347YNo3jdUYkBqcHTq1oj9
dIl7rVj4cSL0MZpAhAtG85z05TPXqB2RrZLu+FgmUz6cImJbyHaNIQVQcF5xDsbpTW4/XOJYLtHU
SKBB/MyHv8vNTK5j1AGwzkgpqF4J5TfEsM7jhVc0aMNjwmEmFXfQ1HqDgvQ/cG3fDDxep7UsiZn/
T6ecVUHGMq0KPBIBmc+Dz4zxD/bp1akyBdGi912wfCLCXiMqZTIke/GcZA4g7EDlLI0xYkX3oS8i
c2atCCQyd8FJ1lmFHGJ+Arfg34JpLQwji2u1JcpukSvh2lQJdAR5ISIM+1FXfX0/0RYCEmoaKnYs
PMUPPlfjrLCY/dCsDuOnkvXJF7zbTOdz4bqaetA/nqpLGGYpP84eFgrqZX5wQI82JdPup2c8oaZA
/G6h6O315btG94LhatZe7rtfLWvdGDrKedJOL7BU1bTxJV5pIWSmEcV69H4nvd1XhW3yfRkqNR92
sKKPN5GEc9iITtMnXmT7j49Vexi6LqL0VJEngsksoCiD1z2niHwExJKUeIm/H9TANaSq7/veVKTg
m8GtPo7J9W9flryJKzg3KOtYFOTiG3QhK4lzuESovf4DLSC//UEpW6fXicZujh2pA11q8dpEHuXa
Xm1SvkclBlyvHR83n6BelwAhRD5AceQb9OZR+7gj0DmvonpZ8dDgRGap7fJR48XLi9zju+8Ax/Nj
i4IGJwKBUhFxGTV83LYWq+yUdYL3pzcGwuxH1TkZ1nHWk/IoqFxNZYKIxEWPLvGAP27SM8nAVCwF
8vSRJcIJBwpk6ODIHFoyqkBbhw9RzlaCF2OD2r7Ps2doApW4QliI+IGhYosmOqSlJ5QNISn5GGWL
hOqi1aXkNobE4a5DxdmAmx2+o9Sx4MkmsGIV8MKCm509r4PpG4RQ0WFlT+FEkyZIcboGbxgMaJ9i
mzHvpE/h8LUNagLVrFinP5c8l4qeToaZuBzZJKvPLkSh1tCsYh9vFVvOPt7aSmzOW+Ce1tnqzlLt
QDOtJ8uhPD7aPLs0CSc97rtHfve4rGGiispNHt0h3zrnarekVympWSARLQNSHoBqHZTn9tNwCMmB
EJri+xlgh5CKqZlSHbEsVAkA/jXyzyH9hS4ItrcK4Gsk/RN3kR+U2UUiV/mlZN4A7A9unZruubdw
GCDu26BzBOx9US4egx7cHRDxxGYiafRZ0EVtpXfh23qJZzZg90LfK1Mrs6Nj8RrrLOjKE2eBW1SA
OTx97T9Fc3crID/0+VcqjUVmKdjdth9L3BlXZVAl0a0rn+4ZZPCC+H/yVaCvHP+PZZk75BgPHHX6
yhxlOQ9D1VQ5i2XSEMSgnpA3eS2vUdrekVLL/agepKTXPwGie4pdCqEXpu9SFsCoD3advxLSejFt
NxidCUPXbrPnsvow+EZEBW3/JYvqfkekKVFRuoEAlvhB+0GIk9BpykeWxlW1xazPuSroBY7uIzWy
NoWNgFnXtFCNoYoFm/JbjDkoOXAAfGssNs6hX7MybkelqUFZIAxlJHpqHCclE8MQVPpwLPUuRP2K
J3bif5rWDwmYjxTboS4nj5VNSO6B1iQ6Uqp7Ajr4crj6EExCfBDKhxhb7y7WRUWqU1OSv9zhbVFr
H6AzdHSFf8pt4BpdEPGXf5VmcdQD0sjK0+gSyR+dywdJ94J9V9YI9T3LNYIbASNU+LxLMq4MOXQq
i8mR4dx2OdAjAzugfNo0ZHNzXUJwSdFKjRCetJFu/Z5KY76tZ8yavvBYqG/EkGVcMTL5mSgfz12v
VNlk0XAgo3/lTMG0K1DDuK41aq2VFSfihLNUkuXAPEd+w6f6JlUFS364sv9/hHCZeT286TGW2qVn
uWrhzRzJAxcVteelohmjHiiSfLYm8LfIXLAaJrr0amoOf/VFPE9M89MUMODMB/n4opaNjehuZJEr
i/wPHBNWjAQza/EaddFI+P6LtoD3gUNy1y2V2Tr8mrFYqOqkt002BEV4c5fWUPoOpG8XKPuvwtDy
46VVROhrzrS90WzYCFXTfwXTgY5DmJY2H2LsoAtW51riZKcYkFkeinSTO+pZDCDRYlcb5q23ikeT
BjEzPyeItXrBTnJ+MAZaiwCXO3gtPZa6iX2BKHF4xAAH2glb9HbaH3EKRrqTWqLgobjck5XccyL3
KwVJ2pfWHS035waGt0ReL6sUh5KqCpjUQEr87JawJ0/cjKSLVM3ot2F4L2cbDyE0ePgGxkM+tSbS
4xbYDFl30yhoffyOX1+NB5j3bELP9DZ+D0qew8sIowybvx0WUFFLQdnyF06mg4QTvLRDYfOI6lGI
yNngH7fttdapSJm6SYY2bjoQtbbuymu9BnjeJSXYEotTMdP88Rw4NZo3S6DU02jmmZr8i6YRAuVN
qsdBQBUwN7Z3QAcix0I2s0Q0AuX9YCp7eGE6SblHlKzvcemE0vWNhv9rRO1a1p1codMZnXvY+uD2
aP20cnGYRvXV3iWrjtZFMbu4NB98Qz9WIbLlrMH2gnpYuqvo/qk2ZgHP84y2NVT7U+bE0J9OFc1n
UMNj+qFJv+8jQgpmwvxjS0tUha4dde85wfsdIS/vayJHU3yQFWRy9htvn/0iVHKZE+JhYO9mBnbV
GD7u/ipN6kCygQNp99seS3hJa1y0TgjbVUWXzNWZOFLCD2WjXKNcZvr2U0FQFFbXHBsSfWXLfptl
MXDqecS8vpvJmgguzaa1MExraGpyyGYuNTWBUiYDcfUZwhelCZUnRbp0iSDOl8kfGvwkV3sKN6Wp
zYUH/uHwon/ZYS3N62E4R5hJ5UrbcRXs+62rFzgtndKqvuCGJOP2MPO0uAooAx2QE3k4lPELX7kQ
/ejKrcDgIGR5BflS8mPaK+BZJAFNulo0DDmTAtlEgzgCLwVahpze+1xSHeRYZhIFXxkQD8dWvMYa
3pzT62FTW+DH1MgNA4CenzYFnR43/gIrik4O7BTOqn97UYWzJtvFU8zbBxhp4L4CNKHtFqjGSsL3
intT8ns+uwT5PudT33vEL8ZU4KjS+x4hTQO5O6dxqZGxGGQUvqr6/FFtrdXvpAKdqdZ1STFctJXS
uD1EVVKWTVECDujGhPMzwa8IPiXVyinW2iKwN1Drrs1s8Vy5n5ZOdtAgPDmh7pWN2nB67KdU2tnZ
iAXY4CsV/6NeqPv8zG+PDOKFF7dI3Su2aCqA+PaY1U9JAM1gro3pLNGscv1v44VnUW8K99Z4iedU
djXrrsrl2wqbYeIc3rYcvzROK8G2hU2smoRfIiawSVzgRwaCOUDCqoQ4jMmIzQeN4LxH+gXu+tdo
DbttOXS/O8S3FKmMor9ENcSUVzQ8pIj91F4PQChvtKLO5e1b0DM+R0SuS9t1g2L8gCC7Y6uhYYdr
PAViXZpNj6aL5GaH4Lauc9rZC0bMYwVgn+FBWuL7ZWD7oesA+4a/orRiZsv/3GxRCwTW6OSwsP1w
+EuTfDgs43u9YyzocqTmpzQblYybBrpCuXKhszIjCdiAYyMu9kroIq/wva1wrJNgm82M25cAqkVj
camqY42DwGvxKu36JBwM72ysNO4ZF3rqotZGKh8I16/EOSxdHZDgT7ZRKbViUV0g+if9S2DmEFGc
xGhdkJzDD4WP85kg4XAGj7GL9yO0t7MtJLyepoBQvKCKNv2u1WijXit3SvcrIcXa/rT5vjOW5xtp
apD6Px0N8F4wU5RQxEQiBKdEJpAYvvN1bST58cPKMQDQ3klzRR8n/BiSNLA+kFmXn8bLl3BI0EKE
PYm0INp2ImsyOCbL1iocGBYZOkRn72FPP5hkE+TE2ZJnlD7gEhVh4qmFoLCutlRO1XyIjwOWFbYh
ajXBk+W/bhE4bkDoUyOeQoh1mvdZOigxep23GcSUPN7PVM0Mn2Ob2HI9/N4Onj8yuODdE5LPItBD
0OJWZuCDnrodbeSsD8Zi29F5w4w8sTe0oOZtad8SEGjaosrCHuc5MSMp7deKEOI2ufJaJW9rxTlg
2WBLAlym9pCmobWBnutM6FnoEV2i2dSwMekV7Zv2gBPsA1K2z6FpAEe0ml3IqK9jN9sWgl4nFS+z
+6ijUODpnLB9EpFeM80Qnka5oRpcb4sKQPiYPXvVfpGqTLT/fNIqiHpVdB5SipphCgi42pzI7XSY
zT7IIPTbIDowJiGRJ0YeRLkcYA6qAz+5xsgHbF0yY5x5LC37HvacoHq1ahXZitEV70kjyIh8IsOJ
mWu30ifpzxm41JaJxrSyd8klhY/8j5Wo8EAbI9E4Lgoq2H7jdFK2YU2rPZ40HWgGXvE/VRtBLLbW
hRVGyz7pct5d34wR7Z8/gp8vsVVWJN1kwuNK8oVM/ZLQNACE5OrG562fDengzogxIBcVAp/Dzfge
CVdIOmKtfLt36fnaciClxDBKi20Gek7g4U/ZAEeTYn8Qj+hmkwJwbSYBWikwAgdtBIlN8Qb1gFma
6YP8g6NBQUFNeXnjL+KThB20pFLLtVsWg22tmGvVC2S4Fp+y8x0uvW/mwYkKkCdjStLrMlKYD8dW
IhXuFQCnuxIpkD3UmqwbhYHUwtwKKpoUi8xGax14MPEjkIjmyDH95BP00LcVbglQEXbR0OzCpOD4
JlKO7UIu6KFSm6raiQolweTSoT2Z/LZBQdvXjldkhpdcDfIVqyPMExP2Ob/8P3PcY7a3xN+Jd2fW
0YgRQyDOGha/rYmNSm6Ql5d1M7ox9J8Hz9oKZ8naso54oxIpCQaY0tzDlRuOyp9oNFgyxWrNaI8o
PlDzIeQB8AMSdai70WpHRf7d0BVuxbnA+socBgjt7zyuEsMflAjkuAE07rw159xz30e41c5uE5mr
MAyLAI7AaHkKPEl964mUewNlXh/qvGIObsrqy3+Q0vvNcWNO0ELDm1kYbPwP3NbkW+ZEc0HPy86M
LGM1E+GSC6dxAuPkjQmi+gbf4Cgs700qlh4pXYxcyHhjLvQQLkbMs5bHtCOWfMrua3Q7lvp2nB1C
l90hJiJMENICANCZ0PjCdi0fFitjeMfkQl0FL0XkLvpvsgHrBwmcCLsI/g2U67O5gbFUiZzTAtOz
efRPhPKm1DSlSC/zZykXQucX2ne47aKMD2qCVs4wgxm3JYZbm23hMNRvqyjdl9kZX3vdnUV4rlKZ
b9hjpY+mcXhSDPryXid2UL/MMedDjpbAXQpv6ZGxwirT/83Dd0o1pDUgPVBQpuYxlnSg9oQrHmji
Ylh42zR7PY3o0ko/rGaiHMHmOGBGad25Ph5Yr+lCBCPImEZwmy2/0hIGjK35jpUPjQ2U7DxrmGyM
SqtAD1kmkh4+ep8EEHS/CCMiGSu0/UvzrjQk+MtOp7bIfRHhpnwCUq8NM9aD8eLAbhMhjEACaK8V
ajSUUMNmigW6S4ra5qvVGTd9exSZ3Bgh+b7TPB9TpUqcxoPEYTNs2mRu8LFbcqQoLhaI80JqVh3k
ECY8krArnb7q+onoIgsdF5heMLgSiisG/hVVo5rYzYyY+vL/c6gyOvxdXwlqkRT8RGA0j2qpb7fJ
ydcOks5GV6s3WPpjUetexPJmsbU13rnfuzJoxAQA+AwLU7i29hJD+9/+C1LzdvXY2hVCyeiAoKCf
HttLNP3VMu8cVEcXP0+dhml1tgEIm0VNG2zv2NS6B9MQ8JF3IJ/B+IwBBolwBAwybcPi0/PM/Asa
pKA2RZGq6I7dalxQMULFOo0vzs08GT6cr8v1eCI3guvPyI8SbTSImL0qJVZxPuuh2n+wGjYjwFEM
OLmmEAYZxkCMQdj/iHYRPks8H4F1iN6uYRvg2cDpFItA0t5wLhfm248CI1nHJkZUy5dATZZx1f0B
bD3tj455M7xNvNKI6L7L0PCp+EH9+t/Yp0URbZ/L3CIk9bh+zyWSqLqXc0bKKchUyhRzL3h0UWMH
HMtTrx2+iELan4hw8GyzvblTrzMyqBGmCF7uDZ+odHql0Y+KjtuSN22IRWdmLU4VcTpBXckIqhbP
IRw2dJcluityUcOqeNNZc6SCkwWQ2U+3y69EQXoYdWSzyRbA/Cenc0RqNbp/ZpkQx+QcPg8l0+gE
WnUioDzwU0KMAHKHFnKhZujdrbFXhpDQlIYL+f9O7j7bmEl54SDLS1V9yveYOv9ateoRFogdhenb
whLTd5BO9BWcXOG/IKQx/r6DBzOBPGAkALe8C+wxW5S1LrNXHWhdYPVq6kYurg/EHo5BMb4zYtlW
NSO3uhreMz5NOXYk6cLtIOrRv6uc+XL39zruDTssusvE8eLqBwupZ8lkn3RwEB3tt2QJ9b0W6OUk
PDud0PtYq+w3khifRxR59RUQNgmtjwlU2hCuQy1R0Saua5b7dSwZ+ENF93EJYLNxFTOmwlCn5/+K
KBTmUWnYIcLp9LxymtqFV7xhmcG2GmMxkK1nisSliaWZgs4hbCpQd5DQ4mVIhr6ZsngwaSeGzMwz
gUe/KASFNX1a9TsdAOcjArPJo9qxYuelEJosLHwysoUB3PH3Uz+gH6qNZoOffdz5YUM+P1NtVEBs
BRpKVNAVggNhZwGVV9+SlDMJnhPuoPhYSj8Tfn+1Ge8IU6W4ql4i3wCfYBq5OYe2o2trNxN511Oj
GV0OKFGqpYLWCrEyANrOomvUTTEmwi4QO+uiWPdRssrbRhweR3Kidw39tblCZPw7o2uSOYEaI+rq
RVBdH6bj/SR7/Cf68DOgLNuuKx5of7nhEAv0W7iBBMp/sPaf5xMCCp4j668Pf+7eTqX+bYnF9Lu+
eq2w/wglWNjLlqjy7UMfmDojqme4/eIDZTYCPZusjYhXroAq+y7MY+9DHgiMyuWYnEpa986Uph+b
P3Jo3/LYfwXs82X6cK5bQXQNGcGunH6ToWMyrhs5sFSOra0KfcMXp2MnxJfzZhftA+whMIoTEqXA
wsBvCh146RFmF+SR1XogvnG+l8VoJ9DjiWFAsW4OJeJwXRK5myho6rW7e36mWmTsdoRiG85oB37Y
t1olenAupo+EbTNwDydiSjhsS9LJvgTc5yetgYA71rpa8oGJyDugB/van6UCinb11l3WCKiteh77
ivVeS/XT6bppNb3OBwTaNJyYAYx2RhbJwiq84w3FHng9k1rRg7atDNPlNeYBzGwRKg3+EgJ/a1Wt
KW69WNomL0Mjl9io6akIYTw2uFEXDGfUd7/AnxyezubekGRdXNAfhxN8J9vDC6985XAuq2ePjzY6
TB7hZSezdZMcW+kWyRV40+oxmqubpXpRTVyOn033IvLXrVZ8C+SlkF91Zxp7aPK17H1xQQzEBRJp
e0IBXvvPh6ILDK9xBdKXBPJHx8/e7nHGh0wZo4DdAg9041/Sq5r1H1xyubLhr6/SioaPBpX6YHA4
75gnQBKEY+rnveDolbxgmsje4RZNAbxOa1wQp+LHNUlCjRt9s8C2gL3w8GPBS227aG9qfgaFJmSJ
Dc/ETSj9Hm/n3XxRworcDV5O3TMz+3NxtmU4idfje7v5kxFFmsf+gA807llpi9AdF8sfMUGiqp5F
lr6Cb+9z1UahiEtgAUzgSt3hZ5zQ6+k97yi8TDrFfUApEyHZXcK3C5UfSk2QaEae2k53TzJZuQGI
fFlDwOX4ghTB1XZFqKuf2XYBvTI/ShgqHoJXoX9uyINWK3GaAMaUl3ZiafHfRcZPuiaFHBJd9zpa
V4Qdg/iaXB8B6EzJRh3V5YuVxjgq74yA+6p1jTnYST+C/2N3b4fq6WvXxKvEPSmgYol3cNt98+GX
9FKwl/isuLrMgVQQUH1vrs6a1CRqI0GL7L4tTXj3SUku6bMOsg0pO0k+vaTUR0A3FC2YxlU6X5gr
+jt4UL6e9mTa7POaPTc9gq37PjIs0h589RLSUQoM7wgp+0Jub9XJwDwuU4y2TNXrDDLsdQP+jhjN
v80WWNCm1P0l0dzKQuVKSid+UDtU8pcHEdMfQDvqefIxsVWSbeiGOMX5ccmPQCAZM36VT21EMVZW
nIs6cB+NNtll60RrYdVtNwN6mpemcPgkbc3ugOVxvf/76QdPeqW6VYQCqmiTbYL7YpmC8lcHptaY
RXaejnUDDIWKgwpX0f3dPHsNxGTpLiF3VxZpGyc4rRZNTqmxfkwX0O5WvdsjnDEmE5YNWU+tbkrY
ixVO95eaZE9A75F2H8rAn0zXqruOe2f6znZIClB9jJxDiVhktmUidB/KfqVaoNIXPYFtMkSx30ap
y6yudVLA+sx3ZcniaG0zDhhhwK/McIzrpOsbaoFat+sH5wfY1pX58mOYnWMMrcGs8HgGXiRD/tHW
ctzvjjWxVAXu6GdU5ehNNpeCeLGewbNLnz8jkzJwTvF8PYYSgQPOAia2zH5zZslNMSKe/t6UoRUl
IEl4tZ9oMR9et4e0S9NFYRVVU9qZXh8tASqzcngO6FXec4Vu8PBSt8Rt/E7Vz/o9967SszQCbghg
2HT3h1t+NONuBp2SHeu1eEf4b81/KQ0mg92ZS0fW9LKUpMFEQLImME2UMd6vGwu1zRsYkUmqcgYL
PEbWgh5dbxLvbaoe4dTJgihF8BDyFfGQ0dqXC2wXHkA737/QDnLwWSyYPXKExu7/O38X/8kjQV9U
cyy38FZH477eMyH4cHktUfU6jaYEHyj6xN7MpDcdGnEVRmf+kGjvIPMFxBq3fjUoczxBVsOQnROd
LHrgg+juDpvnh9VsLZ6FVfwZLTCR88PQtgreg+wLwcgLEpG3d5N8aMxCan2AxAnSqShqs3JdVoS4
2It/FfQSfbU6/ZWsKohIOkVzo6Wt87ntQ6nY2QPrruiDWVFHT2klUMYtXdZYPBVECVXHf7tEP/Xd
r7tX6+InVQtmSIehMANRRFhihNtPoPL+TszmNQ8LfHwsnNeRRjbad8JNnCTO5+eauWKP9KwrTOX3
0FcdRIU5VLbADgn8sLuXExD2ocALB5h3+OalsH5bK7MrGc0RM+ywatE27JgufZIOaT2mAQaBbvvY
AcHAgOnd93Cr4VZBgKFxk6mZVSJ68n70eKX0PzAzod3+vgH6Ikb9WdlFxNsT6MjwTgudwrtXkM7I
7icysI55nygBD2S/ww1tvH5bdoe0B4YI0swD9a7rux0F4ob48c1grZ9PQlrLthkAgnPgnSk92PHY
CmepXd0wALD3dCF+cVBcPWh2sBxEwtaaPwCMyelmTNKMdg7gYq/uCpG9NvIzjzDlC+xrIZWtCg3S
jiM4O80/7MAbJELcBvGlTJWZ7gV80KV1Gv8CGMrhLyQ7hHsI9+3mmymmGA2P2lfxqixIuBmynVLD
0N5S4HlfYo3ADfTRla8vyS/H5MRW/akmvbBh4tBuOloYkVOuLWH7SH/RPf26NloqqwTB5pNAUAfg
tZQYEh1hKAkTC0B3bx3uNhDlnukSIsP5N0uyu9BK5P90hQuJMCz+gHjoflNEhuECk00vASUFV1mJ
19l62dcWHNsh6IsMkAH/v7NtmTtC0Fpi9tTprPuT2lCQt353IY8kWm2PxA8tprTM+nfQ6ylPA+rk
DixH69w6kREKwOCc9Rvx6/NsovxMnixWwwSyI4jOz7KCssi62o9hTnqSL11RfpUwAC0rXnIuyucm
VdfVcG+sE253OqKpSbTrECI9147u1bzvKSrif3qFeHahAD72kvKcr9kgEAxwOi2lN+gnfEv94Za0
QT9EkAafAeSCMbp/Tt2u5JbZ3cCJM0t8MlQnz7z6e/vFnirecOAWpauC3vkSNNqNLOpouMxm1jdN
H42uhLYZTvui0Qnt1rPASafln2BfGQlzkX/BG4kWCqVNgwQynVNdmlYAl6IyPA1I+MwJqSozrO9t
ty6NuhU3kHLq3B4zt/2we173z4gACxHwnJFCizwJGLSdIfri3QJUtqnobNaAl/29nPmTIArDX5tj
UIYK+7jvXWTIYbht2V2IiLqTwAx2wjhUasRLUF6hHUK7C7h/PwbtFFZDCKGmvbyZM19nn0gyMuw6
4rDDinZG7Ip+urKYOY+D0LRqJb7MbRgZCMqUexzIcvjAM6XdX3mD+cIf+9iAqZIVK5Z1WP5Ks5vG
XCRKxwcuwln7LSfLQinLRbU3stwfaRw7rMTSSa8J9lpH9VQijptCmbz8m5vl5jnVj5vRz/ZkTZrG
BbKZ2DAo1BPrwiCHX0OX+pXIP25FCPuSZOXMn37d9CzPJox6LZ3DnsMT1zUi0dMMiNCnYPZV8yDK
1blOKYOKqzLTJvntYpG8+oj9OYRF2WuBdA+oupW8uRBisi5lq1snRq65+gEYvHDsHJbrb3Tun0X4
LS8DIbT6ilYmKbu1mtydjFbxta3Vn0X1VMDs/x2xJhsy9T/9dU5fEZogqU83Aol837jMM7czpSZi
rDIUJ3X8Rt/sYpr3IWhc5TQ299oFitIj1JzBudUybZx8508xn0JzBVoRTZ/qLyJYe4DQBzrYC3vR
14gP+S9sq3Cby2YueyZ792jCll58tYsR35daHW6J87S1cqCgNLpV/vk2G6DaFhhhpZLcrNd2S6Q0
9TwWx/0CigVZo6r/tNMeZMcP075g8ZZi2WdCfgBusSppjEKnst+S1zWOc8gDgFB6JRFSC7/JhB3A
00jdA2BOQjDaNgygSkH6R0tAzX6KGhqLcN8H8gky/5gIC3/plxPIJ8C5EtIuV+QYFZ+EPCV+KjFd
w1J5U3cYBhfzZZwytQ0s3h35pvPno+3Bl0k3grhRQ0kyOYAjMSrGS9HUOFMldq4K/7CXHWAUToZr
dmhxst6F3V2OHuGSqF8FhIPJG3P6J764gM2HP+SVbxTgHDGbxHycI0vHBCAJkdrrFGNie/TIpOaD
jC7bo5xVmpCEBSIxo0M/Hk0FkQa8OLnzrqy2RnA3VHHXubfsBBQs03dB5VzoA1jwmd8GQFgzgmGK
8pePeQoIaKbJjDZvLEHd9IqbVm3gnv/gKhLmB8NPe2JEqYtY6uMk1kU2arGiNyjRAdj8gUOwap0v
rmGvDjYYlLiVg0WBXxq/xzd7QURYvNQN3yp5C5SFQEyEvmhawu9xr/Vi5B5MZWNqEOTNsE2ealUs
svbnSOG8vJ85wRZwDrawV5s/Qo0Jnn9ElnIb0hN5JH4QgfeD+aspBX6cm1bTWY6qF4/HIacYoEyE
vHryFMIuoFdsLRHnaLe4oIOCAtKhkIQ9bbLtUfODJpkRe7q9Di8iJdHiSNTS9WDhkVDBum/L8kRG
0juho7U+1IuXCXDUdiU+IbAtX+Kz8rSAF5f9DhTUVUgenFDjfhVs23LHO2iMG8EA3QOqEZuCL3VF
bdTHxYXUrLi5BLMMOMgTUfsYL+h8tqkQCWdauNT/QxFiH+DSRmGsKzxXfn+MKpxPGNYEo8OH8fsO
iF8+Ok8n/7T4hTThY1HFRhZxA+uCeH4gQaIkQ36EUunMqhKJFVIamGIw9b/puR7yhYCAVQeUHqbc
q6eCU3s2tQBUkGH0G18X8gQJVY0yUNPU/sByIQZFgdObY9J/27Tx5UWeDJTGyFQ7gXJ7Eb9c3KjO
G56ftM3osHvmgdIr5WPrMFily07k+cXsX73c2G4lq2w1VSTTm+CVfTuQN4GmFQ3kLhqlWaEI/7vn
rYRV3NAeeaMSxyYmbDX4ZYH+f7eRPS2OX3KekT29+eMz8bYcRhqsYLCwLtieA0L3Ewn/uU5HcLXa
mIpaIvIRGdB08l+mbwc3gYJ7AEggFisOxg7wzYskwl1BaY9ygdJ28HVrxez5hQSp/ZMOHjO/ctp1
492bf1fLqRvj+xnDzMcFHWAqNCkq6DY0bQlw+uXsvhH+rzIieV8h1SYv/vWIP/UMELwG7ryVRaAT
b2pufPthoLeDkh4p+9oWTbEnvqVqFWSUQ15dx77Q2TnLdwcJpaA1OAn0zda8Ch5ygjLCf0x2pBqq
orMVmu1kHVAP04IzaQuuf/6Qh4thFIpRO3kHyPzMkcu7dJeXH8yknKj6/o42jQdhlSYWLASUMxGT
/rir7U6cO7Sw4T+cgfGdwUxI0LHVa6z1K7AAypywK5HESmyqJBmOhlI91PQgbamx9PX4sFRpOzBN
PgCGzzvmAW9EzUKbWEF3gwi+/1sEq19LwZtQhtnJfAGpvGozEBNsFQF+7/pE2T3uoPTEMs5Jzzvo
DzGFoAsqQ4JkXTDGLtzqKzoJ/UY1J56tVHOMnbgpIdn9oGZUSQ==
`protect end_protected
