--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Tk4J7q5o7EwRS2OWzX8GDGJuP4bao2U6Z2FDkkAiJ75i5DvVncAdxZE+uke0uhvi+wmU4epCAYoN
/dxzr6Hy/aW8fLVScnFPrJKDNzUaUtnc4UxOW3H7Bgh8qMj5ZvwyAb1eOPm++WoIRNCWVzHJdx+I
JeUEwY9iI+RRgUzUG2Yp3nemQLLVU2a1tbI49+aVlBSFhWK0kL1LY2RuwmwlTT6wnzKhLrgueWOE
Zxn3MA/IgNq89GJMflxXlq/ct3kL3EhCw8ikoIC3yiDJoWFom8UenABH/2ZCCewku5mV9zPe5zYQ
fPvwh2PasJCWL6YMvQ52YQ5ng0Q4IWXcyesfyQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="JT6nQjl0mOA+Tbx/lnNZwLwqadA7qOiscve0O5Wu7to="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
NmXEjOU/p8UefIRLfj0eP9Rfc+Mg5yXKOv/qy8dNQvv3AFz73yE5ZMfh2ej8pA6k7Pi6D476Kbsr
TOGze1u2y58si3MrqvEEd7/0jbH3nF2X/iZshPFGKCG7tu//jL63WnK4ctOeuVY8kRZ1kDukcRa6
gNA2lsdpNC/1zsVBHmY4p4nhlYZz646lrAPjdWnE4KDOz3itr4k1yiCdAA/8kkSG3J4muryG7lsR
o8804bc5Vv9Bjpf8aNNz+CbYUivpRwcLkAQMgf9lb5TzSaBBsAEIW1rD8Kjq2vlwZhaiug9enyVb
SF5P9GFP/sOYbqgM3t5/cFWVnU1+JnDzmBZ3Eg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="euB2b+FvxSCiEysz+9hWxTfIsopq23Ox67xidpoSc2A="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
qiU+//6L5qUQ+b1ADoT78uc+qSwBehV3xYwAR19JjkxMGeLo6lq3zh287DP8NQjMWBnAu+jp0OXj
3Q6NoHX2wzW1fYEnAFhppccTVvuhuf0QM/z0acrMsRl/gYbz9xm4awxOeK2iSet0SKcP0uRNvw0r
2m5qDCR9RPrxNu7qkcYJhcBeb1Xy946QkEBxXcaZN/mHEwUf/8FttsVS4cvEiWRL4fUl1QTT+nF5
f22UxDW1N400euwgDekjUcCAkFEtNrViO2WXv/fkMHafehvU5w0kyjVMBUJk8BtXsNMPlCQF4EJF
LFFdan2XD638oc7umrhnxXBOxYAmX5MhHjWf+GKAwxPuCO0lYERNh6ZZSnG9rrPUHY91hQQY/knk
GhCCI3TKVXBIHQcabEJaL2uodhdsyx+0LJFCo5mdIVqnYENAsm+Ou2adxGgMHe0RO05kos/KoiMM
6Mfx6/Bb4dxCbOPDfHiuL6MJyhVmj3w9VBG5zmKFEMHxiC3576O5PzLAnzTgTbp2H1JYHRkyI6R6
rVWnIVbrqZErlHvesJY1jLCi2FDlUVd5UOl0Kx2YRVKfn7F8m9sQ2ubqP+Jw6u+QFo94/i1HM8s/
1DHRrRbxx4sxqFaWQ9Y7/nSa+9YNTepwgSwoE0IlL8xxZUnif0RrjA+96nfQx40YgI8hbCm74TDL
3po46pv70L4m1KNIspCv0zdxmdpWWMagfsgEa9A8QUdzJkXTsSr7QMeiEgDflBiDHXfAn7tozGBG
zjo2n6dG1fqTNszJQb3X3Bloem/fsxNx2t6yl73VXe0FJ8WlJ0oft4eCVDPvB8H8N3RzK6AFHwkU
1uw7V41/gRE4WL8rW5wgWYdLtDSvoM+QomBvaIWqoat1jXwUBsjDvg2jbJe/6+7W0GVWw50FFuvV
MdxO7Ib5FHWucoblD/e1rI0zvToANw19pPrEcVjGnqwLWa1ISsYHqevUL8Zqh6/GoEJI/+lhDjO3
z8LtbCFZIvSxjp6fJZobOAz9e9bnD0EO/RqAa+J9y+CVnPhwwWH0U71eT8oOv9kKE7GAjWr1qUJo
1wCzea8if6iLc0xExPv0PJW/NowErLwQuIFw3V2fiFOPL266yhp07TCa2/Oz+vPM18RfELeZhFg+
P1IbYCWL2IzpW2fanqQY6PbQWYgL3KrNjtVstK7V+Vv41XRDTz2J8ejyTIcyNRe5otmmrRWsJxxh
8D7Ff/RXMSStYaATYOR9P1i5Hz5+5o4M8Q+y0iAb8lSEtyhyAtgMEA3M8ctExXw9NPXefkzrfjyX
Dm9EJ7hS2aZ1/0OoGBgq1RAbJxr6CyasQwKPwF/Z7IuEjMCtnweW0GCPIhPExt0cvAdLT+pCs5Sa
d3j5l6vk/rcEF9TwlaQvMtkzVIyVC5r0jcdS9xGQtXvB/Kwryc/ltn/68/AQswgYAO6cANhI/Dqx
RgWA5XwI49KRtYK/NwmnzS1oMOpfHX34OopxaPGk+iOQV3R4mE/mWL3KkU8eAgImIpchujMTt06m
X9+kgR1VsAI+hLndq2o2+DWn5m/xMMPWZxOyeNlDMFkI3VtVqWH/mlcALir9Er7QA+qQeHfm5uAm
JLDD56H6eBOdoRokIUQ4hV19XEmGx/5rsiTu0oAhQOGrccnrZrGvAm5jz/WH6WBriiks72YpEVj2
hif+DNGCxvaIYNL2y0hg798BhJVCJgPmbxL2W6E461Hm/rVYqTouLqv7Hy46wK43PbgbHplrOJcT
KXJk4crOpLEpsl+lMpHzaFiHS9gOPIO87aYdx/Us2oC8vGxaLzGmMju3XlXc7FXsOMCAVK/o0xtK
wrzCzfscxoL6qFwYs0Ym+2pZLCBby/WVchykESi6bZQkgwB+Zf04pW50DWzrl1JSDqnRjEkAAqim
BbzArqLhCi3djRLkAyeLH+NliF5IRIxz7Hi0P2ukwVEw1sqAsTB9iIuxxHg5N2PeOLsjALcKu8du
pPFh7U0qsi5lOHOY8WBpTRQnb7HovplQzSP39LmakNzbuKdX3/SA/MyW7MxvO0YowKBOo3o/W9qB
PODNvCGTm1ShWhBNDwbph2NWrNGeZffNhyFRSkN1/mEW8ZEtxEElUTC2dobB6+hZepfAl7UqfJTg
SKU8Fz09/RB2RhINbc/8OlvNJTQc0LFiyREgnV1m3C+V26jp3wwWtGz0vS5sDC14mnkhSbZUclVb
J4gQdK59COsXjYsOuJag8cV0Dyn05tMLRL+8p3d/l29NA9wfzt9ZnPDA02lUigQRUI/ko1Y4NBep
RPbMYxpLBs9gLvGCrs2NmYIp3zsLU1RYrnTq7c6avPImaNj+Yf1Mrgrr63cU0pKCHeGsUdw6vpCQ
dW4oC3UqSYl5NrneAjS9hu0hKrkQskycX5Jg7Ls07YY/Jj2xtHtccJDx00Ru6opWlTHlO/faj5TG
ffLqynW3D7TFVvGMDoK0zRQN0qL24h3tsWkHFG/ISdq+zHZtwOprHh0zx6JKdU638ISKcbgOxsvD
S2ntsXzA8VnWRsEDSuFKWfgYfrNNEiWVgmO4bfomED7o2FApJELVzV2FgaouXY0fqzQMdBbuc01u
gHlF6ZY1g4zauLn5HrALVGKKUCsCDXdIZeyuQPtz+KLXif3qX4qY4w+3rnjKMn8j9Aq1HWnRwzck
LtO4m5tlh1syRwjGLY7v78Unp0N6aGd4qDxLzYVxBuQYG7EOfutx6LN0VHqEne59Lvc0BjkPLuWw
3e2S1I9mHGCt5WwbKCQYGHxv/cyzZ/pc4/AHBameG/6cQ2XUdp7IdyVXbS/php1JvvRAIGA1ob7p
T7HxhJon8NDFXDA4NN0QWPi8YWA4rWvHJTl75uMQISFuQc7m0vwcdCNXJai2NdRwjUFVGACz2s2W
Q5jnZAaCTWvd63FsUIYDunDcwJd2BRO+XI3wL6kUcmJxAWkXIPUhXVgnvHNxd5SmGdFfGfkEqHlR
aGGGH9P+mOUkzNZEpmNdjiad7BwL8tyMeK7MfjKAP3s7x+T11F4VNpCPX4ScL6qZqydWyJ1vYleC
urqKPjUw3VncVADoCpFp6Zg6OVOzyhe0y8uzYkUT5VcI83hmlzBsZI+vb7Yq90+sped6Fxl7xCZ9
gXQMPFEclCg9Xbb6aZLEx/VK0gt88fy5+Wc23GTcP8hkv4NYoQKfSG2D5DJk+z7ZdT322Ho+gk6b
IdJ2WRugaloX6cqlEgrcZrnyZsJEbWFsS0LlxMRn3inDya/+OoubedLGzgshrXx6IRY5zgVjqSUI
dB1X5nmIzLUbsR/eKdDbxNcUg66ttcQ2+i1xRkYnYzyiGBA43fVAqz/WANhbVL7+ax7qq52FXQWk
6sy9NZTCjjxexMd5Q0ipcCMD2Hp0REQI/SUNK5RmNI+hNmk93mJpY3r6MOkaUA83hlQp53f2gmXa
+slEzfk8SzIAjA4CyNSyTz2OjXzCVYIHow7RdJ1hg6tOVGA+k6bveGtCYFQ+SPdDqcCsIYHo+FdE
jwR/FHTP835qbzc+l25gg17IX37pLgxlUUeMWp0Xq4zVcpX9MQIWHZpfEm9rr8gGV1z8CJ3Zqk5l
LGn3gbXLI+MFFexBMh5C0jsNd/H1QL4wEFnAwcyQdDnipu8grnpfh3ZJ5KlIMhFPdiQKNFV6u6SW
OEjx0LO4tAAIs2a/UeXfpdGeDF0TaDirxP1ghlr5OsDBlhMAMIEBOvEmX0g1RFBFnuRwcdEeymRl
yei5KZKDFNItSfFkfdZ04eSFd+g54mevFp/XvUyma+6dEqTEW3BJVP087k9QIx5GF6t9IaPfsoED
RBgrfWB/ispyzEwSsJCX1sc75KzG917VITC1mA2olG8Y43UU8xvp9hF/9KJzKnaLUH6SjX8yp6ln
/VR8ZkWxzY0//dgytuJHpiFz9KCjL0KfHOUQZWYfGVLJAZ52T8Dc4v+nJt89Jhzz1PbWdhSu88N/
zPmt8YgE5RjvXExWpwz+H0F00PHgfkDQinzVY1RdCk0L1ibT3fx/jqP3WaVrPtkOpBzk0dReDqCy
NRaMCsm6jvNfUY6JV+TVKjuV0jPX1AxogRcWIxsSUjwNVWP0JlbHPAlIa0bJIvZ07yxZSI4EeHee
a1kfXU8z+si7XXrE1LFhDsychTJs8/EeEVaEmMma/cNrxy9u7nM3BixifH/7nOTD6OqRrte2iT9F
zyy1nuvE5PgrUla1Teg0Y3MLmTK1syS4Gc2OGbwq4HQpM8ie5zY4akqAyv04oicbcMt/wGZmQ4n/
mHrRovfaMZVUQFf+vCfCuboFIbLt43cOFhu/3d3FCCVds/NTAT8DWeqlL+H2YWY5PbB8FsMQNe9Y
K3r7UhKMGwtqRrs6enh2WtjAOmg1PeDEuoaiQpAVBeM5r6yyt1DTh1kA5GYm6Uvy+xvMjGQLpW/h
850GioH7Q4XaibvQfnNiUgwPHbrlWI/ezVwA1Z2kZhyOEJVrl2PL7NGUoC065dccOzow5eEn+SKe
EUo6j8zTsUggX587E83BGUCoDi+Zzmh6n4OtuswzxnpWzG+/A3u9/gRySc4WmE811Ia83pAcfoVU
2gMkeyySN11nuSgQDrsapyBJJeOt/o3ZbP92biU5UWFL7xX8FXdcaW9ZRTQnZWYYaLFpbIENKDN9
ng1wiIMVyJdLbGPVEEsaIRDMrZ6Cja2jdst9/G6t92DOUdaLqB7K4PSgvCH1LLKuMwRfhsCiW+qK
UvtoDVUdMtPN1Gp5ViGV1xyVKvemjlPlORhZ0U+j+BTJ6/SEC2hWJdGMDvLsSN/fFZk26PJUtmzb
oABFUEe7mhLSsXtLXFdTL0dbbFYmNIaCqNL5Znge9Muutq2gZFH9A9gtSR8wQ8LTpShaC68mWJr+
SnXI1eO7k2BYjp/i5CBkRQn5u2XGC5jNUcMWGHeYxOjxZRkGa7Lq6cWYAnGVGEgqNszDB6DjkCr7
hCu6EVbeOOl9s+l2KHvn2KEzEyzw3Ydy/Qjf2IuzwEt8qvQHlFMqayPVaUPfTHqVN2lsZXMPXWo4
WEUzcr0XIs3R4zy0ck0aZ0F0lZN8JlASZAR9PBhKinCtI9PvxQBNeYfgrTkPHH3iqGqCW78VuEjX
jrwgB6nk+gDr9d9gD156WIoybMRWQOz2YNhi+LSEHbokfSRD9sXZKXDXZtYnnpxXvyEDBCVOpW7p
6rJ2eDXZwht4dH6vFpFQTdPm+JXK2C1KylQ7ARNid702jrqzQRbw7sSIrAkRAgch/ShMz6AbZMMI
iNTG4DqVtfoxVsKop55Dz/2wED/6Yqhbulm2kytR6T6YE6WOsuY7VLjA0Ei63GW7IE/COjU4ozo7
RLDi4TMrnGIGULF+1tAd16eweOouoAWU+ZCDoyzO2QSnYk6SbLSYjNKX33NHVsORaXYef3EGJT2h
wl9wkLTWKtY4usiCujZqMWzCnDgEsGvkJEPFt+uheLX6L9dTSd7V1cbLBQmUxht0S1oPR0DKjXXG
gjJz+VOH2dyCkfUjh6atJMN3yIfOqF0PeFFkqHt6Uo08apudbRTbn2RYU2jRys62TNjDjW91jq5v
BUA6tWkICr57Iaj5bxJhNF2x+JK0BqQCc8h7SqWQkmrlDovNfAVWWcxNg9gjME2jsfUTenrjR4As
4it601r29C6DUzCvVnyOpRUJUP5EehrMmK59CYS1OdpLJN+L01S4zalSdtJgB24bSQm+9YdVd5TW
rIcHG81mkClCAJD4mNMlDEKfc2d9Qpw2URhkDxwi4w2kIyju8uqTNUY+alisw92I6H9vFjQ+3AGi
zDDo3HMHrVqToP0jSt2GwAOpjl8b5Po4d+j3j+QDHZFmnobl49V9jKwQ43Q0mp8YlXrupVeliY27
8KhwrmbPenWou4a1h3Kv/4ePA8ENH2e4Mkmf4PlYTtrygAivvrw+etUSeMUGzqkGsT6TjbKZuH/9
aYpsQPikQ44B7nUQIGSQHYmcPiEQt8MfcwrcRamcb1y6v782ra/piO5eNPTxBKGiqmYpbxP8hxtK
OaYNN5svTW5BH1JpDgv3GXo9p59YhWAzSZJKHUazVNo2YeyEaFpUcg70nApELvqx1k8wGYgXnzK9
nFNAHDf1yh/6g4brbDnVy0bGbxesdrcupZMBCU38IcY6fTH/Tuw6h89DAvQoT9XDzoM0zMjHE1K4
2UvushqR/pV9TVbKwebNdbGcayLg7V/BeBpy4H19Kr79KrvR2ZnY4o1GwekXWf4FweXtTzFotYbh
fG2lkqxbmhONBJR0STzFXeSyI//W54fp5QsaQNSQ8ZT7cShRQK03S1qWUojw56TT8nYmzlxp9PUN
NbcSLgHhbs49CT8a4RB8Sxu6o/MPV2lM16aiTUOjtH9zb8OjYu5EClwl76E/tWawJevuaPufU1Du
wpinFdMejsN9gop9bdp47OE6hCTS3eyzNAPiMwcUh5iiiwbnTxl6qINSPKach7NCFcrQqD9Ou6AS
eJVpFgDKqN2GTXq2rxdLd/8DKe9szkv9wA9G1KXl6be+245BQm9xLPaDqr8lzPyqWjVGNBeXlJlt
+8r5bzPsYUzR22IkDKvYYOC8S8h/yRZY0Cz6J2ibmKE4SOVV/xuAtss9bfrEQGdn86Twr9Is1KxN
g/OeAGb18SSzYv6Kad/RgWoaMbA0dJl1cduaZECBW/gwbkrloUsNnk7n/vu+yOiT7wRSx6mpQSPM
xgvGlt/aVQiOCyugnOc1mXTKveWfC6kJbbBeK9f5QfS5890RHNGetOhiJ/O6XFEI4cHuzVrPZSwV
CEOKYz2z+ygCBMjS5d3L0GrimXAKoQjtWTtvtg//lDC1FwKqqfeSd1wupamsVQiKz8TVjCP4GytN
8sFfLLUAVDE1WfnJ0rqrXo4z/P4spm4Ig2sf433bm0FzcedTcPqOcCV1dnJJdEWBbRZoM3XypXNp
eXehjD3dDtKqB2/HVSw4WDU4hpTqgmCbxnm53nwYpsjvaQn4QQ4ippzmi85t4nj/Vca0v2123J0v
/4QZ3FCvvMIyW+gZI+Ac80jKO4fvwg6uYmhCGbLnJVDioGgOT5CXQPVFV91RshSEE8Ux2rMfXT0d
foZjDQFJ8MG+UOc=
`protect end_protected
