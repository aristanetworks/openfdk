--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
F2p6c3xrOSnluAMgz8N0aYai5SevPsn69VyvAPSgNSnO5/42lcYMyLXvNNydCo7EMZ3BEn1XgTEY
cVA5qgCkVeS2ytixRvD9F0o6hI2buDkQ7cbkhFeyh1+PyNTDnMVbt+IECNK1Qy5i6aUeUaFMxIdz
JlF5VgQOOtreFyZSLwAu119JoW89o6tcLteG/MYckLn8Pws4NgPqqJgAAgeI+BX+J1AKz4HUd882
X2o+JAk6ShwRgiuiJCw4FmBcMmuJXgDn6LSpnAcbAelA6U1UaIQ9L7gUgS9iBbR+yYR40UsTSOeA
w8MWlChtMYKiFeVfFTCH6ktKJU3FDs9TFeJ4Aw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="qExAysT/Cy5dRE8tmBbiQMNBnZK5Xtz5tBrax2j6Nak="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
RQ7WTuQMhxjMST89Yr9mFq+kp0F+Yrv8FtnGCZD7YBwoObeJOh9p+E8/HIskItZGx6L86DNDK2+3
RzuYP9mvlYRT1RTE0/FaWa3TGiCeE0J1gO1C4SfF7yNqxTgDPCVROctgI9zhHeN/1/yiSh+WmZ3s
d4+wvWKjpAOZ4NXpEiJnWSxhNWn4LtWRaZv6pyC/6tjCe0wIcV77n+JAQ3jJX7g5ClyXhmxcoca6
JGzthtkLaWXra0P20e88Q4ga6YO+4Y9PNamI6eT0IvBcE0nyVZL+Ki/E91YkcRJtZs8RDPd2vDm1
RjHtJyPzjALGJjRJAuaDaiupNXRTaqQ/fLDFAw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="b01M6e8Baon1Tk5a/o1yyBOnbmUs9CvGefVqpVZdOHg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15504)
`protect data_block
mYSly+PTPV2Tq+WuS3zDlQKUPJqOE/N5ZDQf8xBTT2GKupSlYXD+K6k3z9ym9GI8G7Yf5KQtdg8a
Senxb+T8GNpzsTi1fWez/fINMft+qtMTKsLpP9yVK0QvjbE+ZzlW3uXS1s5VBbgUY29nVJA1wTyD
3lI8k70pWn0qX0jDRbXkNgw6IbKZC4N3DIqA4Se1sw6RzGeOZycV42W09OlRqcTdJDQzeXGX2w6E
dGROZC9eiL3rucnKbke98ix1oa8BIyotUp4VAQUdRCVcq3N69BfgBj4fy0MyotVPi72rrrxSb9xk
MYy96uYbJYb62k+ZklwrvoCbzsFDAMFdjILhYKJmbngpLqqqtM/+TLapxCrFOQxbvZMMMx53MpHH
cwhnAcKQHqihPfm5WfBn7gOcV/5p2Gpna/CUWq473ft265a9h7HmMT7cacvRYrZ62cwhlnRxsN6P
p91PutNsnINzEWOdRdyGkc3F8C0QS6YHmMT8HcPoZTLgnT17psMNFctNMZ0YBDypH16AT8LPBEZK
aj+7+uS47VnzuZn5wnf/NzsI46oCgHZ5QASb+NZRzTmokNRe1SHcyXOVpFA1wxWy3XIOW4Vfgjpw
4/1kv4XxEMEXIiEjuIGswVusSdlxD/GXuAF1MViVfug+G2NLK25cq6mj7+oSkwX6yEk9B3+V3qxR
o6UJcgMcOXDcHl+0X9xOFgWSoLSM58fGeyuFtvg7jkoa1Z1m3HS60iEIbAi5FSlbL9TrpNaItxI4
lvwUXhUIbOURo1g3T+CFLtLPmLEGNFOGs49VWXpmJn1G4dDdo9EsRytm9/Pn7FmHEqeqkzsBqGnk
s/R5/jpfslAArYJxoOptQZfa+6iUxPSEjx7xQxKd6KmHwRSqUHcBpVxC1RplX2jWhvrltYcdpq/A
+ruxpeIdDOoLRorqJdFvCWbPURSV9t/qg3C0QThflbNZn6BrDmB+YQvEhM4PCZrtfhoYbc6RkgNE
L0W7O4bygxwDnfkA0pygsyEn1sFQCelkLqmlKt5/WMynww3afkysC06Vi2OvC4XK/ZVbvIuL7ax/
fbMAFCLObxMPe/VkAs/AeIHRH0ihnzaHUz26L5MdxtenWxxv4Qvm7O9ByCsJjLqpDS9tFlXYqwHR
T0wCqQ0EIFr+7SdLvFvJgchxQLRPKgzevwchH+C6yIyFic+E4BnX7LwwiMUiTDExsgsH6Z5eXEVN
D9F8cleWVgDxAe1irzSmwTFpkejeLxnp4Gisp9SMcebOWNItT/1gRE2VNfis8q7l2KjqCrTXPFug
Q1EQwWeVnoFvHgN6v2yESxm8Ec01uesTzXk88pnVZgyQyR2q99YAKtYe5yVbHg7VyYUoLqOSBb59
OHEjPdNcvytCIXd1rITzwLGJmFUTGZeKYaM5yy6Y9G6fbMAieP7Fcx7tvs3M2g1qzckQPfmB7jrM
7xeVfPdtaDPKdhq+jZ+1ZR7F1WCQSByexy7aVMYnMbvY5sz2gB4OLlA+tj683/VwI7JP4/vrCmYR
/FMiplAM3wr39Omad4OTgSHo18QtyhLf67zyAeSwwfBzFb915ln59oe8Y+Bxhhl4k9F0ElfMv+rJ
PrlQjdSCY9hMkiYq1Qhcn9QV0CzbHg2TkN4lh3FU+4OqqE3Vt0qTCunZ/MUvRX8o6nDTql+0twHJ
gTr30EryVr3MT/WaKwPSBVJVnybcSSCyqN7emFPAPEsjbrOXsInzZHevtV5OpvMfz58hsBQA6iq5
quOrLxuNSzztWQie+OnFNCM0mSRmi9yyrWALkb1cEsaQHcZgfHefqW1DoasZNovBs7WWBjjlxfyz
IrnMEiPCm5xUAOdNzn3evmOvg1OYt+EVFeuY51FEo7wjCUowkUiH8QPxxWrg+Gy/6TgO3mlkiMbv
PEQ2pckfk6Vhy5MK/pXZbYqjecQL8lySR9UyQkQzVt5LPRykx9pfd8MGMvCD1LtNDkGu8ZDQ8cIZ
Kva78EOEAm3OQmYMC701y3dGL+xtg+ST4g1/BtFBDXSEd/74XcNpQUW1YaO18OLYXp7I2LhbbWvK
E3Vc6+/+gvWq+a0YT1B7ALxVnZbbrbMhD8IW+Wt6OmH5tMfUbrhAenEalCcnd54gQSIvRJtqkGju
1HvW5HgmF1/hrt63IqWE+R3M9/izFnRR8RQcsONczEvPXs7PqhM5b0nX8Ea9T8/2M1vCwIGgZv66
Yh7IueagpRc8hQDJc8lmwSgLA0vp05e6vesFTL+FoP7TNWKAFq9UPGXqdhpfy3JhtXJqpg53Hon2
gNG4zIpySbM0+sJUw01j4THxW59sT4aRZX+xSmrzFsasK9MvYwGND+QnG0qzQitsXYt4foZzKJgU
DmiEIe0KkOkD2uLWq2pwfqSWjF7CUq1KX0CKydp1Bn1gkPwuWXqKhZLjgWdDOh+93LxI9gbjsVUz
UAkNhaVmR9zecgUELZSoRcIgtfG2QaYEEmA2NhpRZO4PDEB04DOLwFoPwfdFlSsMv/19DXefqKnj
A5606mRDkb6572ipJgCpvSW9dEWU2fySaPwZjkbvLMtjdzprhetkJ6IvXLnQmBBChdG6Uq0MbfEK
1nhyd7fURbnsRDAm7fUcFLzbWmCi/pNRz8iyX8oMRcoN4EwMulUMiCMFItZh0wI8iHOAiVV9JCO5
o6+Bbj62akkoJwt3cZXaTcEfXeaRqjeMRgDtzCaOPZVxv0ns5iKWdJtUJh71UhV3DN+OlZpaXhim
YVDbGfpH0iTr47sPaG80yzTvjcq+UVx1K/9AdBnAm+uLCWv/Q+VwrWHc7ovmV0+dXyzp9IVACnwE
kup5nxPebtHK5cQg/2h54D9437z5LrqO+YxR+ur8JzAGXLP95KOwoLYSnlIGQd7j5FsKlOchn60n
QckTU2cSZNFarpsHKXqxkUAFGdyDMcskKnuld7Mbs0zCQg5hR5fn7kbInZ3cDAA5baLr8M5bcxni
rs1TNEMBBPdJHwvrJNwtSxydnUjOmZiLnS9uJDaL0Jxzm8wGxkCUxPIsMeXzxvaH1KWbVWAo7E6/
kHoqkcxp0j0mrgjQ6oU+q5ai8uHC4lDBogifYMRBRKcKNJKUl6aY1xxB4fFPx8pUVELZhxi3c8M0
gObDyFWvaw6otzvpY6sCbeYaoUlxmGyeUAdpkPngKMXw1uvQWKV7a2IvQFDn16LX6BD4lbbFh4ed
6pyokabATMTRCKeutXzE5KO+8r61Ri6/Rp7JODRKSwRmrxwtXpGXaQDasS9fxeRaMSTyEX/52EXL
PCgl1ZYQoVIh8hrSehLZOLeDCTYDEdiCWvd42UbrxOUN0z8INmKl/hbfaDtYfAGcTPFMFecUxXRx
kLhJr3bsjkPx9u1szfez7Vmtg+b/Oty0Nh4o0WPB8veGGifdprTdpS8bk9Xlo6kkYa1/ZdDx4BDT
9Hm0vRw4iFc/Ni0LBL1JvlAWHtPvRxD3AbhjZ7BsAAGSQrvZpx0nUrknp5GubOqqPG85C/fA3PjK
vaQjg2mP+AH4fdDhhrE5qi2MNjNp7dvKtzmcXUNA66tvE9f/l3TI29q8By6Keuj/8B3up2k1d6sb
3R2geav2w9cAHRYEn18Fh1Mixia3mPHENqV77G4sB4ITzhp9pJPGojPAY5L30OmfjRigY9TNco7A
OWlhkYAy1uMzcyytems+Rfphqh0ucYiZBkkV2iCX5gvSZUkMoG8aD8qKPH0hWmskGQ5a+KmMehDU
ishHB+hHApbC+w4zhQr/+cOpxpuRfGjIXsHR9nGJU/ezX0y3ZYDJLdR3fy4DInUDlqXLUkC6WjNW
fTrB5UTEpjc3evGvSbZWohklQVlRCTnwTogenkmbH4ce/QJZXRX3vwvtTBK9T1bIW8hFpMdD51Xk
xAvpJ884FK1Sz+I3oGuok4nus2G6XT/Wcb/cTGtfbVRw/Wzaie2b+aNvZlMYFA7Jyj7gNjoC5Bdu
aMqlzT3jw1NrErl6qLBT5FJa9FPxAzGiJFn3g/6Q4cqjkoi9EIUT04gVKRWOgzuj+Jsw2Epf+z/R
v156964drncUScaHl6ojd4Rdyu1SGrL0Mm4/fUFbpHUru2px4tKQJRRjihPxG/yuZ7w16XxfCm4x
lCyG5ZMIKqgWU5LI3k6NAN7DRHw6/FX1eHA1oyKZPddXG1dYh2UDRNRYv32wceNbtW8CegseY/Md
qAkqeZhL49S1PMPFuKRHLUaXQktp5jhOLks/Kfez+4X36qAH75SfEUnfpyd0K1GUlzoqeAimeGK5
2vo/FB1PyMqYdCeV8SGE0v+/6/xNEN39dIMFVQPE7llaQR6WOB+9xd4ShKJ9CbtKYrB/A3vR83mA
S4guac6U7KsufJxyfnEH2gkZAHBiht2fcds2iSdV3187qYpCtokF/kiB2irXigxWwGHmhJyeaa+C
M1avjRLXJcHLX/U4HiEMDZcVr1RWM645OP+ljFWaOnhObcJ5XZJo4hsfkmvYHnbjkpC+gLM9Q7PU
x0bT8NNlczeNB9Z+PiT1MOysxYQBSsUOPFtNbBSmNrZ/DwBKyBSF6qp7DUt5ypcPmkmDPGIAN4rX
IQUWWtrVpCEGyLOJkdYgFYwTMlnftE/HLLrOFbU3eTnKMxoOTYZCj2ZJ3sRCcG1aWbqAoZIU1siu
kS1E6ozmvdLnDG4v1cT4F9iyowl/hMfiHVLsg032MzgVeJ1XqS+dVIFADzoRqHncjTx3nybeYE2P
vZ0s9Ask82nRGMdUC45JawjVTmfdO93dWW2RXJm5p+z9pyTNtkqtuYSvpoFzbEIDxuqJ0zxpk/M5
dTG62b/CV6M4w+dILForomAKpe/wLWcDrJOHkOpyyqY0EUpddoysL7EXIUKPldRHd32MG/PU5psW
LZwAeVlBCIAQy/QgCXxg2rjup6sb5pqzs5pzMZGuCapi49p7uTIfhQ11A6eHJyjgHLE12VzsZH8I
vnY3kWhHYjCIaPx4E7HFMG0kq9+oU7YNuAEqZvvi22pyBP8egWxG7vq7/qp76zpBToP5a2H0g9e/
o+fd6iq0Et0Pn0/l0iUStMtxi4wvxmljIAV0NQmT8D1mzHPcYn3hEi9DwKtVPZ66SlqrXIpMMuzP
xkYRK8U56/yKOcOd7+0u7VLJAz8zQ/pdRXr9WZUQdknlRYMtNP9P7owzAugSJiUJH0SFI5zFOfod
jvxlwVtkFBQV+RjA2jFsTqmCugpEe06JrnZ11F7VGjN+K3IVJaaEkjz4ADN621BmCtNSOAn9cFbD
qOCn2ECx0nzzJ2H/6iwxDkE9TuAMtVTkhkNhF8X6wsJlBdyY3FXP78HF6dwFcXB2Rz9xuvEpQ551
GpQvvZdwHGoKxkSyKk52NJaQ2gZovSQ+g1oo+FbpNC3oIgNyGux1gBPmA/A4q92KO7Vx0h4N5SCd
kbbrmFt5plyD3oa1lHb0kqyD7heskjeQb6nGXMEp/geAO0FzEXIEWSwvBCWVFMdMkTJjZnFAXUBJ
t8BVRsTo36t8MLan2O+cb3JEsxjExkgHUiXHLW3IxreVb1RWmF9EA8u7K6AwaIyFr3txCtP9JM0+
BtWjiWPuBqAS4gzyCmMOqoGvjrtijJ6fjM1upf7zDEqyi3IgfkN25qVFv3pt9OXJs+HEPK9UvLRq
k8zepmm9dkUNcNHKD+YbzKzOZxu3ENcKi5snLUgRf2LrV7Iod2xs6wB6xtt+5Y2Tq5sase8IXXmZ
kIDKqHMOHwchcGH+jJY+amduZ2RyEMPe5Sq/ZMbyAAs+DLGIqGCVdULgHyVR3J3NOqWfGmlm8Eb/
WUPV/+74p0Re0nLg+v/YAfpaev1DXCnyBvVaLPVYVZFCWLyoa+KiI7BO+mMndwWME7acAobVYiJ9
9TJIdvooz71Etdj9q6DXvwvYs6ah1O2V/kihxuLJzvOVxATC/+7KTe3v5rBdfp3JwdeAwxN8qowt
2vE22tb7hNScp3D2iowAfE530GXZhByFX4r5KSmEe98+5oYKKm6KydB3tjWR51Hl6x6TDR4+ckPM
V7Mn7J/K2at1UOjjPIQxkwsyLQMvAx+drjgd0bSrCkWLIp6rQDmdGTtIwcwy2SS/96AUM9UziOL6
dWK4pdwH5kg39PR3zuIJi46NmG8wN0GGmoxrdDZCqbbNALhHB3nNfIZYndN4D08WE/2U8KH6u+e8
54fV2tnDWsRjnCx5pciJUY2NotxH8uYLfqjnzGotPq5gx1JKGuToz/6lLmXs+ahP/3qSBslF60gp
z79YYR1tCFyGmEAJZ7dXyFULswr0LMjAGaT3eTRLRJEzy4KlqdYw2FvGax82ZR0Cpa26RHJ7kMFO
83AgQ1lSRnArdjZ/w30m0rgz9DiUKxTA5yuJYuyKIQgRQGBuj4duD5ZPVAFDTvq7NJoxDTaWbuN5
8NFU8JR7hUtoJjDocZDF6y57Lluj5RXWn2pqo5xBZs1fMIai8ZQJ3EnW0CFbJongCZbdPryRUuZz
mg1umC+dLTfvAsp5htU/YToG7GqLERbWK3M6twc0SknsEV3x1C8zm2CgwtfUJKCWzAxQl/ogIoJI
fG9jgSTup7NSPZLc14Xj6/4oHdQ2gpB+HWRxi9eH7Hz9Sk2fX6wHspVDv2L4MR44UcP3iSy8tjJw
h8Y6hqoZHSmupWeslT7NpPjljJuV9hFthvKEC9uCe7Smfc3V6m5seCc9JPgsYRsy6AdFBdY2URL9
wj1eD0wWK+6X+RfTbjxXHDONhicCDAkGafzaUw72RnD5Gn5VUDF2JwUpf67Z/sUPHlqfwOcZS3VA
aGMwN01w/TdrQRcFC2QmJk9uy8XPOVFwJDuXnBmrgMmFos776fVS+nPnQkI2XIgUcv+SGC9ieVuE
3bKk+oGCcYXDBhJUBajjReGUitI26S1cVSLFL+2qElH+EaWx7OtIgK+ibRsaF/iDWwyh71vMuxmt
wc3RuEGsLod6N5XYGC6N5SrLPgLf5xoBWAgYZldpFd98w/KNQpw4ebMIdg7O2Uf7Kwo2BvctBpJ4
bgvFydMa758oAMEMexjQ3f4RzwdHcBhy0nk6vyTrd6sCVfN6QoyFJFdn1dLAAy4sKP87O98K3dQj
iBNZa6CxI1X4Dxg6ywKt0OuFgPfpB9QtiFaS2nWcHc+o65WBYMDljCYsEU9LEzZC/l6DLvgsyKx4
JVtqbmRC0UohnbG+VpP5SzGUqRUpfKZAmdnpWNxGno1VetNnXiEhKTz7ZoPtyuGBucklXj3jlBzS
52ycjmzc9hkp/4u8znAzdJxjds61XffN9JI7KN707D0rKAQ6Sn00xD37QNW29eBwwVOj5+3qGFr9
2Xlsu5t1gpbivYNe19ZH1yhCXL6pa6PagKuQWBpurEgZxPFDE891WUCW1Q/VWRqj/C+v+YromRSp
KvratqXQatkQRWF5FqhJIK6P0rvEQNFjtZE60YRWtj/pEuhNUa2URHNR5vfNY1unOFL+qULfhebC
ldyyP/s9eXkybTGkKANJs6MV8UMcHGxUl/SwQ20gOTpb9cq4VzUMgwsqrz9wMjKVHlbAz+WckDXt
C7cEXXXbTGHl9HT+NOv6edIj+vRhwy+7s7E24VetLXmOOypxT55LQfR3vl59JWfVbUVNqQBsZoq2
3Qe30DBjDRNKadJo8KiWKYNidxbhGI/a+TBbQ2IIUsCXbANIDuBLDRI6NoKF0w59jaudXCd16b6b
TE2d1OdyiitHYdkL5swzZnXGgUxuVDA1gyrKcXnHgovIMzHWK23Acmqyxegtsw8k+8jjn/4eXLVT
ZzKpSOTSSFaK/rGHEr2X/lgh1XvL9WIYEEFopfS5gRfHGQl4Xfp+hHkoiwF62y7pjSciLutcww0w
oqtrCQq3EBx/ONNFVBxp8WPGxObVAHiserbB/CPpaAr6NjPL4ITnnlsZHfe8jxLlMz4rfxdU+2wJ
rF5r0BTBKmFWHDWlr+07AWG/VKsSeQ0Yz20d9Ip44ZVLqU2j5y1YmyWm30UJWYSCA+U5LD/GIWib
rA851n9i2+hWs9U20gVAE0vKFU7Bl0gPD5eVt+xAcSWSkxGGDvySk2ZL0MYBVGziFP6RX+4ilf5f
oCB54aO7RChJDQULOEDwu1eNo0cHSNqNBekTSQIrCGnvhZcoKy3JMUmEnnb0rewu7IEleFYqIiPO
545Qg+8S9FoostS7iFgJtUSN0Np0l6gulWg281Z1+kuFyFPRQHJSqI6VaMdHUUZFCnftL/Paizan
QJeVxUOJoffS/OBgI8r81llWSriXSqH5FoFEmBxJHpIgX54Elpug4SBrcoJsFSz7uEXUIMxygsrp
DYncXcL7jr8N6SL8JN7KvDyQpyQD7OwsP/Nld1/8ZhbIWP6VoI+Gj6GaH//voVfv0QFGcCWp4mCv
VTuoDKK+UHqaOTa+jBuahtwofnf5RjFI2W/nO0J1BD7ueAMFXvZMAAhH81Xetk7vB/+S7ORnUfgb
wdD+oByl8JJWn1oiJrXAQEXtpF9m7A3RVHm3+PV+aB7+45v888LK6zP+zk4H2lMtNue+D3YSQ+uP
UQXi1TjWD/XBlyP8xT4a6y0PjXt9QBNUVf4r2rxYqCtQA7x7gsnrrzx5RutYD8jAOpgT+0uU54ck
70DqS1BkzkVeDu2byAH396TRWfHBo2dHxudGXXBqy+ZWmCIbND3robYuY66BDPE/9r1bXYryRCwq
7GqDOwQfhMMJt9uyrms1ZQEyA4BjuptTsj3GynQHUZbUcaM5d1fAveRGweRJ6rZYT8ZVzXFPjkDy
rhfQ6nSG76QU9Z47ReEhkf7PGRQRxcaY230HwWujwCV8dcWKovzWuM6WtF7LRh70qUKVPapY4mKw
vpAk9rZKjYciZzadzbr4lu0jaUklJSG2ym+P9vZnpkLmsapsA99udjEAW0Sy6ljSow938A8rUJNO
e+TZyswD+1sRagpVfpYiuZt1VGMggZMJech1VNeAd5MeMANHyPymE8FZl0u0lBKs1KE4HYm2oVFk
N56TjZ4kwiLRUYmD6RvTb3toWH6xLmE9JvrXfRbUXj5uauPYjqZls39UplH1J6ZWcs+l4QkEBa1F
LUxVB2Km4qbqKgx4VkivWXtsqSsOXH0KN4K5nZUhzd49QNZ021Wy5bjpaz8TXxaeCoWODMaHs4dd
wiJy4HGyATbLgnxC2Crn31dl9gQ2N2VejY8OXr1KMT5QHyhS5zuaOOPr8dqMgy/XT1xOUADEqPI9
nmZlOHRtlnhadTkVslb5Zpe9QnQx4XT8jD0pGTwyiFTI6xv09T7GJHih6ZQqAFOECz74ZH3Zdgyd
43uyw3rVUbo0gGrw6bY+7JBR5Qyt9cfFtI1JChgoh43J73GB1RCIo0VxCE1SK/U/8mSgYaRyA9sY
QWn5Vq+EHIJ7GpCqs2t9/+pMpUbSAWcf41e0kUJ/NlG4gvHoHfoB5h65K7BkGUPO2qD/MX/PsITd
JtXL5BbuWimT6KnNd/B5zgkdC7sgaa0MPO1MapAFK5F9DZxl0DS792bEg3o9RQvwyJy4L1vJJvYd
yRuLB5zAmW+1QUE/cYPoaA0Wx3HFOyhy79KeHWoE7gVN4DVY9c+T6Oy1JRqmi0CrsHBSyLhov0BE
sOxUvK34ykWhEhiA0UgFWxy+KS65btcugDe0+WTQFd8YUItFeCbZ5lzc9Ge2Ui/bxoV5uze5Lcle
mY7FDccqt2gBJo8UVG8we5ceOJqx4n+PQPPraAza5nATuG7FWHml9Q2q03D/Bhi+HjUWGOTcIGpe
LnzvbHMyWg0HpELRL7ylpW3cKh3fOWuE/0jmHWA7M94BhF+4a6GOH2u6HeohVuZLjzSK2ErEOmil
cDCy5xhoLulxvIBFo6eTlDKBw2a3TRRCUmdJL93vLyNT2wkHJxL+r5NV419P8lHgIDCLWq/+lQR8
fDmWI1pIQNyjWgWh8BiZkyPhMt2Siv4FzFXxU27Q3gFwHQOajYqQcdTK1YsQDcY3sD1qSLMMMDqA
595yzinQuclQBz0WK3LYDVFbNbJZbln2Anb1v90YVPQAsYsB3IapjHxFtNADJLcpDf4n0bd6pJLf
3ImiLClb90NxWJTFyjklMhPSNDExtWrH0CtrOuYTEJJWDmfd3aZAFEd615tTuc91/8nV3rU0wUtH
ygRes0qNK/M9dufxuaTCJw3tGpSD7Lm23zwsPtAckArS8EqhmjqOzr6dxM7NhGq8cKDgc9Fs8+tq
AclYT81bFtgQOcFpxGYlVsDw182PcZT1N5FFWqZ7ex7JB3Wc4Q59SB/XtOgVMNmqgT7L4hZvGlCg
t5gMS8Wi6Kr6c01BmOS3bkoex3sut8LVR71XQ5vmr1m2LHu5lhjKkjwSd/Q1yN702boysX5b/nta
sdpRZbHjPA3X5Pf7Dm+nWPbnudRG9Lj+cldq2yyBVM4U0i9VUPI+9qNgzN1VJ0KIv1/PoQRNR6gw
hIG7qkiFrKP//vc0BaL8JkzmPG5AWa0eM25oeXsBBRLBC/I5XMu8HW0plmGgMtl893FIS7w5UL7V
OWlrf9Zd2L1m2oWiOlZUJpG5JzQeXg7QYBzREB0i4TpvglTU/D7sZl4G/307t1HJQLO9bZqx1L3Z
wWm3YRQt+ZhzeawwXXEUp5xS2PlUPYpYyBbcFp0IdJSAc3H7XBxVZBrvSRXzMFe3PovibAAJ99cp
KcoxpJOY0vC44uXmI1PO8DuL8UPzii3nYiwNIOlsMS4kN6Ywvnts9RMbhaWprbRmcYcV+iYwi725
Yf9Bii7/Qly3wNzR+NKmAmsFZRrYkO14PRjfAqutfRzMN1Hn6kvnVP3EPXw+ouY44zayzc4iDZMp
yjHWtNavWOjpGQy2fZnvms+Y8M9kdPZ/q/rwYTbUzJ6K0P3Dy+jI1A8pLWmMLYAoGZJdt4OnzgUc
+G8mt0ixvO/JLcUghHM4JMWWszFYpmmnglOhUNAvEOGl0/bse/ER+zVskULFk2L9wPcLPFbdp1mW
3jtv/dT1nsxuGARScUZ5+De57WzI0anMcSI33Z7KkNvnZBPuJJg9LBMKsD7T8ZKqGCpWqKDdQzhL
URy8+3v6OcadnexDfGZVkuSnqett8hZadT//Y3L/FPUmMGhzznDb1GBLZUI+wrrzVJpYEGgvstB1
jBNfqSU8Nww1hO9E0stBjgYrtnV2AAY7Q/xhlo7YKkKVcJPb85uoA9wZd+ut2kghfCOxIoiySNmf
Iect8Zz8iohy8MLxJxxF81W4MQoOlZWhhCjpUGuhQQ2PXTFEejqGMtausmRs4mjRcwUWJ29L/Hdm
rpJxuhWe8eNSGhI2XF5kK0z5kcbGF4JB4lQYZ3pP49aF0dxa+ME24wkutpX4FjyCkw3QVWu791aZ
fgkZ5zD8a8SEa4bmyMp7VYgEp4B2ql+RBABCNcJqUGNkEiv832TXcVefNPzmcUCZ+WV+zW9fluF/
7TvE1SYzTxjSvlmPhb6mADg55k6ysBxr7xTbjW+y69LF7VOvt2RnspJ1gfaH99KBeilagzCEQWPi
XpGBqw0BE9j73AKEeeanfJWFQrkJu2GbWZ8QbGeJNupUdJ0Zpzwh2nbltuhydaZUY0zVRvOxyxbP
d5SC9gB0yPvpWxW2C3/1o9w398mVJX/odkjwv+OpZAJWcj4+cxydcZ3kBVvf2LKKLeW9bF8RW+nW
J2TaAG/QaMZhJgTS1cO9A2g5mvSfcLRzF+0EZOr401qSr6zONE8A07ufAGlA9NUPmDnXHGRjQ2RX
j+DIvM6skEvwS5N0rh4dR600CsEnyTOrpxL9hSOOFjpHzLYKrsdePOLJN6XU0jzWZ2hQvqHPYSor
Mdpd2lTsAi/lOKfilUNQlOr66qzMb5wh/O+N9qfjrfwIBIhxN3CX4ShobpWYq2+jsxTF0OQ1YVF+
gj0u79W6PO+ZnorMZUkSqpc/SKSCUnvXR+Hs95DxiOMeOw+4cSW5IT4JtyR1SpesRJQmi3kUyvfC
miYxUwS2WBtEdnfbcOm7lIhAltgSbY66hHmXqaz8jZBYWe3jUezX2pIu9drcFYwEDEGxi4UWYxH2
DSNC2sI0c9cdTLgE+nUaAE66F8bUy6ZzB/HQY2sEYxHRiqn+hhKzlOKH0rLBPTeR8ueUxazB2iZf
szlxDphYLhBi16WwppvXwdspcFC1xuit00G96wUMrFtA1liXAoOYPlJGBjyo1EsdD9K85PAXA5wH
8tTZ46par7mjvZx5MQg3d/fZY2PFC4R956+1pZE0e+q8DKOLLtn0jCQj9t/hRx2mp6eveuiGUHlU
1heLAn7w9O1FHXaDm5RYMTNsXUgHrslm5EDmIaTvIqEu9w7tZKjz9yNkiKz6cG02ykCL1bjGprjS
Q0CwYtYSY/cNTPivsIzve3JZE3iW/E0u2f4W+1nIlmIsXW263RqTT32q1P6C+sy0s2xFss902h9G
20sThR4doyftcqDJjVO1DmFGS56mMXg3P8U+DE9Q+0BuTsuxlnssZ0YSQnk0AThb6OWLGMsf5T4Z
Bv5r7w51tQGOFtVX2imOIO6rO2rBbKAaXGUwnBFZc/23k1B3W5hYmSQHnX3d3v4EI1jHS1JhXaYz
2D3Xsuwbug0zRPEa3qNVvdnM8AEHgI0ze54CEaDzF5cOfttyAoFfryfQypN5/qSiwpjyd6UZRfeO
vZdzMeIvws0M40pNUHkWq9gKunMprSry3fIP5FkB8Q0cfVwn7eSrF08AzWJiG1T0yw1oZ921P/CN
AItX2hPOMgusleS8miadNfPL836NFffr2IgH/3Fy2WvfogzdOXm1nULhTIUaJKROLsuoHDjFtRi5
zk9hw6qnNgyoQHYAPCsNl0x726t/GtLlYXcyMG8yBbjY0VxjOR1y/d4oTnYuW2Db/WMofZbCWwu0
SlEs7c8Xzrl2J8KooyOWz0LlQ9tIg2D/mzR61rZlhUEv1UX/OTa6NItzKk8XNAOgE0U1YrKjTloo
lPru9xX4mhQzGQZz5/jqMqDT3Ye3QjOTSrCDk6plYZuRTw+j5PB9x91xCW22lev4W8Hic40xuGaL
fD+njy49CkQd6xe0hJCU4RH62vqu5TfiymJoi48m0UgJPiALhw1P+tmIn39VSfJZee6agPBzNU2x
93qgt2qFaA8FLSQtf+g9FVGrOs5S1Cwd/ZtVPnLR1U3SRSXbr4WW+9dlBllP9yOndxsXaP6eIDkP
QAkaZer5/IroFQPDPcdgNmi4W2+cRpWBbiaeFiuLW57NihanJTzGpatkTFohBueDPMEqJxEbgHEk
LYo8eCbRjhwrvbXLVqAZQXlqc3tONUTPU+U6XfH/8nvUgNGr9ZCrBRVy1mpaeIq2NXDGClQ2yZSG
9NywIaWVw31KkrU2PPN4D/i/Uew7KcBPJgZNHq8mBTKRTDeAalDoqfmt74H1pIyuo5lsAW7584SK
jJtudaVOB7WP3eIf/B7Krpx2pa6QFbQuMIxbsR4ivkDPBEQSYMbDz9ZK/8vpved+ZNWVgNDy5h/u
nz9KGYDoohIJnEmK3S8qfQgm2sk3853lPsCuTOheWAVI1g4hnEuZzT9GQ3ZDEuLLwHqkSjrY0fp8
KD6mVwpoTUUoYzQZ8X247Mz6KY0yLWYcXAnUidkhTlcn3O0gSzfA8XLbAMcZVdBdymmUQn+ZeP6D
k4O2pZABSKrUTd77i2FuR1ETzb68DSC8P7qxiXRP7l8KBdL3uhFze4t0U20mc0BrZJlGvuwNKqXX
LSMwd70JkEI71DRcqEQ+dACndIy0MSfYxMQPGcsEC+P1VTBmKLSA5Yt/Ws0WEYKxrjZOBho003JV
yfjb6Wr66wmNop6I8B/rXkfZd93f/YgzjV4K+iZ2pCsChll3T5ndwN4K2vuUuQIMem5ee2fu0Gv6
Pq6flMGMUV5qtGSfRALczZbRqvSn4AFCrXhdqz1N0Dv7ioZiO6YwleX5AIOJaExxRmivLEzbLeu7
FD1cbjt+b4WzkTYAgINCwJeOLBz0aUk24cgZS49Hwscn16RHCmTlnuF35g4z9yFLDrTUN9GW5aR1
8Any855O/3CginzUaryodddziMMY5n2AGc2t9TOHdecl0paKti/gBc4snVtzQh9Bp4mx0cW2lCpv
9qQBbB0fAO1dmHZqXOeiPWRHFJdTM0dt3+ba0ypriXWUsyACgIMQ5TFKq4CUp8fa9wRfZrlNdb0Z
tvZ1jV3cklf7LHxiZjZf9nbqj27DGo71odD1XPWgPFnlHUVMUkzdhlmuo7WcbsP2oegmrSo/wyxu
VR9LbxPRkza1IFsxO1lPSy2nVLpbiGMfuTKzgehJfXg3gbfXliGgDXzQSKNNhZG+SlIeWzbMBsuE
6rYdeKrVUJO1YNWenxb3BPdYkGpuYsjF4wYnKW8AWMo6fzI/UJUz3RKylbvyeLiZtic1iEfPu6pq
v9vIhcxT+UCcsU5fSMx2fJyz6SA9VMA3g9hBmqxoUJjBA2WTt4WeiGKYlCBr2eEcKclzgGMmaLY4
S1Vu+2rhZYDZvgw6OaUm0eXxVF/ZBX6or1ntFWFD4A5KMvTvlzXxxi2XgWbSv5xQZua63j2mJXc5
ZPKVlDhyPIZK8p8NJOAwrPzCSBQ7fX+hKyLe+lG2vS0h7SkI9VWX52KINihcdj9VJgIi6mb8RzN0
4uL5ib6UdbVvdG/GgsUO9LTGE+mk0A19/NnQwJL+o2p3Od++/bwjI65XBpd2+W7K27HH/q/sqQJE
0u2l7YibRqG+FeC9B+2nxkYdyvYXhlf9iblMQn1W6MOZYVRQeTGzNOdJIzpzi80WF9eqljG7D9vP
aB3kneINSg91Y2rkeJ+A4U06FG3Z0qZ98QW0MTleTG9En4igarrF20Cfez4vvUvpIO1KYo3zH3YN
XZGVKP/wvDe64JpL0bZO3Ceg5r+7hzVtPFEFZMkDVO4snYHEmYZxejI5xpeycjKVQmqprK/l29cy
ZTMqgqVifyEim+b1R+rm24tpO9oZtAWM0woxhONc6/hc55fCPMez/HfsNtNVEQekH1gHPasIWtJP
Hs+hoX8y21O3AEZD/9XK6K+BxBaVAZdoggmGUPd/dGUyUVbqT/fXvTWRUwmJFA9CoNShrIn/BH6n
0qrvKsFmg8ku8P5QDG+qajyAXo/90tDnL6653u1pib5nVdo5V6FOirv6/qafXu90267K6S8OixrV
IwWA18Nv80s0jIPutLwyBnYpeGWO243Z+76WV647liPri9JENWc0QBnkH8LqQDg5EZ/+YfuNphJ5
wl+Dqcqacsz8CkEq7YGqt+w0hAKcHeKrpri9cp/NTfUZjPfBl3wz5jI/N8QDVODarg6OLod+OuXX
rwr/98ounOZDefyC7XbPMvJE8qGCdz0Thj+vw5aeRD3j5QTZDeYhgyXyP0nLO1AdgsE+irqOA1h0
WqW4rHZKnEMRGCZt6HonYoPTRnitOKNDJzowIQxoahXOH6qtXi7zVWPJI7Ri/PBOp6zilL9wc41v
FLVSCcNSQ4izuWGAe7RluOVT4nLLuBkv46jdszry5oTZwVAxtFtlYT5he1tdft52bMyud0Q19cL4
PKWrbeDhld0cEJ2LalThifQiIlcY2REepQlwWm26ZzWRuc7PV1x1Ekuv9HkpjW6ESfvAMIqwbf9Y
4b4eVRfBHifWROutpFgfMZTQ8/POhmeAtBHcF+YMX0FFZJ1ORnInK3LwDmSQaeH4WaOexXGBhsYE
0xw+mz4XIZjTYehz8Z1JVBhGBpcp5EUNdN7O8kbT0xdegOc8XwZU+kGi5zA2onZ/RgKXfAgDhgqt
1wGlol7im6DRH0DmiFs7NBlBYgOj0qVacXoZ71NdMZSF4T5pEcGs40D+EaK8FlZzi/yexi/+8GXP
CtmCTxXjcYfSlSBL6jZ1rS2oamWP0eWPj746MaOpK0mntCxoaHC04alRLJZieslj136kNBu1d608
izy/8Dgiiy0o3Hi49anfp+yffvW/qv2Oawvs1llyerdHM88f8Bx2rMX34ogwtKW+TOxgt3C6AE4V
zigIsfY9hW+tJ4bvjKrchVCeDxZGkh/HUbgxN/TsL07JDYMCgeCjtHQGIvoMRtI0TXkT1Ax3xZSi
Ks0kZmGD3DCjNCGoQT6FhqKBai7eoIoD94Tb5R3yjOhn/si7vz0Hs8bG6k7H/0hoOH/KoW4N4FUF
3WlWL1VzUR4FBfqyrlF50h6JY3I57gnwxwfXj67C7cU1p5TRaJ1WA6+ap8dz25zt+UizzFnLo+o5
fbnu6gxSMeY95EU3Rt44ccRAzbckL0PpCxLO0Fi7vc+TVOPWyUvWfeDyyNfcm8YNDA0+t7lE9IuJ
fES5b8JTYw5M+L8PpSqVRDqPptuQ8aDPRAq+Giy+SRcGv25ev40+Jg9/ZuC4+2mdRP1qD+KWu4hm
pUj1V3PPibMaz/mynyzarVOtJPJk05aJjR/WLoOj0ccmexdmvEqrLmVCse57npI9odAVmSdScINH
2miN9XlXl+++be+CCNQv3e89RySC2i6WPb3aeoyJW909psiQHUPq7SaHsU1rJiCO1y++SgomAW3c
z0Cq4AW2WQIsenk3nYfWCH5WavBkbjJC+1feYPDP6JIrcZUs7BTmu08NcfODkSvdzCuBG24RbMnO
VEcT7BhyFhIJ/nlw19Ne0Pd0UDwvvy7HIBhRBKUcieEl6wMiwXBKkAE1S6SRBXjhXDzbCPx8axCl
A611+7wxoVoHmJXO6nJ08nL5N8Suy2/Yi6YFC8QSYmvPqAOyE9NGOVfl/6ANcACiaI/9ZXrE7r4G
NqqicHMt3Q0EasK1v/N7NU/itw3Soi8rEoph6WNpFTZTsV1Weh6KclspooPQHTcuXT0PfxdYmLdD
YpKlC/BWlVj8Kazw3BvyGGswxXrmJ1HW/QhQznXN+xqsd3CGaJpUOZHk5CWUQtV+m54QRHOGu1sI
3ipwaj1IAlD4i3/CK6wX9FihtWzVVzsDe2bBtU19UGjW9+CEhfSpGml2sHs3e1wyKHbW8X/wrCGL
DxEVBqLO+nk82PRHh+T3du73ss9n5sHJpqudUxpm0LER4/fMh5+BtvsX6JQzoHW4YfdHcD9Hiabk
u/8QyNN9mMgSKgVn2kBi1pkw6te/j0W82VXNwO98xu7spNwe4VTiwDj6A/REV7rvw1ZV7hDV6OUo
maI98DkJKzZ8pwJjKRnTslI4KWwrCzte6K+G/oHNEBhTzlZ8Wkg5HII0hluMl+lZMLRcs2BI8Mxl
iRlgPiema1S/W1kU5PTL5J6zu9EvWRnzIeV1dTtMQMGZ4FKhvPAn0QcVIszl3S/wEKk0WoXOfg1c
skwUG5Kr93wObE7Jha48NWGAawvcSIceTxjdMGgE1ObnCm+u+ao4RG1dDtUnEToXUWnqy5uXV8ZH
ZnL3UBfMPSHSqC3ZFawP/VGIpB3rvcGqM+zMHAW1CsWoo4x9yr3jb7/TiGsAlcpboPHEwALdO/Hy
csz/9ABpmowJqzbw/a+hJ9L9A8s6V6n/ygq4QVd5VYg2K1Rd5e9EWlGGerSIcVas1g68MTLoHX3u
UNevw1caGTlFUATaTxzmQQY3rBk6pU3YPEJyoOGgb+qRQfBlnANjBYdfYy7Lq6WWLII/D8LkujJh
DjtlUwfzFYCRAh02fFvb7bmP+S4NUz6Dfqp/lC8vXzVOXhLl7gxicVIaKhsrsiRZE3y4OcdT9DBt
AQM8qMT6bCD4HANfiALvs2STpJaUzvGm1MTNxcI6QHG1KFh11FU68/YS4U3ocB7MjlslpiwCJHxO
SDFpQf9dGubSSS9HEwvuKGQq5TJW4eolbMRoIkw1DI5TcmPgKA4e4HupSwEyUDOFv+I5Wnpmb+6S
MVffypagC50rjCtEsktpmS9nRcr292FabUIzteKDaYF4kEAN39zbCex2yCNDe4j1ZLv7308VctYA
ROd4njSR5pIdcN4vixdN6m4oSxaZiLXCR9EQ6wMBfMeMYYAB/CdgCDcc2zR7ooEdNlqFr0tZ8S3W
S6VhsarptBBXnlXnJthEmvcyxlFfRi+GJGSPefWdT7FHMOgqMrcSJL/QjDX2mMNjVvYg/CCOG6mK
BbOD0Vvfjdee2nvQqI5xaaOuc/Iu7x1kcDIw1lhttf+xVzgbYYl/d35ekrmckxBWjauh6NcaDG/k
Fc+QNZaocIKzF9PGp0MebDB9pAeWYGY+06O6FyfK8/QABu0nWNnL04NmnWxy/eiKrK1tkoyIp4Cm
cn+KeGDlonCEqRNljax2q4HjrPOqVEdHuXWKlPBC18JOToD+QCA9hzQNry3/bAL4V1wWH5i5VR77
yMmMrkIjaz4ZtQ6bhktf5v0005mh+SNtTLZA3kAdfq7q5N+wI7JbfRg7AKA1JPAO2Tq7s8QuOF8M
l65RAegrvELfwPr2aDtAyC1Kf27BvlYe3LPvNxRN2gR1eqRd6NS06Ds2hin+d+F/3iL9ZAr7Wkdw
YGSVzyz86ItRg74l+sKykYpqIjU5Z5Qem/2GQm+jdJrhjjaOOAmtmWlzK4KPmCIabSFb15IBufi1
4pqAxhZxcfl5cghrodOFfxY4P+xPOX21QQowOskC/0QopkFzsmeYOms1Es17EvOWkRGHxcGD8d7p
9SBStm6gX1Li/7tKAdKS+hYApRWzlPg9inPQlhvQHYf+WbJu4EsOH9l6iwVfgONBNmt3EKfQL1F8
QFprd0Ca+9amVjK83+pW1p29tWdIdv8EVHqzKMFD1zinGm2nnf/4J8nxT/1wl2qIGp2oau0WDGX7
wLhVNCR4mCQcvS6oOJRErZMNXJCEBH/LT82kBu6Gm5EBn97d6s010G2cUh9n2qv1QAMozMHqiYAH
qhdMTSkCbgUttySY36egnyFn5/nd6oDOnbcMrZ79j1A4y1K5JHjy2WMAXq+7D971ayQtek9LGzLV
nFG7e7ujvDF/M+8zvVs1Q6QTlsRwGloBAJJW6MUm0my3IeODPk8HI2TL2IQfsXsvAQOKleZ/4NO3
ZwAGygTkbVwkcFLu3eAbri5upNfoRN8BZUies+2c+63RY61I8UhmTM+rPbMsUZ7sOVeS8W1xis2g
y1o+zBEZuSGvT2fHc9V6mhAwKC13EV12KlYNnWODFZ0E+wgwFt6x6F4CBuc5eBx39KSW7YR3fZ0v
5eZNIqcwrOTmnMPvOzQ2YkKYrALOJjqZERJF/QUTxhopsaFKqHv+m2TMFkMGb2hJNQGIkkrfC9SF
yjlvX/BUZB6YQJ/46ejvLHxPCJZELD+HjvHGDvyoTgcTrZTUAyMBjh9fd+ttqrm+SESfAR4UxPAb
ToZJj8BeCrLaarVEbJAAzSlr1c0xMn1oXMYkWmjy11tZcMzgdZK3MLByIUg+ihfxBAxdfn7YvdaL
UWBbm1JrqxXMIsd84Fbgb9AxwVbCh+opTEhztuBdnpP2EgFHA5L7A1eTlcTF/o6zCjLex9de5HGl
Ux7in/ixz47/m3tehDxUXwzagrVkbzJ93CXnI0rboZsbfyioZnDDwzx7cdYii2QOjVlDaC043M8+
RPvxSAUqr1fyAlVJuSmLwU3Y/MERriaGORzJf92LCKLU2BXR5u1q2syB7sXZtSVOv0uHEp98UEw5
vv8fZs32W3BBGPfMz+ETzIxy/Na2drV9rIhJk4VgXHtP8rtD6gw4AGhZzuXMySqJXLawnsTz3zSS
YT3TLcciSUToYbYPskc97n+HBWzZx9b8jTp6L41arAnBSGL0XX+ePA3ACncn92mLSrV0kvCaqwUW
i2bkHiQBTjPY2J7MCWOwl1fEvnZsXtAsYTSEaCM22ZJNUoBZHALsITvNKfZMkFe4Q2VIFd4T1pwJ
tE+geHFGuZ1Wl/I3TLM+IsgvfNQ8alvUkux0AC3aws72k01E/AR5LtJis9bQZ9l9fiI/JmTh34BC
z03YBNg+TFskMh1eBqRke01Zc89RX467rrdbzY/5IPz8O3YCs281jTU264iRMUZAqHGNgZze+spp
T1vEFCbUBjhmlx0BNnd/sXZyrQ+mZUY/QmKPXyuFtfqOADNpOKr1yApIuvroVNVOU9s+8COivdnF
6ZuLqyctNG3oxCDc3I9hHaEGlvHprJOctNAuErBs14+R4Vw+PsCuQg+owOzor05VudmfHaaKy3Ad
8rYEORXcwQhUr9vOGiPGqlFoohh5xL1eHN6WAyZyCOXjCFV69/8AoPsx4LAdmv29ZjOab4/dS979
a8kcQtN8E6eCcQ5WAYtU5ywAJEVOtflYksZ57kUVxOognjpp39/31/UdQpx7STTId4HnHeurC2H2
DCySP30F1Vw9zQc5c9bqQQh5L+uE/XDLN1qZn4hCIdE6umURO3UxowiffsqV37/HZcFsBY/Nf+AH
/du0kddDs2/Z2lVh7Na9FnK4uX1aIRiTXcn24k3x+s8JrB8jFo+VBwmTSTQt3/VVjMvfZQ8Et+M/
4DFJfqnIyoyxNsnc0SOaN1urwegAAmrMOYLOhXG57MVw/Jx7SJapnLTk/RtiWuGL+/tqIjTS1nRU
JJR1xG8FqSoHJM27qdnFgIZQYR2XjnMFB3pvZdN3ygVWTGn8ggyHcKk0Ci2iOmSX/Eco8cFtlQqM
bt7DEHrCuX39FxhR21qcIQqcYRHa66RQS+dNOpsyi7oGclH6nRY5SsSm0kfRPx37cGh61TkWXhRB
g9Ups15Lfxim8rcIjUwDxF0OxKG0DGGzy7I1ude6Lcy1ODL9CQicKs3Ea8VTkf6loh3cIH6vlWgi
`protect end_protected
