--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Q1p53y8C1NvMsO6M1wzN3925RysoganxnlMCKebD9Cal26DcxN3/NFCP4PAEc1uAr2w6L7iehsar
xs48L4rwWU6cjefljZxP7steX9e/Au2RoT3NxuProuOmpefKgeRjJfkgUhA3ZWlvSOgQnlYgWxo/
Ee9jrZ/WEkER2/eTPst/05uccoXcgQJUylUS78lz8Y18RNA72hlyJ8TuSWoGgBcC2yhPER22V9pg
UvcUE5hsQ0SJX7+wQTvopgqLgN6lPgk3loKVMCsszDjg/HKuVM96iqC1JW1NdZLlzwYUPBQkI27g
gppLkd1wrT+OMtV/HJO5ma/oQ4+1FOhwDtSYzA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="49TZWZky+2nu2qDplJPrH8LkAbpBo0TVqkqyv0PVbas="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
EAhe6HwAqy4k6he6HvKPTCI4TER20bAmsnNB1so25XTVc1id4MUNR6bbspZcoIbCxiNQsTyrNm0F
2m3O6J9vNi2ccjgmiXgj1e5PZD29uBjzN4Jwgd71fjM2ZtmK/MLP786O8wQwXuApfEhGbzegUTDK
j8hrylBfywIpiG5KhMktX76V6fKApXo4pHU2l47UdSdfk7DImVZf+tfdN2VbtM9rdsWs2JR9/NDj
s8jeA8OtGIJfSgJiveccYt91TFFe5wQbOkfxBSfpZcRTTqwWGkdsAq6P9J2rd/Rc1UgA+z3QPGFP
ZgntYzGbxA+XO1jM11Qwsgt7Ew17w6AfpMZa0g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="/vvqGf+IwaMtpnIPz61Znw2pUOWOKkSgtdNbQmnVMy8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12336)
`protect data_block
4w9BRObuhQVbPT9+0+wUgt98nIxZLIsi+fuoVHX9dbSEd0V2Lvah6Pzj8vdnYYQqUbgOaXbvCnlc
BGJjUcPeefQ7enfVmLCefdGMJTuSvzjSefCp/WGpNdk0pyXo4YVJ4vos6U5sOoRY04rRG6bakg26
yICEXZg1mXPzD0toMpYHFe3HEpvJCpZxy+Q+Q05AxrPtJVp8wcqzltz6a8bUyMQd5FKM1fYUnO4M
HYrMdLvltEIym2EkkdWxVUyV9LcLBY5b6jCXanCAZNFMFblOLC9GLFVskuR3jeLrQmJi87+FFocG
l/2SsoKnIR6fX+d9TsgqdvpvR1G4hPOE9TJzwIctwBCWTqz5m6ybausXVhTWeni2shhYw+RZPBKZ
n5jKKOEztMAiGAkJK2/B+ptsrqCyIDq1XIj+Hd09RfLI/5CmjSk4XF0MpuVMd+91c+Rx3ufzU7Z2
ndKQ1/sibwB05d5DxLoYpPNmSGZ7JhV7uCZmWG8vVVrX2LN+YYjQsk/3xEmrQYoSe2WWtK8tyvBH
BJjz9ddNnEti6R+DeMVvEhvXjg0kSoKgqGqexLLefc0vN+NiRG6PgzxxpXBlzV7S1C9q0N7Xxapr
NTAUuryab23JEiB+g0KFzrQofeSG8ewRR7/RIdO17Vdg2ro/UvOHnaWyM+nM2UziGnwbWv4voKX8
gilYLsigHUgz4VQmP+YOisTX4KYjOJeBXVM4lSndFHuwmvBzYgUKT6RAz6Gw64iKFCKylnOQB+C8
tDoaoBCZgXYEboi4TDM23LmWLkqJe29pC6Dq53byIbAib7Xl9Z3TvwBtwEjS0LAikAcmxJRQCAa8
BxddIe04pPhSOXHVu+rfCufALbx/Ny5rnduEEzUNdtHCGDX8RvmVI2pIF7gRArA6dbwv1824+Pku
Pa863XtDn2FrExdiwirdOPVwkZHkTgN/adm1Vq7oyKQPoarTD6cowloTLKuTORnfCUzquPy7PFWy
2Lme3JVk/P16+hivXghwjwBsu5DBE/OWJ5c7cAhqXF8GdM57qhhIZIyjUurLAjawvnYSnlU1WfFI
VzFnhzHvCHF96N6kQFwyWQnlwPuwiSmsqtqEfiptl/EtL1v5QBv65d9IHRQYWN++/6Bt4AnM5RdT
kcJIfiJTwEXv6T+iEyRPT4K5BOnozmf0m0r3PSdW9NDEm6XYDa5tno3YQ1lsUI6ZGZiS5pOITdLY
vKUZl/rtT1vf1tWFocXSTV4vfdKAbmleehZqVwRI0MP02WMP2AyirnUC+vOHZTDhlA3A2UngCB3e
3NEyys/hFZVvWzVzxvBvcDjTOKDzZtga8eIfUswPt4u7HgyFzH8S+XVyh7RKx+xHj+ygx30SBdih
k3JRJ/myXIN+wDnCmF/KUt20ExDXcsT0zJseMF0IOAUwoRsj9KLfR57UIOZx6dJM1sU8W7hQORE4
SkFzUeg0UPd9nV3hmzvuPqbaIpLEYB3Y26ys1S1IK1t6QK6EDAPD9Y8bLVWXqEA3wlzFiBsrmPwU
42rNZnxLkeuYqF4ZWJxZU/3//ZQhm7Do3B9xgwloQq97BOUqiDcN5fQR7FHAPUSwmDhYZNIT1gs2
nl9MMWS4EbV+RukWMoK5MfFPzTQvt7FmdJyPWI+skHZszGTTGlcr/NJd338COCkpWRWrmpORne/R
1QDxBj94m3j0TqBAhRF0qTdOZDYUs1PCMNkO+Ko6zMnGHWjkzEgDdUXBGSdFxPP2D3wsL35arsxk
mGfhkKq4x7qq/q2EC4IBg6Sr5n1aTssRhsW1hDZp8Fs6CgguY7xALN/1hWV32nKahG5YLsMOkFH7
Te8Odkplwt7QVkqFdL44RZQG1s4X7F1ISKQHYMKjOUi9NHks7umQc/CU4UcKjfLzBMRwh1+s1zAx
bGeqkaqQ9KhadMoJvfgVbuLDE9y76orVF6ZsLGous8QxQVS9TKrPLwv62myGqsx1XH+dhmAYRIhY
vB6i/xakj2gukHLivExNJnRqMlXybUoblELu1dNLLJ5tqDSzB8e57OQ2gysY9KwfokllDB/5n+UQ
hj3zDCIwY++4t29V1tuSy8L/6e4AxorcZePq0Ksvg7dRrdkkHPshmcOz1sizZV45G5YcS/+jeixn
5Wc96cKIXSgKvb5AxfwS04I1kZKO4+VbTAIbEYppfwdhAuL8qby0+XHT43sRh0KNZTUQjNlCcxE6
ErBIUXjpm9dc8cE+0supK2aV5Y20ix1uDFulQGFW8KiOYwacxAGYf9hLxzgJ0IiyC/zRubclvxaL
DpiyTv/YnsT69IRBG3ENPvVyNC3K8EI+J1cSLJN8BG/+AjVKFD3lccvLeeugPP5bblNxfVg8NVzV
y4x9ahL4R4Vb6CHBRAWXOejiWNia/obCeFUkFXhAeJKUuAoNnkX3sS9jFmHmlOO7ViTPyqcVZD26
dO2sqAzNThvzddkaz+Rcp92vyb1nVAVl4V1xGUcRy9WEM5d1YPZHgj1kkLkZgpKZ5XkZOfm2pa2+
Y+JrDGEJdxdvks2RhdoTYDKu9UPjNQYhL2fW+5pRnVr3+QJuXLg3xKcOiPQlZY6rCFaN023a/Nlw
GaNBuKS5hiHe22Y6s2uDrpIYZow4/LnzpWXZUIzeOnqyeZ+rApb3/isaS+TQWX3+0co/EHc4oNCA
h6uaYXm2b7aFdM4iaX2r/VB4WdGj4iXbLATlPX76DJq96gwHLOYb1vov7yCQEqmVNGlieUogrjMz
znEPCmV676kS9rQjs7l1n5VOkXqDe/3o5HHUjc6PtykXD6aVXfiP1OmkHpzzNIgoP9SABXMelCYV
wRp5Vv0mPC61LzlAKEtTy07hQl/VazCA/OWwV6IlU2Uq+EJ8Zx437iBJH/zBhf2xsAfH/0h9AguW
DRCZYXT5NI5P/G2rBqhLePW/AZVqnNx3qvWM/V3hcfw12OeFDP67e5YEVNQ3u2UxsBQa1REj0PP/
P4H0sCTCSdbvFtaFw9vnP1Oux/sdfzVuYB8Sao1W/9u2wChH2KeborKYvgirTSjBZiQq8npbwu1T
O/Z3X7euv7Czy5C6L9ywdqgb2H1EeDni9hq6haolTwJryskdDBBY/FgiGdOVpXfv1RR0q5Dh75a6
6oN15U0f7jcUUPAxKwfzCRGUZCUrbo3gUQMLpflebsGCPdUip3l01r68W5Qr08lzFFZ+VNUO2A0X
CzHK9r3pvKR4ZQzgPZUHRzj00B1Vn+B4ZHzbn6IsNKy0TefTogEdDVMQY1lg2ILqDj8eC4Mmb6os
Z30AWiOXd6UQuZziCzxQcH67APugbLlrxTxG99OQVrXSGxyew02mBhLiksOjA8j9bETvz0QymApz
aMFRybvY+yDADr80kQcdBJ97rkIddpYe+aE/eZJ0iwfhPo5g1X2RHpxwpZNNK5IHOG3NkJqNzrIm
7SyoDNEPfQO9aNlCarGUvijtyxJfc2I8yQ47BzpGfIr34zCLuGbfTvknA/uT3s+cuU1ocqmme5lq
QAMcQoQBM341/Pp/mHYLpJsfo/i+dzPQ3eNmko9G5xN9AqFF5dV4cHWq7vOTeEubHLgrnObqnNyx
pgj+/x8MFAydC1nOqx/5hpaHgEQWgn83QGrMCNujUUjPZOuX0pKDHJBbfgCYTZ1OGPKy1J6WDixg
swPV7XgFQNELZFChhcKdRKTrop0anZwoBf6Q3ytzJmGg5DvPFAgeKZy3Kzq+ZWG6BJK81gZvQeov
atZxIjAzXw4eWTjtxvu87UQXwsGQfy2Pt8kN+2Al4kZYqUajcc3XY6Qptx2O4cICFK9y4y2yHtDs
dethLaGPvknzHZhP2PZCjdNrwe+KfNDD8mNGzeV8ru9mU0JYEU2hbvkc76hyXLYdztU6aYHsLZeO
n7TkR2J+ZzmlX/eJXeOiovjyXkaVDOGq+418750OOKG2zs+qDTDI1+fUoPf+DNzRSCh22YMGibUn
1ZqZNRAUvg7YYUNX594jUe9OxnNOKQs5e7eENYu+Uki3mHtuCTalanh7v1z4tZIK8rZ48DWQL+Fr
IBnyN3JQgwBDqpS6gkY6ylIIVVHCdtOX/4q24AhdsO1ZAJ3BsDXPEzilMPj8mSvvsXOWI7yrtRO+
5JK1hN1SKqvyGnIJfLstWY4vpZNjjMCLeQUzYGr+Vqun0Ww63lc8XBEaXrI7jIGqnBw13J9s8IJF
FDlIXJmtS9rdLxxKUyuxJkCSQh14rqGXjeZEAlZtIteJLog1SsrfetiP20IamklOR4dhLwwW/6nF
GzaobRn1kSEEIb8PeJIj8a52nQBT4YzobfHvelDWkfR/48ZOO+Jiw1i0ug/FpOA0r7jDLELBV/C7
4K0vp+Vgd/YTdr6SFENoAxxBdLlJdjEagLLr5VZJ0KQGqPfedcUjFR+m5WUj5T82Jg54hrB9FwGO
d/lV5z6rKvmZeju2nF/v1iL3UaLQJ/hisOySzKSSy5UwZvgZWXBiKnOZaUm3A57v5hxu13/kODCG
G1uwVi93yjnjD1NMAqBR9/kGX5R4H6FG8Yarrn3DZx8qGxxVVMYnbkU7T5DdlUSZnkeAQZD4Rm5N
nJ9EZB/+i/jUByngSwG62tpgtuCXI+dLuRKqVHW+QcfMPqAYj4CJetT8Z6oGahPjEi9tjQHtJocg
5LhtKnNZgxAHBB7JQ9asK7ASC9hostemNCIxj6SWt6FRH6lGbqDcvN0hFunJYzN3IfiExA6BOXON
wR8/+rkhgBBZIM6tcu0NEwfSWvOGT4jffOd1zfrBCFfoioJOfIHfzaFEs02aaDOoL07Lzfc/uiRJ
Bj3+baXEJ4R06DL6MDFW5I8OqqMZsagd5UFmqX1kVzdNKm12fItDGFuuQNwy+fEFRL0JLxD+lzbZ
lqFdWQnG3UfumADVt35dSEdzGPRrU/Tw3/KNvClludkl+TcgWNdXUeu3uWGjcnB4O06zO9UYUQuh
OWYgDqbEjPx1GZTXVUSmCDSzJ1hk9TKMn22CeiK5DRl5yEkqPW/+4M6GiZaG1NZ7aEpjHaXi5udR
QadVKMXfmQfXd+wmNBwf4YRrJupnabjFzOMZvy7k4inZOMislsxB/KPmOjKk+nULkaeCG1b1HUWy
fFF9lh4SAmCHZ4gHuTHtQgJC+nsfL2UtSCxjVtM0VzSP04uKPfp9mGuWuZBSRZKU5/Ms551UQ/6s
NTysUPJn8fElpC4xarZuTrqHLcYJYa11e8bRDqvTXlABTNlfNgrb3cjOLmtN0T275JztjBYj7en4
OXgFnPk1HqV3zyoGzu1+mWPibAV1fEnubEwdsYofL9Ny3YrUWkpPUhScy/xDTUGY6kNy3GXPcjAA
BUEbca3NsIy2oNkw1lju/gg7ahti16losKbcN6YfDDun3m4RHVXi3rrbpXqLrwqlGdiGvRlcz8nJ
W9fbe04rqWRVGjPZ6cwdx/BQ/PfOb8Xcc/21r3TRIROI0QlUsQEG+5noWATwpHjYlYpaE5qBw9NY
a6JBy59u68dJG2GU+tPYQq13+405an/AT7Xl+qdVaGqKRvnz6sc3UW/VYEC6Wsw3Mm7uKWG/61Yy
qLMA+RqklgOI/Mg8iz4JEGt4tC06LDstN62tU9p6PcagPaFHGX6lHaHiqb771gUneEimKKbUkxPw
+MDfVOLFHQyCQsjSb8JrIDrdQk+wI/gKJatV4xJMydTczYLmQE9T54CoYqZ3y5VuFT7drEAYksF9
JKsQSJjFQY6chco8sZ4f0JptU8yuMgw9GsZvsqdE0EKE++ZljFex3RRpK+NWYTmfvD9L2C3YW3ab
ufVH9OFsyIIU4PxI7cRFuDC6XzO05x5+rgfyGE42Kll71k9q+h26CLI7ECgljGrx7CivMF21pUUc
RxHmx6aKQQSwxm1GyXQ1sz1qtQ2M4aq7HdKuaGn3EBOLrd5IWfCiXHTdMLGbPOLpMzCoA2VEeo8x
7PBSWP9RzDntaMyYWO3bUVKJFVMjj06jdNJy8yK+HmhLWZNg8pJOojI6qWHwBs+P7ShMF7EqbnwN
cVvZcLd3W5MRrwWcc1KalLm4PsyfXuIOjQSeTl7uEzpLbkr/0SrfSIoxOz8wqb5d7AvlZNxfl4rg
pzn3TNzgicZ/lUqVDF8IJoLiiy5dSlpQBrywgI5GICxE3yMHWlQbYyUnyf28hRANb2XpweHL1/Oe
83Zgy/qWe8jcG2fK3EuiTT84olB1hwGbnr0jK+14+CLpZI81TC+nIxj5y8YP9KyWGer7NdqQkRQj
OphjRHPEnw3XvwglvwtjPNx3TUm5tSagWgorrhUffUPeeTFzo8MrVuXzPJGd2CJp0RaOzL/jidJc
IH7z6ueqkFHJesTQXW1oqkjG0ju5VoylzSKVFQaMCeJaC9WsnBeqJI8MSsBiXZxfev17HnY85g/4
vk+amOtbjvDd0PvXU3fN7ZQF9XPKCZ3Xc0wykbOx6TjBzAejO9t77LiEVvEiPWTw66QnudUmF6Sk
Q/v8YDMfARfojAFVHprWxo1ViYjk52132AHqqUTWtbiyWb5Taaf1DwIAxYsY3ejylwN42tlsrISN
PUzuMY0UYD+8nUXb8q2D0C11bAPV4HJ8HICY4QtCIMNcNZ1INZ9kEttmHZk7Am6KQ6kobvOK4qoI
h951dUtiAMV1RTDKhvG5GsbEeQNz8SH6+q2/H0S6mzxBLTm3G4T1r5/+LP/xEGQGQKy0P+HKZfsI
bJbysvS50PH6lefW7/dIzTk3wJJ9+nOP1smEpzxHorcVBRIDBNVEqLOOLn0LcWw4WLiK67oFrcOj
OBV2GGBwyl5+hcbVL9M2YgFzfO2lV5CzxjroT8LZ59v1n1wVLkHoHjh3Oc41CRimrevqAjUX+774
qShYS7GlNiQzwJKyvNGRQFwMwdHFcqzhTqRwpfcsFP+n8+3UryZ0OJXL7Hho+7g/xQbSNABFSDy0
0crYFDun1B/yl3wAsbxaQr8esuP4ebie+a5Hcy69827/tXc564ck3Hw+3SWjE0rUZQYaaemt2kYg
rR7YFJLk9yfucAri4pyGwwoT4/Cf4GvkzmAY/m4s9KG/s38pK+KhsZhO6lmcWLY5RyVYr1KgYIvh
+BCF1vLjMtr1eYEVXdliWFra6msafvtV3IKmOTnkpbfI+GvLJ88B1NbxonKaSjG7DAP34LXR5ZPV
gu7hKXblmoy50GuEjyxJ/KxxSe5soGe1x67RDs2w6AqH1YJcwnzryyiG/6aOyLU+MQssXFfPEQ7w
1wH1+uBMlZgCNo/UWp0U3z824e+ohrTkfXCWTteFzH5YifVgm8SMjayFGimX72tfL/iP4dG0glU8
rvq6v8Z5jYdCXmvYgU++YI6hFJrl2+sCz/k4HhgFXuRB72dSh4XvlXBmfPtD50XAiVEZmvn94049
A2gzA0a8JPoqnEirowPkEdStnk9WjbWxOfKSG7vNs3M+fGJqNOn6ZBSd/IXBQs1G0WIFzPIeH9uC
lyqCkKj7Ej5DoBV1HRVvt0GR4v/WNgY2LkhSs4ANkHlAV2eQCPIqCzuNjapoVEIFxNHDd6ure0Kb
duIKSdhVy9VRS31qI5qVzNZEF1hOM88xw8u4MkZ8T4eH4qJj7NOQ23XbwQxzvQZQ+NWIXX7I8urI
Mrk+NC7k7izIqIL83cQqyC7gJDTU57zOa1jFWCMzQx1jJaBSoTfc3NKCpFrx76Skhygwx45sGM7P
mDmo3FZjykCBrRlmKoR+cJUY/WP8keqy50k2bm40fUIn02mYEGFksIiV8zuOxndpDVAcxVE51zPF
MC4ocrVW1RXRf7E4oE5SUQsLB78oc06sz/B+YIs1/C/C3YpM2Nt/XEFWC8Hyuz9Hggt/Q9+oYEP/
dIayZd454KxbZpjT/1qf2TjpIdrrG0GjpB3FQbTZqO//B6Gw56hzfq/EEm2+LJK3lk6K8nqrNh7I
CkAALENEjBJB7fqgJc0p/m9U5fziih+iVh18SRRQ8MNjsM6mtFiiPiiGYbZWtoXQRM9rQcXxXmm0
syzM0l9yp4OWOsTIXfbp9f9oHHoWnU9DrgDq6aUfs+lLbTgJ+YQbtvZTmZIRQqruhzh5CNxp/n3L
pQllEFr0oHwZ0AHvJEAkUcL5maiS+jjFLuTZz1vvpd65L8oAkspLRZ3nuUnh6ZUPfOvYAij2i47p
TfVAKK4shzyqctGvPcPTzkpEkvUeUv3sn4ZkR6M4BeLkTTA1qQBKwyaorDGATE8WF7rTTc4axc1U
PZ4kzbVwclFCfE00PoUj9Q0W0LwhFD5C3Z4sYmg7L2OE446suNtFOCDNMCPBoxNFParORAtrnDVr
V+cTOr0ABS+QjH8qaqutbSLq9Q5CR7JVuEwex+TNeU5F6H5d3zw4DbBVrU55Jvdbjrwf6pXKzHSg
TyYczn3u/6zpzauhTvz0LcL5e43wbxu+6/KNkPsUfRoJ+iq6w7nYOXkEiNQBM2aXicWR82KJIPaz
g1c15LFHH9FCTEjYpMZ1hG+rN7m5/ZQO6+4vdmgc972OQY/HMu+9+TX+uYld6TGDVaMNQDEBkxvv
m365BlCaQXbrGjtCuPODZ67AZcZwZkRFfh2D2x3yKE0fxBh4hXc93PiqYb6axS7wtzfeO6POy29V
/wlbxeskOIOsJ6DM3YEtza90lLRRgSJgUz7pNcBSRTQTGxO8OSIYzlAVdYWbS55GH5Ydr367UCDn
3TBsX7YuGAnvLIrg0UjKFKa0B3eKO14jjNqvhx0+fBwTege2354wTedXeNFyF6yM8gdV3HXxuE4z
8PsHFqGh06lS0gmBXPklyjyCV0842/gLH+PM4a7tBSHIx4LxroWhJMSc4VVn5CwN9vICRhxuOrMK
WuNCl/0yaaFZ2Gzlq3fjuc/b3xBRvRrzzvgj65ov1fT1tlM41TPr6TPFQQ9LrvP4rkM/27J5ut+b
LxjlHdD/17DZxxAENMctrQsTW/+983GqwAe6CN6MDIJO08buS7vSgO99kRbXaxRym+ePz+7clWwy
N3GiQFyM9WYH8y6jG+b5YJFWN6FmAN5dnpnbl5hm18VVAFuLAD1YlBLTkP/vNEDDmus5+hPCK70l
aTtOsZpj4P28ACpRtaH7jEhSGFfiw7k+F+rYDBYKW45TaG8BmtASaYXqfGy9GUi9m53LVj+z/gv1
R7z8FeZegmOIFLffmVNq19p9JbEseKMCwK+x2UdEcNBaWBNNv05Avc6mgqdv5NJEtBaV+M/zVBo6
/CZWjq01yc5A3N4WvK4KYWkYwsvSfs+wJAqpTn8gHO/K8gCmtwHI3yrL5iwutUHFABUN2qw4KhQ6
Em/69TVd08REtqPOKjXD5F7up9/dOo2weB+frGbxs749vwNSisFizTrXsYfTMsG/FH6OY/CezziD
TNomj/p/eLCMJrlZi96C9cyqeUUM1nGErCQlRcpsQWdvmV082LacYeoDoewo3nviPw57NG977Uw/
sAzvgADeKPLZCUQ5jup24zQPFeNJFs7t63a/W5MvEJIn0ANPzOuHHEa67kynXGD/etJ+JeCHEdFn
aI9YYsFz+APGtnI11UCcWYudTEYkGbrdNKZUWZhfAVzuqu0+5+c5UP0Loh2DtM20j0sJwlcIuOFO
SkceOJQKhfPRzwaK3pIqeeMNfAsntn+dPdj0FFCyi7COvL2vQA/EojfZT3520wDx0fr2It9zfwd3
0QL27uOpK2u9tf3cwWdh7VvL3FYwOdGE6cNS06wJYwVtVywoANHiZHjZ6Bwk1BM5MuBSqDoVRFrh
/5H5yeW8fNzK7Q9+89rNlPM4j7rSSsxeB7kJ3oxbNEcDnjWmzfoVHWHR1Ccq1Dn/6t1MPd7YMl8H
p8s/P1OBXFms/N+yGcGhPW5DKgX/ZVfIC8aSDqBkeGcTJhjBPmAx8z1jlef03FX4qt5vzKip9lgX
zgH6jEcJNyI8P66mz3FwZNs3PEmXOjZdIm+oPD6Z7NVkdXIoi3mAWWpUkSFq1M2X5FkvkPs+QtDI
gXWGWRB275Qxdr1v0nYH+RH37Y4guL9Kw5W5PkP2sa9HxoWmpSVsBaM7cPNxzrDQKZShd2PHVQ02
69Bc4YFPJPRa8E+lj5Djim1jGO9l6NwiRtwDJ81yrHt2LkoPnwKPk0z6vUa83XYb1K2KI51IdQug
FmtkxX9dW2UCxGFQ7feDrVQl+wS3/siOsSYy9F3zV6/z2Ow9Ldxj0AfhHm06dIvSZR4WZIWr85/X
n0LEXOdS6W4/3X2LAX9MhvtgP2tWbFvYq9dufNCOVpUt6hMZzIAR4ttfq6t+c98zeBptAXmKx+FV
fVFCGjc3Una04X7fpNCLKKEvrr87C8sLrRB1y8SJjVam0N6C+LUuMHvjNFw26UamYR/sHTPlNrIC
IVjya4viQG2hLIt5gl//uuyLL4IBqtEEk3b5WJP5rN8IzJfTkbJRxR5vOmb6jeHMMCCPVIQkux5k
6/Bh+bsyAr4qyxeBGFgR64x6Xr1XUDqSaMPtrbW0d2xfOBxLJx573/aZBo+/3B7CNf531Vin0Uap
UlUrrFWQDGA/wbz1n1nYrkTNYx/R5wp32a77/S3IGwaXfn5/TWcr56gR14U0St6evM5duUJ3BI0+
f4HxCT6cRsKQJrpTlTRHf7706IvcfNUQ59+NMOooiMMa4Dv7x4fqu91e9DKRWz2uSNG0eQXdklkC
Bt3RJBQ+a+ueh7FSc70zsLhlgC50gqQPwPGgMPKRUFjiafWqLPHMjDHDejA1DZ2gVa9cNpWHNfUH
He4NlpqBraAFRmxNVSOad2qJk+nX9JjsnWUgnVCXu9NlyNLrmuVZlRvJBraJkpO65WrPzOO8D72Q
GHCAlQXIZoDmE//tgBAkze2mGrPaO/utedSmk0nWaZk3Wh1WzLUCBXU+1zyBQEcolkt8z50wOyd6
e19FZL5g99uH0TnDmJEn66+LW/Gs5ro82TzEviRXkdAtmup4cycrZXY9Dsdp3YaPvYL/e5tVvZnp
gCF1XJAuPSrMXV2Dj9QRO/jZgnQtu4Tmthx+A5RRrm8GkoW9zGJZ3KaqyUo0/wWqzsaVIeogoY2V
Hrm7auEELG9Ev56KdcyKtTulAjXCeNXtxGHIvaXE1XosqMaB/XAKlDWnT5qYMoQqVC2A0v7HVTT6
SLGNYFQ/K9U+gUPzHEU6wChwpGWSBmwp15VoVc4Y8YWwnGGzHQjBvxBVKgYdQQFSrS1qa/i4Smsk
OoOuaTshGRbF56gJB982ZEE1CamV9TCd/LcsQDCvS0VHt91DwgoK2ArLRHQy+TibQW4/cwWUx2c+
Trf0iTnv4PkOcDHTp6E9/IiV0vVpzGKXdCADM4ppvUS77KtGizOb+qedqYjBM1ymnt6eFsSsMye8
WiFYRi+YAgYVzsNBFtc1MCWEo44nzri5L6IKlCIToupV+Lnx50mNkom47pGMZ9p1aobljvhw8HvP
hxuafoBHLKy/DPkSAKRxhhDpszlTaBUnNYqk+zu5Zt/8RP56ub6hmJ9VY1Cc7phi9HsudOy7x0FZ
T7OYpXdbdgErQqHU+EM9zAVuLihc/TQ+UVYabOryD4ANLe9LHNwHYjShHtUoOlOllb+xszC81Bob
M0M7yivE4TH/I2A7cfkS6aJxbjBom/Lfut1J3qlKGkXumL3Fa+pZ29DYMeIBBI7NBpTTtxvpLwal
FCG7pvknC7PmKSbKy62JqgmSHIUVXuGtKhUNfM7wraFyl+FuMmbH8c0MPGxDO92aDj0/i1O2QEvE
LwOm/4FsDOAbCqoMkbfKNOkqFkfZU56uh7XEujIDCHNw4Aow4L9T1K1jeKp458ptQ8w4GYvXN802
DgeZgk3alRD/udmtoMgdd1XPOIE7z1UV4XBaXwRgTChoUt5b3CCJq1ztouOqNly2RFy+tczBnRvI
gDGpjccmlr90LBz6rCP4+JXVuH7PZUzNOsVRlo5h6xUwUng493+rsv73oyL/ZSuGo4JjMX9lKf83
c93oLs4CYw+afIHUmDV41WH43qqTpZmYK7WyWXoTcDSuDNOZvkbdNXjUyPuqrtO7pA+xWot9/lC7
cZsaSndzi5Zh8f6vWKL4pMnezeNME+iM976quqlsRacJAnas8BlEhjY9avelJFh1w5xAg5aEsCbW
DrzGwJsag1w38k6YdIVG8i8gx2+oEIrYfWUvPDRP6jNNRhi63enOr7h4KgpxUal6J9GZ9fDddQUl
e0f/zhesLnVDlz/v4BqecXPSAAs5BoSrRoav3CGpSOTtgHvJOE8dbds5TUzwp7HyforFikDk3Dbe
tbLN/j143XlW8BD7ERD7Wtd2MlHsXS+sPvOlcsK+HBa69nWX0bJfh63U3GuoavX0mzAYeIVT06u/
rnFRMpL4EYOQ61xxfSwdxD2krb5WheFcL0VGS1JSte3WtPt5XP7RTTw+4letKXJhTD0+/Ca5FlyE
7jv7hJLToqHUPXHh5Bk/7rXS0E5374gTgR7LSNuMcdQyRFd10Yk46xjrIUj8/i+F657KLZ0fGcKZ
e3MTtRe3t3u4gJfyn5b9J/5SywiJdSJh8gO+s5/Q2w1yhqKYOutHJjd9GLyw9YfM/5V6LmzWiz0q
4IJb9MHFRR+XaZGVtRp6IDZguX7QFLQWoDqKOLqbkbXrfOThcRcWqoL6Wj9/fFE+nQofKJG2ca4S
+jZBFwv5Z0t/WOnxSWb83hXOVDj9uQPtHe5QKrjt3ZmkLQde/GsCNczIG+D6XwMqbtRklZZ3gkug
whl1iOrGVn7fHrsL8S8TIlzjLWNSb7qeanFBW31KIyxHB3I1Kwbp/RL3ZfjdVRQlClj8qoQGlPsT
vTsnAFeaH85WmCpnTLLuU62ULG+Ff9taJAcY+tt1YMG0gz/kuYF0crx9OCXU1NgNm/VtLgQNAzPR
xRuf/Pcwum0j8yrufqCIK5EZzIJvNunUZ8cKrPkAWMiPYR4zdkNiXJa5db7Y2ZPYJGMSkj96n9UI
rARkeGjGUfhityMRKoZyP33lmaz6a1D2DhuFoLVL0gTqEArrdOUQURj+001+SASmIOVWN0iHXAg6
W8JXODnE25aDyzaKupcJmSaEe6IUVk+7k4a3HKl9yu03davYqv++lCix3A5GSTNu42VGElnlWTvW
mWftXYeHbR8lI/NPTdCeRK43gPgUn7aPsjLg+z101UzMaG8mwnBB4eSWxOujRQqFf2I/mFcd2E8A
MB2+HOfJTZHjSlxGg/vIBJT5CE+ks/62djVvE5WcrgnEExdMRvsYO6wreGRtsdE6w1vty5jq8Ncb
1ctb36kNfo65wt4r0jJ9Atxk9/5+mIj7xyK5TKfiSFxCJ67VQc0TUM2f73WOD5CVIvSDBQ7OZyeF
cMRXUE4ZYgwFLQ1NWBC1iNBB0mij8SAWLeeQxVJYAn+OGqnWwmSV12PUy+31RxQkA6kZExheSDiZ
aKQ96Oby6Xk0A+ULDajd9shQSqIv9xMwFdvpW/EmqgZpNl6/oEbWbRVyyL/CMfYri1b1wKxVe1qO
75baxbm+e87e+QBst/B9AxOVZvttf10c9GHz7yxl2erNoCU4CJmOkmYmRxi0ejHKf7rOP93T1X4H
f4opjrWwiuM7YZmEGero4qi7vd+H0ofYe4aqvD4ZSMUeVdml9dqs006BTAQySmpXoEpOIkuz15ne
KLL39A2qD83hwQV5zVnHYiGz50+CyBfVnc5S2+rApcqIcqpMIpR7R4NO8Rqlz2/7Z84O3tZkaBEg
uJ8YI4y/pBqPr5iB+vJQERilqSpCgjrTyUsWCP2qLNpDpNTsuUMfmU9wUrs6Jpc0t+mnVzHqTw/K
rGHZWcvJdRw93Cmd8+1mxIdiuzNC7YuLIhgWPt6YAGmeEpjh1WS7lqBiwD5CV2ajtvmwWQgVWuqc
V83kIE8q7FLw6gWddsSmTLOMsJOnzusTgedSfhhAsAPDZylPFBeZeray4othKEnJ1p/J5b1Cmm7Z
/QpQNJuTEj39iB2WvqA9cS3QCloY1SbyZ4H0j2ZBRjnm8UR8mSwKaWUzsyBwCNKgDdRnPPBFLhmh
Vb475LwdKIuP/PGGWgw5HPOaHRd71AHdx4nZW2vyofaT+OvWcVy+VJf4yHvFpL4hqgmLrGes3djZ
VqCMwYbjfe1k93iUucdBo8RA7O1ooeYZX4YnvDCeZ8C100eTLXlaHuZamaKo0bwLpCMjO467HRe5
xmqqKtDMOhpyjts9bLVrLXk3gs9YLeIa/GV7IkZbjgx3FQOByoJVW1h7r2s0awLeSrFHeMo8QlKC
tl0cTcv7kIOdvHfjl+yBstNqb2UYuFYRiw38ln2IcpGvMg5SKycJ97K7Dqy1Zl1aDx3peRoXnKTm
BW6bDCcAYkUPJPF7Xct2bNPEjTJsElVJKY7tkKOErR8DTDzDRB9gOASbkun71ssVwkRpWa9Diiz1
vwnQGa5mPkTKR+wsvwq710BLAMXiGtBCx6ALm6wrYVsUvoMau9Mtj+zRNJvi+AVmHxMWVTpykCo+
UrkYDkq4Z0eJ3olfsOtnIVOoqT/RRMXSr3AG68W8L6ibW+C3o0haJVFYo4aMJK/Y03YncfC/Fmr6
cCN0L+V490raFk4ERW3YDrK8e5JSzsP68v2XaSThPxPTK2kD3yG0blrsk4ZKnbVkMWnxDG5WHGW1
4s2FsuVqDVzDRObEikYVbr0BCJtpknfPgjYoWYml/ar/tswl1E+ImaQLMuDnef6klN0QJMoa5cpE
wEgxsMnvTKM3gFOE4d6hZ2c0Zi2zAdq097xeJc2fZtGkHu0OP56ppZFO+pHwpIMNEg2edyZjfAnH
lGfP/KSH+qcXmtLQVhn1CBXdbrf9tlBVwKcuCAOZ+u3zGnGi38LT7Ahr/HeuQsM8TjM4jeU+pZV8
YyjF7CztEpPPx5e1PnfjKajCDHfMHQffBLPADVGz8o0Rk/epkqotnzWUckMaTQ5gFuK2n21+KvRl
XuDMlKw7WQMg+bx4IOh3SjLDAiD+o3frrElFkt9a/XlNtEV9ehr6iRP93G4PCAC3MGRzcxNf5GCR
isyIqyfEvX36P5rjWi/CDaXcGQfWGEqZ3gG3CTNbGCa16ZDRlKc8yv2O7Wlc+zZsXv5PSVSl7joP
8CN8ElU4fJD4MgBGkMjCt71Y7FVfwKN+u/ou/vkNpajjfqIlT+VzWMt6uTSp498LZ1Qwl5j/zgHQ
069ETHAeuZ/XuoBdTZVS0ySLR7RaxEQzwVUFxM0087w4WoLemi4yfo8YIaeT6MLOl1adh596YG1Z
2qsqmuNMFM2Y+rsnEHBuyDtjb+U9reu1186VJRQ7yerQyZ5gFRIbkTKAamhTuPd89mpd8aRJUJpe
QtcZergFPxQF/ldY2Rssxe9kEw4O/iD0ymsD3Pz7js2OV6Bg+PuXaSj445j+/gvQmwJPPkX8vA9V
rsotXXSEdmq/zlzT+KABSW3ElX6REmXM03PfAAASi4fWhBYgN7EveryjOacaUNMWASzg5sp6b7lU
kmSPTXi8H+YBjxGhuHoxJTPSqbIzM5Wx9dhRFilSMRvt1WXxiya7ElmCfxG4wnqnjTQtLSV3SU/d
Fh2dvChTmUqJox5a8Mf5ahxsd9A/xOzQqIH3NUS1zxWwANF1g582rpkMcZ/+5Du8iemzx+Nszcqi
xqZuifkXY9EPIchSPp/yuiKBgrYgJOSPaG9aaXo06ktu/DAvFD0mSBUuosfGspxoNdhNpp0NRm88
7QvMJTf2HBJnd5Q6uusirKBSxBuo36VV6KpP4ULeIhNYxud5lEBPtcTby/4fatcubJLHkMjJb0E9
40edu+EEPYKrRXVp5vFw2YiDevI7W+TQOQamResKuZmw8Ygcw2wFMbm6Hf75RVEiw6vrAVcVJHDI
OZHSJa2t8LeU4flyengaM0FUDOCIPiPIFyq+/cQOd5JfYDmDZh3XZ5X5wlc4cJcQERIggQtz7Or2
7g5Ex8FKkEIwXTwsvL/cwYDU71th0bmWjdoDoflNxR53r21WUP0BRuMIbfK3dA8Icv90gASYhLNa
Q+Z/gI+oevJfhlM1UpyWBb61PvaaZteR3qqWEpAVpnS0AJHQzFzLDBGsXVyzmRk0rgdDeqFKlnsU
H0cQ0k3lzSN2AzJtZ9CBV59F3zyvlPg4A2+J+I/12kPSYInazMUNKaS+GP5E5JaUtm3wKuUpNmFD
Fme2twr/41BteHPW1ib0ZRXMwiWgL/NcoHe6Qc+XKtb2oNswA24ue2DFP82DMzRf2ax20/hnIRet
feXmCm5UeqNJpQHqsNn5wbcDYwxROtz7z1H2VzK8QUM0EmAZQ0tquoMD40P3tIFgCsi46+nqBUVP
ug2+2WG6faEhW9W4DSHrC1tTWcB4/pBLwZfqn+AI09Po/wccc4oWSeDwEtfv5Ej/FZHv8rpkayOh
5UYCRDiAK3d675EmwIoM//D6VUJAF8Cb/LGi6MHqavq7ha2V5SJvFMLDQOX+Z3BBPu7pvDyF8Hg+
hCIqsWQMMg0ZkTMEHTawFDil/2VmRb42
`protect end_protected
