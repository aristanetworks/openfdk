--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
dWL1rIxcJkjin4Cjw9pUDqXGbt82nGs6PDE+SM9pnNfsqwx+0tpHK05tjY+eB6QR47YEoGyAVz7u
bLKOyZZ3ckvX26EiHXaKvt+viev4MkdA79vTvNSleeWi96+Hr0RR3+zP3lbWUwrHX7IaSVio9RAV
TbyhUiED4exgec3NtEEAgj3PLgK9rlnDSdj1XQp+ce+uz3YjkvG+ZcCovYhkkDw4Ica3B/8B23Un
c+SnT3W1ZpTtVXTgEPY0aLvyOZ65SlaPkx/CjgMnUCh0GPvVIY70FwXQRTrBF3k1lBqzv3J91SY0
EYPa9oOvWXZ+F2z2+JCCkR72oBz4P7C8qH5XBA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="b8WuErRUX/ixUdWxBPEhERz5+LtrNcs+wDBRg/NHp2M="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
LewqjQQW7Ql8Zof7XE/qfggICzSEne2UwU/c7wmwLrR4MvGCq9++qJvbkY0lm8EJIJL8B8gx42Xa
l9t/E3DU1txxvPZRJRQBPIbHuO3uFdT/4w4j7bE6Q3s7hXOcxKpbxKWwfnFu8fFnsx7ESoFiqiYF
5u9djT4YT0z0CqJ8QYxXnp3VBCT5z8+63c0vWyakCqiF0xNaIDaSuLhAD+ylEE54xz74KHDXuD9H
414XZCq4GviNo7fNbH0Owy63zf422UeL4+vh93b1A2TIYxEe18r4DleIvY8U/tl8LnjGAS3/MLXX
yhwGW131Tw2+9uItkoL27oD7VtcBuKXLVqi7Lg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="MpKzBjjOysil71FiEWLVoFXnKqXZluBPeLYoLcSzMnY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5616)
`protect data_block
aG8uHJ5/hUkJI/C63FLK4wynJTrjvfcPm3dBlwAWKpMlDQ+npc5vEajswVjiONakVJ8SdSRdfDQp
GJg4htNJM9bTiTAm5pBfJv734WYyPIdlHPIJDIe1/TWDa40HXwxyksk035dVWwkWhiX+A/8jns4J
U3H5+Neu327gxnoVUsARG674W3XKBiiRJPdE9kEWuNoOUkZM7CuQdc1NqcJ5z//2WChpySdOv0+4
cl4ZPyh8C4EsYSYrAfyIZGrb1OeRUA2Z5cvvg34IyO80RS9UsdtvZlZE07lLGLSCwSkYNlHIecEf
7TF3z/k+/xEu1RXwpCLFQH1swRHFCo8IJMeU7sZvpg0mb62fl7ib+UyKkq/XCwwJvRebw7JawrsN
Cl920XAt94a588SzBoC2Xrw1sGcpyfYhrI7fV19Y7eWfK4YlM96Ra9SVQm0tzkjvxQMzvlOQe4JI
dF3/fGUMVEr/YA8Wy37ZI35SDJthQxHK294rbkYFmyLTgCwzDvsnghqGHAJz98r7ZA8g9i6FQX8y
Mm1kM5ECcKYadWQqBVqVzqU5UVKzhNlxB13859KIbfPZwuYvorVn2C0D/Jt0ek3XYfih1shq0jl7
cen23GbKn0ZdO1KXX2aH5BAv7jjYq6fqgBckeP28NlajpXsZ5vd+Tq+twd4Z98dceFvOr47AJMv7
2vMu66b0FuN1qj4URecXnFG8SsPpnkQqdat9PicxQhp91CTqVBlyMVMsgSp7MNc7z7Xqn10I/QYy
NGXc6ihoIMQGRWz0vm64O1NJjrMNl8HZOnnuQipJHEZS5x2Ci3evb01nSbmczYoDcnpJYojDxam0
mPh8I/5Ekh5hzg6xPZVtT35SUgKjuGKtNuB5DQYYA2wjFh7tqUTbGZodIZMLxGdoSF9Rv31cqh4s
xygFqFpqebW6RDo81cCAQcM2bFPYzd4RapSkqbJ7faC9X42GhwsV1iWTCuAa0IhsunKYcZsBmftj
PqzRAR3YvRo2I5mjEj2Uzac8uwAkbY5M5OZg+76Gs6iFhC7pKe5Se8R+0sEMY59Kr/EFjTikyXl5
NatPd0WTW+WoXDaCtCP9VlAUYGKYLULxMrMbJdOYrI+MDufHyCzVnYcuI0aU9Zf1fTrztku/yZsR
+e2y0oKEGqu4tX1RoAM21TYZDiB24Zbfc8Aw0UY+RCE9qJiaLKVIft1iBULdbeDqZb4BD5jw7ufy
kwKneY407VLCtJMK0h0XJV31DtnmcKOKiOqeGkciXAPKN22xiTPXOLeiRU/nQ/bQMEjwca7N8y1x
SWEBvGIu7UX5UuJMsgfIBr3pvhAZGor5z+ZyEqKrR6rhK/Gso5ekUw9TLnX9XvJZ3BjeTRusmaNO
iWk4KZYNu6TGa7hHDKDBL2L5H3eB7pEghZA+MfzjY9fYYP3DnBdIF0LzwKW39tfUl6rDdAZ3OS1d
a4opH9ZFRBBkrGuRjh11pBdLZNLvKwbzYafsvDVjlywqMOlp9XZrUhgnKW0KxJKnan+jXukDxC12
ik+0S+tyaqmSwivZ3MPsYOvl+PBNjBKNZ/pZj6hUD9v81741JbLwTG7IGzqg+p2KEOlaR3WTb+0E
ILVjgAb9mqpOjMLhMDTLw0tMx0gsHzCiaatffHkBlhgQN8q6Ry2A9l6yVQLTnrumI/gTJhAEPxRB
6WtiFO0sbVoPHMEB1pQisyV4jV+vIcxbZbSPhNJVzeRz8L72RpMeDBnidEL90AhCXKYZGiO9JqCh
zqYP0yEImvm09mqOb3PSYg6zqSeRRJVITYEe4KDe1lwEI9tc8T8SDQ9upGmqZ4A66N9hlMZJGqMy
UQPC8TyaSN0v0xplZxDqx7cFpejS6BhaYGLfsPg2VdGjkLXMH69KzO6EdNW02XlaJFF3i8AzCrNL
ElgellHZqxzRSYdU0lzJZnB32jSLaBPRnrkd7X38lrGX/VkoQf2EmxcQ46CPYnjRIMjUUrILJPxf
RAnHB2UrfleeBRMcxVJnuYD4RbmUJ0/Dfko/ayKm8GY1hSOC0LF7L6yh/NSi9gkDOkV1TpGRv3v3
TknONJ8izWEBAbeMbsS+aNjzPQt1VBSKd/MeKBaBhVmDqLu5ZwBr9Tonx668kIJQKUozX3RLfTfx
AzxjjkEaroBD2W2PCxJ7oFoOZ1ak33OQvGveJChKcrI+/lK5CDJ5apFLdASGFxbicdDVh84fh8Ze
pVxsUpd1GxSmRnl9SKdVeWFFg+Jhg2c934BIwrKHAinvp/qO3jbdhvLeTyd61f4Cn4pN4WqcVFwC
G1ebaBWA+LWDEGLM3q2p3zDwPyaLZ5RwgqT87pPO6jKYcJBfBnOgtDrifd2v7PVy2SXVdqfNdheo
5b4Y3w7I/eYgQmhEvWj0Xg9yLF77V4oQvzfEER0o/kJPOwwP5tVF+yMNQ4rY31XDxmhjZXowxX5j
sd1dNrcpIjAm6lLM7n+Eu3ucuCj/VIUhhHmd/Bg1NH5HBjtz/wGD2rt/LtyeXNEUdKk5dEeB0EUA
KoN8feTWcfxXzsHTLDGNuwGUfBjjPNiz6WAVxGNUgQ1i2Y69f2lUWBeenQFwx17mE9Q1b3LGJCX/
yXZOjdPaMNI5is5M+pWjwNeMy461tALPmnKWBfbYUBNrzijUvBMNNx1uJh97HtMfYnR8hnOVSUhh
cLYLEGOPS3dCQ4PbQKYGPkvabDAoCpEls/OWtQkjSoZiBlH1v2JeC0L8KoM5ZjJtwyJX7GECHLNv
l5HTT/x9ZEHqSIiZQy8ZV8i7MrbaQ17tA943/KnyKvOJGWLsuTAf8GoLFW2FVdryrRaTRe6l743S
63HnLlQebkd0oEqiP8dyE9YXQhmTp0Kmh0XqTYc4qpgDrXuA58tkKnYF7won9a1QokIsOGIa4vBy
4NHwSkvTpd2TMJMg+/l/xT+VA6rR21JsE66K8j6jvLzxneJnROPh59hKf0GAf7DDYFdBd3JF8fmb
L+BmSaVHfBXEmrwtc7M41erA+4sm4kXQGHUiSaQfronBtc2vM+Jd6GN4mW5LjE3KrBt2l5A0JS/U
yZmcwF95n3odw5oLTYqEMaixxpHLMrBsilZ1ftqK66H9+AHiSdIFLq7PvsecU/6CqEIpY2/hCR76
u+wDdtOp/iKSmJy94Xy3rja6naSbCtoALCHzlaaCfojAsXleL4Ho9yNwLowyzxDBpbvJhoZsW9km
ior35Y3NLrLQlHfJs6zAyGUC5sTXgQTKk+IqfWUXHSrW+wCcWc2E1/PjtBI36FOZTOcta8kmwT07
oQRLNxrBvgCtoHZ9eL4UxaBipqVWVXtqZdMhUK9Glqsva6bLoOOOQKAqs/BG49DVTY1CIu4TxO8S
zpFSFnYciVh7QAap2YC21q8CZmTONG+t6a0a+2h9vPRD4r45CKlRMgF6HX/lKdSgTA8cyvkZfZgd
kRJ5O20ah9JJMWToSQvUtEou7H9+prJyLcZoq798HgeynTiwEnwaibjyRLrTylNLrZnK56Kr+I8h
VSz+iQSlDRUk1IkmQGXypvJ91MvtjicVKPztXiWZm3HGbCjV+7+Rzh8bJlgLuGT5G4szVmP8oHF9
qw5aItxyftj7EdxjunO2TAJZqVSYu6ir5ceDqAZcSJn2oH32tofYoxM2+l39GZ34wHLy+9yFcOmK
MzaPA9mGuO5sbdu3QG9a8yi0bhBuDVjjQa4dOa7ZsM1MGwP7dHL5g73jfg4Ey/Xn3j+1tOLoA689
5WoQet3lqr0GIBKggCg7nFY1ymgSix/wtqEGIQLnOA+HQq/a2I9+0gw85Tx7ntZMUkV6/ogHR9ps
D+qCwSCSC6TQ7zH+lpg2lfQW3gagHtbAT/djsGfVDPJDKlL4pq+4UbuNjvLkdWbYTmfk1x1KVI/6
xKsoSkVgGI5SEHE1M5k+kTOU7lhGFhopmbph587EFsp+OzIsJYMiBriFYJjPHDeFLbUc6iW4TS0D
GkrQlMr3JlhfHLjHs1JG9SS7R/mbNbLTXIKiIgxp6ySAIoNeRjIAmxkRHYA4zzm7P5YhDKPWymkF
f+1GbSVAWJ/tQdASpLl01GWuoO8gDWuSHIIr0B+z37L18EfccDYv8iOn4wMW1JZhJmf9Kr6b23IJ
X6fYgvu37sFY8ueTjyCVTH0DDR0cdGqjjMxJh7yZgJbWDBWU5kydCXKTssHxUdoDv3Oa2LYhnLRa
ZUa+fdFNEWp6dLnw7JvX2JR0shohtHUhDGKmpn7YtfxNzsALMQzt3j2AzFCpMIDVCHxb0jF8oJZJ
51Z6rxLYzLy8Xhwaa0Jul/uwHMs9fgyqs6M4fRs9fwPtjzmZKevFpElwpADbGWFKmzliS4W//5GM
imNru4rAjC3L+e8kVgnk6PHHHhKBiG6n3LGblVIifckEDhHKV+aA+Owg9f6eFXpXAeiWoyCxUL65
ken15Nupkt8vWeb+1tN3aWLbmQMSM91CzN7k2nuRP4PKNbd3EByz2b7EJioJnaRG61kgRtnWvKjG
4bJHkHKrkXadF13IQfsoAY8uPuj6NeIDEArwnoUD/UuoHinbIuaXq2cMv238kQOnEmZ6eaXh9vTH
y6W5dWRdDck3jyZibuJ5atS032nd1JPjhjCJ3WAJ8cr1raKTql9NHf3glcZaiQgE7qa5Vg7CHwG0
+WTglTl+82kihL27oN5j6MgACWSo3rz3U8AMwyCBS5+3aJDH8u4ko7oZxAF57vpzx+lRm01STxxc
waHlGvPwFmF6h25TQYXEJKeXlnTmjRpglw52crStlTfL/Y8PHYnLsSV1IfUnPjdfF9eUkjFH+sz0
RFVdQewnftKFCb+wuWWuk4UgjglfXWPabqhRlbZQ3LVBvsDCLH9qmkl4wMWIY2r9GXqB1Gmm12L7
UtlKYKLH0bw0WWxPheYpXG2ca/n3sqPf52rOKqwzkoSRjMgyHEkuoZNLqOa1NWjLGfMuyOU4aNXI
l5JXSJvZ409n7d1q6D7z+awc+x3LI2/JJWktxLSZcxtD7CoaQcLoUoGps4M33znEmCGUCIq5BLVj
voMCIkTnQyMrPqbQFTnOhPSWOK0LrjnDlxRf7ZwuFT55a/PkNtmyNWuOgrC0rPlj4ENrQcu6vcHh
2xqFOxB6jzhS6N9jyGNQhVY231y+/yIhYO1ouhw1sWM0PS4/bO6NaOBOUBVc8nXzw6deMcuHD/jz
Btut1x3SIhsaac3r1SFKTlpqjBC706t5KNdTcJP5lO53cWYDdCiME5wThh1178aPjVAZ/5hysD9q
nkaiy5RBTstHolciz7HmzCCHZYDS7J2s7zfwDRNd+NIQwhUsoBZm5tyllnAN1uM80gY6a5h8Wtt2
FGmfu6wUpC0sqpymaNtnEifIcKRZ2WicWtPXYLqm6W2TPWIluCkJusw+v9sqjKQ16+uklX8hK/nq
EPkdCgidndbAcuLCiReAUvcpfECvlB6bKcdlw1kgH6ChmpQksaSj4NndGSjyKzRELvbedah4SaXB
kR+/iA2WiZ3By0DsZAcAyyjAkqL9ILuBgcZN64HWFqP8e2c+9aEKpGyaD/FFmHJYrlVEuW6ygD8H
9e/k08LasM91EHYWxPRGpLs3QAw/fLeCUb4xbqgnGG2L0iHQd92mJqd1OYOAFWm74WaLAsS3+Ykj
m1SNN0/33+o/z6p0qUB05Z5fOEgwrk0wV95IH36wRQCmVadZTAY8Mv7TrhdjToUb0LPj9HohM9Yt
JL2ykuy63mmYFm8/DgALYnsyMypgmzy4q9mKVh1mrE6D2xHED08qk6Ti/oIoa0Xr71vxju75zoGX
Taz3+joiEWPiojxWuYHd3mFm3f59ZJkT0NtyOz7ZIFr1cSawF3xuYTNslT154oHQinWfY2Uvd10L
W05bhwbg1icaWiqoOpeu4YfxTLNJqLEmY22yTnnMmNTcJ2blxdPYvlZkpJeS/NwiXwzjKIrWz9Jy
N9SRj2BhmPO9j/ivnCYz3S5SMLRvOEjH60DF0Wmpr9gQlF5i6aUiuXc0Pq5h19HzOIv95OH6x47j
Kb4DKhRuWmgKbqYiA1bIfxW5+lUznKejy6BvpjY7lG3B8Mx7dFUtzvF12y6FlqKtreTgkonpZChN
v0V11vecBcM9FvfzQz77Te1Cinw0JRY8zp+WLZuA/c5MZM9GzehoOdvcujbwJKlZ4akTHRn25vcg
4KMKr9+iDkTpH3ljn8I97wL8gkPJehOfdSSz9Ffw/wNrEFF7lWpbYGdBq0W7v9dTeCpcv8gmdyW4
P5qUje8JKAZ0w7bu0gQRncquZQCFp3EilleNei1OUazchyy6dOWti/tfvKXy4rgoIXAOBGe/9T1A
y8JZfwhzKDTzxDqp5Ucb/PX+rXy1ibpsNvBDyiLAK5O+9FtQC3d1g/DaUx/+CI9O1K6q/PEbI+6l
CIt24JIY4XEHkK9tSn8UIUSKU1mhFYFg4Yxuezm3Ql8YbZ42wKxEtWSRarJNwnJDMYpUtV8pXzp+
oK3GMKjJtNa/IWC1TdlExV5ZkhEtChADIiyt6tkzeGq8EvzTqny+8kuTwldeS/3EGhJ7DPNz2CCl
GOvUHYzf6yTp+B8pkbxlDNDZIg7EzQ/tstmj1kNuXNy3CTt83YChPQ6glhlWfHuGBzr4jqXj6Njs
AwRQdPwPUU+Di2nq4iwgBkbaV9Xd7JMJRih0LYVbBvHUigSPPIDVNBRDWs6qpaz1VME34vd6daS8
ma54dUCHiIR9ip1+7SrDJk+dQTYb8vsKSDlOMRjlvcJJMTYDxYNKmfwsPOiTuW2Pys+QrCsPHbrR
8QwnguM4ec2fm+v2BjgwbPn6VA/MUqps4b6OvLeim7OrWVs+PpzXmjYTQkOYkrpRjM0meCNMOwci
odBiW1ozKkvNoMVGpiYUVdeOy7qnMNwCy4cy+hFl/vULtGielMHqcWBuHvRqJqf4hk/kaluYxCZl
lMPj9bOxtRnma00Z3l+7Ow4IWORf8egZzKgkatBtmSO/G6pH6ga3EhO9gR/95XXluZCU0mfygH86
4AC+SNYg8+HubZB6HL41vbvQhM6E/W3eeeYQSj6bG199vuU3wjErnflYjaOxaOVI8T6NIFHg6+0/
+GB+VfUho8fU4n7qWBp6WR56fqN/ChV0GC9xlHClXfhhxxUhL69jPH9rlmz6q8+w9dt58KKEFVkF
d30MStDrKi8UtDwoTWdnA7n4HYPeI3pyOI+XtNoCs7FpA7U98rfnnoGUgFBgotM85DN9wymhYeFJ
eIij9AC0VJYHxTte6uedipee7IIcv6+njTOco9RIWduhP3yGDdxh8WYkvhO46aX0uiPInR4VfVxz
m+pMwsZ5E202QVnlee3LEvivF6+3HhOuKiXibbIOJZaW0KHaxKTaSV/9R0i3lYQeyeNXeYVeqVm9
4hu052wpRTcyWKjZYr+IRChlUOeRf+UPxJVQ/u2VPKUjMgdlF5d1cEp6IK9zoepeCPFaaZAIND70
Q7Dt7q+DJ1NyGbbVc6NtWlpmgyjtCHZmAMqmGujD
`protect end_protected
