--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
N366552fTja4pSEIwSLHcRchvvqTXsSmoLdIMWuVl3lCxhpnBf3+/7USItJPVHSOHTSWE7NVVXmO
k43yoqPLHUgF9B/oWhA/rNektiFfynsSc5+CANdu00A3+OdhUy74/ck2H6cmNw51iw8sfujOJtK9
SppKvOUH4TWqSZ79H4/tmFJb4mO0rCucykKAeKjsdRRRcehHquiLTJqTPqsUrWZGmdsFnSfyuRGo
Piv5Em8lnW0uAaF0FiWtZjaS8CtODDsyoAic/aFR5HW7yYRJJ5pzn9/adZQc9fsZbFziE1jZBD6l
nICyfwMTYNZY3FoMRkJKG+nzI34RevzsIugx1A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="OgwH+CXyt9yk/V3QUXhghXGnGjB3JgUcHW7Un83Cv8o="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
Otph+vt+plQxa6mT2qHuClcmDlbKRgzaFmTapGO7zdkDP+JdyF0byvleyBNVJQLxhilFKBTXokq9
yBQOeGU0Exi9FqjnB1PDIuWQV/ZqRcnh/b1m2TSmdiRRJm2MIALdCTGhR4nGv752kuRYZpJbBeoU
s+BEMpru41CaUtB/vkeGrNDu5oHLq3bp10zUC2fT2pciB4qTrykFa4AkHrIOgFTnUh34ZVvRtyY/
vX9YdUxOfbcBnQkMVXrMBscKN19NuSQvZkEcX06/6itJGjHt9oW+sH/O6/q9W/+HIjgEE51Rpq8N
6Thish2ViTIFJDZd7j5qCeTpTs8CWwfQvVDFXg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="+4BwPfQLVuUU5uXTaMjFpByhxtTSxuVo0ySTSOU7M84="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9440)
`protect data_block
ZnZrEM4MUcFJO45HHRbSNviVAfWkhfk0RoLNGzAzE4D3GODHxUVvt6r9w5j7HbcpxF85eqq7xezd
/C5GnQZEyyOwczkrbNrSeMcB/osPi0/P6idWS02BApimrW7cwysGLX8aUjRJW0Z1Ms0xlR6C7SFt
U09MYaKzn74Jq090YNMqdUxjc5qyGE6Yir3VdXqaQAPTbL4eOmvCu7ImfWTUSEFU8Pixd5Ecoehw
WeQJF2fm1XabmJMk2MUnUxiGfnRK1fzslncHxp/xBDQcHCE3nwniaA2NgqikQdscUrrA/ENGzF1f
jKd0S9Z8EExEasnuSoONCfOnWeMjSypP1tATu5DwwA0y+jCdkDmHisg3K8fbQe3vmiGnsk9ZhjO1
n0JU8j30U7qKtIsrD/Y6xUDYYeBv50pdH/2SQ1+lGnoYvMYkUpeoO45p8vXeZo/T2BtMZb+26f6p
lQmeqODXH17ZRiPtGCCcwSZI2UwGasFXCCiA+OaGBhszQ780pS5R6sbT7we6eo7AS77aMgo/Xwg5
QZiAQaJ2lf3B6RLesWf3jcogU7M6nJwvdQYIgNHeIZpXuSgr2CYedxSpUvm0cxtM+b8fCFll0QWK
EkvLxjTOfrZOfLB5bQCQQ6y4y0k/33rObcoupdYo278lKkE7VDN2YZvf6uGnvcrew1+qi8rVs+NY
ag7eSjVpqGxo2EfaiX5+AjKB3RxEgWW0JAM7QhYTsU08bUbE4aiLeQUIUJoWWm7iaiU3A23k/vSq
TBWvO3hX5ioV0F8a+ydrQM+cRgnG4RdSgSmt042YXPKizSSW4pG4OE26Klov6Fhvr5uxGn3fIMrJ
HJymtqzFaCrzk2VIx03I/WZyGzRXK/m+SFN5o50nRlEG1ARKB/AGjx9hvGN97gSY0Gf1P4Fo7Jx5
+N4KHIz0sleFm5OY5JSFp33ROWMiiBsAlVdHxIWkv4P02+yH6m6Yw6tZWFG3YPvDtJDDRI14atGx
X6xxXo+T9+fJJ3RA164vHh/BF/wDtrDBbnVPSbPenPBcqdSGXTPloxYkeLa5dqfbUM/tyW81+C+c
kQZBnvPcl94I04sXW7VC1o/XQWURINagcBEw817hgk1KElkkd8gERMzRkGd9nrt9aFKgDmoLznNw
rmaxydHEh+OK/rbsMY5VyWV+uq7G2kaZI8GwEl+52TC1D9E3pzWLDPj9kqmXXfA8/UFcXGeEP4aB
FbIx2W78l06Q0LTV4nrfwbXR6IODF/frhLbsXTcVeU/nnf16+YBV3cPBg4XisGoLdRhvg1M+6rYr
M1yoYwSqgpXm4YniJx1rlWsbjJow2gjeuMgVQ1hTQS9VjLVJFQmpxltMqjFf96Ud3wGs6kP7dWzh
gP59mPlBmCDFXgamd605xF3DO6rOyWLSfZKXOeNbLCcYFgQejC8hCWGoZ5hAxXgAmXPkiVlGw8us
Y/k7o+m9hlNfwiaLkhRUBdUiKGo7m6Fy59kH+7c/QU3POIq/XnCYEt8A1II7eBAupKRegH0u4AJL
0npo4bwp0d32qK7OnSMRESOBU7/aZFZWxsMqRRbPiYbFMnA0X+4ol2EhiIQCCz0NTZeadL7Vfb2r
gvfNKhGnjTxqP70ADNERsQhDloUfHzvqKCYdVpXh5aND8GS/6n5bhmUn6rKCYEeKrblVR234Ve2d
pjdjfABc8hLqwiNlbhBBOcaBIpWZss0+c9EWtjgcwCqn/d2jmRYk15FbJAjbtrBKAQFxnxN3FNdQ
acSPZ/0nJro+ZmJidBqpmuH1vDTDFTVfTexCVpwoaTmqTlr1Wf0D2hCKBlSTu0/JLs1fepPpcOn9
pbz4/fdasOLtqmDkGejILcXC5rGoZSbYr+aCYUlpLdUnI3pN0Ghoc6AbrAjdzjnbreWjL/fJ/mHQ
6C9JW0+gjq3x5tc1LSH7GBMXAkaN5Y1dKJ3wUD4K6Es+k1d+Mx+Zi0Ss2PktSqi3UC4cz+GBQyM3
G/KKFEaRMj+bO6fS0qkeex8PTVHdkxf5K8NIlCSoGfQ81bDD7zcmGnmbWpfr82N/hrb4r+vlwPVn
mWLX76ylyjGSP4ws8Wc0x6mFzO1GcuPaDmID2RpC317AIY0W3meI3evWnbsLcPhB06AxpYMSOED9
YfoUcsHnHwH3Am5F1amvv651+uPcutmJCl1lvvGMBd29UGDTStGmIH3rkpp1H8I8QzDQERyP+bXO
5QBFjPNt6fdSdQOjOrVrSihIbGajMaOrqK8nx2jzLc0rdaWP0lvpfPuNxBgXdYnGeQwHtjM6Jjtc
VZ1tu2+xkPMW2N3i+Zv0aI1Jy3qTdjB5EG/mEgeBidqwLi6JXVHuxLJMZRjxFQKoFXTef+DrDjt+
S71HVn0a+8iEivjgvPKR2q2AIlUz+mnqrFderbBGkKttRGlf4QANG8bbL+3hlBFltGSwsi2KJOkt
pkE4LvWvl0SLet8+Ky++8RAbDYFl9XW8fRnTGPLdA2gE2whtcRVKrFNDCmxEcWct6mD0YG+LhlOJ
J0CN4fmdLNtd4bYVyHa4QQFnEHQM6k6rSNj+uCHbCcIZcdeWJ5DdSSicLs63E3kO9bEQ0P5bhtW2
sYgck1Qb7u6EBV2hb9Gzg9+O8sb1w206RLxmdb5KEU7et5irTlH2g9Dc5jLk/PJudmvFEuqo8Pst
kkUQlxhwTZUavfA12maDBM71/tY6w0fX1KIaGr6gBJIExDEvNMe/VRMlnu1no3x30FJy/KX4ngzP
STvd7tQUD1gfgl+ZXG1D7DrioYSGQ/m8pxicwlKyGrUtMWoC26btnq3PgI9BYFHI+Bmz6K6RAsxo
3YGmJ3d554uEyikiE8KPhln42eMxi/Vla39guTsSBxskqmX19zwfq9pRB+GjktYc2yChOwTtvVap
UWzkcm6S6szPhaPG/i6iS+cIvOIBdITD+1TeEru6tiUQ4x4syfSM9d/n3YVEIP5Pf1u9QDI3BCUw
9HxixWCYnT9CiiaW3+WtwJjWXSHHy+dqItGxIlBu3YOFAOW0BKHkykKzFu9Q55gmO0rdmUrZhzOb
SR+SRczSwrQfginsaBnEaUC64y6pk4zrIIlpnfWB+wHuJ+zrs6OaSIFsHWbxvhmfzPEQF4WhPIhu
KW5CPal1mKTpwYxxkRGjcbNfNHiMK3xq4MfNnWiy3rIRAhQAxlQfm6B0GoCGcGg7Z+1gftgDHxNE
8uYqrhM6BwTpvL+MhTxHxVBJBLDD7N0C9DJ8Jv3YQMSHe1tsZJ9iAr9Ejdl2WqdNYFauJdWDjcgA
3xug8x7DpsiWvhQzG7qf0h0UnumaKt4V0eWARvHrQtGd0sCfxqcDa6JB74n1LR8KgtRSM4RUD8LY
s6DrJ1zrkeNuBkE6/qbHtiMecKSj0VZZnQiE1+G9KfOP3+xhHA1T80LS8XBrncuxS/wo3TwkDru7
HT0+5gsMknoBewtTyJtWs+MJd/Oxm7x0IOzdcrKoVOQOAbUTEImQodjSu5CysCe79fAFUB+eY/of
nUbhbHy0aA4EqWuns8p0Hr8MFB4qdVGz7jdwvM5sR3/O9I8mVOG+rwwGZ5zQ05vHlZb8R4mHvIIl
VjZb5xBnJIkq7LuI+GIU576KZQeU2roln2jxnfvOVERbZL4ztS2Or0bulsvLG6LVX9UjyXd4lVJz
Y2eWFT3gMgjP+Y9xzLi+Z31qrzu+v8O5N2drjYY50XINn0d0y4Tm8Z6Ya4Sz9How1tyCfltPZvpN
WKK1dvfYcoyIBHMf/ZPd+y2Rdk08Hu6idG+g3mDJCaDdp4MmwN4+zx01EKvCqebNHC4miD0f64M2
NvwGLqDbRwKa39OPTb0tVA+yzGR67nMHgGBx8o4RShEcoX12sV72K6pbdLDnbMqglXirKAi9uOfP
IUepVGeamfZk5NuU669BSe6WzkIvdVDWAzYiyQm4Fbm61v41CZEdEybSCD0DCwbzLcxIX4lvadp2
Hwm0FRy8I631lKaCL5i/IlN9W9ftzdSI3gFNB/8/sKp6f1JxRzMtVsIu8iNfyx/ZD3OisHNUm14r
mP/Xj6i0XhxNt5dnoXZhQfz4uT8hlh2BMF0tgqNkmN5mimTeldZmeYsRg+NLhQFz0aFV1jN6UviQ
PcfMb17xgFP2yqVV/hVqXefZAJJvExkZ54ryzlhAcCIa72tpAbOyVF90Y4dv986CPIDLgSgp1/ek
XgKPkOCwVw9nQBI/nYcUKRFcbUM30NCU2TWayPYsAR/YVROuFkAT6A7BbMNXau14oPYkL3pEOXb8
WR6opIR6w5cb6GamE5lhaudcbdjJIOHHMezLc/mRd+i9DkfFqvfJ+lfWjyrM9OlpnmDVxqWTCWKe
XGqjvzcHmBRRHaOEPYYt/4bNQsQevDY8/T71/2V7wNHzDM4WZ2WQEpg1kdj5etBQQOm0FKnQY/Il
cVpFGo6bmKZwn67LCz3HlSG1dEWUUisDA5JFhqGc829yloDP3S2O4qD8TWMrSRN/mObyfOpg+YD9
V66+hTzg2LVKNRiE3sykl9y+ZfH/qU1J1LE7uo/H9+itH5zq5HtF8rCaoFCpY3W36Ha9KSXIgL7u
pjezxALsd6BtohZpGUFU7ApQBGxIAzvJXh4q88unfndzbPoptsxTORe6gLJfbmzG64jxgapm+PXm
E+ulnqJwrh/1QKj9SPrZfRe1Nr+w1IrpftycbmpiCC4SAN1tfCI3SKHJcA0KXkk/N910evFfZw6W
MrWyoW2DY5HP8eKgG7MtaAZzB04UonUp30mIgNLCbD64DJPsydMtkCWglqIwvtV0rDlevUjGwqMy
cTO8IExK3/HezCLC0jZNAViy8tr0fbK0jTnFxL+Se4TiPO3fQY/soB7bOUNCsgceimHoQSuiPtpm
aKUPVwY4yCyv/WV8ra8BTixq8USBgr6zLMRylCMmzS8Mv9ejaJ37BdXlQLa1bV+Z8qp9cZvJDmr7
4C+cDBKaYfJvj2sI/Dzo7F5xm9I8PKAvWTv5e0lfJRDcNCLrE3xl14mJg0L+uKtnfDoz2wc4LqH9
xmb7BcgRhJwahzhqfG0XfLZl7V/XraHzAdzL5N20p+Vlu7kpk30JDBfdowcAqUTAS1Zn3eEmSrcB
2UFEJs7op2PWUoOOPCGdjo+5zyePyjF+v6TErIAIcGu3ticJ0vggZbQadgCYOGDPf1vCjWBcQKop
n5ksjD9MUTSPXtgWyo3C+NldBKbbHe8KRTKhFe2cWHtSbamwvJ6NcQ4eMv2jzSZHtOsOjeLJRNdC
3JP62i0NTfGOsCogU9apTH0QulHrPFKPrLuAVuowBZOmn+2X77jgAGad7gJ5Sret0vj+FdFzICjl
x5SYf2x8HwqAjdnFWa7iNSqDfXU+MK09uzWd/wRIWG6NasZVu394rREqW8PcJGFiNumWXAByh91H
WVYFtCaqa/YCKYC2GuLxfXJmgBDJBF95eL269stm/Ci1UijNqRkOPeUPgZUMqTr6TrrXMypchRbp
vHu+9/Ia2z8yfA5zHaOjZdUfp0BlYPY7CCdjKGLS/ziOOniQBXf5FGY5Ux6eMmJHSALfIJeShoa0
cMu36CJLrVyv92Np1DkW1EgBwc1y19vWzu+tAks1YsbJhlpv46x9FvlAe9Yvp1O6IOUa3N+kVRUw
PF9Z1Ood6velGvg/oxRfn3p9JC+zGN7E+/FucU7bHMkp8RrtQakiZ+hRZZgeb055J6irpaa9CMny
nQQtyRWlbYFJaCb/JL17zC0L9nsFVHqKMrbRmP7B1bmz74IGZLJBzIgG6AIY5w8y6D+px0DDsm9w
hehADnmOditF49M0ALjZPVE1GZJ8SD3k+UTiM4+8ZxZ0H19PlJjOIp2w2gAMbovw5BKlDYd/mNAL
iyQ9QH/lmQ2x52rFYfMYd8Dws4oV1DbaM/cP8ZjXYBjvH0wm8ppJUJTsrqw82UMt2WxWZmVNNxNT
rjeji3g5Vxtz9g6TZh3oZd7abo56W64V5maxCV3rn/6HyLxFpjtsvxIVdvQg2D1RaMq1dbCsWJhq
+Vu9pWGzZdD8BIGN8QDCbFmDknCf2M0PNtc3vjL/CJZg6XoBMQp4rXgLw8TFHnB3LSWHDgCJi/4m
/n22Zi465Ujtf3UgSNK0eE/1QY1jZ3TuYGUcFV5AnfdhSXl1Ik0J6MJFqOgBeQr9HaWXgPf2bZXD
CAvQqUc5Qy8IyGQlQBZe+VS0rtJu8RYQmhMfeMMzEWtYGSrI85t3NRhssbB/mMZs7z/woDFL/4wl
gRv4v1i61fcZSaTgwszsuSdaWN0daZr4bc9QuFVEG8fyhBYPq7YE1ROm3DaOLEC2dqk/Efh/V7z5
ucGybiFmiTNw+K2vB0yuNjJnh1+tcxU2wjSUnyxiWSYyRCuagUBHWjVGLVfYxDYUfT77R1CWaUBc
13OAEgeneQemYlAIb5iM6iC/1Y8fNyB5j1c5pv1vgcwyz3O5TySN7MrxxB+FPuKE7cjURtW1J1rl
lKZluke+xXNmc28ShGB/DPlEZOqFDg0WJgyi41aoE2Gv2olA0Lz7gpR/r1GU2hnVMYEmyab+FsYg
3VFU4BE0bMdjR799m9F7QTmnLo4i3Mom1sj755vJbCkntImODhgk4vAX4GySJBgOvQ2VKItTgp2X
vLPoLodjna2w/2NxUHpAUktYb9xe28QoAVDFFz7YwtvcDeMSHwRBzK3liH6dypDj2XMtosOUWIyY
WfcUtzYakLfzCg7c9vhlyYrsmwtKsgCfT6akcrFFKDYAi5y6WFfo6qxWsFjQHBpErKVDqWC+G8ow
1J4hqX8IyE+VAN3RZ3FBXGvw062zNb6RVOkhCRDUiLmnGvFgjst/PFC7d4SCLJIagwiwWNHCRUdJ
kT35+RiRaIWJlq86Lv6EXDiSW/pFXNS+Eu7Pu6gYhm1jXHZR6Tb+wZbTJ1aivCQMqTjzpFdp6p3y
D8Xo8/67DeovJlhZ2VAur7x+9NtobhmAY31cL/xTWdxMmHrnK6VngYqIFQjaTljSJpEmb49Bg/Hs
4xNjsWzoJR0NK/bd1vcRXRDHi7mNs67JOE58f9KB33Jv9JjJ43b5bynAUWVj+Sii+ozwqKpLPEPD
IZwISVi5uUoVSCPpUGST0K/oKlPQe468R39nrDLJy0u+j52nsgQes8xMN0Wy0sSN8N6lzeeRaz79
aUZnggcOBTq9/Z11X6LUTcxohawwxsrxvSOgS0B2sHr4wDe87wMEvPlzdRCAEj1holcHRy7xcyde
LuVac7Az/9RFJ9d/sTab5t/Nt/qNJl55BESQtJwz22+mmHGJ36WDIO/BjHaMWC1ebBUAgSjb1+5J
jLpDlVAkkR6o6Wu7xapIcaNUS1qj/ptda4ESTLxhIGn0TvKkLnPNB5jLuUFqbk6t+/h6SJ2SokMk
/R3zdowZPI/x6JGCG9s8vfT2bbWNCPKQ/czAH3/ztaGcSuR6KXP8gsJbjjhr/wSoDysNKHzZ8TgN
HEn9AtrZYISXrAxVtajOw4WnpXjntqzoZDbFerEfgEhFb3sWPCQcqIIsZEHpFbaQP0UnqZVW0kDu
Aq/8k+RcyWAsvdipXxX6NgFuL9hwx3jA+Y9x1BvTBEHBgc/V+dujkmkkwk0PN+Aj3YVsFhbi2un3
4FtfzGDjlO90nw1pSkoh22dUqnumTejq2G+7hQ9WuGgD1QOt6beurwQgaGjL4CusvHKIQyCLhaHs
64cW7UyrS7b9px4n3/abPvac3AJOK1J4RgtdEiTSdSG5daTlLKefKTwd/PFWrODdak/jNd15cghw
RJ+/OqqJ5xHq2lwc2ju9Zn9PuLPpZIp13tQzh3n6IN9yokNCkeJ9nm43EWpU1Phj/Kfg1mOiQ5cr
zVIR4h/Opzq65QuJ8URz46jj2MWHlIN+cENZs9Xizh2iDmhuJz13q8EyZ9M5O+5it13YubjhuT8i
w2nOcu189JW8y+l1h/Ncm8h3VP7gb00SuJ+x1MHQYds9rr/wq3Jb5zlOqRQkY7dnYPH4PUH4Ipqd
oUT5N0bLMYShMXmMtUWAIyb7tVJsOFVQUIOEXoTefpMW+QBCePy3SobRPBLQEY2sp/6qIPBQHSjs
D8H0RvmJB802XjRaw0PHsVamDHvcjaHPo1/weLkLcr0E83C+DF3ue0x4E6tNTyElyFhiZ0m0WiJa
sBvgyaqFIwt3uTpgi7tf+fMFDNGWb6j+iCQKu25cr254NqhKU+zuiQQD0B1HrgCGBqd7rQ3PjiFY
l/A+18IL2FWj9GFVZerBXfksiLc0++Hh7SmBmw6CrBglTIeLD4YwJV5ul7GGj12KIRpL6Bl/gOZ7
qOWtOh8sGNaJYJQInRxnN4Mn5VsX2jbw4sRmbjfc6BnsC16O1KXKWnpcGj168H0Ofs+rjYN7Bro8
FnMtYVTWEdJGxhXo+lXXwNGV2kcAInjJgN0gGmIIVf2GR52VTNH/77ZApq2bfjEmBp7Nfvr1THtJ
buHubSYUHZmORcDIRVmelRI3KK3W6ZshJVbMm30X1P4O8le48nwACZrWddDKT7GYB8hX0mU2Qi4y
2B6+88UyjX+noWyra0hvDU+ZJfgaeKDsxTCN94NOnTEUQ21+DbKpJ+vwUwn6ZKMfMsWzjnkzYMD6
nE6kaNtaACvyaIRriWfnd+4w0VLE1l+OmRW1IakpRJ5pxNYGSVsSCZV3lC9vlJykGot48irF/SWo
O0cIGflb7qRekF+DxGrvuRzjfAWmr374tKIV1ydWbneThhRaZPxseb5Y4Xe5Llf1k+9oTfhz1tcI
JfRPKO5d9aUXlvYiZoFLfc4q+NWQfA8CQbD4LImI9reRTKOHiyoLcpiL5t1dK7HXwnBFWB4lnsAB
8SXAkRZICu4aLvmYLpMi5kJWflTkPPprRAC5aaRVE85vi4COhHCJ6FRbxhPchsgGO535xAl2NXMF
oaOKVaJ4bgeGoHH9fLA+8ZQUMc4telXN74hXVa94YsbkniA1Ppob+1KEe+tEHirTeP7WiMhTcciM
S7mjCtRDiBADJB3HbmLiVziIYUpBi0nqV5TvZJwTyKr5FK+b/B3YbOmXMekJrYaw4ceIHyr1Cn6o
MyvkaIjSYqZjV9lnAFROxM8vxL7CUPHv4ANwFkJyzmJAXsjGirmm3IyVTyFgljvzcqlPOc4BTKCt
30U2zG/qhtQ97vTiFFZ21v6BM9woSbhJG7ykeNv2b2bn/HxZ1T8EUDFPFZ00f4a5e91DUHXJCjIQ
GM4aeQNHw/YFq8w/mYWKKiiL3DmTluMc2nRXuN85huepMo1ywaQAhonOxtwTlb4Wzva47eHFdpYh
JbgnOh2BZkns6RmAWGHrdvOUBBwomLr4IHIOaGPZ2ZMNMD8y7lO+L33+YS+Yrz/Pjaj8fBNKW8Da
0wefMPpRbEEXaWxLRFLQr6RFP47bbyNaiv69kPuoLtGlz/SnPMyGJdjVO0dgNl5SeOvdxesPldhl
ct64zo3PlHOejj09uirZDHTLJvlwTA3aY8XAuaZEVvF9kMX0rdDzbU02+DWzaYB3f0zyWUi1j+fq
qK9u/M3rQ8blFCckC3l5hG0POvxsTXCoFSZnTyrBloEha6+iOYyB5AowWkgXUphdKptwErnsPbLc
fvOIA4KYxiBS68cDeUEVDlrsJ2AekXF/jC+KONL2FjGd3OliwlVw9/URJejzyiJPF5jxLI6rJax9
Z1Xm0h6RudrImHmJLQtGSW6gK398iSUQ5rsaPJYMlcmEXf5P+VgCHCbjmNFk38UjvjlwwrqXuH+F
B6XumQxcQqWNs4Tk9vjaqsApkZAkPtvisAkTeSVqYPKXsqywLGYhM7Q5A+X1UWu0eGhzzJ/v3iFA
D2XiHUjiFJcIngo/60ZmsmIVg7OZihW3VTdwPK0BIIeHZa5cPCoF0QtkDryR6NC7kFGWIo8thtVH
f5AiRqqxPOL/20fqkgNaqkU4TdNcRNYfArcMyAvTZy2KUa+oYWTrYOC1VHCY9TIq4TE64Ns293GT
5L209dx25t3QQX8OBD2lOyAU1J/g8L88XL9Rr0+I8A3rchDpBD0rN+Of/cLUD6mKuZctZKSuUEpC
+v+3NVTBaxhdhZ9osLZwNpL2rtxZTh2GkIsf/wqiImbQg9ptvB2+hPVa76TxYH8o/yOGqMVQF7Xm
ig6Y25tTx++rX4zenXVDPC/EeQFfd6Q3BkTLJk8WxrOLYtAMXsvYNLrqKf89DxppBivnI4qF0zIg
ElabpPHaFCrKjphy9cDvGnfgGMbl03EFKh9oAKmKyxZ0AqdJzWRhjdTCODaKISXFN8BmXTYbErQN
SS/RojDwhMEuXy6UtV+voG3y2G6ZKQdUwCTeFmte2KrBeSjAcgAalA7WNciSgTcytPaQvZUQ/G7R
W2/MWHIb7nmXGN5ZJzgXxtQp7/BSQj28J0d5taKSh/jAYVfgfrG/vdj+9af5upqwssCZkuMkt8qo
xrVYoY0nDCVOBH73S81eXncQfXwM4GKSWQ8ZfuUgF/5N4jhg4f/WjR9mRUzr/70kmS8SAF/+IMmx
NJu3F/dOq5jJksjbvWxqVHfPMXgu4UT6N2V2uHAje6/W7YG8NtZnD23VWJDabPuYowhPq3hPs49g
qn1sli3DLRw1WV0MCjQe/2Asj4zufx3Z7CGOyddglJbLPgwHNXFLWw36zx8i6cuhr2cBl72kVvjs
0Y5CWG6VAUCJZ+kQlBubrwSkExSH3bVEJOsTAUD9trUFy0JTcSt0cggVmOTpxvIrx+1v+CGg2zB/
wFeqO/yZpLHtI2b0duFIDoR2cLlcFugZnZNWmcjeByZtKdyxdEoiFy9QY9eyt2A6v31vhx1HStr7
xkGLidO1z/ZLzLkGNUT8SV+POdv1bv+suD4/OkripwdK7K3WHyVGiPrJQsl74owusR76PUGGUOga
pUSUDb0F6J3hZn5jq2Dgi7Hb/53vVW4L4efaNGafU1u8AnyYBPzY3dfeB7hBKnsfZ4yaw/tL71WH
zgpYrPPvZwe6VdXiPWgSYb9CCqOn33FYUMGneiXIV2Ag/5xyvyHxxf8Y53QcQ0IhUhMBoW36Bh0h
9myhSCm+UpeNp/yFFcTBIuErzhfSckfgulYnLWlirsO4cIbt1O012apLSQlvCUo6BF6vTL7v3sCY
d0dRila1iXXiWIcCztDetQKswioBAj8BuwSZFJjUNhv2Hszhi15o8zCXn9RjgnrHPeUb68+h+glL
m905mLIlbUg1KHsEQDzn2g9zY8C1pKpNGi3NnfJOYQGPjItFOG6ivhpTgGVMm3exi2TpmUY4/YBY
+f8lgpL9TGzbHK9jmNEP3lsmer/u+vNnBnIfgcOgv0y3PFOTb3r/a3FVBDVwjVVgWd6Lk50wNXgj
DrBPoWHCpLcuM4uxFUBzRcs3hM6aZVBY0CBbhdYwTJqcJZ8jxcn1zKbhlQy/BVwF9QGsjCjGcmXA
Y7l32w8YWIeb0hOPxv/zDO4x1HQAtl7wa5blltOEtQuMVyuuq8V8XYjMnS0KHNHu7eC2OjnbtsLC
ufSRhUoaCtFh7hAL/vtOVOnwmt9jhrJYuNpmHtfCEComIo/ZdkgJTDYTpCZcEzv2sQojJeQIWvRK
WdFX8g538O6iv9LYzDADc8tv+Id5wFI/p78KaJPllAMnb++8XZHHCcvhwaN1NT5HqF4nhB65b2bA
DX8aIyc+nmvWLGtv5QciWgPNIg85ORutsxaSBspnapl5Hi3+es577RZsaxaDCeb5FJP8iGw+tbdq
6WtePrTibGravt8e86DcEFxGsDUyUdm2gCKH8o1ZEWZ0kBJUzJ1kfKONfZExih5LojGkBnlGvKdQ
CSh5QBzpT0/hGrTmPqJZHQDWBFFJvQjUBtVuQ92HVGIpBb9Mc0BSVjuZkP2o0PMO74P2JZSEECmP
oOJMnWvZvhbrc3f4Yl7780X4QvTdZ+3v5I7ZQ38DO+uhndCtM4HPwxL+e5krRNzMMJXeZ3y6CddW
E4wOLSCj3NEs/dG/yYPRX5m3bseCVFI8oX8lYfMAuFndHN1CQ27bk4ra/6w/sEzEGNRoZeyrvSKE
Ib+oCLG8Ra0NFC1WjO4rsDAEgq9hadHhJ8r0/8TLDtlOQBA8z9pAjKg70arBLviiHEpyGvvTJnA/
q9dMNW5gePik9l6C4nXiW9/WyzK6SsE285L3EdKgxlwIm8oe8clNim/7wJOSt6E8LY7lbqZej5jx
gr0uG/l0N8yZU9IL6qmz3ZcpsHvPfcLGcMet+ydnVvNfaQZxGTjJ2VJQ3FrKlt+RJGYNSGbrQEBr
+px9lM0gN++HbVtXBkoCfc6F8tXOMKO7saOO4n70iUqq3FTVf4JzKopJ2QxW1nhyHh1IOcCX4HKp
Z/cVDnYBIxNKM/u7yKq3cbXKz65j2cKvUA+6DIyCNgp+XtkvDoslrnmNKyH/AAfZyMcksTEYe+ad
toDutqqx4T8yGg/hE3TaYMidE2EH9egPaKVEWRUEfiyB03CRMELLKZHUJWD87klFYJPxiF5h05zi
gXrM9sOnpNtArp8X7zLTu2fti+GKyOa++e3blYDcP0l912poCoVjmGymMJN3YBHo7f20CkUz8WEw
ELzWVVXKijyq74EvSLDMwp+mdsdE0ejmBSUGn3rcCH6tr5M=
`protect end_protected
