--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
cERSAH/XbqY9YQwyVdKS3LM1IpMFilC+GqK8D63UiO1vW9Knmu6MSgJgkFTVn7YRdvlSm+gSf1e5
5Oc9v2ZdkGrYFnxBaBNXh3zaih/Z6Dq0ekUmAs8mdeGWwL4ubTJKAygSF+Mz8WUaJgAI/3XT0ysa
i1wiUbOVYlVVU28A7yEenqSufY1V0UyTYuZ/VSKIGvKXsO4LiqqVoJjDqsxnPBPKfV5oluHVhoXo
pwXANIGKbmKPWpnJKiCBjwFJbHw9U/DzULMVKC0XNIknHSzP2pycBYNm9byhOgTgeyajJ9pCNQF+
hYHK3CgqVdFUcCjTgacQLWIAtbjYSebWx5U3Mg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="eFJdpf9VcvO9tI50IyiSyKv6gjtSfxJBIZLsbwZBltY="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
n4ng4/2WYLkWZjxjN7OWioaTQl27QVqE8pvFGT3+qWbT/J5TKSaBUQByM0QYLhtUWuJc4IZZT6BU
ZCCjTeuS3C1BmiislJnAxY3qxFPzIdOh81tBqd0fQdzjwa+3c7aNRr9gQjqYXSiEkPS3UF3MyyLy
Z1PPIO+rvvPrY2FuFw1twzyrXBVoaE765RGsJFiShFaDSC51ndjZ5/Nb/pO3QAVpx3ATC+56mkz9
BrTtKAsMiwM7/OK+/CRxZ+RkHw9dJ2MnOT3qHA3crThS8dY4wtV8AxrN18rEF9WS5NplN0BE9eof
aC0nR+myWwe6pbfF8KSq6e5FFJOXJaDLhwhoPw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="or+6oG++zrsY8kcVN53MncIjZVyLwCBCKXwVNlf+8pk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6608)
`protect data_block
Wr4Gw2yxtmRuQiJgdIOXkpayNgF7JUxUHnGsv966jdXnUqiZDXWtUvHKkXOffCey2fVrOMntw3tl
xLWwFGJ12r8Bevi/LYpfiNmbKUHz1eUE8kseiP2nP5tdPvoisCzPkc1G2oK0RYtizVaMImi8fjNq
EHMDmk9WQIndWQalBAQrSESBpM44ga3kzVtfpdw8deq5VwhAAdfW3sm/qs8ee5FlJ7KZp4gO4TOM
xLtyC0MnNtDICNRdEAvmTXo7nk5NENDWsXnKuwckaKwqNqpybt6hrwjeV7PBMdC+BiDrzd3EApmj
WL04lD7A6nEO9UJGgAytyKjOiX7/O9FDkTwzaopOhoG9MbtD0jgr9vos1vkgTg62kpsI8w5jO5XB
blbBa1W2GIti599qARY+BKYUGsLkJn3vSGLoIZLyqWb6Mv+rccMHBICwUkAqtr21tZc2bOEWWtkc
SMjIJCNjkcXcEqJi1vd6TvYdpSBheTxiVFS3sszMeVdkGWCS8MfzeLhcgJRWJ80M95CWdHKbDJAk
pj0X2Hpti7HHrJYURi/JJKAMA1U3Qcq5CSHJyuLaFajdTglQoOT2DP0QT767hAIC2dbBmzRekS8j
QN17+IOXUTyEdhXlBfk677kD8O2nT0tlqAkXdUxG0P/Iz+kLO0uIt6aVMaf9BCp9amW+gjmmbFlV
hW3k+7d5UjBdEgH5qc9LGAaRmmKapQhBOZgzH6FoEUroRyNte/QmKivAWk5NEBMnDjB+QWu3VEiW
pIkTpD6Tdz3thIrrOwDWMXKwJq8vZnwg8cSs+xYgUEs81MjL+DWcCjZsdlcnVBtZAQO4pVNMGtpA
yoxXacpcMrRoCmHGrnhUdcoQbk97wRutnjpKoMlFU2ciCcOXQ5UNT5nOfVrNZN/jNCDWzVq2AaEP
6wnifSEaPqEegBRz3xb+2lYRCSC+Ba9qhy4ne+EW3My1eC77O8I9HRRHh1oSEfDMG9L6mstJz1E2
du/xXQiCuelxnFkb2s0Ra0BizKvSYe5L7WwcMfrhqIGiDdprC+nNzGW3IpaAWPetmtVbB5x757DC
w2m5x4zEBQ/KmATm/nDO9554uoDGPkpets0bOC2nRQdC2F00MpW6uXeX30iFMzOr64KvmQ8iq/HR
OXCBZsM6/kGbP5VZZFkO8LH0jz139ML53d9f/rS53mUIjShlZrt2fH7kVJTHEzGC05rMBJClY/nn
oMjUajCRIMXEXhk1/yGrjrRJbZQ5M5nMoCPz3KoiU8jQHGzD+itaEnjqRCI8dYPbrt6fSM++ZYmA
kwUUcI5oqDoEXndD/+LBIRULz061+ll2LM5BXjte+vY+LRCVE/Sx0N3fxfpkE7P7NWMQs01b/M7Z
yEOBoiCibS8xTBKza0JyZZ5v6DByGS37JTX8eeYNRE6vOWL9O9RNExuehZxdvdtS+pkXiOhG1WwC
276PuHWDijO/JJa7A1pnkxNtvq/tU0s9h2Ev3sSxDJWsjRiY5LiVKOMbhUsbyIXqJCKeO2lCP850
O70f2sXwOjD8JRJHo7MPurSRaUsKz75dUZVzPynRH9ajuUPUdX3OVZJe0Rx17vhCTscIg7zj08X9
nU2ZPmedcnP5alSn5sjldz+eO61Vwn+B+tqjKz1UCYqMyMWLMUtdSz+1KSGUMsL+3nyBjuY30/GF
Dd61UFgCv4FWPh2iRxS4blaW8zbbNZqt/R7M2R3IfElY3HcQqOO3fRsbIQBpRasTLXt0dZhULLOO
05adeWKnCYzn+Bwm0pCtsfv5Ht0LsgBob2F42hVrLyj/bJM7QTwGlyklVhPh3+VKFUAvCtneo6uE
//NTr/yfDwIaOJcaLN0RpKtrqZKvJtghm8XsuqWxcJ5FGComoFyT+YymitQFZLngCuLsuU+ZgZX1
SAaJnDUP0ZFLmiHmliKkccBdEC9yiJPdz4RZVPM1IAEghuB1NPSMD0+4clXsacUwtQTymLDUNPW9
n1M/BVT1AaEK8YDmJmWOeX0PFqe+v6FNQlqsI4dMBPUtPyhqmnOeaUBoQ9MOBgiFh6tz9dsSnb+b
QCJu9mTXtxbOwJD+IkFiWMapqqZNIUFYkyNatqsb5CQtlRUu2i+V8hwP3kyuV5/ZXYwYLjf0D81U
d3j/vb++IG3jlr3uhLQivOaGGuHq7ZQcT5ta+vR9uikRyqhyCcpzrtRlCgNjR+JJUuNZdSUvZxSj
C1Y9vXwtnEKuxtFrmWGIB75ttHb99DOFK4uh/a76mTAMk5i7sw282UkwbXnLqiYh0j53p+RQ/CJB
BTq3qmCUOZDmtczdA6uGreEYnJWDA/roCv/PnT514FLNg+OtLM8+z+DjqagIcIcuOySolqWAZF06
hSir3Jy1KztSE/+6czy66HhG3O/C6RsncwO1HmG4EnyzC9B3LFUujCeT/f9CguXKeMVXrVxOIahI
ExtCQAtHMMhCPz9/Zh/5piiBsGBW79S5qzbTtiUXhsufX1Hy6JLB2PnKvaZscg+t9InXYI3RwU5P
OXUBvpyYk1eVeDNE7tMGPxdBq0Ac1jyPpQy6EUoQzXVvuTd1mX0RJDJJI7KMXzPTfNqsg5/ccouA
ua4VmImooW9QPL0WX8bkZ53pyTiX3YdDC60kiEkT5zQS1eGK2AgXEduPiNE6afWXqTw1vLvTerhx
NgVSWqp+lYETSP4tlpnjZut7edDh0dDUMRRVEI+cNK7p1VOApReps3KLztFOpQKU6F7QkuhgS0f+
caiJr1oidhhHaXLxXd4wTMmKhGBe59HHb/aUT4K/uMgzjvLFqvoo0R/AeKfZ/lFgOavV+OYjTwgl
sVsW/0Y0rMRWYGShnfr20bYkXgXasfAIGJLuZ2EEdL2gDD1QBCTG/aAP8y1dgKTbyd9zlmhA1ZDb
QldG/wjtSjbWxYAE2AABpaDFS5Ppznwnii/1ddxCe8TSZp160xgWBWwloI58h6V776Dhft4RqERY
AdStTnGfeAopL7YvNicQD16paOkaRcMLOznULBpmFXmczsmTWEJG2Lnhx7GtWKOmU6AvvOwuMteJ
dOaq2gV749+GTh8OOsRdwqVJrLTYalpFwhExzUqR6OnR34+uqzmNe9s36Y1TXtauFGfv3NTR6tEh
6XAVtgJSTbSavlu0IAG1J4iEDtbmyaUZVNnzgD6Omz86Ykzpz9up97/xs3i93fJ97cInTpR4VCiB
n78zuf4ttipciqc/So6tmh3uJiC5MysRWfsdHBy8+6Lj42luETlli5t2A4T/E572cv91Ibdi6WzF
n77Zqe/NuA8cvaAp/wsFsXVfnErhUzAlrSVpYHOLwbk3GsMavDr9GY3wpxcCNudycYSRxyPrMcQT
PWzun/+70ltiHztFEMni3MlSPeDi9KddOZ/6HR2YuKipVOBkKMB63WW8TUt0VUMCmJkW+RlZCwGv
HZyDCHxG0P/19NPX6FciU8dLd2nrN30DjfrFUy0rh3nCT5dkwaOeUsahMyeD0cFr3/A19LWQDf/8
JcM6hOaLmWPYJhcoNQj1Qxe59bjX8KRDG02DzWU4pKM0166sigjniv/u+NF5kFSlE9cX4dkJK9pc
DOfuEal1hz61cB6iYj6TJflwcMEDchve2ItwVH+Vylixfa8eTusSVZBb/P2Nfsnr3KfXNC/rLnNK
yC/wFGAmHLsKr956T7i5x+oIjhrT6q+xwGBC5YSKdSVT7c7qzqgnFyk1yF006U5MbUTyYsvouVie
UdxZS6+EYc3o4GiG5EENdTgWUsp9RwpwDaRKgpvwMB97M4Me50QcOKtVhnL3E+7BFknblAfgxWNO
nS42NCl7ANRDq3na8z/bh4Htv4D+OPJInzL2rJcl6bFMWPV+K+H5cMRuROZGQL3mnF6U1u1/sHc3
AJElZEGzF+j7BCMEX5HQ/Skql3AGpoCQH3N3PQAQLwxsfhb9IN0VOQBaMgheBW1u3vHI1Ryoak31
rtT4akt58ItJ2Tsnprjz2a43oSDzMes+K/PytDiwuxC3R2OjVF8Ad7jvaU17tgoPhz79CSUhfBOo
wTKO0W/zEyGjnZeknGgCflPxhKGiO3lhA//8PUUcSG2Ij26Lu53kiJyLa7QAeiisZKtOKNZcv2UW
SPb/LhZ3EioF69D35PC4VCkUwl0atkoTw+9O3v/AiKJ61fqV2w+BEF7EeX/1cJo6/vfmTkugGrPW
3fyDZrSSPZCgCvIIpqdVtjBMerdPaKW4vdlZUDSx9RqHU1wNOKkQbrJdMWPbrnTyHWWCLiKRgpN7
ZwOuyuGK+pf6zRNHDTJUTTlB0NecKYA+fBa/GyI9qwZpDksvnDE7cRRkmnrtTJl6oM2VzFaEMVD9
sd659qMddAFQaPJPjKXvsoukU+dgod8cqemYMFfGsY4Vr9S2AYgT/PhDfa+g6SvFtR/YVEHF3pB1
ql7WpziwpfcaIpC6jNqA8w12NO+HE6BQLdYSnlwxPHk7uNP/gIiyFchbd8hiFsdkQIMWeaPJSEu7
r1+aCKg9rvoLgziz/qSOAqJmD99Pb/ydgqtuYjsuyKXyB/GbkfbnhSHSeHQFX/Vu+kbDPMuLCP+S
CWOo1lo6THcKBFLhawveIKE5ORgHGJY6JbUlGxMM4W8ihTkE7ie3dsJTfn+IAsUT7dcExp4jJndx
hsHqVi9zz+i4nhNXS9Y/kkdbVQctD5hkfU4fi/+X7Q6JItaskLtqEtjumbqj7akMPfVCSgSaOmx8
pqdku278xIC1mLq2kOtaQWiR/0vXdvZJtNGJAKY81tjvSJSOP2/AXg3Eddd00Ji0OdJAIYloG69G
lDFW/rf7MkW4KEFhWzm0FC0PWr4SvWMOcNeZBtkZLEp/Rflg97kfpt0GqaP9P8IkHJFJwklKoRoe
bxkulaBGIisGF332LSuPfpIF47yjx4ucH7xONHIxiU5ajSr1F572F3rtRxo0a89K72+DVdaYiYrV
IrwoNJrn0TAjkJujREcoIfJMH0SW+utqsi7tws8H/evVxUTuNscmbGoYu3kaW1jUy5Uxpowfw8rH
DTJ4MGhp2FXLxrCt3bIZsGBCSeLm4nXc/1410498l4TGCtQs0gnamlWYSYqY+O34gKlP9rEHFyd4
0iD5ZlYuaM5XYWOb5G5F7nxuIGuqQ/lorx1JVxCvZcFyqMXelRWWMHg4O7jOD2F8yXqE2tvKJWhl
MAAB17Rl1A6Ws18N1mt60zYEqlxvXEfUCaKWT1gVhmF4h22pK5XNeopPn9Q28okDIgRoteEvMl09
eovJ5l3AaIlYAkXba/hd/hVHWsTneGtE3zdE9PqOvd1YRMeT5Vgl8BZi2AXtLM9v20zRuQkEBm9N
2l+rs4gw8VSl280Lo9YXC14hPjX8SRO5VNAbBFLXQqx3y/VRXPHjH2gfemj7orkdDynhH+5hWiC+
TFfruqXd4uWVs4Nkw1twelXYCQLABWnsQOGLhKiq59LAaTJhoE09qA+wHFIR3M7y/ipQnJ1DIO7r
SJygNtfflq9DLJ3oQma41BLrQ4AOINamfpmJ5FKjx9l2TtGkTOPQUPVNCjiGMQ1eiEe4yPB2VnxA
NEZHc2ut4nH9f2JV4j8T+rrjD6ZIEBHbdBqaAL4ug07WymGliOmJMVszoAm2/TU5D47ZyYpRsrdI
TbE8GE417E7n50NoIwRXOi3Mx1Z5w4V/w5lYueJ0aqdGtt403E0UEdLBdRxS/0OvqmJdkOKg47C7
f27U2mn6y4JiyR46ozF2S1O70oE7biYBbxnvyCXFOw6tgH0F6hgV/dwzmmQIacuETfzbW8Kt2l73
/h/MfExVDb8BnUWdijT5aNWd5M6ylawAcc17onmgQCGDBP7/fu685v6qsgP01/RGPTUDZhW2qs2g
mpE0C+VbqRCNV0WtdsZUMbnSuhiUAIpCYnONbf6OrpNaCOQ8biYLjSciJ7x1/HDyKG3jUTJ/kpiJ
QxIvySndK+++A7opA4ryt0BjYauXIpEzSwOtOHbTD5BHj8HNEaBYBZn/RkRUwgnyZoSMkhVLukZG
A6a/LjTVwzzZkmvb+r8BSTSeHMmouzHGVN5lpZmmGy2Z4bcUxzQamvwJhcKSG1ZRm/R669CEH2cN
6O+JliMi1ZcXD7Ndk6TwSSHENcBH2COzf22IwJsYKJRHA1I54tpIxXERGRmUgUBJp3spf3zxw20i
w5sNH5+cxohruxg/Sz0bjTB19tQFQB+N6QQjmDCNei/40hTjv/Ym/bJCh6O1Djax386vTO85mLNw
mJ3NCoH/Tk5PlyccgAwWREnoL1eMNRLFcA8CPcZfgUlYAoq3RjADa+RLl7W3tz825+DolJgLvb3p
DkbIvBhmG2Sq6ltjA1GtFkTgSvLa+Zvh0Q5P/b5WuJVXg9pXxNb+7LSLLMsvcDlMvBa+JBFVptZK
aISkIBxP22vj0XBTHbgeefYDdwCvNiMKNX6QlhVOdXBf3d92fDZxl2EHrhFYf3Pa9ooRHhXu9gCV
9t5f8eiSCjY2g8VTxEnllVyEEA08Ab3i83kcWxeMrFS6mDahSC33+fMk/71J4P4m27Xi8Ai9br6F
HvUK4TcVtFBFAD5enkcHnXlituMkf5JhoiiC3uYZA+SZJKVT4iTXG6g7QOp13CVclRP9yWCtNC4t
cCupXMZxcOk4n8YFIaN/qemLqlrEcFsddTGJtR4vHLBwqgFgfuLaAEtnUnVafhPeazCdYvdo0yKL
1WfhtS0gdW5uX7S8RladgD9i/Cvd9nmDfAsz912h0aIRBoba4tGTq8nHDAg8jj/Lb8AAu5ncWd/F
5xFenMfg1NCadP7HNpc73Cx4K9Z+JxmRhJRGDUipb2X6Zy5fhKSR94F900qmXaQjmKq2w4ttUCYP
Z/C511Vc6J9gST1MmXXuxS+YkhLY41GaKnEdKH4QZPkLGJ450JtEOzweKGVUiH3cbBzgaTAGP7Z1
NHKyYFXd90FjEEIcIqq8C0KLhPMKm4grv9LSvdLcvAV9SNJW1n0xI0rB8o3FMhcB17BC0SppEOuX
LkFxqYFKnZUxCWFWX5zHxM061kJapG1qN8VT+EvYSsn6tRAAMm6WZGad5leE4ef/+dpJXVrafwC9
LOvisVf90F0Z8Xis4kqe0M5xClb0Cjh8okV8RFy0S/Qq+54IZSzoJpBCtjL+e1/Rd32r8nedbG6r
NDlOJCi3er60sln9u2ebFfRilAu1zQADssy8jDaIbZvtHIlhmWfaxtoDgDqBsjtYOzYm+kG7ipFU
EmLBursOJFE2Jyrqamtawtqnvc6cyLdUSzdK8V9YpkERgiyIruVrMjoSXSBOPAUDj/7G6sEQtuSN
aPU3xYBxmCezfBOTEP8P7tiEagtxoqMAmuREdD2RU86JdTyAUJRJAokkhyibkRYaoZfbTssRX+ib
8JU9TnBaEA0YJOvDYD7chA9H3T1pcyTF8hODrFS2r0PSdhudmrg0We/tDLQozcY2XfeccbtY2nZT
umfsNvHYjsaytncC5K4Bq+1MX56RGV3xHDDnoYjbkNJyiYVOZaOAoLVRQ1MuZYEM226mg3mS1pQ5
bExts1/55LKLKNR9GEUWAUkPz1eDugFAiX/OhfoaljnTgAWngNUALZatyodpQeFfr614vRNswvy/
SoIQyITQd3Np3wPwdbY/N0/KczkrdzbIUXzitHDO2lIXmxpNtVzCz9ILNC3XxVRyoxLaG5XTGbJq
ddBT8acaI6dOq42tPRZyqU9tcUvx9ekihuixQ1GuvnzlZpIm9IjuBaZ+rlDdDrynYeCTGzOvlLbM
P6lHmNy3GC7KdiJlQGeASSYu8bMmcgJ1EOvyU6Soix9VoowkUtAsLa/KJEi/noHxs6PcZa5B1ibt
k/XE8p8Br/uUfk/Do+HY+HEoAJvDhduwAFJHqFVzJcmj/k0VI0IYWnVa8ID+0FlZRhY/s9mM/ZPx
H7/sYD7y5vN+ouB97tj/qSO0nn32xFYLhQxNge+y2QZK6dCnicmqmCkoJBvpZND5aL/ODwmqd7Y+
kTeqw70MFEMKpkSo0RKfIDgZJmiuEFbgxomc5SNyhTDtvXDPiG4nhgeZSO9oIyfzZVuofIQfXH1f
CcfVJKvU9JLpp55QOvxCjIRcU6or7ef3yMjrnY1+JcjRkZRNDls+v+RyRqy+K/kCxJOvGrw0DZDR
klo/te0uN3hk2ZxTusatj2sPX467x1iaRxycdW7PDpRkdZdLIQnrM7T7MLeGy7zswTBS7JdiN+eU
PgMOdAsdsa3EtsMD5RkiSjJHnJ+apPYKHAYDXimVFl1VGkloqb4OEOoorBGki3rZt8FOt1CjZ9XJ
w8K0PllaiGQS56uqP99Of4kaI/0LlHMBcql5Vo7S0may855kACIEkVUb5O6DlwSU+K9Rpkrgtq5n
usbY0AnX9HYohXMz1o2aBTGSOfoqypo3AWrMgKLw2up5LC+aixs6PhCqW/XhQygayI/JwsxJK7cl
MDlU3ZH5sv9N7DpoU38Mnc7V1kNDMJ9inAwi+k9DS3bPgo2SCx32YCyIA3K4saHFgwAhFMgqasDL
qkzeq3+P3fgJa94QMrDY6mZBk/f7UyMFSFek/EHg3s3II16WzpKLz+GetzsojVgbRLNgr0IiffMB
HIKkR6R9jrQPfq0yATlC4LwyWZABjZTd/uwNmzlWhnIxgnKT1pObqtSjcblDlWUNbRtreyzK8oGb
ByjDB+Mg5jEOWV1Ktfyph0WOPGlfoqEfInoam2rNHNLGRcqAeC1JmOHH6WAt4dDZ4tcJjWGH6keu
u04SzqX1QNJEPBc9Yvq/JDsQNyBC5zBMI1LDfd1oyJSIosM+bE+3JB6BliBXDPSFYu4gcBw=
`protect end_protected
