--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
ba4XuPYKkbnQXMJH61RDWA+aPYdVRzQbnvPZVsISht5Wp0NCGEKhkiEudiA7bq8oPMCxoJqKp9b/
JMyS0PD5Gu3WbBtHrVpKyZuuGiHUsfvyCCfUAVPNxs17VMGOmHApXU3iAgVueEi9WybcHlNT4F1k
HXAU+8SfGq2kBu9h+useo5zaI3vhK155PpkdNKGsBS31Ge6qgRqiXs0TSoApL1+XpCtC8wdbz+be
f1qkzHn1lVTWS9sbpSMZZn/ZkB7Fa4IrFlWfnCoy76bTSRBPf89mzYyEP2sLbZygyyUFcYOB1lrX
UxRly0ZBpd9OkYVHw3eSlDdoPMrtLnfkwfB43A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="AzvIXimFALe5OER4cVrq34B7/31icvkVSeULEKfxrTc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
VeRXF/o1yjwnxfXHysuDs/whinuR4UL5y2csBIgpKODNCPaxPTtQCyOMirZ9bF+j9I3RpBxcqjKW
V4jskBSquEQNiQ8W6j6IYmE6OrvDeQeWDyH04P0nNHoEmxyD0Z1yg6FkOhm89FV6xuu5p+Znh8c2
kBHzYz+B5bkBGEvB8dFUyg7ZmFS4OJABeOlBCYTAgGsbTI1/J6my3q+fyAULTGw5eVe4LIyUim9n
dtRrKvSU9f+UFJMq1ap3SOWRCdSpS+bs0fM6gjXbLHlKRfZUNlj/Z7h+puj63kH9Pv7Wi9qq5duM
ENG1lYrH7pHaoDolYWHjfhymYBSauTUxzCgMPg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="WHDif9cffbIm0USNOvg66GayPbbFP5ywK4oigTMAASc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3152)
`protect data_block
f29XzMrcaqj/eygE95Xax/SSsn5E5fXublkwLSaLqj/mxlGCUbI8BOe9Nk7WjQEjISd54u6lA1XE
jiZUuzvLjFjU9+v15oF/DJHBZ8v24xKFJlRWpkGiOttzDJ/MNP5x0mcMeBPYociI2sKvJIrxMWpy
29vG1MT+n68DlyDQIWfMuIoplRbn5XDp6mUHGi+OSJkhkG+G2/29Tb/PKzFFbwjpQWo6o2qT5tY1
tn5uG6YwT+/3I4Yh90poIdNzdL+XawBXabD2aDfQ6fKGA8KFOyCCyhnbTrq7TuzkQf0fsHvcGcHu
FP6msUOrJF7pBmO48P3A/IU5UKabX+0wNYfOMyVUmGZKOYmRpSplgXo4wvqP3ICivn8DGFqyNIMy
SH9NVBRSbxl/910vxWjkEC3jBJ3BLx/7RN9we4Oaf2i/apVfM8UELToqevIKyTbJhOYIz9tzCYb4
ABfUMWuSs/YMuC9AS5wqSTMo29FVpivYs9aivydY3ROE2OOaRwSoDl8Yh6AkmS7gX3+1ZOcX+nSu
DLHImS7uCVWLbsiMpcnIGgK/cZhvcq+EdrEEYDSCFToNzMI7b8GbVtoQYjT67x2GuQccRTrtQFa5
5BAdJ0si0DPrtA20d941rdBKa3ytutJq5kWHOY9qqGJ7yTzgUi2TooFSqj6N0pa0ukjXkvoKFHUN
hz6FVFXD6odHCmzhWPzbqo0AYFcmLwkvx0xCG5qYNvbUU0H+IGrq1HmJ67yL9A5lc6yFjAm6WYym
rbKTcyC5NzhaDNNrdOVSqxrGhh/avbbSPZ4NOIkJ3PN0Rpzc68dMJWK0rUR3583gcCfyKO2pe7VT
DVO71Uc5cywtYSBeacJG751BFbDTI9vDhIt/VFr2vR85P0tLrzlpTSUvB9CacIgGE+s/n2dRQuhV
JPBLHlyqQJIzD47QGJ9A4HS1yog1w3wJyqSHr+66Ux9aJpbZrE6pmfkTOOCLV1qU926c/8FFxVdP
IlRvvaWdEgBcyD53MEZyU/U47D4Jg76QF8U77IVjL0LYOakqQsH1uKIJFQZhMcPjIDquU3f69QrY
0VNGVbDcQ+WM8IoFijCSxJ7Dat6K+2tjlE2RHwGGSrCleL/o+0JiRVpR8FybTRtEgxLVK0pcABWp
gILUbHFrsIa9HvdHRFxCK4jjkWTbVut1V+jWZ2bVkosYa/fE/Ucv2eARUn2j8louuHbCG3Ds/3Li
etvBKuawqs/af5tQgRYZNXeGx9OaTIccWAgSBRiA4ydIAm2+VEC7u5mKABcMuVplWMs8H7WZDNC1
ICn/wvF6eLo0ofJh0zGwqENNq676YXs287T/R8lJW/rR5eauWia7/wxqKUIIyKsHrH4fVDDDEJOp
MAtDkBFQasNPp30sN6KtGADAn4rbUGwbrv37wkTxMnZ7eje51gig+PioeGqBix2OBm6Hv0gcnc7R
uMEEGgcERZITXaNLV5kcm1vmxQJFOEm4yfRL/6m69GA6td26C/DpQftQ4tQih49v/shMhha0GkqV
CkXgcNl/4dp9EloMVu1qwDlIc7xwNDG4H1JHnvnMfTr1Ci2hzmvRurOQU02/5kpFaro6sarMHzDs
YS2LBlATtGz5DWWaIyMqTupOF2QzgFwApBX7p8R3xf5qHnV8IxUioyiUzW9UJcZh9cBsR4Qpr6+1
tMsIBvSgvemDW8wBVp7tW6d1FSi6oZE7l1xYowTtGLfcYqPvk9okW8TQ10IVQ5KA8lv1sOMVtJu1
PfwiEioOHOkre4uClQihURcAwOdocgN0Vmr3dA6m9BymnpknrqvDHY0pLiSF/QC3o/425S6eOjsv
2Vf3m/UCJTwi37WmkDQUQsgBDlNuEBxInrv8bsH+59KXi66TZ4PV5ZRUe3pCA8ibTRYoPWht9TGe
TB9uVerOEuDI+slEzWekeDT50dnmhOh/g7YIdKY64Vx5TsJ651BB7kvvT4Dt/iMGFY7ZIFQYVfPQ
qe0Eqp0wTQn7ga+EwJk/ukbEL1pMF0yPzL4yhe6JU1jTe8lL6kuxSc/LboFj1rPpkbh5WnEeqQxk
PciDknfpefhNbiLDM7PLSduUJldNcAflzPO/8SuRppn0hyx+4rNLmFzgHvWdfy9f2qLH4C9ReTXU
CfMi1nP6OqWspnzHJFOJKb7Fv71MxqbR8u4Tpju+hM1Gml7xMiAkMBFGlSTya2SX+81pNvaO9LQi
GwMLj48H+2ldu5CzTOYd/iRTpEHQnib2vrBX+CGjutcU8LvHrGQ661JgDtIdcx5UV/8yI2Uw1X6O
IdZkNBHceXvZr1lFRxHWBHdq6j8CIOdGpJlLf4q/2LsQbOvAGgfhe1yAtcdRxIi9ex7qLVgZDe/M
tN4VXRMjNo64KNhOtxD+1psihH+OxYraNgUxVRQaqAK9jYZWy6EMA+uo0dyl6nqahFapkjBmmHFb
ABQWY2hzVk+3iEPYGEl+87oT5WZXH8A5zE12uGbF1rAYTBzd0qKVNsYIgT0C1x9hTuSRSvw9g4md
GhEJ5Z9GlCrKBu87edroIbjWIoV7vD1NFp1mhCHREk3Ig+pk8Yuk+TeOmgMwh7DEKvAfJOr9g2/X
i04ZYZPdaNAa3ty4He3qxS8MTKDkucmwKf18Z8/smYt702FrVA0+Y9hWYdjbF+OrI9Xq6pVg9sZy
WlVa3MJowY+TL/vCIygWOTFnliFXgZjWj3Q4FyrUVRArqu+1PW6OTbEgs6rlqd0INpXquNo5lW60
CWNhkB14qGIX2/UtTURjEZYwTqWXFldwzyO+Z0KEWwqL6JEj+6ZbnRQGnpAWxQxxM4KUh4PwL5nd
AvGq0WwyfPZVHw84px/34mk0P4tGmY93WHS+KpD6hpwzCciNhXBT1VsuafCb6znjlx0cHs166Ep+
TKa+e1t0vG5chrOh4FM3q9G1HZly6ZdQk3vFC3u/NXn+W8rF5SVMHEmoWfdlNKwGKjgw+liO48Cy
KuzfMRxG6nY95qDo3RhryERVhZ022xi+8K5FuHxxBXj6uNrLMEu5y3fDZuZr+F5vZZFHG07OS7oi
AeHpJjOB6GK1ArZlGK2DXEdEW/cEZpfglJNnv1P/77/BssbzHthCKYPt0bIjixTw+P78XPDK5LuA
fce8Yd9j76tbG2rdW2TOoj+dJIhrQwltfXkIxQFve3oDND2/rWYgkPyf8Bw0FBt1FupCKHSweXlZ
YgEbLB2hRkJ9/ZiQpB2ijYwrzG8A9OH1I4TZ8dv3Gw+h+qw+/xKTtY5QglAeRzKt3cywQE7WPgOW
er0CyQMcqc/x1zVTgzonnN/PRwlAqsFpqnDZ7w70blMXCRUaW+jScBB6MXLBRs4XV8NExcV7lVrh
7rQDhFCn5e8eIr8kZdJ4XFYy3++Dr5mGOGIJbA5aSrCJoaJV4/IlUwFQEYMTpVq9tpywQ/3DJDAT
283to6SNIGxVmakYaN3ROoUypneyEo+SvnmXn2VrPNiBo7QpFKYioMOUNxRhgxcILQ6krxADV1PX
DwOoI/grSH2qlX/Ys1SEKHaVk/QtVmkAaKBoLybX5DFKd6lu9gvZS0/CVDilPE/1+KrZu76QxZCf
U8SgMX8YbCH+96nma/7FeWh7ThdyxhQFmckj6XEAbSXLEm2NOPV4qUDQvRhOyOqNBd/rJ8p0vuIu
f/qpN3ocb9MOMF8927rJjjJh9pW1W7mn6HvOCGDX2YZfyP5aQ37UXy0h6OYgkH/GJ/yLox/o0daO
dbpu5WrL5qCbbtyBj1qb8GcN6xHWduzfN1gQ5lvv09t/l1aa267U2KjjHrKpHFCLZJBvbyQ2RAZK
AUcxEHN6nZNsNXVU8CUuUV2j+intnX/sWLGVUmfXakUe61wdPCPq1gJ4ZpaemrUrvhJxqthHDZ49
CC33epjmRwdugvCb1EjAcsUXZiEZV22J3a1MtIsQQWEGhVhMssLmmaPPwiFJ/d7HVOy9YsSLbhUF
bDtyFxfR4gjK/OgBmDhug9KW1BPlOKVmd4nHvrh3armeS8rzHDRPi2bnoP5ppnJx2KacW3Qw51Wn
ENS5Qf9KeOvpDF74sBAxh/KSSEHbBvvyapx8musx4CEjUoeYuFLXLlhYWBUOPibIHKrSZzAfUzq1
HPVNWctlM4q+pd6ZSBqFgrIwQhquosF2Ea0cyOOrrmehaWwO49TGLdTe1n+jd13I6WnIC/Wz0xzE
zSpPWR+L6q/8VxasN1YvZsw=
`protect end_protected
