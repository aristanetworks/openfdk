--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   duplicate
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
g6e8Jp/8hBotqBZR5Ko0D79ebvirWfv9+rBNC2SLWBNvwWUlCVPbS0Xk5Io0yTIloWRCib7JEnk7
K6kNmz+68SeS+w5iYkN3FWl8nppkky6DvXMHk4WBE0zOGqc7Yr6i76jkkPBgmqQPRO547iGiTjQ7
QHlrZDtMl3gVU7HxX+Yb784rTasLxEFZu8Os4K0qb+9AVKPiyS/p1g10dxJU6m/Ce+npdoyfZT1F
oWYYg5LF2BY5QYFVbevrM0tIGIgDQNA6GXraMiiwui/8wfWfvBEZVRyHTbLVxo+yZDC6XVbwkymM
hk8L2vgtpllNHu8lqsx/fyWDniH9xPWmjIGT3Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="nFSvcKb1p/JUGIDSykWjh4B/cs5+I7Pk6G8iTfi4sok="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
WoHjCMWMfb3c2o3TUMqNc4T4BJkoij30AICq7O1hJ3HCEK1EPtpChwOOVcoOmWm9TzNQaPNSMY3V
ItmLMopwBs64Sb3IdJBv5C8zGlsZy8bGDySXpzwBEc5MS/4vlZUlbOyy0XYDdqkxIe+zO2yLjU3W
wjyw/LcHMbfuMEh7QI1YT7RhAyEiI6F4woDqfNvDTgVlo4zKZVDjMsCC/uUhROULX3t4Wr7bAKU7
0QHW54gxFdHKGcL0jEcgevndwy4h/Yged5qN8KxGAHErbddTnbyHT2QiFTjucCjcWmJpBayhqbpK
bMHvLDIPjYJN9xGd/n5DNr0MMg1uYLU59ps7vg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="hXU6fdawxJjsnZXmkGuoUdgz4SKixjMtmbRKN6y3NmE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22704)
`protect data_block
4++ZdwEBU6XwLrvE0EPbQ+bxEmgcig3gFSm+DLr1dv19QXdDstiQyYGBQtTyW4+EI3wsBRNyF+R4
Uj64FnZRMVqXPwqmSbTCNuJ9ckqBF3MRISwoIxwIm3c6nNAgTAVe3SRCKVa83/ZgemG9G5fLDZmn
JnML/JKCBYkAPQh7qNGaD41UkSV2tvBhsH805nOxjmKNHueRhGNJpUotTw24mAD6aAxIIIRQHsPW
UFUZ0uOPSw/xszvxJYqMeYeC8MBwOZbcvo0ejWl5otsDLd2DdayQq/uq3X8LCWeynHjEEbPmyXdN
Nyq97xo1CcnPVZOD2F634YIvA3oO9HRxSJmh+7t2lejwECRyoLze12OTW7ScUmpwSLUC9pKaFiFk
5OEBUE/b+AHftnNISBCWhilrh/WrkLdlAUV1/llMVvC7ZRi5eCx54n4h9Jml/rJ6ezNcqg+ZfO4h
o/E+iTLMJovRPIhJFzKY69BFBOMwXTCzbPATYybMO525ErD/GxPzgYUshxGgIP71bG4OKMX6rcXu
aLHM3DTYvFStqTp5NDcDeTWYbjUE5n3JGRx9y1nsWKagG5HwBnLy+bezoghmXPdtC8b0n1FcI2Gq
Plem0lTRvPwk+xsCFCw3lQ6h33H8ZJbHInoTmdwdKEfcx51ZkDNu0WY13EjHO6IP8HkWHg8t9E+Z
V/G8kDpg+d2ID2zd3VIPP4BLUxBpGjfYLw7tQg671zAf+iECbKrtnaHMlyaEweMIddy9P3kEgRsP
6KYq6sk+aaPB2/nF3pKhPwBc5coZNBs1wTTamTrqipEstYajne+YFYu9slQtWapNegT+WosoN3b9
vBxM8Qe+gLiXS1FMcLmuKkztQg/9sMPEM3IwwbEs+AOubeURp+i/HW3vIuRmegaG8CbQBjpCMQ55
nxR8VJLzLQb3L8qdO5qfLE39qfEQh4a0E7eEHgux3tgwOVvwcyHglvkpBUA7htKnn+rJpV1S67/x
56QU/SdUAuSsTULAKLD+gO3WJBMw0YCEQ+PSynHIe+s7cITBcO7/rr+mjqhaoC++lbXhrZoEMhgk
NP3fRsbdS2zlNI2Bx2CkkRSm5GGR8eeOX+Axkn2nVqcoI6uUFWzEBM17Jg2ovd/Tc1ZQGpHWImJ2
N0WDctb2CsAn24xZmtbPvhJeXJGKzqRiLaZl0ULRkbUyAuoty/N6IYWfZIuxF7+vxR/MH7aZttnZ
xtJ086ZljN7rSl6hSsxl8xZ1Wy2xz3UzN3KEuSeF7TFOezMxdCkGFJWCC8uyU0T1AOFqFvPh3E3V
XDDeXzukMqoOczRgPSGJ/jghg6YmdZOSBSH9deCQd+jQ+yiowjHC23QFhPAGJmdWtgVxA+rj8aI2
z9kIt/ualLo3rKknBa+X7EMIPpEkryGGFeO90P7iD+STzQrl9LMSF1v5+pvUe44H8KX+JWm2chJk
3NKU3hYNSBdV5tsXMZXKjmi2SBY7U1EuoPpjYum1uj9E+XyEsNHyoz2q6UTND9+eJzvvTiWY7adP
WHncodJ45ABz33cPl+lATRCdcas5BDMNVjBK0/u2f5z24MnAlafACzO18YYbinIQquQIFXMbeoUL
Ux6U+H10dZv81XuZ5LduID/IxIAejHBdsqPSOKKxZDE3G+mg6SitTctzzdRIQ+4ZSZkw6VxjvIre
Qil2UbQm12zuog/iLQ4VQFAuG1Zxc09AcPCfDwz1k7B6H6aaMEcRpxDCoKVJwDDLupQBHrilt9l7
89zkOY+IXMnzmTPYRJ9pay3ua46Nfjd1SqSMyujJ9E9O83HXAuuxAUg/fDr4CXfPIADyAH6nXHaR
BJEZVRMovnkZloYsj59OcgXNq4kV7E8sga49IxQE3LCuInExayH3abei+vvn83HuXSOzuBnnalB3
KifnTzMj5yEVaA+XVuPHwFL5pdrklEwFxoJkHX2WXLOkZ9kB9rW+oOPBTmcWXiifmYHFcs/6R1YA
xaee+9ZNsjrgkl3jD+59VuP7W9ti/buy2BxNUqbrlTznWgzTcDtcxRTET3PmdzqjipLpSSLMrLBu
XJIHRbE1nyrdiSqtBQ8PuL0n+Rx9Ktcvcuat+rAUqWj1F8Nv9AXFaUrxuDEbB5whwBKL57fkIJne
VFygx6j7NV7pTRWnKv03nk2x9f8sUPPcweR/yh9zpRtDLi5H6EXBRiXGcwz+sWOHQoK/uhU35xJR
mMBpvdKQvdKCU+0ZATv8sAbgjEXSgGkV7xHPBST55ET8aneTSyKAflu6EHXBy+/vHHzz1Yy7sDEI
qOCaTuQzkJdVibjFZOxQiSso0SDAC40qQL2WM1KqYD0Y7X9DC0sifqlrE5GcSaWHuAUPBvhpXwsc
ZZCWhhwcezRz2cRGXThhjfgHeOVqSeo3Nm+YPesqIEC2wlVeVe75m4xaRQILuxjTT2aGuacFEEp0
OMxlekDio8elkyun5qUg5I4zEzK5oY76viYlawCI6mAk6q9fVV0tEMVm+LpJRIKLTWmX++rhFjDu
Z4vKwFAASZY8TZcf73NM0VPzDzJeXBw0KJdqTwEzbPw0z2uXye0WpqXS6DzBfSLvQ3vFp0gmmQZe
EvMveacirZYtuwAmSDiroDbf6uVkOVCsuK0BxS9kD34XGEsHDz7iUPNj6SYVHjci15QC04169Ttm
RYXApLH7hirR+lZ1Zwa+53nqdqYb371JBRsfyBnGGBPTqL03cOT+hSoJg03qt7bfPcEW8m+HxAWV
bnl0LtTC7tM57Q6qeYDCJytlZfPjQhjYjFt3SvrXvHj+Nwizh0ZWhUQeoDu066PCzJAA0g0QD7dL
0AzZNnLm6dtNxQyGSM+3faA/NOYEc8PoOEIS1GIk/r0AxgttDSiqPjgS+0GwJmm4vLVxcezjReUS
XTwSi9b+EY4Z/FbYxdS0x+tgD4sM5KCfvgHiupbmxmZKqL7tAXl1T7yeYBj5NzjYHaJZ8K8uZlMp
B0ZwXBHLKyeOJXOiKiPaiyby3wfjdCj6lAfP9vIUtpbfSMCK/DyOqgbSjg6udCB/LI0GolehAnga
n/C6/+pDSPofioyPsI5DiP1+5kyCYwB+RuVNbSrRy/twX+Lst3y922pL5vTRLVn67FzFYHSn16Xl
gT6qHZZGuywgyb5VKVX8B39kdbP15/SsTYIcNInJuzV2P6i1zzJMievzAWTy7ZBs0AZAwZR2iKge
oRv4pQsdtggfdDq0qEEQW/UMJ7LvnJ8AZlZl0+H13t715Zow0TRZ6zR2YwWiz4BCHlxmJyXbJPod
3knwVKbDejzzVARROruuKnFs0gEd1jyZ+51C3Y2Ws7lW0hWW0FYUuW3bpmZrGOtJ7fd2RniVaff4
gpQmGb/STpAA5liSaIN9KQG5FUNCAStxqJ1xpHVhLOaciysooCv0XgIx3j9QKExVEuskCnDpNphh
h09nn939bvD1c7aNN/bGVs0RvjzrP2WymtrlOYqX/vgMkxo+HNRjBFIgqZXecXxeOfgM7SgMQhb3
W+GiYhFIzsAC2LLsyymqspObdZw8kKUzdBWlPPgdPkkm9WQ6i2pZbb/XjepFOkGnT8meW/YkNAou
oY4ETgG7z5HrLnSUPwim9dFT26GDbdbpzAN6zYtfvXzQK00inj8Wanbsi7AwyczvJfNhyBon4j/E
FudjeMi+Nfw0z4p2brj2e7gP37pgnFQQs6EoQzB7o4MaR9oqpC7Me+49w+IgGl2lIkC1D0x6kq00
N+UeRiTv0x//q/1GNVQpd5pJO9c3Te0JrKmz7JdZ/0SFrrmqvCRfayfvfUkyNFzlIaBb3y9gzjOH
WfWkNFs/ts2t9bI5B0zAglHZoTWITl4H+1iqjd3CC0yrutyqvdj6NTUyCWDTIta17PcbrO5CaHiR
lYCLOvKCeeTGQ6LArYYBYgSc4fVeca4gBXc//uUd+zBqmFGnuZyL0zy3in2V2CqfOwYnpZmEvsJi
I2MeNG959/23VzfAsDaCtsgQC0BieLVtD4llEYrxBaulyzfK/kQk2Bgh4q7RMcZtDlVtmv22u+gd
K+mwKWV3FtI7GH8xKxNBriRg7Dq41bbP9a31pE1YgBOtbTlFJme4oppvuzmdCSljAqjeEfk2No3q
i1upUPvUMZhdUGBx1dOjMfyP9z5gHvW7yWMWGda6kPxarX5uWICL0bAbDQhksBEzJ2eaKLNaMhNy
AJzIBa5U258RvdAj+r0h5W7mEqETLde3KPSMdFMnNrmkt0s2xQVaO8pNv6yP/c3tHZZGtQtgQPis
wYPV9YoD4dXNF2pg3mg+OAVG4j73DfyHNdp+6ZBACEEBoXRAdH399ULKXnY5kteu803/MBRnfJva
bHFd88LpWJ+INp8vn/rRsEXSiai24xi5FLtubj5cZaIshbx1AqZ0rfBsDce3S/MaSI7j1zSgb5IY
SrfAhI9fzC5g795jJYPlXnqSoXo8U+VK2ZYq3j4rBxe1cYMtLXELPz0D/YdlducnjTc6odBemfYG
Aw6gAkaWmk7w+NUXWfV/kf/lzDvtxuEvc/GwNzA3RCUlt7xsAR+p7uJLh6v9Vk+j3ztuak/koUWR
3yMGEfWT9XdoqCfKPPFGc3tzUvFrAwzngD23yzaWwA5YwBAyO12PUcYUGpbrH0fknYgddZh/auf/
ADoAM9g6b/df/pMXlKGj2OeNTE8aEzosNGkg8Q5/CJXYQZBfRRTdhOP5pmjM/zySLDr5sClMYX6B
5aRtHOlaLgouANOqjne2MQUhOHow6etCmU/bVfiS3EX/5BtXOlrsQw4anEx13dRgKZHjrnG6ww/6
NLZGUlHhlxRsQ0k8HTeo6ajkP3dVCk1S4gOiPeuEgZqFtX+jVjEVZTsYoGMylkb9a+LlgzQL4Pi5
zRSDhHeAMsr+q+4xkovgm1l8cktSy+8FxdvLXR83YC3qlb+naeRlitaB7nMZW/1TeQvZI/ynuLA+
5CUaXVjfB+AfCAeNolTODVPHwTnbcRCEyknFc4O0HH8XcCgxTtN5GEAVqPgsvslL3t56q+mGvQiV
y7HZ9xaPMeO8ZrK5GPUOij0TeKm0TpAxkx1x1cMRs0nR43a/sYzVmCuFUZRWV5eoNoFafiTDsDsv
96bYVTtH8pK2DY/BkhoMaLDoGOPeisfjK8ThNCLyHDKDlPSVlUTJgw1H5ZIxAksNdMmM4WoDJ2P4
h5UgTqIzwojF/RB9qhORJ+95ZAx78uBfdImISUa7RaD3+Hwg3I8B1HenNKqJ7nTDdL6vANZtphQk
k4+qihNexaFgCPADcag36jBwlYoUbHHdZhb2LNycuXbem4sbxITRx7kptYz3wOPVCWY8QIjQnMhv
VkGWI8Oc/AvTLPGNkLScMWpAqdka5FVFRrxBbR8FnxFf19huhQgQeYjztO+30ycIZRD05KMTFIUt
yjhDzQpDb0DtGgL7NqMXX6NGquWTc3L9dHYuJyICLucIJb0LSL41792cMuB++BfAQjQlbbljO7fZ
SPwx9FMeHdYd/w9rSrAgI2IISR135RPias7ZdeVWn5k1KY7u84TK2YEGt6wsMq/V/zdwKhCGPIgP
2yVFRZgSUcpecm0v+SLDhlv/ln6zGn362Xnd0STppe7F3kRIy72+ulSQKIfmP90ZAipU/V+E0wK4
kyv3EAD7sFq5iB1odUbw5qnqf2wlwLuQ5LiS1K+2Yj+ycvQaeyItVWZGxXYdTsookZSSQ4poNED8
fT4bGBRkHn7O8fXWOGpzsaE0xUdoTITD9jH63k9UY4ox+av4UogavJoFyPxj5IV9qk9OADIrbXsL
gAzxgAXoL2PCwRWLM9SqiO1iFNObt+XjQUCZ7J/ldKyn/0k3sX2SV5nHDcEzBAnYbfo589j1wxRk
Ppgufg7zXuQ7ySowzky1IjDCmqgz2SgyQDT7KieXOvdoELPi4j6ugkZxralP+LGYkxgnoTqg89N0
CscT59mjkkF0UwdaFdEWD4PFCsGhX6FFIyauNr4cWGD3PwZnG0SzyvZq1h+8J5K7zFd4gY1hdMGM
/8QfxEInNxgDNmf2rBrrvK9npVI0/ITscuTi/HQlimcg8tmRoBsKxJjfn13luXYkMgaZQXhOatK3
4L/yTDSXpJWeyEyPEQV1jepDvW8theA67N+896f1j4ntGVazpRBYe0QQ+rp9xxwGm1IBqluosVy8
SpxbCzNIXx/NMQAz7wvqcnOXbtcJquPdalRo0PrL6Ivl1JSjG7mKp+H4+bfgL3DwH0gktbxG7odd
h2YWUYE3LSCU8yIu/pxglWtK6ef3lDsf/5YafTP54ICWXKh7rIHzm1zzbgwLDVy0YjGHdMRzvrkA
B01DxURwU/rqt6gLz7dOQSXKobhMwh/+mhHVFkYs2huM5lBEQhiKvTBfb5GvdRXExywZyOOAlefL
3ZuXHDDOf3JE0iTwm87j/U3wGtyg522N9KYQicIe7ht5G+E5cLiLF+WWOvcT3x1DHcjuYOp0CMy/
XKaZiY3215ir1FMXoTVgRJLvImZMRWZSmfDyRuUaO3608webjW/JsZDcMyiHMJMW19rfxt8D6PG7
PvWS7oHJdp94kJlnW/HBqfxbr9+AIqAKQZ2rPB8pqGt03rkQbK1DC4jle7IffejCROwQvmcGdW0L
Qfic13XIXa3VLWqbjaVZiRP3PGVdrpeiOmwZH7CMKIombc4bjvqihCczPT5ISO7VWbfz7J8XXq/d
hh47/cOppgxBCpGj1r/kO/h00mBm6O3MhGz6Dazglg7sYUFBrWU2Pb2WGFMImGxAnqUl3FvAAIx1
LbEexqO2S3LbpBp7au/g3VlKzLZzTZQDA4dC8yXVrI7VWYqPgEKWwuy8OS3BNq6W+82ggWH4DwKs
ZekalNXa1U+HDVg78VuNtdeEWhEref78jk+cbrC5OQEMcXmj98BRcA0HtlPJN0+uYmhY3uDFl7pC
3pa9C5QW3Zoh1RnHimXPi2vY9p87xzduHd1160HGzwf/8y7nRbOBF2E5z2uy7QmUOMjj8bxItfuO
j6xtrffuLeHoV3YGfyjZHD3E9VJ2V2LYaUddk5rz38bFFgWnJawR14selgVXCZ233J7niQ7o8Lae
3q5tVPQH1oa10igmtZHes6UD5PF3FXGxIVtEUEGJ0SgbBp/g/nHYPwlJXLPlBkXpImdKQV53A5X5
CTsWaCMcQTsKnHtJlb6Pk+cDyc3gGMX4ZbZtR9NAsMdms+Ot/DFjAsOCJR4TZ9e4NnrH8emXQt9s
xf00eRsL2wfU9QQJ7SwKyOXbXM3rzyzePDoDOBnP0NHusnf73kP2wtCq0o+rBztwo3slupKe6lZV
jjitKtt5iVOFjy0gF5iiuOySyCZaCbFU7w84KluWkDA8DFl4h/14J7ZDLyt9E5ZA7WbX8/29Cju2
vSUQOvvIy9MsLqEGxZG1kGZXU1cxxj2YlZKPx/1ws4kNlUApZK5O+kc26ZJnRsG/8BPDbyI8277F
pvKCwFgcR8W+FAaX7uugglBxyuD5v7M7lEKHx8qp/Z3T/VmOcIXisI4jrW+mNbewQbDi4NYL2ACh
4hPJJ+kjOFhaBXmymGKPdo6h8KCXR8xK/sVjEInscor+RF/Sj6vMW6mjBJdE58hyl/PTmbOameT8
7HpDuHm9f6eRDrYOEtl47k0Xj899V9qGSPSyW49Lr7Lg+Sw3J7SRDd4U5Ij4WDRBD5PAFyYTz7pJ
2lx6GcxrXO5J38h66F86YLweEdUOt6AsLfsyrNuZ1SQHK9+WzYbaHXPcNPaL822uNSuT29fNOmra
CNW9txStNFPMF1LdTiDJgMRrhIFekWDHXL11dKCnmvpBUGwE4W5XXo+yZrbYxv+DKP99y5QmoYVb
WuvvGipkHaZZ6ISxZizo9uO0K95Kvxq0T+RDxB4CLvi8tBTG0nkeOHmEkudEqh9pPyn6mdo89EfR
7lc+h98i1Do+nVCvdKPLaUNLszM4mEo3TJTkZ5jgFr1Y/rxuWXZsluikYPO267sGzJCJU1KgcgUN
k5FtKWK7caQCPXH4/2iBzR0iOz5AQfbOF4oRIp/Z8cfP5j5qUQli3WH56O4RghwwMwGFazHyRwYM
C7aeXzP9+J4l1IUgsIkElhHVgNdU0GTgawWBDZxmg28TOzWDA0VPd2wFr8fqnlQ48ILPnt+gnq6c
OuEmnncd+Iu+0q4E5XFLsh2YxQ5s5ETK+hwYMMdzbJbOgx8AJEtnwBU1mNK7iKJQKhsEuRlupqu+
xl3qsXjV9t/Q83vdhh0g4zsNSviMHwNbtVfWNAxB2HV99YA7i7uoEMuY9oXrgiwYaomywo5h62JI
lUUUn/OuKplZ7Idv5gwC08o//sGZkDw01no53Sql2Oln8n0IFtc0qsrgETR1swW7qEQ2NpRXq5fS
Sg5vJwsbRdz15FunxgQEVgJIkchrWldMAxdhMNIk4+XLz9B3f71U/UY+TWY3IvuB7oFM/0uPdCGT
UyFj4F4uuS6rMlteYxDuozA1lDoZn0LhZH+mMQC1Bf/vD24FwLc3tqQrkRxSxUxVjN6fDkzBBWqv
dAYGgX/i0ixACKIa9skRF/1fJSErfY7jAsqlPCZaZlYrigYCrV6xyQB+yCiGkSIggDUqqcDdR5fr
L+O3nhz843sf06KheLpTX728x2msMhhQRuXSjlFhKT0bH4+a0IQ1VCXFBnk8YfyT0kXwQJV98v73
4Um7fMJOYOAbBBPQ23P4cakfIbgKTCXtCsBt1/+wnQKivKvkxo4D+6llL864DPBXYGBTYtg979tO
gdiVPmUx4IMTJCsRu5ZlQQKa4/XCiJ3Cw2uILkaj9FI4xq0Fc3DqBe/PQkImRiCmn3Mf5bpReNXL
LMMEb0IUyA5aRB3XdiwGnhWzjxsUGJcqbxImkl7xpdJL0fAaNmuuPN0bfvrC8RirQ6r6LOF9cNLv
6xiyukwjZpdEgaH2AeiI7McuklJbXmOFYtQlNCXHucR74AVE9pvkJ0cEYBbCmvVc0UrQGiDZGjUJ
TdEJQRTeEPwr2d+sW2XGzqYYchkbPJ40GQnlYrcDeW5ZfTcreKJAz3TgAWO3iBVWbpCNU32aq2Iv
JKZRmeXpGTf+H3yd7HXP1eXdvbct+J6El/vDOTz0eg70lQhLWsA+82xrv3J47VwqPTqu5DLwrllZ
TeW8Vgrozf24LFFT5zysfUIdYuVeMn/WyaJWUryS3UHeeyD05N1+kK36srrJ4ntVeiVABz3AYAW0
hRM+Wo0AM5roE7FGWCSWeNi4qFdaku/+3be18uVzVBW9flXjcC2EAGccSDDFC25/17oUMXdLMz7a
3wSLKAsoeWyAMOPA9SJqmn1P9EPgjL6wbYAuRQzKuLmdoMlDsG5thnhH7z53CDe5XHml9VCQilZM
2+jOB87+iJFsAsIgh7rmnaV6VXwNiUn0uge1HhkinJT/VIaeZJj5qIXgIf/TXabBAJwEVJQo3w88
1edrBcN/3l7wuN0Z04fdvQMpcCxALdlR546PuByAioJHnV5RUPcDHxubzzDzJCt7MJrFZDQNQWOU
3eeuTm2TqW1aHJSwTwbU3OEL4TKA6exMdq5obAr8sdBj79qMr2OA0RfQae5bWiQriLbKzY4aEt2E
UPZ9YN80xGSS/f0dOqkZD6sSofZakiUmiGag6IF2s90QCXcGc9A4F3yypXR+fPBhPCVdOT1qoynQ
9FKDRGKDwNK4WV739QQWA5QF8ceegLqQH4ltxqn3cX+OwYKgEzGiCanGKoaJnt4A2rK4do7pqmzh
XzpBWhXSuarKvsyPcreeTlNPUhZrIfimF4zStkq0JT45Piro7TA7TuEwzldUwM4ggZAoEaUw3vL5
31M5mj6OGm9yxT1ouCZUmWgrEDECuiwWvYAnzdfFYaA0p3kw57sbNa2Ss/4ipbVeuwN+n6j8RIWP
MNEOZilA7hNqdcKOxHSdu087UsjW3xlHBpePr7hQc2UbMVLA2OJFUXJa3ynbDkzIJg2YB1gshB4B
1xs8U5ed7n8K4Nz2AxUWt1Y9MrynUk1YNwLy0y5ampB0vLEFJ5xjN+TTFPIOQHyHMn59Gjd7casY
46ddMTdEKEZcKzcWYMIX5VrWMsRK7bRDqsAOY0Dzh9OI0zk+sWZSqwLh4w5ZEAursmsxCx6gYMKk
6x+LehaqKS8s6NFVGuWmkwhRhZbQm2Sah5RCtkiciDcFFhTCCkSyywPT6J+nXObfCX6oY5K4IzFB
RHewsjYdjFzy15fNBfkpZ4++26BihGljyAM/XKoEKBrTR1NgZy6n6TIwe1V772jnwTyn7mDyjz6S
X7k+Fv7kfWlozy9rqdYXnfqbsA66tRz0SG6B+FewZ8K+DK+JO7ALBVNZ63HjfO0obVVcyAhPo4pd
hL4/x+xPNXJu5/hNfWRbO2njou68dxD3B+E+lAynhRtpDMe+CRP+34IH2ER1ZrX+2FhAY2RdGlHX
UFmH1vZhplPvN3+t55tQ47oLykpDY2H5CR1cjAyLzYRj2l355Utu7VAJwqfKKGTqeKzZU1WC1n/E
gg3WNst1jYnkl5nPKDdqbGjEMFlknB5WDp7gY/ErxfmX57sZhX7Uoh/MCOEnAttRzHF8IsU9bTzH
u61AmXs6YTFeeKdSQm9A6hPLashYR4uCEq/JvwDBtvqsV87eriT7fRLPoEpt6woYP/rOhZfxfon+
od0pfdv8zQsDD/bVkndAMisBlOdsF+pqHivIa/mpJ2xuY55/DMq5y2SuODYXYKQVSgW1OknAyEYI
UkiVFkgnHzap7DGMos51VTegpwC6meVDcpDpgawVmgWoFX34KwepfqIIliJOw+TpKZqRPAj8jFXn
njExhZ5Um4vucjxi9wNIF4Lac2nfnv4ogE0heYWHe1dlDP77sVoZ1NY1Xq7HtumzNMn83DpWqSNG
NeOS+YdFaHmLOBRXbThSfiZ1gDK/XzTVtz1o0+p8Ny0vrbpApbpnOAW3gAU4LookPE3slHsGxCqf
w8YLecu8X/XZTpka5NELj3UUAyEvCteel8xavSvj8syZrUz7LRUqJCvueLnsC7gOczuxi7I58AJ6
WAAOfIIknB9cUdn5Hq+Iu2t5IdK8nmz+rbflytouPrmkrFBeKuByKKqWxGGNJQjp9Z8H+7s5kJg5
hVTJ3qaX2OmXezJ+H6pWKRGFAHAqu1x0fytpPv2TPT3D/V+k/g2bTWHSnlSXdKYoZpW8qMlXMIbw
WLPmSVFf98mHqR4j6nSLMDF5cazKR2kI0Zfjct8hXo/jdFDQ7+JQJgtaHRiYz70mQ2T/sX4rHMKR
qM/wd8yBJmbRU13Qwx0QvApCjOY0vAOUDXkTudGQefy8jaPd0RzsGlhuQS/glQlaNudY2CAvG+Vb
oHsURUSGQjP3LZzjcqDyXp9S5rKCYnjPWy5V03DWLw9aniHiCuGCeHRdgOIBs7cx/thu7LFqpUgF
fmQOblGWKboSwWiR+EwKYXtie9WkKdQLNnq2oC4Cniwnx/02FFBdYIA2ZccnwsF1KaxP7mnp6N0M
i/E0NbuhAzJPBYZ0DfZR/o7Ib7NdaVWyIxr/comvtQsAyKhUVXLhNHYsTOXoYQ7YWvtrZs5YxRgg
gLLQDbV0nmb10uzviHVHPFSvSRkFRoqhjIIgo7+Al2STSfHnhXYJgkr39JUXN4xquqmS4NPMZgeP
nY3Bp5Re2voSWMQziryBNTT27xk/LAzot6G7UsQRf/O6hN6boGBvjU1iPJyMydvwarmaDL4ORtF5
FEj5m6JZ7vibhB2+YLXhoHW+lYxY9cB12nhLBaQsFDYyhW25mQxgsduGOE/AZ56R7ULUzYVBwKet
pbhifoQFw/wtn/JrzTzbcAia21Qkwv1vzQwsUmeiMW+EWrb6DDjnTCF9FQTa4Ye/Js7kMXfFuiFy
uTVRuG5QPtkegE0Igo2AKmA3xCJM+QWsT02C18n5bQ4sQuJ4TZWClD3WkhqBWFtqlgbXKPc3Y+/m
lFlYW6ENX5FTMKLHB21cQlYnJeSrek3gAT6DNRc/XIV9gAEcpb3nbtufsL6jrEQwJ1yu81Jc8/Yz
liN+sepP43IYFzb4Duup2Etg1+pZ1IOegPETtAhuaJJMqPSMn4AhsGwVmeWMvg9OAH52svXRg5bA
sotvceIK5yjT1yqz5oTjoFVBZaUZJtvMIBsuEKossEAA0ZV1A2DKYYb0B8FWBOBZuIU+YLG+w9Eb
Li4wTRln1pZGiLJezFkVo5GAo3wb1Bf/RSA4tNgiA8tG7qNLbUuyn38DRm0HswTfUqgpyPdLVLyL
444vv0b0KZsqsUgBPdhuIVsBkvNxrgipFwBo27m6TeBF6ngOCIj8GUIFImnVWQrQgb7xXnkprbOz
hotLgMKTUCZ5k1GYOUEBTKDPvo6DjUixNm0+/KCEbMufjXlc9U4+fFZA8GiGG2cL83iEsu6tbcjQ
vHWhJjZq4VxEIU4gsP77k1DGoObsfvQaxxPk5KyGo1XBh8DRRFZsCV5ck8yuA06a+A7fbFk0DTgV
NBbKj2Jobm5WRwgbDugpc9DkZLJ1TJ9rHAFRU6y0a0KOyP4u1fc5e+/B0rN6B/fAOGShVYLTv8mn
Mt9zumrgXkIETMcQhqR3jIf36KTmWAcqGsOM/a+ouUVpe908XwBUW3AoXakl/4eJadYj5qI/B/FH
9uHv6fAQf8d9Djd2XdkeZtr5BVvNqMdjEJLijnBJ2MQtc4anidowwcKZGrTGDXbPPw3KilooUGGg
0YSsW1C4derYqo81ak++IKIVE3BJnVuTh7rLjq8+8rXTOU8X2Wh+6wS2Unvj6YVK/b1jz3J0ri+V
TJtqTCNV7gOpEOL8g79NXMjId5YP/hist+bwCSQCN5Lb/GD7Ky6Av0u6AxEjKQStxnOP6g678LT4
tx/TUCVZtH5Lt5mkSkVL/iYyl1Zsyh4Wo8bQgLTmtEWiXEfy3kLhpyO3kKC3J+m3EYGzM8MZkoIl
9Ljkk55+wyGVjnUxjY9R2Kp+dYg8LFgxD9SajfvtGlbqLxOmD9LcV0qSUW8qYmaCQ5S1SOmExbcp
LZ6J9Abm09iqQ82FoCCD6//OOe11fczNMLHO+Dbv+IJZT/o3+yX4Rb/tQrTJi8YvM+PcEMrDoYUt
NmRrbCJ19u7PYyBr377wxgBLl1Q/Nfz0n2M1YWxxC8tykBDBakGvGNUHay8GE3tnDsKDkrwpP/wk
nf6V49pBB3At3p4jKGjg7fwgu3DZZe/m6YiSnvSaUQM2wUmT2CsJaWYNxzz9ilTaLvcDWt7NsLad
drPqSaeJRNLWc1XDEgfCFre8V6QVKUf9eYCqV96CBvhutn9JOzH916CL9t5odNn9w5m+Lo7sfV3r
S57X2NptrmviA55EuW2kv6iJzhhuWIeKjAz89Rd00SKwcz3kYNTfiYcs7eXJQvB1mj+Bac2gyNOv
btnu0FuVYbBAINhXc9jqwDPFh5ld9fIQb+ZepZFU2D5woKpLCyTWNF+IyV9Tm4zSONALQ2TkgBtM
XiPJXL/da6ELixhI5pfyKmCS5vo/wTx75j3SiYB94wKcbiuft7i6XqCstdb9losY0WwjpmVTM0oq
sgApIm4An15U4u90slq08Az8uZh0fg5gs/6/ZEtY9mJr+R8TAeQoXAvA+ziFYR3DtQJWlnwMgAM/
i29/qSOtRzF0eUYEDH2R5+B2OPtNdyWN9DUL1Rezc7u08NBiPeyXVKd23cH1ccKVdI/DPpRlqxNK
lLqUEzJ8vZJNLnSPH7n8uxcPSQ3+5k6NThCTD85/Jde4MeI5242QbcjCmUaXy+nzUcG2e1Tk4yMV
fwBcgLrP+obpUkIywRV5RvS4vOLQk0Rq+Hfn52draUqFKC/ckd/Kvjb2JIg4pH26piHyZChPGXH5
tzocDMHUDTjQTa1JUIEo8RFxfGJKE2yr59SU5ggLEXeNQrNWaJePDBKa9DrLPU3bSi0oQPRAZE/8
WDuKQbcdVwAnejSC4/vxQL9q8YqJoiXfDZxrYu4fs+1CdZtNeVj+e0ZarMMViuWC/lCAUSpFpbTC
m8r1BkST4UcJluEFsy8zcV+yk5LwQbfsEfGel5qC0pDtI0fzbwRfsEoMnDs5Wnc17Rs0gnTw5XOI
3c/ykkkVP7uQQ7U/MmFCDKaNeEYc+Z/E/BWPjBkttyl3pNXlN90MBI2x+c4y5lGPoR5pX/advjHc
3PDnku2t9LBnEiEExQzpOrMxrhOPMuVSnvniDogGxu9gyTDdNrwm5SHrG5KeSbyqiRxKdjbMvQm+
Bhlaj6tekkY7ZyxJXBeiLg+ehYDTjJ/RcgaU0FdkKMevJTZtZI8BWPqUTb3WdZkcj42F271FFBCd
94MK2I+Ng10870qJHUVWiM0IgmNrfCjCxnqP8ASbiRX7hotjlWVm1V0BDBxs2kAtxCWP7qwg8d22
4SmEYa7rXHxP4viw6ayVHJ16Wg6pLkhJpzqdI106JjvCotvzkQA/6i1yCr9dKrv1JhSfEIqZ5vJk
g5sfUS/8K5VOAVoCw2LxX6OlPvACB0iVi+wqA5tBkXmDnMOkbKRwFRGpqney1B2ahgH7uDZprk3a
5tFUQVoMIbcfbIVux04nW4M5Ks9ZpOvnQN3IbYD8h9pxgDKNQxi39eCcbL5K0W17zcKHJ3QV3LM2
tGW3XP8asrBhaVY4ePOtEL3uWpqiym2roAegxSafeP5tWhMBlkT86h7BesAbGTMS2KuoDcLdbSkO
JJP89EHv2PgNcTzTeu/+GqGzlZEz4KE2INfJ7fDsQUoyeoGQBz0ONnHZdQjpvxt+OAb2OHCwIZZW
oOpVYHv6qT3eaEI0008sdMD8c0wmsdIMKI/4V7XSeY5uNt9J0X+Y3FCnWPIBvhEgLMPb1f6wL0hx
NX73J5tb3YoPlFPaGXDQahv1Gr+LYJMeANrPavQ6XBfJskaP03K3lLm4gLbtOSLP4S+FBDrf0kE7
XAA84J3Gr8tl8MngODTDrX89F6nFR5LHV9otg8CvkRljZEgsk73M+tqZuJ9W1yYLZ0K31pvUXLZg
Zn8piP4arZoQMiJbCFO8GkNVmnv6vhkugujEDQwkU69wFb1zwPkwXR7NuS9tV9mPjDEjKXwb7JIq
QM4M5pqBLn0BBQaQ1A0NYcgpPwWiXugmKNaFo1bu6WV6MrdtNGQ8FO+aMkH5GyCqGbfxT6eq6/8r
suyODdMf0Jl4pGiFflsSxoXZQjAGc6N4QRezvS7QPyJGcy/WKbOww3rqVy/kEyweaOhCIZPRwul2
8u/WKetoRBWMD9uj8QLl0fBbuPbCYLng66LASegzHIb7qJkntovyX/iyJXYYD2D7FJPyktUn77X7
zprrT2Vf5Haf/7FPldt6lIHHSjyVQ0ZuzPiIKw5fHyMSlxZgjo4KpZ9r/mbaedjZGWRPSsoQmE8A
iB0VJwnhhGzgJIKWUkq3V79+0/VUvrF+4R7yFI1mZyJdKfMsAwJNxFo+a3be2gDrvt6Mi+7L/b3T
qPhP/gxZnJmS3gyp7q6Wexen7dojJVCH1sny3WJiV8uDrRl2thdyB5jQIXqp7skKloxJlf8EfqOp
eOCRF+behepqdiXY1bBTJf6LSZvPrA+Bs3NpwdTs/Uz8ejf7bg+kmhXnXjN3YVRfd4rxCLBxIBxa
jlb7bAPK0CKj1EN4fF792zp/XftW0mBeXlcFBzEKr7muhvgzDCePGL3lr/MG+CoG2r26FwOC1QLS
xB5Ti+vXKHCLelM/iEzVunIpJNt+PLqny114SbdtM9m9/6igfXQlRZgIvN7iT5bHDTZDOX4BDHN5
RjJmvRkt1Zaz2xrbLmouBf85WuQcOUgS6hzHiLZx1/yFFupWrHQk5NlZaGPzZxnDqenptV8ZqICQ
64VE5sPb5VaScczQzQ0kFD2K1mFf4qsL+hRtG7SpxB+ms4MzDKnceT1NUMWxTlh6cwOLNjYxLo7Q
bq0IIBil12EcZcNJOBqPC+d4qh2pP3ZjgYTbPzHr6GEkLc84udFtxoekDYQIzcNUWunJxjudqNAK
CX9/Mb3zPeBN1GXg6IpnZnOMYOg4WJFpTW7VHZZ/GZ5fgu7dynS8zXm7iJmSp1+RDF4dnjS5bQko
FzYOGKd5HH4JZq0+dM1Qu34KajG37ZFYaSNSF7YixQRxkhdCjNOC+y5U5E2YCIU/FCIaIopOfGNn
y1odd7srld1GSEz2byzSOYsJT8cIjwPWkMNPj83sg8ULvKHfbnauo0b0WoKZXwgQAzJwpUEq+LA1
ssy0PqD8k+PT04cZGp9j6sspT0yk8Xz7NqBPC5+7iSQ8O0ID8qSmw4mLcbxTHK32YFnv+WXUG+bR
gVQwnzeLofYqE2Bg+RTN9plS22gcD9np5Hk3sxYfX4iloURf+V0mZlqz0YYhdckc/nYAT11BkrMM
WWlN7B+hUOnCcc5MxJM1KTfOGYyHGziv8FuLjfTa1UD5JASrFI7UVeiKMDJBjc8fdgNa24J8kuZ1
aXNO0xHKcxyvsXZa2hMOaGr+xmlUW32wcWxiwFnANhOqTqSTcZ2wqeGhe/l0QR7MwCE88dzz1BKx
sBqhNvE99lTBLb7eDVjiWgXzJ+N+lM2On802ySIuPyoNonbWszncrDzPfMN/nfGQ5NuJAtP6kmG2
zgudoSrxb2FEDT9HqfJwf9bw0hodQLesKZIu0S9ACc/y8avGOyXvBsI9IjRgALZ4wsecGVotY+eP
SbFhHMlpOMpO8P9O85EKeWkA2kBJsEiDcT+dJ1O+uHsW2niexAgT/5CZByIolEyYkyggBm3ikjz7
NiyspNw5c9edNydir5J1DKpn4CkW1QiqJUS1efC5F/DTK6tTTs0gPZe+l1FHHjexSWe0Qkuq5IwZ
/NPXbz57VQ1uXvdapeTi0n1sMB9kJ8EMVQAGXx6ZcqCXbybyC3ER2Ppc3zuXCOS1lu4ga3C4d5Y5
XUmZCCR5GoFKyiOmjlpmTqaH+ly79a859ZBUBp7EBW3ktHuCivhFIVLUhtC7pJsE0NUyCP8yuu63
WhRPkd6oawgrjfVHUXnwoVoXq2r6Sq5TT51bcq8iRMamHgHYkg1mgeRWfO+OLmeA1PCETwFbNIoD
2aKkBi3yaEKrgegHI+YtujsIKDZIn/X+SFNx1F1hwAcvFiAhP8YJB7DUtzyotvpsdVvjC97zvr9H
4DEEepX13aIlLeJmP5oGp80ipVLGymTpXFARsViEZEPnhANL7s2kd9LriR5HrX0MxJnt7nv3PUle
/C8kkT7Y7flbZYjl7FKiZ/MmaMsgFebA4/b1fes4hFrOP8QRU15bUXnzGUsbVsthgqc+Gc8yqkzk
Vio2kvBZa2yhOLdfiRGdpe4tZ11N4ALuCWe9fXF2VXgDhp3GsYyM5ldB8rbcIe5mSUmxT+hKDHNo
gOSim0QL9u+80U8jbWRtyt2x3K9FTEmAA4MepB37VpNSPlAZI8V502cHevWgknt16cpJwm1CO2At
LWY4qjdb5VdDay3Q64WfsWWSZvHPp7GOw54mf2xmSECNN2Wd5X2tDM8B9oWYVS3dJqErGlm2H1EV
p1m/BJyOYDgPG1MIMDeOZixXFKRWhurnVU1/2YuloTBPf9b3xOj9S95GqfDDmbcSdGL3HtqQgB36
sXBNOSdFjQDWcry4ByxtX0GljZovOC9+SRO+pY9VEzoazqSxOidUtDeHh16vMlrRhXc3rCLjVcJ5
zFh4B2WpgS5rGNZiQkp9V0CSlcvHqbFMdOLfaq+LE23UXXIZnONpe2218CsN7c6+0ZWv09snONxb
meLMqGtBGNx+SK/3mqpdQirZvvmeI3dlgNk/1ZUbV3l1tsDtu4F1pS9+NQkxlp7U+/HkI5Caydtl
i12xUsmPQ4SnuaMsMFSSsmAcskBJGIZLMg4TM16xPhVVFa7lk94NMPS8lzhW7xlQdAF0HDMThrT7
ri+MU+zt3qrS1foiA6WHzRi6+F7FX6bO9rSAszhQ0q3VsvYxstBhMtfpq+LJdo1myvU2h7iNxQBt
PQ5nkIdlIPhV/9tQ4GdhmsHx05wQYkHIceTAuXuqzhvnEReU5hNmYkMpGIXWw0spSqymchwBa0gI
ljYfMQrldIy2a2VOxz3WwKZ/nzdUbqV1Y7OJWpy5KIyWmR2lBTohhy4xBR49DyNQyTFcxy9c+uJ0
+Ta7yni34B70tgtwPZKp5prLBaLbJQgPP0N6gAJ+Ubhx4zUpgvhlwUNx+eFObBkPvOl0CnSftRaa
WCTT2Nr7w7rYEwabdJ+yNXzyMfO0og+TooObx9SlhKNkg88Dp5ppWm00jc0b6Hvw+O1LJcukT8PL
fPXeC01G8+rQ04jd10vuWP3aueK4Ubf+t0N1FRwin90zqxMZpzmVXrl++2wkm3PuUR7hxrxDUcMm
nZAXEOrMHh6rSR0hmKb/Gq2sr+C6nshHF1LtWj+j9S6G7+FOWqtzQqS1YMuZ0SU/WJOUJ37BGiQG
rseD/ULjiwuVGP4g3GdNKSIeieYvTd7o0O/qlEQ1tIsipxOm2HEqxjIVuCrF0tXKo7xKXcwMk68c
4jqYR5oscwKNhGpJrOWxLt5X6auJBIDxau8fuULaJDhq5yuCUhG+D/VnqJq0APh5WPg1pvvNkCn9
RQHDcbfcw4cOZ3G/0IDYY7qClap/A/FCtPAqg7hUtrF5Sk6SRE4Kjnk5K/BNrMB611lCEUWHt7WM
g8klCp/TJFnYLKa0sFLPTSNv84hWgPVRPEGyltgSAYumEQsfXBT7Db/hZYl3wmAJzmVHe94YWzMg
uQl/wmvLgZrNj/i7RcYYJE02dX+iU3JgkFR/pq0YpB8cPr/BNkn036fxhA+AFh79E0UuCcSDYjTK
QaZXVXic8uc4waYzQRpzaptDt3OrCqp0aof8E7J5Tov4IOUtZ4Gcn3licXrT/voMYEBqBlkifBFJ
vPKTcDBodQoi15ihPmEEv3IV9Flm8ity1y0QsJluDNdDl6T194VLPXvkAPtuaNIy9mykz8GRKTrr
oqHL8oH3B8cJdHVTWpSHaaldhmkjaW715uGKU45sccM3EVXoy9uLMfGEGLXVHNfdZnjNbtI6eVJc
zWJhuFseHs2gWKNfAalWtRZjwFqYPEMIFFg+QfIkav54zNr542yH0jPo7C4zBFnM9tLr4g58QAkx
e7z74ajw6fnqOXaDEnHLLEGlbuY+sXIgGbskw2t3dP2VFMIQw6h1xHzMczqigv706Yhu+7x8oeAx
DFM1cua6L/IuNxjQxNl/MMAJl0/WmITyy/5NsLnFOzNAkkvF58pBUw1XphqXcOITQrg6PrMsxCk1
B1iqV0hdFYkG0pBn5QMrCBP0VKt4+8T0dw8GuUlE11rueJMyQjSaVRu36rMTTeYAkoH3rWqS1s8m
2UB9fTxf1R2Pdzp+sTrUmj7iDC2PJEtXo5D/WbWmBi1P7hgdt9nFjQKDaiKQiq4DAEOnz1JwyOvv
4H1IHAJFP3FSqshfAYsZqgsU/0UCCCmSLUZ3vF8W6vcXDZJvMh11ekkxIr7mjNZqRzKLMuSzZZ6K
XPKtSP4rSaYbF0jXVH5LQwY0VW2l3fZp+nRy2fcQ6Npa9DK8n33nFnvMKGV8NH9EOLEHxc51UBW8
CyOGabnrj+7y/Pqvr2E4c7paw1wHn5LBKefMvAgn3a0UvPye7MvEkP1G1ppB5ja0m1nLvZ4jF1gf
goZiGewZfLL2HJQ9DGxN6jjKGlZTHYhH+CqPAfbBk6K21iqz5RqXsAEtnMQcVGXSpC36P7dweViX
YdC+7yz/kOnmyAJr+J2koTa3WDIsyajcm4WbIgR0bSPkQ1qVOEOZh1ukDfg4xHnQRahxcq30hfHb
1CwJHvlzvmH0xMj9A2bS6zYpz5iiWSOehl6ZTuJW0kuMmsKaN+FsHO5GZsUF7u5ywBWjpPortod3
vn+Vppax3UcuSaheLaWyUGx7/+u2Zn3HRqFE4EQ0td3SZ8p0mHcauY0ru9/4t+Az1sPo8vawlKYi
dCT/Mky74ZojPpAHXjQSLn6YULvSa0vmOl5A9m5qXzLDsnjvrRExVSbWnQ/3c4Hbb5tQiALKp+6T
lTMS3vwhnJlzdu8gr9sba4xnPmdzAGtkyn2bL+HgTukqyn6ao29u3u8Oc8dBaPGlICTKD5khTA27
fnVYOYut/29ChW7gC7ada9PN11FSRTBxl9gqUXeLO0L+XbRfuowlEZ+I1vPpRMa6kJZUoEsZLDj8
gBuMydZQZnxNY/q+yt+SRhtL74KOPZvGEzIK+gwmEl05xd8Lto8+bkaPJWGlj3pmRyB2JGUeCPRU
N7857RG/CHDP+LJsIUq+Li+tHInhvdKT2w6C6NvLjdJUWPnU9yopfsZNpUYhSMthYmtSn3kUATz0
n6mt6NQTzzPYC/0SFFW3rOtJYMo6NWskL2vM+6uBMZ7SAlBLAgBQkyjMu04gi4pqRPjcTHkYU5Z7
GQ1GNrAiknMMXyymYyjAd3T6LS0/9Kn8QVR6EkMUbQ7PdSAIBGXFWYJTPTPmhEgQMHk9ncwCrXY4
CkmQdX8Jt1KT1PmQSl5u6HL8VmR/7mK4EdBmQanXur0gQ2nVXRVCFryU2yzT4msI2i2BrLRryPKk
VwbGmQ7mxcGwRZvHb3SpvWvavgSNOhyE2y/na78c9FjUujxMJSPUTMWz33FkU52YanueVQKeo8Rm
WMD+ln0eSvDqorA5jltsVfdwXKf8eIzw54gojbkl/C0eMzF1oCJjG2Z3nL+lHIyP07IvfDVOKRen
VTClaPgzIb1tO9kEoohU3jebj8sMY17q5Q+vl2ArkMorL+kDKf97kTmuEZTb84i5CEniwlgq9dBn
/s3VBKG/2Omoncw2MEhh3F1QWX7/tz2oxZm1AO7VYmZ/Vdc57ox21buUPkOPOcu4hldjNQEWEcXp
+nJJ1RAm2dmSEeeBiUaMM6UpnM6clGF64o5iC2kJ0fsdxRfZSgO2bh2vone8KAJ+tMpexgGzpQQv
6Lg6o2BaA9w/5QgdDO/05I0jBxZWQu+hmW5SD7HjWS3USknVrqeWhSw44sNtaMEnPD7HsENyTKKX
kUwVVTnFDFmhvafD9DdbOq+kfHUwD4lwJDH0d7LrRlQLye7GC0qEDS4ICBboyCDxpXEW5wPxCqID
qBooMD4nQaG+ZejuEua25tu3NP8iXMMdIR55aGKcxEqXn43Q01AG5qV6XaCDa1aAgwDinuHE1/Ln
jwstIL9z7om8cBg6jJy+Hkoo2C3YJwjZasVgZSBoJTN/eEkb+uyI7jZUcbl1CQ7/sQl+3e7vfB5a
8yA1hrKHXEe7v021Hky635znlnYEYWvWpsmpx9dROIre/eDR/bE3yIfAtjVV8DEMm9xso3FjptA5
n1mwERMTak95VguzUpu1FIC5F7MhTbwkuuWQOTqrN9laP5X3k1hxiiChduOuuAAI7W1DxirOTXYf
su+EpQo8IhvB0p9oi7mdJxvMD6jJKQmKDdRbloYkM8aTaQLbIDxk+4K+ipS/6cVqMI6PU3sxWNzi
GP9F/HkgW3jP3GZPl2PxYA47kZo/sO87dNMPMx1Xn5NNJGVLXSiGbLHTCM7z9zkTGMp9PeCWMcol
RrGO5y0SVxBmfbhdtCppFSTolI/OdejcLSHmj3r1jA5h/m2HhuNqx1G28Ryo3UrT3QEHhzFwzzGy
9pMPcFy4VLqjgN5X6HFf5rY5nOv5LcSVhUZt7nEwWTYXlz4A0WauHGP22x46fAtswCyMsYGCea6S
Z2rcrjeS5nL+0drh/948dIf8GLyRQHcNvCU/H+w7s6s8pwfwr5mJYFZZxIyymAc/VeZvunzB6qpk
5ujFLXUAheCc+3wgT5tOkbwNzzvolBfjnMXbvwotyY80NjJPePDT/Eg0UOscjW1qxM3yh2C62bSD
z7mUnK0hlOt1FU+NdxLfeA/9LjTyuLsM9DbUPE4XHbF3l+4aJ5xa125Cxm0oo5usvy3l1d8stFcM
bacFFeum9JHNbxTv7q234AY6bdTH5Oynm85CV3yx+KFbFwRrOOWtzB9+L0Q7RmOQ2OsRZEmJggOA
lIp+XOMIpYI2zplz1hKHZ4puoLoslyDF2wyu32hoXnIkWNv7MmPuz+xcotReEfJQlYktGalA2Mmc
ckvLonCVBBEuwBdQKGr9K3Xl79HNlnzxlTjbsK1vo7x+8vZH92vZoSN9okQ3ZbDtpOFU4LtwjlP1
81U51P7V7OEkxWUS03IEB9WvRm9cym/zTFiASSp+fOxwXCQntch7J5rElAZ40gCZQ7EckR4Kuqwj
9OeqtnxQZQmwKyzy6D1OUSxloQxe7TSmYzRbQGCdjKUm3jxlJcMPm46VsUVUSMy/wG19P4IVEr2e
xeqynVC3mnmY0FMWqyZv/KGN1ur87EoH1WmJqTixPcq2LxjbnKYU7ljDx7gy/8l7C/kb6M8M+XAh
Hr5GaMnUr3vA5YQVG9g/TFhV7BXeXTWsPxlrXl77+ZfKbxvedep9bGD3IsO8BPCP52vvFUBW0+EP
+vHzJHTt13l+e4r30K9EAp76gstMDHciVSGhYYt4+CNkhLO/619pnyUYJXolH5Cu2riGVgezfr8s
3jZZPEkvS2JNubCaekOVeSDgj097kU4BF6sJ+GXNjEiPUPbNEuN83bdQYB2cgZR1kWj/QLzjk/2W
vvClHalsLcoZMfnHXiJNbUg11uXqosLrUG8nnNDhRCcVQOD3egX380sfCd0bkkbC1f5XnWryYof7
6KQiqKkOWue0PWLO7CvhSixK0GLAxsQBw2ujwXqxfkwRtZMBG40K8bOWHsnv6YgnGvtOei0ZgAQ4
JC4a5ucp7JCrBlp+f2NL30CyvW/IrPea8ygrDP6Q6yf9lKbrgbTayhiBEahC3z4dVAzVGkiof12U
1MDpaNCCOTHo0TH4Q9PgbtDgPe9DOZHR516dAh93SR2nze9fSq2x0rcTXjNonDuLcGwHVLim9ZnE
PGsQGYCNRMTKBDygA2R4oirfMSLRcXI/untfQO84m5FyfBWu9h+LL75PEqibqkYKB+Da41NWWCxl
P5a7hRsZedk1SrT20DYXcM+mT15/E/erx241aX3wWnfLBYvt5JpupW5hFgHNAcpPhnz0YQAwDrYN
RphjEjzTYmKd6NM6LPdUoHrpmM5tvfsSW76PEzdlOA41DWv2MxZYRX7Y5bx9Vffg3avZGPP0y04d
pgbDaxzF7Zbp23pDM9Y/CLqfcr79rM7buJfs+wf5Ao3Qjkso45yfFE0c1+yX2szdT6iEVtqae6c0
hK7RxkLD4+CdpUnNlXK8pojWGxbBEe9VJzQ0IZ3oo2BNp8BXhFcR2XY80q8yXz0/ihF9yalcQLge
hNLd6EWwHZ9WraWNQn0Y2PrnM1fOmy55gLx3+E7/lYqnlDx0SCUYvRXoe+/uhquDuhMqoROHNnW6
RHnGLfmg3Sjix9hg+4N1AbaKU38TVLFvqbAFu55YAvO0bFZc1KB75eJ7KyZGT2XrqLOFRqfh3/E7
fcRVyoI9MDUi9qEfwmzBvolmnJmnhqryV1WLqb9s4dkrQ2ictsBsLKX+OlB/L6JUDts/PsQw15Il
ca0nz7oS6ZmUnJCmLTJMcgPjINekDO72WsI/M5yFVZZjSFpiXy84fM7nP2+jDYm/vmqzqUfFD2Ja
yCj90wIqkJFZTnMI0014c9izI6zpbFTxjyu45vw0nyAT2N+ejnNgi4T5obXcjDZ3otQUSG3B11hj
DSz8ryYYjIbHsZ41ZuVWRDjAfgLbwh7KJ0/6bCeceqV96nksA7zGVU2uT+UxWiF07wZL2v0i99wA
kyOwbxjgtpxanb8BQm5BaXR7pbrf6Qxcoyc16QpOw95Sxq1HrYvaDyPspG6DKmFM+/Hu0tmsltTE
6BTxBu7yCV8KE9Pedz716mPp5ufycqtYsaddeH5nD/fcR3kxCwnMukvPJpGs7tC7yU/KTmWaIbgs
CH01Ut19rRl61QxDRg+qB7nTnBg8IfS+LybPzDHkhYXuVgxIctcG0qvCIbmq+0TCfX5AODTxKAzY
n6O2VKuJtr/gRFsv8mfDpRgThix8N/hPVjKbyilck0VA0wH2eOYBfWIC3q6Uz0VoB5tjiQLH6kDF
bF1jMqgKVpqgfC0NeR5K6nJXgvimhylBUvYYXAtBFMGSi1PHjEkCoxWBjy275aebgZ9reH0ivD4Q
jC4PU4v3oHrkmSqUAQ/OqNEVr0VUUlfvTv4opuAgOA6C0vjc5K/QrQRhsikbAHVQJkVSzLj8GUeO
dPfc+QVtnoiR89qVQ/zHU5c5pVPdCIVePclE6fbsiQ4swGk9LFxG0gLQxEexcm0v4w6bHIq+haO6
GXOv5uQNgKSq/wrm2zegBQYz9UORxc7+VBNxgygwf4zuvGhLtBagmUeI+ept6zrfR6rDAdtIPMMX
iqteTW/MqFrL/psWLX3BXGA8G0PsxG3rDi0uNL7864zT5Vkgm/6HhVnpgyKIw2BWYbYiEB04eqVj
MU0OpcV7jICxMvVDrWJjkb3+pe+zn27bWsOJZ42A1dl4Toi97sUheMTtCZ/L6bkKm1GlcgAAOIyU
b775BPk60BZjl34TnXH6kgpFUGn11V2D4S/5yx3RfG487l5smimypUqOMk4o/avlz4DP4/kWcI8N
nnaVPiMW5cPYtPQ/0rFzQNVZNIQjib/WdTVFQNsVS9UB/lGJVhYYhKG5/LPF8ppGLoqWkt/aCdkT
0wuA7rJufyk/ZISrqbTKQIVVeedy2drHNoWKLdEuSKftRXmXGDeesiRMe6X8K3IivokKRiin+b5i
Puy9RkZfCL7bB6UThXekedVQe0tm/embN+VQKB/vnc8wrfkeF5bF5sT2jNZ5LMJa0SUf4MsBLcQ0
7Ep1P6qLQ6wNVhbNvzb3OF341t0YZm3gby/+VKTZ0/N4Wf0fPWj4qiW6ZeB7Y4fiEWAt6KXgQEhX
WFKdD0ffPDmhpJbwlL8AJ05kyTrj+9BH9WTZVbXvYpQxR3KuLUtyah/8bgOAVlVlYIbNrBXS8RkA
gFmU7/EKURpk8MMexZoPdwj7FXIhvtcQEIMuHOj21WEAkaw7D5MfdZ7XBBr/LR9W50AR3Kh3mkoO
YA5R2ymKtmZyAhAqpRO1/ViwRt6JUereaaS2pHim3yOl7wx55gF/o+Tg8bMLGoJAvCA+XbFroRDQ
FIghl2TCZIhQmcwcU7bmUbhiiUMSbvg0UPoMYk1R1v28Mj74Ld0zKrD4zu4FkTHuru9j7rri+gex
xvteXZWK9dbma2PgeL3/Awf69ylZlItfn+Sf5be2F1q6j2fOHxmUMTtfiz2YUIrFVmovov5I1vST
3HdaLELQZFHS80m2VKdAhGOjm31YlzYa2JmyHfxg21rM3WdAyV66S6GiVs7fBAYXmetZ0qLD4Z+2
xb3Pj9RPc9xTzLcoV3RWPX5KRFGZeUm/2ICBZgwGdaNm07PKM7dyV2XxFDzENYsfo6QEsBV3aUdy
zjoSFmNW5i26OSN8l/sIj66pJ4q/NsaDlEKwAvulciJuYyb9LiqUBIyYc4cFI/zO3509a3R0EFGD
zSKi9O8asLGZ3usqhVMc/s8ZHgTckMtjC1pR9Z9YZa7ddrjSpv0p07G/UIh+z8vnKEPJdin/gov9
0QDAjHT/Ypsphh5rqcD4UUhUvuAT9rXKOTWXmM5w61lnMtiVPnYnO/QtQxBn1Vd5tgs9T9ro7quL
zk/2eG1bGuGsOYHNBMqSKI8Ul4oP3fFu97T3Sb54PvJm9Helmldp/wsFMzyLYGocQ2CLJ8KfuuZY
Pr3+8GXaQQLdDarEh+c0drVZi35vp+w2JAkGt/FuH1eSu1GHBj+Wj/NW0d9sdBuEaIJXDpxQ5XUG
XYzP3XYGTnYR+Bh+h1m3xt8ZudHJf76btUXxv+P3m7zm3gE7E8O1OaJuhNo+fY557QHYvm/LbtiI
hrepOkmCxBTCEB2q/a5v+naZ7y4JsnuSs0GGqnOsgvs6R/LK+B0r/wjrHM6v46PA2BqweWU/k6eG
lgqaldkKfpZ6tUUKu6PrplySc965O0UsnqbR99hknEnvJ5cVqqDh25HESQueHVyF+PnHmSP+BC2m
hknyIrE382BlkgsQRXNSK2ES5V5B0eesyo9P2pgl9K/4rebhzYZR6osQRnJOTD9v0J2FQQOxCDUm
BQM/myeSbnxUK8flQkud8hcBTO0Aanok5TklPO1dDp1JWOHkZyeSEN1veyHYEKBZHqBzi3TBNJhZ
phCuLo5DmFZvWQt4WlHoZAC4TQCqukBPd+LM4LR5T05CSuu2Pi/FrGhzW1tnVdOviPKrygoN1OyU
qQfysr0+TfvcDy0ar7HDlU7wAZbhJD8fkNFDkxyAUbOa9yHehDWrmoluoZY1gOPFDtxM70rTE4z4
XTDU2ev27dLT8eM0spSNGprcUYvYhYrdG2pROP7rPAo1SLe3KOsJ01mPSUzHB1+1kKJYC2Bexq76
91C+Rc5Nj+IIHBQZ5lyqZ2ynDc8/5Mf5eQ7uDtRwB+gtIe9eMjXcwr7O5E6JcCJKaKeBM1BS4NJU
B7aq5UP/SFbnVVFmfwqQCuum6TzxZARJPLJQ3nh2fTRA/AaOrdKU1blZIscEQBhso8jslaOxjEtc
764fY5T6FZATx08RMYqH1gKxRE0qFBtfwCyVv5rM5EdvPyzbu+4tVSskDNOmLC0oP6SCSwZHt05U
VEiFTPdvAg7ICuTZaLakFI9XKy8REzD0FO+d3CAoiXt9LfYo7GcaswA+FfXS62WLiH/BjPZTNEy9
MZSadCXgUFjOLK4CsuNWCZhcr1fUO+Vgej36Zdo7QVu12liTMEiTrrShbz0zSU/Zs1d034EcbxcI
jquT1N3vlOV89OVehaKPWTgz5mf/6Hmykn5maC+C6ap/7jylt7djGK0gQz3TDMUpbbqMaE09ESkJ
uJqE9lCwXJihopKqU+HEhSzGwa58+X7UmnucIJy/5wo9hgiUamZPuJbVXX8jPbrbL3irLuuj+pmE
sooCRYgKeCTxJieA6laqAytDIQZy1bVtfylkh3fCMHl36y1q3Lok7SljsdjzHL7Z8IgCUrso8xLM
ULbxQcAUvBIePLIJnhLUZrl3BpxIqmfyEYGJQdyKmcU5DpOf7VU7fu0sPtRaSdIztRSzSIm2XlHH
IeaB7JVvHdPm5mTeuWOMTmuArxdRd5TbNy9CXAMe+ct+RI1paY3wHWQ45SqZV2kNzKYZVIs+hxqN
PdU0GPLNyo0+4VTBL0Shn5wkfnSxqMBox9rJEGoyQ0d65O8SPPmgzpp0Q6d7EF5wF0BdYbkchLy6
SN/mptpYuKWS5cYug8jwqYgJpNET2gEFKDB4Tu2m1wKK6IXaCBizKnABOgCeBIatYOzbjWCupWQl
mlC4S9ybTQ63jSpSMtdzUBiTzvN5MTGV0iLLdGOOk9lmsNjJmEs990BvSMf1eN1VnA6RJYBVyl6+
IvFPAGHfU4XSWV9jJUpclkWjf/XVgLuYC0mbx0FOLD5cYLtyJCV0r8gnJlwn0IlyjpdpTkhIxyfY
z6rDOZJ1eu3zsFv14JYh0UAZvWZcEnirgrauFfcmVEAmO2tqlcvSzFw0mZorJOd4u1/KbSjkvfyF
5YNTRMaP+qJyqcneBIiehJRsq92G+ivPNPfHxTnOey4DJxTg1uuYZZMPxg8Fw/I5QloehZaaODTz
tt1Q5DzX6nzQJxCtUIOSNc7oJwUuYG36LZQ3L61+s0A8/OCnGypvppjdFlloEn6V4K4SYPrx7BrX
kRccyQxF2FdtvHxuzNvsxzjRzpN1O3zLmk6U4NsoNI1oSE4Z6Z0IXat3s+g8kH82CB6LEAkBqwMo
7zh6k17VL8PcMYejzDbj4rXjdOZ3i0Td//FBMVXl5va9C8Y39TuKWAf6MQej4XqfAIx95P1/zP01
qpRKhIvK11WsrdsdHdiWkBjBWl03L2L2CQyxr4RpUHOQsr0x1gqswfhGYNgIVyn82zpjm6r1dYks
gvt+gRJzeXbhJDe+XcIJsRf56MACbGbxQ/hr6CLIJZUmG9Y3Kz3g2HLPK2BHGGunVlB88j19CPPl
YJ6n3q4sEy4vRgRA/Cc0jvMXSNgWq6VnDkX7wkDPHIu7d3FioxYqNfH+rt/SqeufoKOvDlm94As9
z7PjZeaOWh7+DHEVIwRp55uQW2gf1q1gC6cHsdXZlJnZDVgtfGB/EDKKxFEQ36YXwgPrMHKsHi/M
iuMGOKe25r11cTcj9R+MTShZf93bWD364WGFJBCbcj4jKGBp0v40lSkQ/VBt7Nd1NbIf6hGG1cVM
D0ikHrJ3S3faaJLNw+Rma1pjwELtk+ugK2ZzHW6ZwxpGg8eAw3I0hdryPHF/t4Fv7b0o3gUWWOb2
Rv150cyeyfoikKxcpijkvKA34oLWZceHGiLM5Acuozo+qTWmJIhxftkhJIX2veWsA/8a4eymLibm
oR29ZcyDjk7rt2jgiRZRPmgrJtS5hMMTrtjX45Wcnhb9uhlMV9B9pyKo1GQA+B2AZQR2ljbnVU+E
Z6whDHIqMaSyPqfnmNC43iEkc1JnRK6wvLfRnCHDC51b7AoPryb7is8SrxD+ec/Cods24AKNtWAr
yoIfVuSUnTw/lTYiG6Gwf7kKkra9iTBSzC8EIOd8NrI0NwYBXOtF0Gkz2BaqJNVR728/mq3tJMyF
4RwkOgc3oj5X8qWnwPOcDMuy9/wqG7BeyG2zXQvCf0yKSRzGh/D1IqtW3s6ZYOKbvURjF2fC+Xb3
zfIWrkrcG293N1khAgT7LxYh10ErXkS6VVomdC0k1Ajn/lm6UUh9b6wEyvfccAVqpcvRLPk/c/7m
kK2PUazlDAFpi7YhmNfXtY91wjRzHpKgJthWeoh/F4xnmEmQ/7t/FYP6vbmIALyDo/2ahDyTomQk
5xKZO8N9w+TqA2UiRDoSdMdZCiGZm2l8mwdfexZSsh4/yHSe8JqthXOPf9NruKrV45ad0s7PPe+Y
kPGpygXGyH4MwC8qn8/bicSo8VFA8iHQW2hygxTIZBX5QoAx/vf/lRGPzU+PKyfaCOHlZXXfCdQd
RKmy6sDtkQRoRZF9MJfKohwJhaitC+/AAZAPs9Cz61knCdLZLVRteGXlSZKwrVQXkcfHL/tXkEiU
PZWxQYfJ5L3bB/MiF5V5P5YvLYFF06at6Uxlg9yQtdz1r8FtsGocqwtpRibjPBmAwR2ORpmydUdg
MfLm2L8w88ESmz5e/FLkR6+Q3cSgj23tI7nnlRFjzpQ/eTPNMmtoSc7V4KdgfSltewjluDpAZElA
kQQ4fyA4Xu/n18Rqar9QcQhN09U2zP7auLoRCsDvOuXprMztp5MhsBLjGhID81jAsdnDtGTr7pT5
U3PklqbrHL7c0b6JjEbPnHDjQkDn7+VSIPfbROnKfL70V8NdmhToIIkf41F0Sjxwiwd95HobugMf
tsdzlJPCiREQJeCXmPHyjMmnkQSgBc4iYU71ZTcfFIxkkpUswgQkmza5tCtjFFNoUoJzbOBX1MGK
ZXHEPiBiUXeZc0ZrdlGic4vc964vsT6Xeq57YR0ZSb9/MFJa66cyEFgJPPTNgwFE7lgvZFjCNx2Y
i9hw1H1MzyU2rBi6FwCDV1ry4pv6kwgWtjdnYDrEglIhztaDx2GUW9CORBKgEiWkdcamKC6W2iTw
hiWvMAKfDpDmx97niQpZbgMkw17ks/yiZ7X1sNOBO79k1I+E473srlJMjfPvxERLxKrm38fcJyLj
24KntGHhRXfF72xrhqPA1UoR/hzv75H/HNtzxvYR5/02gDzymuP/uWG8XI8dE+DkpQ9ASE4KMlM3
CpAXJziN4Wig58OEQSi9wV3fiS8ww3ysvg/WP+rJAt1ZO7MBt2IvwOUGa71d5dA0hPsM/jtW/wxt
MHWWUNiwDudWb8Clr11naIqR5xhYwgF+DDjysZlxdpD6BWSGFAFtcF0p6zKVVN29qMoFf2WBDpoQ
jCWWAbq2BlZGFq/kC40TvXU6F63XAzz8cmaPvsUMk7VqwGEXgO9+VBIP/FV91IipG1XlT8ErkbEt
hthuF+bhoEkMDnpavrWJ/jUnLqGZqk6kxDZw7Z2hSS10DE68qBaAgQg6pcDIUyDsdiag+ZkB81E4
Yinzawo44fLAfj4n11NynIxFFASfW1J6mzNv1p45MVhfR0R+0eW/rpvD/H9Vtz+2hJpEuhVUCJEP
LNL+ikloEV6JbxjaUjyNMkb3uBTQaNXor4cghBPd+sqgikWna207PgsbZPjTlzVrO5ZFtQpAQbSY
xjrYlccEiAXAfydPDkf1eDhVv0sK6+Jy64MvHnPxRZoYMuBIijfxiZ8234B4JL8WvwU02EYbLLpQ
bBoTEHtOlIt+SDr1F4W8w4gL
`protect end_protected
