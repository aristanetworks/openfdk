--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
iMN1kZAKVdqXPEADwwMQfpoKHBTVVdAV459fKdDdXzJvXQR/YpO4e99jwEAMIhQ25ac9/JxBIrY8
KpsSqwzggAu+i1hhcOpNq6vl7/STzbuVdYBQichbU7rnpmlpuSAUc2yIqv5ZAIrNHXxSIC6eF0IZ
OO/Fabs1c+6fyUtTwzjxJaR5eENf/nmdlxAhYPAd/aQqimBIbFCoG5wdOEcVwrbmsmW2DQW8ap+v
6Bhx9Pp9EfNBGO5JAm+DAjG8tJz8g3yOEGuxp4JJarrna4DoiZoTlPFv2sxRKOop1qbCHPdgPWgN
gieuBMbKOyFA+Z4SuLDqzUvT2Ne6n7RfSUFLYg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="D4ReQEoZJE7+8EdGTX4TZK5pHiig6M2F8wVq/eSZfKc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
QFESIuUxV/Tmfr6vhnRMBiy67JTgW5WZUAHWN/a3t4RU5tEYa41uR1U31PqwlO+7SYuAdo3ylsfx
S0e5240N7XAQGCdMH3aD9WFuZjNcXRS7PwIsFI15Xt/B7q7bhGeaIPlgffIuUB2QdUyHmnA0ZxVp
VizBwFwB4HYvNDhvNwPBNQBs2N/fTJpYD191Wm0WDtuCHOSNH2G8qZ3/Z7TIaIQIzPGn7/7uWQQd
wsNJqR8lbThE+IvAmr1h6h0+vM/poZSI9nymeqUzAEKfqSbwsYtviFNoQaiyGw6vMRX13STcMhWm
E0E2c8oSr1jFCh2aFOsQ6qPrv861J7seKhRArw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Zbxhg/ZsjwEtcJ5uCxvFo89AUlolXj6p6KxxiEUGNUU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26400)
`protect data_block
/MWoMbn9VeUp8mfnTNZV8nhlstS+5coUYHF17MInd+6aqdS8PuUGb/6+/2ui0INCRXbCPJew00RR
xPxRqmxltcRShRhiixsAM6A5VDoDwy+FKxCg/0XRS0A2v2Eraza00HOhZLg+nadVk22G6cqF/uOY
9pwTAdoxweWzfPs4HhAN4XibJxM7ICnbpEpNZeO8C8wNZFOCsqLS13aiX7klPe4lik1lfWrqFaRu
A8h/v4LxAD32oQ/9WfeoPXFffJHihINcIRMYp60zx6NOPki4zsZR4LPl+N8+UgAnOuJuJ5wxiR+6
iE+g/WYTzlBb5dLPUg6IJqLZmgiK2U3y9J2lnCJ4wcNCxE596iIi1R8lja6kgpnJREutnSfps0xu
pEgl7mnCjlvoZrT6ZrpzmDifo3SNhDIziC3hpa1ekn09OVTOYRVJfiNWA9eSfzAeAsWRvI/fF9HU
0qJSe2CTaTZh1psf+D4ZiLGWQHY/UsE1LWndp+Kxm3roq6k6NhAzf5LLFtfoh+snGz+T54SNGaZo
ZyfMwHFN5aT/XjiZqv81O3sqyW2scWXuEpTp5lXclzPEJa4jjltozTIqZx/1hfc3h+PCrMNF0hh/
CRZK2UYXsgeZxWw16qXQ4F8MNxsU6Oiq/X49B+pLPyj0KVJ3za8kY+ppMLH07uuPpLuKDCveBLvQ
bApg80cD9oBoOMEC0eQiji+rCTum1qQ9hpH7JvnWJA/uuVOkn2+V+76srJrOgATIv7V2xVw6CFyE
NprkfpI1ADBuXLtS7jdSwG2I1WEM7q38NdUGHQBVRx5dYwJlxQDhkyaN4UcdJJ7PW8jDtOSWKdQP
p5XZBdY7fjW9QoAkE4jLnHgBjtmr4+jUr8lnR+XMzM6uCIPTk9tiiLHZF/s5DRpRz6UQWUqcpaE8
IiU5a/5iZmJitmSMhBAMnhZ5b2nwrNPP9p4Y0kY0tGr3iUa27hISoqKw3Ne6V/CK08IiooxsBQIG
SU3S1OgPFYAdcrKbL+6IVL4TV7ocL4kfwQhZq7CsWaThlB/hLsWfZU6gN2RVFgi89GEkYPLDcy/C
EsYHMMU3mk4pxUgF74A9vMFwHjUmgtjjqhagL6VIcQUgmeHF0XXyDXW9KRSbFNFbSpGt2Dk7YXAg
xw5gwdn5TnXIZ1j0PowsX2glYnVgzDJLS8ZRsZ9U/phhxHJRwg4T/p+BQarIDxYruN47+VxDG+lB
XDvi9TqWDbJSAwOV0mT+sXesm5K8rS+LRV3MAaShTWcTRK9IGw6EcS5SSuil/rL16rnIZeO5wrT+
qJrNH4sjRcOpVxmmy/GQwB5EclLxXhmq62hqeAV3NRBS9KD/mPmEi+PErxSlzmHWA55SPCK5e0AO
WU3TnhzrWgEpeTVrlbY6/AzULpdfph6JeBSz0bAvZphIyP+ABE20C+3A4idhHnY5u/tnW4oThEVN
+JAQolRSokPAnhkKSgR7yTxMnl+M7vQVjAUK1G1JvUEP1LzVORhbFnDEbTAFHUdwSwJibYVnRRWA
1y0T+hPC/vDIB2IvckzOKkZu7lFS/+YvROqu1bp1nlD/7BL0cR2heE9Ki1iyL04p/POLaPXma/gC
9tMKvSXWZt9z0XyAQj1W0bxujaaoKzdkuoHvkW/RSdth0KCqoGK/WRo1ynDr7wm0eoVitpu/w6qQ
QwJNPZajhieaxebuVFIMCaoqccFSJ7Z5cUnNkj0ua4sIARcAFvJETkfIN5aeE5ZZfnAomiqjm/u9
jKPBHvk/MZ9JBDAPYcgqkmKhnJEdZ6UEB5MEnAHw7OpVFm4Ch3+E6Vqcsv7c1bNJevxnMpoGI4Ik
2ZZEO/Gie34vJVOvcanW+FBPq0o50Exj4qynY2+4GUpAQwXur390dpLpP7yn89XOXvnlLBSOuf33
+VAXMyuJuka7ySVmvFkjVnyHIavqyDjBRRsrHHiQV32n3z/QZgC/OmASB4gkrpzvG6P7AbTYDAR3
gkdyfR5j9Jjzjj0OqP/ddzEhand5pIAHILJXCO9Ng1VSqEuqrAXUY9O750Oe6P1Qz5sDWHmIgz4B
kYtMJ4PJe2SsRbhiezFemIR62hRDEqaMqABrS1hOMNu4OrBoTKanh8i0aPMm6OpmlTrNDlbCO5KP
TDlHrhEV+Sf+T4FZVXimDbt4RGFdrHU+SdeaQN4H7/E1pW8nIodhkUvV44jd6l/ug2FYOx/kPZWx
hDpOaqa+TK/mcWRWDB/upAV1raPC05irwLqFSZELWl7mUgfTe5tla1TD5r8dXeW0oaljQaNt/qla
mx5mxvf2j9qE0hsIJ88FqwuGc4Wq3tLgDuqPD9txlWnukoT3hrpLBqUiTq7RWTcA95ZxJ/3msad3
Ltf4K5YYd5aDIr0xoFKDVor6dasGcJdNt4LAOX7RNIWa82r2f2JMjVHw41LwpUV/3BZJte+3C73u
IqP4EtginkTwsUPmtdAogyoYxOwtIP+p89uSDU0MmZBFMaPyWlnKozOnttprhHaAC5c0pygl/ci2
94ZgaTE2fwms9BOpoFd3+Gmc1AzrpwEd2IEyws8D83gkDE2W7TkvCcxpNXcj6HLvkSdyyvL8S45U
jrezT9q/HVKDniXTCZXtJlk2M6h8CT3XSCxYU4mCNY9v4tE/vKMdhEAeG/RAsHHD+gpO05ybKtIQ
wn3t5DMnTeVQvQTDqavXL3Ys26gsaPMx31ivpPAt7pyJ0wfAeAiDJENlY+6TmwBG/kd4xCiVfh8c
umJBjZ22898wolGxjywarB9EJzCiMKAe9K2LptepZcnSwQh41JhcgVgtT330CNNndCr4zCNdUYLL
maC+oqPk2emX7BurUrLRNuxk4bFuDu6EsXgRcqquBrLJ3mzvbqxwkVVGiJFqwwnwcQD7HrTXHaVE
GpUd19DPgdeCG4BQxv38790t3+Rq985qqL8KVAZDmmY8NlmS1btNWXb4JkrnXeE++EfhkizmYDYU
pn9n0bDxI0bl55/APfj2SquZgJcb3AWpcIt1lOcEf+pkyk8NinGJtAJOjptu0Bvp1unwyYaGWbxg
waQEFv+4VT2qnQ+TSOTL+eWe8//9RKblnJlVHsevunZGWPjFxAqsfvM0MlQtzxv4C4pIeKAlf7wI
c4CXCTWsMycvqLKklzgix5iBuTkCLEgQljZMV5Rpu8HbmnpGOTmzetK40oiZ4CJqFsz0bYy0ksiQ
B/tmD3s58WJmjyVmy8KRcyUfwy6l2QtC0hIZYWGCWjR4AVLnpKKmjnX3PYlNN/Rhdd5FqyaQ+++i
JValV7rwCn96FBSebVw1BWq3t6E6hxoEcB7Zd2WXSXi4NVh9cTOHH3Oo2zJTCc9RrMKeVosfZN2e
B8NHy7j9vAWlis0Qc7J2ZdpvYLJkumENgHjumkWl6X3iryPnscOvOPq1I+WaFOVg8oRjFvytr35R
2ZteJ98zaakoCZ6OMgr6zZ2BgVxucddQUUlZbvGdstIuxbh5rpzk6/NmpbuOrljLQgR3j620zgYL
KJHfjBMdCY43n/R9kuQHtbvPq+VGa5F/Nw7tF+Ix8JIPsVozChkI4Hs78eh2fM1iuvmQ0prqrBb5
h2jQdy13RuBBnaQmGAv7/tlgr1b+PqPiN0YzF/zQGQ7zabvouYHsszrmZpXFla8Fcjyik0P2THaW
cGsrxWv6a6savYmiTLDYAhJzlIF7fkdBJ/IEwSyFWt+nVQh3/q+rlRTu4y4XsPoAFA8BV+TvZdt5
tNaCjWKcESVh4esUCM1KFsUpyWViFqOu+RjHD9UZ8j8S6tV0yFwYHdJwTtxAWTr/iLXEowxDtmuX
jAC7BqHYEwhTXSmVCZUf2RmhNCUWr6LWl7ynSoI9oAAiVzPYNGDS0/xfEmCnmIWAYJSL2EmgOWEO
3gaRjj6DbgdtX6YKH8pVqAQ5OOXOnEtzwxjr4IvcAko7jcRHd2hQXXuv+XON6S8SzblIbOFc+9S5
FeLtFw0v98DnkHZU939V/jfbHqnK27nIJDqjzi81aq1HN/yj4U0nAS36EGXI2HQQx8TyWZ6HvJvd
NeAdmVnAQwNJIwbo1EN3TtC3q4F32oYFS9KBFb5r6zSiw03LQiPx545crs2kZdOWAKbeaRrOU8ZC
Ae7nZ20YCu1qAgZ3NqmJiO/FpfM7LFuSe4FnafNYvER2YaZY2bcukuu1BBZ5rF+dsgvO/17QwHHF
J/Qilx+zSNHNKFkI+TfioRQH0aCDFGjcarkLgZfHo9lXrInGJC6U6KcJObTlPxP54NjzgsxYnJU2
53Z2VqxptWfNT/IAj67tKGE6towBV69KRgm7gSA5wJIzh4usSgywa6aXOFswcGldDUfba+M/qU+F
IcRMbmIdxDfVvDWqWI+r3IydosWjqPXT7cSIZ/BwWVpuAG5vBbngUbBav/rNnyYxZ3ISTg+ueEIF
kAAH1UrpFfUR+pOAIFZcemZSj7k1VixYlObCvCXSZjaU6Ea9uRHKULYr3hrvMgMXtBQOaZ6GohNA
mi0BjehAwFBkv403c216YpKGAeZFSMz8/HAAMwupiGbD6IQO0F03Ah4AiYgBXWuQvAXeNXowNnzY
HtFBibKTFTZj9skEWZrbVLmv/hs5sNa3wQJeLkJ9xKIGF1D9DBkovqXQ3gMifcnz8OQNFlTEGM31
qfUzxiNNG8cTUk1A2iqyL46n9SR4z4P8OT3BftYkMpOkM3RjEMMleGF6cps1Xfa0aqoVxEhIFVDo
45wU/aKZeO1x4W7/1ZdrkilQkf8Cloclm7iUSOh+NOIaL/TrI674P3LOKOZv9ijolp+SquYDYtse
RqMwJQufsVzGhZyF8kNkfk5WxVS0ZlNcmR/IO2YCwE25BwO3bqL4NVFHeROKBewNw4qfR6XOcdtP
xtDLLmzEf63JqMJVB/VIDaG500Ka4JgP88pZgtXR+o8C7SvagdkWGpwq9ZO0fWDX95h5dMvroCJ+
1MQMP11d1COC2VDFHnsewdx/ykg3ioPCKwT8itBQHsY0C/0sSr/7C10+yk1N+7T7p07RBQQ16b+l
LL8l2KOgwIOeUxMgx7CeZouqyIfoRkyXAMaKVEnQzmhtBMIccDklMubYI3qFf7Ai2LexnSAjV+ef
hDKQPJ2ax3+jO8ymRFuVniNuiGrqZ03/OAnob/Kf1kpVjiMIXGVSi9cFhoQ0XfDAsH7y2IFa5SYF
eOVjpUnP/3Rse19BBT1g4JtbW5vtKRHmOoLTwPqOs2pZJz1L9iqDE3rdzqXu7tVtvs5/kmdBnYnf
5gCjpeyD5kPAA0H93ZyOcalfdeFwVaoex5Q5M1k4qKoyL2CAcgV3RtUp0NF+kKzVdCeAp8R0ipDB
6vhyOak3nXssmTvM2K9V7+sEDjaK/2n08Tkitf3dADaGymT4i3Iu9/i0WAA/QfTqUWydoxdM/JqP
Tn+nyTWncsEdfusNZjq/LBLjc71hWrC6fZusFiSkDQKTp2lUDEbpTIFl9FcCXwk9TclLBLkVasBx
OZlp1Fvum4TTQO4G1E7MmTiWhE3V1kwozIfCp5K+XXa0AUInu6cCcVMWfpgdTlUSBOpY4Qqss4AS
sMHPX2Jutzv/cQNeZwGlF9pLPCVYruQrDc+GT8NMoGFavFT6rvA0VDuvn8ic6rnVb5UFFl+DMI6s
pXPOlrJX4/mJ2r8MkFZMLat7UXUV//KoyUTSM/7F3xpNIw5CbstYnaoe8eEOgUmkj3GsPctsQ19K
qa7HQNuaAFd3mXvFRyueQg1oXzWh2qml/mQZFyNK+CDmxBhyZfHyz2+/60sbLlaOvxnyzkUKfoSj
0wtuM2YgKIfU/4z4UE4e49M+7npebh+2QCzoGaVBGRw4Ew3JvLmKo+52ZeBqMZ6wQe6XlXRIIfEx
hTAmsBMxvUiON16S4Az/2LTqJJN62n7Z6g1Fn6nK3Pqd8jCTSUXawJgQP9OtT3T95p0xrMh8PEaX
axhjMigdSUPOSmXsYApqJETvZNwbIFE+NQo3eyWwcWiKUDq1IYuQ0m/dv6WizX13ezwzRY0tFi8/
vN4T2OxfcXe4Jhc7ZmdPEskfaGVZvDy2NVXR+8UtviBIYkNSDjxdDvDzUrU60G+9cV3aPwD5FoSm
RpB0LCwGJSF52C7DAnOAOlO+hhkHP86PVlZmm+WVfkjiKU6zL2Qrrb8vErwDAc/AQpHLfp3J6tAW
4hxaB4Aqh7udBD2jc1Hr4+bQPk7DAFb4VVEFN0k5nguHrrtB0oMmlwJ8NDend2Ra/aFDtZbv1MmT
w9kilGQDlC3+vNvegPG6wXKG8SlOYn7ggM7LzEZeH0kWnOFlqZMnMMRLTLroq+gqhmu9tm+oAsj9
yysgZPMta6C0a3DMnfTzXWClW/Ggbg0puhXYEalKGnzlH24g2DNvlxcWapy/r1HJuz0cVlx8YGVP
/ViAxSNeivUP0O26V+BEP0hgznyHtu8YWzF7B22tsmboOYBOH5Z21KEHEKhOwsVAbDI67mQIlCJt
/J7UtXw2AzZkuyfYPWAfU1As05nBu73ppBTxSbzzg2b4Ra9HF+eatotkFYdwer9fAdVZLlDoSpOC
2YMrNouUCOo3SoOAM/XQMsCpn8Hg3kBoDZpXZ/RdLsAK48lrGE8ST5XQITwvX9PyBty7kRD0fBL/
r5lAzOFCdHsSko2IyGGzw5F/IONOWZXrw8Xa7SwGqQN/fbibhjY39n96JwKJtTKPGXgu+2eS5MFI
dk46BfcOW+4WxJUICBlxMv9wtw+8kTlYjGLg7pQjfTuZ0YipSP6jlpJbXMXCi8/9/9rwpXJMP3KS
8J0brgHfnsNwOGns3Qv82meH7SkZhau6bPEQvBmBO0kUk7Xp6G4jey/ePpZZon9FskXfjEOk3fLS
KWIZbaKCzVaEKIl5OCGtZmmv9f6lpfrW6WCp25Xt4N0Q80P2gnibY0+wn1WHx7P6K69TPlIor/xp
rMOVKo/zhHa9zm4HBKqVLJRYB9EVUvMCl/zl3GBO7KPdt9PTRWlmu+PIpU22LPQjLTTl2HMCbqKI
ryNzfN+sC4Tmuni4cXtcHvJ09K1+QMlU8bB7OtUCNHSQplqKIz9ERJv4WL1UFIhiWCwzOx3XvhAB
M4N4QC27Lrjn/xhLwbNTwvWWNX2zYNjpIY4IKMg2+xuOEU98rmm/S9oMUKhY3+/2XFjB9HFoblFN
Iq9ENyWRXlHg7KxhjA9APiKA9uFf8dGTtAb1KnPqSIQXUfMlzlwEO+8m0mthwq5k8LFC7xqEaV2p
k++6xpjfoYbWNlk0de7bi+fqmSH3vmaNtkx4usQA5Dzb4vCVNDuhDfZ+Wx8BZBxMM6IXVXI8nxB0
rTu6f71bIly9zSlhvaczMqZYQ1d+RIHhGb31BTHVxCvTgErjQ9lJS++ELD4f0GD8nt0ZAjK8XqcB
e8pVeD5/q/WR/e2c7sxffzTB58YiYeYwIYda9uYD9He42euvOQwX2N0nvg09tKamqIiGgSuETK7n
gmxfI+ynHEPv/e7D+aRQcUdO5r8q2eClqJ7hIxyGqMEWe5yy8NyWmLQQIg15QyGTlGzUJ8tahFK3
WRJErHmScqwlkTnZoZcuVLLn47AXkUSEIqpNOqHoBm+V315UGc89AbGXK06RN90jO7LQ95GkasoQ
RwZZC3c1Fu8H/O9vgUzRpgSigMwQcy3LBhb6BcJ7tTbJbBigCTdjZWhGpwIIVYid5HeU+VFqxXcv
nX4DwePII2X1lx1doMO/wAc27MArpeKP2FMWhCxKk3cmqcKJ0XPckqF3zd2WqFNWuFoZOHp00Jes
gcwW4ico+mJt07NqkCrVKmQPKvWXWv/AzvJHYuDn/Lpos2VPyd3AYTK+WJbKtXeBV4DSs6Pf61n3
p0wFcCGBUXiLLOFHUrYvkA0TBDlpKChNY0faHc4bujnB/G6fzKEXY6lvBUhoKkJQhcKbWHU4Tfvl
QS2WEljfGnSBqgOdRoba+CWxJCaMdg8on12bxG2GtJxz5LIZpOLPXzrb6MDh+DPeie4jsQydZg05
lLrzv9qrXLXlpQes6lTxZbSFndROnBDYa/Xl5Lece8tX1SJa9LEI6FScoMByHkLARFiyZ+VW1i3h
zvHqkUjdcPPleBNyAPbOF0HEqc3z1CYZhpqA1SbKaQSYqPystqjyiEFBBGw6HT5yMo4CFQrKiKlM
nXUaXg/qIzm1499Ue+zcowyk+ggPkgt8xdm3VNVSJfeQNDbDTyaYgEMPZxH5g6i3isaDsicEqRhs
S0O3n/pe0FAkjOogJI6yIQ+CWSYb81eLOXsTPLk6y2tcO0JZ73rAOFsFeaQ7jfFBHfdoYIQGrgNW
GACTWr/yaDKYrGgR8XNggfjtZse1EwRFiAcXofIjMS/kEdQj/2mLAFVK1dtKWAT+xHoI0P2sKbtk
mk7KQBBI/eiyxNQKpuJg0L1lvsf2nG5sIxUIU8s79mM9E3xKe17FlInQMe8yVP0Jnp+8Bj8f5qlx
Nbi9/Polf8O1mApU1CNiBVF7FpOj4Lvl4RJqh2ghI6VPvW4etPIAPaciPU5TeGk4//Mbin8CsHe8
lFIJIpYf69Gd3RpbkmlFuJJAZxda5sOBvnPpPh0txCLJ9cPL2Z870pmaP5JVLtPbtRLTT5VwjwUd
5TXa5z4BtO2lrr8YSAGIdgiEHxEr7zUTrwkuZIt+V+dTamua+SjH0acFJPQRXkYVRF4dSjkXSvco
bT/OWpfAkB3Qg22yZYccbrXc16ZBvf893WQKPwMPtfn+QUNYUdNO9Ps8VnCNLpQusIHAgwkaUR4N
PsWBZgLbNWDCML5N519tNq0p1o23hHkzNLzerbxExnN1+YZw/Q3OTRLX/0S+l35TnZxAvwkwt5eW
VYagvh3h9/z4IHjunBW+OYGpKjkbM1s9q9DKs72kD36i9Xif55DYw5vKj8bXlAYX8umNXoKoGm77
KSvi4FxK14kG30084fp3x/g8SC5tlshjL6/cKLYYtTapiWxyxP8+0fXd3y6hnN1ESXGZKYxyQJ/N
FJlZIn7vy7w1VSlPJ01JgoSV4K8XphpPRL+aEZHXZgmZv5RpK20Z6Otz+c3yD+3PkcLL2iW4c0hf
0rt+ryM4AzGndq0BDFbQquJD7dssBDOt1YDAQpt3RRS+Ek2Hvdfn2Uve4GMKmcTnXUZHgOkX8AR3
97WEPbimCCfgeVtMmYsN3m5GXHiP25UJRQzlZy2/AkncuNG/0cdWJAxjUuy74PxHpYcs1LMoPT9P
sG2UhyeU5OWkN7GY6LVKy6b8A0agFDCuOpEKNvRVddKJOLqwQ7fAH9T+wyILSd9jiN5FpC/OO1Sf
kPatr4YDpLxRjw6hHEZrwiyYUfdyFy6WN+9BEJaKIiRfZKn9fdfIIb020BCLV6HWhFRuWbo+FCUs
Qey6y4NN32m6Bum2TgwnUWDyxCFAHxV/Y35ZD0m8rmtSsUOb6ZhRibDHLftTZKRCcqB+zKrvfZmw
5rVTiTcV/md0fiEDZtN/aVHwoIvL9Gx7aJbSnuT4DdXDkuY7+PyarRl3oPVzm9kMy2IAAlHM5U98
0gSrfN959SuWcWsPW4U1nTWbejpPqt1yWqJUGmPAL5/KZe13tSZDyTjns6FHgw3OaEDIFtbvNxRn
/mR3nK6YAOIZ7efb6pqCpI43DhNFG2IzwzSME5kysFV+mMz8prsSxo29pATMqseMqYDbCM6HwaNi
oOMtm86SV1T9awGbp/W4qUhZ8smA59UwtAdAUkvBBDPevX/2fiAHunhjVrY+gI/ucifctMVlH1Qb
4cWGdGR87xb2C4qhju7mAzZyS3zAyGUHY+J4NBz5Jakcc+rZVXhNs9aSwavjNnEuuXp5aGItOCY/
cMOv1wjSHu1puvKZ6hACALgETs1d3HuXFXpKlhE7s465GgiV6gK8cd4P7vRJk4cR0Nb6+KvQl9Nr
pvyNwXNUsUMOM/QUzx7ugz0jr1OeRgJ3Hjsy+M0s6O9QNqt9B9qLA6q7YERXoP0qWS2KaOvnSTjk
xsjtrnaiZ5ODglMA5r+ZpGgf+Uxv/nTnUU+PAx2xfKdhtOCb3ZD3k1ZlYvu49aXXNgDRcuCOV9Be
kFKZMJz6vBKpDj4aXxZYS0W+Kmiz9Y6U/f2VypCyy4qvmlIDiHNCmHMuqHS4d2jG+hzKBBJgMNK3
2TKhzCodoldINlSL2vX3k6/6QOikfC5tt3KuBhDXbJFhFGpYDtcV8JkUXBfkQ2C7fy5/zixDi9M9
mCpg9wfkEXAFpYqAzsk9RTZneE+RgcCZRRvalk3nWZxmesGgzPg9vnoAmBAn5pAU6blmvDr1vRf7
EqyHjrysVvZtAh6dLobG0daZjaRcUlYYxSZFmMZ3+EhpL+JnrqOCC65qV9c1EL+fEHyR6jfO7htr
cuzGsxe5a2sEVeSciIYdlF1cIvBxHrluxHHQ07NfnYp7liCNsNM0s10voriqh+fqCdjS6QtNydKv
PZs/r+f5kAKOXVf21CcwLhzenBPcVZhvJKzNfaFd+dDS/dZtJFyWKjsPf948YFgb9C7Q4fLkud+t
ccj3C2w8bQshhAnQpvikQ6DNHZyZizX2lPfbiQlWbghPNwcXIXDsX3xZvxLJXXqPp1dp6m6U7JM+
Dfr2cejwSNmW5FiJ8oqYfW4NRUS+vED07DwNxFZgCJyind7SOJ5zhnwGvyzfiV1IZCD3aGq1dlzn
+qqRQuqgN+PYTHDrazoKtATlEnQrCILcRviAdcsIulTrgaP6rsKuVbixErXon52L0eKel1IqIu8+
hlRyvMpISL5tfud02gdLIlwONpVhonvzi7xQ6L2+HE+i5T++a72xdjR05mf7gnype0ry9qWeJsWn
QM+JyeYusuhMlQhzz0NpHfHfg+lNN+D+ssyqtipw71M6LsQlGhGq2WularA5kEAGKWaopluEthIS
C8zRz75B53F6fZWHAH/BYDrCp7pdS6sMsRNkVgxVbChkMU+pUEEfUTI9N5xf0aovu46DdESlBTVU
jWMQ2uWshBEZWrs2VtL4aawCMcA/mg/+TJ5wm0BgKlvUzuD3p1ESjDhKjZRzQxA5AIevwStBJ2eX
C2ip7BKzjyKgSsWnylEjgaHwqRWTIUpcZskDNFgLe3MIKGLOuz5EdK3d9E9/n2KATrNAo73yg3xZ
yuJR5LeJ+4tuB7orbl/aLn/L3+ZVY1xcT41C/5X98e+ox8Ntt/xOgWdZpJE7CyxVN3Cf6Y9Dh0Nn
mAu3LntpalUdvNPfHKFmQfkiJCTUUi9P01FCdgMihRj/IV/4VKVDGdPqNtRIg0ZhnKyZSS8cexuY
4uOib/OgPFmgJGPc788uUolbTpOXqZrUh2jBP6t6Jr8vlHL13CjKS2WvKHrDpFfJY2YXc+bqXgB1
zNqssLut/6YcBA6K23c0J8Jy0zmb+4400a6yfs7NA6+y+XX3MRaupO02WeVyvEEMhjYZ8J4tQFmt
7CImBGumjW22iYkBFMSboOvu8zbGUJxfaQmYZ4Ct7YYtwMbCDHOkGl0eh+xwtr1L456G+RhXsqcv
J7Vdlcm+tu5kEtpDtE9PvmBbB217gIIHt3COdYYFiocSYmOuMgSuaBnzqKe+21Ye/AFSwN6AWRSR
+vifWP3W0gRRZENwCml/X154dKiDaIPCdwEz4FQgp8Lf/FF3nyplnSEdQVJk8r+6s8j2D/0gPK1C
d2KoWD58Er7FXe57QtHhPN+x5IsRkMJLtIUJj5uCKE6qEXCI2pXqCPIWut+a44PTZ6XjDWBc5BYP
jz4lGKBRK7/UWuC9mtDvQgPipIPiRZ4Atmp9WhbtsnMOoTUfW9XLigBEcOMo/vHcO95fAEEF3hx4
GOFriqWngGTMgvNZnl6ARJHoJXz0g75dE5mqURtiLVcvCAUDfDa/GegkKeCPtKF/Lq070GJTQbhU
TdAUQZ8yAI03Mt8LJGJmdvwlcKc6mbnt+q0P1JHY2N938yLGbiTugH9FWx02RFasVJ08YLovGdeX
gw9NXkohsc6F43pQ6XvT2+lPW00NwUvFOR64IkzSuCc45RGu6ODGPWRvhiK0teRhBC5EQTXmthc9
U1h2BedVi6Ru85D1qpckrXl6wkQq4y4fnMvK+KRjFV4r02CR6U9wtDKI/AQbJ+zyW5cBw7DhxTIk
yMuT3TD1+HckvpFBk3ZQsQ7jLA4CBDJbWF0d9ZCcYCT9gpHZmgg1Adk4S54zekgO5YUXbI40b6ec
DbA3/LF9FK8izY4zIAYarQS1RH2ueRah4QZcqQ81HBfdvk4CX1ao0lpd6Q1Z4lhbCfdHdxAeP8sv
Xn0AZx3TGVey/b3aZvLzAaJbR32fN+4wJl0EqZV5YqQTZulR3fuLa+hQixwluVW338h6nWqsQXfp
/tOgyyeL9VvRJpI+M4tat0m5PNDDV2T1lo63/SiRxqiBHnM0mHRDfin1aHJPhl8A5HkwEpBA1xG8
sasLvddzT3K0Z+rBW47NYq4fgonj65E6WnCW8VI45H0iv1vGpVAyH3ItpHST4uPJL6/5WOg0q/vk
F19f14ng6Z/NXgNjgz/DwmtEjF+KAIvbcQoEVo4je4dHF4p9XG1GFhhMR5PZF8ymsziHpClGFSGH
/grvqn3qJQQzidjLzDJQSexBdGTPyaeHIjQ78S+JGwiqLqUQ1RtJlbiEGHpTek5gEoOb7K5knmcl
1c9MBYJoa/vCZ2IF2OOTCqdAXa/2su7lKmALYi5GoXaRfirPfrAXFTJGZp5P76x9ewDZVcHgJHxh
DShDYAjetpFzFms0pvWATYcDy5QEFdR9fHP4Jcw9HXHQ/ZuT0MjXLW0/JxWlF7NlN26oMBgjD2NF
coqcRp4/bXGSOD8rZnZUn70BKgYTGNkfAOMkmDoen2eI120D4WlN2mvAi11NAEyPkDQd8zeuNDgx
t+k9kzhRNiZwXpXnLsFLTxvnrsB6MSsU2FIbSUbT8Zx12vYg1zavJKd+eaW5ca1wYzcVBLsnY42A
M35lRwBWzzD3OVHQw8IKHSO5F7GBV+dmQsbXjtJuVgNW1+nQM+rHnTdfJCcprbUWOZmbPIPTCxda
3Ulu4WZkvhTLZsjy8vSZJBKUz7Jy/SCLaZOzi/yba9o/pklWvt0MY2Wmys4CMshl+hYS9HIwuJuX
NuO948/Yg1pqIJyEzlLHwFBPQuJhoakGhxiBagylYIFfADb2fydTmvNFuW3jNFOo9Qk58h3cSJQP
4Aigy8TDHV3yJBhZ+pYFxUQhKdnWDjEkC69AOTMoSX95gE7Du3ZCp3fmsu4Nd7Jnp8zIO0GP7iq2
VxgGdzxUyDa2iP9yrTQV+zY9W94Tv0QtROma+Y7klCqNhAbboZFG+sKdZKMLJXp9DH0opViGSBPj
rGM+cfuWqXdlxpFzVfLuk1HxiXAz09hu4CrYTJJXH+cT7aCjitly/V5mGX7Lz+ZKmYHz3yUbxjMv
qDbHe+vOtv0TlCfo7/h0ihuKtYfg6VqK89XiLnpszR0rPGZRuJIrU8ToBWqLUhHHiFtkDS2DchS/
ljaGuNahq09/vwTSYOh2sgenL5vBt7uRAvcIRzC9FsBzu+RSnVloTyOZkTGzUQ1t7ke1AWL7P5CS
8JzkURPBbHNCiBdArzSFVPZc5IQPvihGoHIOIACUv45oCLqK3+z20QT6q5mtU5LSmkRV2FrOTFq1
bS+dk5tuFepENXabQY5Idm8gGg5PqUYwVXOai0xrD2W2IPDYUyezAyoRIyfrIEKBAmDkMirLnhMD
c2U4NveHYwMuvJgc3wEay6rGvI8lfau5CSyRrc8JWlb7ggkhm7qAyd1kDAxS6iJk1t60B5X8xhA3
HjRXHpW2eqph3Wc0gGgfz9zm2Z3QHf1jbxrMiKnZpqu+OMK2mYy1mEXUxXNLSwoerEmSBZivoBwg
E5XiNwDQvrd+s1RGsCctluz6geR97LrSBpXVhge6AYYvSP3DLGaVloJ8qwCepjeD04oFp9wVJQMr
IdgpSN4Awas38AC2X/9305I0zfZ45JSX935Qkq14i7a0CVt+E+587BEa4FMfjDSMct5qFeW1nF4S
nvlxup0mG7clE/YLKbTr53abtN+FNHxMTL3HAK9vlfhBoVYQAr5+FYQAeyfvPwfMlscGMqturD+i
Nd7gXu8PPwIa3f3ATlIXaNgj4M3kKmPvZAmv5CllXEOd2wd/W2IQkXtw7OolnpcUfNRsM+DyHV+P
TgWCSGVQSEp0rrUlW0DnPpdSTRGuo5Qsb/IBDeY9KOuckHR47lkPuh2j5AUgP4m2xJe3Oh6Wup9K
8kzzT/1rFPs+DHWveDfD5nwg3p2HI6efpJCU5v3zKTEDCdV8U2VdVYhs9FTjp8GywhbgtPfxR2lh
EphLrSlUZelrXvCuLSOHBtwJy10RX5NzeyYFvWBnrRWV8vZltVkbRvcSs22ZNH7Au9tLOX884qqp
sfgfK5NKDSmrSlkICZhsyvBcvATPIhbPBSKVNjcTT687GKwZFSVX2qkwJDnjVbaU2jb+6mPlJRKl
smDYoRf9/G6X8jCQhl8HZ1jugdz5jgQPiAaw1W9pLfuqmQv3sJOFL/qYRD2lmFcOFoXTbrgxS69k
QJvAdLPmUMDBbrPM5fG7Wrc8wL7jkbj8SnUkKtZOs7R0NP0qyY7DXvThDdCvEq0K2cmL+pK92q+L
cRX5cV0Itz0b9XepNWyzKn8uAOJBgam1p0WXQBHMcBSN6IaNgdLd/wH48mObsVvLGA1NSHIFw/6y
fpdGtn4VQXRr0Kv+YkTzprwxBm8OdvDSTBFGEG4/61RW8HbRvISMIjuKS0qDURiBHVf0EEHBtNbK
/Wvh3s3RenTggEmUhbIgZFzYL9nUg0BVXYymjP8XTUM3hYdt1H0K05A+QS4GzFycC4AQwTX22RLU
xufKJOpUob9jGcW7U1jw2j8e/05vTTnJ0nb4Xw4T7HBx3/97UrHfBmSFP9nBUcQVJs2284LPXlfK
H5SS5f1vVKoLKuGPNcpLEz6o9+GeIdhFwLjl0gj3GNayeXPoi3KDQfiuB1cd2q37NJKuzhu2XL5Q
0hy+J/KrB3sywNVShx3RVLzzIEq669bQTzGwz4CsEahp1nfTt4QZ23ivvPEku5ApPywjhHTBdcZe
wa8FKsPsU6NemMzRUWE9ozjRFJJYjgSozFnkNmIKBvAHRH4VL6UiaQaj7c8/xHxx++z0dXoY521O
hWSrElgr14+otbTBohqgfQYbHEe3Qcs5K56m0X39eygKvbBXT++k9ahNPzpBtDvb8zwLkeIyBZsL
fhUvmfCzjsGqIq9Oq6DVXhU2wu9qqazbfNwYSekjRN/Ncj3K1UVfdPEwgWwUPBplInuxvatRfdTE
Rt44DhLuJQuWsOWQ7Nel1NtK1Wcpm6xzrhF/tdU6zUFexOkBgMyqux2J/iUaWPSv7UfHLkC8fPI6
edBp5LcF/zRtR/dB9JY/W4l8t8BREtsRLlMK8tFJuS82qzXe79k45EGye91OBCch10Z2fC03eBcv
Yfnm3OsN9Ti+HIHQUCdnf8+HyN06qyQ5i0iVeU5wSlwgFrZd0w0MBEBeXtxCJJpN+jwNclhaZH8V
VXvlQqc5OI3LhNtK8mw1YF1yFYSA91GZczh6dCygcDV8EESj6OgoLAbLNk/xZfiFHo52DomaPial
jYjnr3edRjyLXQNb1QbfaDTypdyjdBGXm9a973gbn9vKCaiLyJKEy9XzBI7MF3yJiWndH74UEmtk
3OqaMjOGtb5iuihMRkKaHkwtVMD8xvFXvuppe+9ONud5QOgTSZDOnvzGdWCZuk4f1o2GETxiVWBk
th25lMLn2ruV2kJDLIa8RxQVxN8Z8e8Cic3SI6n4bpjXeeRCRZGLg6sopm5obMHs3xKwmUmN1tda
fHNxmALM+1VzfzOlH4BSLBvaoe/uVN6Qdev3g20KoHyZC5PXZdoANPN3FqvI7JL5TAwXdd3KHdcv
xB1i0V/Cw/V3LxCLSDuxeDKHiRp2q8NOHom09K2xUF7ItypJy+UM+F9sewItxqqWx5WDU9mWfslB
GERN/7rMuq+7OLdu+7iguyYWRdflIroZmhUbEb5BRAWNkRlJ4CkNN6Z7UDIfKwVugX04Y8uWXxsp
0Caf45UQebJgp45Xuw5T4ZU7Ec4IjKEz6cRWYCe+yQ0eVGvZsFJD2OEwtmyekCoL4xcEcsnCd1OI
3AwuW0ph8OuFfOuaekiUdtAAbzvPTcyCZzxA4a2kZoGhyB/P3tBDfaqCc8RXJytYLo1UoAVKc8oQ
9mdQrIGkKkONcn9SRFWm48TCd9blNMYUW1Qv3JnlOT2UJMeWgBtlv5XscYdzqE4fs35z8OzzpGyM
j8spbTtliwUP+f647YdFgz7uCTiAPkoqMtk8JxhezXrKP9zgUMTO62i0i10Go+u+Y0TUKqJZML7A
5YAJdIDnIeDWmgasaLHEF2OzZ4/SeR/86jH6NHoRv9JrfM6dwuT0LLSHYoy3nympOu2jE7pY0bSV
BYuFrOl1/R3e/IYDgZwB4iKlsy46va3PGmZXOrbHGR4YC3UDPzaMM2sg62pgHY7ZaeimaLtp1/AH
KSri1MXa96DEHLjNhNWBKNz/uwVgl4c18CpvixH7DxCGOcwkx9cNj3W0pZfftmCYpnprgoH8gkVu
Y2jmMY9uQ3Gyi6alGBoPwDOVN64FWMUtTJh/gRxnE6ZpaWMDyFe90SomT8m5PbFft27EKkYQlbBJ
2/qPYYygHPMRLO92FTmPDJJBOtEOSivOSVdBKsGVO/UKjXeoYdCTOrL+d9sKGzcyfKXx4s9DiKbo
oSjENUC8ucpzBqc6c0AVThcHrGy/2eNn14s5xqew8kA5ZWWzgNV2By06pxw8/UlGIKo3MFpzhyHa
82Qa4KmgS9PjMRJxIpwAca35lKV6RTrySCSOLqjPC5MbNHANp0w7b0xEUSeFpMd/T6/2b/ycllwE
nZLlT4bu/ih8beRtpQlydPbc0RTE4kD8KQWYAmHNyYpUOp3dojf6+mHeytkqwh2TV6NJrgFP5ig3
UiGR8wZC91l18seROnOYG2SKDA5uwSSXPSSWSxi28WOXM/AyHiECfj0zg5pRxsmBLL7vV5sCWPeZ
LeeGYPnHAWraKXASLBiCTv7E21tH4gUuGZw+lJ4CF7hNldiEQzypx510lctsa8lr5RI2ab3hkr4F
P95MtAAzToAJIcKVip9UjlqRqkPSpfytpaHqISMn3cQpg/BZ/Ta6H8hR8ExtKMgTrWw2y4gUfzli
mZaX+91C+x6ZxOIP37gZTx/RlmWAUzG+6ULPnBUEJ3WSKs7lQ35BPqChZe3rBuMWM9aRZHcM5X78
MzB52sfZde1uKzfM1tayhNSY4t2sxnAe1ZOQ+BGefIAvuJabLxNiEtI+vyuOMp4CImekrP00SpAx
X//BZcxmBfOcGN8HXBoPUOPeur/5A7NRKT4TLszHEwSEWjD3i73UN73gaDyl6M8XUJ8tzJvgobuK
sn6YxxnJQFJX26mR4uXrczsvco2A2qhY0v87S9e94EFkfRF0yd1TC6xLBnAsswrJmw1ICPXV2Bb0
1hgSEJMsRvYsArvfx6G+IAi5bYVAUYdrZ032pduI9VU2pxI+v5yJb8iF7BGp6SP619/c/6lGZoay
RorTrrc75dSnFSh5Zu+RUayjXm7pID4dE7h6j4zSHcgoz8/vqhr/lf6fV111oHHmO6MDl08J5DhJ
Nn6rd7LA0rwA1hpaUgb0OI54CE6Ci+AJEecBxGDBkzPS+e2JhnEkLz2m3YW66bL3v9FQCFDbjDcI
IPBUoAqiaY15Nbch3ykGA6mcIoy0ARB1WM7j0PSHMdPfnIYmVrK8QJzr07jfPJ8cl+vlCPZTVKci
OGC+3M+vl52ZvPoroaowyQzC+HBi9baXE/E18wLTf+Rvu4CwE2zpdC6j/y17z0wyG2ZcSrzPpvqK
jh1QPvsEM8a9rSR+1LsasgHMmOCAQ3OcFDKnmdbVUOtWQ/nRiSOj21+py/Ysw2LD2Wl6ZRBe65UU
BvZZMflBzN+YsZIiT3jGJ53RqIgY2q/SP0/uQZHoQWY/9LbJTuPQDeVxyzpIk6vzJc/06qxs8zgL
RIuP+6hRrxE6CjbsSK7nOr54cdm5p2KwJXAH0X4z+pU8nyvDIvVz6ok00SPGDF6bDP7KrM0mMAzQ
gfhWWM8pGdNQn5+oLBgZspcO30xEc9jvGW0YNF4Vtd0pbFKiQGcMjiq4t0go4G+XBYpxXFmPHRLK
dENU63ryWa5RodEtE7R9M1v5fQxq58GI27tnscEGTrdafxRKElUHoC5eCmLiA5sEqYKZzzDC5rVO
aLwUsA64zVx4/jpfm/++erRF5qCShUZs3+bm9d6mlvWYou0RVKxF/MJFU5W5U9Zoyp5XucT9qeDg
ek1PTfFF+9M0BVT63BQJsxJrdGRCB9Yrc567utz9fEIFEG+4d6KfzLvDwc9itE6GIYtcXMsODNp4
tpt+ZMxi4fWmkEhq/PU8cYCX8x5rIHx8d1ASShmtzFpm8+xMLwrNsKa2lcxh3CbAcbtXcRc0ls0q
1L1WcV23P3726lxn7c6mgu0cp42+I3W8IducruSGSbF2mCmVTDS0WNEVL4FckJG+CxLfSdVNHWpA
U5PM9LbuVsY5sOa6qeeTX6zVkmbs9YFt8LxxxWkyvvYR4pDCf6abxu3V6tRKaJxcOTeHHuKqqVVz
cv6ET2NL8kcPjKWwwRdnsu78tS/le99lrEeTmpItvLWEBKV2RQn60dGY36OnBheHOdnokc3WrFw1
ali0BZUoOqtaMnAkRS/7eJq4t9pV7yinoOQXyaDkcs8z7gxkAYXL9dpTUXQxjprwXlQ2yDTCn64u
zS1BL0t2Pm63KcHhwx/5zq9pjKAncqf54WZiIEN5uxRpeUZ4hpLLwp7bdAZIJzGfP1ensVrm/D/U
tHVflbkSN000RKeJwfrqFAZ33z6tR64BUvu0xRUlws0u4z7AINJ5ZL82M76Vo7Ke1JuR+w2s/TGU
z0LEzwOYuq+sWHU0XWWTqwqyDXNxuqp0sAANGci0RvIgTzP0QTqK1LYzpAAPSWupoGMi/pXXTJur
XX/i56NROdvdjbLXs7XlskwajeVHvMUVbklEDCbuEhfgK/CZzqAgPlC36X/uSvzFaYq31Eea02Q2
StbkEm4Vd7eEvblF+pCFgVcQDUMR+IRPbAGdAzS7gC2GSRip35LaKwCoZZxrTR/vXPrO6JipPL3c
43eY0nuKDp7lnwCy71+X+q8RDrvpZgzyO/iPRZf6mLt5MBnnwCnn2+kY1F7Nir/3PWb1lLLCAMo8
wpu1Ddc4mICfExiEW01OaanPRxk39LoB6iQGw855Gh9r4p/glM8LiseFtSeSUOmbVvd8LYF2rAio
RYf/9UU0RXvzZ7gbfU/NBnBETyhwMyT8QCYhZFC/sgUuPVVSKSNng9XydYLlb8RyoouYlyLz74NK
Ekkib7Ou0CMAoJ44Al+cFk2d/WCoyCBIHOLiUXJ3D7NHY6K2Kf7L8bZlHIdRBY4qxA9mfRWbqoae
s5Lt8pafWikhSPpJwUykUpstCVlrbinVSaavPokjMuAU0YtdDGEQ35puG5hNeDeFHBF5CEFUScja
0ak3dssOrK7DnK0vgUmrMJ+UQpaY71tSnLi8y9j31P6v4MNnVsPSmklENh6snaSIu/hi06T3KoBi
EKgyoW/DStp//qTyaNLEl86t6XooLmJNEfVJB7eCgjFt/Iem5XDlLvlHspYCN+OYBtaetTK5eyvA
2UT+qmqxVXKJoXEWs74CZ2d3ndfZdjbCCZB7UaKjBpfiV1mmfVUkbzC5v/yl5dxy1XsqeAc8mxuQ
J7MeaYFGM2e6SpJSGGRq7NNLz9+Ky1fbrNm6PiXIBwXTQvmnmBqVnzJcsE+6zGILRbjVrkVNIWv+
qm8sGJPZZFq6NOqHw0stToUl7qFWQus/fEtHnwFgagjp5iHYLI9d2JsXWr7Nx5FAeTDkMdvOQq6E
oiq1i1qcfYUS+zTOj3Onph+UIWUPJkSeYgSEpB3hYlqz3bOZbrrQXPu48ZwITEOyPNkcLTU5CSII
HZrj/CNJMwj5twtABjA/pDMkESVvf0nZnFTXBGijM8Qmn1ZPiNro85gmcDIy57hgQobOjmHxHcEX
e9GWV9JZ+YtmQBJTdGISAIrtwGjnyWHS2cVvg4VbG1zFyLwvb96mBTiUqMXWwzWfw6+IngpFSPgX
aRUF3jKohXlQ1i/tvK2JpATr1S7PRWJBAgG75kDZ7D9BTrlESwB4oxPQYUWgkao7d2Z7ZAd4neeL
h6lLv3bol+RuvstkdjpFINAfo+JASQOYAV84DM4euIHv1nszws8xgkEmm4qx2gTHcMRRZ6vM/AXP
HE8Yp3tTEFIdALBPLN9ccgKB6JzgkGEpkdti29+HOwSzr3msTMaYXxO27FteHqNvSdJvEXltALqT
cywqnXRioQNM4NhWegujEkv+5uPXYpr8G3lFB+FlxBuz/l0Yrc5KrWQ38nWdoZnrr3V/3exOFLnt
BexS9XVdopyHM6aavGtxpwgfoIyIhlQjWkjInN6v83c1kiMvtyCHoq6KipGUjVXRh7Ds2iv0xGS5
C/C/2KwyqCM0a2O2aYfxYCPQnt9OaLae4e7cuzWrB+KRXr8YZpUBz2/arTpc0mwhgozcMCcJ33im
61joNFz6RSStQCuPAVNtcfAy7NuTG8nO3xiZGjRfIdQct9a13xlb0+6JmsY6arnnDKZo5jrwZYTH
2Z72EhYni6HBwnN5hT5GsYoJIgpSsdH1XBK1MPRhIkGjR2nxgZsJ45+6k/ordZ1yV0SENxpP/F0r
XIEjCNlPlHFC4TPfNDMDis98xFBL/k8ne5WlrPpfL24VkZRAA50wVMv3bAPmghtW5imtQ/KiLJW3
P59OL5otQS7wB+Vs8rlFxXPkEszdiA3ya3Ur3uj1kihQOzqWljBq0kXqkaUwg6IuY4U/Q1L4XY+b
UZc2B781IyCcezykbpgFv386swmZSBYa+qoaUGA3MdLcLn3z5Cd3W2B3o+Hlcr+EAi7SOh/9ae1M
Pmrouw0lApF+J6IkyBnjYQRN+Cpt5GuedJEzCv2e2gGEGuYmOlMrTaL+WlpOJzytDnEdgpE+2ple
XzlnYhZ9KRzi7q4amVFkg9s3EsuBBhgqeYGrO2Rj9MI86QYXbba0JhRGIJKYHNL31y+qIWyfycq3
O1PwCi1zREBwZ3Q1WzLvIWpZovrIasmRxM1ZfRyYI99tXv9qPcjQt8O89yprE8ia8T8GvYaxdy/N
C9P5l/NO0bVwPz14kzJzcy/EZ77+qAwxab2HV5KgDUkEEELvWs9Yh2PHsmqSbwFYZyu9CJV24HuK
kWaNlu59J3PrdfSUaAmPSEVWgEr4ot3HTV1BYCkC2SsX/v1b7wLEkNvq+BTg7H+rA5wQyBf7fdxn
fu8OTX/BhnTclL5sECt9vL/MCNQT2B9KgFCQXGxbdGTH5eCggcNM0VIGRsRedxeUeTjCOwyerL4N
Ay+PeIbFjQ48IOAcD2j12gGSv9ytAzbTc7mr5BplxlE5+grK+QRM522vLdDINDB0hswCms0F0X5n
lOi/QCv6fvftW2I1kn6DHKwr/iHczMY8bByfMS6cfbzGmiv/JayvDPvDNlDNvQvBC/8TbdDk7osv
uqqNlcXdc50RtofHQ/1FIC12OSMztcuPfEv7FVoWxcXkj66ni79h+D/Va4es+7mQOAQCFKvG8JIK
k0BjlNBcp3ShZeMhZ6Gol7S5ek4njiOmKbBcgVm0OSrQyEPhrackrp1L6j8ZP1pH4NdoCRYbMNs/
HWYsHb0ZN0UPw217lc1SM3SjisTgU9csGEy5j0yeLXWBZnnH6MBf68RTGwXWXQD99nbCqRbo3ylo
I7xT50AgOV5XDtylDncNqFx/aRQe2+znpILOpcK8re1ZFX9To6yc/8j9tYGKJeljpVNu4o6JrNT5
17gmnq3kZBt/Q4f9+SleWvVm0yMXIH3h1N5VShqlUtbBKiRDilUBDnyo4kqtqimu9zsPhjicMsiQ
lVfBCDV+O8evsvdJ8VnAQtMNB9Bx64zCkEEiSGan2mTswaU0k+3Nmj/cwRinwqiLB9BoGhMZVoYt
PYpTyXprvFNnqwtLY2IpFIYe0Zr3RtFZn6yXWdi2s3ebMwlX5QFpVWRX1kQV2mGwgjvGxfMTnFMd
oAdA8BR/CaPM+qQR3pFYyW1sfjqTUEd8WeZZQRsgtn9xkNU77V0oisaXk+xRX/T9Ko99LXrx6yLe
q9V33dzLca+rEZWe/6tDsI2QoxMpZkgigoj0yiShSnwzSJ9vyVPVGBpJYo+GbEpKmyVK8aCx3ss4
N8qMuW+quWUAPW0rw8MOhfPW0RFQCCcb5gszq88HWMrvOhpv682ssyZErVPoXwPPOrjkdKUN0CJX
bPoq/5DSNoHG56n6jMtO+k5aSLpRkdOnGrpizXRAmGF20le5lTtYGQiUHWudBo1m7G/iTnKxONGP
2oZDBh8k2eE3kOGXiOFt9WaJOM7Ya3UZ54K8FOOd+gW52zz4qXNksiyDoOtmFO5jzPKQ5sZ3eFtv
jzUHmms0VIz0WfnxeI1hyVP2D3jp3uigzaJvObdkLZXSefw4Jy0RSbIZ01wJGriTdl3+bMsn4xKM
h2GaH+AnX0qGpROwXE5byVq5xNPljxKv5XswH1FIOeL4+K4AjuQpAKCtVnI4s9ds/+glJ+dEdwTv
d0zMqsFKlkhmdS3ojafbPFTaWjUbd5JqnRiIsRzgwYcdu1TZw3Qyg8BeyQjmOAVUy44UV0Q0Z1Ju
MXn5ncnQpC12kcJbDjLOQRCKzWiLn1WCpQWKgQAZSknKxGlQspUKFwH7vZobR9BkpH6kuEz5bpHB
i6Fo9d9vzYHuK/xSWQRuxvMRdiIFLWOWcsLP6ARS4fqjC4Y9uUaGNhA1MNT9AZdWM/+cCOGMFoIj
grVxnNkI0p70rHUInfOWLfUUiukgG6RBMdywCmqn26SdeABZ0alJPxok3SZ5nZI8i3wbJ9cE4loV
GHtRAVO47MDIBnczXVXZ3sehbob3qUrNXzfadAIGjZrjwgBmHE5k6FDbyjIn0ZTxdab40tJ6OdV1
UalHTZyxSt2rYAX0UX8Xqvq94zEgAvV3r5YcNRvX6AFshIfA0w9jlbhcBSSCc06OLO6uILiztXrz
MFbhWEYS7Rst8wCI8Mg9b2dYykD8rxhzHSeXFt760ji9HYC6ARfxaE/ROax/gxYnxS4G7ioiq7nT
ydmypR2Rd2htVL4IB0AoM13t2QRpBFSyFw8w3hfA/6Pst89fWKYfE15GDBe7jkhRj3FrenszEEI/
VjLr+33Ak0Eba4FNDMCco7wyPABOvwpftWvOHI9RPQ2RtrKawct0iP27C0aWCVvS9PaTD2UdvmdX
Zy1eeUhX3TSecqHw6mL4uykD4+YPlTcBnWkSFCQH7RlUUUQZ+3TqVHv/O+UZmTIvpf2QmLsjS5Rz
2KJR7QhwSZpopzQbq8WWLCX5OX4XF9oA0edSJEk0GjUN1Qgs1By8R40lEE+//45x/oL051ffK3ZL
h9evPQb0yjPk+teDclncC/FYHnUKWFQyiGM4ga6a6JblxfNpzHtesOwVp8T6tFBy8icYX3K7bY05
S8sFHIS8m9+t3cG86MO/72oDqnx2DxBDETxi0KWYEKGNZ7vivl8QvDQKcomydZePpqbawJc8oZXy
0XjupHzClmL2QhaNNdgYpQZaui12s1SB0c607JHndzZSfW7BuH3RMczq5Os/IX9RpdOZ9Xnfl/Ev
Yrn75W3mOFspKAWlX0+azmR9kB0w+rDmW5VHYOOm3dnEYKwymKisk4gXwb8lHN8jHL8cXg4CO35A
G96XdRg5g4p2XHrZ9LmIAdjIzR6IS1EES+5WUP+xWLDPTDIP9bRYnPqf4byK0r6rZdaaDpcxCIlN
eUd7kKPt/Z4g6b74V8K9zx7TLhkrzege1iII+nTOoOkruUPbLF2rWqhoB+i/mjNz1VWLo7XCXLCo
i+GJWelgWeR86vYU5B/l0I9k7vSVr+FsWSnxLQ66gtJMBS4BOJhWO8s8/eGL22i9QusARY1nY5sh
ngxL2+fQY+TiZOPaWKh8BoFDDn6Pvlb4v2GFkEWbRCKf4gltAFGfu8Pp7/kK/TQ3sOt8vl0VexF3
olZ8xrQl9MrDsMyL/b77qx7kH6JR/USK4JLb4n0vvH6nTgEiAkeX9WX6VGJaCgIKcb4/5lr3tayH
ZpPnY+A4uQGWf2NMsRAqVZQVZtvW9U8DqrJ7ayqDHo+BJ2QpIuQQ7ORvGDHXu7/19VzrpqHzoiLp
yuN6j6bKdLCBfOfAELVpwddyHZgyED6+h50A2iiE0KX/Rp9qIHQjo/j9wBDwH69ITtRTgVzrrtpV
YAKDO2iWDuwbsIxvdFG0FUUOet0BCqRS9Nrcr5BfUl9D/NJls6PVALJlu8ijmaWsxacfYeEGo7HG
gSLWt1c9Ap2lLxSvPVHBNzJ77X1s1J4SXBZkRirXauN1tXhbMlcaWjFoesDvBQtcVlNHA9pRvf2+
7qKVeatlHBJKjYTLXq14lVZuYyW+wurt7B606v4AmUA3QVbcCLw1vi1Xgpj9BecpWgUoD/R4mSRV
ZWv+StkumqI1gWb5DS98gzSncLCBY5RcDhDdiy5ds9vB03/zzLzMD78dN3lY7pcV0Lel5yCLyMEj
UH32zkA/0EpsJmi7q6nkQdtzkyZVC+z/hgb49pvHqt1UdFfC5aPBMH0uzFaS/oZxgAmd6xj290uT
WMxV4cyi29d3YAP9WmbnJg+l+VyK0qKhfLptl+QGOzGOp06wBRED0jXf/oGfpq+IRbiCnI19Wsn8
keC1YsBspBymKbVOJyrOc0W0/3ZvxlOrsDuBVihjCGWsshC/pu7AvBOw/esmgplWBr1UynrHwlzJ
FRBeUNmMGYKsgAnLMWW9XN1io1tJxBDpTuL0p54CsnCYlK4SQSxlNC6sRmMPBzgAo6eR+7Jns5Nx
SZPveVTME4aLYanHUrchjT/ixZUML+K0+Yg/xcGn4KlsRelUMSQ0SOfcFlcnYB9BF3b+BJFL9TdP
GqlGF/T7LbvtfDh//kPcoMIoJT8mbXR3MIzAL3uPsH8A2HHPsItQefYu/dQqoI8jwAG+H8BI8nN3
DhXihT0u/L5yl6xH0rfwQIitMD/POOuyTbTEf2mud2k83hV6s567LSz9w9yGe5xvM7c3fZslL/BI
+nTD813clpdSiN+CntnH/TNeZM87PITSr3BlO2DZ7jXoXrQKgcoxJUouExhtJyFFAtYDM1cI0GPl
ZdoUvmOdseGJJ4j8aAOmBU6N+IQ55U2TLLqUHSt/34m54VGfRcYzBF7C73U8bLrVCk/0JlFqdgbc
9462ippeWLVhSPKesfae9JZhPxTVZjDhiOFCUaHYrTX9uFADjEM6L23vRuwbTcfYfflZa3ToSsUu
ooZuP3+xrJUbNkj218nX79X9jLJmwoQIcjGBfgWZnofixyTTFmVO7s23bgiPE6TIktQr/OPtuHG+
vRIDZE/gZ7yYdNIHoCy08BljqfGsUIg4BZRvFPxutI/gjixCNYDhMkTVZSIawmjIu29jyushzogu
cXGh2v3l/7JWB0le2kEXSpyTM0YQglU/CzAqoMUGO2Jwq2D2AjJTp1UftWDX+CMxryws1dlLu5+V
TzvsK1gEvDqFOU0g4NzK5xkLyH5KXqZoj/IcZwz/tEWh/UpTdj2lEgwW9zDORIjUNuf9NIjGwDfG
rpcZnDs88FCKX4U/uiXoPEK/e2i3DVWQWYEVmXG34RD7ZY4b1hHCi08wp46VDH+Ig9+k83ZfKCj2
J4MDVI3uwS0IJUk4DuXGJONoAKef0V2Mp6DFIqJMnIxONeoiaTvBrfvhf3iipjfM8j6JP6Joj7+9
UhGl9tTgZkj6dDb6maEK6U+Q7+sew3n7Nj67bEw1pYDLgSLohbW317lcPuYo65GI0jtwSP1S2QQc
0CuqAtcUV5TYsCmvCvsKdbB/SW9hQsEr30lC4GAuvgyvo6duik8dZNoUqeef/VLp8HNQPbTQx6HZ
996wPBNYBUIKSAMMPH4YnqIBi6wJoQWoD80A/GKk7MVhnjipYllQwCheCxFa/eLUIz+7MrAwjwKk
f65fVBGtd47tOLV2pxUh0twEfInTJoDb7tKR6war4kCmKoJ9OdwyTcfEBdOr9j9LVqLYPwi9i53E
rWSYpUuJMfuWNrN9UOFqKTTbpsCyu5y/3Qs0E6xvm9c3DOArT1BmSpkp76xEI4XcfJGLgoCZSnRD
6Yaxg73Et0093Wp3M28O60paRJjRmdX3AyPMEYG50VxspEMnojXdnG+djasxANl+26zrmF4oabPR
rvjcBjkLRVp2dus9Bx6FdIuvOMFF5HUuyhcvTB6jvHOM5i4+P1k/MndGhWLMerUu4STz1NkfeBFB
a8+DUDfk592pvraswnM0vbav58knh/YZA7uKUBq3ijmiOn2IgZImjkbTRG9sUjP8Y20r9QmXTHf2
RfQ1jMNReWE5NUqgXLLCnzaZi1p/vTMrRkktY2bSa2C5FxcxojMggjP+6ci/z26fLJBIdyeW3DiY
lxFmvHD2UEyOblbEehV6io8RPFxB4FgoquuRt+PMD8T6r+ZaczrC7N1s16MQCpbvPfLq6DY0Z3qL
yse1GdfzLZXU1tRZkhU5lpOHtc6HlTbDUv94yIqX4Vj8Mv+Ci3cw7PvNBxAqBeOLq4oFYNeKtEka
yLK9SNh3R0RIfvFk7XGjZ9rB8v6k4B2olQZAh6ViSoopvB09M6XsSW0UwLdeh08uxBCV6iS0YHL7
Ni2YBRweVhv7Ds9pNofgKD2pp9mFKkGlVOji3d1SDkGv9gXifvcewKBcOGe3tqaIUZmZ4kQ3fwJG
WHTtbNLpJ/AVMWuqk3TucBmpfrDzZMiQALFMFosCtxxJMqT1/7URn733kCD7/qjuN6OOsVkeb5q9
BDAtGjaMGha63KCHu1c4lCu7VD2HFUc4s9MJJQSMX5Ow+tnXvgG5vYXTG8MR/UylrWWpy/PxwxZE
ZVJwkhpnlASYMiwqh1s7KV4Mz6E7h1SBpS+jQc8Jda2f3SFLIeDPdB/QR5wnEi+5vzEAEMwmcSj7
oc5PSKPSMVlryenhYUvX8KPxRbVsx+VhmYyr5Cv+alDida6i3jgIPEfRzDIN60cLcbiwAtUQATLm
0Pz9ujyfX8rGbvGlsCd1RhWwB/9uC/98Fh2kDZT9NNPrnd07ibjWTuvZyWTPSr41DlO6ugweNeRM
0sb7q+K7/Czoo7dmKVxU7zDlHHDtdebi7R2iK5RWVTuw0Prb+BHR8hZ8bCOjoKzl+LsLQnYdHW5A
0LJUULisj7pxEiY64h22S05LvFi1aVLLzxTjPnGUeOCp/quUfTp3aBEheeBCwqQrvp+KM92hlgJ8
A2nU2LTw6eyaZ65aMB1++5SRx16f7eB0vo/c3/R1aumavw6TeAnbtKBVIxikd0bUsQk0bwVWwrap
hhvCEhKeWgr0qimi+vQ4KWENopy/3DC3FwklJDwumfJpzeSgaCJcoTp+hJNFJhTVNLmPb8VREBKY
a6qsDZ4TMHY7Rn+OcB0Ja91ByIDFKtP6ZRb3bzzlXJzWc/4XFuzD8UTrdiI+WGaELwFt6cbhU1/L
LJqrwPhHxCEGJI8EJoPMBnwUYIg1W4wxfo+Qw22fWucYWNOgvnpDBxMhvcnHzlH383rBtImGW6pZ
elsas6WW8XND7bN52oiv7nO9DeEumg10MhhyOd5xncv3qkb+jMh+FjzqHQWH4mBCXVIb3MRZjgWJ
K+DTnvIV/nCi7Fg3zSr+VspobVvke5gpSewdcBaLP2AU/nI3lPbvvX45fhfsfCgCjUz8ZHLitEC6
6ct0xz9tJQdQ2t6roT6i/hKgZwojqk4OFbRL45W98j9eY36bULA7ch9YG0vCs50qspnNtVQVvSVb
MpRDy5cJq6eWGrdSMxzezfbA5He8fU48H2HUbqbr18MxKTILlZ7jQjmQv4Q1/ef8HjTGQHfmQ/0a
EyRjgNcNLdcQA7gJYnc3+1MRxKsSCkzWcu7AUK0065+TTPjVJNit11lcqz5jhOO8EZAlT79AmRdq
Ov8Yf7BZKWkfP0wyT9U9r2oZNPnhJYsHmV4oG7h1drnrqOmgcxIuAgaI1kpWzZECETPzoGgfH+wS
NAOVM1cEIc1tHgDMvomglDrLoG9kG4MNlqEhyp/rj2ox3lVtm40tQAiuCM+DXgrJVQBUA6xYlzzY
OQyjYSXjUZO9Gy6NMDy7jR5m1aKq5k6wBMEUHqL8uChCmRvezYuTbj8nPhjc2DeKoQbyPLZTWfxa
bozwpes/esAuvpATjCtHp2PHpMfv3v3nFd8dW9YGNDFCM/6+VYQSGE3okdYZnpia4KZxELlPYV1i
/5hxo6+2oyCZB3kcKgVWBxUCEAHoYcI5nl9U6CjfvYsTbC2Hoa6i5eKzs3yLVbrnNTconEzGw0RP
CBXL9MUKv8Y/qGwC6P4WTxg5tLRrZfvtiAvl8eaGMxydRPeLR8ud5eRPm1rKd8Bv4EA+ZeH338FY
QWEf1td1wlvUZPtKOcssyrEvw6410udB8LqtMMYjQ434wRE8++3QO4OIUpjZnBsGZ6UDOBlHmjC/
f6u9/DD+VCARL+hdRIEjf/YyGeJaC1BbGwpjb4jGFzF68d5/bP3W5QbZttjoekpXI1K6xwV0STPd
tMWxmnIeDLoa2XQzffdkLGoHU8WyY5NvBLdziL+MyL6GhMVCrj+pL1rx3vOIFFaE29SYpm9jXyy2
17dnHDmbUfP3RovA9MlPk0/WmchKIZahFm0gq260EGM83GO306J6LLpJCj+/8lSlnBHt5z+yDJ+A
HqosugHuMCB50jbHn6mFfm+w1yPn/M2MB9WLk5e0UhPDqDvosZVUaDRLLWl0r3Sotp544p0EnydT
NcB+UOrjLBQ1M5NNQrZh4scEjnXtEVl4v58RlXauVB7BOIP9EV8fPsppqoVIJwtcZ5QTK8TI5hhh
A9GXS+gjDy4PUpGEqh+ucCVgefyPUEbdHWVj5vkr1QA/n4KqJLwRbXnKuyympt2wY11WMvecqHca
twSlxvYrPTnQty2ZJaDJxsTZ/u39hTrv9RcvNmXZfyV/jN8Th3Mx6RDECZhGyPlHoT3RrGF261UY
2oUcgO44nCHw4neWKuRo87loWghWySOiI7w+7HNZR8AAJGMoUJOWbvVxJ/1sLQNsJXU5tgiDbGol
yI2hvCtrtVSaJWHgAzkaVLL6jJ/LMJP9S0Z4cBVI3guGcJrvmzfPTvQwp6ic6rBaBupqrn7mma8w
TJvUHcagGe5rbZKRg6Lwe377nVbe3rZzPEre1JcxTsXIowi8Jlv+669nfwx2Uig2zqLY4402bFlG
wPJ1qqoaRz7hMjPxBKsw7lO9VL5OoqejB2uivn4UiixHjhneKpix94hlbnmuMeVKo2mOo0QMDJvH
dXdOtaOW9SMUjSqm9D897UMxcPnWeCJn6XEPkxU/BwEHW6/0glx6RrSRIhKCjl0h2+V6y14nKMz+
WC4dDCXdMsz6OGLfIqygQju0WTVP5KV9Pra7mfRQEf24NBvPMjSG1wNQsiqdas1NhAMfAIspyx1F
P+b5EPhchi7rJ2Y52OgMazr+dmLwfidP48t9CbrSLy/kd3vwIS0LMxxX04N0kAyZcsHO437RDo59
op58QYK+uXjiW2FiqWBlgu+NCJPDFnrPDgsZBNsVUK0fN/EWIiB2SZIDSSRil/qZNRamWBjVD6eb
cJJ3EYo5DOiAGv4xRXOt9XvaN3kNVlakjqEfIoofV+ULZbnbrd4DL+DaZy2nKJ+9ml4Weh/Ff288
xcgX03CuvD844hakBt3gHEBFixIpF7kTJIdUE2ElTpaKOAdf9GustDoIPGqLXEPcZHYAkcH4jFYT
NKtbIc2b7d/dJjz6oAfFkL0XE9DlibzL2zPUGCJfuAsFmRx1jmFTZc0dFUVlVlGNBogqAbZdOBTC
K8sqAuSmPXfFCkshVWIMoBThMasIThLSuLCYXChUdrLsTgm2Au1CtD1KtY0nDVRTZRvk2BdyPxBP
z4jeD5ZstN2TbWOXyb4J9H8CqUoprp6iRB9o8tVBy+av00K3tFH8KfiqXZNoxH45o5QoLCFXBkbU
AmmaY7Jq6zq6JiMv7FNEIbpWf9X9OM2KLYmfb17AhPp7IdlWAscuzLA3wCyv80EObtZslu7TNtWe
X2jVbYRVCzRspdyZ0v8RgAR9cJaGGRq1vyB3gC979ki4rAht/9Eg4Zoemf+kQW/geW3jAPCmTg+F
lAzQBT7YscuvYmZ/vx3VU+S2cVqpEgHGxYwyit3rbJmmWDrpM5MoEsPq8JMjBmRwarwuSBg//uUB
s1Ot+ZEUoe+1pn9RXl+DVTQwqRSW2xv6QTbnRtb4HOs4AfIZfsxSSqAlrGhPL79Ct35Pw6mcm61N
5ds3doWyiNGkkcwVAjtmBqj02TPwtj98DoOVNkAZUjjpNmBv5jOdNLbbyYq4mMHSbTcSjhNaHSfp
DTIFSAKYOZDkwzamr490YxDnMCEIA2Batbv5qMZByL6n98hYkTVNU6qdqGe58EK85kzuBGe7GDdE
j6sgFPD877Z0ys1pEDhGm0xgwYtFT2b6l0sSKSSyLY++urFBaCFZQt/ygYIKA5l30qcgyE8IIl5Y
R090AJ5g7lpYRmV/qA5moRLImd9fjx3STWh3llZZ/r2Hk6jvLAAhB57MKrI6V8k2ZXOz31U9/D3s
frscK7kHj/oJq1HzdNSqfZrA6aJ0MfwuZmKKH0RsGQaKNHJNyVl/e9htVohNw3iHObtbG0fg0aoA
Vkd5Oli78uItlC/ZANhqGW4pLQL0EFKUVsxn/2meX7J0N92FVvTMjLG+X9CdVlFAPAhu9qzkbH09
pbRrHuhKYXp3zIxQ+fS9DoF4ChyXDI2fTe4/puntjAfXeEQvwvkGZTltUIR2ymXRcgXRcQrj3Nes
vABN/QnheME7KDXMAbG+A3kVIVQcrhhZtIjwrIQJ0yZeixB6Zr/VePnY1UtKiynHNvEWb9vwuy03
y5/dKT1pUQ10HSzqHfu5/clFpMhZ8reolYwtOfn7jsJVKEpHtACU2pCVxP6TQjhzdYPif+XFRjnI
e9nmcFOhkFHNsEabMLm/+hTZdo3nAYQAcHkdOfpWfTEjz8WlRIP742u8H8J/jsTYn21TSU89mX08
D23KTVK9+WUAbzsN9DZ/gZF4EalG4C/jzXTFl+yy0c+PPevq8CI3njsbDAlzdVBce2o7U55Jm6bR
sah5XKU5UhU9s+o30OcMRYstDtmXFsycrAbsHQ+eFLoI1+2pWK+3irODFn1aacFN0JSMht9k1seJ
+MfsEeS+xbTo88RDAsZQUHqfvU3V1E9BSwPLqxvDVwaDISjWi3SLgTmd+7UABAUupDDLwcKr5A7s
cwrOD2l6O0kjO6tGTo2jpB3Bblo/9mqm9dGl4a22QNPmC140x5xGD0bfCLUU6DkBUIgMhdR0Wpel
iP8StOLokCejgT9OXfF35xbReVKjli6k6TViI6r+Pz50jexxCnKo9ej384rYDd6VWidkelLZMUO+
LtBZ3zSFzadMhBIEBbcd6SBAmF8tIEB4dokC0P3Wu3hEUzKDBGQ4sINtjT1w5WeFwsYtRdQ8FHQ/
DbQoLgVy82DvS2/SnaS78NBxFuIiz3eHfWMfPbax4U4Gx4ptCyEzgi+yf2jS8cHk24i3jFlQs/hV
OnFnig+y/5cIHlHZnsSSshtNTLSREp/aKHv6NRXyrmzC8dJvG1hlo0jzrp7IkqtvkzScX2z8DJGD
YAanUQ15MDDSAC61kM5tRq8lM3vGReaTuKV/RqZaFuNJgGbRK3vMffXr2kE4s2ME0pDzLsQD0rcW
q4dShQVHnLsdKAGYNxtiFxFr8oUP+SNL7Hl+LdyTNghlSrsyfLyhXPUgVM+K4eNKwS1CsSKIvDgZ
dK9TopYNCdGK70dZN8bi4Cl4o6LKMoYRyQYKRMm0g+9+X7JgjwtL50hZzh5x5oFyQXRz4nffeeQk
JPAqi7DLHr8SqStNC6gmHEDlE5AEwkSlc5+nsdiAcnQsyx1ZdNd7OLSvkLz7twXIsKfPxxibpk/j
/WEZi7aJGZTBK0bWnpMvFDNQi/X3L1lcciLKa8LslSgxcjkVVKmRFQ4ed3NuTymabSgTt5yLVOj/
MRZwjbrs3txcDvLwtKYtvlRQ0Lm9aH63GTASDi77LwpSQVavWA/FSMoBW54yxUnTZL6uJO5WdzV9
guPhzc8om411aCVTRW/VSYz5fSLMAgoExd5xZOMbaFc2SOXsfiqz4OcXnkNgHhOdGxE8dAUFXHwk
GxcuV2dlBR4mx+3QRyKdCms06aW1F4ibdACWFl2/KMIGH5LFzHswrxf0rETZOxc2tawjnk0e8KBl
m5uQR7XBHm6YF4hgLkfDkbKlt8GfigGjit/FXUNZfHajKCYDNeu/anUPXF8KQs7v21hos8pTLkbg
4zjpjBsNfpWSDK7OqenG13Ny4No+V0TAYNN2CcKRd+0WHfdAOEBdOpEAjBUiKGjZXMoNbcyT+vhT
qNmxvbjGLMcCaTSWaqzHaAieJKxBUBejlNl675PID8k02vv1vBz6C2vWm0Edxhi6Xpd/gLOrqFTB
QSlEwhM8mm0s1XTerWmvcZ1lkvTAtEbt8UIN3u98j8N4cUuNjoNPpiuUtn6gntFFrICAb6cfVlXk
XkBBqiZj6GVxpYLoZGTWD3uVJ983kBh8M6TLbcwRte2hQKVdCxiokFOtU/dw1e6YmG/04AAV8+qa
17gsYzALtDmQp0KpYOFNGxfAL/XdUS1BzuOPQ7skXVrgxl8+SFrgNncV7GY/wF/N/LrQdHtbIhRF
Eh5nJUF/ZX25VuZSWlXwICTFElQzHU3Nrtaw0+CVCpQhOiI90PepMaIZZvldda9awJdz/nu1BMpM
oO0C1VGstnU/IrS5rzw2Er26hxWruN+z/HwCp8WMBm/rE/b5r5r+8yUEUtggdM9sw5Q1dYeLDVSL
8BqvWKL8JJjcRUZyS0Hfrq9rv+MhL7XBFmzrD34SUT0jXtfTE7DdUxofO1ZHRpINnHvK8foA9+fe
z67tTwvS1Gxqtf8qhwaAJ5WDFs6tq2l35x3CqysUifYii71Y9pPUkJJfUfw1C6mi7VxwfNo5bI3n
C9u/IRaI5byIVVcq0HOzFgyN8nQFuyLNT2rni3kmFPkHCNL3aZugAw9BZuUuy+S15jizJwf6SDiZ
4Mr239vArhU4o0/d5M11Cc9oZ3+797c/J+VQgWRqN5IDbqHO5n7EkuRjrptZYmi2C/BLJUKhPNqY
rhVxE53QfpIOGc1/7iMFGvuL4kLi3RGnFDJsaIe4RDPKuyfOB3HW4gZ5m28pasnNdUmOqp2SX1w4
Wc02Vulm01znWuzeK+O4hw8I3hiGe94a/7ouDoVUDjMm8daLfPufHVJk3P5S4zlXxK85vOtSK1ol
eef4Gl6BRQa7ZmnX0OQ2rOoh7FxDfuMuryrb8bxp4Wbz6ks2Q2ewTBMPyVZkrXIiZjEso/ZPfIc/
Sf5MaOs1McQElySlykRUVgSsxIooy7ZFuFz0D2sckwXYqVVfxoFKASPrrR0RboOxw4nqD+a8KDwX
QQhKMvmUJAOXbUVeg+xo78u549cHoNTuL3ivtB2lX2nbkTJH0tFzPGzOlRk0e6lw5XADRMEXqx/3
u83gR2GsUDj7/sGJJep5ZEwKIvXcBORp5psHvrzibzX+aDVl4/O76QHuGbe15dE0sAnpbEKA5Sw5
t4O+c/AW2pT9oG3RwbUIG6wdN1HCQr1FkApYgvhsKEcRjrHK/EyOt9mC6VgLYnlXxmyv3X83hNmu
NxLPP2CAmZ/K+FZRguJZqYY4n+c2JnByDDdW7lKd/KvOQC5UPeQtMTDK9T/xszZ4cem7ohbEvwPz
jAo8l3lem5tpIyeGPffIY4Q+31eo/PT38KBvANOXQzw3h/x0wed7o7ozmpstf33uFQIBQNi0AioW
Ag/4DVlkWFsZkAFrGw3tvplCjRPQGZx4dWG5TVi0sSHrHHselnLN/XtEsTMyJYcPwBqd9FugRZ8+
wrrEkqQumZPoftIxPIt/xbrRvq54K96yCu94bC98cboeilpkjzha3uP04tgV9cPk4HWMV1oIS+Tb
blcoxmnAHRFgi/UAqtT3DtAPwCe0zt0z0U9P6ylc0Rg7Zw4k8u/8FRINAkuR3eV0s3OPrUmoEXu/
oR7Cz0v6KXvTdUJfCauGjQg8axQ9a6KAmwYwkmsIG3EgDdxD1y1Ot4rAGYOURG+iQJP3xRKeQQOr
E0+097Di+rXOho2jv4BFegoJSi7Q1zNuFrQLeg9pIVlYAtkySTraQRNLNUQhWtZNZ5Niz3MXwkZx
Q6CQ7o4pdquPl30EO2Bk9GMu0gFp3NRsc7DZf/026UJ1Q+11zWgYlvz54+Wj7nRJrPmO6tJdxCvd
aksHI0xCWAFkJEIMi0AnCqNMri5ubWesDw8wfj2DX2l/nvcXu+lDKwUDZXmc3vaGMrjwQCBL9KBt
q8nzCrheFeMiMzCX9c1GEp2rr2fCGXQs9La4pWnM/ldg1PE2vcnGW6+W92OQYqQ0RIK1lOQpIz8o
EJwr6bG88TvfNP/4nHs+kxZAKuWw1GO5M8kaD9MInfGrMo1btLX5fV5sjcumOIS3DQMDwWfLbhph
8gQQzox2HUOLlGcxGdvkN2M7/XhXfABTl68OrQpFrudShCc19IsxnlkDR+hJXYjVgsGb10275uu1
B7nzlHTIF4JL3QwKmKk1e2XlTfiq0i/gdk9b7fFx2jy+J641w9FhCPhue6kVgV3PuUPZx2Aa5Hew
WRO6bxUu9JbJ/B5vt2BsLbfbsZHbCUMcZvcXlOKMx1fTjvNwi61anw7BgVgm9ZystpXB1aRvKTwY
NvDPEmKVe524TXT6zCeK0O+eTTBncw/I9mssVHpYigT0gRwXyf9D5U4fvG3cDW9VDvCAJ68gHcUG
XNDTzA0bA2hElqJu+ZekunSIc3kSvw01IxoEHblrCYyiQoOD0Zv8QaPSg4DEpQPS/nbKYszFxQje
BR1zJwf8KR0wJDfvqM1/OJIoZeWGqyhYuFd//JmXq4FnsmfMc3q9zK1ejaGnwTon1dIUQZgvFmHO
n6rBZuIR3ToQkaVy7patRDfGJnT+mjV+vaF3dHCl15vKgtufS+bLAWcDsgQVaSbxKlDnqXgwhvm3
j5tyeRIj2FwM
`protect end_protected
