--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Cnj6C65kDnG09ZrETCuYW8CutMCurwHXmW5Jejvq/uV3yas+0liZTBkYAAZ3O0xol+pqdk6IkZQp
ROQkvY3Loi/jKs9LCsAOl3Lqu4M/4kngGXBf5/G2Y6UTQXlgcsMyuoP8WVikj7qR57UZMqLbLtKB
b8Gf7VSYFTrQI6aUtxAoHAM2liXsxk2hdwdawQ3xpCWjC8eA15qE+qlkXpqJZmsbs1B3q/8UXP51
ZSEYK1xVSTRZBvWET5066yEBXwKzmFKNUXCfQonjd+0RxaPUn9JcmlJF9/e//Wl8g26aUStcj0RM
aj9+8G0cxFopEJkLKtqqM+R/zFUlXkQW5PWMuA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="D/DN/WhAZoQ7Pjx2XbIC/+idbE/JjudIL7nYL49xHlw="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
HXItSq9gimRhy+e86vquwHRQIRoaXt/hHJa88YEEisB70FBvplFCM+feOh+67h8w7nts9l59Nd/w
ygMQNtnHoPhLj1ndSnp8/Gt2VuHm/EXJKtgg29q9IlCS49337zkskLV2hTnoEfO7O9MnVOJIvWXr
Y/Qg/Dk9ZTn0PlQqaAAcIYDW/Op/Qihl1WL2p5prAT5ZRBMRNypY5KX//txbPtDMqeRyIAvEPJBr
+W1FNX0rCDShmzff+iOtSxZE+i3VwyaNidbJbZxF7lxhJtprnpVBWL1guFkv8GYEXuybipDkuMog
IPY4i5pPikS/OaYLwG4xXDXylq/tZ/9nv+u6LQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="hGlxM0nNA21VoNU5X2mRZgKFRPqw6Rtc2+TVVZnzSTg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 61728)
`protect data_block
m66gPbsXGgR0r7zHD4W2fWYFSQcqZf+BbgCuKMyfwiHADummecBG4Fo4Cnx05ctd66dWcIZiyv3/
kvWu7LkGTcgoyX4eI2FcjO6oUYVcwCbMEihaqzOo8dxGsNiCyNQuRBo5JYqqfNw7xLg5R5t8+yEH
m/XttuxpKW58a/DX9ZvWMESM7UW87WR3BHvzeHWsW+9MfAwOROII8Czhh2VpxSVNrK8QIq/kgUc5
Z5YSQL/aNXt2dXF6lqNNim6nHVM7L6bnrhTGW9nsthWQrJe5XKH74GFsn7YW8/O5iFJNN9FXVj+E
NdQ1dmcx6DjCKfzA2e9kzo7jJDTANUMSPH5X/sI1lu4eeJOVKII1cZzxOJSrbxxxMGVahcsgnpm2
XD/22m/15mAurXDnSzyDo79OsD9sZMKA5KcuHDQzLA8e1S7u+Hyo819LznyhNMei27RZ8vRRlaRJ
mryN3TML+Fy1osMsbetq8e/9mzIPRGrb1dWmOdZULcEH735aHRvfkCxnCBaoJsN0Z8vop9M3jCPv
pgbKYhb7FT9C5+Qk2rfIkYD15aQLwElLJtBurJT0CeAZ9PzMyk0V858kQMxaOtS+32i9WmHKpPOs
17qWLh7tVVHQeCQ7MzsVMHewSM080fgLRzt6fdkJ4ZV7ftyUS1Om1H/IGU3/ikEmnFJyBgxcG4m3
Tir1wSISPajzQOqQB0suODaPi4N2U0xV6sOr51hMz/Z8Fy6Ncl4uxukDqdV2MNmvBPRSRvmawz8Y
DgLsUnNByNIF11lkaSw4dQ1Ck2uH9se42oDLNlwsRg6Uv8ZkC/ZzpwFxmOPm4oZaKS3Ho76owe2m
jfUoefDqc6nk4mOfdGA/45zaUjE/P6YKr4Bq8ShUva/cY7xG6Q4zzTA/3KfcUYC3Chmqll1aG0fb
lZNS0B86oqsRGzgCpy/H5lKKAfS0+y1cAQ8lad1wuWga7HG6wqpTWRUI3FWPfQky/V2ED6yh+N8q
b2xtnLAAdFAJ+H1vj0hZw4TSsnhsjOrsRhSFu7g+6QtSVK77N/vQxYeE70SrP/AObthEvrjYOIeO
Lgl9FZcCe/pXnwqUPc1xM9IlzxvTBm+sq2ciAh3K0gvLjbF1FKWGD9kW5DzBu1ZjqWOJMfnJwohS
FmZ4lE7k6k5UBKUVguQUKeAMrPgYpvOUUjKvvMDn+go2dxnHo6LCecGPWLoJsfQg0xzyMTw11CPU
o+NlSgo36jGFKMkscT0y037JXHlBYAk+33tY1QI0+50LwiLDGE9PRZtLARWPmKglYijj6W+D07+b
AsOAPefJV8zuK31G+DwX9sRHhZ5YOGKJxTkjUORJMquAJfGWsxdKqcdIu2/WfGDhOEFbv16robc4
qVoeJskpbMuEqTjsJ3b8dksLe0M8b/sTe2taiK2ASD3J9OoojJ7i4Qx0glaO66WyCpFbrDg/rsXm
RljgJOylINkTkvUUCNbA1/6cHiWrzyfluevs2dr+n32L00TuMklFctdU1igBCK+7ELjIdOOlQb2d
xY38RGd4Xn/HsicbuCEwoDJ4GIxvfMYWcjuuUMtSzOqHb5YhQva6A36XkvP3nEW0KWVUra5805CL
lm6cqfqZjMrS6/8NkcKE6tb8QaRjWPudKpM5+Vygra+dJgdRzatP1PtwuVd9Khgxe3yA6qIj25hD
DrrMhOIwaGqnbsrHGwGubZD9Rubzyyl/K0VxUXjClrWuBfWxFdqtSbVendFbdx/Uq0AfH+4LHtXp
dGKl9FZqWulKwBR8kQ432jPwqWbwS1XIpT/AHgY0ERm1KMnVw5t2PVE9ON6xLJ5fYcLGs44C870S
8anW+C0h5MDKvuY0Rgd3VWOGT+MS8ohxIb/4LQhBt/UNykzcL0afkZem2rhsbwcRw9vCp8kUqtGp
YmyjWKorRm/yqYCULM5IKOMWXycRN+zYnN48rP3ra4WhUH12nkLyvyQEHYzqow8IOknB50R6iCpH
5qCxuVYeZTqIKeYnxgodciiURiR/iWHp/qeobIp6VZZbjT3WQZ1k3d4hwxQuzJNIIR8B3+Nxh9LU
fQdCTBh0lnlEYUZW7h3UBxRmEiAFCLdhYAOOVGpvszcFO43jLfy1Yxdm0Ol31IfhGkQ2pj170LL/
AuOeAQyxSVbplv49xMEZ1JaTqW0mLzLlCfxi1U0mNzTblpElWhqJGb8ZfmBa74KaGB55xlWfVBhJ
phaykBbvBsFZBCH3GaSLkY3QgsHjxyhq0WB2pdWNe3Zkh3U/wxWG/TR7WTqQ5p1i29WpH5iHqpBD
EOgGQ8ug0u3SZyq8WO5RTMVxClJ+3VmoMXm1Q7Hv58imw0I+GtenT2d0jElml8zqiTXCGqzCdFJ1
A4nMTmGcuptrfekubEIP3zAXc8eiHVawEsPvhkd4mN7bI2xvPZcbrmY3G0DebG3lnCp3qIy46bHp
UyJ3GPS6B4SHir8TFug97o6ann4c9oA08fZOPdx5DhMYRzqihLU+V2TDyxbDEeSczhKHemj9OO5c
RykR/CdhomexEdvXlGz6ip3WlyQR8zxxXCeDj6D6mU7dEf1j/762zB3zWU32jTT91iHafoHQf2FC
+RpPAhUUKJGroXBWfwaWJ6ZD9/XNY9/MqNJPWytUBTJY7lza9EevFji+3Ui/YV4oPPcCAAqqKoj1
Zyxs+mNlymWSzFYBbaI2th7/kzA++8D1dqPkO6531qpx/tDkbYg9XBzw6x5JPfTJXlkQHA7JNGUx
XRiMo7d8MQQiSgXUimDIbzMIDPs3YlByUpaN5oX4Rvc1cvaDTfoef2GEFNw/TZ9Qt23ytugUP5Jh
1jME/m6OTS0Md6MZNlysfK/2briV/8boIG8MdWa3bh6EoJNKA6UKrvBKfAVNrTlGtgr2jyINu0qN
RLtKS1eV2P6eFRNhr3TBN5WRekI2G6lOjO8ka9X4Fgjy/ScSiFgZnPtFj2YYEkPLncxOwKnMA7LE
NtExfFAJeCdHfrmAlhINrNSjyDshv8VbFVZFHpk1G1rpgITwau2XPESUb/VxWO1I+Ys0jV0T7Roa
K8YcaFPS9kltJStvG7FxwAys5edlEcKqBfLstgsG9aTg+YLkXSEgQNpcQjvz56903GG7bZCWiolE
LxVSyruUpxHOxXBgUb1NlScRFDzAhI4KzCgujm/lLDPTaY7BYay2k5v55PPro4n64guOCLDF+tEG
w/Uryzn4AfEIfzThF58sc9/skDQYp7tcLCVhg57KREHRf4FAn+35tEI5pWsysCS+pe11FzXhNFhY
cc+MuI7Nf+kMCLCAl0Co6ouqMDHwTt6VGhXq1wIxIQ/ZiSYJOlqrZDMc163Lx+Y+Ym/mPPTeLBg2
O50KWwrsW8p8v8SBWbaKqBHrwr8mpk7jIQKMRzl2A1cPhyuUjVaFOOvD9qytvbGqsvfSjEhw9fY/
zgiXnauO1i0DZKqFTxOVwU/B7rSbuRbAxWZlto70byHVTQC6G3boYD/Oga9+dCCX+Ct3odxqISwg
lGbd9FYcxl2rvWeo8T080/vTXDuwUd8y+H4KpVqbYtAJBTn3Tl+iGKNgMtSSmrrNU27+i9W5gqaS
qmIygGQE343RN88foffC2ovylA/pscjO0xDC4EY+ENg7QbWBQCQ+rUtw8/V/szt/0NpLhujhoPUL
OCfd1EsxasPRSvSGmUZvJ84SbAgDl/EyPFvpCIk/C4DSpVtXnaJ3dz9w0cdkayXweGtHdvF7Q6zO
zgWdn82WorBz1+WPQLv46Qre1dErk8iEwRNqQaagljblnLLYHpfoyGNPhBlwbz727yBcVXLQ6yzq
QK+9BKbtdfxlUqDZWbl7OJXsBkFhLOKTUf5r/SsiNgCuvZWg2CMSXbI3U4GCZ2lykNtGc1eWktxt
gyRxy9Szwijm9ovUiCrRSUijh/mWbPvMKUgkmocCBvvwyGdSEELpKAvy6P69Xl8NV/QJPlnHlP30
BM/seZmMqrop/i8or6dgPKpat/iQDjdjBUW1b7EAxtd1Aj5gnm2H5XXze7mhW0Uch/DmYYWooDND
/wliiXtDkPBe0LBqY8nWoI7VBDE3u7897HQJFgfotvURgm8M3ei/+JmAK90Ur237Q4cjMzoxuLSf
3tsI2+YUQa2ol7pdDtv55+C151t3Dvv8cKXvQJAx6FHeVGrgfiaf27ngUToDCm7C5Mx5NbVP5TFK
eVAa93qtaoTtwKmtM8BrDvpFlTcCSPvzcHm/0xjoSgmZo6tDtrfzNSN64I800ls1y9jlfvQHyxXP
q9gtsMNHmr7cMifuamucIesS2Z+OoMcwqmtx0iKlsYklPm0QCc3+UyPN0hCi9XutQqv/HnllMwwL
MDu08F+hiKXa4PjCxnrxvDZPNUJwUL5I87US113+UIyrOaXykaTOlAEzczCEOhyuMjKyQErUm0cm
N+tTtZQLoR0Dl1VUl2BZA99ZrOGJbjv1rzIxQEK3L5kQjhT/9i50DmOPYvFCi132u7Iy5iG0EYA0
4Th/Ts4TJmcCIG83ltP1ydj+9OrueF+lIiQFEMK4zU/AV+DII+J9hXawv1fEcs3Fa+UnVBqdwKut
tR4dtFUV2AsndAEkSf232LSyzxBG33TNK1FuPuS9OrDZOKGx4dTCLUTn7ALJtxtPDVQDq2fP/9zY
G+vyqvHoW1GUioW2VjmYwTAsYYjaDDWQGsP0vpkrOHtvl8XDU/nSk+hF0hoWeUh1Mu/8HaQXfzeC
sxoWmLHJIbtqes+LY+fUzdjY2vLIKTSFRn/zpKn++lCNowNy+U3pIO906zgnvzLhgQWqsnl1V/Eo
3NHiHAHPUIjUfKlqEebpBTHhTejY05v7Ut6JcFBxpF07fk20eVirxzkoCIr4JS5ptFLcqj+hiMD0
qamR0LOE+/Pm7NpR9MPJ2suNpSC5lQPyivewSHyoNBv/FLCalJx9d5pkePcWuBiPdM660S/NGFX/
gxUruQzdkl5xJVlhmIg/1CnOkKEkxHC0WIqr2/57gxfyfdpL1kGccFpZxc80L9xkqR/Xm/bIq1FU
rwyfafGRjg7WXmUWyYUikjH7l3PAQZb/GG7o4nlFPj1crEOQz/VoIeTr/gr28fuIj/NEz48zAeCd
+o6CuW4jcGm394E1bGl8TbYlbLXOQMSrwryP29EZk5ltmRas7/LJJdaZw6M/HOiubzpzCuZIuonp
x4ikyGBkR1NuuH3RHiVTBbUbNzl58VGc9oL5YHOA/iHI3euw3xWygw36ttayrt0tPVGo54enEi+y
fceZxBsgrzV9VGV2HsviMv/vRCQjan0BTZMzI16s39lIpYMy2fDrghZngeuhpXGxLAMQ+XOGlAXR
pqNTaQlZhCRmaFLTvhpTo6G/rs4IGffiWTk9KZ9hugPPTwg21hN8isicAhdloIedSD/NlAj3AjeR
rkb12X5+H5MLVig7MJnKXu3snvfPrNQOdcCv9vcEeClxXEUGMukB8NnZZjbDSAGtIFoK80VeMQm4
w4K7zoCId/Om3URZ6eaxbwlFaYgT+9cX+uB8/zDnztvo7ruAuYxZ2IVq/ebLvgjZj4FJU8iXz3om
uRYlt5iFWHMPH7iSMq4ntt9JsGR5egEnzJqZQ6wp7xgQaZcTWc8xgCIEF5iI2hFyZHdVWPBDIBWv
dw7OmgCPDtpj6bxcjEQv/HmbwjYeHjUviZKn1PuVes2DfR9D/duw1XlD8uqE2zzfwdS/dkzvfYq0
tWpwTABuRwSnbnBcy7HvJPHphxacjLRp+KihQS2xKsTp41RMXva9tjMd7mUqiQMnQHw1tJKooiI2
ZI4O0xnAy0DET0uboxppe75/SoqBK/0q25S3YHvHLNMPQqgSadcaEcG7oAmoRiocLVyGisMAEMU/
p2amO2ioCG4IbzwQEvYgvCSqn6NMRyGtKc7tSyTlkU1PANcyAvtmx8lBjjpJMrc9uVcIjnq51kcY
Jh5eP2iLvHv9WRpr7TryGq9Je28JtmjtmWMELEu0o9zXosXAowap05rDDDMvF98w1Q798duvpBI0
fo2czf3NWDqZahlNPQXSZ1UV6B2TiObS8YTfHhWKmryALVyPr0XTlgU5xdVO7Apkvz2HuvU/YSA7
g0PRsWdr0eLpsH+Nb05Xmno5T7FMiV+Mv6jQmKIjsw7eBpR8K2Pad/fiNH244sV2d/HTBPNSR5Xk
Ld6d8yZLMaE4Hn7FgqkOpZmvNKSCp4JrKRNfOZ6ong8D7mdpyM6LldxHiUurkTJUUbMQw5Wh5KZy
+iJn+6/DU8oSAuHcK1o7A9Vn5H8voPTD1GSluYNbE6VsVqCeU5esBBgTiPCRbFKmrmC2dKTseynL
jwxE7k8Q6ipwFMuwDSxf/zvK3vn6pseRAnDyATUc1nAIpypaBD48JaYdRJRmdOeDqh1Lm3iAu38p
a820L8Kt/bN21gH3UkDuEKdlEO8do7PnWClk8MtekFW6goaHHUw8t7+hqrLr2p1lbs9KQ1y2hNW+
46khn5CjaZXdjv9R8wu+3Rwbhx8GvsFtWqFfzEGWBpKwFnvb4NW0GLrSAd57V6o6V8+t3G3+QG+f
xnxWaozu1ubVuzCQmjNGmK6LfuGOKjfehczdIEvjHtzeQuKWwVOann6rTvmWAk4bSxpLiHR8EQtt
ibF8WvgZP8FQlqXPVP+YNWEioN3eTYJkid6qEwfEXXNS0o98o1NSQ1l8cI4viV7M8OL9nDodxdHo
Jam4gvuNIXU7EWZQaekAH9BBX0lXdSMhCVRnyX9LUtUsaXmceI4N+d/17SQGORXQM3swhZRedH73
yUkNetnrk+USLdhkAufFzgTszehvDl0wq69lP4OYdxq9ZtD+gh4dDhz7clCGBUcNn8D2XE4H4ATS
uEh49Y+vcnKRymf9i/17jHhgzaXy+jJdsHXbiydeScAWvJJzNM9KhPZKWcyTqFzgcIGU5hmDHYOb
GFT46lwT04c0Wf1GXuyKPCP+a4KB6rAabZClIsQpIkFuSv+CMfJngo8+hB5jwgj4b7c8wnwueCYb
m7t2/eTtrJG0QVO04WFDQ1F31PZoSLdhZDF3hllA4KomzNkvceSSBXjLXdzQpn6sUpMWxI/xx4O5
DVFUpp08qOQ0U/Kw5fL9uyVAmwoDXaCAWvgcxs3lT38OagMpxvABK/k6+pdP1fXBzElOfjwFysAw
9JkgBjYLyCuQbu74m2kIztd0mZQ+fzCGlDkU5YuNXncAg808myZPghjzi49KW5JOW2zrPQ3RtEHE
G5S3LlCRTxHLV6GPwQ4mUJRaY+pJyK+QjyT+c4f9hnA0id6TFCXtgxW0+l3fxu9N7U49t7BJajja
LKp2rBFhre81eNr0+l24bRZ4Z6JouHu9wnxwfY3Dbrv66rCSRp+JSYlSw/pEcMSHMVd1pm4aWpRN
/68R2ik+FKTLT3fpjALhqiDjkfvFjfz1EhuJrejAfh8nmShFK9k3JR1y5absC8DrePVCcXWWFpFw
YOImyw1ZHdcq7tVsQ1m5ERS+ZE+NjZli3MWVk5WFdcoZ0v/NPWgoDagUAr9gSO5OfJvQJq/TmBMn
zuifYejQHvLBy/2qH+ACv2y0YySlttBk3kxyK+svJUEMrEAlFOOZjKEjL75jASPLPEdFIil+zwFb
qB7BDmPHqN2aWzr4LSp4tkqmsbayJEeoNgtsXjkAh5U0nM8/THaSn4+nqoAkk1/fhqazDSTU9M26
E1dk15gF03THi9+UWgRM7frAJLhHRM2cYPEFRyEuDDGjMkEf3RRcQJaX4vWiorGbs5qmCIM92I94
2pOan2+muI97RgjZEu+W/op80ACH/nYDinXOXRZlu/QOcHuJKjnAt0Q7Vxh29w4WmN1dcathQcAs
CNzX8x+LoKgFrt5ZuVun24guo4SK8e7UMalXAoDd0pLyt4XtSFFJ1VNcg3Q2yyUjRSEuUAdJn8Nn
on3n7plaa9Jk/h/lkXB6Mqd3pCFTkonuRcQ2gU5p4cCPH/dzOVSuYRKDBXbyl4GS6bl6m3VOlO2s
Rqb5Mycksy3xCpJhJ6MV4YI8A7iUnn7/f/SXJ0zOt51QRorWnUlQ40fTShKFtycwLcZ9YwMK95EO
S3g1BQ8HiBuZSaRwtVggza6VcP7rNERk0JhnSvETDOkfSVCQHiUYOUI3bUR+6CI7h9lbmS4rI8PW
dxxGSzKPIGCGvGmmRZY9zTuQKSNuD1HzIvE4rAjaWiOKm1O6uPKl7a0T8IqX95p0io6w4AHTXXXD
uNRY8FVc9BJ8S5QvpYmDRITtRyngOAA4MWRgVXGtrsiiudiEc+MrQKe5Est3tORBik0TXjY2iXZm
oykxf7Yn+Ag1UAmuqO6t3o+5M+NntebmOw7R3oxV438sfIMrOR7Njb85jXoM46IQ+Uu/7hUJ4dAD
gjAYM2WEOMWBCiao9J4puciX5mUhrZeEbyTP9agojUD55DHLCgEUcLOR2eWltOjD68rS9pkKLv5b
8qvbakJtTtK29QYaNmlRp0tvC7G2b5fJPRWfYVrhkflDgRlsMioAS2/UQPfoBRn+v4y17bowj5Lx
NQTHnZ7qpduyUEpIq5NSFtCOeWiDlpSVueOQlvV6pc6x+640dBicZn1KPhJj9ecNTMQdZql21xqP
FGeN37gZxyCLOuaYFOxsPXKRq3ZqcUN2ftpONHVmLoybQ705xyfGxHsofwn0rRPifgSr23dSF9xP
LrvLS2bG8nYu9C4C+meXMa1xD6HyOYxbeWz9jaBr9XTwhv76/6zOyWSBjgUvnT5RRABmrqDm9ozr
kOvhtlPbXeiXKTYS1AcQKZMBQHQcFjrixM4fOq+N+xCmu2L2u42jmDAC5y83ahGF/sLOEvi7tr1+
VJo3AI0g1QdL5vSevD2n3wH7bVvt7HW04DScvwpEs8irSIqA9FN9coiyc3IlkTwvlUhiEX8U9CoH
PteTF5RX7BzMcBOHxFIf5fflFf/6YQet8X1Ieo6ovMd3TNG5DdSQi7/WVyAWvxG+gOgZJ5UJ9iWD
uwxjfr/EMXeGwCVniGXoCId3hX+aQ4mvj01KqW7UkTR+4O6XozS0YIDdY7SX/MBYjHuMK6EYCf1e
zwihnF13M49/KAfB7bwjvlmaNd57A+Xk0PbnNEmoCTKsSfyRDrIiXAUu9nUZp45V7HYa15kCZx3r
0DX2lP6r0f5juos+Llrx/TDnkcr42JVtEbMI7eQ9HSuuv/FR2xtM/K/DMShNdy1SIY3SQNC+WKWR
xBceV3HOhG4KXAaoTi6XGtWTp5/Eq6QeHRpGVvKyRmaXzBtQp0uWLZHQISUw/yn+3lbPl1vojJeq
f2OY8K5oFchcdazkwnR4CRpn2x4Z45uKV8X8yPgZMD7N/p53Nl9hxm6zS/A6nJ9IKgxPuBevbWki
v/1UjpyDczbZ9BnW4CdS40VXR7v23wAQwFeLLh73thUQ2YXpGTuFHJWeX+XhbGlPKM6X/+KHU7Kh
W9mIr6Y5bJzTp50mzqeptL6bCXjQaKouIW8Uz8ESeJdrTDZUMKPLxCXkAEe6rnDgwJaQPz2IlWr0
EBtjPdk1Sx7rQzbuBHU5v8a2nxI4nQH6AZBdflLuVNgk+83nAlPHfOb2ODDa4T4Uls6YGxhZbkGs
315IcHh6++3p1nMx69Pw4P+SFOS4tHOJiIqZPmMMkOZk1FZpJcO9Iu3h9dRhhhrn9/1q9zzPW50B
fLJmtojiNkq5d8S+c7dNjNJ9fkZGZEYLQr0Wu4FjUeWid0GKCvwupuznpgYQx1NDquvkevy1nAHb
kMntBnYO0QVnQaXQOqA0YO+X2uLlQplrswQqfp8V6+b0SxsYe+3ccBSwWZOTduIqvr1rRACDJxwR
el7wOrDqCQBsJsDSecgG69O6LYw7X5fXL7lXBTVjn0GSAnGHcxPkdzReHAXupGixqwoXZlHZBv3q
xpZ8jkkHX45WfpNa1tsQbVYlwJ6yBbh3tCQE6UVJgbNYe2OAwBPkLMq72+EVthc/tkyAPMBHUR5d
WR7M91mfUuznHjBIzojqffuJBT+1ld4QtvX95lVkulL86NFZinHqhhMhptmio1g0ZO6kRdMRhR1f
8iz1rDATJqJD8P7X+waFLqsKDjWn6EDZUC581ttnHT17lOQ4fCYyQa5BbcU2CLBm91M8wGBTQFbc
+l1p+5NaMw2FNiAmTtPM50H9JNDgS6votGopHCbByP/RGfroV9/KTmlMNNzbzky6GDx33QXeQCMy
ntwHpImAHPToG1JpX9o+boc7xczjsmJQbnQcXmXz7V7r7r8BEA+KGB3jmsi+mH++fCETkKO0OwXl
4UA+eXzq8CPcVsk51UhgMk05gYWNvFwpzmJfRB3Xb7VpItCkewf5lQvXhu51axnrN9i0QhE7rRnI
MvVBFKse0Aa2SGg3a/3nvUi3WbxxNozoZ383+PpgtdhHB2iUpzSmBfZYnQQG7aimBR+vuCLi6pys
/JAvq1R0yErqpfJUgx0/H2K/wupkh3JSh4ReLnu2A/pydNMKTLbFvk9m3BtR+gLBv1osJxLEy7+U
UJBlGg1YFB79DAWXN85rq7f89AIBOrE5PExVvJ7exON8FFRmG/EpF99yTkIdPsDvySHmlqw9vmKq
Z8bNqx3VqtVB0YDE6+OqXXeTKtlN4WIKMkVl5k7gw4IyeOqlaQYuiMUfuG8+79scGx1O4kDvJdNH
eQ2D+JYeXb/LGZxLwQBWBH19+CWk7zC0SNNM3/oYeQfAjXjqra5kR8ivnq3DC00JcEoMs56+FzIM
HMp4V6EOdUwler5GWwCHVcBz1XID0RkCOAtjhvn0RrvzbWCKyI/Vnor4I9yaCUrRnlZrG+1N6+4R
PhJKug3HeKY3vtLlOs2HkFtO+McehijM68o59i0A2r2n5sqCU4vgKZSiu+NGPdK87Te+TSXy3nsX
DPEmOjVtKLG48nyrOma8YfOc2LM9sfczk1k4qWH0Abe00EqyWtj44Cg4ejlWJSTImClbP3edsB2n
xQDW6DTY80+Qq6NcEm8zRZU2qkz7dqKZ2SDLSDswj9R/5XmMbaxSnpSqE4nAfzATSBtMYd2pAGFy
ikJ/2HZQEgNbtjBo825OetoBFsmPmIKlayo/cY+m73sdASHp6BYvIvmwdkj38DfSHeZz+tScF2+f
Y9zUQLebaPFuUBEAUsVvNTdYLH6jsaekFJ2iN3beGzIrWW/aDLd30oQ3VtqZt3+0VVjzql9Rd7ZZ
bjnIjl6U2QD7BPEtS0Nu9QbhjEFAorJbuVsMBcJrrJzTaMhDXnHue72RsiQE73qNcDBfh5JCaxx8
VwxPlY8CoMW7m+PGPOu9r9ebwdXlaccEN+gkK6nkHwOKiS7qChO/YS8gxcewJ7AQOKQUb+DgEe46
FfbvUvaeIK2yunACfeo9XMxFDenk/LIitZ/OzKLqwy2j8demUt4eBHUozvRXpjpjX4QoB8dI+vcs
Q/4Q/523JbIecq/cRQsySeVG9KqDo/huKqYiewWf7LnjW3hA8QUnuH11Akm75ogtxBSrb0evR4WG
eZT1/ANo3dm9FpeX1XOm/mN8sELbEkqPXtaJOSIwQHDPELQPExhCVDS7NRuN4XmgQvsyr/tyia8r
0CPEhZhA5bQ1IdkU0c7UCs8+SuH/MOeoKYlvxr2t4DKcR9MO1Wo0MC+wpwjKvEf4VGAaVEayNfrg
qTQ1tSlaAq+my9a+30RVMCuSn6aGkCIsxjh98zQtRgo45siFJsa0Hsqe50q3T4ntuYQjewLdx9fc
sUBRVJD9MsVPiWjWhvk6X1idjhwoY52MJc7ERrCmzCeNIkOL5oI/iiEPko40kRjjZSmAs4EFIxlc
pqHYSmAx0glYoU+djKALgglEGqAoH7LwPlhY6biZdoxwRQ0M6F+Y3zlUOlxsUYfrEqe4MZ9nD4CJ
OGMR6EzJLF5/ql/yGLXV+ee2vv1XxRYP8tblkNUBaWrEZTxFK+o6NzltgDYFVdkxEw9CCfuejrLL
z2iO47UPixamzkhdC3hl2M32MWMD1KHnEftCtZpPXE+PTw07m8PO6+eivH01eFeKu/6yScKHuWar
12fKxXMYXP+WyNM2KrgHTa4bONU4UoJsewdioGFB91VJN8tBIRHRMsTetV7FTrp5650GdftSKIYq
OaoME7dQAJmk5iFGFtSYfvhYxP5zqN9zscY10MHp68t2ho7uJWyChscN++dWGuQf7krMq3jeK0IG
o0mDUF6YGTmS79+H/Fp6A962jmNLK+l23Ll70MmW5sbUT+A68HiS1UDr8buVFMQfkGff25+8vpAE
YhhINDvkhswjpNfrmmV5g/+EqKn9+JH0vFG2XWVABeOh71Cm/maUn5bL29BhaIBvDfDsT6oLOr28
gOIoelcFMsGf5EszggkhtTJF611g6ruAZiTjzvcHAiZIEg0SRBlbk64xVzBgpVt8gHY6vAxw2Rcs
k8ez+9zd/D5Gn9tMjMbpqKxfcCovPqOxkttA8c6CW/ezx0ycZNzw0QyE6UtN6s7Dmpsy+KaCQ8IH
9g3VvSceGsDXzloMIiIHe8kLc14y2Ccv8xSV5mhvgkkwYCUzUnDmjhbhNaJqdB5IyYqdCLAB7Ms1
0ljy5nlFtd/RUaGOgRm/UQatrJ2bWdgsq0064IhcmOq1Zb03GHJHc9WT0vDX1cUTphi47L0BmYEI
l67zlMSHs+zzyomeSYStRCVAPhNLvwz7okfE8mWia01gPnsp93cY+XtIoIyQrEDsT6W9HkTTKmWx
xmu/QDMQMdeQlezUDpZWwnMnbpDw2AohSq7wPgnYIb5ryg/1igpMehR9TfmhdjIc55BK3SqphjsJ
hdJJBlOi4z2XxntgtwjfzEAG9v6oIPpswwRDgvecdaSlbHAco2yle4cPbNSaybLYxDe/sU5sejIA
R2ufU90P4Mj6XdVjSQ8bgWf0u7Zo+iEVUjGVFD88ughgJpL/WORivRpv49oycwsxn7V0hAFBdUYg
m89SvrPMHBKupA9FizKVTBBoqS8Wk//pq3nLbF/5LNmWMUO3qbceFUX60XqzaqkIM9B8OTrLXLwL
sr8CLvjdaBWlr4sLI1nZ9PMZVhiV1bI1/BV2ha6YOXwuxmW5X1JGJV8qz25ChcFkXPrRtY0IR94E
aNN4zvN6DwBaUX5CYxS8SeguGyjnGnoT+fCHfQj/NgYWeUBaU1Wqr1YeW1dVNBrSq614OQPEVqx5
fzg2kzsFNv2rxIScKefyT0PF8mZz6mmpzt+lnhbdmtSgzIpFW0k4rznDsqlTDwJkU3jtN3y1Nva3
HElb818uWhhh25oL366ii+s0Qspt/HDT5ExBUvtXLjg6NPEcyek355AqDPUGOnpoPUqr2mJ1+3Kl
DN42NmwVtFyRFMsc/MsjXEAduYxMkgnO+5P6yr785GFsE54XcAKFXvPy9vS+ZZmvCMNzxNFHuHe6
DxmPAfsXsp/Yv5TjcRcgHN8J6COSELEOwZSHEg80jmbtYejn80HQeFMr7PoqhWOrpHRJqE1cFz9v
JGHC58r/tw5WzC7gbK+cPjLEtMisaAsaDHQ43ueTI2mtpJ+O5ip72sDCsKq1rTwICCeO0x0W7lbu
2FXxPLlIi/O6lq15s9oBFpKke2g+2YSul2gUENGItw9aO1KX9rxLDnLj+aG0lIvgAzF/j1PaTZmZ
3V0ksalbTHr/96IkdQO60i1oEwtZJBFvQ1G/l5z3fk7RtvMKddPAyOeyIlzd+jAlTdXl+YMBIrsr
Ptq3/BcyW6IfbzEeAa/T87a/xPzrWqtUM5bWJ2vBaxVQW29G4HYfe23p0fRRwJNAjnW3JykIh+1e
94rpW11sl/V0cNJxioKOAX7HaHKcexDR1xsu5HFFSWTQs5GkA5+YyNecr8RjIYgLuTdoLKnIkqQV
R1vXs1Yj4vt/GURGDIXcLFXN6tMMOgJ/gO0XoPu5LXRPucySPpDgkkqRUI0L8z0L05GTy54S6ss9
AGRiFB5xbFMp9/H7lMdyxTfurrPflslzfZoJXeqpiBcLbVb8pa5cc9BI1hrHEhrkMUAavkbYavy5
wua7jpyWwttc8eNi0bVxccvytr6MdxJHTbfjnPPp3agumqNjfzSaKT2hwbhaOUTIi40TcjFjZ3Oq
pDYqF26XD+t1Wfqjg3tnvkQn+mRGU9MNPK5Zgy7NkbCAGNnj/14OLiw8ZxdurB95fgkmPIewLqLL
MRr/ZzRnoQb1solWTGJft3y3Zz8ZvOZGABugBkjNIh5qbNxy8O0ECwombT6VhpQ7Gge9weUPH5en
1nl3HpR695AkKtOtXMX0z0z3VP7OfCiJ2n0zCupe17E7iyULgHCu2ZwFi7cEWvHsRosC/6oPC0g5
0L6Uh7olcm15cSvUrVg6XZO0AmmOW/F8oBSkalEyzBL8rdKppoyJcwkUvIj+O6KwSVk7BPGdeofR
LcU8gVoDlse0gf1xEhY21pOZ/g0Xs60W54Msh0MgP+cRWlykOj4tIIXy/dl+HZvSDEXBy6yWYvP1
NB60bhTr828rI/uQ6h0Etui91614rrJNPqvIX0jJgDGLTWSrIUFNNg+odXbhxte53QT4dmi/jhMZ
Bsx2l0u2hReiz3ZsnQCHLdOvpjscwKtM0qgpVjALAqsqIxWjMavD5w6f+BHQGzuWPQsTBj7KCDJR
3mFkqKA0I05E5sSKSoGjl/VbH43q6eDI4IiCM7i8J9dBp1H1MV864SXcm+R1gQ4R2ykOkEcqjIFQ
y/cyo5zVSeelIeT7ukNTZaHgKZckHc33kqm4t+FHnPXFjbZkwqxaOy0/v7H8KcnjxNIHskl4SChx
A6ZJGn8Bjxe3pbBC/kdEQsFt6aLwzINYDHfXDrQyjyWDJaJu1oToKv1D7DStleGQGlwKnRb1WrxC
iAEVN13mrVe0bGxuKIXnB919VJlDSFFzWX8ldIz1YiktJV63JUVIgIGwtqMT7xb3iCMH6HMK3i3+
/5EleE8gRqpcWgigFQOyB+WruUjWj8l3DfmKmRwQfpeBhMI3Wutz4E4YeJbCK2yO2YXGUFrFCOsW
LNgPM0EornLPZw3NGJZmKNlM7Exd5nGSySTkNQbc+Y8GSR+NqfqYchv8C+iUv+AvnQ1CB+X7jLYe
VPoeB1m+KeflpjAFcr2GTEIw6lfegxJ/C1X2mTr95PhZfAm6K95WOx0iDiMJK/EZTvfedy8Ls75Y
Xstsotyly0bUJgnYj0sf6Z3Ey5IaocVQmTk65pBHNaeqyW6KRekZ2llNwJVAZUAUaCe7zi6ANa8n
6Vi4YwatoRe4wkQpvRHU5Ve2gSf5F6Q9E4xoPwqBqlYaXVrpgCc4pB/Y0Yv8JOa2ofjZANAt84Z8
4OcwRf/bcH04wZijfKOfxzwMIraaVgYj+yT71nSzL2nl8W1lAbe8mmcf+BM90KYOHLC8BwpimZVr
Zofp5HVjN9jBbsN1A0bmfQCh5rF1X7TYo5U0JjvAiWkOd1SmBMib1sqc15avI4K1jjolDJdo0hyK
l+fweL3OWq08e58VR4JP8SSX+LE8QaA8Flf/eVkeDVjYIfH0GS5qb/dBNqB30Pr0p4g9fdxBjHJL
rZd/Fircwr4hC1c9k7/xx8gByjpqOMht+y84Fcvr7yuN6fL0vxri5R4JWi1ZNnpr/41BSZTT4u8K
m2T82G2JG3/bMJqGADAIBEXrwRVxnQcfEo18wQtmPiZBa6+ghuCRFGI8g+jqz5x2/gji4SdiVt/I
PKAUJyV3kY58KyQevmq8ojDd3nmXJAL6548xue9IuFqGgxn7WbI//Vzem6e72X3m1BS5MA/JsWUh
KQdcgUcuevKqAIyVMhSZ+MlRd6/qPYlA/KfYSqsTStfw2hZYetrWZFrmfXjFyWBU2s5SdrToNe1+
tyETd4hirKXti2BMlObnouFfpJT9c2LvjDQFNI0q0SHlcOJBPBdHf89iRvD3MbpTsblzRrxLcgTO
QCERwxSMAZsf3U4mo3p2H/FYxQY0FuDLlIv6NaeAGleLJtQVuyL8F8+UPe0aXZhfoED76wF3RUlW
7Zru+jyZ0BwBv8OwWCbFJ/1QUCcyGUcht1VY/Nggjih91w5Dcn9BBga7BBKxKpF2OLtv4cy0ll9E
YbAgv8ZTS1mWf8tP/+EJx/eftnOKDj+8v+8SRLzgUp2e+mol+BBakgdtSYGIjmg0m4RH0q3GxWTs
/0diMrfK9YwTq4oht1OLxu95+hjuqdg9FVYmDumLkL9MZL2SaIF8Em1U0MFiocPdLmqsUguDPP7Z
r+hevXgI7EYPWzotCWVnyCAdGywRp+VHK0I6Xte6V17IslRXOD3fn6BTBFknIaJvRp/nE492HY9Q
FlH82zOQNNxqZbh/XOSoghkMjc7DPu9/zATRG38Wz4HiAYTKxhITIKY2VZCWHEWbBaB5jbCodIB5
LkKgI75mVkkS6lQlAo2VNdCkYPBsMxe4B14Wiw45t6RMdrD43eoaYL4DabJTMPQpwNB6lVF3LvlK
QP23Zx9MPfvcKXCarJDZe6Qt0daa1Wi3TQ8fPShKVzSl8DuSocYgf1IuM/nNaSqU1NQC1egs/ihQ
EAoKJ2DAt5jgyxqqb8FC/QnANfn63WxU+O5DxwkQ1CUZ1YFIzsfmLw4B0I0MaScPiTCY9BZqA5FD
fNJRv7OeH6OJfoanzSGOBzsCcVfzC3893Jq3iclx4Vb9vQSFby7MiAjPcN88FZ+W4RZUktvLoFlq
0sdvWzLuLnjqSGNAtil8dT0Hh9skt+1QhshcKBR2HCHjLc46BBfvOGIgmRq6wMumGm9NTzPlwc0j
IPFfIMqBvhuAB39z+zO+QWIkJafKnd3VEkBdWDLySogCSiJsEJG7D4zhIUpZ8B1mHE5oY+0X0TYW
dDa1vFKBD2CZQz/ZlQ7j7gX3FRoJYuyaFBIjauHVRtBzl7IDXI3pBNoZngCweronetgBeFAbPY4W
UT4pAQP25Z+Zn8IYMpPquvi2USHWNK0UzqBRQcWqtunJRlvMkAdfDr6Axmmjpt/T7FAfds+9BMst
UWnQFBJE6UAGZgSMfsiRbV9K4r8QKQDPcOa2yapV0hKdMUJCM+dLPieBKAeDrIv6H7N43K0AjOfJ
rG/kV+5HuGASNFTuHNjfiZyDII8eOJ0ez4BGADEeQdc1klNMGsnIHgYEj5D/TnWLAm5IP4OqYgig
Hp0ZB6kMa7PxoqlO56RiN0ybthheVmv6pcegUxbOpI+kY5WHWGZMw8nkAkWNzdGHoAKC6pwNHCwb
j1LHbaREpNEuP6jsURW+4BzS4t1b+iVmq4UCQJFH/LTw4wDWHaPNE78lNXkMfyAs2Vh94ooAx7Ch
kI/ccKy3fCgME3Om5PrbaaRxZVABTbEPMppoZskwGuuoEUcP33NCNxNXVJPuDdWiOqkMzRX4h1Cr
oLN56QkN7qfkb6x4+E5+nLb7kgx8QlbVGVavzVmVbcpdSM0cge3tIBGTPRr3zeq3wlR2m4g21g2I
Rn++MLm72bYqm+D/D6scrTSsstv5lbUANndo0SsC/jtEmCmmxZdclv9+oOzp4gGLmbYY4TdblECx
Adv4Br1Tf+6Kq7VEEt4ZjOWuQ36cgozpnrblrAJLVqw0oqlytRUme43CsikFy7rnyPTP89iBeTeP
PsRScbZdixTYYbLsa9auUNyd2L0O1GJCppYUD63qrX+kQBgHsX69e8P2niGmGceCTN9j3bnLjpiz
sJdqR3pFnyFuoY3Q07Eh0QZ5MVHOhbQ8sOwu2gNot8YiREHacNtvSv/715HdOI1QE4Aa46SaI2fY
ZD6bxz5CWq/ehYKvQZhRXppUVToO4hhuTQ6wuD62UICZ9BAlNWID32ppJyS+xEYdAnQtqG8PZT//
Gm/n/SeCGg2drvi/OmrTGGRZikOD9kw2IdxUwHtuiK/9tv/8+lHZKUsNp66ctbYv6BNqoia4Uz2L
E0XfTRm8fsE6ezz9NulUCCUqe/3WN+BmpJlBWdaxZyH+Ew9uattIwh9AgFOdLbWKRLI3mp+y1Zy+
yNxLeXN9vaMT+wbpJsWi6Cd/EHrvr8ktx3kIGIKXivt4nKGPRtVgTzpoSaj/ZB7yUdhK/2YADtRt
XECWQHBY1s5ZIeKW0XdhlNfUKhd3EpnGZDgDvhScoXZ6+3MfNF8als+SVuQ5ik7ulppn7L3W2Vhp
ebGKQvIUNotlaR3hEl8J6riCI0KY3lI8B+UXnGaWWBOK4dm/+aJ+az76WSSBp3Em1HVH0uCExB69
8vv4sB/ri5ORGTOJWzyh7iiEM+gjxr4jrh8z9zt70zrkIj6ncJY0nSxxeVlGWbDB6fdyqKd5QpOm
gLSPK9zfiLe5wdpArJs/LXuFUmhW7jAhyWrDg8f/5L+6YVeMYnXPTT0+Y/3PfYpTMz7cdCrWlL9f
vUqwqQePGMA4ABRu4E62E/Md5T+whanqwd/2Tg6HiP9DmNlkLpWxAFaGDwzclZM8Mm/AObMiwZuS
pQg8COFHyJVjQfuex4PJFIq+4hQeY0GX27r+o0ozPrwxN1E/52b6mHaG4nIButjVeHl+wkqSqFQn
z+Ec94U1Zf0wls8jX+knEeo00yP+gc87nHiI/A/Aj4JnWSg4aCcCXuSYYFQ7cL+WU5YnCZteWDXq
MnRUpbppfEXBnP7ncn9qVUN5amHM2sw8Pa3IXjhdP2cNgpB1fYPZFBiwy0Y+RTKhlSAUJVfpdF11
2YoxhQu3YmVlvivDo7Bh03DUQPjxpAi4SSsIaX3UBtlDS1izpF/6FMkPb1pNxt6dWc9VPOi+5svl
MJjQhBVMuPdbJ3Dw8XtU3XRhqstuLrHiLMx0a4673WtCXrGIkSVh9+6XTAMJx8WZbaESKRNbEH9P
iZKo4Rpp+0rqKlNMgQwOepZJ2+yYm0XB+P/01mPQtkpDVm7x5Hq8R3naojgF9+h/JC+BJL9flv5G
JKLoz2M7v6ynjIRUCxgJl4XosZQmyRtuM5fcsr2S/NU2Oyp6/hImceaefjYWUP9UBJZN9CyRxoif
JvDpRgKv2QOsdFguN5Yr4FWzfrAVab4Qs55Q147vap/kMd5eS62nduO4uRWgRZDqMcOzvcstqZU7
+yGZDXjTRb8ysyVgN2quoFUfEpB6LwMfExTmWK8gQB7WZlEQxAVZ40ytMIx6rTDmHmL5jkZj22SQ
q0ZGAlDlPAnpaMUoTWNgPdf5LqDDnCqLbSVnq2wYgQ5DwQ87r/7r5lAEQxz8OMQ3kg4MNEY1Bm0n
UTkEAgGCr22msdfeqfDy0f9Gws8GGwLekOoc49mLI+5Q/yC7woSY7lSYFF1Z0FfkXLiEQjT+Y/G9
kl94VTjFHmRIAPOB0GoktdNEYlZvxdvoEz0lgMLdqUI65jT81pUAgJwF0qoo02VTR9U+8ERmpoDh
/u5zwDZzebnmroQurhM+U+SxibuP0SidizZ6h/ChS0UNzzJcRCqT6aLF7EK4Wyx/2uIFsmxQdvnR
NbNiqmJaXyzDwtjKNzPfAA70iqTiohMPgnXDAdt2UDXJrka3ZVGbmZnqW0wHo6oL+XKoYvOM5R82
pVBJEPYKtCDNf610b/Kwu63iKA2jgNfwKZDri8ULgK2czGBxiObLiBkXcLIlzR3ltG6/1nCbQvzq
vwZJHxERsp5D5BbmjoLbL4EScMRmoQW9zu1zrPINjAQwGsHp51L2PJlDjVzT6Ip4UNOhYFGuEWpG
jtIAOHM2ezuRmLsYrSB8nprfaHUkKDbtvr6WXMoFCy/Ri/h8I8EzZXbSMV7uCADHGQaPyYJWSyiH
PfCa9001x/X4PkPDgJFEol6cOyO1D4JzHH7Qzpg7ZRy1MZzL4d53F/FcNRKU2VvpA6oAvVAPqCut
YBX9WqwTJjdS3SxygHk4bJSpiLUsNyoz6qtJYKBV27rA+EcMXN9WHuGDQYX9qI37Ru76nPcVfkYy
eJakUJnQ5BeQttIbCKV4DWfkl+ysJnIzXCVfNLW8Pqp4/nAv1stxgjvU8699qnm8G9ULV6xtEHPj
X5AaGAHbrm2zL2uzRlNqC0AMjq13g4iPk0KGLAQ7qvqythQbyDomEOTvvH3R8nCqU7GTGwmdiRyA
dxg6uR/mOgp5i9msPNb1zUtV/h2t5ZUIpy168guDg5BQEH+b7EX0BmqVzzQROkJ/scRrSy6s/IFa
/23sIcnBlKrRdi8QriImH0Qw+b1beo9UcJBhZqADlObouxZqGghyyO/uFg2u6aFWHoJYvVlDWARh
j+FzPuooPBJlW1qagpZ+drB1niPtK9SDgovBcW7N3VfcB+sfwzvbKbQ2XU5fALHRhDAvJfGMdRUc
xKv0HHuOyRZg/Va0T4XE68n+cegRu59KXEOwAA5NSmCnfvPfxRe4TLRqCC2LhhF5LX1NQKbhi0Dp
HYNKfCx+ozAgPUCLMiPD0o8MjxSotQ0lx1kLSSwtr2d8lgKv/jxFlkViQJwLnF/RK5PbOz45WmYU
zRLY3q4ntbvWhBeZFXcnH6ZaSIGn3x+WHmeBzfgZDLBOkW0pzidnEV6h+f//GNOF16VSb7mvnMzG
jmx9Wv7GTEB9SGD/DSMphzrUVDcOONCLkZ1egX1k/PF0ygTQbDDORhBkln2YVM2Tsohtz0o00iy5
WNoKBhMF/yyjaYg6YzjseLMBPw4KbeXZ3nHZ+k+7omzRcUdEc8h3DJNeTSe3fbkK/mQ4xuHFF42i
hJIgyBkX12pftcy8P8XMdfNTnIFHffnqBFt18jKzKBqvfjy75d4Gr51qpCvb/xfYjTpE8SQrSk46
ao6nqxWmY3eQ9mcZmZmYnGkQowFSlIV1f7Ctbp91X3MFwp0lulIihBSNPrCQekn6PeF+SpUoEhRy
2y3Da5tbIuGsGDgdA8G3oI/azku4RbhTKLy4ygYgmq2Kiqu6Nl1x728meTKfh+/Gp+LOekOmgJBb
9hOcfFhq6pBVQ2z4F6+CgHyktq9nN5We/QJY9WJQvOTSPnDL5cYoE+GxuGRiO8WPJbac/481MSY1
s4aFaUH6xChooRlAx/+4XIrnR8iVO/P9ekt4xFOB5t81RDtvp+tzB2LLdW7QloADJCQl40JK2GRN
aWNBJmRayhY3MKCooNW5Txmz0QbxYn20rmPK5q4r069wMH9W9ZDM/fzU8et37RFcEm1tST5NSiA/
gez3d5cG3QjJdIjZhlJKSfmqAHo9U/EaOdJLoNqSkv18ohlv9PonzOlg8NRErCiqWWQWnsEp1oD2
CqgY8gIn0IJ2/Dul2ohH1EA8xbqiA4KyRsBQhOp7474rFQMhR3wXyzJNKxNtId9tuYLqb+OfN/GN
QLSCiZ/XzKJEFjtn68xMv5XnhJSK8SAfEcmfRN9nyqkKHckXQa4nzB9nqmLb8abVoy85+209y4aX
I57B9NP5h8rTmzDgCk/DwFU2B/dFWlDM7yszIsAJr1vL29Ei/m+7CK53T3WkO3Z+Ozl2nnM2p0To
tNISaxfb26A/vWJi+BCHWzUmZ3nZd51hsufHwtDW4r3/A2VTHXSTA2urikj0bmBGsyU+Dx8o5NsO
HUPMkLmBAshqyzAtHLC2+BPhsTVc8ZL1fE+7qk9x4iV0/GMsI6C3RvYROwBV+aJ71CxD+zLOdRsc
C97EJ00CL27dZ8S+lhlwP2qRyqqitD4byhJEglQCvVk44cN4G/cHca0pZc/GxK4P2tSD/yxllTMD
VQh8X5uLiFejHTrMhhSnWIYq+cwYEsuTV63cEPf0vDa5YliMvH6PSbR4cMxCKyo1saP59dfbeqP2
Jx6yK4sbaX3LfUbJNwnbyiYXTKmUU6xwpZXbcqklIcgGt/aMhDN6nfPZEv6O6UhPe7xLhOKVSsQR
bGa/4n8nhIODin+9QvdcHSOw9hSVwlDOVL+AUDuhM+RBJF71Crrenygs4JSjnsByXTKMxR/3XY3i
RBkAIa4mmsTLp9SuzIgwbX5N0QBtljx482XqvdXlGUOdZnRQs0dQN365ZurmdZkZfXVd9ONxlAvX
gM2nGHGRfRM5XOM/4DTvM7DYl5xm6HFpFCisg8RHpIF8inIEK9yQNa4MnbElNZYvKh1VabFM9YQ5
kptOskHdwkKWp0ivqgQ6FkMMMlUgdQrw3eFLIII3NIivSA8PnxtIyuSsIiATLHQYHVrLAGcYTuKF
vpeCeV9U/H3k/1nDXOglb//sWJ5ycfUGQmAJvEBWO3GX5yxh0RVwtfMJhguYGZWBmGVq3KFZVJDZ
l37nZNGlwGdOPdAVYbRTEhBEsaS/c7kNl7l8X74QJcCRRnm5d3n98mwoUq5sc5JHnS+fFmyBx2pu
I8ejroFF7JpYyjCwOu77vkRKO9VA03wUYLdgnBwWNwwAhjprynFxL4uZ6PJWHbsD62lsfKUH0pcT
JiuqnBL9s3X3XnnmANf7gWFesUvh+MzKcrUeVf8MUq2GBBJDWaXqJWFwxiuyrVEcD8IPOhClZBzr
hgc9idhc47/qxyxsG4XSwlArGM7UE6F+xPc2vCjPlyD+s0k/BDvE7grJHe390ju69pLKwD9c8nOG
Iu+HW+lDZg5ae9sB/iAX2fohIApXuj+/j9l6tJwGENhpIF6/0sL4yMY0SGZClEr5h2iI/ys7p0iw
4+tyadblK5qmQiCcxlFWcPsLM+1LqMdQf/bHXG2s2+2pGp+JgVzwOXAbbcuo5ij4K/9fOe18uSHO
/lt5AHtOksxaLKBLDHZwm0ZCHvvaTG911NECFxshws/KAj1PtHkBw5mvj812udtihziHnqVoaOik
oB6vvSJsA94HBDqAGQab001FLf8FgxobgqiiehKJU+LNLtqtvfgDl8a7CyTiKThgDVDq3hbDqcpw
KfeyMRReMXB5sxud7/t11Y4gx24cFIj/HOiEx6EJmdUVLjVXFTqa/hXAU9syG+NH3d3wp9J3iXNe
zi0chvO03dVigdPWE//fIRDNd36+Eknt8wQAHCgSG1fUQ4vXK8SpWCfHUfoICbn2wHW6+atuGxwz
mZEQXfin0+fmCBmRxTWzHucXODETYcYu+jU5+H8KrqLGFl3Jw3eu8iwsMlh3oJlwYWzi9LnIv7aK
Ch2OGE/ltlSfGrai8N3G5AOOM/p6wJEiMd26YEy2zGS2xqaDMDS+qoldTUoc7HFJVrItsdcEUlGv
FOBa4RsGYCaZq8CAY+Uh8QFO4IhAlvQYbmaw5hUlv559zXxCNyu16QfKojGudKoSE9c5Z2HwDCQN
EUfW2+tHFFHe8W1palTkCjILkdvRzyANF68bR9wqtE+qII3ETou08bLUcUZQAAwaMz+SEI+j+pm2
g9EeW9qklLAtLvSvGkkcEuvH7GYPD4kIevDUA/kv6cG+hfp+xu518AYOQvxQZjPcqsHD6xxq57JR
ak9hhXrc/kACnDaZhAKJqdegPruTjsVcKIIS6IGZMeNe05PcRSJxR1LUxAbpMpEG12K7koKfmp8Y
+wGXiqVvY+BL7TeDKbRtpDsGmWGckbaf1dQjO4UrYK1Rh+TL3jp/irsG78sRfH1CNYtlvoRtOgrB
eFJaO1vJJ0wHTzQ+0FdXrMrguIXLeUZV1LbrfJqivvz+6G71ip0zo793AD4KJeb6E5LC97BeQArs
T3NDAZHwbnpUJSopJjQPuJWQLjHDZokLm1NbLM/ofQFRKRpuS/++W/0qybFMGDo+e0rO/CYGv0Kd
KJpcyiA8BSa0G8QjHTZoaG0MAhEURaOhCNZryaReNXNRjgmvilaOknKBs60pqjZeQ2+eqlub40Fr
MSL2vCMKgKtTWKQ81Vpr+WpKTYx+D7Bq2yeGKyRLtvASHSQ3aAMRajeYgh4c8a0vycV5EIIyOgPo
TlPKrz8GsqXvZY3mq2rViKmS5Aoe6fHWii45mvNBN2lBXNfgc8IlyURkas3UOmAbnff9qWigFLaL
IupWfHBk8JCr60AcKKg6l4zDttNMKL0+aUPixOalZO7IS7kYt27zu9XUlJp4isOdYG2oJAZACKiv
aqH4aL5Z6WLIRyjLRX+9ildw0QIcRV6ZfJc99rmq+JaWoKmmhdHC7NwVXJNGG4C5xCLtcqPCW3oT
OIy9Yxe3zp5qTMK/9EFGmT6B9RgKqSKUX0pvX3yw5fS2SsyDXwCOdSESagk5ISRL9fm4/LZthvGJ
0LNEC9HYGFkGyEPrBWOYDIird2+ESzBsGKLu+2w5DvK8qypYRw7dFYH4kgFEmjQ9K5s+HTwzp+fK
0OW5RhNUnTeiVJJj4ZLthNuQ8pe+NEjQq8xK7eU+PRW/WFqXwZFx3/z2JgWu/kkrLUly1J+kAVHe
dV/JIDa9pTVV5k7p93W1ftBQ+uPXDV5nEPM0cVcKZyXeQSknJqDf2+MAsUpQoMT9TJLRnjSj65cj
mJzBn9E4owfPl2biHTI1jMHuR1S1I4xDBX2kM7w0C4g778ZzDhk21DYDxORyTyLyKg2B9Y9sZTUQ
ULsOWjk07Lic5EGaqqP/GCGC83uGWczD6hapn70CiNcsyOUgbBUNuDfxpQwqIi6EDGFs+u1wOgtE
RLt/gQ6ORGkoSMsxJRUxRdRbqrU0oILOw6YCJ/CIx50jzgUqnE1HGlVdQmh7Hq3XIGkYhrK8r/74
PM6fzYYS5pTL5dFERuTNonaRn+EAiUGOHL9jZws3b+fxfLEBIXt4z5stHwuS5nzUm+A5NnMNbCKY
5gRhHj9DKd7upZqjBycdDo8cjlm1rpULSRGtrm2YbfzBOLS6xrMLsgiYZBY/l+aSyiDQxmjKRtBL
yqTGe7BGWtPZaeVRblm+ZOfqecfk9ArLgGVwc812b98IFjjHhUrhgRH1HdHYhFJJ21kXMWNS1wjD
6xt/+8qLqnP0sbNOiPU0A6uOjVTdzHz71WFLVzVtdNqzkhOfoiLgv+Iwm2cXx14+XW08VlWOCstQ
4OxA8fdytcMt7T2Uhb3+P9HiSAqntFPOg6S//8vKWum3UAVkVoZoZi05IhRs6OgXZFN+zB4nWRze
zzwesZiRH0ZRaQLK7adqLpV8irAnmrQZux5W1jlV9e+cwPkhMFI+zFbPqepBwqFLjl3nPlaYChic
hkXGYT7xLXmVo9D0V/LIreREl+TIWOa3Na0Ryu1xhBEWqzPHIfr++PhRL3KkfApz8NDNdRK3f+Jx
bK8qU8P81NUwghv3Cxrd+TNBqCauRyGLHvNhJi4dE2OF0y31bK3HdcjMLyUrpROdJ1LAtqycjZse
19LAlCmzyW56gZgFJUBuasD6vIavVvfrlceR+AtW77ldPFvzGBkV9kWvKx5EaaJiX4TnHp3Hl5wT
PRIoAgGfJ2zA9GoKd1WGnl4O7AVvJmKX8WQaxwcRv6cfG7dRQSirBF+x1wM/GaNAagvm6OGQaeFS
CjKAjeMmktb/L8zrOi1oszp/+pMX+3AKc3toRc1+lAxPZXAG0hV2nsG12FL33YoVsUs6/guGidl4
3DzIADlKoQTUAGjPPwkzAj2nHcBM3gg1ogAJbVvZyeplc94ViAoHqmH8uIpCLUNlu8xkAMvL2wYL
r8TsgyCe+rK6lJys3H+xHhKAT6NeJyewr8sF0j3jwSWS/kP6Gmf+wk1/SdJgPM/HL6SjNnCjb3MK
r9Cfz01voxPL8uERl/wt+ZaahgfeLL62SUocTYw9/t6I6PV+9ijC8rdfknCZSgA4iiUOEsCIUzf4
G8IhEzH+CchR0xmjTsExzTf8AEOXOKbVWVUY/VU4ZrW2ZlOfSxu1yU5YDL9oJSqQ4twqixmWiUpk
l8CCg25AZxGg8aA9MPD7q/l7ZIosaxXdDfm57tzOt3H4CxRi5ZfNDtQmyR54hIjJ//VKFawDc/eH
SVFvtjfMysfPopHCsW0katJXS5FapZNZce+zIl993H4XiNG+u1PwJw02tMJBCJf6q5yXZCbo5d46
KuLKmzjXGKegI2jPjT3wDejAPnLInk20aouyWi8ZfgSfiyRftKFRcO+XP8GUPuaw9PdoxNy0Kivz
qDZPspPkmoR1qsYdcYQZOtJn9OQDu03bJtKCF8yCdVjvYbVpVnPY+71jW22iShs+MmAPBdEbfFLZ
eHXUThuEm1sNo2DnyLElnGiZTp2pL+NYwIandMuzflfUSE0xiQLi0+/HrzBrUILDdYhS5BW7IzI0
TmgYeeJPp8EIRBECk8UU5y0PPs2HxowWTHvNHY1A75Ecdhaciwj13QUSgLidPljCIyB0AW0zSIvZ
k9iv723YcL/U47RHAZK6Fh6SMnclWMeJO8r4Gu583WO6db8lYI3OzfxMZlHXWEuPUxJ20Bvy+6Zn
UVXnjW3aWqcZg5wu2L1FB3QY77G+hUrWQKyWSpSungHwga5GL35ItYNPVSaQYqaT/O08zQGZR0RE
UUiaM/kpH5MbNTRPWSJmDsAKQrPoMnYiH86tF4bQQ4xgZnaPNcevnR0NsGDg+sZXp6B2StwIb8UU
iV1TW4PwyoN2QZCQyA46umV2oNRVuUA6T/k1Uqskkgg7PPNr/3tfKWYbXyEoRQ7PgEgthG4YnsDu
zE/Jq18xFSTALtoiGAwoG95SrStTkWvbB2+0DTD/MyLIIJOLhExQGP5MPKkHaNhPzY28mGvCOH/F
1/eUmWcvgXwGq8DbL+SSrUsygNyeMqedCApqDqRxWpfapBoJ3qGK38I9OA+ctU4WhXxdvmXzj+8C
Y/EPrd8KV55bCiD8s5+kdw0+q8fuuV/fouZA/Y1ayzWJvJGZ5vdNw3+zklpxOf/s9AcLXfyT5AeQ
G+vL62LmZ1mE/hn7qY0wgASr55qjlPpBFTMoUML0MKwxs2oyrWqbcDhKN0s1OqRCGWAg++J5s5LR
jV+p4CfJVV7XSW5sgwiGclboGwmnS/NcZv8gifsd6YQToQnqteP4NhdPvcorbVkmuEvl0JPGw7Ec
fcJUmEDrFheAOh8UjOEyf8WnXVxXz9JuIvtSbeOx9pLTIiNPjqVTEzUl9NyPGuKBD+ZtPFAYcU8M
tylsf4HPydcZGme+VgNhsaImbGfAp7EfwHeEUBbnqZLaCP/1j7wMq7ryR/Nhu2lhFqO9l+K6EIfH
Kphw41w2kcZWmk9KPe2NjYK8qv+INTixCtCPO3iy7Gjxgy9C3S1w9y22I3yNv6R/OULjYEE/j8hw
/aZZfeIiVE1hyYtX0g6ai6Qv8crIgfHGJIyI/zptER5GwV4LnM8D6KqOY+Nv19asHw1CwRWbJOwJ
w8z0ZTt1y4L5cyVHQjME1iteavLxz+bnUJN0DJwCiGIq2AU1AhhL8d0aP4x4fQi0lZgUcake01Pp
6ryrSG+hXdOMj9CvA7L+QeXzmjpAU76ImtUh03yKoW1hlZUcxcHi7vmA183z7gnQd/XoUZd6o5OP
3QCpnyGH+g6xOlG0ewRvW9sBZ5d4lFMYSOLCeEhhI/yQJ0XrrpI+d5y0X31BIMx6MVov5OB0KIsu
e60Kg4Hl1jvgIH0GGL7EE+mR7TqlaWx6Y2U2jv+IYKlW6z3nA9OAlXr7ol3qbPY8EQaF3XUYnVLu
003+4VAwvwVGIBRIes1i7xSK0r0OSjANe8PiYKuqjccJ4jwa2BVKQrQEZJ+3hNdh7JmFd5UQgbip
o+8g1bBiJZVN9Bm96IEibqsdkGgtMyfk5Az55pvF85tj6/n1u8CnUY8IK1l17kFhj+E1OxUS564U
epi1gI197gKmUQmLC80n8nUBRX7OADTUGLcGxBaUMRUW1AtJOxXwhDCqrxDfYvKPtdFip7ZZ+y9H
PHYzXPgPdtUxeSTQeLsIrkgJUHDkjzCWXOhpBcVJici0i8q/ej9On86MmiG3N3/34aVuDLoGQCar
jqAK/UyxhG7D8GsEKAi4RjnlnzP+sPA+Rb1FgOzOI0KlbWtWPWJ3Kv6tYvaKAfTynlaLMjna+VZm
C0gMHWuH85GrD/jbQLv6CojZGWXe/5inkirPyHLbECB2CTVGwm9hf3FrXHwQXPvM9LQxtLbYSUse
fQOoZtX+6zAp9d6VJuKvyrQr6NF2J942wBM5LTxou453UbFigg46SQCNHXg0XLZ5Imd4H1NBX5XC
L9yWKkJKwZ0ekM1Aac3amgxNR1U6F1cvnF3V5eyf1eClsRH50jkg79cGrndYNpnaMscDjSDK9Cl4
Poc8nw07i0V05PyPhE2OXYg3CZ0gm6c2yVCZwlphci/jNf7G83c72h/4zKK1vU1tMJ/3WeoIb1+u
7FffWRyXiob6EOqUTFUy3lOpuTB5Qf0yoYZcLHrtV+yRsD6E1WJE2u6xxYc/jgeB8zpH5wlTvHn4
uAqN0rs8qEpjwt9Xo5c08XsP5Y7XTm3z4LWmaCj1jQ/XXF4bKBu34GcVw4pL0ah96SSv/lC0njCQ
RPuv+nOrdyGwKpH96zllhFR2ps7cTOZsUMNrtEl+4GAs814cIVvbE6kFTzQVgtH3LziAS5bLmB/b
rdNOpODWWug6wzM22zrtS5esgh/qN8wjwACm8CAOJrjaEBlboeGFAx3ZfeIK4hNhMSvQqU74BkZL
sWDTRqqpPLNwW19ZIjNJny2HogNuOXF+HpDHzJPKSpjuQEw/ldaASusGcMdVqxbWmJAsA70L+vS+
8ytr998E7MItikL0pBVvrE82TvsIlCrL/GCIQDtC2v1rGfLAcJjNS4pBU7bG5LtMXiqO/1bGDfpt
jstRkMwQEQ8MgI+kr8cDeNp6H5W/wVrjNAtVMlUCLxfn6I7dumg4EJTzSU+NoqNOZXU18s80hIo7
JMNZ/+4PYMA7CUB9HQMi3FlTIR6LN8ocJ9IjrU66xt0GV5j7+7gu84RezhE229Ew1sb4fx6jsKhz
h6lPsCG1RVIy/aDMESBrhAnXXifAj3eAPrBE2SzR+IJYGXiAwPolgU6HwJhbyHLDCGqzGuqfRaz5
5jg5Zn6LJuvuscFPqZUgpkc3F66WHo2KQRMiKId8MSTsg0dD90A3j6kDk006bjr/5dEGrx7SWxhD
REh2fjWcZLrRJx6hDJAlFp6z5+Ps1K8x/Vn45W1mN+NO9XOfbxulhuwCzhoT3fQtz2wgiccymMNl
jS/+Ryl+iC7trwcVMnzZU60OiZHjmSTjyYeeDnJZ7U2Q6R4wZX24dnKT3GwHH9U+Y3pNtmcLruat
X3UmxtkXmTHZVVp1Znjap3p3b9sTWLyWzxuOmlJyxsfDuaPsCkcnwyKocKD/1S3Mdr7dSRZmUkT5
ets+hgqZxh4JuYMegRXE47RW54lHnHwiQ4U9fyZalFjmE0blUuVxmwY+QeXdIVmSpm9VPaxY41Vj
3Lfi8EiW618syVYdY/ZdiKK83WIVsZwN+vgAySPvmhizIjd+fWfk38jjcZYB7mIF43f0flQT8ZP1
Xa/oEgfRyCYRKgNN/figar5J8tonPnaOXNgislisplIQTxn1nPJ6SKqRmZd+i3FvrcpGppBuopUN
jlSUMVXjs1m1VeBtdE33lbGmY61lIauLrpey/yyMXwkqk8aWps4XyMOKbpS9dUWtb+U9T0Z3LRKv
Jj8F2a474PNhcaDfB3pn4Ob4FdXJstRbl8Wq8AZE1KxVZWHRx06i1aY9Ky+WwjXwOsx1AepYT7EG
gILuLO3sYuC/vdtPEov5UUVUkwlpnmG2lfu7eKZ+meV0KzzuCwz5g5CjjmZ2UUR74ySrp9KQkk88
rF63zm4S8Xkap3h9l0/YdYy7rM+kLC4ixAgrtXGJIEWxU9IetHZcPCZTc5q9fir/4oj4bqjTRDkz
ccWsbi5patCF5llvfYrFRSGmox8Z6IVlP6BNWDy5Mn0pgUP1QbqiwXjNYBnGdYkdJCqsnt/Zp5xk
jelLhhkpkka/C2PCdbMvpaZIysTy4w++VJ9BCaQHW1XckopZdfVVmYFTXESzT2HBsR9ejpCCXnpB
0ZR4pwXbDKs5yn7X/MiXRwXUzKMI/Wg8JPUm9w01qAbl8/YtnJpGSRZxrsmjbOmXuKEWoTZokcrr
ZREBfDFGX1AdM+hApd76/jsTnQDkdS9ql0i5jOZKWz40fu7EPQMkZ8QqotKc0mOzq5XJHNLwdWhz
DEp6aD79fCeVPdhnvE/Bzs0IyYr0ExTbMnIjXptwoRmB2YtkZoVZFcfohwOH0FxyBu5avwtI4xWX
vmNOz8qv+JFwtBZbqz7R2xQXB9shLsML0gR2qeZpSyBvVlWaCA8rl+Bweh51c70ynLZsJ7sDWA7i
qaDBIOD93bM9ea3K7zfgdjm4yZSFdWleF8QJrwyTwnejEALqs4JA7Gps6KR/VsQQKWKy7/lJWXwZ
Lb6Pm2T1xWZkzxINFbaKHGvymhPDYi0BFwyYI+iNq8v+66PMX1uKee3j8ZMJ/Wd+U+X1F02Mtwb3
Okw9plUzpm3kBVbbGsa22KcIQ2hLaBp/WWSfIZ2VMkUxvvU4nioRe5mE/FQ042/DmIMyr7mvEj4B
KMMgiPOwdlT9chTtRTd5PN9Pnx2F4b/AZ3igGitFq+Q999X9ppiJkICHMcb3cS+o670CEIVuNaC7
ndPjrP/539TXjoNAV88q7vB96IrP0MKgdwOIYP33dgIaaJVsSfXTXZW1TJo4GCi052VmGgwyMM/+
YfVtB86DO/mq68d63BRhb4/PI1UoSqrgupbNN2HnCqTwmgMIXAVIpWK+Fy+6P365BZScArNtA9xu
83YX0XUtodzFYOcH387w/FDf7wY0MMpuA80+23mVJkffj1XpwBSnrQWxB34k5uEzk2aE2hVFiO9D
puggRoiMXXC+lqqUURPx2FcTImEdiQFaipxEsFNBh9+eCJo413i7pteRM8dKJdte/1dzcWbi+CZO
jZfIniETRt3LrqhugT6mNc69/6v3hAq/zdleMz0W8BLMxh+arslFagBawIIrJWwflyy6TeTZVw/n
MU6uGPep7KBnC6lT6JYPjz5fjsqc4ShBVO4uLVX+uxzekaQp6b0xyG9IytRSlOX2wINOn31vHRJs
CTg2xc2G43ZMj7ZTcys1eBxoXVqTp2SiZlr539NyZwu9yHmqucmmCBvVhE9YP2JX3XYFq2hJ7OfS
auRTGkEgfov8BSK82Kxl+k/zRR5BHEM7ibrLDYBFmnlf529B1WwbF81xS/rolnwxmmPQ9/4I8AcZ
uxRjLKlF8bL4nof2rtTbFGhZhuZiUirYu2hIkYpqv/guQWaFI+DbuO5Ycbm0QlVBb0RINUEALhwm
angtXEV66+6ZxbF9WlwjK511czSy3ch/wjFCG2wpAhUFfqi4ktTM/RAGryySxCO0SAnkKH+FqbFG
KVzDtN0Ua0dSpgQCTwSDpoQ12QNXzP94lNEAXsJZi4beeyZcDcLhqvxPjJFJFWyHkRFYgvOU+YFD
ORnLuHwizkQSLNhiiAHV3PiUj3vu1bK9seLJTxh3bNqWOy5POcNKUVj/4ivejbTr24SXi494vB5O
TdXBE4OkGFbljVdOwKqz2bzjYyJicdL9DI2K0ZSi/X47350GTGzfXn1nAwcIWkZWP0dBDqglmuzc
k6IZkpN9IDynJwNHyAyUhkhd1dQerVNaiB0W5/Mzm1zjN3TGdPBmbWOFuZtFEvunBdjWalewnVsG
iA8oWtErGdt/n1OoXPcRKdEZlr9ufgDP+HNlIybFjGo1t0JhoXwZWQGtROaC2xmpUDpObX4y+/TU
exNyLG3qTjhZzASQjN+j3OU0p+dAMJdc/LIO+CNCtP9gqSnXLnxkE83xhOL5TwhPNSRpoehQ00PO
C2HozTHwHiHTzH/RHdPbzGdoiFzktbWY+4Gyufv/bIwqietkj8WgIj9gRqQlKJIMrY8rBLu6H2Pp
rGuu3IDZxoiDYcDs37lmfdP/cRRu64vS2zUoPzGIrLObNTKOX1ZQy5/XlEh8L6/Nc+0kDOKWIAEN
1Kt0z8QPbozgNXPgj7O6VpMXhXkXPvYagfL6nfldt+PvDxtG9YMfC1qSVW22TstIqtnW6kbOEIKu
EaCFhRzWp7sIY0sOkfVsC8Dvgwj1qDddWnUofN0NTIp41x/Xj5fF8z49XYOVwFHtqK7h/bzgtSoN
1yGb3QXpcBH2exoJVlNUH5IDSEqgo1+ZJ7rJh53chT91g9cnBBz2SnuzGGbHlu3kKH+u14ezqa6Q
k/cQcyXxLGHKzaUm6L8vY87fU25io57htARdhM5uPqjL9uGid33GNRbM8jInjKcBsG2veOJUFn1L
YT4n4dX80FgarsLOZ+2tllknLQIXjCpefWO+4zMLR0jJYFhvSvkFq4z4rFioCLmeM61HeyTiu4eh
RBJBitlOzyP9s5ilh8GFPYBVM7BVG8RcNml93ciGajURc67NDOyY0fJG5P+jUAI7HM+rQMU0NAsu
/l76aGHR92VcnEnC9zKduo6hGIiwdeBXZ05Bc0h1bmNROb+Q2cw7oxQODFX+rrky9dE0Ww5Sq3h7
S8Hxx7sA/BDpLmZSCPfakKdoiTnGnq22JZ/Buqqj+f6cY+xxDDRvhHKWNsxX8Y8C4CgCB9DTZB+k
oQXqzuZSHlbSy1tvcM06PBDtXXQWNVvQBj6CFRBaBu/KodlIMknvEcR1kCCk5QKcOEVUw6rLBxxr
/KZFQ3Qkyx9hKUjO66RQB2qYiqVUwwAkTgDsKqjqButKyHrlJoVsNAugYPXBlAClAJLvooUbssar
jKWfeRtoF+DIQvGKl/65+jOjHkbwcxWKGJMMJDGmCVCSOHBem5zQ9Gxy3y+gBbzuYh3SL8wqU7H9
Jj7PKDDqSHHApSBYdyiI3AwxJo9jD4RbrQMmIIl339CvdGIdv5QcoVSn8H5DxvqnO/LhoonCOAut
1v9YxHXTj/1wBnfiJtR8xA88aoTHUM5yfNpZJBhvKCVYXOrbn6pkBjJA+8BCAMwId2G/QHQ2yz6T
itMa+27FeFmpPLWN/P7hj99lDZRFVhSXjSKet3VpH2+xQ3jMbS894/55h0z9o2DbdkyTu4DKcIbt
ZVvxDo5raje1duILVPcDGv/CfoExHc2MMLu32lNWX6MAbWhxNufEEnitL5WdhgzTjRgKQwvNouIl
Os+PtSt6QWlF+4PWMEkoypWXqquXi89r29C+krJIYtZ1WeCIE/F4jt8lrdO8XP2odZ6E875tE7HP
o4R3mb67c8gRSL4+9R4eUcp1AlfGrWsu7o/q15iIvBwgXLRN5/O+D8spV/l/+cp9hzKtM0WCUMrL
yRRrJuSEoSVTiLj55HP7CaSZttQ47cKYhn5g/0XufJN6MzreeQf7bHltb20ItFQEXtARTUEqZpA/
/ZVHDpeKUoXNhL2bC3unVuEdLMsVsbAFV8EVnCUAHY2KneAUqBWjU1iTIYFBAXvlRGod8pGKgTpM
HUdyitiGyPQQG4S/jkoF3IK3qLD1kl3mJqcr9DxhznV6GJKgZE5Tf40ZVZSdU73dvqESnNHz/1P9
BbfOJSJ3ZpnM+5tF9bO0t530oRtUvO62hhTKx8XgeOYspEIvuO2VBRPOHJvNN4OnR63QBYFQZfiM
MIN/MxSb10NpzORRFLh+Z+Jn80XfJpM84VYKFWC96Jpx8HrBfCk4uqaZh5JLEFZPQT+f99Ex3pre
iWEfS8MR6V9IgFFo6j7Jl1b9VjF8pBUR/dB9frT1ILQPtJy7DeFHd34pMqls5gJrOO7NFoeHbfl8
LrQJdimakxSc8pqMMLf9MDn8CUYhJx7pQHrYxhUYUfV3oboNNLG2aJHt9+Q5N9grH6qt4eAYSOgm
MJQPzJLXu0T57dTMIpqYNhTnE6U9w9yvrnIYIsbfu4KNMD3bC0tGzfbnbYHlMWuvDroi6Fo1GJdq
R1IC8Qd/S44bOeRXGcN6UdCA0/hHPLoRU2coT/BxGGJ6lrrD/hzLutcRTOsigLiXZRAx1+Vk8haf
2qTmXWeoVT3bGU206KpLp+pd/7AH2X0RGFcLy5RrBEZpCCbVGVndJXFSVtbzfIbEcDYKbxFSXnrg
0QUJvUloeWCvRzgtRMh6XPF9qrTPwCLaMyMPLnE5b4/oPBSmhDkvLwa/A4a8dVgNpGv8CJWY3FoB
Khb6sDiOfMRMeF/ryNRt+TvWqjwDHPuQcuken8JS0KJVsc83cVSOGfOYSUT/rNwJ5ZkxJM87HS26
aNvXsUYpubaU5XFaFmgaFqQ4YFHHkoRWQuyuUmq87QQ/EncAUGJrkp4Pql5NdbyrVVspmekVPMzY
ILE4JJwIGCoFpBVGm5jjY59k1cw8AkSnRMzr9n6lgumI4rpOIAMBeiZbUDeQXXWtcnyZ9ghTKh9h
8qBcMIl09RXc4PluP6t0PNhaYW1H79Y19jNBbxaQrh+a9Fs4Gi5x/BmheB783aSA7pHZ94E8hpkn
SkSyhbJzXIlWtz0HurMjcLsDMzilS1WYnv3Qk468tmoE0i97evY6KV4bmVFCLubOcpSJOv1g46Pu
XvB5DPwK54+kjZqpkN5J3hkozoahDgj2jw2vDqYBzh8is5n6bUv4HinkWHcnISND9Q8Ow8OpC8+8
hcMHDEPrlTmh13Lf58usgo044O8crFRvDp1wG9GbJ08pACMGDgvW+KiaIivx3fGLvjRVr1Dpdz27
b4xdKQ4QG9JB0nQIFYc9Y9XsOULFKdF+R1OaZ8at6pGUtQ2UmgtIbj+t5JyNZRnDFxvujkrYm7yB
4bofIa+t1P1FAQ9mchL6QeeLGNtcz7qj9X2Xrw9dE3UO5zKY5TRhkFPDKo8GON8Ex5h0nR0Hu5GX
FiAwud0LMM2RE2t/OpN7iMZxstjIuPouk9mUrG5l6YY+9A6KY+XTUj/7Lxcx6OulS6gVhCfS/NMY
9cWFqRcG0+UItzmSs3RI2J63M9j0CQKB6vxJHFs63iftLAVUJg8zG0qxINyFaaghYvaPOUGx+d0G
sErXyGhd1JStxndmjmo1OV/HPnBScHdIPmAdT0IfwkKUGxyf0EMIYG9jgcPJufYWx2k1W0+X562X
bOz2CcOGJr78vXUgjdlc+GS7lMBbJ2LZAdb6HkdqsPl0VZik5kuuqSUts2yUCBx0+Ju0jd9k2hnn
B4nH7Mv5abIMHG4+DPzanNO73q0YTFMjviU7uwu0SXA/+fTNDsIq8HvFI4jCHDARwDVtEErSMVbT
G9+Za6cK+GsD7j/ENRzYzOLvitPqArBS3lW8zEFYm2H2CfzA2E0rxMD72AsJOPUpJldgP4G4VvqU
C99g8CGyZHHg1EO7vb/GSDxZvqZu9pkM6yL641+OA++Y7elVluY5feFmuL9gEDPew37OkIDY7Jr0
vagaFLKpJd2KAQcRFNWMfFFj6najgNjGAvslQFsOoWh95mLWTvxLbbrwJMqEaJ7M8VlVehaTaeF8
T9DMbBb7ouXRP9jrfD1s5J+xxMxkqj8YuPUFHP/OirFG+rnyn/qZsVt6SL4mIKwiVIw9QudC6+CK
/S4MDUfDufYCSJKUyD4ron+g2vwYb1qbK2+tRdKKu+Bm6M9uTpW7F9B1vM/j5a0FjWnte+furnFO
ZSbZWoIeJAQq32yEnC15AgOZQM/Ygtqcb+/quo5IVgbOwkw+8SRtgBmNfzbZ349SvZ7skK+KoyQw
wkyaTsJChSIiz5007bOwRz2mvji/l2rngAlpGvlmhqe8zlNcHYZ5fyVPkNPfsYeYqeKhMnATBeV2
iGKnRk75ixuCaVvw8CBnDDXRcm8fRl6WuVCoEIuvP4H5SpbOzweJm7w693M9/D+8uOTl56Qq0poL
aLHgVnFtO6hgBuDkgpr/s1V0UEv0dTExjdFzLrFM58IWe9GfYoShE8+qaajAs4oewipRGSHjsowI
cSwAYTJwWtvZeU/2q0YjOEbS9gMFb9RF04Ujbw5E+DlJL29BrjlA0HXgTAJJHBh35Q4m5s2+NmJ/
UpH6AtYlCHzFUY8/Ncq3EKYXwtAUpxqLTKqZb0cgOTjtgD2q4Z5CqwqLxEza3OhwEu9pZJOJooYS
xCEdrtNr2U0HlcGGZgFL7l6u/rftTvn/tQgZWi2P7clNkwP6OzlInQdallm2DsD4NaG/4ZVWtmgp
yZNlMXhvIAI41tNTgEc6iA4p4Ald+F5hxa6ZQHMQRnEP+CexTXzbo3f0D3Csrx9wGuinRKXglay+
K0lhIAhGk1MsKUEomDOdgfurG5ZOr3FjWKw9cAd+JSUZvKIWfMPaYPsKjX7wZLg9tqjn6GPAWUkb
mMmBSNq1gKEcaFk0ifBq+F32/zBZRkDmqxNmNplfL850XeO+PKIT/VRVOBAkMKClBwQaa4lWYMFb
Hi/d0hIVJvt7rINdaziZHNdhAgOEOJ2sVF+0LNAgD8BsPi682vckhoCncYfk3Cc6P8rQZsYHSlKi
r6TwVngNvc6u2XFID8gmwDzYN2zz7LCjcxa2PVY51IXIpHLu8mgUp26IB3r0oimdAeVeTiALlW6U
1H/kDM3aHhpQZHmkO5wsif0OBpegMXLe6p7Eb+sC0yG1XUPT6vpnV52WzmCoYGy1/XDomhjtV8bL
EsboADe1RmhxQUP54tXYSqvnFPborBzbaP1ah6Zxl7g7SR8oLZBySrJg5VhXWTtLHSit8+Fmcifb
i+V1pUH1+WiWjyyV4qpkmbVwPnCP9NTQUdzHqg5gClNltNWhpqpBfHqiZZUSgPXMV2zedDr6IKOd
VahHkyCgRdfYuYbj6wNNPMW0D/Um8X/GE3cDMt6uujexHn/hOkBYZNMWzQInMsd+U8iGwRlVmZXT
B6jRqvCKVn0tUM83z5uSp6ipsik+1wn9t8TB3ZopBnnSMEuZr4xWyDRMK7jH1qnR1RCAz2E4V90j
8lw/j4EynBlRxeH/eVsD24M1WWNNqd6Qjd1j9MjYJ1vgnffpVd6TANiJQZAYA1VJjawdcKjc3VN+
8YXhzYhropsC72oaLrhVprQseh2jzIqHOV1dklJTGToTIsRXonQMDFcGyKThaaePa3/sMClZ/pf/
LiwjWZuW4Bw1bRNFsly6KVMcUaTwYSHhkDpe3jIlm8EqsAhVh1RktDVqMUtRQjaQuzTJqpQ9Fond
MI4ZkY8islgczLole/1QCmPo9Hy55SGfmRHIU6r9qdef/KnPDML1HAXWLy+b9lcCy1qIQDC02oTR
QQbTO/V0DKLLUL68I9bF0OsvSd8k30oqlhJhsNzFuNcRxzFVFKwxHuhNgMmyNwuvggKfn3KkGTLA
znSoH+IVGNv8Wt5sSqvPrns2GyIPr9wMvyjY15KhszEeXOWIdnr4N4ujpcKE8i3iRbIrS81kOlc0
ZpZd9cXfuiR48Yi0oxob9/FrjITpEPH49bnbilTWeAtQ+pTOnKNwD6GGjaaEIu14aCc/sDX79Fmm
QlN64R+1DPqhZaCVOEUrLWP8XIJCGypBDGWaP22cna1fFploxbV1yPyiXzrrj/kNAyK2Be8Jr9V0
Lcta0hVJGlPe6hdI57yCqOokoJvr8nSJV4LkhyZbsZUnxNBQglkfBmB5Yr0HTu2oElfym46tO4b1
3ahwKDwLdKMvNREqsfxLKpuuEWtdVBaEnQQawHdn+8KpxiwrI8mLpJvJpWnS8EElz7EVdNEJ+qEu
hpX31kVgC7auenfgMTk4N3roOX37I4EEUo16yn0zfIDvjR7Pe4lOiN1cImHxmCUFP5cj83gL/Arv
0L26NXIY+OEJ3NSE5hxcDlDCIC5ocy1KUPmsczQQ93qRHCocuu5SloGrBMKDQARULftP8Otolaff
d2K4+OBLp5Cu5MLTpMnOp8Bp0G67ERwre3gKFtt6Wa+cr9e3z/7UK5i+kY5NsqYFCuIhqwMsb6vN
bmyA1Sd1KRC3tFZCn5cYMWzQV59om5dXoemCIZnfhjNh+fCethTpPF/Y67YgnFJOJDLz5ekKbwOo
69VzUeO6T+e50tn5xJxaRVqh+Ru8nWrcOZtmvDJL13/PEtHPBp8gQb7QDVx9RhfiNr7du9dpIIRy
BfzBLVkmmH5lOfRpQ65Uf6rp6baKCRSKsVT/D4Q4AH9Ak7P0h486unkiaiUHAwfZd8tnsEwvKUY1
EVPniFYdLwdKjkOf4NpKJXC0Ubd4ZRuW7UJ6x2zhtbU3NdvFkH4u0mtbdlk5GPNBN1SG7BzLauny
NgxY4gCSGV+Sh21H6ZUI4cs1nmMaY9ngXgbbY5VcZlUi5xBFPjAjXC/yEtLzr2ImY0xkWd7dLXod
6DnqhjZuUQj9zzo5bkcquD+lkhlnZ1o6pRXdAgX1P9x7p8UXcqGMUnYOM3xF+h75pau1DhfWwuM5
x5dpQeumyFcXy3AwbXYT7F4rm7VWjJEp8fScWHFcu6zI8lrrb09sGC4234Fm3xr7x2ajQHSDmDBx
bOrTp3Fj+L6/uPsbdSS097UgFp3CefPq9UYw55JgCbZh1vogQpMK8D08uI06HcXY+ICHtDNdhRVv
J0f0hyK7tmXh5S50zyosEssA6wKCb+KojSi/C9HbmdX+/PjUqV/3WYi9X3XSSYSglVgEgsRTMtDk
Jj8F7y/ClXULeLbHJqY3c7eqszRC2EUfcYSKRP7U+OU5h9oLDA7bQF60yBgBhyDHyFH4OW9UduXO
Ldn3+ntj6XVQRevfd8zwEtgxNE161AeNrA1jk4fUFAeTrkMAkQKVy5wyswWfwnvSq6xkYGRiZZHY
WoAhag7oH8o60mb53ClqkRVnpaCxi6BAGKp9Uuh4iQfsNIAMpxuJclQgKPwKQ3pdqwCp9SWwcbo/
7IGHHz5jf3AxvCP5EW07Uc23S9LCmOfO7iEIaIY72qrz4bn2Gq4bZ8FkuCX378gHuSp3xmd52RSH
IxYFaTLo57TgDw5kHy24G7ionBaqQD+ga4QnfytuSzqW2NmvPuUUtEIIWNMuRG5xNlx6WmYOZ5qu
Hiu9wjBk3yikWKBiGvJLlH0+vNaFzgi9DwsUqmhNZ10nIPROJ3qgoneOVe5PcBiyWyg3gT62epQN
zXCYnnIBm/dmVIh3Yb+r2TVeU8bLSemM1WWvUIwT7S5cggG5xL3Gl8vRPnv6Ai9jTsKQ4pwF9aX6
GPUz0Zr3FRLru0jIj+y5M6eRHelLSS1MqQD1PQmW3XKv7+5VS92Cyp1gkuvM7REFRzyreb26Gm+R
G9MLH5c5Rcn24sDYVHCbIzcB23nXMRqYZazKCbMdfJlhCnIbei602Tt4TOt4CuUy+8rhJJUCu484
nW8rapVdMz4HsRUt58xhCb310uou7i66Vz64Z57mfn2XFI2AHpNc18eFGyruy3ETvj1FampQo+7i
NNsB3e9tsrVyuisAcjrGiS6ZKm0tIGuyr/51RKF7NEuix9dthjIvh7uOhKoTzCGVkFysm+EDPPx4
jZwe78WRpV1k9FdkPnZ6keuIUpSoLrwO/GGoYtG26d+Cp6PfPZ9aXazCXMWB8DT/41MZWydFm0Rb
TJbo9Lx9/uAXJMtXOmDZxWfU3fnMtwuANUX2cMtZvJXNh0Con0YRhtgGdnaDEXPCQR9/P1j5AY3C
i9lhpJmiHY84oRA1VlmK9pCUxvmDlX+cnqQyRnHk/gI8PMZck2CdbAPmX00jn1irLM+69jDMiCH5
Li6lYv4yff3pVYEHgyRBRl4upA3g4c5/V246kiyJrGmZb06vakbvUxEQhBnBzNqfRHUE0mncgbA7
7US2Q8+epYPEx6IfHG7aiWwGylCmH4vwky3lxxhXIxbVFWTyKTxzEhp+JuW6JhCyHqsMkCzYk75/
OmDKogGuCfdsXfv1HygKipI6b/mc1SU/7KWbAHUufJkUedR447EaPGn4/VLJJTQgsgMz4Ngkkahg
hpAhHCn+SiRILZjN+9sUZz83M+7MyXNozYznh0sHR1xYspnj3gD9kmZYk7JMVBvhu5z7ZboHungd
UyiPLGdC0HxQv+hcgCxXDdpndT5793nJ6ltPUoWSeB9w2N7ZcvkcuJkAml2zvv7SogvpqhzAsYzh
PMtIgxJl5i3Z02dSiSsHfxOlJW/ZLhfb1W5p7/C+jjRvfOuIzj4XGXfwzLO/VRNW25/rqtu3JAe4
UNi58PZ7u3p27rpMX+1ssskPw9vtF85MVAzAGiyOgW2hDKEO5Q122j7XVI9ti2YjL0EMJPlcYQPf
4X3Sc59sSWDP4TLlTPOpp4PLl6AHi8Y623e/37p9OcXCNpuLH4pDVV0t6D13aabVnq61HLwioAl1
gwWWcKaRpUCPuB08VPhbSVNNltQaLTG7ATAxMqvorpWg7I5cz34O2RVcM7LKAwLuWrXKvdBg0I1s
hWqeYYt6PiCcb9sixEoDKBVRFh6WQsCHYUOxPa2mHImtAN4LTNOd3JdJ6TpshH8cfAPSwVdaKEnl
gMEDHVf9uLq6QAHGV92kTFW5Uiow8vFrUG/TP+vGYly1AUZ0RKKNfYUq9hOSbw8ymOk1Nuzr5iq/
i6Fdxp3R+u3mc8MofUzt43YAy3wqXBA7g/riTr9aooGyTRmM4GHdmk+AJaXso2jMtrtdrPGlREOY
iaw1Hb5Y7V5LNNxT0wPoFIeoYA8dkIBQ5e/GYDGYH/voA6oXdkJukEh430gcyah9ww5sPRbVHvPA
exgZzmX+M5Dz1AzssSAlfxUB9nc0r6fu5I/GAiHkF+a8gcuyaK5xEU/ga1TUl3dQM7BFgtZbflKh
ygEBxpp2a99V46AE1jLKcKoXvl6CHcjml+mZ/2j06Ri0wi1c4XV+mz3NRUbREOHExYIDyeJaLAyK
mOdR0w7r6E1hSg/AJviepJgj6OCnBY9TE8oaUkXtrHeWCFr+Jtjji2s6QCb5tvpGbvg6zUG1OlUc
NmSFR4uDvEDDjnMUeQX3IWT9CesLPoh7JA3We33yrlOuJucawMqGichPVRPFbg2K4fSCWKDMLRr4
guwfFy/Wqf33/zECVc+hKgtFflhpgcno+pLqQ17xltbJ78Scg70r+18T2sHEyBn4XApmKv+woApA
mRr6yo9fvHqpgRGAjU0zeAMUmE+yaxDfrRkqYsXCQJl7a9RfopqPB2NvkRxfM4wP4qJPzTfz8DFL
9jiM/wgtgU4sN4Yl3TJXsbQmKt0EcREPHmbPc5MZtw0gL+71Dq2CliUz1Tuct9IaQeTSJDOV71AX
w8HWBJUsY/P+EMxbC8yemV6BbpZDGQsHi7vYyPqpzLcjN8MWmWSx2A8YECi9G7cBk4h9CYgQR1c9
4VRPL87ep7eeZvIpeFTFw6MZrXLeMDpZr9PXqbAEMjFlIZ04KcVmseqow+wlKJaWIfVVFhtXJXdK
ePTnRPYHlQx/KgTlLQVr4Cue6HHygLjdR015dF4wgbAhMdBqaNp7MdtyfycpwZP3Bxk93ysEzZgm
IftEYYRja56c8kM916ZD6eHH3h9icVnaL95rTEVYRsxFyUSGfGOOMGDcfrdpIKpo5IeVYZcyIhCL
/+NPSHUcqzLEzIwgN4mIERbU7yRN3hrWUdnGk9EBSfeodsun0oQ4Akd8bX2XJ3ZKI+nj7taKCVk0
HFMta3a/CQ9XKN+xPSHH/J5LRMYnc36ZxjnzRNdRyWXOf7D0YRuGBXLDMHCdE4K3kffAKbE9swXG
e26lT5NltIx1yjNjRvXBVxFSup/6OQ/S1Nyr6tXD1/jyhTJ4mxsmSs8Td62fcJFNovVljU4e2OoY
0KRsiUyhp1SerulxAepYVoCxFISwiW+p8Q77vRYb1Yy3+cKiaTH1mv4I16Nut/sjBshYnWg3cwtX
pqspl6fBV/AzrK+FDJzIYKMv3rTJxUJAAZ+deuVWBHaF7XC7fYC+IA28WIUc9kTm4CPErdCXWO7B
WD/qQWzomHbQ7ULDQaqTudaYdhWbdq5lKt8bdS8s0E2zXDFwBwFYaQ7BzRfXYFxRbYXezH+hPF+j
hPSudIhTCHSPHUN+KrslnDz6vtBfjrSazjFIEHcz/fImrfAgOKZqnAvLMnfip1sSqaHqDYQvsjyg
9ju7xxGRHySAxe4AaIGg4sxsuPNR3LNE9J9T6e/rcY9bGN8mGwOR/6y1J7yQklTcAxGtwBh/cBVE
VYH6qfX2+cLXlNoCE9tkZ1KMytn77vF4AvfTlNtZQ9Lzvlwba/qAyK7ezmHt8je/Tp7tqCe5wbyW
3Tur5V5Lp2OdGZqukMge7lhaz6fVFxEZEhBp0dYKSjSQoRa4HMD0fqpBv2ww4IjzaOsKTjjAaWnG
9gtEMmPL9UXlro8c35uyoOaQonlP1NXDhXDnAka1fNyyKCmWDe4ZxixpoGcgFOr1ZAra14RLojhz
TAz4W/hHJUIGtoY8jUPpKAOp+n+5VRBuymhZz1C0YVHzjcry5DuiV70wQXJUXwW8igxmO+JSPWRR
GepF6TJZu+OaiutDu9TPai/fxgBMdP8vIhAIGEnTGfmYXYzkNfesM1RwRpRVJHNxeg2sXDFYHKi9
JsOohshnIDzImqONURobx8uvC6qq+BKk3/ZowXCFyVIfM+/rnwTdl5GBriBJddhe08j4Ca+zjbUc
WKly5qPf4PvcrPSZXTlQMza4SxeGl7bGIv8WyM+POsyItgz+wF/rzqp+Tjxk0Nga5a4+Uf0lC7Wo
2M/0AsCWYjdJXZ6szACGn7+UisFspeVThQ6yww6E3y10gE306kexyMXcZyc6fStg8P6sB41BuUfD
/lwnaoa+GWjvnvETutfEUxLFGWnn/4LAUGz7laYVu5ruFq+cvc1R0PDjI7uTsFxdqpGJys3lroNY
X+/64zPsf1SaujXnOLrReKowF53VN7uf2hILQiSNFAGB5xaupdLzqb+X5NTKq1qpKGWtSiyUGx5l
Y6uZfT+vOISi5CmGxEPAXLSHul5p08GeL/ecSHIAz8yK5HnrPdrmyQX367Vunqs32mmM3hWwkFO7
BrfLPNOKZuTA0z44KF1QjUE7ijftO/5gap3YtmN7DeDL+fPNu1zquokCWu/4u5qLFemxBqsB4UA1
XziKH7KTkMvm+sLWw6M1fLaYFjwxTTk6A+AAH5bui7ETuktL00geOHs6cz4W4X5xCiOEW4HRxrRM
WWHveKQxe7uLm3iQKV6JN75gemI+GAxfEWfu7AlQ+SFN8BE0HVBDPCoNV32DbAJeChrnUgzgY7t+
cAp5clt3nwue6BLX8tGDkdz1cj2sR8dDAsSOdQd+MLzeQlr4H9DS9uHU9yfWGEh/F8s7bfHuLq3q
mlgnCR3YKfverKrWzvoL5g8lO3WvWDDDCT5nQpQ/IKdShROrp/Y/tFfWGL7PZhOO40PA1oAyk+WW
XBOwAceiDNugIe0fRGlhA1APR5JDr9HoLch9J3MliWUW5WhD0t3/WlYC7YpYNVxuAov3VQVyy3ET
8JY5Hv89YPJIy+ACicV04deUHWVjjK69rdSeQYOLLw0dnoR3sD6JtU6CJV3S12iOG1sVszJvNnJC
wHCIqea3xBPfv8ZqG6rhdzFkcyWBDDXthW0lyFM4uAn9x4S34963sFPbLiko095WEgT/R8YgXn2s
V/R9Ecuz1dgzGkzwXG8BDjFIEK35hLZ1aZ2Zs4BKTPM088eISit5hCrRZWgvKlh96+XTU4UXDxVS
GIYvAzbCG/muq1cSz9nh31C+wLxRXIecSsxEPXu/Djo1vVqXUuUFmTn4ZcENO3tuv10xl1pLMd6J
/1y1CmditXJ4EDQBjBaumy0TWNP1KGOERDs99LcPp1awBEHsxOTiugXM+dHXu5zqO+j3cTCEhgPA
PPRNgXQ91t2RGh0/M4Vyhi5j4aJHkDXE188DobgYPCVOxoV0zCd6B1P5Dvt436lHxaOFNInNLbds
VyPnaFn9hBYhV6Y+UM6ge7nghG6IGCDrUx/uoJP4SVRyZw8t9MHrQU8YAwdLDTOhL5ZIxkPBdkPg
y7HdBU8YKkXGPzHMZOh4owkeWxLJ8n+sB2qclUq/jzkmhD/r4EIkwxNsaYs/pElyJyuj07HE1bE4
FNw/9EExgM/aM2BdMWHunFM1OUfrl2MMueWLBcX0iQG4+gG75ALwerWlTcAEtSNp5GT3uUPvFmAu
ADkFt42zP2iZuw6Ln8zIy+NdP+nUOl3ltaM1ZpSFhjW1WvqMIyCmEtrsCymNYqKZsX8LMo2kNyjJ
iOhvpUF4ExTeEavY/8DbVoy72lf9Rdl/OeWbTouDT8GoRi3AABlQUx/JyhsnZ86hW69ImoMZ3Q5P
m0i3X6ajPqO8XL1OfHZ4ukJ//vm46XmdMVhEPxoC6nVH+W8J/P+bWVHJvfuXYzOWUz5lVu2FWgNH
8oz9v3+ENFBDNaA/cuI4KpQeZyTEAnVyVRyLPFN4S/5VHPyZcdjsa4B4usbDccsXqdzTmOoqz7sB
c1n/eRbCuzLULYbrFlee9oM4YLAvO8tl8XKm0NevL8SwAS6Piry/vehMzFJS6tjSsUagl4vwpa3Y
SzurzfxqtpdYtDu/Bvc5hiDztPQXFLmtTDLBRZves25RK393obeCwcou5SY0ph1Sw8zF+12sLZxJ
+OTMwYqmtPWLghew3yzyIkbhxyBXglqDXCYht457fe+k5kzSCePxTxwVdLiKUu7UhPnWoS3BQtiE
q8f7+7A/SNa5oGLnyRbGLynLE3olbTkexVWBHuvrxMJcHru5DPpBOh1I0wPCrbJ4tJyQqks5JfCN
DZ9VkMJTQQAi/SuIjvOU7/2y7PdZxmqBDseDQrdT/nqChh7ciSAzNOgPLdrKFmEW5PMLYMwbsjO2
IeYigaUtyjir+vBKOODcSw/ZoEBhhNQHsMWjP+ViKjqijzzQ4ULBulhLkxVvWdxUbXvr0tVor+wG
zauhmHw7vY4A8uubyx+7W07MGBvTY+UXeiz+o+m27sKbQGRWBNI9kcLyeLmh9Gjh1KfshNbNdcU2
LrCgjiYVy1AYYytS2gPvULVhMMa7T5DgXzo+gD+kTNgUgoNZJj9+OkUmW5vEZgXHoVyRRw/GJdl6
BShdOCC5wMizSxdjEyys/avf5nWrnBhtCiww+GJ0ZhQk77GrxFo4FDvLMwtoHyDv/fBu5w0twXrH
Edldw2g+Y15uFU89F9TKmKBgB/U+F83NUk4mJrqXsYycbT/mtZ7M2po3NiMoLxFGuAAfxEZfAw8E
oboBLRyMZeydxNJuExSeovznhOZs5bxwzAB/Ifl/9zP+DRGmq8i2rhDiUTRpl9am6hOUKag+cigJ
0X/93E3W4eqTMlvNAaR42euQNAfpw/CAPf7P545dujJa3z+NouWoNaKv6o8UNg7h9srz2aYvPA7f
BCwyc3IFkUakWGf3nFDXiyu0310rWH7dc0mS2miwI/7YbwT4QkmJVrQWFHAQL4WovaiJ6QEpowm8
C3yqat1IrQ2VCfDcMbNrZuvFJ/FGK7wKcV0h3PlPg5K8f71nupZH/Y/BbX2MeR9/XZTDWGPyQ71A
Y81X45cmfg1VNkBcvP2+zEONTa4KG286wUiRimGS+xWC1f526+n8tnJAfem+Oo4Vh58UoC59GlSg
1OjUi9G00F51nDpQY/NoJavlvMdfBFoLGbmZAiYpwhXyZsxK+painrADlL2ZFK8nc4npaje4TNjQ
ybToA98WfPpXsaqpLqmbWt/iBv8cZrtOa7olCELg4yeiDxCjUHHMHrFqTMKEK6B8hXc6XtPbBr1h
x0jvUsq0z8pREil4Q0EQqPcxcbSMY7Y+cLxwrCQhibs7aJPx2egJ3sCdfqOdQ/jmM5WaLQWVlwId
hvqPsDgvm4wtzDx3L7GwQwTKcWshorzBKW9TYG5zrBK9OyebzhaUx5vCqcYkpe7D5MGZq0T10tvU
k7OwtpfKqvU1d8GdRL4JffR51bhVOXiEr3pUWMEORyLMRl9nhK3qe60jWqox9bVrTqgp2SQPxgkB
idaLgxcemAiAMarvBFvSGX32d6N1ix1vG9bYtFXOqKTsv0lrpBXA5fe6JPy3owWKaCrRfE0UVGd8
065+uiWRXfQjTAtX+gK65CNmOB5J+lxdrwEz2h3gdLRVcBNYGpBSPqo/ynrLvp77ZlO2XED8gaqJ
6a7vq3/hDAcG9e91lums7QiWAJMlu/fgTapcBA/ijgD44hTc0ClcUsIPv0iGT3ah1IlpH1EACzv3
6Va6nBptHWSbYXVHCMeYhI/FraBKzbMHtKrPZmatPT8QNvH9VZOQFtgl72x/C074js8V2i9pPOLM
9fURHzhYFfKN3Fq2IU2LQJoaSQUrS1FSy3OaOgoV90HneI6p7RL1qZ1wyOshD+Qx8af9KSewXHVm
jsddqLBgsP0AN74AahUbTndmidg19SavOBcE+yx6Whu0098ntf/PB9kyh/1d/KunAr/JPCcbsaYs
tegUAVfu+VcA3CRgOkEOKkhpO9L2I2HbsHK0Zk3e7UC1H9RsL67CauLo4FcEhA7zG9iNUZdBqkwU
ZbxLlFMtH64kLqLQohHR9jQyDwigeg1eJEHE39yZ6ZuAk1OtYjQIh8yV9EgT5ax50XNpPRy2EfUi
6raphdGCQyMI+uIjYehSinzBMpVtu6vtnYDojuN1ZwjyNlktLUTY9drvxRoWn8SwiJ6T298w4F0u
uqCE1UOdukR1ToJ+vk3Aa0iBkDviTW5ED3hYDUGzKzHZ/ZaUOG0iDst7TGlfH3jvlRatPsU77Ygn
bpqZUA5eAQqqwxdF82ge/ypWnM871nPswSwG+RXvOsPG+wXEtVI1UGGKZcgpoRzn60yPdGFhBoYq
7bUGR4X+qgSvNmWRTo00ERfC5cpsuTu8qESexXSKKguv23CrLm/K4+DBeNYLV+MiIqVx3hhPmLRA
nqBeVWcJqSk8a2sRIp+1EXmIR6nY+g4Fi8BpRK6Wg6/AHGNFHsxuwV0q1AMMuZ49fJDQ8RaffEUk
aZE+5UkLNZH/4IOL/tzEhE9xjFxLreKZY1RGr3c9VpsQi2hi/QFC6TJoTGaAyNT5XWjwuygsIqhr
+J/fSJpaswA/KKbMJ4FL5JO3sfpec4fAWZFotflI7JijXIOJJoBa9kWotd0xQbwdJPcJsk5AED7B
1la2ojGfUzOWfO9anWctbE0c9G3KqlNx+QcaDF6dTvKoiJWhs03WqqED98yY/rue1EH74ekCEz22
xt5tGIhy2NFQDRzbCcsCPr2vYpWLT+cYFzxTo9+1RcZWcI+CjnMDJYpADbXakHd4VN5T13/TOA7O
dla1FmA7jsgRArfuzehuYe5YRK66D7G6tFcbzYvLZM93yOqwc0GUUhgiH8XlF1PpwTJz90Bs4h3y
5tbd2WuSFPYxpOVqfkX/IK2imo/0FvXkdiatDgMJBmOtaF/TNtYKuJ6NLChrztijVA9G6uqqcqjW
pZ+O5IF8fsYBr/84FGHyXFuwSBFgagRrX7WjSO47n+BM0IeAP3Ta3KqcCHpEAUe5vt/whvp4na9A
CA8bWDkYFGn9vzsmfNd36beyr6zqE0hJ4c6YeL2ldm63Ovbyrcaecwp4GnZsaCQGrZpXq7q0W8xF
gpF1qWCbhwZlgmxhc5X4EhosbqmJ1t7NfjE/UDIFXCQsO+M0bsE/EMRnP0j9qpDZTizetpAdeEDJ
SHYZ96nmr2eSIVrNXm9fXQxco/lVR3RSRb/ZrYIBogLAzy1f2HER6ok2h2z542iwhmVZ5ACWJodB
ZH4QO4TNqnew747ebRDX7lPNUdEKbhA9jcYa32+ypvHaEVdrSK/Pb9CWUGVun0ZommUKHiCyHApz
pdLF5aSAUlTPsQq1rq8FlB1qTq0n49pwlioFa0BSvmH4JAZIurUZgMRD/gp2ms8cg5hTdrg31xr9
VQecv4FWjmgTuMspnFCRI0umA5V9x+71wVao+V5y0lTsAqmCfOz0cxCEAN7ZsmFLFA/Ux3ABF/1G
k/ZOYU2t343R2s9/tNrwN92Z9eaXosh7ev2huSOV9FEpU1DyVJxpEEOkdTEh52IHJrl5TwhJlaYc
Bb8Kh4isGfwHcWvj/oaF6rzq1WLefR91crRlcOVNPAsN5esxFOV3riC+fJmI9KRbI6gqsV1eSutg
w8R/SIDT16Evg1NEZvbc6LFXchcmDZ7Xx2tBfaVbPXjnaDJSdL5A1obdFwbfA0NTcyjfRNekaiPd
ivjB+gV5adQXDNxxlK4mHimMBxaA5u9ewmEXukmUR2esPzFuEJnOQI+Tg/cXGEyioTKW4utP90Dp
exxGTQQfnnk8+4OBSqDgxN8geNflfhKfRfPx/Bm8KEINWlezc/el42hGECN6P1DktVhbV0P/p3aK
yL+LzFRbPbd+oqJ/NzWjmjn8MonLMOp9cUdmlD3XL5JqplWAHZp+sp82K8Yu2CQvFoOGp1UvpmL4
+7M8oVhhYCx3Pjd+f1wwEfYmYhCOy3VSuD0QpZ2HNX6d9MrBauHGRLndl6cdPSvlftecQPLGGmyt
OAaMubgwvx94CkHzxx49nexjpXhpBEWRbZUgedcI0LE+wLpENlITDr6NA0AMbtRwbySa3negl6jK
yyFqQ9kYIqQdO7C0af89S5pIvdVVyn+AE8umhxX3ju0/Rn+a+SmTwAuUY0EMuqbNMymuYpXWFD64
FBZ9deNPXDCxNPCEOhYLVgdheyqy10pdq7/8cobhc2WdmxKVNS+e6Jlo4YQEP5I64Wx5m2r4jaGp
kmM92Am+rrM0YyR0DeT7lxc18daL6OxjCtbwLORzzEongjONZsceAvOKsXIYHcH/j9SReudB2D1g
O9K8JzMpJRdxHj6lYvXK/ABhFXxyAuy4n1a/hCmsfi9BKHMj/PywLHNYMaDFQzqYEKFWlRc+rENA
ua3u+plTSvirOK7RkNT6kvv7qA88IIVuoCHr1JUlwES2143mCFZLiC+ViGHLaC8D8A3zb8Ob2Lf7
oC3uf3PU9TEZr6fG/B5ayY8ysTyJCQVCp1yqsExhiiQ+mqaqOB25rGNt52ZHceTdgWdgmGSx8+w2
UdR//pAJT6VvUxRcq5u9V8T0KHAA/M1d+8UVomRHyfYs2dxdDxHDpyrD9jTJUzM+YhEiwlyiHLaK
gVUHKA+Im5kw+leHiVEqx7xFnFhdpkV7tHiUS9mBZtbZOutVAw+t5dQs5N1jgqYlf2cSi2x09Iu6
by4Sb/isk7T7SlDqwxihBj2Dd55OcP0s51lJCYCmaEkZgTeoSt8Rnj831L9EoRyFM0GnTH137ncc
yQPPFo8J/awG6GxvJ62i9wtdr3WhkJTm9dXujsn7Ro24xm2G/iJnae3Bgfn9dIR15B7Fk6O+7zeW
lIOb/Rz7SwPM63a/eTcK8xVodjxMKMVJwruQk10BLo8ruWXJE8uxC3vERK/Yvcz2vs9DnnQowUwd
5Yji939QVl9hFLkDyRifSsIIDph+CW3IYkBqnAXdf9ELMtrxkPVWj3gwZ/ys3VqDYEeUxvKb4Bza
wVd2tTnY9c+ER2ekuX6/ndFuGocwBZmpYq/dgaUwQeD+Ocg/Q5BbOiXEZBJl6xh1tOM80ePQV+/9
XKU9EY0eMONVXgOWSIqF6YPP1wZULn7AQ9NkpHBblDlab+4Mhk7X3Jcwn1b3+e8VDDeGFagzjnSW
+we1C29BNivoI3vgDAFgI/1fEFZvwPk78HWMhuHqVR0Jjg4ev41cU1dmCVIpdpx5cpmmnhPZzOeW
EaG/njwG6tbPOj8PkYzZ1vXknNQewstOPeXkqIkS9PnE7cXp1nMCN9bCuoIx7FtmSE/aJPJZejJ2
7vVwcRDK58ChWm9KSJ0nR/CGo0bCJJFZcOKMOCfPg1SbU8o/6W3uDCMS8t933unXiymjce9YoJ9D
wdM3iWPNp7q+8AIK174WgWEXcjyFiPpY2/g615M4CX97is/Y8l0Pd76w+P5BEqqmxYDZ83Ifr8wf
PwkhOX9Dy8TXuCjhWhjMUBjNUrjkPTyyqihK7otP/jT6ohg573wjOzBhfP289hx7mfKSbWi80Gu2
FDwslQq/BKLwQhuBYF85T/BFB8/cS8ZpznXNJ68u9YuVNwLhsiqM5BL0c3CiN/lKOhd87TbvDDWc
W5nX/eD0n5vQiLSn6CjzwusUObC0f+7jxsf2IIUWFQlh7y080vpRNEjPIG14mWhTQXeTfCVAcC9M
xkkVIFvR87xlXyIpwyKFjQKeTgtyLwUbTt0NlhXvyNLwJ30fHEiiNrqEDjpoIAgiR8q9wv8FvOA0
bhBA+ztmuwMbetlKPA9J7mScJnz1fZmVJN7jthRTjMfBLgzZTn5Uw8erBLVTHPiDT1IsH31/WlaP
G3/mEl1hxzQCi3vRx0m1QaTaQXfe9pqJV5P7XwHYxft5PKEOq/wsYbeRZPTkCUXedL6WTpyQWJ7M
hVk99NsP1/xpfSXRGxNI/K2Fo5/A/4isXACeVuZwXO9LNDDgB8uTidkjwwlomz3lrhsB4qqZuyk9
kgaxum+2374TcqsbsgEn3vbB4Dy2DgA7zJkYK3A29TkszPCaViGWJt29M8fu5sHDFXbO6acwqgeg
Lfm4idrnU/VuLEuasnkuRhKag8wDmXSWgfwDKamp5Sc+608mWOo6nBQ193ezHrInLIckZB6+CjpF
2kuqiXzGaxmK26HQAivQC96d08G1Xo7g3TBWu0sZ0n1qQW/l3BEdMDIYn5FoApX0J4i2NkgvSfaQ
G9WEh7XQZ3XwBrIf6fLMfsgqV5wZWDUOJ8X1iPYKql+KPs6CEC0O3FkmgkWhM0Fr8Q4N1Rs5pzEq
mwAUlvlWyf15slz2IYshuK5jgArIII9H5PKBFc4ehQ1g5viJMUTNUF8Hn+QoIJAJ0MMFXMBtf9VE
fPdp3pMnpHoJDiIs+clEm6Sj1Q3tEit9mEWo4d8LMvwHq5Vq8paaraVMzNfud4xJCK+9ijxoMsYd
e29FDLjYnih+VB8+X6KLa/bZikrF7rBES9nBiQNvKaolqwS/TpgU+/IvHkQ3reMnMJUeexIb9SuX
o2nDF9GQyhTznJuGqGlTmJ6XNfEAIQeWOgflPeRS5GV7LRKvoOh/BVKXWAhUZmkZwEIh+8dTDtxH
JOWo8qo+gDgV5axVjp5jMFW772UncpGmiH3L67OjVWqk6w5fT4pfIFZMHjw4GjIns2MuFMkPbJpx
g85W3EDMwm86SdSNp0uCG+nnH8gpzfiBCqkvc2gaCeIvZt7lhecwsLRxi2y/HVnK0DekipRXNZFX
8lRw5kafJgIG3rihvLBbwjMJoeqpgHBPnOEEnpmh7xcqtPvNwVfRSnsX2V6NrQ2CCdbwh7ANAR1Q
Re71vL5rcJjS3qzGYSw83UvZ0ODTUelgPYgCbHAOvea3PUIK5MA4yevaXg/atdsvno0MOSv1xiNw
S8T0b8qMZxEjE7sZoylbIiVRcndF+cZca0+UEoheuQ0hkyr2lfYyWkrJe99Zk1HaSZ8lqCHsWZzp
JPDLiUtc9iE8QhAfR/LqnoCfifls6ZgvM3Ggnw6bNPiK51ZKKKvFaCSX7Ij7eYtdX57/HItLY31f
Bxlkdx7lMhCc7scz9G8bCTMaXhLdishSYwgCpt13ool6RZVpgPLfJtSX1XAlm1ne/+lRg7+TEpd0
vvGuqkAL7kFlC6yxJbI9eTPZV1cZ3xNjwmx12wbIdn49BbmoA98dtFobU7k2ycxcodCdb8nNtE8P
u89B1wHhjOno6j0A86AhdY4tLrCFS0aekpP3v1R10F3/u3aqvo7e5mpm6yq7qZKXbOWgfsTC3gWF
GeZLu2nSBB9eRSwluMJvCqYVMlh0nevTTC4QCn3NoiSWnhMgDhFSw3ajhmL/SDoemY4Tkw8gJ8E9
yMUGTOYmmgYlbPXyyvsEh8WUOkF9WjfrI08/xnJILuClKDfrmLtSd/LrYGjqPA+6x0m+0SIutDsr
f8l1DQovm2k19S4Wmng2aETAwaBBcQ+K7KA/p2NLZEHs+VxNiYPydjrS+pZzFBJFKzHvTBhYXO4K
4WN09Sy3xmBhwFUu39+8M+qxMjZeWKnRyCSxHAgn7RHE7fjRi6pvTe4O0KzPZWAd4LHg6d3KDrYZ
TJfh7A+a/GEu5eEm4QTTWRGZQJF2GildAZi4LDAg8Gx/55KYkZa1aywC8GVW6/fm6pUaYe7iFyVC
oevt/4GGdL/rwyZujmKAwuCJ7Th99nhkPBrVCkpbTI1hacpTd3Y2tTkx2/vMBBSHyVdwSCs1yYuq
EBAxmeCayxBy/kR/ctF7dJAxDLora+S8BsSbXm597aiF7WBXWKZcTeFpO6vt8dYM8JnXiRuFVMPw
inbHmQLERgVv1CLsCAJOH4X4Wh6/EEXA+4PsRMx7QWIYonIZAoEFSLUJnLTi89L9XZ/IoBA+39K3
gnrE7JBAtVm2Tix2Ugnch9RMZnqvYmXAwLlA/6ay2+gGLGCKH1nAO2yAc6jjIipnHU/5fSsKTsFP
TqSRuMfq310BQqpis4FcRsu6wWsLCjpn/RpYmnkqYGCNSDQRde88mA5AstdYv1cpX4avR9ndBqPg
q4a7cVii/yJZJ8oRSvoq4qlsvzGi6NEa2Vmyo5lx4W5LtABzSks41kuNWtoRAlUenYVfFCgpGhxE
ms/lmaYLW5gvb+iXzTr/P8xujtpkzv8v57H0gcuIkt3qinq72+w1oepqUtU99RveBkoFKAkFaTGD
g28JMuCOR2pHIjHFazW+xMZ1plvMjd7r9xojkcYefyLc88DQevNtum0DxjcCFDhChSokXkrmFkm+
ShhaWhkOu/DqmE18A32qwFsXsY+TBFOIHVnMAOVWouCfFwOsQn0CgTU8a1W5pSZNJgJX9BF6N7aD
U5jLNZjKOzyYX15vGivcTa1A6dovV+7cPk1DPDUbGen6PnTU8prQt079EiXrKIN2aeJ74knTo2eR
Roi757ZwrMs/yNFKUPZPORc3spNmNhlwJm5Si8rTHJgP2pToFrU/r5S9NeGqWBkC7qJc7aNQL2LQ
h/YRss7ZW5yf+Rg2OhFYKT5FqZK9FXvsS9SacEorkApywSOwndoO+AL14nUdh6tvSiEx5vvnDA7C
5MkMM7U1Km5uFElX5gEMnWC03op6exQMzT3tpoR+f9c+6S4Rg48q+dTKzqMnMJudWrwc8OP+AB+4
/R+fIfPEXMPAgJIzcVQCphiRe/9pxAFgFmC9GsdZCQ4b3P0VM9MtW55HsBSrrmjwvTyIwzCcf+zR
3KIntr1g5lwlL4l8Y93xD+tahBVcTjJjaThCvsPfE6SBfvV9Hd0DsdTBPTVU4vXhbk6glNIf5zcu
MXw5yzfBSP0MIfGLp4e3A5TOZu2xLyBiEr2s3PGdQYbRouQk9Zqvy0/0opFrkvqlXzyu4i0/abi/
8rWu/hYAOCXN3G6E5vXxxzJBA4iZX1FiB952PyKjFHP9jiXqY7wGX7DRLDfDuvSzvvYmP7j0O5uQ
yAV7+WUC7AR6bOx9FIaqjc0JsBv2gCS15pgFvjqGr0+iSXY+P6+4v/dnOwvtZlqjaVTIxz2udKty
yvK1AMIzyU5qlqpMkcpneb/h4P/DLYbwERQ9W/UEpy5eylje9q8M5XR65OrkimJpvAwKyFNRayrn
Vt05/jqO/mG60rcTqsQ/WWUAtzHUbTKWDbzQKQe42wpG97kr210duDgDEw4uM3Fvcq903Dhv9+2V
7XPORexYLmo1V6aXdOmPE2iqAmx9M70DIwRI2ou4XJXwwY9Fpf94AC/C7QY24A6LR5i9HIPPflce
hiFJoMyOnmT3SziuQ3pAt29XWnYH/BGeyapOATlZBnsswHZVkRmIvV9iYNFS223QSqXBF1nT3gAT
1q7teFF7oLVnKRbL2WXpKX1sfQsTllrDbEsv8JHifC9FaeYQbRMPFaizEXbaIprC4Fq5TQggWDCC
Y0m1mVTXSbwpLXaCvwBxdqIyVmxKuGgC4XO5h4c5lhu/deBKNlJDmeQG7fxA1l1owy4o3JJjeIRY
GS+MDULjoTPG9kt/hjl4D+ib4JAm9y3094RG4j/aQvIBDwp3W0rIM3fTmYieUyxYHqHRRVECvM4Q
sdcolW2Lek/w4f7U2SzSZEuGZeS5qnXbLBce8AWZK8ekqG+yIqizFBL3Vbb3jMAgQ2mtNvRQUFEb
zEuXe3dGqsMcmDk5hcAAZNMgoSnQQtQ9CYCJMiC7lzr22/hyFg0nM3WXBwpyO5ItfZyY4iKovqf1
2R9HED8Q+CWlod84udPtfhihD7/kvk5xxlcRfAelKkRB5ZVhjsVgongFVtiTG4TgIo7TwSY2n3g+
fkm3h60tuQxAs1XzD0KzbeJMTeK86IEviwuV6JzRuS+Jujxcj1ZIHuD7hFLyYfeoKfe440N6Bozw
yB0hodlPtv8FgSUooMZQ4IN8RhZqVKHJ5zUJ3yNh++k9/0Kl9d+ATYgcB/Y1zpUE2hXhnT/0x8Uz
bUV+LDRit938J6jMVsvTWtlPQaNx9O9pkiS61f7vFQApYVE51EsTKxPD2srzEhXiR2Ilb+HjTg83
eAP6cZ3CzqXS7BXG3K8mtHz2XxojShr5SBM+EIx3z8IytpVA/xjPszGiltyXMnkcopWr34Zbl7vB
hFL2I3+GX2hFJObby1PRViXedjkDfrVFLe/2XugKnup6JfoVnL64KM6IicckF+tV95Bjd+dDti6b
bMRw0e47cmQzUSsas0+D7u8Eb0il2t6Rq5mCyx5E2av1GVAG+8XTOd3SDEA2Dq9+vT6nxij31/ra
0jaUWtZ3tE20Ac55e0V3zTwnlTNAICF069JrOXMS2sMmkVcUEXsZusattlb6Ig1Qwo5j1IogFsW5
wR0Nj9IMwX2HFu8QEwhvqw6mjrH1nSOqL8UREO/i96NnjHNv/pnALnSxKsIzvYQhsbiW3DqcikLu
rt7nOtpTi7W3/edg5buIsHl0g3QNw9K9gMfAO707pmcyIR0Xc0xjWwDJWxwD3qJkZp03cEWWlGu7
DHo08k64cTEJpjeJ8IvZT18QTyDB786NrA9+GH08sPLu5PiLhPfVn0sG/p5XDqpPHcWaNT3Y1SrZ
vhgVYb7zkSKNUQ+U6NS0ZNjlhfxtJyB0YQ1QYUYddvzb0srZPxkPdvmXMnl54xvNdKdphHs4wkiy
KkS+kOEb8iBOYJWhhzOhtA2zTjQNSnaPo938fpCyu3TPEFWaLo3Vt0kExnq2w1xv4rJG8NGoxc6H
vGIC7PT9qzb1GskVYsLOGJvN6xYWqciPDPWtgBUUAqp4SDqb6s4FrAfy7HaGgPY0GjUZe6xiNM4V
fBG8EzpgsJSGhEcAwkfJz94HqTBEbZu3YrsM6oslxP5oHJzELK0+Waqv1Ogh1CbV3oL+J0WX4HEs
4e/oaqBjO+mPPrKhuvYaLo8MN4WuJ9scqMkw8cN9f2IyZcbvjSdE9jmH356rK14GUuLu65XHkah5
wVB4haKWhQ+ZEHuf7vbGhTa8YcgR3QKd3aeONaQmFP69245d3biwkmfMH9782lld0DxkP5Bg+8iV
OATE533wqnrjffH3wlD6A0covUxs1PmwP2+ASrPXpaACjgMUIXpVaD1AKPKfBpuhItdyi0J/FfPc
M3ZHZGPsxCHZaefaNmKlk6RVxVkU11n1LcLQPdb6AI6wcxsydE0NphgqOQ16jBf2egaCUffCbAFa
DV23ZcPdkR4cctWmDNCoWdE8ai8PLJvbEndewDT5EWpnhSWe0HqOWutgt+PchQ+j8JIkqzRRGrux
tWnhmC4Vbrbo6RR7GAfforbjj6bdzj2JV76A+uachF1ukrWGK9nUu1lD5+VawoUKv7dcKGT1kfo0
dMLISLMJSiSoFdf+ynRapwc+4cTRGL3H/j4ZtxViP5U5Ewvr25hkFO/8RbhHR/7mP7LLc8ST+arV
VxtdYUcfgfLTt/F/VEsRpPIjXdG/5v+Mwwk3cbovG0cU8BdDdVpX+yA55KYEIfcGsrnd7zdLbtrq
f4XvrgPwbPFNmK4UzPIUNX/2eGQA4EyQpL/M2HF9GYmxKF/QmYZs1Q1DGncZtvZrokt2psTVpNIx
E684meoguZRE7enUzeT+aFm03GFc1EjogCqV0ff83dHHIOVCNTrqtS4s5moKJ72RzFtgE6lOESH2
LtVU2S7mmV/AJHMLGuf1YSwERrwC8Or2efq80/I0Hm4+EBbInT8tpCVlq3m2K2FwDfzyJkarCXhF
nHETj4IMQHRERQiQeHSStWMQT0JTmVIuEBnPrhtxG4sK/wO4gSdUYNIUV4hcL09GBY+XPVIlN46q
mVR8mieWUpFITMs0bexT1OUsG6wz9osclOe1I80GuLzipogVmutKmXy2FgCmeH0Qnz2SBDMJhyf7
zEMKx8Zpx3+GbZQORhtiYgV4QaacQUyJbbAYB8TIsGc85EwMKTH9kW1ZWrx3Z8IoDkuU43yB1W6L
rVEXebdmFC7g8ykb+06yf0Ckxdsd2z5VeaMtO9Q7yDNveWYLZJWrRwZ1/yZ9RH0SBRQOqQkik2qO
IeSvAcUK5pp9BwEek/YcoWSdvfRlw0yGZvytkm8xQJ0zue3XU53nXOaUH4OauFt5aHVe+6Cqt1CN
4Ak8d3spawYcKSA6YdVaYTxaZPPbaZg3KYX++H5f02zR2rgjBPqTBZ9Q7A2yhEOPGiHnOjH2EIee
+IxPTtH6tMlFsC3BRZGR6mflcaHEABbsmZUofS/aMmtU7NN4aDzgwmxAZURLtH6RNVmLVSCSepSN
pkuYMGkffXPIfow1nNJ9gtM4veR0pMtdPvyMwXvQwb8YUSEtuT8h5E0dQZgdsSU/eJ/wIp1OqE9h
tbMn9Cr8ELhE8gtvTdUw771IlCoMDDO68tSA4ysydFtErQFda5U2kwyhCmHLekkKhk69tg/L+GRe
C7tQ8iGA93cgklmWHpPRyXRfZ0JQ7bIgJhfL9Au0OJBR99Tw4pZ61h5404yPi8l54DtWl9iJZJyR
KDu7fwcXtVqdz3IvGRzKe1MOOnetI6low5i8uF+f5/y9sY1ZWka5EijdamFYgiwOxRquTy/YUtKr
uTku3EUlUn4eiZ9XWlZlDgWPZI+7ntesmvysGPBzQo6ZvwBejE1dPg8Uk7XYnCPsyZWP6EG707td
zRZB+em61/GKMOG0ye4p+lJ6qUY42jN9GgJU7oXky78avDzDCfsb93yodx/zQYAOlU5/s50HY4Bv
kTFy5OkOjOT9hTjDvFNUOMS/5d7W+YZKRGWWyUx6wLF4m7Zs/5YrVOSrsBT/RZVSStLjCLdBfr/E
XN4E3JtFbEsX/EHHG5bMydi8Mvp+W7v3ENTkg+05zRz4wivE3mg2904Xk9yyvOu59vmyNU33ypK9
nHqWDd6iu85MZwaDG8ArTCvvD/uoyCkyUnX2ZwC0oP/GNv+JDUwu6Hvxr1i/GXEf+W65DBgk4Wie
U3X1bt3AijDdmW9xmx4NhSX2Sd2FWyOaaNWpB9PtGn5u7Z1qHNyzgMTOn3DDdx3HRyI4ZmViErCh
evvhH3/rH+uTVGpnfAaHQwknwCyGv3cyxRv9aa1FmsxLgQyi0Lp/OirApm0ph6dv9ZzdB/GoeAX7
RoI5iqZGnFKU7tHYZ0I/0DJwx8KDGc2SoA088KLIN668pJDd/FzbmZ/UkMXGnp5tiCcYgxmlrZgi
DK4ztKCxZ18rWfsWANcvtO+PoZeAhog9lazFivDKH2uNACRyTs0KKo2l4oz0kB7wRkxOWF3lMtMS
l5HqVXJBRhU0F8YN1+kWXpF7aFR7xvUbaBeYgu6tXSIe+10mDg2U6+2N2rugcYd6RZDbYVlKaNik
ofK9jTTQhXpjZ0yErYCiP/Svr8cKHg22aLWHIHTgTL9QxyM7s39KP+WknlTb194d7a89eOMS5ovl
cHWF/ox/NPQ8zLcULnLDfDxfShYh9gVNBo334M6dYxdymPGZAMYOB0FU0susVFKwN6kRDDZlsl36
b845VI+MSOi6pR6qULIMvaYGzmGaD22VR1TcKuATevoLd04H6+cr8dRGXn3IPR5s/OEszAED4oD6
12Ixht7p5fP4ld8DwnDkzLPi9B3QaK0IWWVHUrCpB1OikuW+l5jAQFoeiD3/C52HxX7q19xnZdVi
ln/7quOJTEyto/BUWyndhXtfpDD/hvRYRlOVSEekhY536WiAD+6lqfw8GqnoFKebb6P90B8f+jgF
h01qE6kXr0YUXEKOpd6kER5j7fuBusU9UGRE2YONt6HRSG/pieOlCfwI5Fgm6WgOixf80h5wnBKu
jdD0hok1fDseBp3VIyDXrn72AN07NdI3P2iEQK9/vzGydxSeMkMR/caqC8PwkrjYuBPv7+XpQDxH
VmW0NVhi5QlEH/6X8BsHZE5T8lWGtgyu+//yiJmrxmmlTsULK4JivMyOUXHEd1xZ+7t7kT24JRuU
chk5dL5HyzpguS1rNrY9qK1rGJgcDxV7RBd8yxE6dlDjkSCCSmb0ORh83uXYZsSStdhZQacsHY5F
xUfAXLE2vP2Vr/onCp/NCq/I2+LVuJWqLSfmt9QV+5JrwsY1/SiuhXTfdqPNOtFPVhPW0YIeDd3n
DvK/482OoluKHAoAf8wUIieWMuvnrduiSIracBkdYqs6Z7GU+KejVs61+XRv0kxohqllrd31ta7t
Hs3toY4V0woWa3COhXvnyCG5gt6pmU+j/BKZDiOrCkQIfFj9JB3m4nMVnsOBzFVXc37pXXd0z0og
SIWDw58PB7cKLvZqggu1OIMZxcRMmiVG83LzcsHqGrFsBJ3CgwRy1l5ULMZ6eRELSnIMHdzzjw2i
TZCziu2oB1jcqnSQT41eTyqdCHz40Vme6pLJBTO92/cqS7UYv2yujSvkN3VCriiviC+4h21NUnsS
Cw8ibitDslMMJ3UQagW8INmc+gkfSnGquw0Ice3GbPIL1Pea1UZ5fglS+lqjFo/AV/uiEy8AIiEj
BNXJ6tq5iAiQXzXDMDrPsreBm3Sgzbou3EMTTdXsTO+h3OQjEutpSXMlJZ4aAUD+srivWOts/wul
62px5rKyfcmaIniB4aMjrzzDKw5buwBuv7BeCovvE4BqkGgQouDvPuOoBrJRkYMdO9bufspEYpKD
1WE3aPoJtqeTlsAtI/c+wweTauPzpwQWHA+hcFh5n834WNUxRl2XZ1EEKTcXCgrcuVI14e2bW1mw
UeryzSHsRXOkZ8dqvk85Y5/G4/H/BezFs/Yi7CMAadid4XdJoa22acnksBedBmBUULYAZW2JieHS
WG6DQGWJwUnAdY48Yg3bX17WOYoxE5xP8I0Xt+oDzWCjpnQvYFQfh0/FkXpdEThHei0Tf1VndBuY
HXzmTvVthz7V7sFEhBGPpHjUOdoaI6jgShN4a+tyuyoYsgspXsR8v1iZtVhBgMAl4ap9pvSOJJf2
vtbunJMEyCiaLufUygOPsA6Nvxx3mUsrN7Lewt+jCjT3aM2/BYobmrzd6nuSLQzS13wJ1YWnwyli
mCvC732YpQdaTnMAtpm7S9mUoYruvsmKKqP3LEncSYPYzGetnOxZWBZBh88AXhKI5hrpasTU9WJF
SHpK7qnVikHvEjlFVxVM7yd/SMy+lrQfEF4sPhFvynMgkdE4N7+JkeRFegBKOw7ABDqxF+wEdIGR
HziwUNFYxK9zChT905yEmxuGeMDJbmH1tavog72AZJqebTlUkFb2MusxuCpNf/XC7WPduvZcAcPt
ZDvF1Xlj3nB+KqE6yMbSxXeUvjrOCe880akTrop8ByqprXytEOSC/K4PfU6vLhJVreFlW/tVIxLL
U7PXBZtFrZquBngEQNvuBm0EV/37aXVXpQNJoTmKp0AeCAragrrmiesS+EQPwCbJ55h+czkn6F9H
9z/dwFRJAi/Ws3lGgFXo+Sw5ZmDFPdX704nsKyzHh6B/ZaLEYHS4G5cyKLZnD7M8gXvh9UnUBFGQ
KLWCLhMQMk+RiQ0uruhvqc0UNBzfc1gD+TYH7GxtQen/tVeC4XK8ydzKyAp7/7SFyA8R7ZwPutco
QvgNeBAGS/wxxdTMmV0T9jAzV3oSy/js67QiTeqqjJ4kHglbePLdGkD+KMZW8lIFvEl5Px0TbW5j
xykArsSyqRKDXuoRZDOYRNy3NV+eZWYY7jtyabYoKen68/5PM7R8jTYFW8OPh/Jv+8Ys9M334DbB
n/Bg/UTSGhC6ZLDM//L06mEtJ9kL8DsUpFSEZzdJucBwCcjKkJez5jG0mB3mKhAqUj61T+s+sAEw
FgNELD4S0nC4NHl/volv9knJjN4rKPD4jv8mUu9E4oZf9/XbRwv2Jf1UVwDka4WME7s/AfzAshRc
ONGqhU/h6FPToeQF66JdeasdFnIjsX4LloiP4AnSHvF0/IOSwdfsexZm8UlclDwVDie/lpomQw2O
onDYDKmiVvX279tj5RqbHH1/kfwlRgVUdmbDO7MpOeikb9Nn4Uy23lLcYwfJoA/uxIuXu16p4gqm
dCGU4eRpOqRkSO+YOdtjRGt2rO/sRcIv02rJIopz8wziqwUnRODcZRlV2zZZPbgK79+PUp5xI0tJ
SjA0HefhbTXC0SYLjL2kiSR0smPuf3ybWtzLZ005Iq0u1bs13wwyU0uQVPKiGVAZLtq1XF8JYGTb
kFu/K6RHC3EOJadQyxaqxwG4nnYdq7SJ76OFpM7xAG2679pu0/vJs79uW4Hl8tMQJISdYrpmdVjp
wJ7ht+9ZPr0PWOsBP5ZFMt5dautmkx1NJ6RSTma1zPLMgmWKZAUvzrCDU1gcc4S5sJ+pj1NpqJ/b
ZA+NgkEJCdwTNLXsC6DumKOV1RKcqZi9IjZ2+UIY6rExvILFTzDKWpFcE2WK+b9oq8a6PLew14wb
XhQZOhPVGIuPXL1dqK+TyqqX5sfbaLLeDThvCr+mWF0ZC1t004BhR8Kb64VJ96808pV3wxA4IqTi
YXF046d1Nvt7Q462ueIqiymAfDRpGyOl5T2QO/64KOX/Pyat25P9Z4aiJk0j7GX/TeO6voHdskDD
z0FZM9Cr2rs54EkrjNewAwqooZ31Gn/HWzBGkA46HdPruqnFoPp6io0eKGZGN9Li20yLmesJqMp0
6gTDS7wXtpdmCpvVfKx4QeuYotB0RqjtQpeqmhTvG1v/55Ypq0ZirKsL6BIJev0DAtO8YCKFX2q4
D45Bk/0ciJ/HKTnmacrBqYDfw5oNSIWHNfZR+szUDvFW5ms0QcNT8KPl/44RXWtI3Zs2dGdYRBEt
JVV3E49RCbCvLUs8F64CCy9n56FldC389V2whJk4zIpJA2uzuIXI/ZaguMSMnB53Md0P0Js32gkk
sSPgElZjAI8TBYpmsZhUm0EBEgRC9wwoUy+IrLeQ8U2f23h2jBDLC2xCLRP4Wbvwj2/qAgKihoVf
tmhpFwET8hArS24plUCj+2Ld3rR/xpisU0AoiBAcUuYSgUec+BugZL6Lk+/euHJ3Lrd/kYcW6Qb6
wXnO1JL1cGrrPcZBszaAdYj/qDm2yLzUaHeT2gDZ9b3FcdbeOS9NfLOX9yjL8jYnnoV/YtnwIiLl
iS3zSxG1GcvNCWyd7su6BO6c0O44BGEy6TwPqRNQt7Y2DwJD1Pr6lOKNtO5HMuM+nraQeyiw7PTB
HO7Tbg2+X5cVU+iL4i/jSx/vR/UySimNCacMH53syk5NqPnHZzw4IXG99J7hStyo9PE4h/zf+hSC
w4Mwnvhasuq89X6/pS02azN4aKtIyGNtNIV7cjBcifD9da04wwYMmRrh0Ah6LORhgfLla6qDhLiV
0cbC9iFIrpLw0+clefTFvbulnIPaD3inGk+GghN4A3nPvaebChBptxZAp1DrU/rzT0qW02t2fF6O
bzUA9A0aUHyQQnMwblQg4K94lqMiSZctp/sKERByWBKb0M6fTm1lam5lRvtVpcUrzI4wd9SF6sDe
yb9yZb6qTrzjfPRmE8q5uv7Isl9lFNGUam60OmE518ClBj/TyOorx2PuI57xhQFGXZ12GPFT4fbG
XBYptFMbWYNn0tjHH4S2SOCqtTybAMMENS6dmPjCF18a1nAg5+MOmjrii0QxPBqZHsBXPngUvd4n
zF+jIpcU8YQoQxaeaF526F1mS97xK6jH/RBrQfSUI1OW17uX7/BRJHWvcu+JPO8gzObqvvSmyqcG
VYGXp42d4uqblZeL9t2gjwQJb6EE2JyYs6Fux9nIgGkzozqpFblo45hqcVrpXPwEupRB4WlA7jrp
FpbR3+SXG/Ip0TOetRhCgHrmjgq0Y73xqOL5e+lCAHozt9bKiNqaZiXmmPpsj++bLU+CNvxmRKXT
+IayOgwtqWa+KcbXCGCF3Y6Ur59afjQyyNuaO9oWqs9lS5WcdOxSJFJAV6V275EDfL0r7ieyev23
5SdTHpWIh6VltSJp5seWBznpO+7pcP99jZChrfZ5F6EyFtySyGe1Qb1h1gYLgDkdnnR2RlM5u/am
0PIUFY+s+0AAFV+04j0tqUAM+IJnAKu3XQftDtLpUH+r9gPjTItxjozJh/4/Rld9hPs6zWCtDK22
OOsYhfAxtM5mqARFalq2ncyyB05Mom5seM1sQe+maT2pIoVEqNwkNG1K9ruUXsBHUFOrjQCAx1Hp
0jJOPstvuIvUy2cS/1K7CTWGmi0hgwtjzYj6jBS1VmRfQGL970Iuwahd81NSQ31oRHEpcUGJQpNZ
Y7CFK6ZiOgGGSY0aYn47ZwzQRGEjK5UpLn2kuvbqX8F/wNkh2PYHz5ZEgAsvZdkHx6vQYFZMRNHC
UIU+5THkWGCJ1zhvQGEKBWL261zlh266S9la50GnAbhqIKUrvdDioEI81WobdilAQZcPEKjU4Q71
r7mc8jt2incpBhQsPToT58QrbTWm6Ct2lCKDAmEWT/GXlL+JiHhhQ6bbj1Yt+fCW4voX3y9shBUQ
lDYIkhr7berJZ+HV4Md5fzzDSss7FocqpExL2daDjanhY/1LW9BDCIoQdvEswtrCjAnvNJz4H0t7
GFZrlaYZVQST77n148T4TNcEUC57PMlFKzSv0+BdgIq3oztelxTIqZEBS8s45ZIBEnbnubOl8Ymr
rB5JGHUFHyMH7cdl2/co3uvniyFKRQUehWdmcQoToh+72iCBZ3mdJTY2F0LjO5pUWjYhNsh5zJ8y
Qg9SKqiETYZzyzpc5sbNgMth7r1+JnQG5voXzqstyJWw0lCP+gx+6BqT1g38U1R/wm6PIeThC9yT
lfCzCevL/iZPY/RwPXkdSFUTH5lELN9xK7hpAuIH4MZIEWpNwRD4grAVy87RCeHLLbYKgSLzWJ98
e3mtFRclSpv6KNhwS/AToETGT8tjnwqzR2YylAb9tmDETVmrYpZiy5mYlwgNMhxiTTfEByZD/b/T
ir5gjcj58J9ru1gLHNijcyZom6jWMeVvMdTUSZdaLlBYLdtzLmqzEt0Ue9locX+Xzu/iG6sqZ3IT
FSEB91G2TJO1OClYSQrvoSsose5zXHDUj0XpRuQ8bqmF1RFN/X/yOoT1BYmhKtKXU4E+QBnW9fGv
PFeGixK0Cz191YfsmZcve4Bp/MeUCrQ+te2Hi+vjK74EOV1bMmCVnAyCDwcc/HvKwNgpLVIMevFH
02iX/J7W+uCvI3B+/3xYhZG4miq4o5zy6WiLSFhL+35tLDVhoFRldKp5ikNP99uw60QGvS0e5DR+
Iq3MlVbfEhV+GOTU8aO7TQN3ouzi1q7tMT7e1CxInLClEsPHcDccccva2lOLIDkqPpa1UK72vIGH
uORkj2+xTGKxXHHVXoAegeMd5pdwY4i2duxPiMuz+81oMV5qs5yJt3dJD5qCR15FL/3wgnN143FD
JYqcpiUOkUmnaU3Qa/jXcaxll7U72Z2L0H9TvXMv03AHKmr9wVAc+w7Ty8+vPnxV0va7mKbzcmRA
OIUPj0HV4209owOtdRZXncRYflfrGGpIpRWxFNBABbjvkLeJSM9OzNXZdKkzFtzFMcrNy2EyhR/5
OdnzwLcAKeY+sIvm5jB2RZz3VxvdBdulu5G8OAgYNcfnSx6wy64hpmij7vON3fLkS2quKD8VC1Ff
5Y0weYeCMi0IZkcEMDVS1McXz6k/omOwn0bcT7nfoX123wuIqK5axAoINr1mWrtZpPB2XaJQWjHz
PGR0vMHIFFd67D4uEVXWi06WYCpCG/tgkehZooAsThgRpe5YXo25YWveq1qXH2Cp6NfJF73GEXs1
+AXO9AyQJbc12EN4dprL7xPrIPK/Rm6iTa8G7t1JprDmEVksFn7XuJCitb6rdqeFpvJtdy/dG7Jq
hVUlV+j66isqEfNu/PxX8Ef/UxUvcvdEHEGdCGH6mXT/aTGTihc1eIUsyqfW+hnWqRJHVNB3VxS0
WHEYTcLppvQ0x3ugLCQ0Gbs8o9D8k20EVxz/4AIQDOwVD+jdZKl3ADpXmvCzrB0Pt9M3vrdlPeHW
fHsPtT4xh+bq7BDz+O0dLIlc7eEz0qM/PFuzKcHRMT/+zWQDs4DlqXaNzV9qih9glfW54HlSVyHt
9TsbS6o7ya5tcGAwWavbbBEDoxDcCSCkw3eNOpOehwTjxChqXxagm8OdDZ80q/coEApgoIIVvtzZ
xNRcC35szCxCiUW2GLqo4VMKkdIbPa13hzofTTg3/wCj8SlTkxOUNaNY5B7g7Ly+/i404RW3vWzN
ViFWe4XgKlXnbqT+S3yM7/ixRpibx78FJaN+Z4O6wPlQEXi88iUhFgsHcXBugHhO+13f8GPU4h+D
8nAX7R6NCWKBbjyxZWPcajRp15oBPNYRV1hH3gy2JEzGcLfBt7G4fRL1coa2aqvc7pHreP9Td+qM
dTPUcRUeusSUvh7780tvMh6sxCWRtR8HBIuPzPHJiaOzqBRSYUpCOocOmxDglTs4ENMA+KTC+XWM
z0/CRs3icjQGvfE8TG+rhPfKBJg4+2c94Ex0RMZDqRoLjBF4LCvJsJqGw64SBPQGklrgZ4WpJZos
3tbuUPKLQWAv4FonQTL1J3upkLzkaTZHwzlIvNw1+3ZbH/vWefOZIgY7eTqfXvgQ4vz/Wyogq7MV
ghuedoEurc0KBEvRT+zvmIw/jLR61zNgE/IJbbQEd9YwdNHQRIk6W/m3z5euhMmpDo8nXLdw/6n6
CZOIHaQgLKtxsii1OdZX9faL62a97jlUdfCyXauRPwBWY2MEkpSj4cgw09blBQRlfKfyJrEDTcnA
wdnMoUZAlFbK68wjS5GC7QCfzuUxkvhlNDAIKmgmV1mgLgzN34kchsdWIwtDnvS91z6NmnSvU2T3
q6gfbxMuevNinWLpnUjs7hlJNvywSF5XHGzZxzqe5L0s4ICPJZvrKe+nJhRv+NFlVAxbb0yb4w6d
EejryRRrgL53KcTEdTpHbdylBLSKfJPofLdERoI/bhbkXOgc8Wtu2WdyvNzpBkV9sWxBDeX8rGyX
52vr0ZXg1tyc7v3GIc8CpBhdpzCP807LII0jx1ijlLycUcTbJF37o/c6/lQpevFglENJv+75M9DA
msYTGNjkYxo9GJwp7sQigVaPv2/fATjy8ImDnJc3SXN0xM10T5Qku/MGjx3m2Sr6ygVExzwsf0qI
O+hOZEpyEsHdP4sL5p8+K0IKRXegvCilG1IinsxAXfoKtzrxs2ILDVO9r309sK1IkCDl1j78IyVm
92xHUUGXp+FcoBraN/ojPMZAlX/1C8/3aj6tHeZ0enCd/ifma3i2CbmVdRexE4+mbLkBXKuKq83D
5aN7QHxPWcn+va3uGTQUKjKQfF7ggdXHTSMFCQtGdDkqeUtRSyvy1dyUyDvCyiEly5sDfIlpanpV
ZWAi/5t7SDml7lWHINm+x+exq4fq9zBYDYjZ3gpEL5iawJNbcq6O+yoYkg9cp7TtSRcA0JJHzkvn
ud0jisKjiQKcjq/BoxOA1WhVFxj7hcqaWrMgq+P6+EdTKygcq50dTvSUfLuFOUrzEEuK26CjFo9d
bX1uVgAId4nTkE106GGxAPXpjH5qtRhyMiFLyCm6f5BHeopAIiidTNfa7RJWyzEQCd4+Lta1/Vs9
XaR2ZZu91XkuKOlpzMt56nqNktzhLtE2kRHMVxbAJMdciMWBvNMs9E4IOmgaR2CRKb/cTbQneNJD
pjhenxe4bTTxdorD+8sZ/iziB8qWuBzJIuz2mzVbgQekLPnrven5Vm7UzpaIbLBUcnMIEslX15Dm
/p8qnJTvHcAYzrAT1gQMoeFvj+seOxEZAbgIXmw++VE72r0iYLjCq9ws36gK/wxuvelFLOiLBIKt
jKkd6r6WDuv7k2+MvkLbbh7o49DKrzmGL9j0Ox3HSN2vvGMK7x4rsaxz9pbPK9Z3UZeQF76cdPck
HWc/NiUd73huufPD7+yMBRvo74I+D7+sAk3H+ksHyMdRns7TcgmfnlumDt3YXdK12k1Y4h/GcKs4
Mty+rdxEw91kHsgv4K4rhjOoQFNXFbV2JS7sT/YUbX5a/CDkeJdeN0qdUAZy/GAXZnSdSmnBXNCz
iXdNiiC1xI9FAycMr7YAuw+h3AH+YZL6TVnDjVJfxSVfdebARmA9pD5v6VkXWKY58QuefeoaLCey
4IPrcqwr7vgLB1aowNSXMPsYFYHTsHfmHSI+241gcFgqvBrpxWjxrYOxmvcSGVVRFlj41lHXF5SV
WVy9ac3UX22Ymg3UCWK8xgTPqlw1ccG3L/eKXCJNV+xKvath5LeuX58R9yTMF4gs3WbuColDYr9H
cYVQqFqzdEP3lfkW/9Vt0JYjO4dM/84zuJUE4laSIIw9IPE1zDcdQtcQvCY8i02MEXdvTr+VAUIX
Ji4Txao6fwNlKhCtm7AH1EUjWzAHiktHfAA2kDe7HHM8u0bu/2Dilb8RGrESICRFcWMFuvsmGiP+
doILdVT/L49mWDDcEVk59zyBnikTbnCPP0sMio46+dzPqssCmY6qM4IXoyXk+EZdzjWAHDkt3Fvu
hydV9JY/oYuUd308WTFaOrDHYJ35G4g9BSeoEq7mhP67MQh1Y1+yn5ajU6U1knu/Tom+xS2hoO0e
Yte+Whit2YMrv9QXHg6m5JciBqigZRBUntCzXJ7S5z8/LBbyfrb7BIpRJXgWCJJOPeZwf+n9mz6j
zA6kB5lupenwvlbtWRrVE5idlBS7nN/fFqNvnFYDaajMYU+D1Qi0NCXWwUC5Ev8X0+PUdJy6JRnm
hinvhlHs4AUsdPb3qIT7FHf9smUJdaFSqiZXiPcPiHRZRykDeNgkF4vbDsKE/wV2UDaq/mLPS9AJ
VqsQX90GOvghZ3qOywlI9CodAeW9GRjq7XpjZ7WbGjfUONBY5xSHMqFOsC1v57XXUNrOje7TPxOu
sQ3vhdTzIqLsrWPEluVXZt2KHvR8Bg0lnGXxUg0G8pYldQ+QRVc76HLsEazINwWMBVB3ifPMw6K/
NNZhYlvY1ixlAnCBwLrG/1WkTu/jf5nNuq9r5B2DMxfrQhrixATD5bPh/EXRQDsvT1FO+WeoG8H1
1rYp4ZSEUKDZY6yJ/OMWlSeLfUivJjoemA4V+GnclQ6A7YeGb4dJ2D5ElDIFD/Z7JD/bhPVBcJkm
lBroVaavPHLO1BZ2Hv3E7ZpSyelgWiFOozZCLm9TQ3X7xpPD71WhEoLV+mrRFtzEI9deIr1p/rP0
ConTUxBh57ofqyNJ3BLZ0OewDbgbRSxM6/fvDb9fG4/sjSsq1hxu1ORdyffC2IP2WCM3E7BjZVcN
pVuN/AUG8omzdUJtMEu7ykUeRTIsMVceDKBZNoabm29M3Lz5rFFuXtuHUhp26LHmSc21y1xtVTWC
uyvfW/fMHqA6hIeZMuneFiYocrxGcfMPTd4B5AjxS7pgGUuZJyWVKfozZJrmh+6Or1Cl5K/MY/e7
Mi4CXPminUFzyDsTpVTOyz9za2eYL33p74a6MrxqD5ZNt77ILAICSLDddcoP5fs6EsbcyLwsLCYo
ioORP9BZS5qMWUC5j2VclfkVG/RE4lG2uekXgQcVNU6/LqV19MIBXAb5Z5weaDECu1LW6I5H0rEs
2CXdvarcI8Vm9Q/wDbeYpAS0EpP17uYRMCR56Y3pTF2eCpShUM4e/OXrg41LcYpmyA3ykA/ZE6BS
+UfA9nUL9n7+IntgJuC62cDiINa116E6R4DkWVhc9ep0C8FxT0qq+MgcwM+sHHlJrGtL6h2Ra/a7
euVNDiGKbPoH5pEZiJ2z37cu+Rp3oU7TncVxjZeW25fK0k/ezuTEjscay1plHupdjL3s1F6t1du8
yMpQV7YBV3uyxpw510fD6BXJ9uR9ii/4wRl/duhxYikaktCSgOMIxo6E8OmgPJgPfdBei/kk9qYP
cwnMw159w3JSM6d9dV57jRPGuG7taRrzZ491Ez6Q2S47uBjKXdcRbca8GXiUI5C4HPgggycA6Klw
1PaNexPpqHJiqLxO1BRn6uxTzmBayztnfGPm5EqSujsTrslTewWpC/Clx65JfIMv1VTPv+C/mzIy
QfYeEH4nmY3ZrSXgA+L+YJXyr2Xa0LXJtAHF1AEGS9gAFfOgUHLrRMPmXu/uhQ+VIkMzkFzM/lsn
9aIaxp6sCSb9Yr1TPBp2doRYRt+WiCBG4N3QWe5ZOY1uHClRFx54JJjQuDih+cQ8jQjpSt8NTVGV
QutP3l0UCKi3d96nWlW8WhDHv5+FOQMzd6yENO+kSzqITqP5MjJbYbZrY/kGLp1KWaTpkAIEHHqt
ns/igu1wZ0XcIAyMyFObDQMaUsPNnHulW8No/eaAk9+oNrKk9rMdDqWprSsW/mjwaDGbvvvNq+yQ
SKDBJvyYbLd1VOEWYyxkdh/2Q9aSYLgp+WvURV0DDjOb0zM7vmEOEPDCIHEtYpU4nH7njjbD0+Xd
MCXSwQXvZn/7Lk1K1Pi66xMacWhxK7BPa37sHdz9jtInunRLVZIYHvrx1uDZg69cI1eHNU+gcbg7
GfPB3EMr/idggbjdwzUlYPqDDanLITiOmQOvTz8Fa6ATefgIx+IIwK/d+paH+MKkI5lNxWyNPNdH
drmqQpCqZqhJSb/IfHTPgLC9j50J7AvvOyUFDHSXcq1whhNXJy4qI7MCcZ4y340Yhcs0RbWFFaXk
ecykEKJUiD6YIrwe3tz32KRhmD2SqzqS/VUZtY1EUV5z0AJw5rMrGvRoAM2e5oeygXeGZaf7okD9
tg3LZ3SGnjSMu8kvMISnxCjInwOV//ZM0Vc81QIFrgbBn/vCrpL9FSlO/ES1mQKr+/UmVpJZcwNz
pNcMVi2cUsSzLcrVLZCWM+R8l8R5M6rMloV92g70CyMr1V+H9AfLODUuO+EgO1r27G8ZQuiPvxU+
QzLGT0iWhcxMXQ71N0oGk2zxq9T6D8XZ7ILBG+kAhkNSVB4QKsp5G3S5yqlOvwutlc8uDBdacE2t
zwmZ+fUvG5gGtvBrkvG9JW6QjypapnBc+E4+7gHKYaL9P06kxzVIWtAsRK+fLdFvNONh14u8m7a/
O1vGVntlbLvzjVB75Qd7Su3J8K5zq4Git61u9QPjKQVZeXwakF485sjT8pPuxaLa2xOsv7cWLE3X
/GUAbKlKBk6Pf7J7fGTla3DZLTJ8kQlSZo/AZUuD7YrWkKa0g09pqRZMJq3N/JSEAIAvLox8VU1H
oT3Vx9T0N//WYgRUFe2iRQCp+cNwsLeT+zAtS5woC0hfHE3Vk9pB4zmpPhXhMC7XqtIu8f0CZYWt
fw3LrGyMSGqkjCgueDRHEp0IiMgSGZOK/pT3MdN15wkTvNwg0ZGBJXGCVMpBwO2WyNll9fAFnq8d
zqUqEbLxXiPawwb7wRHjIHs/hffvyevZLahvlKoJU2JasPwdMLY84HwRk+smprICddDacQpLgW/1
oSVSSrJ/CmsDxD5k+9ARs+t4wmPAdYB7PUn9cZNDXDTeFwCBLdnuho6pRk9gI7DShMrKGnNMNUOo
rNNjS+KweA+2i1gnv9c7Ge+LJhwRs8TLl0VC4iSWt0T2ovK7xKvp8nkTw/mFNq/0jc3fTaiFKH++
CZ5QOnP0u2gNmM/ihaXWzO6J6Rx78+xpq9GnchrxyCLvV++3+zMFwwvK2Ybo6GolW2eAl7AI4gmB
fascoCRxLjoBdIKH3xl6BAR+8cUirmlMZ90NdPJMMZJnUMXwkMMSZkzKQ9bVc8ganKN9PTRfAAie
b8reDBxi7L0TfaMO5jaO4UGRHOw1o5FF4Fkje1BE6YdlJEsGIpiNiljf9pWhg3KV9ZxQvhqfywIZ
tEb8F8eXFKJn6SGvf8h9Jmk+NtlNss4ieMWA9B7aiwR4y4BC7O/hqUIvnhjLVlLRuCUSWtIBuw9S
43W85qSZA+u7TxHf0VbI5zqYIV7g2y9dpvmcPWAy0g2KaHcooNto3LLyo7gxSK1DS9cXGpnkfGFA
rgPFC46/gMyWiutbpw7gUVD5FGinXf4cdz+dsHH2/qXbxWfCKejfZqBXYTcrmJl+b3MKe7cEUFYD
UiXe9UgdIt+NwmSXmFvz5W3iHO0XLm0m+hfO+fWk0OXzO21IruPGKX/2lLtghLatKqz+VBfe9G9g
FoAsAZy/pMe3aB0D1HcpHEYAnKzSXL2392RCmL75MWp7G+wSHFZysSdc9KMX1A/I8aDWc1xOKdHM
R9agTVy8FkJJD2sMVh/wd5GLLBSZhdSBNaJl42FTTB/Gajq7VHK734aPX+lVzElsGbI5EsvWxfzT
B+yQrt13BV9yWFxcRthzV0Rs/nvKs+exEX0s0KSXY46Hp6pAFpPV+KJzLi/NIVbZ80eKuR1imX23
xNytd4OACoWTA/GYOpzotD9i1XkK6BtvwyBLkgRhlCAbFov8n50joqA3yvJDgkJ6i82NiTHwxjBA
j1gNbLlNXRe4EAOznYBG+NLShpT/XGWe/p2DBZvcQJCYtK1xocgajACbR+KIpnsvSQ5jBdtme96N
ra60q4msfs+AGtfCjW3jbnvO49Wk7j6n3NdUniynKP884nWhERop3TKwKlHD3UzerSI49vDBueqw
snr9VjZQwGUDE9gc6z2eUT4k0XgvQZw4gjNe53iH36K+tlJWmwkby8oUnzU3/B+uHbtcBjhRZ2EM
H8HiQMZQmFr+SKZqF4IROCxxJZE/i0JPhRjvE5ffIhdIw1gpFzpQ0kFGNLSdZ6xUA2FO8QCasozw
n0MHWYrPKowOMZdS1Kx6TPqZV3JCXHonkD3/ee3g0/o2QFtVHeqBEfHiD/rbDOpGTWtoThZQeS8Q
zlzaUOqM4DXZP7W1h+YG44+9UvSO4UvUEweFWq25zZVzIp9C22xbHInZEYOnfBXxI1sHrlw4eJfk
AJhSpAlKM6o5CVO1wFIYdTSoMfLq3efOpFWtRfVWz6yJNLbekPFcNXWNCKxSENy1gSWB9aje6y6Q
4wCWp1Xf1czXnitY7uOUZPTZ4sABUIcb3yc1FcX4nlyLh4tkplKYj2UWo1yHdIsfhtBVaERHlUlM
LEe5RXA0aWSG0+HS0qn8qSkDGNYwPCfBYjjqFpNArmkxUbzeSngSrgJoIFRd7f1xifsY4zZwEDOc
9VhOhNWwd5bP61cCKHR5AEKAf14SKBZyG0Q7EaKBbDR8CY2ggsOmgkVVbgiFlHToUkJFq70fZYmD
KtQqZ/3/dvzR8H4WnWJkXaW8DZj4ncEWytccK40m2hr4t+bMoFGs5H8C02LqFKZqNbZmKcpwuMRW
oXHLJ8MxywrEi/PTcnAOAE1vUolEIVu04sFh0fOvHKfC/+3+TWP0XSykWByFBlKXKwvry4rwZ7G5
Ea9Lq4xkH+oc8xzWuQsL3OoNmniDBSB5+Y7SvctpMWpm84zTKbJxevR/oRpc0V0xa+AvHqyaoL/6
XmCoLZQ+3uPQzi+cexBCllhR2TAw8DOkXe3Ge5g3IIl6R5NybYhnxY+I+3WV/wvywJJhiLYZgjTu
JZsa//qhCvOIYc7HCXNi7JbltbKSNetcb+vz3vca+p6LpIyHECl50LQJxIy6EsKvjVxKbsBmoh5d
OF+ZMKajH4h4RITRIECAPfaiLeeu5u6Yq3rDdbWA0bgdnKR3o5CLio7loVfSt6U6NnJVmviHYw77
Wpoai2DeHAporn3iofh+zMn7L6x+iwd8n8OISzASrmHIPo+x4+M51WragisocgxlRNwnYURl2Y6S
cZ6X8Rc7/Efwt38AibFY3D9E4jrS59a1KkQnLf1TW/feTrd+0H5tKQ8QvwYO2stDPRjUjaSFqc6D
fP17T0TmDihFNLpIxJQcw4yvzig5iSxBQeiAmBb3Rj7IRCnxx3PmBlzofBtpfJlAcXZDBYqlyUjC
g8fpwFKNk4ya5vvsNGU5lLa8Pc+2knmXsve+UjTXTs9l+AG93JTvK5DngzEnw/x+9LebNUpwC+wc
1KhGVuh6h1HnWL/4WSIxktrMaPZWhQRiagxJtrws2vPhgO0Fv/7O5q62bTANSrOUzqXiJoXZK/2I
pOMxfK8h0HldMo0k3eKeSUuIiNbZmQCzS5NFcTOIZepE4NW8bvF5ofZhOv+mlmtTk413PEYFlCrF
EKVseInV66qafnx9uzIxV9YK3EJJNIuAbWTchdN4Cygn1daYLVrWy+217So15lomuLoszYITKYgb
qSokr7a4N0gZBOXmldRXyFqjoABuyg5wL4hGoJtyyRJH8FGl7smz6+1R6fT6w4F6dbJYFLpxg3/z
zSxoe33JH/hV6swXRx0kKgDnYyCFXTOa7Ms2Pp2Gwz9s2oPQPKDUrCLS8ELa0XtRGt7U7G6fHJ4h
MrQWXXoK1+ZJga4yjU1f7OEsi2vX+o/lOj52Q05EB9/kQH9BmUMvUgJiEBBTO0YMDkzxefgiKpPX
UBCs1tBtvOJ696EUobEhb0f6VONjXig1aae4ggxvgR6RPODl9UKTxOjV9GndP0vM4wHDEJ5abW7R
2QpkyEYd12idlfv4ekyZqZrev/guddhjJWGptamWTe+M0D7mIUBVDFYea6GREZtUtGKazjmIIO0G
G5KY7G8ZW4BLQcaoKRvvr5q6YbDs/blYmHZCM7Fqd2WpENwM+escOSWjjtllcWUCkh52VtGlPHH/
LT5wyzOeQl+zDyC6xSmqkec5X541PCzeRziTeXcrKEqVBm6YcQ1qZU7rvqajPYtYg8qL7OjcouCQ
YNWdQ9o2uPlYCcSMfmDepDuGUFhGtYlQFZTBkZQVmoRcgdkmKLU15wZy1KtRklkH7eMeges/R7nf
VR/sGSRdShP7igM6+iqjOQCP9njTR+N2tvyPEOKv32+/sGOgRjputkCltrg1qBGp5FRqk1S2t1Hz
CQb1nNdCnCcMCnviwtTwlUPpfKLpGQUxLBmyj2Fpw7jylXmxXffu6BnlgLAk3HuI2l+67Wa+9tO1
K2OCFOu3MNo6xyYWOcWgg34HWbf1xjlcpla9Aiysm/s34ttIqvSzYaAF5dDexQnJW5OCLZ+L5bId
Dr7SfMLHGIKe83PumfkwPNq4XpsF9f3+P8Hc0jj3jBnHbKutq6oxTxddTj8ghi3eaCjHcTqFL+3w
wKEkt/2FiEK+Sc5QvGX1flA8w6a+1EU40kE5H9xu+zqulLbwLDx77OuT9XVv5j6EoBb1EgD4qcL7
Pn3Dhcs0Xi7AvaUZl8bRgYG5ocdyBcNPrQA6Mvx8wEDvFC4wJWFfSNbEkZSpQxEV6dzXDRhMku9q
5bX+64YVotQpubXGPnjUf5ULarwUFCMNXfs06pSdKW8eXdFD+8coPhDPuRIdb+RsFgV7x8Zi/BVV
pFbKX/BUYIDLkoCP5HV/QhIH4V7LsTwDsdyWopnQLlSDZkJAWqoR9KMpNJNOtUccbapoVcvif4o2
Cwc0LEgTvyUr7OmBS4420V2ux0GU79rERa4Mm5xvrWEzTyQvk2JzdYqIP+6F3RVSMT5bPJbL3GVi
NEaaaxoGxPMpkQO6fjE3M4/xJBxQfOHK2OxS8lbvK2nHrBbI1zBovxmsSaQWrrv4e2SzW/gS0So7
QAR2lGN1gUwn78GF07WLXK5eTttsooaMBCwFouu+H+fOAv+oAz1xug6PktKkr5QExgEMc+f27OAi
7AgoS9Rf3tO9BVfuNnSlqPsdjo8mg/jhNYN9Ss6Ezzs6LCd1MEw4GjxOWl+2aly4GeIH1GgmLmet
9/1UZl3nAna1DXr6qc6cfBlAvqZzlEpCwr3iDEbfQUXjiDwi1HEqE5MsN09Naoc/WyFJpEtJu/Vg
5M7/MCIWonNDZkhghlPSkrjlan9pMWq4tDSYR6MxY08ak1jvTVEQ23a2Diz2pzlmv8W/H+xRjHUW
u6AgT1XNi81VZ4MWrgaZP7pwh/i0G1Ay8zI8JFoe6f5RFtuVpQJ5rfH57qnE+jefY+zvYKTq5rk4
IJcoZNA93IxrzERF/B4K+uzMR6rfDmPFqU4E8/tVGbcWaXADLsND+rKqCh86hEji0Y9eU7N4kPYU
YlH6jmUazdQ+5nSympdUEfpJrPqY3sN1Sy18oAfrBS4HeiqIgnMONOT+LYMfy1HEApFFypfxlZgV
4FQFyVoAo+cfqkG+8nnsSfvXGTpK0Xq5XAC/tE0VA5Ek9AHAstEKrWR9pa5ze8x7QfaRwbQsGA48
ZDwx2O8vEQ2S+QDOaO4K7zj1/Dcp5rgXMgbCrhVKx8/aNOzSieRiHzv3S1EBAFh7ArfxSLMWuUKd
W2j9JP7btq+DcptaLjwpnMttgbVvg+CKrmZHq9fPNV/RufdBnFdvEjZHlL9LX6O38uptdIDwTclW
kfyOu6EB3dADcv735ALP5F8KNDNnrqJbpdXavGuBmCzcg/6A/8AB6/+bqgnE/Yt+yY2KBl0BFDfF
w1PWBsghI3aAiBumKn3QDWIWD46aSRfq13/GIoeEE+XhXz0Olqn4AI4uovu5RUIpCi25/2wgUd1J
wKY/Bq5PwkAWpJE5iKzEOwLjKRdzXgjoMwmCCfSqxgV0Q3bh7H3h7EFGdgZ5BB2x/bon38+RJH2e
Ts8gpSCr94iylbWXcPzMYpBzpsavJdL9WJ0gg6XrrBVyWLaz5raWKgi7Vpm65zSdZts8FngWwfHn
VMk65UZjD3FVWl948Us/h0zbwtTdX0qOwLfzQPfu5aHc9oj1jtAoi0eQxTj3F0V12a3+jrEhn+x3
3EfGFvHJABDiN4ut3wRXJbxtRPT5FMD9Y+iCso/D2J7KKx9N1UJAN9H0I+FiF/pdfzUZhSxj0XcT
edsJnKFyQ1jo/CVT1RzpTOIgBABJHfsAqRUBK3sWZ4ASfsZOkWsnnCOD54XzNZfAk2J9c0w/oVI5
4I0d3w9xu5bIp0mBjIWqLMGT1GBBXYKjjAN1uS8Ui/c1TtooUrHBoLkggna2EuBYPhaKx24gApQx
RDuvrqPUqnbejsGaUKCYzrQ42CH7IxqGXB4/byIRrPPZZZLkj/bDeics/Vzh7/RIy8KG0Uze4WsA
8oIPDLbURFgnHUzGcJhNsixt42J6P57CTXGRqOkUXw83P8gjg4ybUGRqhUiJY8EGEp+61rCPgPi/
poXxSSUSkF5Kv2/KLlggnjietmZYc48D9DutDJm16Wk+uMquGcY2It8ykrzsK7bI94yQHw8jLU0C
PTN3yia/GUvBlM+gRCJ1Flo81fVx0tQRFQdlzG7BgHp6LajjqdGVcDJZ2iYe64gbrMhNIe6p6mQL
8FbydHRdjDNaTJGyPnnnIjdPcMj66NW5c3oAYsdtgOZedasGJ7LkDqYzD3ar6k1/P4Tw+LJgvwK7
psqqpvf6vtMZ0nTbM6ia9QMwVx2XVcjVydIXLXcx+aPpSZeMw2HBa4ZaTwHPCCb34WKTGCubxHtb
sbkmKPfMpr59jLT2loty1Q/Gxmm5KSmZD6rHxtOAN9JQuMTfBdnwQaDsJJ7SpTQSwC2PUdTzkzo/
w+36Hg1FS4S6z4hBmpvvCkx6P7tUYLzeGDMwkxEigdfrtTNAhB6fpC5hnB9E5XpW0f+GRs78xtbA
dtVybvtAAcYTWnY7x3+saIl7ruAcbH34u2/nNPAKl+rsAYKvgKDrhs5Qj6sfi1dLGetdZKRtMuA+
Iqxe2HtZlMxAN6qo5g6oMT8pv6K5+1kg1au78fHfG9zFX97jnAnu/L78C9T26uQKE2Po+Y9h9yoB
7tSQ73USV/hMzTLUbEi3Q+6Q5iQnrdrI7lhtA2wB3P3xKgnDvZSbecv7VYi9o0K969yfkGqf0hpv
shOzX0h+NwsvwZVD61woQL0L4uzJfSL5Hx/+vRz4N91ktGaaZVvCec84tn0A6PBD1cZajVNo/KOn
4h/Mu12E8+2HORu+rbo9H42inUYTuquoEqF8im4+A36y6SpFiS/7dKeLgyo02Mi7QdHW/agYTEHO
WswhtnNauDo4xF6MVVWyfkVLYcpmg9JW0ZVwMtS8mZcC2s6WyJbwiEDKrPDVX1J/EKOEZ8IJzYX7
puY85a7VYZAA7SEXDk/Dxcc76Cn26XfCojn2jprXSx0MbVCazOG7fZLb9jmK30h0DrU30YnhJp0g
kabEhuv/ptmh8pM38eH25jGY753FW507fAm+mhsjB43iMj3BOaHqIbFTUO5hHANp0KkPCOPDFCDA
ikJqXJWIerVV9U3NT3z1qpS1nttmFZIONjoiU/nBwm08O4l7RLEiUCZ/Dvj89XXY4BK44IlJFxXg
wTvmSJTNgXqcIZ+e9iSWBl1vJKjV87pIQs4YDIxDkueLf608FAa2YGicYq6OWL3H6wWiB1QhQSxH
RnxX4Fc7C+zrTYfEGUS2oRG+KSfGQgrHsHDFdqddIojdeSZinwJQ3ds4l1mdp2S/jkiJXePKnwFt
1hDfSiQszTVf/4WLrKsiWMLkj6oL0vJSuZ5Mmkh+TClWaV3LDBrjb81CO8bNjJjAYEtjPSIu3pz4
hF13/SYJvSF0kAri8tWyRb0cBFE/YjUmJ0v53oHa0todicnVEMOTU+1q0QVPrWA17JO/l4QibrHL
uCakDhQiCdpzvb2DtMOT2cWr0/Vw2AKrj9/LwOOqNYF/965JeDg57uy9PdrJ7/Ntq21VaElebydk
DBHeQobTlWpMXgre48hjp3lkFdNq3AKqjIDniZmF1HgLP83Tykr+mPAq8Fm7uYDWgvuGP9fhNw4k
SicsPQDWOqs3UTXyEgDPhLFb5BH8hKb2N5XNM6i4WzVd693rLHo62m6PZbFcRPgm/0m1W00HQj86
O9QfsBx9oHtcGybZVngAkVTcBi3Zm5JHPofXpj/065vAWmBEFsb0islX+frWa89WUxLa+V9tRlfF
nuY1hyOw87zOuV0BO/zgWAevYOIqMWKNeZxhVlG+LLf4lD0zLMZHKvVb8LMhrVh0XxuqLx1bgU69
eTUewKqnINOoJCc7h/z2+HcchYzN1ym1TYWQ5Dr8/1ffVTfcRgBJsJcDG4NXcM6k0eJwaIdoQayH
LGfP08VDTIHj+JbscLNEkIqA34qHdxiAlCYa53O5ip3p4Rv1W5zs2M0MmcHylSlMJVQZaldI4uVV
ysYsSacbEKvApUQmI/4efpTLlvWWZoF2VCKzSiAbQWnlUKQ/RGaugsOaZSvyvmHkys9VvylAXp2k
CLe2ScxrCF4WpgCm5HkF6o1CSlRRLRe1vpDflF/UG3yJi94bXxHGtFCatrGqyALG/OiVRH2wZQD6
yoJXB95w98FuDIURS2NSxZ6qSHc9uvZtDUN+zn1k/9UDKbtTyMCfxAvcl3TR3nudaGpuBgw4ECLV
v3ACARwkegQQVbjV4+UQc5+qsV3tvHHRyRhq8Z0zH7fTTd7tqjWE0MhNTwG1vIT1pOYKVyTQHA/4
GnU9ENsKZZHRDDhin4zgFoun64tfXdS4tVz+G0i+uW3IkhyuHDYcVOfjwAJIkGoz7MVk73FGLe9u
4G/ot/8VOArA6sJiosO6ahmYZQo23voC/ZrEXUWvCnLAZb4nFnZx8Z519R1hNcKjMqd4gz88XXIU
HY2IuYoB8doYLizWWQUm2pgFzRrVlSSvz5XHUEbOsieOHeczCke6V1k2NZK68N4lEiTtH4cOGjaU
rMqQFGIUmvzNRwsD4MN/tTsFyX+0+V+r3pwptinVLOXH73SKt+LbgpU8w4D78DcKBYoot7Wd2E8s
vy8C4gBakAQNnpe5LpgWDlF5oJCU80Wh2lzE13r62h54O249KuYHj4FgrllxX+V623OulsADXsvS
8VIWJLQKrOoLsrCOxfwgRZyRF6O6Mgy31dmTMEmRbqm5TCMWWWjqAfwv4LdF1RH1QTkCe1rRao0F
n5F7Z0cav+cyGJ2GslejwsTMCgjTOeA8MpddDx4QkzZeo6CLJbRyKLkMhWEJ99zsYlJOypCFJHIc
3o6UCGnGHS5mquVLYn/DNzlZF4VkFoZrKMAPF3a40rGFHuJ+SylbqUVRk1AHcZInNk73rDDXPwra
U/TlG0YUTCFOuDcn7DUyLFjagN3WtX0DToSrPYwxdwIPBFCIiTwVOSwLzN3Oe+SyqiJMLTHJ+FcX
rthwDQnejRdy+x6XmxAsWwLJaGO3uLXQZRmFrl1Qqy9+H43banCd3XLJbfY6/6nAPYuLQJNPHVJ8
QBWHR0kCyvvYm8GNm0BFWsxp/XOCPkLv1U++uwHtKTPkN9lHTuZ0GNEAO0YePe6TJM9gDvfEhUry
oT5e/4bUXKp9d0Y65DDGhg0HqEsZp44hK9Z6GUaGzeOyiI1jSr3A4mp7eQChepQPVHi+Fr+Xaz4W
TmMmCu9xw4SsGxekt+T1WK9tiv/Oi7buJcoQf7agrJ+4gFNvHQWfCbf2qqJfzvHsvTND0IGmtJLx
dOBUOzqRUAvxBtnLQLA3RKpn/nkex7DNX6LlKuot8jExG5F+UpfJVGJp5EPJO26y7l/0KaF3YY0G
QU4sqXfE+oraH9CGVI4dWGIvoMUQ7vrNym78Y6Nva+UKbxDgUITrEoFrZLv5R9FVfIeM51xyOxp4
2uX326K329c75rVZo8UgBFDlpUU/oPhkB+iiuXN/ll6+apzts6xQ//mxfuHRgNx9YUgRPE0LXtgB
FARUd/iFbLLEBBb6GgF7L9ignVTJqiDNECpS5pKN4G0tqMClStAFq/oyUSYevLFX2SR3ZXPcpeSo
MyvWD1lXf66x/GQktp0XWkPXH+nk5p1wP9uNhj4KR4z6JLe5KGgyjQIxc2ED4EbVqbw8m4ieut2+
uqm5DUSYKYScFvaOEwdAWP2HURk2jOr/Eddu1WVnKWXlH8qEKO8YyE8z808yVcPRSb6gsF3CqW9U
dpo0i6LOovHDAqhd1WJVh0s5BRC95Yq/ybumxnPXy7H0FgTmYlcX5zV1PNGeC/MySDbkQqN+lDSs
txld9nGx9BtiVod/JA18h4iQnofxb8toXW0jYX9RiQKtWp43uNfZrVEdqjxGkeV+SVn39CxwdeH0
O36+PwQQQcayCF1PEhZJksZ8rnOxkAJ5ifHsULa7VknxqzyVmyA7T2In6n2V9p35y6h/qmxWm9uN
ypHcupP5Bm0/Ca/NcAQpgUX/3zs3X6I+ou+ZHg6B8kJT8aaqAop9wYt4lmyEkkvcaoQhYugdXZv+
5fa/9GjFMbCdk0+v5+RACoKDdlxNZudV89ca79ph4gXKPmY+hlMOXp+stAe5rCubFq8ChyQ4yJYO
mk6IGPkv/fjpdRwlnKUqloqbUZ8BbWBiJbBt0kGUqlaBqLkAaLdkRWVeuLpoDV66zmM8tgCYp53d
2h3LMr0ukAjEQaQ+w7PQxZk8/+T+K52A7zJfUtAsigLoT0gZtJYp6Vj0hi8rL9NuJyqGA9hHeNMg
d9xDkjEfDPJbv7n/1BhXqaXlJwbIuKdWIltstSubA5JEmpYWv29CTDJj06jiABAWv95xxgwJ4xLF
zZXYGtOm0+vH88v6L+sMqPTxMrts3CVeNvOHZcKMoBvMk/ElRd2zIWTqkRU6OI7dOqAujJgS/8It
WFMAzk1CDOyp7b3xCysaZWDL5y9j8F5+hy7lqhJT0U7nvZwwxVxbscutwsFPDnb25QckAYx9b2Ht
8LOM9BMmtIfssk8CpJbuCBgsQGeTBB9N1WRjoZvXvO8LI6+yVzY5MUFhPq95j4vWWf6ddfQgEibK
QjdSM3lz0xlyvBwCHueC8LpZsaU7fbjATz1k3exKG64IAmDyEww8EGD4rpin9CYr+P1aaly/RaSK
qGpcje80u6oxwhmBCkHGqXXrO60ZL2RY+bu3fnBQxwefe182vir0/la/COPfuw8cDh3IVUJgo6kj
TvGttsLAzBzkwuCKdnzMFRdJvtIWBlhYsm+h2PVyOUkXVG7BJPQ8HKZ+OvLmYwTiO5F4GZPmhoR5
8uFDVGaES7weRI2k+ZQHUPYkTraidSyitC6IUx74pifJIcFpa+Ndu8OfXUK3gpXh32xXXpw4mlat
291n5pAAdrkFrpY9CZUUjFSi6vGVFayQb2be6oSCQodAhmUHSIggj9pkwWANpVpE6Wq59yu5g+Ld
jcRnKrJw1Lv7gVmEjYgpAMrM8cTtheOKIFujPJ28xUZDXgJJtmVGuMw66LElvNyMButhPYUF3DxD
Hruwpex2uA325b4P59/axhL88nnyN5FreaBaKIeiSCT4kpM6d3Ha4+u841Nrdd+sd2TjWO6Wz1mc
/gFFNF/fj4Ypxt4HCYR3yIhQMqGQqn0fOSpLhiYYN9kmqDuOa5NsrBJGF5dDYG31JMzIPTJYVnX/
laQsEmoVkKorPt7avJSTUpZFdPCynWTg9tD4reaYIgBiTb1JqlTC5LbMF9Lub0OEfeTNu7yg5hrI
+OI+wbXa6+XgMMvNCNaFKKNS0DKaJKjGBsiQtNiphwPDbU8NIJ1cJ5jRU9sJe/4nzLhgX6UgLOtb
XB2Kz9Q/Ybed/m0wA+6LrpRoD8JiiPbM1YrpfvMxqXy6SdV9IXlDR8V3oXH4PsVaq+FPnUigXjyx
gHgEGzvCuOS1ZN3w/QG9kiEaw3VaLV5yb43RWprFrJ34XhRywXSGuaeyQVpz+Fh43PNZS9UKt12m
kzHTOrm42W/ZmyVypuiwZL52PtneFDdOKcbyGK68/zemacXJ1FW5x3GnFI2/Yaak09ZSXByJCsbg
JVxsiVlzD9Joo7C7DTtJ1DAafjaDezujfZjxeNIJ2IdlD1LlmI/uB0wjiOfyiXf+FR1Iz2l3v7nN
eyxJD8zQtxeq2C0gMdn8kZ0NowrqNqwBpPca31VleYsdT1nIGEqohjGM34f+lkeVNDQwMEGBVprH
GPP/BQC+Mtyv8TSKoO1/7FkcMRVB5ASTOsQF51g9tD7MieWdJ6dSe1GX3unzkTb7l6+wgjw61VXR
lHboM7R2yzDAPEdeVYcySFJQAtWVcd7W8Tg13mVLdD5qPUxT5iygC3cD1q65pNgF+V9vPnCLLScJ
Cz1MrTfEVOfpNNGqPY3efteTJ78R1VeVHGrYSGJr/zkUOHMpoLGgu251SGy6X0s/W25GZSUTwkEP
HbpL0Fx33WU5BkchqhFMwjrBzE+uNqzfyFFKK/DahUKMmPM8JpaKTn3a+WzJt/8g9IvaHpY7MnWA
k0tdME34w0+Usx1CvaklH4sDGpTMtQ7m1Y2bHu5WfJMhLmWfglQRms/ZcHydFCb7aSRv7b/C3ZsJ
I695L23qddLlu38N4gfGHwleebAYSNDs2i6W0h6zqk9qW9O7tr8z8OhV5pJ1nndld0LuXuJ1MnVE
n3tbHzOAdKpD5jTfDsY5G9uZk5+AUdxAypv7oZ2bBi/lz2SeJTYv0NfOQyKn6PEKCYyrss64Na1U
ZZ/cOZeeDeKVv0TMXYDPpW6CpHOEMH7pqNrzXAXBWpCdAifobdGyFZH8drmXmJSIrr0cR/p/Fq8z
6IluGhlEy3VTbGYLcAPGR1SuoP6AN9kXiojmeZjEybDXod+m0+dKHmbLaSmkT+UtPUSp3yESMT6g
lSYlEEb8TbroMxTxdZBuY7GB8f0hNmRCI6Ou5jE+q7yEMpv2hw8BiSZbth1/I1ofui6GpTnWP5hC
mrIjkJVv9HMd6YW5WWwKPj77QhN+cr3sncaPEt3fNFnBFvotdK6wQTBCLzE/XJ/X0Mw/XlVcBodk
FqSRDllZi65YLXZzFwzk+oSioUIHCdBu0AxkVeLwh0OVTIvj5SSh3ypLXmIkHKpFDhp0y3aKZLAx
MgTaX/TkABpPGVbzzo0ivhKhd76HnQeuq8oJVxl/Ebnql9gqipJDjT2Tpse/sBVYgW3HVN/3E+jD
1koimuFPcpZ+Lxhct/niB1sbxU1LBzQqk/J1etpxzJ2Tmc8v1BhP1uPLam3CZBHsUDYwym+i295n
7uax2lgLg10lyog4J9yVK2ksqmlMA5JtOISuYn7/QnoFoYjSdw5AUzVx0lCpkovA92aUGaIhElDN
oJvWe7Td8018aJNYhPlARnE+RQ+VdhXwb1+4TuHP90UQcQwhBSnEKLjac2ndNOZDsuK0G8HtX5Co
lz/1C2tXtmYnEHulgq0PGszrbEJBD6hNJCOdWby6o5aElir4SFIbhyW5CB+B7LwukcW7gGsktC5X
LEX8VenHLIbdGBjPhIBGBl3aOW3ezH6Z8Ro6J9YWimd3yYgdD19xcpD9WmELwLRI1GVS//efjJff
rJxKuXMTa7fspdmQEAfkYeyZFmSewqktsJYp5mjKCoVPLmHZ4TSH0pzFb0NO0hJwN3Oxtjv4XEaE
MtWF/MhgYj2+pPmX+Ark193ZUpil1PhYznyHVjx8hshnWLp6nnJmtoaOXvCCA3/Xr2kOCWf8cgUy
+AA6E0jXxJCKIRbNDL6j8m6vz+ObZoROORcP1m+dlLer9eLjJJmyUVSMg/uJsYrzT/W64buM8yoZ
o7ptAHWjRs1sRJ/q9wkqcyHAg5gXosL1NrT5CE/1fZiATeEGHTKIdJUoVQpl7trI00qHEvTH
`protect end_protected
