--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
oeNhiombBsOKe/H2eBlrbrVqK4h2HoCGdTRp5HX62xoizgCdKYR/LqvrVWcsfP3YKH/8rsPoo/X6
7auJyUCXdA6JBfVneaxxD3PJYFuIrniEPAVsDobF2BsLjvCYZeXv4/55NitjVgVdJiao+mV83ZKV
MxFCOelgkGFsjPdPzYrAOLV/ijFRzrc0Fr9GHkHupPHrIdZeRciEro0FR0YDClUv5cqVFEd0M34H
fl20/LMEcvzWq1E338yKaeTyOXocQGh8h2YBWox3Nw54CouOqwQn9ymiBUvoTqBtBn871FdUU6BX
rA6tWrQjLOmqn++BqiJ5rjObugH+Ka3fI3Np3g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="3qlMxVcP7HC1kHAtxQo0gzqvqEKtUX2HeB13wpQ1nMY="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
SEHaohkk5zLSWvXfEPyDvEm0akm4GP9iRyM80EWf9QZSDDe8hQ1NO+6aVSYzvKw3C/N5TuR0lB9C
bSzvtK+c0zegsjtxSGVtlQyDujl/FsV3yr10yo/9BqwypHUIIBkmnsAJsYvl+vd8SG8YMa6QdTjs
ZW977JF4uqNy4LHmcyBzfSYueqlJwhknwmgGA3Uzw0cMIbuWYyRGW2OGUhXHnfVYGGFQpEDHcy5G
QJYOyzVNYGXKO/C4ZdfyOezVwF4kgmSpcCYCzrCoc3wHEEp51Tx84Lt7tcB3tyj+1yAlVJ5D3Lch
zzQ49V6vyrJLV6zY/fZQPsR9bsjXoLIa/u+RFw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="H1n56BVWAuJSMxUlF0Tibi3ZmFjRQQ0uOhArVq+VB+g="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3152)
`protect data_block
VGFoh1iKUsJq/ZAq33iE1XIX5X+SVPtdI6OOafbj+G9hpiyfO93zyaN/Qsukv1ZsCQTqMXdmm5A7
ywCDtcz2iN0hntGeovrmOJTzcvgcGdFhm6YTI7w20w9GKZgcMQarY4eVHS3VEHfC1sNo2sXQJuGG
d3DAjrmTtQAcQIE+2DgdLFSBLjkMEAJf87vBuWoXxHJIigfZ+SHAOaYti2VgsYLN2yxLEwHeoz6N
BuqxqkOtNA2RSk9A9NgMgxbEAmAZ7/qgyabxLgChddegmGcbnwjGyMWyyd+pVBUicTPiA3Tg7pXa
uQPQWFY1Uro2/Z86T/v5eGnFsRbVvWCbxOSsKnSe/jM3z4BSiBSiW1TVdNQVlgqq+L2+f/X4KuuU
yk9o+goT6QcCxxyCwffo66KdwaKo4ZSrYYqolo0AqCkclR7Spjwtg+2JQyyVxOUjEPfEKFY/15qo
LjHwln1UiRslSwK3mINe7D6nR3wZE1G4UlmKWhKgxermlEPd37l9eHSTGZjE0VI+WX5BTco5MEtU
Bg++Kow5j30m3z1z2FEIBnx6GG5vJyJkrWv0Dcw88IOsiebg8xPpFy4FbfrVfaVFaDfFPuAXledu
jAvQMVDDDJVcPCgGA24j8jiSZ6WufRClC5dP5j0mDsWSCxgEgp/DyRpZcDME/jphcWWann/qY4HX
u3ZVXWGxFOuQBt4rCHP6UoPunBOyMBaE33jMZx70CQo/66ZiOyHORvbAJM5nfONsjtFFsbdBWiIV
cUPIY2nlNxNjtvIAzXSnP8VHTVIfMjPAOgifrVaJScEXNhb7PqKg5FVBj7GCw/qrCy+TT+y17uOK
NsJnB9hI2faVXsQBgmJOY8qAkD2ZZjUdvG7wLGzfrzgFc1r3L0GZ6YEq3UltwrveAag61/HSM7gb
N7hIvmY8/iTjZb3ewvJcYHInmkANn6UlIWoU8VQ5B/sXbWbCcP8K7wLydHEhbGCyJg3IGv5eDCqh
RvXS5Q600DT4rhh3F3fr/dkDq5MnCB9Rh0Ee0wDEjBAB+hrjBPcEQdONlh2nDrxLbYFgVff+K82v
mRAwaz6PtL30cMqSD1rGS4itczGbb2x6JkLm10B1HPRvX+g/zhDQy7ndeCXLHtNbmIm2A/5z8b8j
FQ9NBt1u5HGD/r/rVKOxbleXb3VNqdBc7wTGC7YVNipmQCdjdzJ6ZJj5CDq1wJboEeIFO8tUwkXS
0umFuJqZwFQZzcoqikeSre5Yhfj/nR6EWLwr5s+ReEUZ9K2CZwe0cZBWlIQuuYNwnl83glh+HWle
7HqF6+i9shnojfEEEZNy26A0++5LxxzYJBFzCeLmQR2l5upcISxo8Fo0Z33JNdXLLa0K4PUO6ZWm
zeZhQer94o+UFRzDiNIryZvktGMLUW1Z7O2zZsP4WhyyCEzpiSNloX9ghFKzLaDPrN2kVIlxEg5B
ZszGHjFH2nlLsM6sHMAkvpkvqZo29aO05fUEDMuDMCDGZymi3M4CD+pxlNvHJHdEA3gsIwi+wklA
qiCEsYIlrh64Y6b27r13lWSRUrOK7icXkmMWIU3r1M0UfRoXqLg/EMFGnZfJNt4aPlLpSH6cTcfD
y6VhOnVn4FApkeldcYas+s262uMbO1LJwRhk8Lo8ZhpsKZ/eTUcigJ5qrd1GM0sAJTcHHLkvxKTE
ONxIvXdblhumLtPW8b6r/c+GFVLOqXOoQIy7Np+gTFumjMZpnE4mJtSDFyTly0pG/PakAz/pejup
orD/XU8OsAhx3ibUdr7Ak3uN59V/TzhG0uVoogiJw/S36Nmt4EM30+1ZFglTrBw2nPu4oMfDy2m5
ldL+ePpe8poR2DI+i5bVn5y+rXjq3FsKuWIQ+AjfEbSATyOutW+YB/+jR0by+eXXGvM033qS+wuT
icHLebObluIKZ8eDoYE/DprDAP231l7aOGfG5zbM1sEgFm8FPu+4r4JOLSK1qv+rCF58oJgcat04
MRYOXry2GGhYpxdTyNXdouRFqj1RFFMbe5Mf6/1L+bfTipwcZBzMDmjrUcm0t/LIdgG0AlObxGFv
bK45mTzQIzfgikot4DhqxAWHf/1ip05HNZX+a9/gWbMDwjWtFqHgZtAfeQZ4/AEVZIG7+9C2/JUN
17OKWHfPJ8hpj2IbboKverDh2JyLXJHxBsWjowPuYjhmm3BG/kLmJS6IjLkGDlyqG3vnZlcYYIzo
Z5VFubR+M7SGC4SsvxHbEuoElAd9D26ZxGA1eonDdvcD0DzPX+GGHxYMqnR7RDLOfMKrLvZW8+vJ
v8J3zlTJNkZEZE8gMpBC2qF/4lG5N21TAxDVCRGBhExy+MJ8VuftfjNILTIwZ3ZJMxbCmNYyvy5z
V2Y7IEZi11iT/wAL8okCch+cVzmrS/EKSQOPuOJUik1hIENmpnh1c1PF77galzG5CGzEwj3GXgJa
oyqW6N8xiFnTo3aFSsWfMXt87vDujxJUu4FocBWUOmrnhAtOjp+VpyDFr01MFWOrGxyqHZzmFkms
bCd2mW4yzfgYDsOJ2U0VC/OBAyrefjrJK1H/OyRi7/Uupu3kWOEbz3vWRZZ3YviuNNFamr6ybpYx
Me+1g495LOsRREotn1eXBrnyVAhBTxPWAEocKm5LNUX9jOXcq9RdjAGueSAiRPUCwHIMbCzrauHF
C8ID/WnVZRLXXIov+eunRUT3ZieWqK3+sIREJgPTXEEgQnYaVpEqbrItfw3qKtAqvGlYLoa40vFq
84oJd5v5NLXEwD5SYLGizAkr5HIUwoy6rZ98o9PHQZCMiLkhKcBZ/UcaWzIku0oyklcoEu3o3Ebe
EdXZdB9PNw1z/P88JXApyU/G5qSDyFJGvz/vMe/9I5ZA+saoGMIl0N34GQrgwq2Fwu8NNS4kENdF
heQntVGdze9ZrcbJEJph/IYXd/4OS0rcObPLp3FnmEFgk5Oh2B7j1pEDjq5T5olU/3A7q3gcfZ1f
COamLjQooKqOv394R1irkot33biEU68gccEKRpZqNNJD2LixkmtsY5ON6da3WppFAbKuHA8eSX0W
TbPXOqF79QAeS0yuwD4Zk3OFOSi2nRQc8Y/3+NBDWHfPhMoLR7g/ax4qQplbJwUgZTfngixvI1DE
+USBypRvGE2DN9zBcvan1fanNQckkx3qq78GkamO7N7yGCGa7t0PWCEJzaOWSrExO9X8BeYdriXI
LRURKiCuWmRDmO6xHSCoQAyPbyx3k4G0vNZq7ZM7fN6q57D8aNZkGq4ssr1YRNAhXo++TWmlWy6C
sBmzbFWtqs0XxcfHytvlpzCFWfy8rKW4ZA5xmQL5j0IOPSvDIA8hLUb52M1z/FhBAJImauvapdHJ
WDZI3jT6PgjAJLkCVaumQ0mkPCyaLNGz5YXNAEB6kuaG6PKFRvMe9D0IqHFmL6TTKEBDFvnA1jo/
Kp/UN5tIA+dD9o2ywpWObJF6fP8YhEm5jlll/uXcXFKLXv11PvJUlv0vTrJk++cM2tq/GMkdhwPI
Dj7B+9yTibourHsXp32a+ZNJtqxsgGVeWpRASt4NEow3myOfViFGhzVtF8TXzhUVZgQCJZDl7UTZ
w26+rB/hUP6zpWBgLgzVnvVFxfTFJDux6QlL/cqXTh1h6hktoVcCcGKWm6IO1fDYmrNEbyxQqD52
9jMPYJt0NraeNwCs1VvhlL5YPUaS/CHunAFf9LGuvQYpNpuG1mYaSkSRZ5xQuJzAqgVUkcODiQSD
LFNzh6PgNFbrt7+RrJ2UtzYKRPmN0SpGQf2b6FYWnXFoyOOXeAKW6bPp/V1KLwAPaFJf+Sab1DoG
zi9aTjQIZbVcoW/Cr8ciRQMI90IhmvN/ASxNDiLmmMEh3j8HPeWnHqI7yhhM+V+0y0dc5P7yBp62
wwyDfaV9r/RSE80S2kJwWMIB2pM0F7czBExfzjiB0BpTKPfygyVk0Uq0oSt2PjW5NESIxrRG2rq5
c9WsGgUDdw5Kq5kU/AsoihLobatWKAGdKQ7sES++y+mq0MR/ZJXTiFkxV5g1rWX4m/ANn4ToZ+74
WbspQdk2pd2Yq4SvVjwrqZxmDIOdNsJ77T79kWzkGWG92hV1jkburPY2ZXqQz2EiG2+opbDYsN+L
w6tow6xShw6lmOfgMYiqfIV81voZj1rrichOhixySfQaMuzwpNMZY1GHmMQoTpgaiD+iBtw79Jlo
MzMd3W8lY2ibxYuD1gNuu6U=
`protect end_protected
