--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
UP3KMAN2PfCTIJmuYik69+pXDnkGP4q4EWvMNeKD32E/l2t+ip2s/kll3urKMkIx1j+oOWjQ3OoO
re6++hJdFUFEUH6c2moQEftU6f3p313KUXBedyde7QxO7wv73bxKfhwjUzASitjIjmuA4Hl+goXL
IVQXk7mC9cmQb7RJjt6lZKM+QIpZ1A3iRaM1DFGvarlDLRyScxChBmxijhv8hilrxw6zVMoteDeM
rM5rDExHxLKLuBvS3FfKQMjYUmvCgQREEJmIUfh53RMWYADTDz4wWsLyjbU3VjCyjjXJzfP/VxWO
qoD2Qq3jZpSxNt08CmZAGQh1+8zhf6NQjd4szw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="oaj21onTA4v1jxP85pUc/IaNWqY+gjwD2k8kSjaPxuo="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
fcpX9XesL1rRBSwEt+LpJtVktEWAPstYCLEcoBHjfux7vX06QRhncRA8G1sfZkcnFg0ffXt3o76e
fAVP7tS36HfbwGPSvIYc7lG4vK3YHwMtZCzW/aC+GHQaxpBL6aCkxoCNB2YLx9Y8ggHSFEfo72/d
phfpcccKJcFOPExZ0Oqn9X7h6DjH4VwlWNIM8ElN6Xjqy72+NJp1hCNsqsRJr+Ht7hlIiaVo+Qqg
66iFKNsiPSvwAFypBcLVF+xQlEK7Jw4AlLGyBDoyNGmFQUhX4LZ9Bifz8fLSAtvEuRkQkPxy/tS0
5r5BcZkdVliJKdEYNdsCgqfIpXtuWHQNm/v3kQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="RQ3U+ZF8BpqzL2U4AqThNx5/otb4FcjBcPKWFcimP4g="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13888)
`protect data_block
9EnDLrvlWSW+xg8GWCTRBmuyzTNuY+qiNlwBtaKzMO4powzv7xPtklkh68H4LziW1wlfJjihqaA0
lSpQU0uIsEQlArUbOnOAYF0aH2R8K7FnGvDA4k3esWZiu7TT91Wxer40FZMklT28d6RF5OI27wvt
Fa4+f2yW+3fDu4KUEQWNwXWuggyogiW7RgERt7cHW2PkdjShH6gDiJJqhsQK1CwXBBvK49lKhaMq
VLFe2SqRQXZU1hb5XWMoLXKc7sUYezBOfCIUdjyVtW6i2UE1I4lubkz0JU4OEAZSyLdAAKVIiRd9
Ln0khgJyXVsWnS9rS5d3pKOOWy1DZam/cHzG7priYZ3axvYbOne/cFdgw2ihV7Nlz+k+zrkCSEC6
uNr9dY9mFFjauJGYkqZ3bI0apjlswdBBRZVFmvZmXCf03JfXCjtudk27c/Rm55EYoa4ygL469VdB
Vuc3GUuHDNIMYiRobb7T+XfM7atPpQcHGmnqdS0kXdfY5Bq3gHmbjwl2rZGcNzd5Dp5nNAV+gdV3
njEWSjYjMKGabisCxwtN56vPrIvI1muSuyk4g87UQwEJK+dulqtPI0jXPQueDxlgsYBu3D+BfhVT
1ge95wuzjsjoge4ZKjEuIFksV7kK8hv7aQjFB5XSeFNdA4ob21Z70K2Rl8XIZ/Z1wa5N3ZdmR8jw
sQME1l3pnhe6HtLJMYRoqw/U0Rs10UT9ILuQ1slTdzvLZusDb2LrbeW9yyC6UlQDMaaGTLwJ7cUU
i89UHgtyT/96QaJtcoLTc860bypL9XpffjuWl/91lSwqfi632eZ0FCxZwGB/0X/NzHUI9SkOJvry
Erbj+CSpQN7rIRznWUON0eUwTMwtstbOlISmNYPCYhBgOYhVvUDedjuUL8xQvSi1Pm3NP3wr6beo
Dd6vPZXjqR0JBasNuvEaPb0ry3qubTYwJvF4G/iFvG6AbkW5L8/GZrZEJN3KyZ8eLPWBMtQw74M3
QbvYQ3Rx2a7SC4gRwmT0d6A6mDE/eECUUbgXVi4G9BlymcL8tAyhJ/yIdBj5LLFt4syHLLedoW7r
ntGChVKwYMLNPHiKP6k0Je7oOS6SLkzwBNX1CAssz+CSIupfkq4IchK4EB3saXETGe0eLrg5BUC9
5w4QLtNuDbFYdzdOUaCH3yjCHwMNcHk9xKxaqvqakIdi6JZMqS+sn1QmBpJJAW7mnID1I6pfQEAm
fFNNsIjfg88O/cteXt/xDj9q4gowzzaa9GkVTs3/3BwyK+9xQNJOF2IOyk8Asj7ET9ug+9pCpin4
+00v6Naj9ODObg6gmfJNvPuhAOI/IyQKcoksLBKTtIz4wdNWDQ+SacazmSvop+x0fn3BpwG6B5rR
JlgUVx4cFcmrt7q/KKigJDpvMQd84U25PTYUsmnHgotkD/fcBL2q6fSIzWx79IQ+BuMI/254esbP
Xg29q//H5cuRUi7zdT20n7llPEvk7a7jGfUTrxcqR1lD2LumlmU7WBBQvjqd8qYQKiVOd8+BLwJB
/fJwtXnyZDAffOLmWtv9jXN1qGz6z1RluZ/93O7V0MvRkm3KvJVIqqR2f1aqNgzo9ErR1GUSybL/
Eq/OwTOFCV80x2eq2dtevtMmbvxVqD4tlxxB/EDnI18wB4HLj/ddLSLbYEf3X1nkaHi4Kyk1u3kD
TBiYWaS4Wwf+ePWdAm2KbAOVEo45raCbeM49wx/dJ88r0++L331HkJf0eblKa2nI0kFnJPe6emhI
rvQG1yGBHqRbp4CZJbfMTqUb9ALQbpJ81hzVXSliaGL9Ny1Gqev1iSGZePIfyk9A/7yI8m8i8Gwi
L8cnuKGtiAVycsAA1V8aXorHx/bFIcDYDY3IfCdaT6jkaqc2O2Hp1BNcX5XD/VU7lpbHvZI5ypwO
M4X8KguguGcT09ik1RfqLlVFuHF8JCyCoRCT5x+xuWdWCs4L+ES6rn1CQCW1gC5xk8As+IB9UoF/
DKUUvPj7X7TSHyBuenuwCzsXIYh0OBCVa56pdvlTO7D4dPokU15QeqmhRMYDRldpJPHLguf9NhER
GRzTWhABW7LYF9oDF3J/DiD4AU5gVHKQsFig8bWrrt/LPsiLNcaB5rp0Vc6OyOyqzEoHWa4r5tp9
nu+RwC06s252PsrnBbxDB1xGRhVZJEA/xFwrF4gDIvo1xYeGEbRdSqztz+vAfd54su0VvffHoHBd
3X9O3xcyVpolR6kX1HuGKsqJNVYIYb1RBdaM5GrYspo3HM+yeWdsA/9qLc0QsXlTvZE7fHFP5lTu
9HR7A6WiNUOHc+zWUnXpuWsbHprM/Ei61SRFUTf+2ZGMKXaYE4jYZ8em8n4E1Irnmr8wA87RuMyN
WF5yTLHTsdKB/e8VJvcoOONyaE84s1gV03+HtA1fnPnBRG4sMkqVG9IkKK3iK2vEYD2UdfsGZUCa
/BXWC43cimabDJ4XDJAAUAiLaY3SJqVNMaFdjhssCL3c5qaT3omZNoMLGdjQG+XKK+c1hphCT2Ym
USIiKNHbUMGPjW24N3AQgwtNu1Z9pC8aN9qnnLztI92O20k62Zl6K/wY386etmlcS3fab9LKe5oj
ISsruozdQPSeyDMasfk1h7LcOkyyFyh8LnUCqK031rQSw5ZEmBBNGjPs2CMjUfH98NBR5d0m9Sd6
iQsWKsIIhSR+jPJ3/UFPVQlySuQQ7G2BM/ujasyo6ILiW7fEzVfI4jpE0vkey2nOhU3jLmM9aklT
e7RLsBYq5lysgVQWMc7mSw5fAruhl93Mr+wB3au/6XXoUIM7+0dWgv4rNh9drp+B0x047rmnLo/P
vb0gPykIooV2uh8a/eiuag/RHheimlQFDJp1n54oKFeH1w1rDlYduj/ccBbmx9rSSbnWZdjVKpMO
FnXzwVVNRP7K5ip43Fbn2EisPccVNOSweeRGTsxeDx564sh22jDh17mXanQSeesyNxEDkLhclQCg
ErJEKvU/RXZSLHJPuN9XiQ3YSz9gGOSd//SEHjiiUM2RYuEZ6XB71ITa0KOvq6WbieptWETj+crs
fOYTFhbDGxQhF3QMhFx7Y0UM65lf3HJcM2etU5pKfxd/o66DzWRbQAp3hZpjbsXic71xvavZBszG
VIm8jSYDjZgN1SGmlXaD+bDS/848d306kxnXGUB8oRWR2WDi6HnpullEMU42CL2SiogEsnlXY8Hp
5eKUPMlKwEYRTD9r/9J7l5PkKrBP1tQr4bjgSGiStOyCxQNGzKOTDV48DKdY6+IV+sa6/01L9w8Y
B3MD6yoQ41WubMTrSFZCdYEBMbjztaqSck6PzEgqQAox6avubUC8Qk4NCCSMU+1MZ1Eht3RpzFa0
DwIpLYge858FZzIRu9cI5ITavBQgiZckycS1hHjp6HMHacKHpckis2JihZu2YElrdjAV9KUdFoEc
bKXWaRmflX/VXNrG/FOBv68hqGUys2MnstNAZsrEdAoDlbihnkYP79/uAhhdmJL/Y8OF1ztShiUG
C2h63QKZ7Ohf6jr0PKIzdaglNfwC3XoxIWjwaXjHPlR8QJe6tU9rb5ITBfDtiBRrSMbOwV/6HPaM
jf8vBH9Yp5d0JmSJUSMrWE/spma3botYa3qHjVY3z5RNOTsioW0WmL90Z9GV3LJWnS6hY6bsK95u
k6OqEt1qrXzKUhFn7E4hKymxZeDe0JfbfDuvfFfgLroTt+TrPp4eLhVKOkzx5Qf3/Dq6ltE/LKbo
xqY9U3qWHCX35FNLsXmZEcU/XWd7Qx2Jx0dnQrWnCDDLISfvIiDYVshpetBNJ/Luo8yNha3w9/lL
/cUJZe6j+jCKexJ2e9dDuvl/iMIi8pKkkjia6g04z/ZwL/LYwnxdc0/UIs+ZVARvDs6z0qYCG+0a
6HMxJdFTNqiaIp8kY+MKknL0hjPe7tTYDXZSWcDyUc1y4QI6xkJE1PgYezYJzbUg8q9xzkl4n/bw
NnHpBEVqS0Lt2rj/uo2U6frV7hsiiljX2CYh8051rt5Wk8YJss4FsjnKPl28UGO7TItXJxs258J4
S9E+YFpc5Ac4XO4EkpYNKE6aMtt4/LAiSMguqQRoUSAJakvxHVEWg6KQ11Ow5UeXc1t7diPa6f5s
bdYjxvASmTpdQ2afImYBiro9N4LdpZA92pgc7wg6vEKYHyWhLCt04pSuJYulcJhYsZnT+qMS1Z1h
9+3uZt5wefbSX2HE2DkEO5UaObaJHHLyQK5cqzw6Bl24SFX50W+Er2shiwoTjBEJ42UNQ4gFfHyN
aQTG5Msxvga/RoEb8X2nQe76b+KFGflDY8bQ6vBlq9Dv+W3ne3Y1uVVNtm/jbv/0wxg4X1qL2nEq
5g4izwjfh681zNeW9vA1bYF7PnPGWYmQBuMjTc/4eFbaUlcZ+ONHh5jnMfJVej5TncqNFAC5HVsC
mPARDhQYORyWo8ZAH1IgLd2ylYdEqSItxjSAcY1ZMd9ZE5e+PuUaf5CDPuAEZuhrEgnjMYn74XZw
zr0kFVPYqZjpp7BTLxHwTglCEXwsD8PKxsefUYd5+R8APKIwLz7a4HFBtgrpGg80ur3W2VIGa3NE
NQRziob8yPWRXxNs5wO+My5tlRbsajMojj5PF0CBnxjI6M51UD+7xQajP2gfVvQh2HfO8syVGKb+
1MaERSMbkxjL8AyiVnMZbm2H2rAM8Te6FS6lfHkEx9JV6I5HPqyipmoOayxOR6iQrNji/WfAJMnt
BDFmCmyG7Msp7jScLgynXQOEM4VDzYaFPlDunYLM8ymW6+PLvRfIAKONaMAehrXImAeL5yQfn7zm
In/gV4//y91O9+m62pGfbqF93gJL+8dPkZ3pZ0U3lWS0I+wckchl9kvvp3fQ0CDkXrDhmA5ux0FE
3c5rj6ehHtZxLouUrBZyXHPG3G+4eCoWrdqeOFz9lBcii9xRJtrLIFN9R5i5GChKxfRA1UudykpI
t+9JwnEy6z3wdziIhouq+hV9/XZOHHtBF64mzIFCP5WavGQCuJcWcPo1QFbLnNa+PKh8wRlVtlf1
PU6EjAxeAU+L/n9Ox+Ljq1swM4aDyo/xA0qjW5+sDAb+eO0cu4i2b/byz976a2m3zhdpoQA5GTaC
YozdzHxtBLftg5XZmNSHDhkbbXgYWns5+GVsBQ/QjiDnbaEJU8ghHaMRtEjgi+ouU3X13OwvOBz+
6GSNgJ6jZ0Xcyj7IejQOOxgDN06gckjhlgu/UOZTtvhw29MzbeD0wYCmqs/hBBRID8dY1QoGK1hp
y9sSJR+gEZr2JO13OqNDc3lgDje7v+7FynQU6DQETzYvfx80naAsmAE+mgflAsExqdVPLtjllycm
IkWGXdHU1ps5231Y1SyGC9kW29qiHAhWDvlahr4tUtIe9StPuL7Z2mCvovIzoaDGd/bUrgsqb8mR
hNUoeHiAQfEWp+KerBoL/7sSObs02xeWsi2YVlA2dzJFOB/w3F8eF1gfcCp0xkI3VgyEWEy8qW3r
+UGhVfvigioCmBJnvCcTmUdkhqRndPzUeXEHNVA5qBTW/DBulD7sLr4Kyd2hQPnMnUCcCN0YUHPt
ZyqxrvbtiR/3hAqjKZ2EHUD5xb4pYLqTtfKd66VGMQpiAHCNCOdLyBIV8wt23eeB+xR0TyCirAWD
5p7ejH1OqQt+d3ta4f5JHpmgRxPVngwX5fn0FwGWzaK6Fo5aPyZCj9xs/VN4d91Hove6nwn5UyvU
ftoniJupgyY7HdasqmjcZqzxfXCc+V3mHbU800EFciqZM2utyeFcx9e1rZ9gCinNstYoBsA1rT+0
wIt+H1imCl2ik6V/BytyKz4DrBn7cMCQSSTDv+qOBeM6u4WIggOS2/sn8EXLycQTiE/L9jdxp5IC
FvKJbzwM3MSwW6TXVKmVv8MjI56GAjFv7rAIe2tr94XrVcv9iRFpOFCOxN1urqhHgtieTknxTx6p
Hhvp2g1aQR7RlfQ72wPky6NqDlQnRTKbBU7I7S/i31iKOfJIbK0NIl4BX/qbz7UGdHNA+my+3Mdw
ykfDYLzsrEOUQEEBLFDt1/GG+I7nNg3LpaWyNTjnF8oz6ar13/tsahwqwUlXytH8t5Z/EU2Ovcsy
iSSvD6DhIfSc35GuIPoy/exEsKr7whLUUtkX0kb1Nw68LGd7f2k6VBBiJp2dpHwN88PR+zQC3iC1
jWN1R1ImhFcwor2kOt9YWTX/rq0Ih0EXZX+VDvogogNKHK1BOtDrgikeTWeLFSW2BMdxOrgKUWwX
Ew3c9qukyDy8vMdpetWiUHVny7B7vg/JRVZ1iB/nnelG7oNKzw6TQeNTKZv5PFnAPJ7sOmnkdn3V
6fEtbzZdEWWLku30P1MjucJrQzU3aOK3yVyIPxcCYX2UZ3IrnbdFYIPQOCbGwsglqyJ5gIOHoDDH
P/yRpZgK3+blcMEtK7y/wNeh1LqFgrcC9VzMYA+3ULv7+90tcLZmNGXyIXGyhoz3/XOksl5jGKbU
eUtoJqBZ6QIItcAq2n8OIli+8FDVjtFLjJQSINDNTT9UfQeCvVWoNeTSrB6S5QkFDx3UDppSY6Op
6CkRPpcIAMOyMRgIpjLip7NoKX9Kar8OazbhX3L7FzjuMBUaNKo6uzlC09e/nBcwFmJrIGw+GbdU
o2b7Pdofm0YldaRrcLC/U/wozdINjtlK2sB2OOnlGuFJ2Cd3DFhgRpwKKxQm52YdW63XggSE++wZ
H8qWWR7JGJUtoFK0Gywo1H4YsV2zvNjTdzCUxeTlLaKj2u2bzb+enG8Kr03EN4J4qyj+fPdYUd1H
pmGAuwB+glt5qDurQQ/8MTUUQCxkhn0cu2Sk4qPHZaiB1Vp9t0mfJ2sqxDD+0MNpAD6X39ks9vA3
Od1paYEJW12bKYaJ6yzHSevfoNAxO95f4xJcj1XMQh1rvvs4445YZzxvvy7hCgzok07e9miDCsSt
f/8vEP6QklFSios6iYy9ljqpj+UqSdmnjpEeZDxcoUC77Arx+wLsQ+3XoIMHTn+6iU5uI9/hrYqT
6Z2jMRmJxZbFwOcVm5vDHudn/QRgNXf3vI+K5uuiDOyjkXPqI/mRjg8XnWLEqVLmyIIw7MW/GJte
pii+FfLxys3QQCskH2AVAQe6EB0d1L7xWiMqPf1BqKsy2uyGFhCG3CNdEpSvZJGKJA5XMEDtGGje
M6+sNYphYqRzd9SNZlo7IUyauQOW4V33W/GYw2LqlkYVQXI8qoWdH2IzeVcsbSe66HEIrAcK6fvW
Z3RyqgurNAtXavlLNEgNx/iTt0QhmssJX10S6adsCD1YBVZ+7YsuxfbOsDHFZSTKvEVHdAhfgBrI
3DE+Pd39SIi5vK6hTGOE/WtQOC4qfakeWiQi3Ap72FdF57+J6wIzAp0vfCXFy4sLZfFwfqclG8bK
0AtaygOxa9fWt1pisdcV+EloTbRHU1R6c4n2bL3LrsvAUHQH45ZmFY9B1sKLBhJZ4xjtIqUnoPVw
0mLNsNrjsEposEmp1rf8lxcIh5GXJ3eApJq5TADBgKgCv3FlBFk1qPmHP0n1/aN+PcBvwc82jOeM
bQye+iiKsxgXvLLyCnCkKdipUobBLo3q5RF4oZZK24pTAhNuoj8i7fB3MXtktS6FmS4nqM147tWO
AUsHc63J6yi7FKYVa/uXVW9Fzs+xxaalfuqjnybDLvEyIuxedb3bXdt97hJhFtmjKAjaP3Zq42P2
4VQ+Q3x2jROJ258mVSUVtRvryeCnVzrk7O2Amign+VIHO7e6wBJe7RohGnivN7ah+awqIc8miOLE
eKlX3wzUU4GARaez4JweJnGJZ+QcDU3J1/0IvEFlA3okyNAAvoyL5DOEqdsXxeop1sMsIKyXXo+7
ZM3D+gEj9sbFzyHRV9aCsPBJZVSikZ8tyDrEg1NysBloTvelXVWRC6niZxeP1aVhmU1IalToOTOe
GYjWYgQO7o9ut+Qy4sy2CLjh0UOKF4eJTFYGvg7OekCvvbN3C69YZjl2p8cAn4jzn3exGovUBhlz
bze6w1vjxNaqRlpPpQ0UajAzDcSAKEkBs6tv850Xc/MG8xtzhzmysnzyL/YwHuXeNBPOaXF/twOD
w+CqIMVj1mNKky7lXxsvj14zPLQ9WJLTMM8BrMpBVGkv1AuF4bVOJhXEmWbi0ncOnYoH+AY0j4T1
9xD/8sX+IgCqAEBA5XYUnQY7nwxT6iCW7qEY3QXx2fdyePBHlu7KLsLOm/6hdGziX52HQGRzVODl
Lq6HY/hdT4HUKnp2bNtilPEyOC27jkVD/UA6+KTrFTL6E2IjVhCKAeBCOFaf9vN29jrwygoZ4jtP
ZGfF6MCIjO9y1mTu+X43kbDxP1It4yXqp7Ut+qC+u4wr7GmMe+rV2Ty6jOex5dt7xkmztUVJo9UZ
1OxeWFGI3eZRMzjXsvLBq3609l0lsl3tdPjDuSBRpdcz9Mh27UEKmsBHvH3UfWF3wS9FGKKNSshp
3kxd1BRx9hwWRx6qsQWuOnRWKsiqkgKO6RsgtjtG0NP0cO/9USH/WngGV4RMU4JboWSMJc0S3xTf
TnAL0SwN6NgqzYnAB176z5x0QBnijDpfzdec3fwKSh8K6jtQnLjjjZ7IJAbWYd/t4s0jOwYuk0EN
aFLNZFcUlfjD8qafiVhX0zryEjtjWH/pPS4rOFOOzO68RdtFBIzLSJ8eWdQvyQ+70QiPLzqux5rJ
LtfyEcuSY5XD1x0RrB7YT//LIzJhK8JskJZnXrdaQ27usnMja6y4aAKkAY4yQMmT6b0mviBm9E0s
hXxVyO3lET+NMmoMlPEdgyC3CfPcfuMJ+m0yFiNrk8AL2S2FcJgoSXH33pOOcBV+vk1Ez84f3R/x
Lh9/oDbWNhfacbPzOiLeNPeIh59YRIaXofvGWUoMSNO3tykIbElS7/tKYECfYSimI7Xe6/mtY4cF
habVYID5jtFZde47MadPhuW5dU2QIDS4Vs+DtSfkjWMRYv/i+DPj15wbwvMROWoVpeSvumOaCBNW
zvf5OAt7itXqgZZPzpwUmKLoYspnuuwBd9K7MhzjFzqz1424+r0EdpjAYa3oANwAEj+Dq3oK2IVf
BtQ9NcxlFke1g+60c94XxUZT4bDLmtcrob5WrouMOcZEICW8sWeOrZDgS8+JB3asQQKOzLp9jqBl
SdVvbvCTrJHZM3juF7ek2vUSCa4MD+OZoQVGSgeh2beMVILviasuNEtcWqHSyTdbVIGlKab//Xx8
fQ5/8FPum3PtE3qc8nZ9yxXvgAvqXQkMqsd4WsjIoP5BnzgEFf42tmJOJFT2PIXtbX4p0UV5JAMu
uYU9orBhJjte1YJg40ggZu2OtjCMb78cDE5NoXZDARBYW73o1PNrPWp6TDoU5C4oJ5Q+QzhscY89
0r067Np89/5BQt3zWo0Tx1fiiELDTrSllkF5GLCOpsLEEpG4Y7KZ8E3iSj1F7UqUMKu3hQfLXwng
UxtslwGNnUwyiLtr8z11ln6osc7InueJNT/Kg8N/inmzREbQhHgkqAucGEp8YpvszVPFUg4Cg6L6
dHEZ5fTyV+ICFXUhIPk6uscst5AXPgGjUjwYZ8LNgO9kDsI+ctyd0PDUevGEbi0bTCKpI+LaXy1K
M8JP9nd/VeuUv1M2dG8i8DUxGxRf/7gwXtFZtYWszPTcPSbsqfeVh2r41+LzVA5j1xJEd1ZKQKmk
yNHkyGDWicFibbelQ5v2hLeZa4pEr0MKwXzSTCzP3vh5XDIUjalelosVqgxpJsNn8CkhnPTdyCNx
TBXu8XSIvkYqtCTD7xMLHLVklTY1VXAIew4mMMsvqnYH5FD9fOVkeaMO7PZilxMBNoa+7hwuL7JM
W8Mb//hP5jL9sxiG1wFDW+RSpLl7aceKIPDOHPKtO6o1MKixDJLUyygMIT/+1gdEuKvHoxfKO7Nt
na1joh8Jm3hBs1M8XxZPggb3ynZw50Mt8Z6qPlKV2Q2U8mK5MNorS3SEh5D5f68uVH3evESEDclo
u5HC4n9Xxd6WYTXjTUC7cOCtdI6e9KWAG/8vwhX+5frSKxqPiGDerXkyk4nN2ZBIc8d0YrjIBjH7
ukHJEUjUCujxOOrBNCrbQmWNe1rWZVGTCn36EDKQ99KA4Y2cmr95A+6gBQiAgbkC6zweRIwOWIti
UFyBbOKJYHefgkP/4oWe3odVVe5UnnjFQG/rlaiK9ui4PWlb+fwE1HHOfFrA+le05iqJgYX3Njox
1ItAwmFHNMuO3v0FdIGz1QPYI8enspzuj1enhKifis3HXzuvkiIoglttPpw2AT5+SJ5EhKFO0S+u
GtAuzCR6m0da6Ekf76qdKP9a7neq2ji/w65wckPurMtWbGeZBLKLFbFGMpHKdKiDg0q7VZ3HFOe8
wf46cpDrOs7sE6mCYD3t9FsxNfVaCwyNoW0fEIN3zRPUT/6gauOkFBv4fY7TqRyv0AmqJhKAKuti
tkdiAvo4q94aV8+ywdFdlHpCxIYz1rRTq3QLnsMpfomQ9smvZ3fa08amzGBJGLvyhuRDVAFva0Sj
ZURIlzDa/X7+N+VbPLP+J6dnMLJ+Cu9lYeN5M0YjcSq2u7njeLEhkwHSy8ZlLlh43K7HlZtTB/Yp
MqH0pcpHpnzhG2o3h25r0TmGlDhYOoQTHmaH7H1x0Xw96etWw/lS7oTaDx2JxuG6fp8eit3ZyoEM
lLECg4zXqERK1zvPXXRtuzQaTLnsPkaocId3wfO2/ilU70Hn/8uplHOWFLpKxV9V2xkMSTS///Y8
Txg7eafHY62CiymOskNEMK4eA0ukFe1+9dVg0Xw7WgzcoXaYGHtYzBvOxWXOa57zRMmTTdMfplQt
vLzK2asufpYaNW+oFk7zdlqnNn7Mo0aTLslhOx7TZd6Ldwxg6h0YaL8nUl3MPG1lYin4HOL3z6Kl
GehAqFqvyGK+XW/QPJsLnp6d+vVYvOVwYCOoti+j2LO3sXEyD8OUaEcD1gE0UW/+9t3r9MPbWzxT
VjHz1+1wQXTeneAMDpTGL3SE4773Pzxj/l7mXOadcGUeRxjztLhRqdZLA4rtDhoKUEw2s7mAm8vu
e6sLON4r0wgcM21aa8o7UOG5UqUgY/aup52erF6i+vN7KzT3heBbNF2GdQT1tvS1s4u/7RZqNcx5
f+thmZHNU/3VhfxBjsQSpAzaOQ8ecbnNhvSPan1tSvscWLYNRM7M8znZWyKxY94ywTx6H6zAa9tq
iZPyBdPBJ5lqiJtPDzs2WOwFmujnulxW3bV5vBXFgR8CyjhIMHEtyw7IH+kuVM3tbfbcQFoZb3rg
h/So5pmgOXuJLoF92i/cOr3YrxP1KBFrvbYU1bReMRW1NmiyKyQArDZSNZ11ccG/7q6suEPkFUI9
A7duJxC9rT+XixrdEj4MIWyS0INHFn+fyrkMjequWOYvPu8O1e8gs6E6R25GXHeow6omzEYIbeSc
6w7Tp8V4uTN/T69FRNNc++xzM4UZTcxu2+Mepuh9iReVEDHq7Vwsog1WzP9wgK+oP2XxAxjix9qY
N4qbKx1obdBbXlNFiKkicoxeSz1q+ciYab7EUpoYxVif4fxmK8qCTByK/5lVPpX4/iUaWZnsckDM
5eRcUQcMGW+UiXrF8Fn6jE/LPrFWIXvDv/CvOccIpMBHH1q0VQbjRQdoPIAZx1yY13C7iixg0Xj1
AabCtlLAR1gOK/ZBCrgq2HA7H95O+hWNi0vYLUdY3IxSvIelGTBUU+4VKbrht+1BlpPdsQSRL6lu
/TgKU7xtlChV+/TW8HzPFcjdv+JUkxvtw9LAk2sqQWU6sZfT4nX6UQlIrqL6ibufBaNwd4IwXAw0
/UBdT2wPOqOX0LKFUqaWDDgW5kdpZJyavXhi9EgLl6ukSOxPawSliPrE011UV9KZURsEbtyfi6uX
JSDZck9mQ14nJwuvXP7oZZl7KQwL80tVXn6IcXAlZnyvepaPltJ+aVaB110ReldlnC6RpwBRYT3T
3S3G5gIthFuWgcJnTpNOIPZTMBA0/7Y6gmAJt5/W8uBkFWsuUusCmz3jFf/UuTMUM8xZjWN5JqeW
UDimBCpa/gem0f1eB6g3HolStJryJGOfp5jmm+AHQR71myCW2e+5O1U2U2AEabVTFNuZ7Y1JDdTW
GRleZEHTVrNxjH8+m68Ewq4yLCaZERauTjijlTXk0W//jVIMo6ygAtgTT2q4fFndJKGgGXfVj0jk
c9H7BfVOl64gfV7C7AwApiBxXtxkAc7DuzpKQ7PQybhpI6nZNUJZwtJLuz+GxQnvgWE7WN7ZzcrP
IUCVxuLz/i+HsSq1YRbjIbCi3qb2YQ4O7o+Y5Bvk1NBQlWMUUaL3mijlVQdlsK0ASCR/n4NLkNRo
axpU+1G6QiejHDi9jA31fsWoNRgsxuHTzXg/TXp2065ZJBO/WFGvwI+QH28BZDCi4WhKVCyF8FlS
V0PwdsSm284bpX61KCGRm6cqXyPKyC8YRyLLtZOt2bUrRgp3b94lur+gECjg3dNsYnTGMZrTuENr
KX08UFRcqKPWweKAQEXJXorhAlElbSZvbG69NE/HCEKckTxjCjzDEoqpalWOWTEwttrZEEyk47Qo
nJykucGfwHYmg9DKMkGXThEZ62T6AXzp6sVEIGeZF6r0qCPgab4J7HG52s4iMJuKDgq7sRWGdVHk
xycWpHHjo+cYZdoUHVfFuYyhH/i7TbxrgVjceZxORFwEfp1B663e/lzWwl3l6ni+//pLM5jbYf7I
9iTxxzBO5dHANegEUPDlzdETlGf9I64qvbfyAlI25lUXlaEy+ZLJ16j0lExbwhhrMWtpRIeZ5jfp
tWNotnCAsIqFOlBNJNK4jaoVGDCphsdAmyz5nnfcsS/7HOg+IrzKdHhBXjWylNjnOvv8TrArZtAj
O0Z1TUveZQnglvU+pZKkKGCFw/0sLC76MObCQHH+IteKdvSncRrd3cBFjQO8dlYKVxqK1BKR3A9F
vqZdQSCYu1G5F/j/B5BTQNfZpM+sZESnVotRvpePjIEfqgj34A6evEkawJyNSpBgoqgP1m1svLqb
duAu+6ck0d58gCuU6EUQxrra6Q7Uzh7EgjZa0gHnSZwReIiKCDR4c+pWqVMj9lXvZmZFy2Usvmy+
k9mnx9ApyI3MnTi9rT7GmlukBqlJbHLrzELXkYR646dtbdVs4pzlhTTgUEPxfzf05M0cfCGE+exT
LkPm0/IXrOTAzLETk849hVfk5rt8dBIhQJ6Iri6WS+vFJi7lRQkWLiIfOErZ2c5+14naHBt6tJsF
SWKyzV6Se7CvlgMU3XnDueraXCVYr7T+qbmQKR4zU6LahjhZ1DpoB1EC2pvd0tC9K8UTcnYERJGg
c2RMkH/X+DQlbg3lYnuxrsq5e6yxyPnDzlff9Z/yTuyoupDzsQJjiwh0DJHJ6NICF1EWun2j3mXR
yUiipkuGus1cNa7ckCHn/V8Nozh8fq3TeYa+ErGwcyUQZ4gzNA5kWpltr+gy7G2mdV2TLwJgVRJj
a/wFH7FtPIGa1nXIwbe2qOYtf7x4fLMzvWiG/lk1bh42numZOO1mCVNbGYzyAdDdJW6k2TaKoq5g
NAxw+NWIqxiKHsNCi2cmAn4mjXiyXkm7ZvVnhSA+XR2YqVJX1CLCUSk61JR2Zqox4TYPZALUqjj6
nWr/+6vpXPuAP2yCo8XTYahaRBeWJgVIZaj2XMQ9Z67zuKexhbahXqDcTYT7SOfeZM3KT5KEJDM6
VMfZrmerf+Q17Q7i04ynKwzFjlH2FyeMfi3wAnBjQfIZr7DhtcaGbebHE6udiX/DbjpMtgdrupTc
Mx5LPq3Zq8sVh7ZtVO4lBPln1/P0CS2A3g4BWnM9hwkR3WkdtArIPa6j4w98LWiPmavSfEHq1T6a
A2hOnJK2jEUKLOoX0BVNItVqZzAQTp9ewYSzBZ4KUnEUl1Pe8gn4GQiWYPKHVyusX0nRwJXjLi0w
PldK1jnICohPeLuUAFZkFq+gCUtqGpH+ibH1zx5cdydw8fP7d3XgNXrTLCWBITftzwAtBesMgTKa
mNL0QmDoYR27E411XBuO7WnDivqDk/HEtPmWPFSKDFEcJFLUL/4EHREMR7FtGLQiCn1sC0/nspMT
RMQ9Io6ua4gkdWbWVnvNCjjlgRdm05WH2eo0fY4HJ8SCjtncrwFQcH+oWS2yFYxhqLDWOG9SzF98
Due2pmNc5lKPmKpJJSi2uFsAyT357H8Zr4w6X9UZFG84QeFK6b6v8IB52WNbJ2zTCq4dSrJFE4HO
wsNNerPrZDphyHaJrIVmDpJ3APcVL3OWTo5L+fYXx9wNmIPwAsjzMMHb1y6GI8FZcURPF7EIMqyB
AtoMjLx3WnOyJuzzIpaQOgPNI+vMhaPZAqPOk9buu1HSilLQfohwEfhQxmaRataP+VJij+yxRMgd
M4ZK+KkU80DlT1TEIeZxo2ggLiV4ug9EHRyGjJf2xZS8Atb0PfToPfLEX3gzlRsrv5AMKQi+us7b
JoYXKF/wM4QFiq66Vn2FSE7patxgwUn4qxyp830p3cNJEYHuCmgTk6xrd00wB8MHbIY/6jZWFPYJ
ehl+/xWfO2GF8aLvHpyL61QXZbXD+VtC46m3oCwgJSPw/Z0MgwIJaUy37qnITqVt3QSRDSqE4a/f
23CDZt0E6BIZsWayGYhiIGIsg49jlqklKL+p1s7DwCFy/ElTORpyRkhJQAeqGhzpvY7ul3XtXq2T
ipER+9LQsP399AZmCsrzz1HQcL8DUh3srj6Jd3zIVEGrvmv7ZVriIPu30R/2xPVgkib3O1vAPX5R
F+JfUZv9rKwuxuNJC+jaPLKCcUbT8PdizjCMPUYDGO+y8H3NVgTHPVpk/xKIiZz9GBj0+pTp4Z5F
3MvbOX6bizITb1ct5gxRhpuyhPeHcsIR2U8KjWMjXmGh6VfwcCjj64wL+uKLSP6Oi5FKvhBfj9OD
kk634lkYjHBUF1ClYDkeCi1FK/0y/JKiM4++vQG3RgWk9UlkqEr6X9unws9FBP5pH8DGgRt1hJBK
mVBvThB1oidKz67kynLp1NVjkLBiJl/o/RD5KFEF0vVdBUMpjM1CvVDSOhApPxKgC0NSNMkPeOnI
OMEDOB/cD5KtHhnGvFVyiW5jDqYklIF5iM0K2yvh9pVWG8fXW8qPhQizJg/NekM9mohWB894s5Im
YQSN2XHXXiPETECFbPCW2INRk6k+x1VsV3xQZk6PQiCFCu6jqVPqKhSInVe1TDXNC4lM5h9fitBR
J+f7972RPxXMLIt9FkGwcnzDsi5boROFjSrm95mTb5dhIgvjEu84guUviot+mAzKbUyMID23chSQ
lDOzaGne6BzJyPok8jUfp6DmWJVSWue11S/ke937qGxBJk4d/4GY5b+TCKV4Z45n41kVJJ3Z6BVq
3xqjm2VaNkFAXMKlcMcT7LH3abAi+T10Uvek9MewJOruFa+BoFU/viVRatVB+dDVsLW97hrPMwp7
19/iTCfqFy26P+htR6uSSxX0StBP9KjpVb/bGwUAsaaF8RB+tv68xTQH/GXqMejDbiRuM1uOgYEF
qDNnTwH0M2a4ihIEPoEucR6ECnpeBzISlXQfHs3b0t3TtjDonWliPpoIJIP6h43kVKqa9zFtbgOY
+582rlkR0uf8MqOM2WoBIrU0wilgtiTuOin0sbgaky2hRXZr9Kh3q7QgAcZSsNXrW+PrdEHDHep/
Mp/BitRvcgdTtaG4BOmwxjsb/a/isOvtbhR9TfhQxMm9Ea/nj4+TRYVQHAxKb4usyQzFK1USpc+p
WaLVSl3gMdCeew+xCqYejt3w+t4Z4Mb85oi1PWul4npVR9let2lmXfk9bF6aru9MgMPL57dOdPFm
ZJjHx6l7p4vH4CIixYjcD6H7otkKCLiBKhBlBwqG0Mx1kQLhVGQkUiYakFmnLge8lzm/stk2Q0Fc
y2gxSleWTSaeqGZko4X1mH7KF81/r1xsq6AkTm9lOjj7LV1fA9B+vVrDy/TeRwcCTM7CkAADRGos
ro4RIQh0uUIUfNqG5blCjo1hWCom5ApBfYLTDKGJcuWRXhYM1KPF3qBPlyHS2bukm0hSn9v/1uLZ
/9LI+K9RDakxzbdIQf4wrpvfzdELjFMLXnvQ52Gdf0Y9FzOIKyJ7SZvybWU8/g9K0as71HRme0x7
GIXg009hXWSxCVQuTP1I00Z+ZU/CqH4CZ0MlsidaYY77KxnpcSRvIBtlLflF2Dm6gUIcmutvbGL9
ySDKw9PtWfLcwWnHPnps64vaesUrGMMo5b6cRdmrzSxevpSbtekybJ9YYXQD3l7QocsfxZcyPaGH
5/09nU4b6lvYPQl0XHQKUgzZsZFpkSVcA5i96tfGWdV5r75VS1ONGfkWmNZ2TGkuK4ONaeqZSJzO
n83oGNc1N51vTr65uY/OKaBcikSnFY6bris3U9j86b86uWfARcJhC0R5as3kGMzCte0rbwKFCFKa
9JngoL2micCAb0hs8FCcysGJr6NS4+sSeF+4vFFnaX02Fa6avONMQ7j32FzWX1AFCxL0LEWRfHqk
XdvtTeIWy2kZAoKl7Kcx69wCN+E5Fw2GGytdH5EuLTJRwc3TLwigK5hruvW1QW+v1Wk5TRubYMX5
t2PVqXYr0sDzROPV2iGkHuC3NmGU514OysMj8LAmXPT6j6bqrMHNfdIXeUdAhbfkXhfNfvaoneOe
NeXw88OJKmKOpz6XNWriJf+d+ff4Mg3SbOE/0b7Fybpx0Hgp9dvB/irJkM0sITCGQbJykIdX2O4p
O+ruli92DSgvBAoas61ctv6frGMMP5k5ZQtYNtDOLLlc9VCYEjAeuiabRRx7lx+ODol49lKQ4BEr
lvrmSvqeolHFenkTRlaLrq+u4e/iBjhtYBqoLfjI9gs1ArfTzUJtvfI2asCCdQTcRe6ZwQuVAGyg
r6+nuXMTsezrZqHVjsCG4yEnHtra/Us6h78acm+FLkM+cS2DNzWaZkv9vg6MT7FITqHcZbSQzVi6
3q9yesLwXbXtkBKLujAYunSHjzzxMg3nxpywFfkW/YE5HNZMpeTfkW5Lb868uWnmHO5a2iaWRQV7
vfToSSU151/39+bMxr/xBSbKR4ILXOo2nGeYBMBZgUgqCZPavx/BHS59NNv0S5Dvum+9g68DywnB
HV//U0As/jaOoh1Ny4KGrW8Rrd7b2cMQGrn7Pykml5vE8u6g1AKpTrysh0DWU3VLqjJCiwZG1uAs
wEajVAg+5wnVQHcn2k/Vvua1uijOJS08ReiYnp1jkYvVTEfbzf34wFBY7IqB7a0d6YPxWHcXiVdr
vCD6VtXUOwL/+m6oRtXK3W31/Gby+bz5mCssEDgVs1s/geudJDr8f1KzScqp1ULa7fh4VuBJqCAi
XnyblkNv6XO1Z0ArxOBAKqEBFCwB0pvU3ERl+FhaxAtiQkpg3WYLYED6YHFC1w4Ayq/ARJOqunyE
61UVmCTkbPwj+S72YA+JCznS4sddcd05Ewoa6NNdCC78aIb6l3gEzeNNhgOcUtotTUu40dXeHYNg
Mt/GQh+SlQI3uMOtB5+kM2Q70TyA54qRhPfsmbGzO53RxNHVz5QQKb1dz/xhrge2VljdB/bs8W6u
6Lyftv+Hw5T4h+TleiM2folw/YUa4SiGXMJ8iEJxGDYNSek6q/Gl3xlMADo0d5p6b2woKD65EYKk
l0j8bvce3hn0YmXHf4My7FOJtB4aulwWSCXeYIDmvnQU+TDIejaJXdcnT5Ip4rSOabY5cnOgT9BQ
k1Xr8zuLeYt/O/lNpdvApCLTfk/e9gmIamDqH4gY5OQsfdY1vQOxEdygo5ErEmO9aUAs3iMINYlM
2xgTpXSk8IyBJo2HK0JuvUrwK0zF/dXx+8lyu/t1cMhPkfrlY20//HBMp36yAFjdL9sDXkVveQeD
DakhaZJsCdqYxHqHH2pN9oJfAXbudyYpMAGV0klid+F+QXLWDn5iCR0u3AEU3opVnAI46xT2Ef0h
pSoSvMAkvwwApCeCERZT1rUmI5gSEVlLxHSiWLEeA2bYj5GQ0SZ04HPQ8BAaIc8NJ5Jh8M3bwmvZ
CcKKae9JPQwJf6XELudFhRpc6UOpDlHZDAL5sLIKWooh027BHYRdf5FMAU9rWNZoGPzh/MYu/T9R
5M9wwZxP1OGhsgOEhGDK04w72zXRCSddvHAvrezgkBEzJNwr7uGV61ZeQ2OkKFQmC01slPeKGcr1
LFUZlNzScFd8LzvqbgOXvNOb4GsXpMLf9+DpYNmwkm4ljJA0M6eVnXRZWmvaLJ/eyIdjxSr1pV4V
ztOnLc+8A4xITGh8Xtxf64Syci01Y2pNN4lpA8rqU1yEEsa+A1YnHAEuDZ6jy3sSyh0Pkk75epvc
8HZ1l18D70VXrjmdl5/3jbjZWPPW2HkOTF1Gzmv7+knbD0v7RDeAYVhx4UbVyYN73iqKEgsRBpRv
NYo9HYLvkVc+omzVm/B4n4Zu8UWaPkNSNna6OUkLzKdZX6PTj/D8Iea1WI677Mxb64rMYfhmB6XA
B6PTz6Ra8Ry+wLZcIiJpLv/rjzb71crbuWcvGwlIACyklrHCpw==
`protect end_protected
