--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
jSlsPL8yV3gY2LPmylA0A6l3f4nXuZ9bf9xYpGE4u8V9PCXmVEYpq9OPunBROvk/D/CS9QvZ/FWZ
QsZqhDYR01InAcof6j4cBWVIHsqO6gZqWpDlHrThlq8h/wvFJIUP1MM8JY+zT/S5wVdDsrNE9W3B
hzjyw4xcbPNJvH2JHdmune/hQi89SOuFLlAdbdd0OPPhOk9R3Wf/uX3rdvXRzohNwfskFqPQHToe
l81846EHUBUDBAL1lkUR53vhBmyln+2/mlRs/dlc+G7alHwQkSKq/jFlUDnEZWYd9nKEo6yLjOYh
avvSeKa57LX/qflDDhURFNhXuIStSGtyIntCOA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="7qC1iOjyeJxUr+MB9yKpK6jI14ITAtdE1GvAK9FrXps="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
ebLthU3byWCGDc4xwm+i/5JnttV/6ueSHWUJMbmbLrtpUtDUrXAt/omHqfzdEdeZ/0znTf9eu636
LVagS9NTANho+Uh5md77czCCKwpMb+2CWOlU4jxGzcdR9tJOHkarwzFMs8HuE6Ly/n+AzzVhsYIN
aAbJfh+GjpE9Uno+DQIepHWvhVBlsixrLQb8rjh/9EGfV1RtvuuCTZQWMcjaq1Ixmxc0J3f7jViL
IlrdXIipSAuq4wvh143Id/VE55VUeUhFemkr6Wcx7BTGNN1FCypqzLWZwPsBBSDfA0uHhooYXcu5
l9wZvUwtNkMQD2sRnItLPnnhZ6W0jASvkCedFg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="klbEYiSYKSE0IbZhW+oM7ythPFJFzd2OkilO36DfmOQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10576)
`protect data_block
qLQ+DsV8q2+O6ow+pZJbRUt3CF0ScVHRpWvnx8C0YcRgjXFK0xaHq/Iz5lgt5YaSZeTxaL53gz7J
En/MKKOUYZQ5YA9GeYvl7Q2Vm4CgjWhSrYSWPGJV6V6fiymV8fue76fP7Bfmp+OFK3sNTsy6Rjb4
1XqsBB2EGAb5J1XP8wadCtLTL5/fWWESyZ/C35c3Ws7g23NppWknEGUR5/eApIMdU5bJoJRl0VHS
euwFVoQY2maGgQN9S+5g6YOOKZVf5+zrxhj7yqOAmlksZePaVt9IX1A5G8+yKKeJXIi12ZM7RIZ/
0ePYJMY4DGItZBc6CVawczwvEX/rmPCMGfwRe2liravQYeT3gT0HAYKWVpi0cugF1pidz3XKvybV
2TbAUuBaS40/YcMGEDyvsSbDYpf6eLh+BwHMscqGCRUIEFJGa/n5AH6z8fkLugCCUWckimbiTRXa
jxDYmhGqdPgBND6FbSES/aB7JFEwkpJtA/IyljiIaL3F3zWQZbCAqOUoldJQGLdWJ+tUrgLTeN18
J3xF/UivrWWcW4o31nJ8gGAifW1MJSXWj1n4Mzc+wMhVmgzOFAKmgArtWhov6DABPfH7A4dTgYap
EWapOPSDSuTjN4jCXQcnIsEXgf4bfwWLNKcgd0idaCNYFdp/VbHBaLMqTRtPPq/VZQkohKiDYZuS
d93Qn1DgKZz9Ms3p2f6GiBdmekLjJ04CfAKTh5nPNrJp0q9y6pYw0lZsTKBzyoOYp9JTLmtcWRmB
JjJwc8sCgpdr86b9mlvIWjIBRlTaa68YjIBUoqbraFGIZ8D/9Xoyurv71EUiRY0BtXh271Pu+VC7
Phu1gk/LLH5yfDv9/FzPGtTnLSMB1kM0gkFilK8UDk34zGZai05FZUunUDCEGVPsnIrA+JbqcLw1
jNK9O0dCShwyFMpK/buslzWQqBOq5Y2EIPQB0Gl73FdOSmxwOQ6PiSbVTO4SvYyw6uJxjeF++nTa
vfmBkkVqguyzapoqus8DlSwtRzZIjSV98jBoYDa+J1uabKsbmiZSgXqWw117mJwKNhttjYqW5wug
tU2XzMGK1d+n64MLEv658s9ubXdDagN/7YJFW0oZbODoqu/bjp1iNG0uMinS+/Jv99Q1sF51vIFR
GGDEGXjTya4y8uR8CEq5Rmar1IllmzArE+liixdTJ0C2qGB2nSLlBke1j0+8eTdRzDWAZ7zEbmj4
XbG9wwjpMnGJ9jMTE31v9dbaviGIyi54TMCKGqh6MYYSjzeMXhQDRy/bB7sUZ/MydifDhsmYmQaF
aoQBQLEQQ9yVNli6AIM3xqE2/UXZfZw4Th0oxhtytzONkdC8tvZaqdEVSqd8peN7RuwjgWcThoq7
dtCzuxp/geDVLHhcb+ovuccpnJbC6JO2N7xG+jKqdci4EaHVPm8yKWMUMrjg/4FO72UU3Ou9L2T9
3pCBZ5ctWyaN+5kidbyOt0jM3ge5rcv3D5ev49ssBuitafPuHvg5d/5zx3oqjfpux7XNnv0dZhCP
AOYMrTA1qirGQPxqUs1eVtv5sG6qGuE2gKHLzF8IkRi/ubplGO3x51Sa4nn/inrRFTlH9pa6vTeg
GyszfVvBLtWet8c91G0kh+HUk2vIexQLKnHtT/1XMGU2S15766zdjqgUgynLNI70VopIVVKrW2j9
yZHsau11tQBtpDL07o6CyzKjIHRxRvwNTW0WuV8mi6t8p32oosNotKulCs3LybOrS2WidqbSb9FD
f/cSx+00QJbmMItLVkgMQEnI0ZYr/AolkTE02J6NcrhegmOlyxQLxaZfM7mdDpjz7uziKXRGq6/X
nZ75CLCQbY5t7aicboEebvyQb95FRa5EJ9TEftq4jp0apeigzvIO2BYZNhD2WtCFTsfWrX221EDf
4bkrpNVYDhxVViL8qLsIaoE+Oyz7Q4OM/2UD0ZOk5ibXnP59oONwkd2TjIKJ9+EHYg6PHW5DAomC
OmnQaIh1IhaWHSEfXmnS/sPOxCcsYQgILkYnkd7/8XyR2vHtGn98Lq9o9G98fVYa4smgoDU9UC6Q
Otq/otqk2HIQQ/E3vS3UqFLlTojiHL+px6eywFTixJlpS0EtYAwhBpdmOpqD3rw6xjC8G1BRRDio
6Gwpz5+O33he9J1/fvJfQXPYXZPhqZCc2/JwqyVPJMP/eXSfkRpG5gIO38CFGLXA564Y0tJNfzM0
lU2k366/nHAG3nLJmRb6HrhPI/uhgIGU22uo3UqksiHs+r+27PP+7C7rkT2QCAYRE25XBSdnjGYH
WzRtqY3fbmV4Z43gVAXijwaiJ15gOl7TWkpWOSvQBVSRhkIs5k8IR8x/Shm8yaQ/w6SXRRI7Msmj
rCcylPOYXY1LBdk+P+rtQ3KnL9zMgbMnYAON5mh/3hOcooDjh0umAq3XFVMIeEQ17HpFcTSPELAR
QU8JVcl++PboJzQmFV9knjnOK6ny+mL45xNcy9BI3sktHv+pATwvc0StJXEsBR1W9PFJz/dv8llP
1lvBwEfm/jpv+Ckh5+c58zNCGK3k1rHRsus8t7cWA/2eV2Zv+zRsDCt/Yn+1pbTi1kxtpQDQWi1c
PJREr+Llmc+87db4XFPcKq6S281X1wFHcbQKDBl7Jxd6sBq3nM4nc4deQn4ZgopadCABHRwhRe7c
3Yt330CUEJRFeu6xzT4gMH3Pxf7hIqd8/W87Cs3cSU0nqG4y/JGJLB2krbf4KxORyE6s04FKchTQ
MjkxedZm3GB3hKh0kEIjoFAOIc6Yuh3CzZVNTx4NWFGxKFQy4g34td8/BhnTXLTFtSMybB2UGuPD
23x6PdijgzI1hZz7PWWBzg9eJEYGXd8tvliOz7vbw/uXNanPci7dLeA8v7V5l1+W38vtIlBWwimH
k3w0ZPY1ZmOZShfLBKFMQHaDKM44QEFJxnnWllyS4i9rU/rX2qdcBvXN+oP6avciuwAub9EaEshb
CcyMQr48z6wvQefx+o7CocKecHgdoHmj1HWB8dQ0C+0O9racwN2gTNiGH6lgG7ugcaTfKd4qjqNX
f5P4vkzS1rF9Q6PPKY7Rtbh55bD0Nsv20YObpPBh/nnII7rDkRDU6rWc+dIr1Bq9Ou/ggkmkoTyi
dj3G/kLCWJ5M1zxTOh03iYrAVDk32dHAmVd6MQBnDCl86IXZITUR+qw+2g5fEf3UdhHuLWAE2E25
sVN5sDio/K0GwuIw73zAVbwP33tvfz3kz26Sa6p/SF6oZK1Yem21AQr/Fi8iTcLGHzGWhFp+tIY0
xUQSVpKySZWox8qwy7YrqJILF6rLF7TBUgCwuQ7HLLHLXj0qqDGFVcRbM3Z7P9ZsQBA//F8Pp24o
oOO7JaGEc/VSpNzCa/972V6BNhnsEZNgKNKuOFSts3K7+EhBmbm+4+5UWIPIdhsc+IQbJwuTQ6rT
SEMWjHTXp2ZePqQIrynCnQxbUWMpwoWbXvvxL2nGEM83O5bbd0VU5+ZOn5/1NQCoXa1aHQfZWROU
kfasnS5nydjZ2UHZKSbfP4bMHwit6Bv8XC87cPJJinYj05ntUNRmMN0eYPCjI4ZiksUvzeSjaWWh
mIGLg7w8lXR7Lx/NZaxCPNo20D9YI8W6f2lsMoeFxfffxCbNi9HziuCDb7hc+Ty50WcqyKUOt81w
KUlfDrbJQHK1BmqZYZpW/3JwSbct31veZ/0UtyrAg3HL3L8iGBExUn3JF0IgBDk3TJ/GWT8X4INp
Rtoh6a0q83meVRm1QCpyT29+0LMofrcM3R0ewXgSqijG3N02L6rXqsMoClk/3doa06db1upcC+q9
DrsVETsd0XwfINnvWue+R0f0WF/Jq8QZVwC0Z3AnqdsYvh86s9LKGO/LcXanLMivLpXpmO6Ti6kh
lw0hBma2JsteOE5BT2I4BserAS2DgRPt9k82NJnyaIsaPV6x81/xIjSlnMQaL+BD4lxgV6BdmOFC
K4goZhZWLxLQY4FbjfG5ebEMoVJ4XOjvgL/gRYZPuNKeOxeuvU6gDUgD3JVFS+B213bkBCSOd7MR
moBhJqmlQWd8Ul36CzV7sFzdGr6c8Dq7I3mFZW0d+gTXXy28d8XJ6T5sZXLI0amq+t5TMXqOPZ7a
BYUJJ2Tm66do4EwUUtqRrf4ZVyKZzBlHUifhOXeIAJRGszXwlicFVvynf6zdt7sOjN9e2qFuSQSs
9Z8IaQhE8u8u778S09fJDIBSR4iq8XICHP8aatiJmlJ0dx1yZzeARhFpeOOGZWTOa/svcfVilGcy
cz2kL0hedjPDFAEAsxUv7u/hLwI3fTlZJU6pZgjBHTz+YTPDzjZhj+cBMo6Plnk9gcogNaDmJutq
Du7h7So2qRhKTgUFtv1OrHPxL40lyXY4XIPkWQQW8+g048OaEpbIKyjqfmDyOQ+F+cDgsxlO9Z+Q
8bOkuJjGYvB735vl3NzqgFNv81QcWrMFCCr3TG4X+WtWfxguOJZL4juvB6ewLPL/goqHE3DK+XkX
UTjHiq44oh7YTMbqkHrK65c5acgwM/YQTRyMgyJwFCHkstELnKtWgrc97P1Q7zfGHjvqbl/Ppkna
tP56hdDodi12G2l7bkoIkICu6So22axCyTg78GwRoyFLY7KCj4al1ooiGQpxOA0r1imwgFMafzrz
lWMgpJJUjuvujj1pSas6nvg+iGcM4GZ3J/ky3qJ/2GFc/JJ4dLTHguGoxbproLbxdU5nThuUPZwm
Hyu1WWp/eDs6pISpZzQ3y5E0jraS3n8w4Mf8qHsAI/V0MR/dljcnzDhdcIhuAaeqKm5y3vPtQg+T
GR436XUqepsxCYhomeiXYpGmBG+7fmLSYBvypi3wiZAiKOxYzmwKHQR6s/vpgQbticmXRWc8thYL
8bquURvq8EWwh1CG6K2R1TeXBxjOx7iM/HnRrGND/KM5xh5WKyueMBCUOLgXWxycOqpVddEkZ3fn
hMN0dbTRzyXsqHOs1Amml2YKYBR+w4pFgDrue7UmX389o13cVDvAcCV14WSZh06TBFvOb7f2J8aH
rMzrbV4FigSEyqlfa794YzRnY6G8QV6wonTmTGlIT4DxCUyiO7Om5hnLyOuLVOCp0QJMv6vnzycf
ibVfYdJnjQUz+ah8clP4nUxQJc23ifVYuWWDljCXo6TMrJ3LxsNDua3Y9nrwLgItxHgzPDE2uEWu
ol1XL/g5Q+fz/919bsEq6zMhI4RgOPO2OnpFOnVtwDIA6Y3xlJMK/If/lBNz3oZiIdb6lQ9SxmzN
Q5NU7dTACN+xZZlawIJwdiHF1HearASpauCAl8rCKht+6XwInTOfdlEV57IHuxbFCurI0OJEnpMX
5U9bywBvCh9353NIxBNeNOIl9rs/TS1lC/G4eCOpkr+tLl7RjBzNaS3yUhB7KC3A8v6SmLxtMvm6
sf93piIkZbp6KYXtpdAdgOepTWTp3KOGjOb63KoO1OZrLNAWxuOPDUwRPtW4XyIBcuGCsrHUXjou
XCwTBcwu6koVDUg44i9oLQ9BnZNe+pVZF6yXqTXh0c2mYhcuZDol5xTnRAx8AoHd2wBzClACILfG
nRluuY/cpPg/TQ3HXCKCE936AftGwTxSF8Ry34EBEiKOI/AaoFqkTc1+4cjHyrLXrBEY/y4jsH9C
JTHJAVKsJ1jlgeKBtLVMgTBrNmsdSbLev5flG2u04ppYbXkBChZAT/g+FT4Vfsa9/N6hQ+wjARNM
hqgpjW5w6VxvbeaOpohE1umfiArCdRdT57usZh8zwwafs5fY3RTPXDjv3DHu+dbBZ68fR4XOlTBA
RcLI8FmTjExWTeDr/PnwX30nOLZ0dvb3COv9Ac0UUYOn8JQqM2+V8Q9Pj4Y1TJGBS5RHxDYdZyhj
ezcrxNWaUxvNMCzlZgXS8S2tWnxk/qhoBXVlmC95v90fFcrrNGJiedR5Q2U7wi/JINbniPkpVQGQ
nBV73jRMdRf2O8sCK5sp2vbimZ6+OXD9BkORV2tQLae04r1jfgLyOtq8IPHFO926dZsOxOvINB/7
rwYpBaZmNXRJR4Qf9n8NPAtCsoSS8Cf38jDfoP3zQjguQbnVA33wSXikkQ3nLLJr3TrKwnOnApKk
nK1K014yQX8Qu/lESeWQRI9UVlSk3Gqiy/gdStGt8vf2sAu/LwPWvDil/Nps5F9qhAakByPrVi/w
3zK+iLr3S06HQQp5qgEDCg49d6m6XZxd359swx4IbETrIvYlIjFYvwvXs6UAtGWoRHZVYWSeu+vu
n5dJaudqp0HsYjDLI8vqWPnVqmHKbKdByoT7ndXIen1V662VdoLmOeIQ8b2wKeJvWOnZmgQ81HnG
qKqOpOl5tD4ljjLH318gq07YqCSkjX4YK03jswtB60X8hfonO+dAkTe5AzIOUOUD+dkH/D0lygfq
8WoMN4cx48OCAQrWYQhSyVwbHWLdY7AEkVzdUBVOqfLdPNoZSXM432fGC5wamkiTLkstOrnoVyiV
M4QRHk2H0XCGi/PG14cSpCEMUvPM/BsPC7i36vo/KxPJAp8QXKEZELLxgqujdIQgPsjb8t6MV0Mk
qW3obKmZuVlnQq4H/13sLl2kdOPPlQCLPeXnH99rbZaFv+X5so6Gc1pSFlKjhsiPR4n+BvNGAoXw
X8a2OSkfcto49o+9pC/jZA0lB/P96E7BLqYlPy5cpXfIOElyr5sgbmRPPlz7eOQ+1ayXGqpcSU0/
Jw2tp+Y1kUNhYRKeG0g8xmWpgTYfYq7nS7CBOAHRzhsrWWIOpEDtkGUw6969mZu6tgonsTzlcvXp
IMg1H8/fUSf+D03BAFz1eP8iJWnSjl/7uf38zlnUVeIskvRqrvs675bVOdS9mGevTb7QBzIio6RH
ReeId6iejZFQvAU7irCtM4cbyMhxpzjEGQUTlzeWfRB87EP0ECuoPxm4USPwWyMUzTRL2CPvz2/y
DfgoPookOJLDoPW3IJ3L2GHuFAZwZwGpvU9gBMvV98cvTz4AZjLivvgdoYKw7i7/kpSux64uTALo
+8AxhnXgn0AFCEteNfgm4luNTzuVP+A4hoVy530i+M3apM0k6o4b7Qolr4Ugn5+4XNwsS7XKr3l2
jjwYAPtNCi6/ORYRkvv86uCjYCXkPL2EgaTtRfXaMKagkS0HX27fY39+C+4fz0qXovSLjxCXChFj
oetWKexOITOQbhwrY/KhJbjepxKxKLYsah2wnT7t8S9lxNPJMhPZm1eIEIHhW3KVPVeMke9s5mxN
sJnMdpXQVc3oWUvS0JPo8tpA1pyHGhfmk2Rzyu6VGK7LzvUteNxJp42paJnnkxTygFEbPrKzwp9b
x1IBl1ZJVwsrwfj1WX3hDBx/1OX5BktRQcig2lIhIBQZJRQSA45kJ9d1jDrse55Vw+V4SikZ+pr8
FNIVlkxMl6m1vnYtSbd3Jei0iXAS1VcKegfvjM7TreaphEcgqrzpDs+NQKdZVh865tw3icGhJr4V
TO4k0SvnHLlkZTXLZFHrIQYNUTbJHb19lvzkzWHUKFhJyX7+P3OhvO94BkTQz6kgCXVfTa1nkUCe
5x5VDGdR9tRR9uoxq5VqeZLDv8S9sY0CSURytZo4vj1YkgLrtneZ/AoKhN/Lyqk6Z2oRDOC4tbBF
Dm587QClY8wv8y8bmU23iuPZCCA7o2ZqDWQjlc5hDmSIKNCTR9kg8CZFqM5IF4AjLPd4mqCbG529
SteU3XwMbN5vV0pSr8GETj53qBNsxFnpWRJHMcEe02Zvsy7fVnVyRHD8HcwodEWkV2wrHAJNUUZD
F/pxPA/72ZB9p7u6SdwXf53tECTh968TfP38xxZrq20tCuS1xrAxmB7dfQ94htnOz2uUq060sw8N
fwRGNj4f/DmF1K6PeX+t/QUigTh78aN9JSVoH0BIqDD5WTE+5jwEU2lyRZGYycRyEdpuab203dU7
0blk8fHcbFUyCOIVM4UibU7d04JCAF8h7B8mb61Kt2m6UENkF621aOEwlAJVXmZ/uRez5nWckUEE
jWtdIO/DFQpoPnVVxm1qJLce0XtiISu+jIND36X2ThUGXQg/Wi/qr3ZEK2SnXlG/mi0dUA7Of4MT
o7Dlm5hP5GE7P/74AjA4jXOA/8zwRh61NcdVhZScNqNHnKEIxo8RkRBQYvCn5gmTq/0lbfOQ+Etw
I2PRDAZH62eBXKmDgHdNpNItC2+IyScD725F0CsILLYAkbN4KrTbB5FhSKdOm9Pfbo+PWrK373Bg
WsFvlKfoMwjloaeCdvvJOEnd+WYoiA8JOFmJelCnx1urcj1dV//cMwSjU0T07JRByjbfqvtSTcQv
YVuOVAoYNC+I0XR9mnDO5HwP834M4EoARyyAtdupZ6mONBJw0TbEAOdBVq3elqDuakSGPCeSW5X/
432oOPJdPRnYR9KM1J2skGnilsIIoQo66lbt2XECd41EbbtAVBGLHdju1UpkmaTlt5Bt4ANhWeGE
hyIKndXn8lq9jIdu2rdagr/lnmpEkIUtJCxWkuYLfz9m8WHo6t1K2nicyJN4BDcesNvisZNbVm0O
j7+hsWg6UaOUDdV+B41adTASrs4bH+76FrSaoY7Rdpc+a6TkuPZoSrwdlAKMEZ/l4l1AEY1DueLq
Zfnhx0Z/S1DdzR+dFgYLKo/b/mR3T2+XpSZLyq10xnkIMQNGMal9xaHSKEEu8lYdkA//OK8XeHT/
bURn+tGHYKhlQz5LZvhTMVrl07d59ocyP1tMzkS0Uxp/5CnYRcPNPIkzvMda1IOF1+hjloEzXRff
9T302Ivtlg/LIasNE9BWoB9RG2o7QQFFyuda0p48IxG9EKUKwuFiW6mNqWcbdEjdJxEJcUCnvkDj
mpIFoOyoOXzKP83d2DL9FTP7EW/wV/XsJPVrybwfbgYO8X3QPM2Q8qwEKwylJe8XsrvD6qMOAKOm
09hRLR1nr4hyBU1v4E/GzrKuy/Q0UXhtQnyOINp422O3Z8YpU++1NQM4jSZZgzpIMOFsyUyj98AR
a+Lt8xmwLR0pWwNq9qZYL6qF/T2NCqUNXo6u+uUF/TSyayBqQJvKLU821tbMZjnCBaNbknMXwbTs
RIFO2nrCf5Lz1cszMZsDpx75/HCPeW6GLBd7efC72HpHiU9GfwfS43eDbh3+aVCW1YaqjTM+uLs/
Ur/6TCXRs/IwWm/fiQ/VF5nDRK9e2ABSTgXXjkinl5YVhfLY7HfoVdRIWjQUeKOxsjhPJA94eDVb
ixEtUvTLfGvF6HZdPrZFMB/u/qlf4gGG6lkiUZs5iuxX0T+bfwMS0VGtEd/TbNYQ0n6K860XqMIO
L2TP/ZnWW7Pc5ASUyczAWPnPhhpdRZBjQz4RryTxWRviaX+kY28YYt886Y1FPiqQI7y/TPZa2inZ
M6hWiG/UZiAejacnHjH2oja+m2QCR/GBYupoB2o0gnDPqA7cjdbA7QmarK0v87HmNI5AGe7osBQP
VoMlb8zNbqD40ttmexmdEd/XVOnT6UIeMqXKxzGoNB2UI4kPjbiS6hcRlOZY3pHaPrRW1J92eqOH
NQvyL9wv5ivgIwrQOYDm2RzeRGEDQeAr3Tt8pC5y2lL9xI0rTWu+7Y2SRo4IGSNVP8UzUpfCb1et
W+6lBEQvPwqMDg+N4jzne/qFrObQdpYiLpI12sixBIZHZtn1wPhmUfHvl/dgw50zF8kgXq/OrMF9
q7fj95VPfVnIfWpm3BDFn9qcmu+u56zPPrGyP4Lqs4540gG0j0lHRHx6hGWz8VpEloCXlGcKo/uB
o/3Baok5bvnDcifZioa+81SG3hXFUtPLPLYlqsQgREKAhYUli4RB7JDDJXRK5Ykm+VKtPaxF6wpC
ClBWvfusdyLDUnr8Z3ILA7qiSrEu1g6m5pPdn8UvkyUvQi+bB9wWIsEGmEVtTIpNN3iChZzm8sx7
/sC2Q34YHFqAAGyhST6hEXdDXYscUOtMI6cE0SY0k2xx7LuLNGqpljzwhtQTim7a8spwH4j85hpk
hgVfYk6BZo+ptvUxDtTxuO8xOnBi3P3eWZ28JkN9JytLxJ/DvDYr4VS7Afn3mwYE8TS8cifBeWW9
sIrn0Q8vUu2gNWG5FWbYKqEt2Rvn5i7qfnpWWzCpZSz6nOGK+IBDqFdOtFvmfmBn2orlO4P62xXq
+3m0G3QI1BTkIn6vcSVEM5AfHMFG5XPPluGEQKNk60tiVLYmMOyRnT0kqHOGzLT+TxuK+IkYqbsr
6E/c1xsE/2cYXWHq8VuBqT8/WlC/mfJw+pHpcq51eP66hEezOlHU/RVkZU3TqbW//3SVhdtiD2/9
fK/O9ips9QItEP3C4nXBTT82B1bSPkPINbdYnLeEsF+Fb7q5zkXPCqKywHm8sdoe9Jki08YlsbgA
MBMnpkR2lfV0Ocl5Ugb4mE0kXbQO60IEd2sKkl8jSIykRD7y5Pql28cAj7kvCc1z2PEenDdoqF7j
AiaHcQqypaD6I7c3KESSYOqGIupJIjKzAFuL0a7WAQ7BoL7ppop1NTWOo6MuLjQJa+OORSln0c9I
31/zAUYSbeZo71snPNbR4K13ip6TFmsfB15b9DktH9PYkHXgpyDrrVIHlvGtGMyeh02Q8NgcJq9Z
prGRGFOzDHm6BH8Hlge32aqsU9nhM/oKbar5VfNjMGZM6v5NkljW9jcVz38Wq6VrKAEztIaV0MhG
qtzYWCi6wE7X7sw+EYXwFqNEtySVDm65HBxC6W9piA+NhXHU4g4sojRVcRw7lOjlx+AJ8QpqNaan
EfUwxtHfU7dmEK1h7zHTHYqEbzPoD4TumjNoHczYW91/EtfxRc4ZBhULrrGgmFpFu8dd5WCcURho
JYIMMSqwIPUOMR5ccAE2L+n3bRtzEWAIDjNmNJBAzkCyT1MsuKpMFDnVtzAX/TmVhdG2E4HtQl1v
H3ayiSYwKEjZEJLtlS8h/1Qbpkbq7LvefAwQVlnF02hz3dsnJSatwnv8L9rU+WuVK0OKBj3tbuK8
P8xAyxCsHUeS8izAzn+3350fLNVF+a+mzt8M3Go+ej4pMsbBjkpopuUlHYb/OOoVJ/VbceA20Q32
DLeigherXchwFqaXS1Vbb3OcNjs6kOHTNqfRw2ylXhzgO9Dsw9p5eLGJuINPyRKOAjN7UT0LKSWi
zTaMOVM1LcxtY9RTsxjJ/ZnuDfgx7ydP3m2ZY6kzSSL1JcWj45yMZYWCkZ2QDt2CXnoCroLpJxep
5DRnGg1hM5T2SL+OWo7xUqqMbfTP2nJ+sPJI/osIEo4ArI6e82SE+xFFE+S5CL/SBXmNcJmcDF+e
kM9n9IZxOA52N1KiGYtNqTf8iKOYTt2HEA8bzueCfcV06/nJY+9RvAghxw9EjE+kx1Eqqjc42A4F
4gx1aklQSnr8yohXIL6ozK7h5Pn6XuDE1Un9LmQW+IivBv6KjpVEHswIKwpOMPmH9C6OQrfex9xv
BrZti8hHYRVCf1d+WXYrGZsyeeTb1zGG3fz+b+q1BmdEZ2E1y8lVP1g82YS23Wk6PHNuayNwLjx8
Pgq+tokM/UK1K+AY9tBzTcZYZvigqD9x+l7EOseon/trU3RCJQPvEvCny3k6rInQtG5QCKsG0bxc
k4zx1asNbRCBYPCA4xNPavGX3D+oi5tj7k5FtJ4osJE1M9ry79sAYD5ButcjOfTDTNTX0f3gH6FG
I+5yJJfYO/EUNVZe2DOuTlN5YsPZUqPCSwoiqilsZKqutimEmw4TE8wlAkSzEK10e52hmKD7dZFS
lMTZGkP+46fbredZwuYLSwUojw4kD7v1cwvIRHvhz4I7EK+nb4eoimw3P7htGJ6iKMIZphlk9a6z
qmI84MGyr08qIx4H6yeQBCPbPrRYeItsSb5zxsYBbgImGYiSvarYy+ZAFde50VJJZW6v6iW8wH3W
SiEBGyLzSy5qtEVP/b2upmE7cs4mbZME5eTvbOJcDtbf+yoIjJyrHKOCBn3DWUa92eJyOgBTn/Dt
nPE7ZXKg//Lri+OLCwQ6ZXqWd7Fbi1qbr8Z5bchoKJhu5O/+EDdymiCnqzpIQ1yJEZy9L4fVxbJb
mY4GHGa7+GfoGPmd9/Hq4ySbKuuwQ+B24sq7T6dWvyHQltAZLW+ac/AoX6k+xI0lwErS+4oeZW83
Y6xSybPmme1ANEEcx5UXMFezzzqSiU/r8jy9gUZnbczc1sbCxB3bemC9dbNXwCBdukCC2tObYRcO
c7cWtNKKuTPlw00/WSoJzauAlo+oxBTP0QG0Ma6yay+GmbOkqiesg2vbT9OjfhvEDj5nzzOmX2aa
EkEGpv0HM1m/rFIv/9KL6hBqpPheeIev0Iz5gwV5q//jnmwL1Sz0GbPPIky4UNgNb9ZJeRG5tWlh
tx8QvHXJtJXIxNaIyzQj9ixIR72s1ivJ66Zmii7/7dk5SNFCo4fwpoG37kqAWA+qrChUrP+mp9d0
WOcyOLZ/YEp8vZMaK9yfYTrTgNlZA5/p5vOFD/e8sTWdR8uW/GLKQ18ineQ88ExOlfWA8ObF8Zcr
fjFH/mkWVGL7ymRBU+iVGMUkGOaS0cJDdY+Sd7qq1paNNuR3dqpMN3NmRAqch6E8F2tCfsZUcc8x
0LVN2mqMNiwgiTUVWAZBNw9NiTwWbv8h4+vWswcCJw/rdBL4my1fvlxrAeTb8xHToLbeV0p/4Y96
O2qh2HIgqk1SroPsmi8C7pmthb01wcskdrfUr/sdlGsYlvpqsXIllquci7EZt/OsqimDt8alx+Dn
9w1n04HqZy/QzLuhuGM6E7Ol531YGDQI6gK2zMPCHopIqJxb2AYJhlMw4TnKnqs2a2hsglFMOJxT
UmrTk1cxA32pUmxizmoE2jKhN+W+LSK15/6agNEZvmtNQ/24XJb+xZZMtFtjwLQPXewALS4cu8TL
OGNeYT3HmEBjkLqMZT1kte5z0FbEqe6SAsb1YaNnXvWdeZn8Zz5KAX+8iukEiNTDCZRVtBKo+MrA
NGU29ygvthJuSWiy8pxcxOUc7zHrLLNWywiizVCfg6RZvjPkfaBsvxmtgAf/Ewk/qSWk0d4Sge7T
HS+UOzkOrKHJOvyNgR6ef5LH9OapAPzLPHTH+iPm9wErTv5zLqfq4eVR2rDobWAvXL/q6FhyE0nV
HzSxadTt55NAQeP8WCy3GAwBgwPI7YFMzJOIsJHWHvt6FCocj37WpGtDEswLmr8KmcOOErUauOrw
ArmNx5hsRyg/AIJZDWzJJk/AjZso+y1kuiC0cl2sRRUS2zKhq1yhJv/ZccHbmBiysDsZZHl502vV
rFK2sLY1Eh/x3q2gGpFG+QrKbZQDxixo/UtLUmHrXBcktMytcb6GKRI6vaaKC3kO+DCSCgcIpkUI
VwmQdpKUTzzmVpeB3sfqRrvih3erOpcvfEhclYVqWXBxCJrTcg0NmNTMxFmz+bmYDT6PyXdND8R3
vGcPf0nPjdf4IMENV6D4gv3eGfdR4Pblihuw1sF7JiimmOOzdY4gigR+l8jXIY+4xzvTFeW7gOJj
BNtm2MICKISzavR8kxJhHz6XvL0fCiTDVeGB1MTo2aqwxRwThUERf6zf7/fsTfD6g5a34qTKbJ+T
7imdBslu02Wl3dH50yxu6HymzUcgVA2QLNU1eeHQB4x4f2pZJqXXWWTR/FHyoWAjkHDa9OCx98no
aqQ/fRjBn6nnG+AA8+K9gBlZwLM8r3nY7O9SkizWeF1q54mExRutx9hqrtiMRJqfH7YZtJs24SVZ
DcYPa5O5tJODE7q1/V/TrsXTzLtF4dLSD/C2IMaZ5SQRvIAv4w1UnbS1RU7K/CTPlgzPcUWOpGkB
bDedgli4t0e8CeKqU4TgAWcK7wWhH4qRaabAbuTyKlX6Or7uZGgS33DTfqHHigr4gEA9xAuEDhWt
daI5xQfq9Ok90bS3g9U+nftvaCaMrwlflrbY+8+WILmz1AdJYQGDUefh8vnUx5vzgtKIuFJmjWVM
iJ8SoylPZ2Ag2Z97Yua1ys9n+1fRyCZ1RFxJjlS2uH0T+b8OvqCgxULKmwknKHiZeZstLDFAf6lG
KXNAYldhSOULy9JsvCicvzPwTxux9gNvSjf57bNFVdK0xQT749IRVwLfWp53tX59U8zo6/J5J28N
jAXBoclabINvb4eIdKKMhVaQHD/d+LDUClk5M2/Z/g==
`protect end_protected
