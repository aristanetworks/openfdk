--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
FRqhk0THtAvwBm5YICNyzygUKxgrb6iO/5Xms1UO2fHwl1XH3z9mhCbLSw5MXnE56NEcRjWwhFwE
BZlX0SWL2jxb30SRW6175BXfgJtsGqeIJjwljQ+dIkYI90to5kKP/2KRjyyfufnuTypWLeK+dpcs
VFJ29+CpEgJFWllUAN/dXyk9F+qMPNXeSUb1e2p6FfKULaY+Z2bVmBotUrXvI4tdj+QPXvtNwbpw
0Zl+qaYqXSHx904w+/tVLSpfaH17hSmsaNonAUYplt0TcGhhl0X/wIDGXmf8+aWB84OR3FUfDtF3
ueIK1GLozVOIjL556erx7RMlEVjQfSDxBDcM5w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="NFEfQ6PIOwYAZnVb8zHYrA5ekDCpOZpYLJwWi0jSUuE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
U3XBOY4VmcIdFVQb3ANneoRTuHblCmJNAq9fg06Gw7RdqO4hi8t2y+3a3nWWzsyUO7vKtL32VG4V
qopAC2j92B8JXiKKj7pj+OgQqGA55e9qOCrhL72czkNUSGEJddP+dEpjwk7spd3Arm4U5v5qXJkr
TsAM92Dhg2TAxk6ZAeu9HXlzxYoKKCwS+lzMbygER/raaqc+m9d0YNBl7949h7hcb5EqursRJtTH
gaGPdVk5DSBcTxayCI/OKbiwvis27kIpFfi0h0V1nHwA9ngEPEeOE8ujWwmyszSe3UPyCqS328RY
Qi3RUmVEnzEU9QWAbNvreLuTW7ZGuHSEgpKizQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="eaepvvigEjImBIr3Me9m8Wq1Q+z7+I5YJzKAA2VMttc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2640)
`protect data_block
WpCw/Enq4ShwpKQ18lh9pm0SY1nGdJrN4UppIliJ0vcjVnwc4Ig7ntz2oeeuchLpejlryWQha/l9
Rekl/lfePqHhXXa6SbWICHMGtfcXVahvINdUPSUvGZSf+weRvUna7UP4o9uskVhPRZJepbDwaOCv
men+UgbOGtjW+sdb+C6KjerSVInC8JawqPJiSm2vN6yOHxeyZSDc65jvHAaNa+RJDvnaxayzbT2j
39cjF5HFdkbPj8v4xYakkrB7KtqOYC5qlWRCTS21afj/nl8IR1qeBfyoUBFE7i5jHm9T5iZ9jp4R
aOQG+Em/F3UsS1vnq2X4rqjM6Zlj2VaBD6dBBRfrOCxrYZTDNR6+r8xtGvEuOevytImWimUOIbMa
kLUEXQF1YTcCjRxLlMBAndkSWEZtWCTEVCXEB2upiCi7YBj+FgL+nDpUjUaoTa1RDoufvnIOk+mf
CQfjzmmSRIIAPpHDFFB3TDaGYiI/PAwXEPMpMcWWCJiM7NzoPazkOHp2G5I+Lb7ipX9nCCY2F5gP
oGB+OIEDzmm9gj6C1mSft0G6zw2jTzUtp6pnKCyIzONeouh3EhbdwTwV0Yq60Ak4dzPpOkIuCuxf
Unm2UMCudSwW92glOYRl45oZNur9kYhKe386Hfs2FrJRRpAPcKLI87CUx7gTO62HU85cx1zUIs99
1LeRAN8BJ2AKE/URr/tVSxGm7uZzYXBVOFNBBFiBARrKMAaOFVYAk3WMMWs6S2ZthuIq1VoXzS7J
eDaJu2eo8oB7PfpVeiZJ3Zz5dO5DTqUG0J1/Bir75qYEkI0g3xbBbC4PHyvjH2YGovni0WhNSvtC
NZ9TZ2CbiM80qqAhllE0ndBR1Z61xmHy9AMAXz5HD1IcgBUmbNUveRhP/HHfjmjG2k6SMUI8aYSN
I7XMk50OqqUd7RPQ6hL6IhzSJYwE1MDztDxCtNzw9EQ/yzI7GKTNR24P1+WBjlzXGp8GztXBWWTj
fod5ssaxnr40zZU617C/LcYuYHQSBy49hk1l0ZkrBiDbphnfU2PG607QgsllTJsMc9r2wDLTtc16
ieEpAaqec2BpyTb1q8KEuh1fdV4fKfjNlOmuh6z0u/mUamMobqqyNfVcp+/lEpfedrbw7NG74FZy
a777krscGfgGSpbkMgp8/TdId8yGrEGzvgZV8X5c2kxTGQKCvPksKgMGtfhikbsyvfYJEm+kDu8i
i2MccNxqOGUOqO6NDooQkAeQKqVLMgBefchqFPIIOb0WGkvwtzxScfszIp11DgSGnA+pRNxeVxKb
jjUsggmSKJxSrSmow8/ewCE+a2YCVa0ld5FrkX0kove9+SiMOKv3m43AFkiVuRvsFzrL4JzHsc/m
txAkpZR0YKRE9cJYjOkfWF6pSyZNBjhyUNfZOWW++RlOiYq7PSkgf2P/GqzAsNHwUFjyBCgRTRgQ
J/HdeyI78ggpos/Og5pZPFDVVR5YCjgfU73nC3Dw6AjgnfAkZ9UdCXVAprZjFGSVJlnhOeY/p+k+
JYc3t+yw+aRKLA2HFzL7bSZMPpMcRC+4ippTJ99qip6MSlUewNjE7RFpZH1lSJ4chqlaoKMZt9wE
6YtcMLiZxdyu2fx1Bkuqx+tj0vWQxBIwbwL20AXEZT7rrsKGGjmtVeqNQvWMiMppjAvnYTQnJkzk
qvNPmB9FRItYyUzOuKchqO2Y8pEfd0SvaqiZ6oklVnqiwX9o4rN9Uq6jbXlqR+wj1JL3y2KbWejz
Go8y/y4iC/an0zlaZ+IRe/cB6yuUa8myHaFccyhP2UEPlLuqvhC+TWEH4Y45Fsw3dNjjRdVFH3y3
gDP6VOGsaOQhzDxMjqSkejegfKh+O3Zdj1wdIGMcrJ2PFM4eyMLFzP0EJairkDcHnaN2tIGvvQWZ
1AToW8kXSmEhNd3ICvBhHiUNsbX66qIM/wAVYd/ZnwHr3NRUMfDkiaragcnzEl3Qb3ZduZHTYLTr
enQ14dxwvcBdcRfQJpX4O1ULHaYOzp+OY2Y7x8UC0yCDmODlgkLFuFQufF6pe+zk78Y0d7D9wloe
LktbVL5HJKQk26usuaB2Aj+rngzFV7R2JYbPM7T67TmLagpMuQiz+JLhiTXPlYWfP217Eu4ee2Mv
cQlmZnHC+lz3Z/5nhkMfeQTmqxdM5oFLK3WsTJbQYyusSLaiKt9XNVpuXu8Z4h9oOAZa4X2O4NrH
cTWPlqFi1mrGUielXddQqqGDJHaIorC8M1Hh+TXOT+MvGyZECbDqxgl/PxGAmOFXvLUb82YVBSs7
iumHGB88dLH6fLmkxdu93b9CIwwSWwIQmN0czipYHVXSB6ZbIEF/K0KCF7sQZ97V1nKLn82ggRBX
isVNU/qeTUqkTqAXi1rQRUe3v/OLnUymrJwaKNmvNFgSVw3LFxGiiJXiYOm8xqhwDqphHz5K4sWE
HxtZPj9YfNWr0OjEC/4roxmtNq0kyoqcknFzLJhbC/c42tio+JDAKdb8kPyivZ/6j1SvbM1CPqLk
B5At0Kv5P7qcnk3mdVVUjq6qo1JXxTyi8y44G2ayrBCDyWX2qvUQ7piHQdn3NAoMkj7jUTdp+RmP
Y81ywETWgXJ7dhKx01C/WNbwHvXIZ/HQK7VvmWQffkTQvw7ZNS/oNsrV0Qx1aBlrmyVAD/Q4GYW0
APeTL+XtCERohvg8rN0KUJe99x7cebC9pzf2zTn/7t3PwofMUZ1fJuGYmIUTy19bu3BFAL5cQPyj
jM1/yN1MTDSC/ZaorHzt5gEGWsImjnYxqheo7mnNWNXByxP/E+pLm1Hw5oQHg8d74n7gER4/ToT6
sax2lcbaUdBPtNLeJTn3VaxqL0mAL1J0yKeVX3K1YRY/BymPqkHFNTjiUfj5R2T9XCLhsXFbldyZ
TZXMsnjSlmM252DZ50Gmgj5tUU47ulEj3xOLG4GkVXbmOQ4KxMnOSyJWvWThRrQrMfTpZa3JKs5O
VlYPAj6yMc96va9jdIP8+HFHLPq4VMjyeT82V0dXcoL3uoOa5b6p59kNomhaz+ULsG7mmXw1dXDZ
X3G9ZMMfW1lBUXLb+zfiAx0vQc6WxVLOc8RS2zfsgGcZ3N2R6unLs7xVev+vSh+6dEM1ulq+GIWg
pSqOnXrhaID7xLtOraU4IBJih7j4ksYk5FKeDD2zmbHnesTKxOfiV77AQ9OPvkfCQDksChTi3le6
iiMMvqxt2X40QjIbszZQ3HrDJOvCcuxUpffscgf+OB9Hx8PKT6EjVeEnMpHsdg3wvunbSze03W67
pDVBc2JD20VgMaJ6Yt9huKYg7f7ghGzNu0NW8X+4v8pDSk4EZgKYtSJdEBx4u3v8pbMQ11EIwJTc
obGncHPV1q1iDj0xtN8va2PMNWwrdmoz8Hc668BkUpqvVaLfGZZTSkJykz3EBlMaO3Cige0ksUFI
nUuOSRrQaiHkLh1h5ox0xWZPPA3Sclg5y4iN6LHR7hBBWE1LOiE6AzbSmeiQFEfCbUDF8QAyiy1c
LJ3cM3z44PlvQHsXgr6bgBM3
`protect end_protected
