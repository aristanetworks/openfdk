--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
PXHchyXrnUVxEqiQWEitPjPJ1WUkn/KzZyt6qJ017dDesBxCR6ubkNjzEsrD56j0aPZ1flU/kzS8
kArblJDJZqT8yxAkorgGdFwUfgqPcC+mOug3x+n5F1SGHQXvCulVCUs4PZPzdTiJ9nbFQN/FspbJ
gnh2KjR1Hi0/rh8XV5DR2Mhp9s3+w7bB/zXe4u+8uxtWV7AXPiomXQve6W74Qjb93mKTnsTWjzXD
/VWyPakoeaaFwUUo2HsTV2aoeCFVnq4R4BSibpx7BHMXPBP3vI/b9eabGmnM6T+vsOm3oIlhjAt9
uf9mm4jTIc5Mq1Fbn4mlWW9jAsTDG+l24Upl4g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="I9FghhNiPrvIYGkPh97Czc3o4DMdx0/YP8gCrpk76cA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
ItwlaqObFe5tCQKWFOOEaxLy6QaHSADq12PEzY7UbB2msdcqDArSupJmi605CjY4nX4QaNZP6S6Y
sh/SNMvv/pLsOFKppB9DErflDgUKKovDwLDjEjsDSxGauOVI43poBWTRJyIiGc+4kHnFpd2/dFwE
h+dH0XALrL51onVbkMxVpcF0+9GVWV9mGu8uZ2dNjA5X0DNUG50+bJ40kzoBrZdFPd6WmOvn5xKW
1mM0z5Hmrz4tAoR49hiZjFmQjx7BVfzjqXidRBGJaGWExMnysGU8R8aHBOO1rOGM2MOyLF+b5lJv
w8lUnllZcst3sGlOBjQ5BzfyFb4JMHeR8bUiCw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="tgOU8R5YiNENaeJ/dXr9R19vYlZP8N/UcaY1VsMqjro="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22064)
`protect data_block
uYMioZ5ru5VMf/ypYQc2SJvB5AzqqtlCsnbEvwJlcC/VI4QvjTQQKJNLrkKQJfvMUgw+cxJj3jpW
SvD2JidxWvzyiSy/FPSG236sx6gYAspDJ78z/M2MLcSW7jNDY60O0fq9LmzEtx62Aii4ACJIoVSG
D8voBi2iXmCrLtrTbvtPNb50e0fphmVyonF1RL29Ll9YAukTSqm4i7KmQVo+PgE6Wyz6l819H/iG
AKOjiOMBljz9FNCFvWPWNGYwjc6kUN9RiTK6kDmQqy0odRfw9tswntgaFfrwK1r0330huyFUIp5h
FrAgk4y8+2nUEZohu2BlAl2uiY01eTeh1gUoLoHI+KVKT8GIT9ZWCZsxm+kY17PSkwDF8LsUWeKj
B+CTKSvnTOYNAesa3dD/JGepujSTCzCmdiC1L9w5cER07ljy/2pCybdXkxZzpYiyk5p/jEWyvOI1
befCAlxX7yRSsNlKkbEFx1OqM/nvPfubOpLEs1Njf/eY1NTbo28nyyIk9vDDrWGskPTmeLBqYyAr
isQ1EGEp9LDvTsOFQEXC25xCx01/v+8LDMv6u8KMw2U4rIOWGQvhAlGlDYPwEMS2jAosHOCXxvZF
SfdYppZJhDg14Ue7YkcTh9bYy0rRJoR4qiI0NP64hUik5xGo3uHmBAE/ZhJQxky7u69fsXZGeHmg
k+8xiXht97R0tc9Wci5oiS402oVgQGFfWMrSKNOc5O4qA78f7iYHOCP28MJLYKLTGPtQtqp5Jc5U
NXdMmiWQU/i6D4TF9PYB6Ku17LiUgHpzaG67kywzXxzGgFP/ppJl8ABdUDz1MWPXzBq6+6SHV/Hp
nV1yJQevedxy5MvoQh/d2jClpHRS6atuqY42CAcl96W9N2MfFgIAJwS8lA8+mLXp6nM61EZRihZh
0m0hAUFe84RdId4YPXzyTElFzCqCE1VxqdVzX7pNxaAFj1y5dYj81OdJywyDh/1P+K0zKa5xsaa0
kBKu59uJMP1UrJTiV9QaGwj6gHnS4Y38aIYlyerhokzH+Zy6kjhjqTL8gRov3DqQ8Mz6BB/jmTT8
JTiemd+5cfwHOM38djM2ZR70o2T44FB5fSDojBxC2COIK/Jc89r8LqYDzedzRoj4CQr9YZhhuB6q
J+19Omgrmh0fCJzqrcc+tDY6KKlIcZ/isHb2OZybJ916shX1FZZp4wsS5mg6ccKDfR9z7+tnvOnr
uYiyUlQJu476EXvgZ1t6eCBUSCmw1asOWfJYlvICGtYuaQCOevK/R7O0FebFlZEl9F0HL/QcO2aX
+zHUhea4ZGHMIlEJ2pvGHJ0RWRSIQ/aEvgkQAJS/o8OIWHEaZ93FFGY5h6e7HdAvge/XtGNXK8e7
vvLYz+NIGgD2DKJFCpGEs4OX7whyMl0XnbTvMDr8xvVrRHo9QbgVpXdvjNnOI0Gcv3D8HFiJWapN
ENDiZGhGBoFbjfKohdzCPWMomLJt00ZkqEwemFvqrbRCI1EpUWfc1ZrZOYfFS0/nb9Nasj9ZcXuG
REMbFg1nWDYCwOLrEKmxksYingQaXymtoroz7bZxABCGZn+7JKyQZQn0VbdhzA6WQ353cAJmFJ0K
zvnqwoDXsl8hX0VxR76bs1XnODgd14CM4vWJ7DgHO22+YbVlkyNbAbrawSwNWt9KkG7UkfJCRZrf
kynWS5VcjcekBcNIC8wTGTnmXin5y62nPzILRSeBvbhjsqTGNJ96Y/RZC1WKhUWhMg4VEmfg445C
xt4pYM7EA7r9HvLFRzT149j7lwr33Zeug+G7IZ4GDR02+Xre/LIyggDybpfGPY0uVxP7LbzQdxXM
HKumMe5woJHYe7YQDE7EvbMBbbCi6jO4hKE993J/Q5g9sKUkRtGfLahysWRUiCmX5Bf+JVpT5sgt
TskrgLE+8tEVWZ05mA0W/XrAvPnrw5MzEq0SVqtqFUmAwNJNA9tsLyDOrBAONw4p4ighs7qcF4Jl
xBzUpNNo2ozg4KEyX4C60fvOB5SahzY1CI1bAKrseRzHchpbQeXCiNgEzOCecB0xm2gSuCiZic+q
a+Nbi4UlENBpvFQnDUx9/K2fYSPuk3G6+RrRdffKKxUstrIgC9QmTPNMjrnvLfI7Li6ndYwAhiVO
Lv5uhTKMeaG0dw/kif857SS3Rnk5X68YoRx6VpVjrFNpZjCFCSQli4Cggl3TIHUP8zbbPpAGh//b
oQG6WdftQWPBF8KM060BJMICTMdXanJPO4h+9f6kTvANEkvsd5ZJkUF0hLYlHRmoXrPVZUu9wRM5
jXSzFblZpAjfHn8QKbrLY5uCt/++1JWjZ1oR7GTMDKtlhyWPNVYUhzJyD21UPiXwmFCjgbFqdgqB
dtNs5bfGbEIlEfCvbV8O8GJ70meZw4aEYEKrJmGCn3LWZIuu60v1attpms7K/lbrca9SjyJ0/t8Q
fz811i+jYtY9q0UMqDrjvEtWeYMr7sYBbJ6KGEhTE4TRfseBtafaOX2BRE1jTqJCedsqQy/vSeIH
Rnj6npDcyJU7V3XHoyJ4H+wc2lhvmIznY21cpcmWhte/lattPkOx70LpiGZiohvPO1p4rXcdUM/D
sh8FLHEot8v+ruP6zx/BT/B6inLbjrVowofLiQwAwTawumA1IxKKLlVxdOC1kUr69ekuc9n/o/aw
R41uKgrcfyBppELAJzakjgziAJ50YVuIUXY9GfKIJDEWHlNHDDqOLdfDuc3tODc/dAsE0I6f8AaC
ic6V4iZ29ISJ980nst09OIMrHkFdcuv+64LKNPA9Ps5A0F8rxIjfbRu6ZEkg1b2eGEqohqKFkjY7
3/pzuuDzexAtXyJmlGJ0X2RcuhuQbIyZTGayy5gX9fxQMo/uqp+psYdaTFX9QB+pze0xB27X38Zf
OMVXLkmKs887Gcv+TFLhtmhLpYrYkOjEIiwtHs2kuHmd4fhDc10p9x2zFJyutiEkf3r/0kn5cjCc
Z8xioy88D9cJWtlPTO8oWYaHkh0Lyeg+syNdszq+euLug4uOXMn1LBqcdKKz1uiO1OXb2DPJk/Sw
3Pz5KcKg1PCmvws+s/gsQokGb2YR+JX3bTWL62KLnPrONfZBa8uI7S0FVKbcjiZFl/6uDSjG75yD
dYnoQLRvWb8eG0hmqEIDDo7H1hXzs0nw7m667O1/lnJziFYIr4BQkvJGVXdvd/yBJivqruxkLhAe
X9ub9WyVYiBlEC1v2mQNdyWhhqWr8ft/oASUeiqnkkHOOSQDB6n4WGzyIGhQCfe3K4f32GBJQeA5
Tc8YAIJTbXe9uFJh+dtQCp9q6MVfp/qqP4IskGjfkxr8EGBo4I8cny8EUx5QN0MfKIgu1hL8noBl
aZ7oaJl61Ps0Na+tYfVsQ4uDJKJ2w+f1cfWz0rNQjBxOkRd/nMPmlqTy1wqmautdjBEgk8EqJhoS
/xMUZEab9EjoyeHB9sxb6ixDCuU5nZISXVhdXbtF3gdmXop1QT8NwXXVZSQ/LWpVLuQFQQKQQLex
ggxztkfD88DqpES6zUc3lJKTVl/VrNPihHZmXrKtVrfsyZFHMHzs297jcYT7Zv3nMMn6WYs6xtDQ
ZrXVtVXgvEyl7JePVxrxUI1Mq2O5D+YRqnatsiudiXF/PgmZfRU92kemmRuEEuwPs9kbjKGw60zq
dPjQuCdXPUuamqrAiHc+VVJsRUN6K8Eb2oT8XTxJii+RHmwZi1ZBFS6WdUlKtNmDO2o3bxunQZX7
cSa0Pu/3/SUm+SbskdNFQ/Utfr5oH9aBJKJcBSeRIbUfDzxErsLIsm2/nT2lO9YCouH6IlmkyJ1D
ii/DmkzsPFFp55RiJpGS/5vA9mhBVb/P9Ye7oR4fd2qX60ToztX1PLhJ/1IxWwOS086zbqTfeQ2+
Dt8s1Zuw+DbVHaVeA9pJ26rJ2ImiAhb/ZIXnZPXQ4DnD2Lc5xIZos+OCZ6Fj5b4MH9OAhtYBBy9/
QTNwGeR9A3Y2VoMZ14hKHcBkZm6l/uJ+C5k1E4p0LKs5IFMneJikbZ9QF6hyH+BuQ5pnrcuYMZRv
fjAVZa/Lt9OujPMrsr3PKi9dI3Aa9WR8cBfZn00F+BFXdmnlKvSH0iHVnFbqcW3sQleipqJr6Trc
CJY8ZbVlBhLyVTftsasJZcsk3fuUbmxMq4mqk64LwJjNd3aB4JHRMvbtapiQrih2kmMGoRGTTG/C
gBmk5P9zAvGVDlYm9MB62tzZ2+OZy61BI4i9l8rI0X5M3USh3xTNtr7m+ZcqDF46cdtAoGo5uoVG
pWYziDxCvOzziJyYEgmNXp6S640klmd9rCz/lU3t6FJc7QmF37CEF9rTflU/R+2vxM3KF+ou30H6
OsncfO75/oNCabZ35te6YTfy2f0GgTJ0tR5gTUal5+wBHpdp4bPaptP9QQfoUpfiMkzaeJtloqVo
u9YY5X5O/vC1Dv6U9Rn0vCzemhPMuUyA3uBbsTBjP05bgYBPazcOz4iysTvommZXlS3gSqU5nIum
91sBlPoiHFXCQFxh8mCdrfClhvnQmQZj8Cri1GYlvhHWwlBkkgSwxZAh4EGLgBcZQ4t5aDyoDfc6
Iry5UGwArXKEPO68d9SRzUQoJEco+hdfc47/7lTbBHj+ea5mUDWWSo63BxXG8kASauaCCEhN7FJS
iIN0N0W1tNk8wrAfC2bfCrMyVq+q8zQoVPP2C9aVeraYF7Koc2NgUpHHa0ArFK43lSjO/ChnkmxZ
t4hnVrGVmTGLBR92dXUlVZ0u9SHjgZ0uGfcqqgsAQv5tE63a6bLzGH2C98DT9dpFLpsC9X0Igy6h
LkdeI8oNC86XIOonFHKpp0I4SJD8dVQ8MyMzB8B0wau+7DBKV9wqeih14HK5JJ+gZzSMfzA9YspB
Cl3gVZYn9Fu2Zl59ulkTrn6W4Q+zxgmSExnphGPy8yaBC5eB12AXViMmF8j+ekTwf6ZRX82XUFed
Bg+5+bZJVvJ+je9b+0ynUoD6TNmRm0NwLh25MkXRtA+9F0MrRZxO79Desgr0Vk0Rf3Kp0vWc1OgE
wwXeQMnf+PJRQ/d8q+vBczcNBHP6vyRFcPNR57yN/SrPVWQ4B3oNGha35/rJg1B/7kh3HvEMWX5u
iE/n4tl9u6q4kAELgt2GikB3MXkA4hr0U2sZQS16Cr715jd+zBTeGEIQcUdB8DDNfiDWvM2BFXse
SWFPIYJLIqhqSQUmK/nCAmShdsFtnelCWm2MbQtFZW/hxMIo9KsZ9RNRY+tUQzILovvl9W4M42Mg
3s3KOUqEFbI+3On4jvTjlL1tGBR2iJZcDSKNea/lMfO7DtjIHeRMOv3uZpPljQnxAVHDxUlUMfyU
lrZPlQrlZRkErT6AHkZX9KIwF34YDNMD6Ij+1uOIOotndD5haXlC1gHDWHyUI6vnbxpyqnx9UDDu
IRiIqEC4TLNvydjgfZP2oP9Fdkr+FkU9j5uIKllYIVqsfikgVntwRR0FVQzCcEy58vLMP+PcL+py
7n7MDAIsWfQoaPsbL5cxTwp9yCDBPZpMfDCgSDnjOOnFy3RwPvn/oAE0jIXODsOALrXXJxnsamB0
vcdGkuLaK+ua9Peqm4dBvThKkeEMkDFQUmn6inr0Y4+y7zIj2nJdhrcl1mP6RzU60tlpX15g0s13
S0zoVqtOAS/RAqvG5cGXLJztPFFZWYMGHIyL1pSfB3JHfH+g3XGeotjfNCYUtQkRvgpJYSyB0SIs
Q/YF8oRuhaViPZck3+wFN9ELx+YVLLqWbgUpaq0UG/FQep+f32G9x/oYkOhQek9V9XxGJA54uSSA
UMDraUsve3lEZf4kQyMeT3M6hwei5Uz6vSwqXFpHylzJu6HUmB8uiMEKCtbLtQdE1ye5iBhFoiOQ
IJC9YIWIZEI/QpcJVJCyGQe5v2HEgkidmyCSP1N5xD3OcHcgw0aWvbSwHf6dW7WV87rLFpvu+8O+
dowfmF02PlIOJ7NaVRnuVgaYqJl6vEcpQwSDBo9BWCVnNDy0WbPfsXi5lYhhko97ZPy/GH6CYfHb
zaKAPUhWdx9lxf3J9C26HvJvpQODEvpbLGXtPg5BqmqGSu32GowK/VEjI7vFuQxDX3XpaFmqBm86
EPdK1bKa7SWH80h3/ja8J3FJQORumqCB3w2OsuXclE8nrIh9P1nZDKiFYW1kKKMcink6YE2MXGt6
Y/5O6qB1xkYqUeTSomtcuj6CGyIHc3hM9jkKyU27TC8OuYzrOftYIYReKc7qFafbmwWhTAztx4Q+
9sB3ksjZzTxAvKtI20lFIYei0SF0eit7GeTcj15XH0UW/T42dbKgrNNebl5hVr2rXaGYkoqu3kn7
WU9w3rcFSCv3YH6eA3cjRaMsM797m+eJQTJsf2bz16HXtL9uEOKuXvgzlPP16z8m89tosXCz1x9r
sAiHNulj3w6kOkRBSTqsj7IBszL/5LkWCcQUQiFIoMerhIFNhLj+jQI/qWDLsjIdSpfyyyQ60ZA+
xK3te9Tx4Pmzc79MuiscZ1UzaMNUidCnwn8emAxZClfzE6vgi8AgoLCTtM4X/lVtLlEItepaR04M
4f8BOxL79st1tLl7+qzX1K0WCAwnPrCpr+iRofrZlGs8MpjT2OorrmN7zwxP4YFhGcZIDFq9gSzK
C1nUk464pSXVCva1mtJdAuFOEHPq/Y12aBE9bGzdVITZx0byj4RlHyFC95zVw65/MVngaowiAjAe
1fwtQMwv8xXJYnuF5p7MeizoTuzJtHTG65QNinUrFawevaruU8oxBEfqIZVKeOH0XggPdJKS3vt+
D7cjxxTlDFVFTaQmFG5l3tlYfcRGI1/cqU7iwmo2LTvGIrrcRFLA/lFe7FavksUxkG/aXHV7t22P
X/abq1/FK4h5Ffa/E1INfhJoM1HLQ5lSUOf5Fj1CvvlIQc37J/ky7nB8oOj8BkXSpafA+wLmKzw/
duiAbm0sJxipVUcjqde9UAA69/WwPyHy9n7PBcxhXfdtzK+/+TZy+tmGKOake/b8pHCkc4c5WOtE
fOTxg3UKMWrOoh9HPDV7LbfMO2fJLrKAT91mh7xXSd+SePFimO8KrFZAq7TcihTd3zcLut8fw6Jy
wWExB836cD70dGyJgm06qpJk6RKaDC2LTss6NFlmUKNTlu0bO16qE01ddy9lkwIlYP2k4J78yIG2
Ghqkvzo3X47LbbRAsCdyb1tD7HLMHp8mLLWN5u/rGhsM+lg7lQGI4HKtNBqF2jV87FD2HJm/FDg0
aXU9mL0Kbff53w+qZZeYgbICiU/1LwPXe2cNUb/NO1K/u1QtFNHpqb5vKGp1cJe11u/hnuPsysnN
ZuWMhiB1iaChJRwoipmkqQPh5uxFMqz0Ea0UNhLaoGItY9JbVM3GoY8lf3ILtc8OT9U3Co0Wyrp/
45yROreEjH2o/QOcfb+Pa6RWeiZWTbqCgcnCo8RSJZistHB+HvL/aUTZVN+9FYGHmt1BgXfrCvPa
Hgd09F1dt7YrvXQ5cZhRuAuEbzhbKYj5xFHMazxMcTHKtdYcrAvk9gTZt+LTT6QVoBOI1X+1qlIF
BYO2I+C8To6C74fwVAvqCPo1nHoNDXBg50d1Wob/BdmecrcPXR71H0gWF2fQEWNPrZ6usH800r+K
HawShHOlRBts/fjZu1UJ2SmHydDU6Xz70A072k5FT3Y4G+89qWDKUUX29cbpaPUJOttFCP7k2tQk
WduVPbYsNmvQ4AlKn8z+Y7Mo3Uo6VQAvf7QDKhoPDMWeAFszRY1vMaPDPyAzZrYIdGGgqudh0RRG
nFGHQggria159IWXsEKGBuHJ/UokXgufZW2W2s0fCWj4rhmrCxeiXtR+8QTZmUrBhbpi3bwvI+4n
oK4z0yknMX2itg3+dUoTQHmwCircXDR5R5qkHSaN6q7CUozBrr8byYuIXkOSxtCRO7WfpItlsvFU
2zDRf9nEe9QDsShctab7WL8TQ7hZAlow92YousTp58nZOJWUgMS3DKqXVdKaF1Fr7vQeQVtyZOfU
1NmgoqzcifT6m5YYlegoQs4Gh5A9CFvfOU3DuqITnD9dTUEnvv8N98i6Ce4AUhAHRPSeKEKn0u+N
OpNgGe29ufj+Yh0U0X6OaD7ALyQaozI0K3/85b2MaJR7RTKoZgvdxHdSx33f7COeIsF0BFE6+kmx
Gk/fKBGKLfurHRkxggchZtQz24TPJVHJm4ykyqT7tc22i5pwyvHCEgX8CV7gqvFKGNpXkeIBIYUo
tKkKHwWzylLQ/i6T50icWWG7T1CVl80MCuo33H+EP3d7c0+GaUSHVTGDKsWRv4bDjTYA/xGFeroj
VrY9l5fWDtN+OnIymNzIa/lQ/ZanoosDq+5IjS4pg5d1x5Meyi9z3snIKCXf/zbPkSkVcKMtuAQf
UjVKFYZActtGYHtT9yyUyUrQTHzh/0sLIhVabz4sKW2pS/i5KbV5hqHoqFDbelZ8IiG2EiDg1LzW
TWDYw+B5eama+HB9rFIK3hxXaNkRUkc8pL5GLe3t5b8DcJ3mkQ2GerJinABH8EBKS42GYZdFPBh4
aCofRUv8GxhePdIXV59FF5LcSt4AZybgyv9miw6TZtvxQCJXRnte24kCduvCi0ve1EPdwHugjgAp
QovcEb+ogq+PxBPbfOtaO9kjzRRe4ArYX6i7wE88sKy5fu1CUBk0RAOBLy+sHLJP3eig4UdVsupD
y+q3fhQ3guxDT3UU412yPdbuZ+bMvq1ED60u22kYZq6OmeI02NsAHhzWaXk8zVYuMVJFSwuFKwkD
+2UOXFsUyoR1bJ/DKWBC/oYfWIjOfSnv/V58+qfBSskMaMvkmSwBBaLLhZtdixFNwzO9fZ6qAyxh
BtH5BuEXhmDMttMqxwPCAVqDXbFIduo2rtR6OtYhAg+cNc/VT5k/ibGLEgrNfiQ21VchrKe2yvVv
0OKT/m9PEagJfLASTRoWA9B5ioJm5MeGurb3MobkFOvt+U5sDFwOcibKkcuxXzUy6+x6PfMwiz2J
Rf3bssOGB4uEBXuUI6U8E+pW7Qie48jvReqDjGNnRJxMiHFC0neilgwpx8vIidw0A2yud8K/+k48
UsWK1cD8S3kuWpx6+oYUnQdHq4HpObIodIlbHioVyLDuPfrPA0NQ6e1eNwMLkDoRLP1YE6WkzuY+
YoTJIN5JXL5dcpt5kP/2Y1ds46o6vgWVwMXxB0oDb6z7TNv1Ub7WneiFGq3NIoikJupGBtyxZ/bG
wumPrwSb51mX6DBk9ok5yFmkMGLuEMX1OcP+hRqZAGiHXIXyHgo3CJ8DefCM4vuTvgnRWk5S9EcT
D0OXXMvif0btjRaeyhUhS1c+kuLps/okydwL3+EMrTW3KfHIggbcUJhuRnJR/CxBiAR4rg4jEJ+I
TwJEFoOAPz88qlDnDvjthaIKCmu9CAIkv0sROSY6m0vvMrITZo/09FM87Aq3OATxMCYX2a4b0r3+
kVjv2Q5cTVOwj6X0HNDc6YqVI76LNo4WST2oM8Msggw6PRq6PPIyqPj904am1dSOblaaYyUhqvsf
bHBIcboaflTMK+2/91OFPezbvxokna0l5n5Ur6BTbw6zR2X1H0BMughLvTLWNJbXYaWVs5FgvWPa
FfNQ0FIdRAQryD95DQXbkA6KPcJcxrw+Voq7zt60QdAeCwN6ejAWUC9d8tRdcArgOknrML/dNNjz
uY1o4zvEp9Vo22/qn/ZaxKkfg/ryGptxrRQ9ozhQMYWrPB5uqcT1RFcKkIf4+rFsMo96kPcbfXYQ
CQ548TeqBeTs0KrYUdr4GAEfdYAAHzlRKyzjoueEQ4wKGLJ8tnnSZkGIysvfyMZ1UbKylCg3ywgX
kvmhrYudMKJkKAAm+vn/+qQjc1mum14VGQ54lOozQCoXxfvg2Ye6zkjQIxCPYGwRVebigOs+kRYQ
gA1KQS84U29CdcF3RTAqiJAvIlVCCcCfZHuJE+YHrVOAYaWUMr86ufFimycIjGoKZHRT/xfUyshG
ck8K/zZeEEY5vLPQWkQViPGWEDf8PvafapFhVc6RLh4hGygYPE6jOSbBWybuwKUCLVUls1zHBzO8
bUlEz+ic/nsyxGdHdfKhQtyKT7y7FFPzVGEGvnxrjwBXYe6++9gZ9iArbj+UfHeDi+flmBU4xz3a
izb6gLxZUhCCq5RDpkgwhH+cXTK/hGPWI26WBrMskqRJIRP/QHsHtzlQoXHrngutuGq4gL8wbuKn
VK3KtgPutHj3mMeuLG3DU+xrtAo5lMWaMQ7NgzBGOt2qanIRe7TAxR67Wqrc8LHVkBHB+mGodkLt
eEYpKYMycOgs/3cBDVaPV0eEwK4k8fA6B0cj4ojtq0IwyWTy1mCfj27Pnr+ytubLwm0/g7CgEVIQ
Owm6lUHy7m54od/Qxe/dnG7SSayB8XjQYssSV3FQNUHB98IRpMOoYYjpmLe6gFJF/F8YBllrqqP0
oBsHpHUHNCd4S+D/VeyZ+O0ShIVbV5wmOo9WZX3t40AdxsX2O10SuLuLI4Ib0IpKfBjJ/do8+Yfw
S+05V2rIgYuF1q2F/eXlTLRiLao1L1QX8U98zbmUEd9lhwAfp/+afF403P4FgIIEDwUIKaZAB9y6
REk7O5BPnHknC4dH6vb+gz6iLKsqzqeatPDnNes5NBZvDfSyEiG1VXmlE0ZSQ3ZEJGN8GW9pZ6nT
+Bo5vyFcrwpBaqS1i2NQIqqRpWpbOjjSVCb1hrF0ne5qTFrBOOjl6cs2S6yt0WpeB+TLw1LawLnv
QvgTmm0kP54Zz/z2WHOQ3MXQzaCsYp03aIqVl06ZSO5ZKGZbTXTF5JH4+zDVdUbB6tOPXAcmJoGo
WIiQaTYNwsa4MCvjarHHtsWZ0N4jWOJ9Jc14NQ6sQciW2k6usBeZERC+XOA4k/AOr+98oF/i8d6Q
zHSuLbTKezQUcEFYpgcGIrsPm2dAH+K1LeUJGhKtCIiF1SZa16pTpKsginkNS5SIbXbYYmOE3i86
EIp3sMTgxKtNmOf+XCw4P3ijMTghvrQBdC0budb7EkxHpeywiLhLffPX3FngbCFFv/MWL9TSPwfV
oyBRVCo5uGoJJ80bTAuDQ7uFoseWrxbG0nMp3z/9ZS609sWWLjicXTk3OGQrE+I0ZYFTXjV49iiY
OeswB+woCesKwIdGK/T/u2OZ4mJ9LWJA9twAiOM6Hx7VcoA22CVTo75azCgMBVx4C9ZeF59+ZaIy
x9fw/jlyc3Nc0kJONtjqC9fWoZB/KaZdjeipAUUwejatxRpxRsliY9SCk/H8oQgt/YyY0+Zw0jiK
ALu/yQiNlG3gBl98G+vrMwaVnAdH8B9Qh/O0IjZcz4WTUX7Md/qUiThy11ywuHeBZ3XJovAdJ5Jm
MfkRxacpJuW4pIpuOIkGsdvK0qqF0EsM8udXyfviJ4Mw+n7IXyRVItt/onMBfl9pBkRdkiqayOb/
CQFzzm6tdxDGIf0/i4YBGiYJRT2Kv/I6WBM7MKvPfXvgnvCvMZhLCLVo6xthf9f7n/GzabGcBnr8
lBbirYLkZrf5ruP6EDjtKGHuJPscqh8BsxOBaeUMIDBmwqLpfxxsyhR+GGcv/3LhlK0crVBAPHKy
V6AvXxe5huVQhAd72S1rxjBL85JS/Ze1MCMF2R8QE+iweoGfY1A4Z52sixRsiWvsQ9vKTWi1eYPd
9a4p6wXRc7PEi6+UD6Lx4eoMJbe/VyNc0BAvJKGEl159kPucH4Snf+0nzVNNWpFrfIpXsqJ74ah7
8L109rZwU0ybbtVvY7qSdTcUcaGzMeILq4Wk8zyyMGi7EihbAgZw06cXrIv6/1t7NUd6sBEtXo5+
0hUcwbUF12mtMeTEJ+edg1Zmpe1A0J97t3wZEJDBx/Rk9him93X24qcHPMxcyXv/aANLnmLQXvsQ
ZKaZCXAvwdMxEKdaVMwq5Kgze5X2pz0FeJB5KEHVdCf5sK2yp+9HQazD2wYo/QC0fZL2AsUHWeVO
f/KToCzbooLMIXMbCaqXY5iMqEfwWaVf9lpYGGt4WqEIh2dfkbpbPHQcEUbKIh1wMxB1jg92vvvT
rm6MsJy5GeOkBR1ZvLdq/CKv+z+0p1IPbvgmKxES5GTqPpQT6FCnG1WxoZTHS+E970silEqKOM2E
S3nooVArsjgs9kP8nxwZHUAgIc/vjgp9g6wj8DRtCJaw3qgk/Wv/sLoFiST1z7sbKIy78nHtO+ag
ynzUKIMp72OiCqMepo2tmACqfaUgGb03bKVYTwkz/p81slUcdnDxCql3axUZ1nMa3dywVRnckfO/
opcQwk1wTllooKv+dZsqaomGREyE7t21VvIgMHiDLHE4hD8uUezoRNKYtGZOg0LvHO5GYsZ5eMXD
Ry+ad+QwwYZLy+DgGMYUSlWIZG7z+NlO2pdGFZO6PpWz3cneO4qIZv9x6yNXd7XiJJrVMsMFeJTo
iy5G2/lTQrGOBzgcQQR83ihaP19aOrrWGt4++i66pCYMWJO+mzzRLqhdst8gvYHVHK1rE5HQonjm
+XPSeDFESJjoNfc25XBmyrB7e7f0KvkXGmXtM0FkUqtddxhhf1Mei9h4ifLoL6cgKtr0M7Pt+zyD
tPabMlJJhEc2/zc9mAdpRr5EQkJDlKT+/p2LEpB+nYXsj1x+EB1n/M1Caxzo5CyhcufXlKLJqIN5
ylaD/WRAKJFKXmKds3UCD8nUwqHn525fBS4/JO5CFofA18hDZSFUkdKdZEpR9CzWYBsf3YSKOGvJ
w+s0SY3xDsccE4ZdGwuTBmuhOSkdNTT5prlBvmula3CjFjdcz5Wjt0q5CBRPsozuBCga02FUUAom
7nlwMRjhjlAL1jGDMlk7fJ3vws3QcrXknSZ/bej21Al1bvt3AqCrb23FdkmQGM4VynlTQPOGu7+1
OqA3Btzs48+5vdvcNJSpz+UlG7UQdT0RxFYuZCxrjhIIzXYi8elPiRvFOLeYajA/9t3JqeBU/uXK
OnqzNGEmUWODVKsCalk2JSwmMg+NBgXv7WzEADj4NG7PLZe/v59o//Dsvo5LOkIk9KVoIKTgfTUI
9D2kxSAwnXeWekTAcdPGTDYmL6PNYrdbSGr7pDX9qSNmGQ8xfLkl4tm9XDMsDVTvpyXDYGAugvxN
i9NGn3/IMVvMDkkDRzeNCug9pXMiJbObKrjSooUtrvF9UJP1zH7K67qlNigGi/rUoVAvHmGi/JuJ
qew4Rzj/OFpw7km8I9hoq56e03j80V1sIMWsw2dFOWpRHqHUsuNJX/j45KozjpzlIGsvZv3/xeNj
3inOWiuw5cV+zvm0lbSez6/waLSxYW3n2KWXiXJm1WVwZy3KRmiRDmDSwVhYN5S/SpVRmWHESuls
geFuvsEhkWFq4MfdiXqyRHAUbn0BdTK+m/+0o/ibhdNbHYNV6CO01VeRqCEdAOvOBzNFSFbeyFBW
czyNkpI56dglaNyMpXm2uxcFNIINHnG+sheN2s03FleObwNb72MQXUsg7AFyPE1E3X93Z1VRNS22
Z/7g3xlrhHHyvC1iSKmWV8P9PNu8Xw7bIX6lhTrZsfr0wlYV510QNavYjcdef923HD6qvxhpZZw7
BwVK4yNpxVtCCJy+saR+WiRI6fGPs9DDkg4rdJ1kTNNr8ii8paM+2YO61LL+I/Nq4tCfkBLSKMyf
HPNTgrbdf8cDFDnXxJKrjKCSitO6gW0woreytEzVOTGuygeDs0Dybj2sUMRjQfDfo7BvYZN23BJ0
1Ym62LRkkwW+rG2zqYbEQuC5APu7BXTbCkcxzeXSdofyeRxPjuA5uI6laFZxO0VUj/1KgQKcux7L
/U6SNWBB6f+O23aZWixZguvNi279tv8/Hpntpp7OxjU+bHDRUwUSdpoDdaqomozcuFZ6lE8PD7sN
Voh4VKw7ntp1rN+Y9uVt0cghgr/fCTYDSnBCP4CuRPsYlX4eiTUv21rP+xO2QH7ikN87oltfNoy/
0iaHYbdqreo0tTTnhwnU04DdkMDXCXn0MOc7af4tTiTlNYjIvmW2fe6KKdeNFciW50JMnfyxZ1gz
II0yJl+lzB5zIUSjj8QXQrMVNbEmloBKeLDwC3GSTpetnCWb8E+gejzK/sLPNYAahQKkiVJMbteZ
JaO191iU5s7Hk0rolZbkhmb5AL5h/ewE4LpM/NweF9b+BZU1lfMkivzeT5/Ni14E28Gan78chISk
U6chb6kGbAr2OaPg9qEGlhkGZnMLmo6EhZcRbvW97LDKjsY4XF4fdZmQ3JliTiYp00AqXVPIX+gY
m+LzBpG8ZvEsnQnjrttuQhtn9nBHbQ40O891pvqn6i7N+0s3uXUSxIGjFJ03A9BmfXg2RtJffnRh
UlDzEIu7ETE0AKB+eYWTDqscrUGYWYOnCIcVOQ5ayuMRExctcUAqRqL/5VTM0ISIrutwexLewHbd
gdVRTzenMF7YpwHAssdgIhpYoyWRM/LRBH6W3UceCCJ80XwO/nbZEgpdx4RRLFMQbih5K37HACew
v0PjtLYhkg3bgjiYvF1aYiWD5x5ZG6z0qyEH0WiMboXT11iwb1UiuFr0TwIE0MExccxNIMfTKYCJ
psnov1i8Pi/vdvQS53j5McovYVal+/bOYzAJIB2WuR6z5h+3MfJxvpqUyYTj1xkAXj4yFQpNYsu6
OKfxuKYTlcidSsCCye8iV3Er1kfR1sPZy+c32/9d4S5yndoobvOt0tFTlWE8h+lPZnD/aY7Kz0Jl
zlXqt2tiyxMadbKZIJsr0R4mlpkkQP5vYc0/Ux124TWdeT7C8NUX1L7mk4RFEnuy3S6IBefUSI+D
OLEy2ZRBarRpwT8INYggeFuOt6IOKtjofXRibqArcv/P6uUOdo9+Ht025sE7ZcT/4N99dz0dUzK9
VCaTvM9cURQBN39MXTbw142MB3wUGehkVe7hI82QrBgOW0zpYwDrgsOilZJByT+9s69cFiLqzVo6
U55BDDtjoAeKrBYdnlkQ8RzEcfhmNgu58HBI7W+voNrVqUew37ZYhdaXrnA2Cfxr+Cq1lfZwjSu2
32BIXgXJ1BqwBAUkhomeVo53zqpXWvSTUzFevZto1gMgPMztWL8WPuFEEg2zWMwxdzISeDiGjUXZ
+NdDkQvpKVxlvNiQT/F2VIyk9ptaWwwW1hsWRbmWSzwaqcy0KFXFC8LEZmDHjMowpXlZZjXu3myR
+9XkQd/ffq3uopLsRw3056u007PdIrj8ndpiBm4Ef1MJVtN28FlakKFurZVyvBPiNmcoxo8EcArG
es0sTfcsodK+hG8qEk9qqfBZC5n+LM4+b4zJxAJyB8DQAF04J/NQloBQm8X9wmr9anByFPgsMhDh
6tknFfYRARgArec05gC1HXnw8dePvnh1XwfCyw7f8cVdeB+IgjicH5s8xCR9hdXmuYOLIYMzEUHu
zHJ7UQFxx4604xgjI2cZYOZejCS7JMDH51gHT5yM9WT6GQU3rgGOphMifo1bNMI+Zl2E+7tX1h0I
au5bHagItPr+qOSVN3QiyVTA4TgUOo2XmtybgaQBZj8MXwIhjrreS7WSUk7RhZMEjzIA1KJ9wPb7
8f4XGTvjHkbbJ7pi3eG1XX3N4nVROQUYik40SSdG9qEHS5eHePbpkho8d6swdKJggNjPaoBJ+gX/
Oh0HkbB8ss7XVWwJshbk0bxSgBEN4xUfAZWjIFlcZzL/j/hNi7jPzDdLmh8D/zUSG01PpuRTQdcT
g8qoqr4WfPASi5rc1OnN/ULBRFNefQXLLS6totrHb/YRQnuwS44Nx4/W88Q6x57mbMmdEge3TXxj
olFCcd5+49PNG/BE3jaabhaICwnq8U7+5bQTruwQtG+MnT1IIsZ+0ynuHYmn5IUm62hJxpaw5ynG
9lLy06XNymtaPrjfcu0QLFl9zoayV2LgVhOmeVRiRrUQYflY4sfzzvYt2jCJ1/KW6yZ5i4IxA69I
M+JMD6kgPGqs+woy6G6QxVyWaIKZLgY5OqolUKRM/1Gvsn4swf5zl5OFu0HfByPQ8W3iW5SDooUq
KQb1+QBKhwH//cc+OyD9f2z62nOyxzpaSBrLGps44Oizyq+Vif+TJDD7Vv98SjAvqi6bGbe6QJDF
/f9fYiD3YcBuT1KmOKQNrtcqMqG9y1F2UN22FGzN9Y6E0h18Xcz9hTqXWbUvJvYjovdEHt1oRUUt
JKlB9BGZQ29yx2MXsH/IZ4h5vR8JcK4PfFcSRMD7j/ZfCTNOyuEBsVcdrbZtcj5HcKG8PUqsyzv3
xvteOILR+FXN58Z7OfhrI2eeVUmHlZynl/umqIAKCZsBOtTGzdCgvyLRLas52lwfhA6SVIbzBu2n
8ZG5OI9dCOjcGqN+gArGWvGSAZ5fBRNWntcn9mR5E+q18DHj2k+UgVwWqWujK/o6YW3XhcDR2BlL
cGKNJgo4fZPpKlw9U+GvP0xIi5QIqiH9HnmYBvboDVuAMDIcuSbMkVsOO8U9JgxGBMty8f4MwFAB
+sERyf70m213JIqKZP3G6qzskQ1EsaJD30PV21A50qEVtuddCW99R59ZD7ReURrXxYsdiEQFphbu
eq0istfYOGzHVDOjHaICinyBV+tzZ2x4w+frBYNSWKY0imgVVEj/kQSpnlJcgvaxX2GLbN5uYWkM
zTB206vu9hyfuUmaC3vN2eAWSX43PYPAdhQF7EobOw6UlwUBlkGKOILyn4+FBFRhJHcqA1QBn7OR
alKYO9FyCmOwSnBktoaJFRmS7J0CDsYMKE8XRWRbTrxbB9PuxwPTSWuxWtcUt33PMka0VvwCzeDQ
ixSihcFMq2fYeLmwf0XoQHQJ/W7ojKCCPSkK27ybxCAqwz30iKPwywO7xtO6r0wxrr4Rw+p7MSXW
t7hwG7CCSxgpr27LX3OX5LXHGT23HhTTL2/+9t0x8gR3iUuX+yr970X0UBnga8aRCE9cD4Dxx9R0
FxMXWUxtfoQ5+pphF8VuYNvnroqkD6LZNE+Tf5y+fD6qOXjR2nwlwLQp1B3dhE1q41GdWz+u8c+/
MOVsKnaEH9IX/hlERTEoMkV7eo+aAW2EPeyW6ASEX+hHL6MoN5mp1l6s95hYNz1mkz50qq0VPXHU
swpuhJbs8/jpMx+awpCQ1BsJuVTN+8ks6OfoLCc59A7ac5V4aFe4YZ8l8pk4XtXtKhspVP36kseX
dQ6jSljhrgkSm3Avxr7a8jepQ39PNCy192SZRPFYitjTZQ610OR6emRtRMI7HainIcGs2kNIKhdc
XXSGuqTe9A30bzcRFFBQp+epOviYLaptUiYPwVlMmEmvuKQ5EH7PabB7NU/8VjEFO6kQjUpFkTD4
J8B15UToIQ4oT8PDwik5aWymDrMbfMLaGu18cE7hSm9KYT3gEbdmkq8DJ8g342BEKPA9rJEKvUWO
bYZNwAzfJq3Z/N75dVd+ulsokYO7JH6prmML130Ne9cPf1z8thTw+p5q0CywAQZBpthMrRUipPtX
WhsAcyeXq9H7oUFVUHa+9y6qmYppil114/k2lJy7cFpGipzKAM2MvGrHdxWgo3Rm6QhgFgyA8ru7
aa4D2AspKwwSt+Ac8H1mtOQhCT3kdxfF1Hr0vFRrBW+bqkeaZR8DHCAmIu0aIb8NKC1TuEuSRqVj
R0IwmTwevkLgYauR+4ZiqWx2sLutr+Gsn1TIaHwfaq4L5ADVG8wCvoRx3MR238hsgjOlru/TMsej
SX46lcwXSzSagq2doJtMoBRz2vGqeEiuwtANyRgnMOlBnaMNVci5NGIV0reGdG68znQAJqIrW4ZZ
02tElefBYyFQtNYZ89kAY1ydT2GKJYJwenyhDK2JWs+HyiIHNQcBIud7eMcqEU+hoMiAA2TTCPDh
7Ayv00PBKpsPWFRn3pIA36TMjxLYyS13KtnX8q5Tl8x8lXLNOwpYefOmvNkWls5ptLeeUejnixii
GacY0CuaRAU97Gk0Xh47lHlNDTT4T1bObsxhNv2qz5efaX8RqkmzTw4HicfIhi7A5cn8IWzqOZjh
+6ima9hX+APoCIoPmYHhWkTGOvULmyaY8xISRbMrSfWrOaDQFKV1ipD47QuYB764V7aDTvfTCqgM
ASKP87VftpaLhVDQG7sQK4tgJrsyxmzc2ompa+MmxNHTBW4MevP2skILqZ7Md5GbzG3jvQ88Vvrt
Wa+knPoW3q6REO7wQ1ikouJGfgNyHDmuLCftZqgX6A9PqWIJwo5JK8Z7WF3bfZOvcMejyDRxH+hA
c3klrP7nS3yD6JyhgRY0o53vRlVvLuJEX4CuOHGi/YMf0Qdep77oaTE5IuCMPat+4Wiae0L/fO8U
eAbJ29a/kaFnmXCt0QK/4hKfdHAXJwplf9fs/4EZgWwvyRQR+ynTFZySX2KmYHjYvfkaYqfGHe4V
XLmg5PxNhO+skcdLzSj5KYpBX21yrvRmvmk/27FjNlJ2a6DBfuMHhc1Jyz2xgC/8qY73X/VUIVnn
m7+zM/EXCxsSIauCxijbx5PfwB3HWAxzRyj2ERtlyBBJ7EFXR3vy8ZHSymNms9rBb0tr68lWhzGa
aGKWDBIsCKA/Y9kq/WfSn076RAAWNhOunSWZcp4d8KKdaL4gy8F11s+B98HbqkSdHLzvUxzJe7d9
LVGxCyyAJodVJz4eEUvPKmSjn9Zk9Cl49rKYAJEx1MgCiC46HnqQS7CmJ/+dofjv3mwt3vkDMKLo
bz/tJBEPJ7nqVBmEW3XrGNP2IeE+DpApCBYgIq1xQkhnq7C6465l5C5FpjbncRkRQZ+Gf42DCquy
IIFaDByM6HT4fICQ8ZscaeVqG6tn5m+naTT2YrvI4cRQ4h9Xy0VPgMPZvq0oOMFoU456I5SzZo8C
2IDGgYQnoIzGbePIKVkJBjTiwoYsZGVLefbtQ5usSxI3z3FW20GmAmqf9oLTLA1D77n8VnSutqBm
rGNVo34GlrRsPworlCWnXLH68rqcR7luKGOAmxQvf771weZ3fUNdk287ZxQd2pHaz2v2LaktN+Vv
DE5Yt33hbzQF93K0zzW9Nk8mBpbamY3cDxiGm9veoBtBI8IR9F7Pi9tjlfl9RX3DOUJWYDxIBgyk
1U1UZrnch3k8mojhqqOgfvfnbdy0a+O2Mme8bbJq/l2auxoRTFFpnUSrcry+c1zjpY78J9hjeSEh
sWDgofYw8tBMnEDq9aV6yIczLaH+nx3la/Twoax+eAGaORni8NNeP8Nx7v9toJT+WqWOeGvfZN2x
qz6CatkR6VBIJ14If6v/2s7PoNLJjt2JeOGryD7KhtJYeNSpFQIRCeiCJWCvyH4GwUsfaqYcSb0T
OSVhV4DN13OuqbtAG2R/x9CQrEj06ysJykWaG68F+XHpkha3rLzm0iv0nugwhwM6jv7YEqBY8Q7k
ZQzRDwCGPt1DBxCnRd8H9l/KDUKiUrCul/NXkaiggm/CKLDHCokHIf45I9AGT0MClrG2hGxYqaud
k6Cgvj/foO6m94jXrC1yhHSuR7V2QdaH6wsV89nEUYaJKRGMM5blxhReFGpsZL4fxb+yfoewacCC
LvWBPhMh2KgLCIu60JLyn4UVJiLbaP2407mkGxMqxsYyjF0wqV9ohqTDr/Ym2EtaeFtsB1sAEscr
F6Z+BTgbv0wqsCk/0rRclgzEid4np+n0y4O8DA4m274OdclOZWCxPo0JSeZ99tvjJXh+RJqxLIHd
NOi8X4i9jPJOaVLsyRT30N+etdMa0+olKpWg1Ja11PAyRbga4oHhYN8vhdgWHxlrkvllfTiGP/Z5
vFW/ZTsm72pCPQ51gVIsjr2ZdvIzVf9+azdnkw+B7JBZ23rDg9KisnqMya5+Tdlv9yuc/ftpNnTR
Fczej7hwHFR9OXE6KTSUUYfLKXAHmjciBso46bwhvryI5hEFm6qPRB3Hfhduw5XCOE6sVbBbZZ1r
LAu9DnpYBYkk6IO1JmAkrgmzvIGA3DsEj+KP7pM32AKEkTuZyBdjyrdxGWAL64U1QXQUIulm3Ues
0OdNU6pNpU17sYVDsDsrSkwmhyaqWJdm+TY98A+Ja5N/ZauJ8MLaSyzAffRsAo9wW1XN5ItCfIFf
HxVvzXRCNPJzyR3pDmwIK5RQbs064Qh20icbqXVlb/iqHEWJpd6veX2h0MrXFq0mSWkBA7LISmM8
HjAx6uqM71meaNJ7f62O0QilzAaCxQcv10PfNGx7UD9WEBspom5/+8QUjUeui360hHggaqyokhbd
fQ4x+HLMoXLzc+uWyeZgBxEHEHFz4qgFnTI3INQy6l9lbC/Tr4pn+qmefaDx5MAdtygX2n6rKDM4
thhMAyvSMoJZ0rPO/W3aHBvjR/XHG3ApJSLonXBllfRYocRKvBygL2Mj1o62qLtA8SlmBUJnqhmw
vXNwx0flL2k5k1rtiiFw2Pe/wYCQ4Lv4aykmtLsVqD4PlJ4UO2FyEfXekxsyFvkuQGPeIapnHVpB
Y//m45FntfKX0o0FRiiWU6m09Uo/OgQnlIyuZsMH9IMPN/sVQxt+H7wzssQwa71eFTgY38XWlOVE
uj5X7kp9rUh/HrihLQKx9QV6IJB1FS+UTnsZxJPfwRVdNERzfRNpzFB87GsH3L+OaJEjrSZJvwmC
TVwFfdmGWwIhIXyS6QvmosqPdRTWDu05qRUIW6xKu0gYDMg300WQ2oYaZ3iVv2ps9gucxJbjfdp/
wWVsRX65T+LL8skG/TiRRZ9twjou++b6SW5nQJ9D9B6gLvGN58c2CP5krRJ6FReMdz2JLSVEEKZE
4p0tOKLb6eXHvA5Uisrhpv7zbMn568VLuoC7k+CoIUCN44sAvL8HOxL/9BMYhS0/fiTIkaimg9Nu
+mh5MHL0PfUV8HcsI43IZGz+ua8mYyaIt2lz3uF+b1Eqz5y2hAkZ0W9PTDkW8SzRrdvzHkZfqgNf
juvW/cKYWAR2qh3JoTYkwlEPMRUL3gM0QIIPEpsiSTi4af+zOEqFhnzzDEFZjz+VdFjxz8+OhbFG
cGyDmOFgCNWDA+uvQm53jj766cQC1ww/Xrg+rfKIXstSEjS61I6gNh7x1/IY7oD6F3LU8OJiZdIn
hYq6IEM/5UhbPcUNDg1f0dBIH6xBarXpkOO1u9zysxeSs2UTAUNruuAWy8lAP0kB/PGmnYWX0PEj
v85xGwD0Dn1LBqNTq8Ja3kNSiNFXsrRNwUuH7zatk2ZoplGvtNdFH4W3ySxUm40VntrB+mjJsIWR
bMdSaC5Dlu61acpGiy2oVWisjeDkZVOP1+XEnHLsHqK/xSTkTe8inesF27Ry/EoFC/TIZ9/uGN+W
guCuaBGLIYAHmPiif4tEKfwoVV27daDg6utDtH7N8IYbQR9QmNBnTrjSg3xlU4WGJ+aSuAQPH6RC
tyaFQ6GUq5Yp9/uV25kRVt9J2LUdSXshQPQUCnBuGl/UcRXYPyLyRFEkBx+nk+paFlMivzhXwReL
7Q2pB4mleDJEpsoKbY00WEWWAZ+jDX585aatkMF8ym71qMgArXWpHzefmQ+vSvv4I00aiaHOpKIS
jqfz3b/EVoA6M7zaNP3FFTqHVuSj9gu/6PBsD6hsSz5v08buP5chGfRfzZMJ5DoAsSTqI7AO+oiB
gM8gIOVTqX1Ytlg5pg3uX3DGa4FZqOQL5PG3ZOwSenvuc7J8kz2gGEI5rkHYwlhOG3itCYTr76hj
xG2G0zevDWLimW2D4UnYv7w3fvi4KFVnXJ0CVf2CuNbPRkCOehR+sNy9xR+ub7v2zAJzk4Sp2Qip
PSsyhP3fAO2/TXqGetE2tPx78Q+BS8NBOQHRK1LRB5Zz8IrOOmcrMnJJzIeiZilH2E3lrT4sO28G
okZ8H+woH8LBR6QfUuvkKJWoIXfyhfmNscYX4tz7ujak+jn1HXupX0cjiBS0X22HmEIMplLdG4GW
G+vbL8wB0oG5DKOUnKfi0LUhNvRi35GHQHzaz5GCSwEPFqecFE2BDxaa7+l2Mt4iBpTfhdnE3tf0
XxBMCFyeJsVxUbjBilkhvKjbT1D5P5t0jDPHP4htbe4faJm2y3bVaAlYGaKNc8kTt6L1vjuPB3Dd
WrBwcnu4UcqO0vCXDsT4+OgIZ0dC52uLB3qlDe93xMb1/WoyXRx/zrkNNInAmOJIAxDv+f4z0ira
jA2BRvwF+6JYqGl67DUX35MjEaLGzzeGRULq0MC+1SSlr84F7VxU0WtGBBSpfY0OskEosAxYCKC3
OtW7NqH9V3QehJ8RURRpAMavguZjQYuufk9gGHas1eeLIoYa34tk38y97qN3YiAhVeQUrLZSqIPx
9U1hjIaZJh5Yz/NGA/FYpA+tl53wNtT6jw1IqY4uKQNASozXcLJRKSZXH+51llGQR5Fg/TRXRnzH
nrdAaRZIGHnMmFcqIoEcpr5QEWJA5pMqA9/mqai1N1PqpdLpaD5XnY9umGBp93eV6QpND/NKc46h
djwA42Ds6X7Mckgxu1QQRGDsMCmbYBsFdptUmcysYd2JMxRtcKtXD7TUZP4dgGSfm4u2dgVWbchN
CdC8792Xudcoa0kermnnuNCnSYhjUgkXQeKNe598iYSc9VnxVjGKnnAVFNLwNTeVOcfw8phjoHzZ
+Nu3tIXHMrAvySUNI1iCYt+HWgUIJtuEnqqljV6L2JqAqATDUF28dFM5PoB8n4v9jfv/e0N05Tb+
u40w0gQMxlpi4rmodMFxm2IycXTMlS530GKpCtkrT8PEB7JNL8JFJ/iDnk1K2nA2HlCMTrH8ctNX
OZKPZAx95Cfe40+8wn7qJB1S1MIzhalqQxI1haRHslZK4AuCvQ2Xu/0/lD+o5vJS9PcOxTxEA3Iv
h25cDZJEH/m/3SttLHd9XOPC1UpeUkN/IQusqKiMy4WWzAkbdQNeT/eOjcB6+Secunr56zPMOxgl
+CzNNJ85DaSS51Lyvvr7cI+50ApUCrcUiDiyOZ6/41lzLoYNI8Ma8Prs3Fiti4RArWuKV4RSstG1
cQfS/Gr+OWd78wE8K/jbadT7e+6Ki9xwBOKynLD8P43TTv7MwJkIfet+KeKW0OZFyWI4sBG24cyq
fsUTNSHqKX94lZL0K8s8eM09woT8v00W8UoAYDAggV+QmzaG40jiO1lYsnYk2sAEaXLuSeBP5uoE
GNVMAU7XFQr1sGxypnmoWE/crNfQu75wsyR3PpIDvvG9vS50Zdfc8SWizOE/FRGOqIl2V0bRIO37
j/B12Ds0v5QCr3aiJlmnq/nWOB6bnkOCjAXIByyNGNVtv81rqvkhSMfI9m/dQi8aP1rVjlCUS1sp
dJ3vnNtAfjQ6BxcKloo9IFN6zqrNl66z/Mjm+AS8c9XwsI0szDIGkorBCbQyKy3/TfhWN31rNsJp
/wkka9YRKkOdeEyh8B8nd4RiAyKHOTmbXWMgnKou+xHFUHqbqfSGvPMvb83ONhFiEbDBkM40iRYb
JSUGX4OFuJ5z8a5Py2BmFjZmmisXBbviSswADjfll8iK3UNAEJ5hqnxivm3Dgud4KARQOWsJe6FE
u/n+i+yTduqKM4r8xj0Kk2qH44n2A78ij1pjBsMB9D/nr5sm7kyUjpKdg1WU8tFhy+xecsmXONGE
kgbEZDpM7AW8qZ3APUzI5iSkJl9wmZXUkafHV4QGIUVggw198ty7jeLzPGWoECbxQF4dB8TBe+B9
vPWiCDkj9ACC5BDCbazOwMjj/5FNz4ki7deWDgL7kwhT6oscgmSq3kskthcKz/0sRoA+61skE4t8
dtp39U+YuOK9A9RqYY23zusbIC9BWBZ3FDCvLfTdlvvm9kAjGaceeUQNV8DIJuTFchNHFoQ4rKbv
yNXPFxuYdc9IdVmwWhvUEVcJEJDWQOaMXB911hp3uRg9EqWcesBOJVwEp2UvkhITyTh4eb5C9c1g
LXLu7PzV/5NykOJmiwNmVki0hU2Fvu13uZZ3LOlkVwIudjWBV/yJUvahX3uYlq6bsg6HyHP9P3o6
pqYbc+ce+SCKhwEMC8M+XlB0OFdeAXu3QBXVrtT/pV2uVtLpStWbh5IUEZoejGD825Ao3BIBkhI/
oFnn/ZD2h5OVWFRog2T9x4bFt6r3TWhVbjBSpEFSRtyfIvnbWjuRNmm6qXA3TtSlEPSmUlaGux3U
1XeIdGv7EJD+AtoUxbUqd+u1Aqcr6ysG20IuiFVUXtWU0bLXPoROuy94UkmuE9fktqvb2szPI7Ej
oE6LemaMUCbnI6Szflq+3GxYNnN3+I2woSG6usbItxe6QCYbNdScUfRRvozqg8pJQd6VZwsP/QO8
k2ygK9Eqc6VD5cvCL4KmmhsdS1wVccLG21Piaj/GvSuQWhVNKSyY//8i4VP1rrLxo5hWCBfzFzrT
YTo95to19dmwaBJ4zf0hnvqstu/sKUcfAiQa46zjRVtf2sRUo5QRtdSOsJDbFIy2wbD5QYeVd/xq
TUyQSV6Zdu/T1/dBH10EKVN3ZHXwF4iytni+pC0VTlvE//b4PffufN1dDyVGIZo/DYp/pkuL2pm8
vr8hYQi6y6gws/OWjmZdcPgYGTKzWPCa88VYPUhFTDyCklQCxw+3au3Bvoxpi9Ullm5qoS8kc29u
KMQTmvAP9Mr32/QUxHqccxatvFgTIWOaZpNhskA1QulbHr+3yLPm0nL0eGlRraCJ+MgFd7juH3gc
HZO8JH955U+o5xtvaGqmBjQMMR5q77SiV/AsDNMFwePByYf0jFzrVxJgJm5xNElOxjmcIANYJMTb
uO8osVxWKBPJDdwGEu+h+ZECzruJ60mplj/c6VBEuOZl9u281WkzDX5OU8D6X+Z9wvkEOeIKE3LN
jgssRZ3BrJTYwn0izQdCpGgHI4iXp/eZRtyZ1+TNKNG/IhGVAiNx4V3jHw+yRACo6QH6o3ngo2UP
70dfeJLn7IhlPnqVlNz/dtrMEM+K5Qb990yPvSX1ZQmg+XIeSntInW8Dno5hgXTapyyV+cUWM7jl
A53dkSS4hODBizdi9NmafiQOW3Y2Vba2IjwGw7uUdb9oTKWyQTsQH35NJKrfNZah1uTRCJ8mL5Ox
G9m5ioeHWsiQx/6wXKI1TVFE55ZkAvUhQxR3gQb5Mh0vsdlUQ+QNsgJV4Np3/gOkvbVUxQlqaUUT
cCmp19e5PVDJ/UDn05R3i3vfa8CK+Raip2CJxBoV5jB34aH+07AF96r0Po7b1PCBiNfTC4ncqTqg
oDp52QfdWCc0fud/BWv93IXZTovjVEcZLdxWzxa/AYtqcOi9tDq4n284rU6fLvXLHKWTrPg1icmN
AzG4yJA67mM8/NPyfA91UULZ3xnTi+uMOWDFRPiT615i0ZkKj+eWBhKFTVAULlhD3be+wThukSnN
/UWqXy+EO8ogeczxL7TVMfLFYpZ9Jqo7ULvKT4wOIlE5sjvhql8FIIDr/I6jZElLpR3DDiufdOlI
odRJ71x7Tcj/QyQFRXrLwgfPFGy7j+WGaOq2ky+Z5J9tB4Y0YiEm6mosxrSjEPr3RsdLLoaKKMWW
CMYwpIlF0g0owyJwaYNH0tfB244LZ9D9rTA8rnkQ/ySafOM77DkrT0lCtbS6E7J3+sfrKjxZgw6x
2f1JC6rYkSC1vX9o6aLY1ZrKnBduJcYCvAz+qwl/ZT3P8+7EHmIxeZP7usYPYM/14bjUWatQjeVM
C4/Cqs4E89vHRw/UHzvTTYGnjU6m9jbxwfrBS1uD+zx+Q2a+ShfLyDTwILwAplrP/IqOompEn4/P
4ityMtExEBPqeFE1hMEIDOP3GpQd7TttJnwkucqblmYhSgqAvYtQDESh7oXc0/nFyvjlopddRRCy
1zQO+vJx4+atsgQHoURcH7BDMjU4X+zt6HCbrQEeE9R30DT+tBKZKQs2YR0Sx1f5fPc6s939j0iS
orKYSjQ6BsUCmatvvfm0jtlHd60CJxr8C0a5EznAH02CTwnrQP2L2eukwy2iXmCnObo3iInuA3UT
QdFf8cY5l355j91KHyvmu3pPD44LQop+pT2HXUjYWwxaP8jxECJSxl1tgTxtFpl+92B+588y5ysn
n1pZ6GdwoDXot7YD+s2CbEM89U9QUVFJvkOpoPZx5uj910ATwf4FnepPR91GZ2Fk0QbNPsCtn5Z8
6UlACKt8549V5GaGAlTPPwx8i7ER6yLbvKd6mMPalvCRtAzaw6ZdFblxoJFWhkqlkN28HUPGXBEp
K+MuNkzjh5iduF3bBz52rSqXUQIhOqmoePt3fQ3OWtvDAJ/V4yzLqFxuBdVz7bSkYF+DMDi2C+lH
Z/L8KQD/yW+RS83IgdyLq1TnR5K7pRSbnHNgfv+3YAuTPAgf8GcYtgmd461LkJOIxItPCbcJMDhM
KEOLXrheF8plXt0EqdofDswo5UYPDCVgzOHTq2/7ZUc3sHv+gP0SfoZMg7BTdKgKjz029cBHIwFe
oalJIwXwYZ364d1GKVHrK5dR+xlH4GERX8DK4bNs+xs8ZqG5PAbEfoD4eIy+6F6HPW7M0bOcKogQ
oxzq+Fq5mTFtTL5y9+jT4a3CR6oupiedhjEOithrmhX8YX7whKByALW9IJmqP0jMVGr/pn2ID7p1
wqYvvFrbmdKoYHzsqznxZnIotNLvv94f2sAYeFzJpJOcZO5jpOAtnBpC3Zu0mLz86CZVNA1E/mvm
Llkqb0d7MzgAqtmxCMWUb3RLQxY6u8Zadq17GNfx1q5BPVZ4RI//kX17U46WONuEGIa3AzJVC3oX
t8Gz7cuUadSbPmKPpRe6GvkwZdqUpmGaWJhOVQ+0SM77sUayj4sxM0waLz9nnWOb8iIKeWsKf4MW
2Pl41OWtGvvFLwJvN6getrJ0vripKLItmEUuwtxgTwkYtF5VcsLvLBLYUGP+6YSaPzIvcfqAdObn
LJ1+6bCadrnBlwxlubux9uGxpVxPPGFoBzAv3FResjXC6LX84dC1juDs0okGYUBj93qvKP1Bhjwz
FzY+pIXvlGH/9/AkqmA86xiFWRIxTRjFIwP2eDbpAsdu2K0Rq6ObLcLZY22y0XxPExeCPXcp166X
uM1GUnVmABgSVcGeI3iijloEYodnowDJGBC6VxX1OCHOfeZvSnlmTL5mOmfpBD97pQCpQDJgW9kd
VkBvaewqsH5JjNxLmyLP10zWwmYhWttQewYKF3SwZLe7TjsLj4YLpbkYEaMUodeedmgmU9LqQllA
NuAR6Q7ByAmcs6ooTeL4tVxBnzS28ppDq3D1HNoxCkUo4Xvu0LhfJttEyOeV6JcPnS3WpqiRW0aS
wGLaYEXY5Vf57yM9Xicu2sT+Q38rT9PzUuJS6gcj+OQaZHw+mfFMfyUnr5kOnKS4dVvZE738WsVt
JzMFhHtFVBqyfqokx7SGMg0q+UY4DtR4GiH3JugxBqeAz6W3BXDLxiaFMKw2QgB3n+RbJoQPWzSY
+vI8C0hKSoFjz30mh3o3uHtDCSe3U+sB43u5d08/UjU6jiIkKg9dyU8DRbiJWwzbGlLaSTHU+gtO
NuNErJWP16nLfIzZjX/Df61w3S+Ca9nZ837BwUY8noMWGIXaqGMOMFr9Q+TS8UMUEQLiV7FmN4ji
BKEqwD43nwBIga75k+fzgFXUtH/nakhP65auWBeGzSnJU+T48jXaEtKBpVNcANqOYOTkc9+M0dsl
iGUMyo1TehDA1uRDrxG6oeSfJnECvJ3ZlrCaw+7DA0ZPo2hqbj7H1erRRBdy0PA6iBuxUYpkJg/g
+Xsmgo1LZNiicdZn9VH/SXZhKz8yKIjoI/UqoXSvZaq1DGxXtSuYZdgcK8V1Mjs8OGM+0uMb/aJI
TN+cjW224tX0Mir/648vKPm7cDwj+puz4hUfKHRwL5UM7tfFXaBKrQVjhQGPymeaG6X+a2bu5pLu
AwvXB6P02ZXv0DW6EtNblVGU9wAy/QzFhJOlUfEczjK9ws0ux1PluP8UNzrMlLBfgxake09sI9rL
15XItSAKrnLrvZsBiokkiOii28+OS5TO2qcIiN8Z+xQsjLPgb8rQV4Hv59bTZGs82rMF3DXFw50f
NXZT8vimKWQgJ3dv7q3JKcHCRJfVuNhCeIuKj9QH0/HWKIxI879oOhM9zza9WxslT8E+Ox+9RLY7
KxjHFfi4Zzan6dINThj9q8NFAwF6FPc6LVF90TkM9lfPCirVdv6mSHvflHNJlHMdsW73Bz0/RmAm
oOpjHBfJjDOQmql7Ay1O8tX5Pn9mqNUZFHBejcWAh6py16PBXM05rdSeWyqTJsj7+qGxKCxsYnE0
t2vanoN4Gd++4Ytt8WI62+OedkjrBZSPE2g6eFIDwVo3CMfo8wmQAbUUtJ0LERo6hT28jv5iMzr7
C+NyzGhDos815vD14md0QChcqX7lbK/xxWPsgARXSmclVCQm9zIjZRG0oGXq53CuJZTbHCMJT3TH
R9oa6IvC9j1ZrNzX7RPADLEIe92l5fEAckvIB3cVR59rS7AbZ/2QLyxOHUlQSj/zoVJ2iG79NtLL
tswL3IDS7tKvxiEL5DSB0rsOgFmYHRN6QSMkDxbiKVBLOSjIezWVpz7o/EA5fqtkD6VOdo9g8lLE
2dDaRsjtk84gSbNntHI592/P1wvlcrJsHd32sPn8OsEdrhrOvRVLg4AvIoE07h77i+JIkLsSF/X1
GJoTSnr+0zY9WGkQCBqAvU8SoPyGlDQGWwZwqqsRUwU7lKLpBt33PSqa7Ct2A9p1i3u3M2ioVfcm
+aiTMl7t8RLy9rXhexUwjyfcgiGC/kR7GPDyI5D8xgMv9VT4PDYdLdXYFtpci0uPrGqGW4FbjtXK
jjdPwqjsu15yCDospuFMtIMYlw1Wlg9vOg8CBxNYK7Rc0AbvSAOABB0XZL86SdvusVjMsTYYQG/S
q/MG18XxuSsn53JHnQrNP8RzCnk+N8Njp5disoqKl9OHZ2+HscpLzba4TicwpKBLc+lIWyeLHQME
jKqsOdLEsCRkJSUvREXBSqQ3kU0pe02jAkNAAmeLXK3tNlIMqAP0y94AS9NmI4hqIooJkfvIyP17
G3x5bZVQTe8VX6pQ128PtJ4/I/L+QtcjyC/oaO6GA7Ia8dbDz3DPsCvn6Omg3W8spNnM5r0mjKLP
5QOgAVksUxWMd6jmiCMx3kJPHLF2ussIRxWbVXyDq+DvkYMe2SRJfMOrUGNdfpJb91tQoLaLpBXB
048mp/Db983bhpUi9mcP4LxXaNIq7uPlTLHdBdW+2oxFME5AbWSbZx4A6vckQHltNUxB0UOSotBk
+h/cKE+/r5uYPXfa0HSXjX0psVtpv5eFye65Sy4M0qkdI23OchhfbAdnDf8J3zYrtPqbzYFEnUy4
5/50ipjPrKp17OU243seqrGhLI9v0HxVmZtXswnZfIfgR6YlHaNBVv7WcKtFwqgNq8J65zWxhu6v
Ed6cySIiLUh798qGRw182q2WWI2ut4y6mURlfnH8Y+HC1/+hBibjsy3K2guXLuvi+uTSS1lyDp4J
3wn+fQSJsk1N7d9hOJc70VD2/4BBDLgnLW1mjxmFq/ZLNw5r9jUOEJKLJFsQp2FgwIi032Peb8Ht
Lu06Wz4=
`protect end_protected
