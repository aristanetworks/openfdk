--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
EloE2MldI+Mgta3ZWnol/tkNRxpWmPlImQlsWPfVVtZT4VxpESgH+HvIXewBMaQhO6LzJsq2f+Lp
fvLi6VWs73YfbnNg1/RG9t+gMf6t52ODQprOGZ6nQg4wT23ptXQsOWrwN/LaLA5YHxpplLsecF5C
cScRqoFZtRP014QMdU0qIjnRqTIw+WjJbHvgKvgk/mIOpM4pewAAkfkm0kXWQQSxsWkquN6j6Mae
ZVUWQ0N5kBF7rFruqDFKTOY/6ZLKIdgyF2jYb3T3AdbRE56kGDX0g1Hs1FcwEH+aSKxzYIfK4x3J
LJ70s6u5QgQXnJJiHb31c/3IHCJpPqqGffzJCQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="UdZHQ9FDvrgwQAbQvwMr4zd5iLh+KLaq1WSvl9abqb4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
L2F+P2kXpf75Q9bkgdLJfmuZjuMmZNY4/uP2dysy9Yj3oss22/m6HD3X6ZvqLAOUpsulr/8/bzLh
Ef8LNeIIWKGm7xzhWfMu6DQ+cs6TiSSXOxaGVf2zs5vBC1Mc7U68WkLekGXiG60ghCrpI4t3W7I+
ar/KODDGYAqkCvZWScBTSA9JtQW0ofFfKlHLU/VCIP+5AMHNaUKwiC7gPSnDuyGWz3fK7mWiebLc
wf+hYzdAgqxORGRqG/kC3kZPYA/Bd1Ow2tTqSGIvycyruHJllwh9kEuKRoOqHd0Tm90cp1oeTFtt
IN83ATTVjj8nX4YwwhQeVPqrAcWp1jBWHDM+5Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="iv6OLauANtBb+Yai8GtlAE2rNUZ72YXU6YDLdeuUjDs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19424)
`protect data_block
eCDmS6Bq0Sfk4VmVNOhYs55B1rlgD5vpm5Axr93BWN+vQDin5+Y/XCf56MPGOKFWzuHquI3TKLfV
xDfL0wvg80jGOuDTq1O5G42oXAb7Zb+Q+ahN+tW2odqnDQXW64dxenVTk+0W7WOXA0sK/BgQ1vMm
JanpxQ+qfK5lAwFLnGajx6xEck6Af84UcGOrZ7SOLjnaPt2R4FDeDtITquI721jitYbFxS9WLGPB
fxFvRe/JsatJXpSHQL55oCQePYs2IyEaxdtMspNSZRu2wZc/R/nvtkmAViZnTUFL3nIDJHsqjLPz
7lh8LymK16dBGcufbaeSusw7mVF5hLBuArhmD2ZdSna7Vb4uOMseY3mg4/GTPG2m5R55HlLFxfqt
jdRteJbuXXJ1r/YUnA8jkhWtQUDkTEzAYMl3xpgz17BxPxSH5fKVwT73vZWSaMnsSSfJ1AQdPjwp
TgigAVemKWQVA+QhDw8ZM+IDlU/ToufvPXquMFg0Zf7dqyDTw20S6e12d0Fu8ANcoqX0asESo07Z
fPt4Dlu9mWHtS29vwHaTBHlqb22AL9lGg4QECaZuTWiXvrCitydngSw8p82c2WvgBwN8EBRIgafc
HxOM+GRoRSW3pCdd25Pa+SA9IOLKG9lNlYHE/fybsTZUD6/WGbFVTBpXmCBnyYCOP6jNPB3KxUht
FfQBG1wE4RcuPlJzBbYnc/xwJLqc6m6MoJzyEz4yr/NLq24dWe9EMMSijZwtnxpq/gGw3exHQVoN
xFeRxKIxNoi+wysYgtBfWLkWhbr3qfQByq9hMCnNd4wkpgcZKk9PAn1feLg74AVXi+uovIbxcdSn
YLa4BBKZUV3bA+7xOtFKQvZNoos9/65UnM424p4zoihEtUaDPcKjc3g+ru22wYPzRej3anNseBR6
k8XxppDgt/+JOgsTxBFsuCXoTMqZASvEehEe2+bgy7IUfp16GLea1yUWusR7yaoDJZbmbUNeWyz6
NwdJWU2S+u+IdseyQ0MFr5bEjYuZL8uYxgHdAOlbPZI+eGN0MKM5dAi5CZtWaX9eK75dFp6U73RP
UONhxCdRAB8A7xOk5OPcThJh+wFUOoVuHHj+rB5K2pbn70K6sEZDxCBqlHEMljnY4KTGGox7KjWS
FvJ+2NdHAStT6rOMxA88uOPyIaPdY9EfBIsUqoosQUbR+UptI/k2EnEE0rwer4pH/cxcIMJ9p/kH
9IhWjEVTycwG7xORaSJ+dYTcJAtuuvXOMlOcrqvCIk6eAZKbtk6DoqLg59KDwYfBaKExGfWcY53Z
didtrUJdfxEX+c3yIqhCxHiq+PMktgI9b4A0uzCtm4dpKghd6VK64Oi4b+d1Sp12i75K9gv8Gp+j
xXGmTDnymGAqeuAVD0ukLZXXwIK7PE4mY/1Hy+5tVQ4p6EIO1KCKFa/Ta+jxNg2ecrjvI9gzzuhN
zmpYdtSmkMiohR4OHmbTxu20eSv8bSKigLMBMbmjB62tf7jVXtAVDrHmbxHFt75O5czzXrwHro6t
RfNHicB8Ih5eyD1exv+r1vuhpdhshKQ57ul3ZZFsuuR5TCkQUBDb40Kfb9SVOeJSjo/GdRQBB5Bh
p10EHRUFB7HgWClXvFfte4QxsbqETQSR3PcgmIBM8zOdMygZlsTev9l75dhq5QqNIXBrQ305y1w4
9hEajBtvNsE3aGyBGgjLri943iPUnpW99CF/7CUYCTzkWch4AIrZk9BQDREwfoEJ81adqRp/cFHY
DcF/lIezdGYxOmancakjnoPKAbmf5uacBwLxSK04OkTywyDa2cV2iImBKUVJ+eLeerd+x3HHLxGq
MrzwEgthAXwztgEagA3Cw8WC6mkKRXNFp1eUXLU+xxi97SJ3tDSdbRZnoKfgi7r+KCXnc7E2UvJZ
AeBeo/zEf+eRn3A2CWkakRJ5vmv//4awqOJDIg7Qvk/quVNIQdzsoQbIHw/2zTJDQ7oxHI+nmCiI
Z6ly7rQOACh7QqWwP8peW4228HMhuZuj1hdDUfdpWOG8pFKHMityJ2Yxn09+KdcXo5YS4Hry2H5X
68qZ76rr6mEp7oQmYzjVqmoooL/l5CsXIOPSRNDSjHZyPBHGqgowdqAARnDDQdZr0DgUxcIK332N
XGrjEtAmYrEHSinOlm/VnysEjIzGysWk0lO+nw5QQhz7kDZ8pFwYCQF0dSoPQfTEbkaHkRumRAkn
wQmf2wP2SMkB4KQ9timskFZNuQPvaYx1vCuZfTDnxjZP78d2YwbHA8ObuNlJ/YULf06t+8eaFBzf
ISGzXWIUwitiZMGizZw87pm0VoG/0ZVBp43Pf6/jj15OWGimEcfzwV/9eq26wcDStY3vn+0KdFR3
rkKNsIh/HJniHWEu/DIW40lXmk80GLxd5do1vpiLj0g7i/ep6sK5df9paBhj9Cs3kIecUQ1dKmMS
Aw/QTx6QdoxBgnKCHYA3+wzmfCml0YxDy3ecH+Ws2YZP1hB5CreNBb5TE+0OSqpPxe4E4NAKTOhd
7Vy3mJxuiVuSh7jmcmZpfjLTjeEOHTMk5N7GZ383Je+jsFfg3YsU/jLk6Qw3lpYjtxLY54vs3Zdt
Mm+/w+MR7d9q/wu2HiCj+B46iRdtzOmI5YhApymUEAypepVP7eb4fB4GKluSOd+4EE6dew7ytP1W
P9j/o+NKYkZZNubUxGnCPpFE1wHECOex2ykF82tx1UHv3HpXdt4HlviAvbwzLd9ziiLc4srj6g95
piGbCrXY5LiUopZIV6g1PIrt/EWlfmNxXY+kO8LwTkKBLQLeAFMkv67jr76vg2SlMQ/9W+OXVzPS
yBQgg76kp5gPFUgh8MQ2efF+6X4j1pUiR9z6FSdU3ua8N1fTaYiyWGYugIp9cM1Jbz8/v0rM2EWG
smnaL9T0PACpgxOXnsUcupi9tVn2UnVXbyo24ckyBya49JdZjIxD/4kKCvdJHuiPbZoBeYnPnvpF
JXFCiBhebW2tw1t7CISmklcnu6Q9e+c80j+21svZZlJOuneHuEUwzK3E9kWxcUaFAP6XpNWcZOOH
CdVsb3bUOtdBC6kECsKeV2UTDPmc7W8w0gcR/ysCEGAswwKWuGSNFb5vf6ip8YBTZ/cafOqZ1N58
WAsF0d8n+tiYD+xojjuQTX/67v9tjjQq8fL9wDmjP+AFedBLMMWabenUO+HmRVDR91JeMcwxWiyg
4EJfblwC24TQIUYkPPTZLBnSyTHE7Ob1HEF+Z4lptljqvrfMWB2vvsC1hjnhPjEH8aW/NqOsKSxR
YlHBIThdfEJxezGHJCfiKhAKMLNziD6dq2c1ksPOead1jk3Q7+JPYvOPnzt34HRnES/UtQrdOgHJ
RIftsKcb5TwS8UAaah/w8YyFV3cUg4OiKmQvve1TiBrpXKIH/GCNrYTbRBxmkvLkRFGX+oLbcSvS
1EnCGzeyXiYDSOxxUlPx/XScYbQ2q9NFneEzdUvVaeXWInBlBiKI6d9tV75FVtBnSQny+LBpmNmH
LZgf1JB6Wh8TJ7qoZpdF8nfOs8XvdWFdq7bHSbg4BRZnIqJiONzYx8SIcQmzlIPbDpm/yS6MbLbh
IT3N8WOWhg0qOloky61lcHXT3V02GdwWCgWAvIkmMoxl4387NqWrZdL5TO2aCyk0LPPj6Bsuu3ZA
9fSEAq7S+LOzomjbSE4as2qfvgGkF5K9bezODFDjVp7akjsr9CksAkdhQUufn6P1Ws1w9bBW2I1/
NTpYoUpxVUQdCzhgFbpfPM2xhA4LQ3G4cQFAxglrEpdhVdC3BLtGGWBUHdOKhvped4oSzT7NOzAr
2X3kgNbpda7z9sEyNGld3rPmN5lYBv6x/CtbZy5OKrLfZbBPHgmzimQRTXL4M5jDSbMKUxHyFKwN
2GQi8OPrwvF9tQwxKNHDcjhW6cP+iW0nyf88tURZp29mA9Em4aSjxYjgLX9I7qGeGHiPTCGrZd9v
TQVDjxhHVYaLaVPGJHUxtv0GtSXBJUhdMWhlbB8by8SeNJJSklmCPFSk0LuVIL2kliuM6TLc7T7E
f7MuwJWVHhMyB8wYsy3HJLzAr6oRJlUbVVP6xW6K77JlQiuso2XM2D8eosbyfJc1nCECWnUaO6UU
AZ7CFBe7vN3g5jHCRt7Yg+HlfJdHWZRfPjs6Vm3hjYekAba2I99bADw+BcAxeTDUcdD7U8jylY2H
zroZWb2SLYlelbvjbCzaQ0NJE/0t3Oy4RHQ2XfUw+UODO64h6HDPjz4COGSiImeT7vvZNLGcjGez
cWqFPj2XjJ0gOio2VhuRH35cjM4TDQtnTv6r9kyyz7vF7m6qdnciBv/8Dig3vvw3+mr8K3n50uBf
XFWbmBMBV11bKLUd5RkPb2WVJ4snvXoKn6i9jt6f9hUZgrkNGwlaGktrYgmqFP7FH639oJPROeq6
GF+E1oXo498GBiaSx0ySerD3Vt8lDBpka/Lko4DFx154uq8HeppRCqgUJmUcZygnb8iweDsCZZkB
9me3IIpyJfqMY3u09zC7m6niW463JfzNs0TODze77NUTJjniE5Efhh/rtEJBZkVltprxuuTy+Zn8
CqNGXfF5/oi0BhLk4JP/a11ZzJoxmR2UmDr1sIl1SSTFhBSt+0CcbPj0STAp8nFzjJrFHJ+lF+4K
bdCBCZV29LYzfRFGGoY9i0V+TzKtVKt9UpKoNDbUo5E4U4L31dL3zWhnKK+SedHVnGyJL1Qh/Au4
v8WIz5YY5RA9GVs3EuxlUjctNnaJ9nBbjuSpFlUZhdsuHq0YObwqSMT3VTUk4kwM4301kteVsrcQ
LYOQaq62KzOhE2TZ3lGe00HJk8mSUgaRmkKGt2IPabCOz9iumBOYKqtPqqZEGHIaWHpebyzfE5tf
d1hTc3QrB3lTVcfAQRP+7oQwl303/My8SbCvxqac7goQIa4rhHLCO/24TrEV+UBag8fHeVbRQfND
hRX2poaQkq38C+XPLc1kPE3lIZdxzRyA1/BugqTIBvBaoyi4y+KPDKEuyDW3ksqun/dLQrYvg1Hb
9Avx1f7hraQFPLnBqI8NvpttEkYCIIq6d/ZxfqRESUbL8s1dya0mrDm++XvL62HwJ7xFdmP8u2uv
slO88J1W6v20mTZoIdSbwLyBywibvBTX+owg1BfiSi8eHAJcSo09covxzSLKxsz/SpHq8vLVu16n
aQYt8W5V0deqdyFacrbtPeDCvAFLH2+Q05m7xQGjksi/yweTZK3M9s9x9M/AV/MBx4HVW65o8AIH
Yx79Xlat8y33uJxkZKa9kjWOFTFI8bWm+4kAKrJo0ZcpbfO5ULPVi2Y2SuWBnmyP2/NqD/0Ubtkz
i+2glQ45s8VxkKp7b0RAauLp9soJOUMDgpdSawP7bjmgUBjHzWFL+xYiXs/6GcGgHUSa5zT6H+X+
EIrE49z/tUB/bjv07TM2KNDCE8xfuSWhafbDBqF8nkPil9E/11Zoqazs0zu1NNwfBGfIpRrbpfGH
vHqkR0K5iPiTegnozcoaIFxkUwzOtuJjdD4yavWaUGNCuobItlgMgciig/jMCw97DICgFk3Ai1DT
+BUVtgRbY2dHSnwbRJvJwjYW2kDTkAAwqUsjxpPuf49CMTtwHliqzDFeNtZY98b0BKU0ILwhaU3n
eNRXC+0e/UfiWKNjwCPghdjcq77Wwh4JzGiOfjNJP7Xt7TNki3olYnB++/CWNbdDTtzXjrFcx/ae
raLKjgmki1dRYoU3XkoKHNzm0Bf0SuecOfcWLO0R3kWrRDJteXRVyPGCeFLCpRJeRnRmN57XoVKt
x8dInJRToON5O+X0O2P8JloZ81SNirb0vMRWEYbE4/eXfzypyKPverEgJ8gjZDC0lyhVywFLH3L9
gBGyEPFNYjYLdcyf/FE4oruAzn+BXXnuRj5lFL2GZs0ckklxDo64fFjqqEMSm3WbLoedSKbhuesX
uu8PKkIVEU70PMbe4xpZahX3m1QtCdbY/fxHCtuwbwR4gq1UF1ZmgdH7MKPHMMNrGSJ5PTVvSN8l
iDGoZiH8KuezKarlHzvOJBcc7m5xjrOu3J2NtWNvEyMzUadlzmOy0lUyX9NkDfNwMsz/NhLExZOd
Xg+pN0U0L/BlyDukZeNaZa7As3HneZ6ktRWSCA6qie/rIux262Oyq1///iUd6PLXJhh/h+3baeA9
jwrUjU+xdX/SefjJWdLDPnhr90I1lLdUDrzuqYoXF5zHzRDopb3dUxZwKB1Al6rh3p9QTKxp6Vzf
ez/NNTeuTytMOMAiFp0xSMDClbFBFqZfMmAO4T3eIMgKoMFLeu9UW5NHID9LOPMFvN/0QWiRVijx
kuhnPgepZPLX6L5tbSmdevEyFC1Hl0UbfAecNFiqxjjDvpILXKk6OMhFsUb0vtbfvCqrzC+lQCyD
Wiy2B2MUuElz/XmoyjCVS3RSvlfy0vkow9RqAuBk2v8JIFJoYdlBiofO1ZZpwvxYIiN7dUnPsH0/
TOIYMTe9El14ZNyOKUc2Bh/KzcL+OVqY3M7fagSYCJ5Ag6Y3Whvvdha/tLPN4WjNb1sXepn5+D58
8KDkFtkSERsYG0umPpECtDSaM87v8xtrC1u5yuq6TQ1J1TPXBTGfuCmT2PuOG5vc0bilRPjJTra5
uPYWuf5Ck6wymgs2Y347rQ/7S810X7jyAcIY7ekP/W+cJOgl/aka5hePs9F5pl5+mEM3sbDTu4+0
2jcrbz912NdcRAnVlihM1xi9JDytjmz5EyiilkM1PuS5CEgzlZQjsWRp8oDu7sLZkre7tTwcqA3f
A2AGvfznrTwL83cLdfT6ZfEHxVYges7KG0qqRaeVBd69fZ9D6PtLzIFR5aK7H8lKMUPkztoH90L6
/73/cvi+lIL4HX73sWoldSfljVGv0j4ntKsdcYCOobPyf6xg6+rba0YiRfcgb51iH6S0PYQJEK7g
vF5srVGGABIYaOhQ5mC7bnozh/aNHF9vrFspDFsXl3POTnM6w4XkSrd7tFC1BGUQDEQ6zsz7OYZ/
E9OOC/fkDDPtg3VyMuEKpC7a1RxhGor7o39EHhZ1n1FLoigf7j8XG6Sj3pMTuPP3kMqeV7u9vnmI
bm8xz4ADe2WYpfsnW5YDtOctTFuCWrNGZUw0SlkPqDE72naE3il69O54g/C643He8iI64bJrgbq4
dN3VCeMCPujum6kJR4nflC48ubvglfY0EuTq3RvbgzSNkZDDhKvcc3laQEkYNeCdE7XhsiKGwVtQ
cjYlZAYCGPtggJSYYdqf/dmmNO8Bk/GWtfknmXJWJ1VwZWgRGF2pd/k8CVHe7B+PRvPli0MyuFsZ
xY/Z+kmANFJ7MBYTflaJjJzJbzc5B4HE7QVb+IAFRJUjodbqJ0lWcJV39Ss4UfMr64nnRzUyflM1
VOAaqZnzZyUkDNjc0F+69Efp/8Akhr2kchh2oTLCf4ZiRmHqZErapfGINbCCZVpIfRfukMgzmdLZ
plXB/+eKQyac2j4atQ8Tl3Xm10ZsNAxCXgmo4baUBTemofWbfcZBE+e5UQl3Mi3VM9GlmxW+j4KJ
x7eRX3DLnC1/ff31qsDGDbIApar/tHAfwBL216x3FofQ4FzhOXDnkyxxPx3oZIZJY1Yfyj2yfB36
WahNDWPHs+9DFEb/ca0zervAgrwaNC2nJii1Fot1tuizWuO+hI2lSmWPMbKdtj8bmOiSp0xd3J3F
YNYdk/PDwkd7DEr3Xi/gQ5QxIB3uP2B8a6RS/gbmuDEqHu7fC8zd4arXg1f41m8zJbQcRl+eQbb1
QiDI3yZgwGpgC/77fxBdG3o+9hj57l/bb+3LmhmDY3x9/ChslrMIJbOBz2o20VM9+PUu1DL4eS+o
nuGMV+HT0lVTpIkoByuKrTuhBWzkFBeJidPuYqBZY9VNmqpYk1nBdzOU4NC4SVzGPZ+NQPSP05z2
ARKJ500hpUOegAynfkJSQ6eaJOQzBD5L2ZsPTBb7P6LHHtbd5ilRF5ksq3mmpV3Hi8PbYkyG+iNB
+5gGLdC8H6gD2CJrPKkgZX7zA5CoTtV/x08Wdqol1vzEhjk+rnSFOPARCD0hCx8c+ZgvSGPmZXzx
g2jmWmg8gCTi7pAz4F9KEk6mju8G82+uX/a9yeGRn7G+Z7tP/CrMalQeLcCWtMTM3Tuj5fFhBmTi
KCmprzMgKanRr4bMrB3nR8iWYAX82N6vh+anIV2aAwQUzF50dKOG2pfQWTeHHdKzfzqsNE8pBI6K
A+DQ9JA9Whfqzb0U2sgVvrftLKQBIKCpubII+yzJrCAv2bjbBsGBOMjkDP3o/nWu1X1FMg+Qo9X5
BS/48nTmw619O6L23CesyJxgd+bvXMN2FaBOzxOvX6TDsHJcbsazYIP0vVtCuxw/4t2EBGXgmB1s
aWJKRVNq56HmCQn/X0lTom0iB8trH5UbpwaOPa26SQdZXrCNqDEr3DaY6+phCrMOyH91UVeX2b0T
SsW0a0JLvCPBoWwZCdZiAeaVpr2Z+6K2JwlH0YmsuO5lLsfFB/1/6Qx04Vofkl95scltIh4cvpCC
UjgxpKhDe+D9jOSgsH5xENIcdi8Img49h9sy/K3WbSmROL2vJ5VIxOcZQq9kCGR8dKwUi40YPRMM
zkAbzE0c99pTW4sC1sbtj/T5ZEoFNDkImyYhOciTz+ZPcww8Gf5u1Y63tiU8ihmTf/8h5YAu9kg7
8gYEWG6Iliob0h5KcX1L4WOx97K8KEVCe72M7EU5oVVdvf5BlcsdI29yAk1NTarIqBYPgGhZsYAQ
LJsWTmKDieZ/3xodMARlni0iXsCy9E9jHSedhIC728JkcVkArqWSwfLwurvSrMy2B19Q8W/lHgMG
kr9TldFZJGlE/yTtFXKQPZdwxLCmReIqxlgmw9HalwkpD7SnECuB5E5cF/wjcope5LM6vv5djhz/
G5GJA80RNU+z3ihFqcdEdV6eCFHaYQLPky5GSB6Goy2vX1L4N3YdUmZ04gfDhaC5Se1zPZCZKuNO
WSbcTkIaI6VjyXiiCArtEvvjrU31rxxcyczOdBTE7Bo7zFGusoF91eS7vlfxWKMZIIdLqM/SjZR8
4F5UfzECZs3II86UkPL0Hc5DxUEbObKKYL0VIeWT2lb4jdKcAjEvB4Rwhrhh/ufF6qA0zHOrfNJ9
cS9S31ZXtlHrDI5+vnasa7LDincS8sEkkm3DbCFJdoJUJEm4OwJf8Z7dgM1Rniq1YU3wgwzDDu+B
+GUz4pIlwdI7/8HvreVJj4Zb1y0WcLHV2gX3LPGxB9quQO9KEYGH/4L7AnFI876wFpK3NrlH6JEC
JvI/pjl1F7NxDsjTq5JZ4qunwQ0VjKhG5onILtH9YTXZyZ5/gmNutreC760f7+/ejNqIi3fTx36a
nvibenzwSrrzaABF0pK8GjbVcED14Eg2OFpdkaK7fihRSvrKY+HU/UwQVYIThqwwpSeRIoaHg0hQ
Wo16lzcRH7SZqD71t7S19r2o9nz2PUusqjOI2jLAzXn15ON+fqSLdXGDB5kHfXVm0FZBxiCdEKQy
uGG8kb4T5oW5iwSI7iBbf3xxtq5Gm7uJri+zbwNWpyWhZlVfoNGaHBOeSepnm/RJB2WwXazMmNeq
Qh2LF+Ki455GJx+Yt4mAR+6cyikCd/evSeShdmR4G3onz2uJzCxhmte7VhnB+JKvR7gPNUmN92Um
eNic0eZ4vfPuN8985Xo9RdRHfh2rF2sANea+16G3Hc0j53cxknaDHjFwMxqODVlYpBmAvmZt1Whu
uPlS4cJehPoAgl9m7Ry+rb6Fz6ftMAdPMoAHP/uagKPttyNd3dv8nNUPHYpqKSc6cn5IxqFtSzOh
c0H5/wGgJQwdq07+OZIOqDyDnsfhWcRfuyXtVf+jSET5kj/1cM08MiYwFoqkBDPrYhtOOj1KatNY
vB51ah9qo4w8ixKDoeg7AO8/erwj4AiFFna79iBIZYXjOSXXX3spyGGIQGckjn99UgrP8n5SvTjD
5yDz+BjYqZUq/HJ74AZDnLu1zSNFGIqm39J2AjOdOQmW+UYqZXHDkg6g4bA04Be3FPaUGTRyIqU4
FPmi3yoo9PNPFo6LQTZEC0S+sB0bomY2XipZoqG4Ezz+swvcGdAga3uleaSeOklWKOAsfm0b3+SU
VrM0PtvFnOOgCngXtrVp8iyQuXsrAAAWtqR4owgfXtGaKl0rPCWtjiTEx9u6GbEmhfsPUwfJ2V5A
x4lrUvJmS1cwQdVGplQJ2GW8/VwNwV9wgHRgdN0Zwc3BV9J1s43ib/AoerZUVaG7rqTCXdXtJ1f5
IaAXlK07fJOeYkh/cI4MYjKkJbbt9P0/3W9x62Vphw5oKBLs02PhlL94mb3UPfELPZsFdY5NWVHb
5kjc/7CCNWz/kQYiUGoYu4HqZSpE1UsKaMbPhsR6ptWsdh+PeVZvWHXX6rg5gPHjRJaa7R+Ba8se
d0OcfQmYmPipeFAhEpmoMK8xZ8uSJ0aXWi5Ti59Z2xOE1Tp5UG8i/Sn5dfWUO1p4VpVrOC9XGiPg
f4fWfzkuek0or5ZcaLm82JCmOt4KMxduoXsT5gXQiCZpUKAhx2vq7PK8Nvg7Ng13rhu+jQm592XH
W6gHE1wH8jDRWAsO1AOYQpjbP4itu4vuxvRPo2h1r0IYg9j/Ni91FIewjMdEUuDmCl8uXOmpPWHi
fPvvXLAr8l61uR38oMy9cdtW3uIYvJE5cwVbKTmSbvrz0bKzUyM9xCrB9KhKU4yfyTHLvZwqlS3R
kE6rz5SfOh5nUEn7sxbOx1dl3+Yx1NWo8aTbK2tv+ExrnEbWD6rj4zpZveOTOf6k+8yLjOL1kmfc
ZXqQNHNu9Fa89YhnsPQfoAWIPLWgE3P7Pwz5ZU+HRY5vN4qO6LvDg1mvzCCs9Vy+a1kRlufv7v7G
/F/2FgicfWgS0C2eoS3nYtRdLcGnGqfsCDppRAlN4SUq9TmjbOv0o4xwr7gpD2d+dfYkzaAqKLVJ
WfxLaCM4XeA9Zn+i8Olu0JBQrGYPjEoRqPcWKX1GpxJX8LsJMSev6zlS/fUEZL9hQezXCln4YCtb
W8Z3lCyYYA34mUMsROP9+u0G0d3oYkHjcLn69Ps/82cIeNa9Yqzojg9waNCv9xATBFoDaK+Gxmbp
mTlGQnlautYdqXF9chw1I0PScIgahXtJ/1y3MyIvYyqEPw4RMoBk7NmYpeRKh2a2Al/G49qJAtto
ZwsGbZrQmsgk2cS3KY2vaNB4wyyGp6M914leg9YG2ccjKcVpD/x4+9yVEJCK1VBW9rYZzkyXU+GS
BcUyHpfisTfDGd0YZjsWzsWTANn3J5pvThW/ftg6v0lqXW9PfZH2Dw6OnxWNAd1O9W4lXVSXYEcQ
ZD5W641YOIFCW3A9heOkZgnIKbaIgsVtC4QvqWv9MZ9lTPF6c4oV0Zx5HRPkEdWuiBbKLmu17m5I
MNp8BjI2khOwAUE14C9D1CCTpEKo0AaHjeoOd8iLqxEC4L5qR5FXSvRs+y0W8/2KEquCsBYzYIT3
L5eR5DiTJlWi/c4wFuIBbw/7Aw3m4p0cbk9I5Q5J8JSU6UXu6lxG4+Zyo4+/auMxMGhdn2VtH5sY
lvOe6pWCr469utiNoqQ02nl2r9Q0sOh3rfBjXQjLhvZznDgbZgOpTQ0jyWhcFz5TZAqqIkjV1AIf
/N/E15YGePYB1zpyQQ9XGz61ql0zHuHBD/kUrQlRTcG629LdylLRzuMoLd9snG1TPP6kX7rQ2mae
XqbWy8LPjaKg0/W2LxMOJYeDUOfLay5SfT+JqgOLHyX5fHqosdlOQI5g+wCZ5+KJM9V6cv7fsEAs
goUEQECkVOgA/QYBtQ/dmUBwtmKuDmonsNv4mFQrGX5krz9Irhe7mhaPGpkG1WN6HuGC9+W/alKB
gKPogLzAoKDRa6zQLhrB4B2xpeGiwMzGvivD0jPGpHiJhGAFx4ZZMq1Vk3pPRtm4spgep4FnYsjL
2jhjPcDnY9pGqh5Mfgwynth7hVekJsLmRPvYYmUMB0WOptEPW6dZKB/2sbh75Cdl71wNFyveDNng
ylt22ZakBR/bI38W3FQYBEo+pX0/rU1L5ed3thppLtkr5LNRNwGrgz8rEooo534Mx+ztuTAi/tpW
7zdCpqpaX+xlUbh882QiQljt52szqfAnlBFNm7PdBe/UsAP4nhCVTOWQVnAKsgMJTdFOhC5PJaFg
+p6vpVIWyQ5zrIVj1Dbk57I2t052sWsmI3eAhMSFjVIb8Hm6OPlwU+7Jg0MuHdlUeSVySYQ0J1mX
aDf1IkJheIPygEFbgvONWcZfx0vs4fMf3zBgoC0q8FfIhZzBQAGJgspgfB5XiBL+KxOkEo2JF7zT
YR2bNymD1WVj+EsoBz/Lbjm5ehioeu5CxbapDzQe7EKbX9xQ7pWsxu/k11qt5PZoHnB65KJZd0qy
qV8ZdIV2q85+wV7L2arWF37+KJVtbkftLzZieqi3IvxiSd/AEk0PT5YVeex/oc0hfbydQXRnW130
KQQRBs+Obvt+tQicI0IpZn7/IH0pQTjEuDe/0CKzFrl1cVqYyVOdGrwLdfwAFiw8XwpLlfXFS5r0
8x5Ana7z2fA1h14zrCz52r3OLIN3owXhiUCDc6Vos4ouS4hIydiXEwxKsApuX/rABk1UYfcQcPFb
RYvpciJ/jBxGogR4SitXW8/i/eWxLP2O2jm9dZ19Bl0DMA7R9wCPlO81Kaf9NaTkcD2PYdepYrE0
s6pAzmFRV9NQLZES8fT87/bKaO+oJ+6CaQk/bbL7XIUKLGzkfERnuSWig7rP+z2Xa+HpgclsCjRU
QpoAmowFCPj6xFRb/YdvCOLrZfphwP3d7/A5B+3fTQyJWq+HTzIfsYM0/Emf4rPs3btfmRNan3vH
433R+eBhWJJzhLC/OpNkAjEgGYNIRVH7d56k78QWnS+7A/iyQjgwA7ydel9jJ7UFoMVgJcGSyshx
78h67UcFZs0nK6MWhEZhvur4i0FWyD1bmpqEYkT3kkl/hYwlHopb6TtIojo2HL0cBm5hpV/X7XZB
CQc6w5VWXyiraPQ3uxGwR8xnsAEVNghUY6gyXtRnTHt3YOovb//q9uEJQ8KzTtY+x/NxSuzEBg1w
htoONCfCYSTMtBjJvyPDHld3Ic9IdQ+T8p0LmOw3MfKgPqviaitPgtyH4LgWnFxXqul1ZLu9p5BE
vLXQv50Q9J36IZChDMlQy/U1cKrb0xvOJHt9zBBcajwRW+5C6NVTvhXaYUZw1r5TiZ5CMRkNHRgE
J6E1wq7uf0eQoO9qMCoRDFXNXO5akeSDm6b8fRIPDNyDM3VaGv7xfb4WMvt7QS7xfRrjRLzdqSWg
ppd/08pxH7O8QafJYn4RKE5r5jgZmD3puLRSWimIWW35CcJxMbmhhuH3dwbNL138ObM6Fz/JNp0H
A+rF//aoYvdjmP2Wppfc0/Kk+Y1Ore+wMPzEXr6VSFnZ/nUOsdOYfvDSL3oaN6QCFBlLbCisySqJ
eIw3v4xiBJi0ZeDNvslk/aThMrg79WYe6jbRSK0wSU9KkM+Wge2aFnlEtjafQAROBFluFU0ztf0O
aGmC5Aktyr0MvbLX/i+Lu3VLxHbLee0RRz2XasCeXrr7JGB3HgnTKZ1lH5FmuWSYK0PVGqpiVuWL
WZQc1NODMFJxF/KnLoBotwl0JHGYaz/4OPYx0nrfuUdWH5b9pu82l3V7r4Eb0BMmUvzs2AhJGOFW
VjyYugqypmRSmbj/xkmBq79mCk10mNPkS+AjaPrBqymen4K4AXfODgkF2dFgk1OfMCRebxG0t6cV
blln4PSnZragIlzlXlug/ERJozQ7yLWAOhwyt4YG6N2rxMv01hF+rowBlUKf2td0SUmFgKa2i3bF
BGRm0S7wN6Q3SntydaFd7LYrvGA8W4pACsGdJnVgFTBwmNNod1DLV8TSxf0jY2QMPVSJgbfy0L6B
KPzs/hOPyE8YD7YgAkzkgvox8SwjeJZgeZ0CLbd++nIIwGMC3UsR3FGpx/kYezOuTT3aHYoHTQv+
vsk2X2ihiD0PZqWkNsy45OenCF071pQLAek+Tj96MOSN+g1GQt9k6XFSGQnCaQbBT78vbymHekaI
DIbt8kGnfwsEyufAYN+eQFDsqhfLb9sErad7fN/HQN9pqTtaoaowhjHzy5nH/rh3/vlnL+o0e6C7
TPkvJ+488R8RS/RlsIyu1/GXi1OJnkEIXlsnnZR89V7HZvFLu731ufsH/y7y1g1XFokd1WIuJ2MB
A4HDqrsTzMtmtbnph6f5gw/xOQnlincbcCFve4BmrbAttBmVNO4F/wuBUlSma2qNLUGMPA40SBen
9qKQijuWxnIDS6UABAPHTMXbAVv+DHSg/mZy3vAHukyhbi7eOuw08RJoxJ7rg9OpxDPAnqxlOTeU
arj0rCFzapU40FcJcbADpeRgccrhc72j8nZW92Qad8xhDfOrMRwFrVsNaBdUNbcp+yP6y1qIRaFM
JM3lO//wNFbc3xgG5MHjcARtlYxwvTsG13btv/WrrcCPFwILGGVyQ6vWGAo1m+Nscxko9ubiTznp
AKyODKX3g3i5unQvPBrXem7zJkCbOYxv+1Eoj2qB9t+xpcOyszZ2haNahILBUYZ5D4PHnyDCUpyQ
wuO7gnb55Bh+vTFzoyrypgvzeaue4rmwpxaROCsu83fwaBBKGfVcMGXCpeQGg9kUIa2TK1aDlnIv
TZt5trqtU6A5VHSMx/6+EK5hQI8ZhrXvIDV/OPy4RidA3vx4taDo4F+QCgbfnuVNWBjIv4hd8dKJ
QVKPrSwkorCOXjIdBgH5St5YrKhM9k+LsmeenrawuuzAnpF843GmNtsOLpwdbSxLtGjr0dQiEnZH
05+qYhRCSadqOs56WN+y5Ktlie5hlDDtad6tXkAZf74f/3PtVEBvOEYiXgwuPEJ7Hx7ZmFCCTSjy
Mazx/hA/HW2zR7dDiDbiAXOE786Z69uW+N2kbBD7QliotdOTi7112Dq6QAH/lw1rrF33oopHOVtZ
XkF+jCDrnqyYuXNE0HkISUU6Bh2GTh9vGvzDMc+KYmx7qi49uvlcbMC5VmOTo8VrnKcqmTK7AV/7
IN4GkhHhctBnhYzcABNx90cHFec6rUcOv5uhpRlDV8jooMHDzizRU2NqMNjd43n/mc65ngrmrNFa
+i+6kKi4Pbayp9aP6DQY1BywhIaQh6DSY4S1wEapVHTFXBD8tn/X41+TpuuaoG4IAY9O03YDntJg
X6eXahle/U97p5ZStPNBrcc8DPd3J5q0UzrNw0W9RBaV7OYTCuktjyQjslKCLjQn8V4c9YohrtLM
egyOU0bhtXB1UiDji9yYYaq1fccqaFQ0Bhl+/aiv9aSAZNaHhEAyQxT5+eZbvGySgePnsydj4yY5
X0Eg05hiGFGhOkux+DkEOIyBGMGih3oQqigvN31elDrcsSwNBXlVeXTxpk/MGpaVPdCn75Y1N4NO
6qG7kfmcf+RsdYB82J8MN2JrgIJlW3UjLkRtTK3XJfnE+X+gTKcuBVHKgYeptELf90J2niWJ6mig
8ROHA5zBhwy0IrE4wX8l51W8DbJmWqyGC4SHc7GEntd2WYY1FRYfJahOUt6iT1YapQzKyErZViDf
JsjUnywAxnoKcd1CbXzYqbakWxYSuQhxzAuS3fm2divjQFlpjOKD+VBuiGNUv2g77wDlSQ7Uj64P
yeRRME333fJWDJ0XcUftiQ9RWVPcir5Wlt1eLXPN/CSmtPkfiYM199HLE5e+Uucwr/rOAI3tsc7N
wPL7bBg/30DHgw9sVRdnWkI/m3xOG1Gsk5HmMDGWgnwzaYiZCYRH8A1nvp96lX6RDSiHjRREWnoT
/jqy+oyOyGw5JUrqBRNQmRDTFA1q1T3trsIMllKT+zjDZoTAKhZm+6fYKxgNUFJesOwT4HRzv/Ko
icGW+7Ai3TFQFXKrBAUq6lEA8ZKl4JpluuH/AZwO7TzgI3mWuTJN4OxRHZ7iChYmw2J6IUZg+Iqn
lKT1UKGogXjTNEd4dwRBGMzgc3vLrA4VwdX5Tv5OAnjdyP7V92gMipF3rn24L5ebZXVYNV4fXN9R
XIoJqEbYT6aTbtvL98GGgfWkOPnbisdf4nxrtPxeCRNpQ9FIMutsXNYyiG+/Voxqj4af6iy7Cv/M
op3abPXEvKM9vjerUZEdbtb1REPw7hlFt2wSDi+qZQCvOjbuC/00pwTwiXmmRUzXyNfv+/9QHzEt
zLjTw0TcF67Oau1WSXF5OYAjxSnTv81b/up71nSRgd9MbSyJ6Z4CdjCD8EOzCM5zxjU1t/A2/Ju0
zlyd8mRp2v49JwdUlt86Ncs94XAzfijZ7ufCkGWiCFXGZKtUxe2ShuhiRAihXoBQpRgYRxCrrtAI
72gOZJPKdhMIvhCpDKyF4IGrQeTy5ZUliGH3Z6LDaf/ha9Hp0jPp/CspnaJ6vvFr28toL4C8ifmo
2RwNYP+bwohRCCAb1+dQbTLslm7ie/2eQ8hlPwdUP4rVL3QQ6NLUgQRa2rCI/v97MgRvnSng4WSY
HHwXdc3p+WM799Uv8Gpp7BWrLGXODXI4SQSMx80Y7SMUfuhGuRa48ti8aC8cE5sd0AXr1szGkC/r
SeUPdgVcIsIRdSCTYN31zUjYUS9dJ2rX074eM8PgbIFqsNm+8774dXLNR5kuWFy+QXfva1wEIu1H
6Y73leD7zCrckcgSu+rYsSADrl+Diw/r9wj3/xqGVzvWJfGrSAcvIv7PMYgZxkfk/gxyzI4yegTd
dZqQ4YO4fiJz0XwrbJR7nB74XZ8QOPhaOBJpG/MRBSkZVwPTr+q6u736NihBQ1s+ChGdqxNZFqrK
Xa13+bQ0gAt9RdQe8fIqcdlckm3ML5mr/rDwZkpJKdZJBkR/hW8b0lyp1KwDW3ULPo+f2ynvujA4
ovTJ+X5h6VYPSnMGcRIuJeSkRinyLVDRxkk8YIACa7XyIof5BXXAN7jLLwYiIT8RbZP15RDJwtgQ
z2ejLdeesiOeWauFjXi6VA+mZieCLNx3omJmDkFTxV8bM0sO4igW2nGuls00b3yWtPoeyAN7GfFh
XP1B+ObjVjZvfrc1NPqsZ1Qd6PBgPyLafkusnu7Tr7PAkcmk1uE4fv3NaEa5A1yiKPwIcw3Mxp5v
XmusPULyNIapxp0QMiDUPn4CF0TO3Jf5aV5EagwmQArWjbOJWke7jTgulGYOll4AMIT/qW9q5Izd
o69TzcLL8OSouvHHMB/6o0pKjqCB0UmX/oOs763Q4/UnP1jOpiQisWMqGU0+p/zu6IIPM3P0hXoZ
Erdrp8bttNm9Yop9QDCknJhby55W8yZhMorLUPnigQ/7rQsGXy/UR0HfhqtPLvM6vmwsWz6Uz2jy
W+6xafMD/NRBLjdnCrL8VbcpfLe6Ln3p1rT2qQsmGEfgF6CtEsR9uKKUICVLFowfLblrIXOTtBHk
i9iUIw3PBwYL8PUwg5cG5m1TzibIGPyzgIzUf4OeqW05wsNOVgd87bl6cDiHf1UMirRq0D6wybj/
IH27x+s0+pUKoBHTV+wkC8BRi84V3RaW1wjhPO8fV+5Js6KQBIWbmx1q+xLsQuy61+WDhiNipb94
pURgmJDWcnr5jm0MD6rwTdSTrNAGx2g+4h+X73rGvZLjYOXkRUjtsSdMfNwPbOvOnDHYyNYdp6u4
W+TVMCIs+cq1wl3v0UC4zkjrr7SfF4IC/hFUXg3e1XPblFkaxgytjkPixLt+n8QtzeI1o0MV23lD
3NW6sXSDK1Qk114te3ATM4K2Fb7HOUzt1kD04UoevgWLxbeG4iXpvnbvg1lzL+bFimV2R2mvNai4
qL3fnCE/LHdFzL1FRRbVgiBg5BRGRSUqz8AUtSweGcn0xMwZwMQdcvofKrD2hClLMSe3ifZ86zbN
G7IFon+GkyVZsJ4Xji8Iz2YaFUSfU3eeStC0+RI8jvXPTdOgqK04hU4Vs50bwkjCESyp3YaMqMWT
yGjLoyWtlFqgLEosgAkDSO3DYTYnkSZUIQ5fX0Zy4iZd0At+uneqo80PVI2PAeSYbcLbPbO8CDD+
2WP8GZ81L57Ym0dy81BXDTvO0fhX7+gB/runmHcDrSl/NJ7ckogTrL09Ay4c82oriB9seLXcSO/o
bG334aEaK7X6mqev1S2CbZGp1ZG5B8BJGbgpWFXdK4iZd8TjJJeyR4iQQhFvg8rNLFRyuXow5nSU
TejTWaBywtXNyxLU9t9xa5PSFOkygyjdbBe+tokcYeL1dEiffVWiiaAnGF9QZl/6d7PMa8oRgCvp
J6HzMtImslMAseyp4ImqVJnxHfrxyGhuz8jMqwZuXDNcU4Oky9nWxw8JdgOmLKeQ2nXZf8QWEyqG
TuJLj3B1Hkcs5N3FrYbWCNHDDB+iH3k+Se3ES+RxrlezZ2i7JhV2FPEVRa912xVBYesy+DhzXizS
wi00A8ToIsNeDaUeCqihAZNHqzziSTupTEz2xM3F1DkeEV+gb0SdZUrfNFK3yu0UmZRxna9CTbsz
3dJM/Ws50SEUWS/dXoPpF7kXAJvlSMadDSodSsxkpmOHdCOCTA79JXYJdAk9en1MYT3vsoJuCeOC
jjiJzpid3TKqocFf6b3UG5z/1xXYY42uPiFGtSYOfA+rPHMZzxoPJQOXUnLwOpSOGEpWUvo2Q/6e
0ksByjtuWupAN+K8AmytYsQw021BujB6geoCU5vvw542RtUoK59gBVWNHVLEvo/I/SOcySbaXmtv
uRdmvIX9sEgGK/mYYAx72mezIzpkm2ImDMGQQC0WWUrC+hqPnsaMk/qjRO+iUX/isvRimSXwvOlD
4ElAt6QIRxvX0Lmj+byBH1ie0TDiXNYdPitBkYqwlhz4qSw6J/Ifzke8K52zOVZ94x5xCrM/oiPq
Kxgs9VSco1CDDyyk4dbeZ/XUin3RiE9OPqh2hhfuxmWMvrajR+bm20PYrWKEWa6utqpUXSkwyfOY
uOiQTGHLLstrj+xUoAr6WCnf33niI1+7bjAUbrGpKh4Wp8YOG/up22YyV4yRHnJubV7DkeYDcisq
YUFf0i57larjZdLtVG/4wAiXZBc5felbqKwEdlX2znzLMqhqMchgxYATT9VbKuTzG4RKMTNO3+y8
pLBV7LnNPYNrm6ZOVWmUe2ZiSKe1s1Ll8lENHmTd4o9d6w72sYQLDL6V9LZuLrmHfXqAlIgUf5pE
c02GTiI6oe+0DXdATDwlJ6S4I1iksO1059xv2kwF2g8iwgYi4DXIlmRQxTPfpC+LmJtXwxriqqmr
I867LEuAm9Q48jgRvO341cRb8pqN4dDYOGB6mBpMY1RGym5tMFnj8Q8jVOsWWCfwnlOMT0o1Qfsc
ip5xMISxDl1p5WPNccaImwwYsqoenwz6w0FNcSTXNigroMmYZIzhRv6XFew7RPUQneSo0l/tlZt6
o6QpGDwwBR01mBqCSHs2zEF06tSnkbxO0y+pWxyvXg27dTK809ndFEx7J4ezlk/itg80xURk4sxH
JdRHYTj86wb2lVZWiu+piGglcO0jhw0ao+eDtbEveIX1F4Lh52yfhXImG4j9IiIBvsrlX1P4/UUK
kPEAYhdbYT4f2TNxs0hNUV/SsZARs+oykoT3fjf86voDlZxwk7ttlbTs37AaBFYHZ7gr/zcfE+v4
ADDYqYZlHLq3loUaP8L38eOgwZ36SOWQYXou7fqwrPFhreqr6A+yBeg2Elref5W+euBcbBq69Vlu
+pxmfZOO9pmj55n/rBDcnTAQvnD7kWRzd2CdB/8b9bOwJVQ62GTg0ujrRR9uxoRUsydtFyb2z6zH
iuHKcVwGNx+hzIg2ClrEbFSogSzUBnSohOb+eXUkEBJU0JiflDYWc1nbQYmiODE12U6O4jUp3lUM
Ej/9TPCRrSvTjX5BmYx1Q7KZQfOoHn8kVRvC2Jc5eQjyztfinSTXWpfg4IUM9aA3ihZWlCn/O8Uy
UTdsePqlafXQiuy8orQd9znIPxHR2Zdo8ugdOTDGFEQ+E5GKHPhbStvGADwYTJo2IRYvxi9+DHxc
HePagaxVghe76bHFbEMmEfD3XLzz/W9nu4V6gZ4bmb5NrhymZ+UCGkDez/iwYLxrb5h375ZD9SPi
e7zbNuFZJ5H6AabPWgKnyAUgpJtByzDC/Xo3pwamIcuhhkzLHxu0u6Omg2FkxBjm7tBOLtrmEWYA
2FQxbELKUWYS/dw8nJe3R79mWh7xgeEuTThEWX/omt0q87LmpCjx+EqmjZb85YHMU+ZAgmJ+DFXf
75gKTPXq32iBPxsf7TcwcDRhvRziR5mBUpTgwisgKNH3WuJItOdrVbFQX42Ct4Xyn5xLXTEdgllg
BexjWUrHeLhQl5uZx5+D2MEQwGbWprYR32nNZagAXZDYiaSeAiqDvUXY7Km3fGSpxYNrdnIWVgCq
jj5AXtnCwDkKurK8vhlu7vsJ1byXj9zo7alhgHsH9yK20OIfT2cruE6nzZwlDoK2lIJi+7Cm0k4x
HHM1OL6JuV/5V+5pqdBj6OwIDZDK9v66xD95CCbNUxgDvvGbZ3tiUPiD6xnZI0puFyoVx3+HJhnn
x0MTZaFO1r1ZcGQlK4C8rIfH7QhAGXglisOG+R3G9+XpP7IKO9GYAknka+3bFi53cVVlLezwMiBe
2pC81JI4eOmR1e1uzkPHN9LMq4sadZ1V07IeXofUYs/faejZf+m96KSrVfXh6+LyEr6iXa18RRkT
ZYlJDwdXqbmp613DM+13btovkdvzMYB8GNWL76kZTmTdWa8aQbOBz5NqCmk/d7kKzW7i/zM1NFd+
3oiK2IeJdUfiQLdWt4FwnVQdWv93fSZ9rPPfJkaJ+wzIUpjvFpBFLHblnu2adqY/3oivuZ96A38A
sWadlR0TT5nWBJZvW/KOJwnbRfECErpGVM3cGDv4Rn4RgsWfHYJCLeNFT9YYZ8OQ52xSjOm/XwUb
00kpeY1fAY8K8gAdLID4mwETNo+rxdxnqmfjMzeC2yKNWM5NqqwHXTkx5jwPi1UX4tuKROcHoBeY
3THMCZbR2taFZ5Y+zziDqeO+2S+IRTbSI/cd4fNXo6vbnFuYnU5hSgnSrwzhJvPOxXJUV5Wn7D6c
jVHkXOQxNaLDzWUX92nfnLr9NYDiR0OlM/yJ+Kx0HAafYzylla5yBWz7Rqz5rWFaKD6OTuDd+XGn
Oi/n8YftzqPT6ejJJLfW7lSpEvCV6lNcBd2ENfy4C0CmqOvhARZVTiJNMsDV7O8etaiDndmPKMyD
N4PU4Rhwlr3FvklRcv0MaHUp1ozU+osAVcIQQq7xfbqlVBvmgwR/Er5PxuqtdCI/VWDPnP4Gck0e
7SnWfg8jtNvvz0J4uuRxtMpgo5hl59HRyj1o01sCF9cADzthe3ae3EqFbH4cCshndw4KixwaoqZW
NIeBh8iMxgg5jw57A+NGsI7203gctunSxkjWMkeGSqQzeKCdv83NP3MBrzYgL0ijhrXcHQNPAGzm
2nr1+pmdgda0nPpB+fzBfxs0JGwwpTt/KN2F71QZE8VaTvH61XsJ5Oo+AbyI+Je5NgANUmOeQcrw
IbX33bhP7W+jNAtzWhkW//wIS4XurPjfYBG4eN1HMP2IyFUxNkkV6i1Mkdt9FNZkMgYK7q6P3PQm
WPIJsyd0MZE569dj2QCM16cn5F7n2lIzcDXcg4NgnxhxXgAHe0f/UJYqraF+xDKmtTeXqwb06EfR
lGZJ02tbo/0Bd/Z8EBIxV8zzRRdfX/aj8nEUtG2XZzpuNwoxmypQyF2aw1YJaCY1NRKNFM2WcLA/
Br5WfrG6pQince3Dy4pBpd0cpgrxtyh1G64EjjkohTScwMZgS2rNIfiFCX+34tFlXNshCwJ0okkO
SM02+J3p7GqVhMBziPIBIMFli87uKD+i8Dw0NXiKQlxuAoT59S/rhSwoXv+zuJp6SaB39MP2HVYY
yMFR8Ay6EymV1us3oJsYq4tooZFW+LYUje51xUR2L5lkTmTPFmyDzwcRXV3azoWnVMDojGwMJlwp
Gq06JQBChjSXvcs0nN0ntNaO41ZPO4IsemLp1SR/VFqxU2rdN6sKIJaE08iqF6bQhjUXONaLJeiP
IEvPYIaQ0WIu/Wm7GN4v2/hjnnhDuJIBXMQoFCt8fDYlStBslwKD9vMPQPbFVSl9uw8FB/Qi7TJm
/vGavPJU8JJPSkwqZHiCPcxf9k8YirVphNFujA0+EpHInr9X49MmYXvURCupTw2jlBFZ9x6aNitd
PuONdeXRsjVJgfz6iAHD9B1BGHMIUG2/zluNCbUCd2UET1471PP0afSSG4zG0PMNyKgTdWM6NNGt
eEFEJpcVD5E6mLmsDQqUSGG36I4K0UhntPhZ1IY4j3t7UfMAVEYEg479YKSKB/GIsm0Zjh5DPrf2
b46zok8rXt7AgUMn2KB0BNGOnEGRVj60s1F7DrCwfF+WsmGBooRGRz1bCM+rXQGJuPcu5gFcjruL
+h0jxWbQzs7hmOAj6axhWKWrW0Ugm704FltYVWu6XEq82/pEPxyDlE1LEqvIn2ShtNBbSMIju4BU
oo2Vo2M/wddE+3wJaUkYqj6hNOv57mbBOpOBBQwhC6UcKf3Z/cTyYdxYXBBBOgpUXxgw/A6U2Qr1
AJyGNyMdoNB95o6rD8eWWBJEKElnr7AC0Jnhy3DTxwN2SACDVRpUs5etm/j48I9PM2G4VPF6KWyy
YOYnq62JcPYcmLXe+xtrzWz7lbq2aaMjTFX1p2YjqdFvkY6v7jMSL0QMtp1AiKGjP6Y03PpYG72p
z1whIi5D7+b61AIo8pXMlk3eTFXix9xfI1PEBMtymadAnF4nXvHPkQKqRQwh1nPZd8G1WdC+B9Hv
QeDMA97HThONSaZEBbmb0twxY7/WyqbIIJgccoCwNb4APnNnEsOXj5QBWg5DImXH1tBQQqLTf4CR
HFGWWtIe2CSs9I+uq/hucShL0uBotzsHmUAcqOpA3KY8RoVkRhvm630mswg3ipxAf92rDLhnEDCr
b2Oo7sCNuHXyOjp5pQc1DHsXK+oSb5LEvMbf/kmqMp/M1g++EtPpDOVyqbnE1fx3dhfe5rNc4nuz
FB/M3jDf/KXjke4X8eZOh554S5YQ00LkBZKCHxldYgVkKimwBp9dMY7xwK2GoJTJQ94oijvzbR0V
Oqm+eVQxmQTTvSmDZvdVhou/B08+qmtop1e3DCo0WDsXVhiwMvTun47KDyaNV4cw7JuLssPI1rN5
ise66F1LfT7QCJXURXW9lKy/ct1tX+Z26HzRkAUM57+pRgUlLrakr1odu5VGDw7PoDg0ohwFDycz
j9tixR0z0oNjiD0K0coDNn9RlOz0HdbG6uhgWjokwg5uzEcIUta6K0/ycp5ayDDc0fSySvvEuAyc
y7gPCdNOWg1ttQNzfap8JhhT1of8+t3C0W4si2bmKzNKuVTHuetkuIY+a4hwikmL2wO5J32pELmv
tcEktgNbMWnx4Vw8UhKYII/cbJUtbCJXD4eu1G4pZlGEkTqfxribyzG3H1m0R80J/2aJCRemJH2k
uO/W4ZtDpbCJ6X5fb0eTlhRi7BY/cMMgKkya0KK0040K/Ia8kofvsJBWL83LaWdoRFzh4PcyAy4t
cCJZpwCC9ry75V5PclT7RW3/skJwgGKHQj8167TWpzJqPgm5WtAfoFcx/9CkWsrBDz5cgf9lgOSm
LTgkdtZsRwwr8FqG2NDo2yQHtYzhguFi79AgaYzNsNexp9nz3xhtiVPy2TSI94ArpCARBlz8EltP
rCzoFXle36y9z3s8iUgaySO1bSS8RMMcp/WyDoLRHiMoMansOXfcwl9N21PRKKmEIcNw1SgiDnz+
HgYPI5HqUaefmtjARMMqenAs9G8lJ8XJCzJd3vjtGLKBJD6Nnr0Pu/N4Ny9dL8SIO6U6zeOSyVgD
g6T3ks3IyaJsryq4A1OUyan27N5M7b+idwa2FE/kQ9d5lWv6A54qUDaOeQFTrI1cvbxWfGDXSfa8
uM61RiENduuU6beGw+qeY0u5TEccV1GZh6KDgNt0z0YZUS068DUXWqC7W5JB6uBtjKHxljZ3+RWY
l4+okou1Fkctx2Cs+NOrThULb1TTz5qAyaq7D4btrvHfe12OeM3oPDEw9Bnb3g4aEkouUjAPCb5X
NteUdvq8QhVBTKNUFWWbwv7SX0gUgpsNyX4K2aZpMPJsdGImwv1EFxywiW7FTUZ9pz4ARgS7ievk
ITBYms1g5pjo9I75G+nOASu1JM54cD5w2aI7MtHUOoUguOhLAAdM9txNsgB3IVqXMHvSnsDJJyi7
knuTT6T3DkTfqYInTyxje+7wZ08BpCO0/Tbs0UmJZsoJytPAT2vN3zl6MMRO7V6428mlu/1EOrmX
EnaUUpjvGT0Ay9zWsZbajMDpKuQ8GOsx2K+DZzWzJbUbyR/3oFkNY8PhhY0d9g5OrCL+CNZCjmMJ
OYotU5CWpRbOYUc0XqYju1uCVCDX8pYTpPInOUeuTiEvYxE8vl0t3LXKOYmcAT4kzTRGhCFdU7bd
UE9tEqysPuGU15BraUDnR1cL9BucE8YMvXCGAugfRWPzQc3Dd7AwRkK1LVGT5cCJ5bcrFhuqAltw
BNEIfFIBhHVxp7did+3hEYf+CGkPmMUqVuIiR/nLYqtSVCub1J1q5HI25XMg7ae/1IZko5xr3yLx
K1hv47kkTVhPaCCPaYMCNc/7YHloDwqKpuudqXjEE006M3FO1eJMDcIeA70Q48tEIamxfKh41xbJ
INcBKzGaA23KWcoYK+Xl/rIvHTZTMKOuN28BErwTxbJRjyINxfiupUAYvz3l5SUSJPjTa3JOn+ZK
vSZJSkRMB7DNZNpJBFn2eU9D3jO1hm8wJcfkD3QAliCECoB6fbz2JS37OiXglhcliMAo5B1ufO5d
PB1woh7bc5Lwbk/FN+fuw5YP+AuPfIq5GuJM/NgaHu/y008VOaeWkLXvdUIQYV6Y+qCmCVGh+Qna
tyldvAKX47mzxWQUDvRhB7qMTAD2yGnJifze1FejX7/MImzjBG/QcMF+86WOPXYUHwpmpJiNcu67
xVvRhECpJWCRfnWNp7SvXvcOfLizZ/vHzpwSFWuUzWqoGJ4jlKOOZ+ja1DV5tuKuMYAu/uj1M+lg
yQAr2rCntvQ2gnn8TkqcU0FUdycvBkgQUAp9W8mecDAfI41vrl1R3EnoqMFrfyWjwB71OoWZD1oh
3OYR01ms2qXpfw+Q6jQYXrmLhOxJ/T2M54W90apj7/V2Yguu3t83AsxL6W74mhDNOX7lPRNELql8
WCLjcA6ngjGRjq4fl6uD0Tnqf7bX0wqYy+8P0DLBK9mXRoMB2LVQ5GsNfysLK10lFW6GF2Kt7YE4
vSHU6Wnq5WC5ypV6M7oT5Rwu7AMuigmtnM0ErIs5koJAkrOYMJuIKuuq7yfy6rzzb3eFWZd4JqKm
SOVUJ6lVZM/Bi9STcYplPaDm5aPvMz22n3/f84UKuooCb5karO/yqtZj3Y6GwyzlCYGdiNE5Y/0u
3VrVqJxmvC3NdlyqzeL7Vf3W6YeFmHkwVyoA65Ok4u1DR/0n21lzFBpSmtNqAFQ6pDP3h+hrxbkU
VuWiuRhf9aGBneMpcXGN1D93qQ3DO99RCeU/zL353YHsl/gsYC1dktBkqr00lFnmSke59xgSvck4
SYoeuVL0Pd/hPAWGGHTXngzj43pBa+v5O/B94ZfJBa4UXVkCDJdWsftW8NNDMHH60UawdakOBGbh
B5Xy/e+kbFU1mUvwET8E/W0z1hQ8rg4VSuTE7CyHCbnrl+L0Ui8/JdKi9Fxxfy/KekWAGT7qB4G2
BQE7X30mwYkrZXlSGzqoiRBqGpyiAFZyDWYAZE2n+K5D4al3kmvWZnT2m3hAQ5/Mez03r4uiwBPt
uMPdX2Smc6TBWHXGXQ5by0BmBHb2+puYNSTTpp7j2EUONnSnOIm4/m6Ofgw=
`protect end_protected
