--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
CrIBTvawiDCvcFG1ygynBtppYBZf+/SK01oDPfjqIqRW0f3vpQY5Xt7O1T1vRCCB4G3tpMejowh1
YIuN8CJT9iaz1Zx2lnrdbJEPVjiftJyuNKfXscXY9Z6LQKlWuvI5aYxC2FimE4JQuX4zgOnEXOAe
Fh25tjuAfty68hRTHTCsj8vyTGiLzMjFiO48Db5txHihjxGqbrF2+yw2yP7vwHzYWQxNgVW2re2K
fekjyt6I00CLxqEJYi7aOQvDqGOMGTXEIWfhZ6yaSYYaFSFEuFOdwViR+KFeCCSv9YI/4DdOGGLB
eFf68ZSxXRwXPFHZcVsUumCMeF/BReod70bn6g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="P1SCKA6T+U2k1Iykm/tFEvIy8nruMSm2AqVeXG69e4Q="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
BfWACa5ZPUaVCYxDUDhM8JKFfzBiXRKP5bOplWF6UeUzzEUMlVfXQZlgIfxtPW8blh9JvNQEZhZa
WHLPaf/N2t+9V5oSl8po7XvvI00lbjjt6x8MQHJCXi1UCxREcHZwrIPk4tJTSFKs0AHamITx9ssH
JnMmFBO70PwoiE5MfdlGJCIwb6Z04Bv6ESXJyAgXFwMQknso7BbV1Yzi/E/EV9xR2w8jyUzfUg6b
dV+GCAz5uldu0q6fYGgPy0PtElTjSU6g0EhXrXSvfscdFfA9X4hNsqZ0p1JmqUItGP0ZKv8tuN2Z
1usTGzGC9YRIQfoERMMKblzLRsVpTil1ApH9vA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="59UibiSNtXOzv/KUdkdarutbihf/1TyqcZSbPvR1Ld4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2544)
`protect data_block
Ms8wOdBIYumGIkrG7dhdBRK+YAK9y6m9tvD39uJJM+oOKyYchNaTH0EZGGG4jlSDcYJiGQbK9rj2
nz+ug5VgWmWSLFjJdH01TFiFYHB+Y3OKB4ww8va5/ppJtpJLxOQp7iqLiHZJiHu4ackxFh8tw9fI
LnI08MZWEUFru96tcCl/iRGzuPzt/QMGOdwAjJ2uaOPyV8X9Sb38MmhulhqIQ9r1qu7Y6KdlNtca
rMhAlGvptLO0wMeIx7fInM1s4anbFrzeNBYNidkHsrshT+Skrqc2JL5TYxdUx0iUGHB7SdVUWghP
FdWg70UbdAbEAQXttOxSUQXV0Cavk1XVZ3q/qJYZO7RL6meNja2QQENMbcjw86ISaDYxfpHsDFkR
UJZc/1BsyQQ83uZrOk6vvZbnSx+M84T/KFv96m3Pv1bP5tfEMmlQ7VkFHnjln9+JSzJznszZeabr
/BRwfZNO6UO2Z5d5LXrmA9nyZ0htgSRiBXN4MRFOFlFq7fK4G5SU3J7VefiUQP4fyNY4SROgO6aC
GbfV0K8jduuoEcW+UNtBzX4sHnqm0UtwvHdSxGgUntc8Zubme5yA6odKuf7abamL4N9Qz3DtPkC0
Wle2Bkq8d6d5X6HLnOeqxWvzc08Vgm6kTSj5tu0xwOs63cAm2rorxRz64M1Nbr1NAzbpFgASsiYV
0AHfYScJogG5m1Ymv5RHOHdr3gUVhJixQ+5qqsDAJGJtbJxJu/ScGbjCQ/qSS584Dl+brEmv4dxr
+Lvc93kjryGeitZ3/KwXpujgCkqqWYjlMbaD6MPl1o3wA14cdlujEvaPnM9mfIonF54EE5b4Hz7U
68rVdlZYc1bdiXU5/8zZNiee4szpN4XPETTpgi+vOSPKFfHqI0yD5k8JHbYQY1olA6Yb/DVzpJx7
/rMQRM9XTmcEtWfJrPGkxbmenhZeGHm6dpEcDmuniHqTAjN0PQFxouglMSlUYwSKq3usFwV+VKMV
T95fF7e3hCA3NFcX3CaZeVwzD57ii93zuEajcMZG4iW35Hn5BxEQ+QbseHT9z8cDNhA4GnZ3IBOn
yw06fzpKa5XVqe+c+Nnqn8DBTwWzC76aHX6C+fr0rRCkpzbUnH3H2n4CIEDK+pRvONhGGESnq4KS
c0NHo00Fj3R5n1IcCKj7W1e9Y6JsZy8/4cn37QHZ5IAvTlq34e07Hu4ceOSdhgLuVSBY/Z2GivQ3
qpe5rlhU4Kl13HnDh12lr3YeDFwgHr1HNzCAVVZKgRWGeDrCboEmzB+nXSxNpW+02pF95G7Z5RUz
sGKgQoLmmhBbN4NSRa65XO6kkGWzSYLZavqAfSuuSdqYo8rNWyGmaiSopNCvHDheympVbjbsakvi
T3bxjNEzfEb2O+obxgpzF02zgcNP8XiBYEXgXFQ1dcwc9MQC2L2oo7PlXMqvrvORRY8+oC2psgMH
+QlWsWjYpc6k0eaWYooKS+AQzhSSVsK21JDTCrjZnpNtSTjzoOY0GcGN3JlUenXA0uB62O+P951z
4qbQ4E9vNhTmHIYgqXCMupKqAD4cSWdLz8G2n+MqZ+QRdF5UFicvu0w3cEk93RBIra3LSqMUegIz
39HOj7IYymP8NrLHL19eA4t1UTvZBD1fLfhi/02OY8VDMk7CsZ+/tuBgCDEXYvV+1JNFyCLt/rEx
vMMb4japDEhTsjgoTgSsdCRxJ6pgsGTFpqCulvJq4AO2/Sne9fyYIP9byLN5fJyKr9SE0lMxWsTY
8MgBCyZZj91ocsjmakZNe1rXHV6PCnaLvHP65x1v/V1arzyOqen3opuDStsH6jUM8TMBan9h2XEw
hSjogU9dOztc+kO/qMyewzywD0Aw+IxSNaxBwNn3LAf4ARQaabm5ykCHGVFMD49yGQXS588lp3QD
Bc+cvcirY1lgy9HJELId7COKOXB2HLd5NI7IdTxp+7Cfsfv0l1mmX/nESqkfFvlcN1rbvM6eLMuz
GK0qEs9g9pgEI4voGYiD1/JJaowSr7lp46Rk+4K6/Bkbt8sCoYa6pgDtm+T3eOWPnRNJud7zTjjk
pZrVb7mjYpD+ofL/KPHGjZFJqByn5Hgg92+Xoxg6dK9aZ4/MwXzQZfZrO86priwHBgPJh3XJ6SRH
vs7CFxSuTpA4kPPYJx1eGEN/ZK80KTNuCS8PE1E777x4OAvFrE8KhDFmvIZ9UM6zCsK8eYw06DFU
gW+7rarTR1UYXPUtRmZ8z7splYP0Kg2yiaQZgHIw2MDYf8FfaLfbABFoUVwoh+o3hHGTIDS/c4Dl
v7VvaM31OgBgOfDyHU12n9wx2sWvqCZc6jH/VPbTLMTdJA2hZZsm96fTOaaipFwfu6wDBqRiQS6X
Tr6PaZuOgdo92iXnjDw/CveQCvyHlnIJuJcwxujZCducmtvY/+pHbUjMMVIrYREwSvI9qI0D1sc3
E33mUlLgCwHH5NAjRVAF4/OiUeVFG5kIn8QmHumVBe5ozgDQghsd4KBEszkjFv7aafZr9Q7OD9dG
MYQx//UdPORyLS/jrvBu0qt81Le5EMej7jjyXImmlG1e+ejKj0Z3vj4sUocIDTLKWEiIcNkdz4x3
WJRp549L4LZC2ZMYAnDYEPGUOicrsgKWtZq4VPkRtcxeeUwLJQSEBwZ3u0hHSxm2gCu4SMWnKndq
pXOBYujGz06P5qvGM6IFZyYq7YN2F7wZoZ6YMgvE+kemAzssohzL+dHxiO68lXipNoG1Mix3/uVe
EhyjpXkynEdZ64DwR2WZIr/WBbM1UrY7yUWLzv4Mt2G5Ee7rKu/Mv1l7vz5UIhVZ2aKw0Z7E/dqU
/exQElzcFtaYARaQllv+8Hj3XR/zU+4kbsRhwA79ofd8lQb0ugkipFgo7iN2Lot7Roei7Oa4grFv
06Wklp2EwDvE/FviOQqw320f6MSltglL/n7Pu9mi+JWtIMQA6v515FagBSmLMHIKPocbC4PJRMwj
vLWDE94W5XrGLwooBUFgOtnalWHtlbY19rg8tskNk11vt0v+6sUcIzTmJIWPDCZNeXck8GBpCefo
EV1rPs+El9lnznpkjPDbFHHo1VFVqb+Kk0oF7pQWGdpeuOuClRqhryCXK1K2HYcTMeExlANh9M7e
FdxM6TCJia3EKabQzkkhq3Rsqx8Ctw1Tjaj4JPUWsyq1MlrNDpxXXsWr6dHRX+DBYzYxZHXXIQwa
iLcWg7dYrt7MabvPAzgi/o66kYi/1TXOfbmzYTLXXt4DW1gBj4Mzp5GSwc0OQaq+fVzlfScRwkSr
aMsfu86CwpqnOdOhjJqQAFUoyoQGpp+ft862PZkqJ2GWZH+HVynRfa84V5vDNKauxS4lePWbTsQn
ZwdnMLpm3vmcdlBX0UZJzBfzXfwX1r2+8IVUJVCjwqCcGOip
`protect end_protected
