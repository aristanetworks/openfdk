--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
iwhXmrSfLBp93Ni8F99vyfY4S8MZ71Vw76JH3uwUYFV1qBMGw3sg38lJkydN2LAz+KmBlx4jhApn
tvFsidx9v+OdSLq3FYz47CeOO8HnWXq+8H8LpyEKf11rG7vhGsDO/Mi/g1oQqBpECL1qH6QLcy/j
UtUwM5G3S5t/EgV6WTu7tTNGlZV/bymR+kGP3TeM7aTh8XxK9a1Rsi2Dn1KiWqw+pY5ORzkDw8mT
fiWg2tZK8daaL6aggdudkjrbN4dCnQF1qForiipWAAAdnAwSuzZORtpzfJMYuEI4lx8z1B4D14Tv
27O0qhKSKw0oNnbblJmlT0t5V8m7j/K4ba8aAw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="2ikMHMrWaXpz2kQ3kmLnKJQ+xh9xWHIlPAydaLZ9HmU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
liFxthq8rq/I0BJID6mOcH0ckwjVZqsyoDvti1y0O001mV5xMi6Lxv/aFwj8t5NeCkVAQfzJz500
sC3k3w6nuOzWMlpKUqBSq9g7sxn1Ro5zB+wngfsDSqDbHqhFY2ECM0MLQx/Ywu6UAK74qY3vmKb7
uB30D4MwFMsb7pdeu8d0GXLq6wRXbV3AVPs5e3vKEWtGCqRemdRXERp2e4iqfOqCq5Hp6jKeJz0E
+OlTGxDuOfZsehnU3qbUPAVHbdkBrF5MC9Z3bkup7u2omJouwF9XDjEBYFjp/ySeVImE7wV4T7ok
9sgVFDPtzEBkKj0fH3JGrZWe01L1aGmCTIDL4w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="3I/EF9kLWThB5OUd5ZPck6G7AZOvPaaI+/mlSWTLaoQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8688)
`protect data_block
rudPT2qLbid9efcB7rjVTuSTwF41I6Y/5NRhSdI0W6ZtEqvKLBxgjk61JMRRkX1ZuEQ+tBIlPLh8
up0xkpB9b/9eU6etf6dA8cmcPSig6XVhvXK4C2ilvMJzbhCFjRgGklVRl/p/lIFD/ikR+wLjKoBI
fd6Bgk7oBu6PFMjLnkcTD45wnAFNrGwA+NNCEsN+hyAH7k9crHA0RdJqf2EeohNMO8+X5R44bFOc
++HTNo1lV95ODzn1MweTnXqc6XISKrYg+5QHrc4itNuQletO2odzcP+9bCrYneP7oqMnIFPs04j2
oR1rdLOzIB6H+4//fiAQ5yvVrDWcXJfUadnn6WbOCERkYewFaWYrTB1sTjG7h426xhpEPuIB6Z5H
C5Pg0HMxhI3dBzHhYmznB5IB0TylIeZ/j3+m6gCZkOGyskcMn+3bjLzZJGS8eTGsaLWZpeWw+YJF
41JjQjhgc1ZTuWbRw0IpfH/Sp3JXyGKZArxnHtcEysa4gXY6Ayv7yZlsAM1F4osTHErAIABLewHU
Nyx0cnyJljYCcGoPgg2c0xXRWlUGyWGzv1Y/b4MtZccqCkyheqOyJGmHR4NG/bnvDsM58vyLooR4
tyAflr/WkJVis9yPAFdt9rmhQZO9V76BMxJYDW6TxnUeM6BONjxZrxkHwyoRA36q0zeGDkyCWCJg
CqGrA3fBZWUL7jr0OUpcR1iLSW/j7/+pSDATV+RhiRGejSCz/vErWcBhCWehUBKaSc355UFuXtp6
5v7txDQ0oXgpAIG8oPODFPAqIIQ1gwrhfplc2XYaJ7kBRYOYjLt/S3veqerT3fEUJK9TyqupM/KU
eiUdREJeOV4wC2Aj3i+D0w016AK4ngNvGVu6punitheG/EMqy2kt7n9EDGFRRM06L4OOOsCWL1QE
GWZ1rqDS0hg7nciJhGdjNwWsBKe9T9vcg6Q5Iv0P2zirDM28OOKYb2VwIs9SEnbhemQcU+8oZpRK
P4xihzvn8v27XvsWzlYw3Y6pwwudbSA9wxfJBfab0+Ytd5W6ghM/0rjG322f+dgR3IIMdBTaFHVV
uKbsmoHFLBQY9ko5af/GMLa58u4jDIRH0oRwmXOF+bHiUc6HegBUxX5NIjsyazTcR49Zx0Tb/RYV
TLrjAWaAu0hyMFFPjBH1W+vKNtKMPrkdrO7Xguyw/u9GZiZRWWmRiO3UVdYAEl/HGtVex5+T/Alo
DS4wu9WEG+xVGuoxDT5PeCLUl3sApF8dblVDD2EXx6ayrVL3At+Y9ahz9OjH/zDQL0kc0YqrQAGr
isOP6T4852+s81y4Fvi5OHhfEePVhX7jyZFaowbc4O75cJyBhU0dZFliaM2QA9WcA3tNEidqatjh
NGMLsW7M61le/njpGe6Urb2TAYwCVNRWXFpZzFoqw3vejqkdQGLLyyaSqfXSUsPDQ9rCkm8RWvnC
CCjaW76LBYgzmqCZjCI9azadXUtTlzy6E+mKB+8cB5tHyaO3LXha1UBfV/gQk6nTFquS6QsYP1QI
mMEp6HOz/vCsv2psCIPxurLS+bBT8C/N3OfYtpmdV+dDsZlGuhStDyc6Uino//3fisckqpbocA2S
hyySIqzknLJuYUA2r3TaOHlF4EvY40AO/nJBtJ/TYirhd5Yw/HWok/XgERpagWfD81CGbMVqzm99
eS+snhwuS3MvYUWSFmNiRDBiv0PVw+1DtZ4R70siKcLp8hfI6Aiu3NK/H+CHnC6/L4h2V/18wfqZ
dTnGKH5JSuBSTk3WiF5jmnMxy3lsRQ5qsMaxLIJYfkWrQQG0vU6Hxbq0f0wNZMZrOUpy7+puNL6X
TzTOpA5/arslFOUglpyliRz15A8g3uQ4KE3Zc2/QhAi/YYgd9fgYGgbb9OUPlk1TaooCqUG69oiT
oeB8z6Wq3YWqugxUXhmMQU1CaOjObQImCuBbWnltmjBHUld0kFxc7IZjuWyEFHYICwdX3HcuIMP6
XFbz+dXid9+S8qw2rfMqgFDt8Kl/qc6suf4U6K9hTZ8Qc+svZU6/r16E+aK2kWZ8zUkriUu58eS+
npvLKGOs4ilDSTtDmHrqmsI2QjfUORfUHDl4NrDtAZyhoDDUFXXHNiMYD3wgPrmAI9Xzmzy09Apv
7BB4HjuvFxSpTATOU15EyXzFdXWssoxh4ue9Lsme+bAg++KgkpuQMXsOGLn/acYoszMhVqpt6wQv
6w4kMsmkntPhmpUdEBw61E4Vv+vVSh37pkl6XGPfgdC9U5nT2qJXfIPZsS9e7KkgasS7yDA5z2NK
k9FCGXZi/mRiwJX1Kjx51+lwTynO/x9vG9SxPTzZLiLmmc7xcSuwlvPbCSYsVwKh2h5fsrbY385j
rBiDsayqcNXaQ3fn5f4/kMZEvNND0PX15ykd5Kvc1jJlaI7++J990dlzsSvVJZTKGdkglxYL5fbo
00yfYoYNs3oQtTYcHMXlYH3fgo/BaBrQgBPyS8E4l+e8NHVQ4EKJJYHLLo0PsUTN2bHx9lbgzrcX
Q5zimfdYZf6pP0XyYRLF0mQUfRH23DN/LmJ5KFfXP3LkhOC59Qpb1cOsfRPHzb8dDQtfVPKQz5Wc
k5nZ7BiOmMQK7xoFh5+Hoc6aJLccGKj4/mzBCRNQPAPTGFvxMdbVcJ0na+GNDQLEGOen1Jw17xOP
Uk+lmmOoHCGvWAF4AWrhibkfMcWiX39sSTJCFi1sgbSnCsMCLii9GyFQjGZWQnl4H/qGJ3/3nNmQ
so28FPzX1+wwOFYGIlJCIiSqa69qDdu0E2ayX6Q2uHskY10z8OcCrfkuCiXtddyCbGUfzAqJUOdV
glvPItCpQntdoQDTtr97XxAH15pQ+CvIFnCBBzUTQ1yAa3mm/etG0ppRzzJF/GJ453v3QCgx38hM
PD6yIULIBtG9KUsi3i2pAflrIIDbWnON7pR5a+hPBDRePOuYKmjlvjmS8Xi63iwir5c3DVXo66BA
csH22SJZgCKYW4k9+PnIEF19otgg18v5VdCKWHmKTR1P8ftCMprdm+a9zRYeMUOPG97JWgVruOyx
WbzwE+nEXfH0BjllW7Bq/9MDQQAYymd7ZAqY8ZPkKoxEM46Nh2ov2g4MFpIVL1WOraJFZrnJgkUV
2S0EROfDSDBXEyyq6oS4W7uVZl9rJI5DcT+qFAyUoBhD6fKva+p7ubtDXWaAGtLJdHBtX+kWFwA4
83oxGs3tFxT9qsEfv1PBuUQO87aaUlMWm7jAEZlD/kswAf9cgYhdK/VYXrzNW813BkhsfWfHjIBR
2R5H2wfONfR9HDDl3qOpsLV59cLWMmA/ziHQeF4P0tN2hsmcvaa9QyiTA5aC8DFaF3JFKh5w8jXU
3bGq0hDhIBlT5jDxU9o4Z86a2r0vQAGrhz44/+lCcybntR0XCwSUvvPpyoWw4PY3tlZZr0rZXD8g
H8PrvXbb/h/XG7X43rFC5Dd3oxdpo1J+V/BIsnwrbBsYK22axNe3bchyL3nQQU3R2zHR1r3//yNQ
M+H7+V3nMB2OGNsAnJplC1ph0sd9HBZFb1T26igfxrqD8yMYeT37tzSHyP2RpCFjIrxmEgojyvAU
ki1/mIAr77/YOvL+bHjbpJMxP2p9u9WP4+dQtMiUxjLFCVqjM5XAJMW5EVy5qKT0JCnCrtWWlSot
80L1r4IJ0buY77NSljnMyj4LUJz8c0T/NMSC9Z6UW1iCaxwF4FEd8vXe4winUUtiAgC9HoPYGf1M
tqRbQ2kB+bbgFLhVZVIMGO2LQt3BYnMaOy74gPDnBNa1NrDTmu39nVfZUjVE8tWYlS40H9+GqksJ
3hbxyEPN9XpF8eTdfoTtl4b7DIe2qwQceU1nI6/ngaw/iPhTtN++mieK8G4n9N9U9oUKyCli5B3D
FaODok+hskHQiaKB3SOuvnINFnxJmIALrQU/v04oFBoqY21RylH+vjpD3YU3kL3Zu0HNOrYIVqWV
xJ4fOM88HtDsEzyhk9OQ40Tx900zlS0m4uh9AjpG+DrVoy3h+e0Ey0M2emElSJ9d4FBi5KTWW7dJ
gS76kMXsdW7Kwm1PGTMzdbc55W5mHehMIPLEVKbCkHKJ5fZ3WURRMrUDGVMeeuhB38C9dLdAaIPQ
VGVCpBA2ANGndgyoWfXNLhV4UEZ1NQr4uHwuGPqddBM4xK/XugvxfrSEps0SlsX0fUoLy++SmCzL
VRAE5I9mPWeDeFq7i9y1UoJXm0uqo0wxFm8q4a1iS7hD46slZZRMFDF2uUf6Wy6mE7VpnX5ABEFB
zF1K3vLNPMrj4Bs1IbIcT/K/CeeItAl2djXq0x7YKo75FTM+70Kznw20UwX4jc8ye+xEFdWG7sHd
CScsbkCwOsE2FiFBZrJzvTlG2kdkYH/RHtRQRuN6niYa28DsQTCyUkO3SV0ae/khASWXqn9o0Gb1
lM2RadW4uKu7cD0E7HIx6NKpR5cexBhGZritTENY4lIHoszF/ApqaxgdcQHMx0AERQXyJ08NWkiV
8iYhjG0ORjcswnESzDvDqgcxq3DQbIP4SbrCuSkDO5qqLqCha42stDVdP6TD0CfCo+qJE0IQ6uMN
2Wzfal8xvzJhbSBbCgtN6364YIQZZSpKrsilY8TwBaQglfVgD3zd8A6BLuap5A1BQuPhA5C2kdd/
k4aW8dWu02cNQrxx77m8eeAR8IQeYj6g9x0U1Zb5e20EMsIXRKpX4q813ojJHeEoLhLK0Odqf1dT
ofsxw6aEgWaCZgfET1xCCdTdE/mRgLpPZ+2IjPW8bg/EdKGLBU4wE0hE1W9c8gFUtMudOU6Gwqhe
BwNYF9AK0hOhsgUYgyaV1q4uCJGX7DCCLyaoo7Vzr4M+cYnBwHmI/mn4iS3ObvhZGTkm9JKpXosk
+vAxjj/uU097uYf4TjzVqdvjQ8pn0HS4iIqbV5z61UNpC/ygrYHMecojD75zu7bVhNozHh6sGR1j
snxyzLNy1Jj6gf7ZK+qWMVct7y275DPDhosXW8h7W8Xt/CDVA2c1+Sens2bZU6UahVgolqUZb2kp
N1dPzjAaa7xYf627+MAMtYi9FUJp3e9hr9YOhh+8WQRv/zFbmGDS+GUxjVXbDBcSlg3OyUqQbkZ1
KD9x6AHbz5YcLrL7hiwyB7dfn5cbAKMx9OLFbimS0kFRYHsfASv/v6ZR3qPIfs26S+MtMrI1HUdO
4IT2+/f19dzlHlVhW0Wl49WYwnG5G1yZhImW7V2Yc/EkXmtqlKbJMvqGR4rmKiitGYAihnssG0LS
ztKzf9XXUAWjHxhTDfsqUHUcS/EtLmQkq+vlNCz+R90KjmEXItLYeyghoi1Sr+ybIjw8DKLKolt9
NBMfPepveNP5JecNwIZ/SUSLBP6MwqMnJrkm3sgjQi9tDN+if158mKE0FlH9hVmoWZ754JBJq3Cd
IKYNDeg3nHrwbHkyY5LAzJMN4RxDccjPDbZcXFtjVUgNQ9xdi8NUX5XV+uwVDxqWD19POK9NCdg+
+6RiQAHMnYN6K92HusmlQQSGxSrSK47FvQhE1BTFZtD3OEgbkToIISyB1Q9Aj26gAi1KhYGj9wpn
hfaYMfF6iqnnc6VYYkRHwXyqeN2IRoQmzasaTQS/wyHMxepzApuRRq+6Dqj9Q20Uq5BUxB8wCdwV
2LP9lJdXkduUmFdvQyWYYjktoodFBbtSPfKx9lEutEMEHotPHXyubKk6pQdAak9fRosSrY5e3i/3
Nk7fZypfov7hKbIveq4dcCN3lE4RxaD23bEbxNts+eqGLMosB3PvWYMcxI8mVxOFl0snoa25wYoW
VotbBpOTMZTn8obrmK+bfLxZFpsQKhBT/hFMZF8cpgmEyB7Ds3v08pFafSQjc3ZduqupInASLFXT
2DdSbQIbkjwKneyBR0YLBhhUsjBcGmqvsT5OPXT/Mvryod5ZReepVTiGjqCNDdtzK6b/j2r880mc
QS9M7QAUwsijawvIDRMeJJqE1BDI13dd1POFwiWi/iFPfV0Z/70rG5+sT28MYuFXwDMiWkzdHVBY
ohSrd0pVV17hIaiEZ/YMXORhn0lgj0cUIPK1vh7qwLG8Kp8u31fzHEX5ZNdHVinm4XozLbUDR4T/
l5B7Cu91SimM41jqGLuxxPS4+T7sIsmJthikoSWliml7s0wPrND88iN2bLetpKaKQqRrnvNFEWos
aqgWYKXQXfAp9woWkHg5srCQzUaeUomeyIC41/Z5KdfuQbGqN7smw4y9ftFEl84i+F2qPXqrCCfW
MGcnf8R13hpbVwedH4atnXFtitfv2h758+qRIAR63aum4zcxXic4V4WM1Mzds5uN1LoXc+l1v+F9
fOLDnrjLuFASsslitvG4vCoah9FdGNUTVUXaWkljbuPE82g7lpO/4ptpjRJvkx6Z2JtV3z2RJGZg
tf7ekLdVDRMCedTb4h8NPYq2LnmP8PWbPnZQjdoGQeVv2BdQD0B0/OHYFi2vbn7b98l6q0oyQcxc
XcB15NZUfdAKVv6IopKsFHsQ4h8v6OCWf2V3qeJKhsgaq0bLc57RbcRZPJnNOCX/eCCnWnT6Wn3P
yh4xJDdqEn2gviuPAD3m+f8TMf7i1gp/c1VgRthSUnMf8NQbB6wnPswi4x8QG1RihyFy2aK9ZsyA
PhuQQ/mtcEfqSVOnQ8nXXsuR3tLKlclLfuK3rmIpdMVfdwElCv7oGCVtx2Yg4ovM0eng57g97/b8
bayOyrMNbg5dEl4G/mmZDjbQbqZ2UstzxE6nXLO4sXCW/pVZWgjj+0Na/QXmxo4Im8LpxNevOQN/
AcIga4yjVOole4SDliKa1bX7WeVvKRi1KLukGezKYqT07ve16BaQZdYP4pdQl7SzSvAWkWvG64Qr
XxDu0XURBV7FaUJXk+gYPFGdkfwfDEzLQIe1dgDsXK1ROR8KY5DI05itZg0+WWLw0zvkCu+gADAe
RowbQ+HCPnnyIOzIXvyZSORRQ3k25x65NVAoD0SnKK7iNIIF4QtZi5NI52XVVLXkx1qBp2HJXHFQ
wkdIHzubw06dsg/tmz2mZ3pdZ7/bEgocPQJajI4HvZYk2PfF1Mpj9adlV+TjJEFG72zak4CObsiR
9C0Bg/6a4i4gtKVVU9JmL1D9rFDXDhANHdT47S88U7lpGJLitdbppFLeqZoNQs3fJZexOHk2vRM1
v2lHJwKZlbheBY//Vy0QXpYBiwwMMWT88awoiWKoP45/eXCpTdPMx8OeJ4WbYNNjctnVfl4Vcjva
vvsnAj+5Mw/Ad3bfxf6eH3QTAhtzo7eFwcEz3BzFO3NUpT1/nHhbLaweaTjnOPbSmTH6GLiGOZq4
TD1lPSIymRHjnaK26jB/CuJ7z3Yl7gKUXdrptpnC7gjbaNnOXP/GJuoMC0QX8MsSqsM0VvfsS8LK
v7Rz6H7ysKjaY79XZ4sLsg152EbE5T/CilziIR2oTDUZitV4b6b7gPVyb6tITx5fVUN0zCJGa4sQ
lpAIWwEzF3DqTWPfwIk9ZMWE0+lWFw/UAd4JikQBQSzYR2mKbUj5JCvKJS/qc4l1fzXV1JLvp9wH
gfw3gIvLLW10KKfpH2uxsw0BX6zKPFSxyIr6lTaNvxpfSLKgqqpHa9p72lZTnuAYIZPeedoryTRK
MoEgy4vZNi/6NkbL4UQ0836e9H298P5kILXZgSUnHSJi1KNFsrMLyyAL3SqymdxMMnrOb1HTGcZK
zZaiQfnTj046S8NXZH/FWJEEHPr+bCZig17s7+mCSgCdSLPYxw469419HYGNUVVK9CNuAnseJAVM
JW62NX4drNqkPxII4DWM5OldvjPKIqQUrZilPKsU+OUeU1D7MxwYGFTfK2mfTuHVlRlT88N/VStD
TF+52jbNIJ7hHCUqDlaUEKSBeAOVHAJYpFiTl4Rd0jK/+UDqq6ifb08+m/Hlhf6rL9MiQ8ikomv8
DTzOS3f0SG3XIhUExjszclBcQgQDu4Pm/IbAKvqAhSKkXgyHA5rPevetWZHl5GdbPPRR66V69Jr5
DDqhvY8ifTrQ+yNKn+kVOmNnlTVgUn2VIkrZaRUiOPl0CFa/C6L272pohHzKb9zBRpI3xjuyVDNb
bnO2xv20W5qx3zh0Tqp24ky5y33Dy+GYYFFK+h5cuKq69KV/BXmSEJbqGrz6Gu2uGU0/jakZmD+b
uOME8PIdB+3bvZqxtAit5UHMccyLVdufkPVC79I/4/jOjqkysRqWeAoXsxRV82uzNLDemIRw9CS1
9CSBt3V+mfAE/KoY8tgNvuVAbU8dLeLeO4ydVNie+IRe+JZTP3t5/S504oNhqzb49Fn628UCcdVd
30U7S3c/O2IP5vW5xJ4Gc+jgI6EN6uXghwjEMCupXOTbPjTmyBqbm4G88EJrJdn9wI0rQ5Rv+5+w
9ciYY+OZcPT/EWEPaOnDTCYatXGQG2Zs+A3ua2oDO9f341vR6iTnyiJDdKXwy7a4Xf4raNzxygYi
Z67OH6dsr2EEs8w1hp2Wp2f1JGPG7K+QfpniAG0JMzewcjxJrcIDnJ63fMc375j6r5ZFAn/Z3JyR
UqKtyGhk3hdLj/MuV+S4ihXIG0+wS733PBtsTjBh3k6DVWKAiPE/InJj08sntSZFdQp85DJ4gW/i
wNpUTW5iB3nZvjfFEqlTPwGpc88TYrWwa51e/SLHOW4zU2KK3VxhuFSZutEBC6tILAEcpMYnAvoA
wx3T1JH33PYf6YvrfKu0lWSSPi41qcJ2sJpEjr5ADMIzst4aIknkLXfeH4E0L061kQ/ULvEnUMYJ
z2p+sC9L7sDmoFVN8GonVkeFRFtQjkWxl6h2ZbjeVH5VO2rxSJRdOgafhWW/msM2XzSx0NOsQx0S
Ye5dUTkkqHAp7Xku/u5RonVWio3j03n35q1tc66vngCITiRNOMwAdDNcYwX4r3/yXkkEEWR6OctA
PQsgCeJMUCDJgnYTWh7yprAV3v/4d2d789uicqJCXMzvYDOMuEjf6FsScYVul/oacRfXRxlzn1g9
Su0R0xJ5RlvOlrLANfNJ6M4bnqv9U6qnqyO0oomktwlLhNQKW0qao0JUc4j8CGl9KnWz0eSkTXnj
NroSHLSwz+7XIh4CGnOP+/jYx3wyAhtxit5D3Q+ZFSk75puCo3fgG8R6aVbrmcp2hTScu4TwYbR6
ioq4iVqqIJmI6lXVdDcwTU82riq/iiEvlMlSC6Os+x+v3AzRnxzs8mxq0i7WTFSu6pR7rx/g4/fQ
4HJ7rpbA8IgZjyVPjL9zqVvMfgD2q/2w9Y+flIfv4d/3EvBG8jqxxuOU0IHSHNM1MpAMLrPr4Q5n
BDY9snaUcFKV45YY2PqS2ThU/rhwlP7mAF8WRAJ+9U3Tapt2Kj1YZDdp1gdz2fqP13vfRxyCgsGD
tFut3aMIrH8Y9tdzGbqm/M9FNLEPsCnwJNXdRxNdU7xJ7qoYWqgU2zfYlQ70LBESisjUqkQ8oWpp
AX/I7W2Gsxibgj+dlhI7Tojx9g152UGETyoS4vHSDzViLYGi41ZpsMwA3e6QzKpbUPzOHD355R9m
XginaR87MeWKi70mTbS3gY5k3a8F966KTe3ZouqnvoD8XhueffUZ0592fG6oLQIimJiNJ9fTff1M
K8HMdgS7Qu7FPwednnjoJxXPBv60r8gBH/3QVnLCnTkaPqK0ER3Lla89/kpNt0Nt2Yjw4p5PiAaY
zod1XYwn0sSiwKfZLe7/cCC7E/1suB2QcFnS2AoJXO357Kj/InYjLx+0AIxF8A7AyMkzqw8f95x4
BHlZMXT4pg5q1ZYmWbaouXPZ3y2oD3yrCDHCGsPbzK10S21pQDbPGJMTgQasK4Ef9jj6BAeo0ZWh
RUssJdHLLe30bil/6sMxwRC6yoKx+4KTS3mXxXVnQsPDVLVY1MP4WWj+2YQiqoRFAALGnulNb/LN
p5XxoByhGd1xoVFGNyAtGDhwW4sJnIw3CnlwB4Ef6DmaDC/1SIjJ5oWKXtTNr3etfzk0PFWNDC4E
rAvu70RTzhxpGh1DS6jgZ1dP0xFvJLQZbYbEiVvb+3cf6VxIk5uK4BHMuQNuASNTu97tAOZnfmUP
OrJF/+nRjvXIKnWyDQjm6cASieIzZ+RXDMFACpPN76AfaT+JOPobBozxS8QJz2TflaoHyVv1SFG+
5UsV8/nok3R+iJN6YYQ7fRwZwire+3yT7ZhMSTxF0vpakf0cDtmZfSOB4VRpBlPN/X1f/tWM+9gQ
E6bWYnTJfx/bkjQCGdrpikT3d7bRRfrM3Xq+Qz8lXHCFVO+XkSOqa7eZAiEJt+50Kv3u8r63Dfmm
ZPNrTZhzEWJB+w2taSj62LCBmUpn0+IpYIf3kkCmlxAeEbFGlPVRmvsV9bYKaGE+ZEtwiIX7XBle
5OB9+pUVrQi+hWkXdi+JoZGZWnr5FTNu8xyEsEfNGNWAMOq7gK7CciHs1dku6SWpUzb5h8eyofQM
xHt3YRvvi5b0HkvvW5PEKFtqUnZdMWXYi3vR5G22tnOpWmKVC1EO2rALkgpXLRqTB93gw9NXRvwo
Iec4CAJYK16vG1XztMW6Ac1xs4gcMuQGUZuctcOl9FDFfjger9z2nF/N1opjejG4jbZmiq1TelyC
sPQk3EPKFcmNl/5RcTwd2+0HWcbipKXt/x0WArwi3IGFDTnEA6SSC3Jo2/ipMlByhx6rmdb+wWh3
vvRWqSMaF2IUpUZ7jihOcIlxzu2fAEhuQuXiUrNgWISRla3nScUurOa4mwACoTwyP/kPD459G9WO
en0izpuYMrWYna58fZZ1j3ZlwASgWAzhuvuOIk0x5chOmjwyeUa0uX0qt49MkBe709QH6pW7Lzcq
qXct7LO+Ps5LtQJGiTmDG6aDWL+X63Tq36jjvkY/I3NgOXJdPjAApqLCZqJ4u/6E8gntq5pF+ys8
zocOOahwIauMFFmMjPAxYA3Vbk9v3B95UmNuBpybknKOTJXUBv0HMymZ6UwQ9fPwKcozjw3XFhUa
dSrdGUKAmA/bCpoG9ika/c9P1ZrL46Ly2/N536JjZUyhp22lGmCEQ2zSXw+5Lw+fSC1KhcTFPQhm
qdxBNg6iB+6CR3n0KtqQL/AL9CseOKwpdMCVZR3KkKxKcXlefQs/LqZJYUAP14tl7VPpf1VXDjRC
TyN+Jkxi80JKgE7q2F3XoXlkF5mRa6syPZuMv/cI/f9KXmkZscN8aZngzYU3NawbBn3sHEsJ84AR
GeX4XQ/lPq3EeBqMcopqe0P4+dh4PFvtWdJXfJByAlwEv9vxPcPSIT1GEiJNqo/pBML8Dok6lB51
dxwdH6YDz4EskVib2akyEIOd33c84Itavu7V0JjUhXi+7VjlOmFIp6jRHMlOUEA+CUruGu0jZ3ch
0qjc6qD0VCgts3HBia1HrvG8aC90IgD0xoUuBZzQbgKNxS31vcvyj17UXwP5r5/QD3DBfpjcmt5V
kCQoXrePEq7AGKCzOf0A/PfZNsa41uf9/4Q2TwdDUEHlSR9+bpXgyhVtomF03WWlrMAjWTm2ymuJ
lZrqF1qBjBL8jPeWNWzt/nsMaXL+x9l7zje3SI31K82ASkX03gSDkSX9CcGya8V5efvJCC0x+0a9
8uBnEexUpQYuBeVW0JJfngaimqJs1tCZ
`protect end_protected
