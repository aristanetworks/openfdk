--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
ELDS7gcYiKJ9ZI4w3lOC0X8NHwC41LqknMoKj+mC5M8ss15Wg/ug3+x/BADOxlFICQWNlGCBy+P8
YGwqdWN+740sBXUlq8lIMqaiTQ1IvD+VdWtdn3ukKRhqv+iUUlCI9ySrHatGowMjKSTDvsFkUba1
h04ub+vigkYeXUUPKR0ZttQszSxJRgfU4V+TaFd02T07r35azj6OmHr1HSEJ7LSYyIshN7dGLXNo
lHQESqE2eP7wuSWe2LVsy2QtkPdS+YsfYQlHCv/nHzajjM/egTlSeIr96Sny8PdG68sV4vzuMTFL
rtb50kDncberqe6UGPBi//ErOX0FdnMPAgNO/A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="f/zIb+WB2zSb3O1HJM5sFEh6RuM1UWO8+xDBnSjmT7I="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
CINpgblLUGKEfBPdrnvMV2NFWq2aMKMt+0cR0eYl42K8j3osOfTePGVQbXub22H7UdzMp1IZlwmx
Cwfz2RCbv2QmjU46MorF5tsRcN7HQtZ43t6Z3laeE4uM3Skq0z7cBlnsxnJyrf0Tap1m0Mkr5pRA
mLvvq3VtTlWe2CHCS9shAnbcRCIXNbaZXTJ0CDXm4AjuDGp1Y0nUuk063LASP8T2TzBqCzUajtXu
bR1jDa8Ag3cdXooHWfMvKJI175Ig3NTQSxVXWfe5ifKospCdGcxbT3dp56ms0YVI6Cojz4yvMOK3
XXIhydkWqiBC/8mt3JmMmtCnpgmUeOoiME2SUg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="oINpJ/9KOgOD6eDyUhgcDPFgNjc9Lm4YFCV6ELdVLcE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2544)
`protect data_block
8QMbAi5y8K7cgFmIexoJNjYOj70jmi9UearpjJcRni+XZGOYe1XUqJ2N7irer/4ZSOGfDOeY+xvI
uAuFryx8LTyMN7/Y/Q6AGkdhxYjftDm4bXNlT/dYBHBuh6A61Maze/28dEt0QH3qwtzm4q+cg3tq
+Eg60fT8s752uh+YeUCAwHHyata6S4dGAWDzYkEduVMICgwKWF8o0jYTp3PM+RNUmJ7UJ6auBiFQ
dXGBlyaZcwB2zppaLeYbNmJgZcJY532fy1j/tu0EBZuNf6Obui+S1NwVuXVGlAYPP96hNMdFnKMK
uXaGc5Agl51oZSUjV9h7Eh1mvpW8C/0dlb1EPkZzNoLJ5A9peFZmBLRcyVBjvQNnzR6WnDB8hMsp
Nae7pUuD/BFrwJH2rEg2wo/HmwL+msgiU/5HsnZVCS6IBTV2R423qe7nvNgxO0pzcosEzELT2AMe
IWNLuScw/dnYUyKtdrLKdn42z+ukEeizVgYa7l2H4/mUeeJn4WagasZJ8wMkbKorEWbFQRpbKuq7
TWrAe/2HTJ4KMar5HBZlLhnH0KPJdHbx/fWoWR5SJWBc4mbd2DXW7z8cowU5UhCYHiFXu65NVl7q
E/OSvl2oxxvzoUSKLhD7b0icUeDCFexCVpNqo0f4LUZdLe+wzBaCEmtapii7u+lPEAIeH6YhYnxn
bs5vJlHsa7yHYXAz45Qb1KxNDOjCoNIVii8CNkM0Zp0DIcVhCA4s15mFGFghtsx5lyMR8X2rRSy/
raIJIOQ4jo9ARuFlxGEXUc5+pzNcaHU0iPn/VS04xnRacUdr4MqTeCMjDSwRTFjGzggBFM+9qaf4
V+P9QvxznjKCXCem0EhHxGMEQunxSdQ78+Gqob/XUkFZ2LbN5v0iS4Oblw1CfctbZbqSD/kyIY0v
LJoV7YA5mPSmH5IJ5R0QJf0IhFOQkqzfX45cyxGnr2EvPWayKPrpGfuCKpMM5Xt4mfhtr7Ualp50
cP1cVch6zYAzGUl5TNMq13ASh2reA1XMhcIeN5+IvqtmR+QwkT/zvTHskp9V2sSQ3X+HriYLH/ZM
W4/5Q8goQ8zf2UkUHcW9u2CibNvTlsbCJIBbwOOcsk6NawCja6hltQn4SFLh1KSYfg76KjyOPWjh
g5d77VpC8RZA8Xi6MStff3sSeVpSbHUovgckFC0K+KHWjfMF5HYHwlGscl2CYklhc/7K/qsVHPQh
O7fIG0lZo4yl8zxNEEMM/kfMukPLgmJUqOiKGgwM4qEgqnOym0BpIgFjhvjY5A9Ociz198jRKyQA
lDuSiegkb2uQTtaYi0d+D1qRa9MFM7q2fV9udA/f6TtzuB9Bw7EGNJHBmPL2xizOllzpJfeXCWou
E7kHoJcuAu3bE13B2OhPnIZtbLhg/vJNsKujw+mNzFtoHt+Ue+sdkOQzWL4GMlqzBCjLFigGekJG
co0MtO2a/qJRjT9ff6jPIb/N0Evu84RNYLmTDodfpfIMgM3YTa+l3ifn1YyVkbM3/9J48VHmM1af
I6QhmLZUte82lifipmbOtZt1vuuX3a0/7EukQIyGmNcoaJwQNP5nUvOKdGfQIuocXMowzIH04KqP
BM0K6QiVLR4Zl5wvXFVvRidsfWul9JLvw6+g7e0E7Xk+pzmvuLABz3WurjvKHKk8KQZCL+8wqX9O
0BGhNeuqs4JeFU+OOoZtTk1DjJmLaKYTSRoXHwoGiSMkhrGiFE1GgfSb8R0B4parcFJRe6wyCpS1
/IdhfFkTyEpRzvqrTO1CN9VVW5kW5AXYOBbaeamCIhPPviOy3L7JH11BGbk0K4Z8j9H2BxKeQuhw
UOdeugqNoeRcwaw/ssMEFqOiVRqPre3qJROdQOcK+OqcEbHAskuo5U3RtbTEn6Y7CChv/DY4oqwo
FqhJ0sZNLAO9lZs0UD7oKpVWxLOxUO+ePg2Rkcn3jkkirRzHbqOXuwP/QDx+RV6C2hoZhWDdw8EJ
TKnwNuk3mD+wq+RuXXo6aPm4cHRzcTsgyqoeocWuiHzl0IVPYLjAgmow7bgaaPoMYRYTlCH8s+lK
pAcFNLp0fe+dzpqaiqNj0rmJrzWJgDMaZKnG7Mg9K2oluxVZBGCLxVD/cb+/FdUkmGOAEL+pgGls
A6ms3Kug29Ru4qBcrnH9WqZdkA6qpw0+x/ojrnogxSqxtfsdMoU8bZBMcIlb2DuT2bZl8vNwi3+m
UEJdAAB0FMfg+XqBerA3++KK+fb5/cRzXh3OADfRfrTXlBpu9UnxLP+Aes0x7e1PZj4NMbQFkScs
06awHHGf0Tpj9VbK+UqhC30flXm0HzB+TsjeQi33Qy7NExGNIBOeq8VcrvSzU36ewQUUGpGsq18j
eRp57OxxzHJpufWEsaw+B4UPdFFoTBj1qq8Vn74f0hCE3YEc+Rkfs+MgopVMF/H8JxlkBj4p3zIO
SqFjZA+StcOvdvdpbAXTQTE+QSFfEIrWWNi/p9iCVUggoZ+VqwPvhGNtsA+ZSJL1+meGHax1T/Ym
Et3gC6YvA0crMhekmp7qZuXpkNAa+z9cKM8jztBbe7aVJO2WPnk6EJlXdwOh5MfuNJ9brjuy0q3a
aObLC5oWW2fb+iYEUdEUS8mxrz2L2tmbo5Jp+tDGSHm6a9G8n+qCz8SoPMisXNjJfjyj5HMztQMn
NQYDciupWhcwV5EBRvGsJMXSj+0IjBasfaOxWWrWkUmJ/kNnIJ/rIcRZieKo/1WDndBX3al7GaVh
qtfVZQmrX2Y35AXUKMJpl4RuGvihI5OJ0dMK2xQkDtdGngR5YruEBvtTvyiLnaLkDGOTLri/hCEr
Rbwp+Q0GhP6OfZfyxMG3Mz3l70+Y6UX7OFepeWn018dTMpgqRJwNEVj4ipFok/QENALG+mXJh6cT
Lz/BNgevrB/lX8kzTscgsSg/Z6TcYvezLNwUNhci/fn7SeLtflg1ifZUx3jQVQAVnojw6mII9EfC
mx1pU8nl02Cu6l1Ln0RHTV4QqjoW24NUdwH9x5crwTwvocHhR4+HFdEHINUIJ4DPXnLcc99iqDnS
gai8PF+lLK43JzSYEWhxOzv8CIYryTw8s6SGQF18HAjtZUydSGcj/Pkqa97J5VkgemLZ2NkxMwPT
fYIiHbgFdszv98lRz1psO929z7Mg+whupQyin/S9c334966REHxIdwH93PHO5ypE7d/ooy7sD4u/
bIvtvnEAWTOg6ThpSz1W+M6gtFYuA4mRZp5zJduUO346RO1pW2XJbGqhcz0lzEisPh+Y5o5CFKwt
fDA5isaFMfGubrbi9GicLVjd4iQ1Q8HHEBNJ4Yl0MfcPYIK62Pm1YV8kRUevKJ95g65M+7xwTGi8
0a+r4LOCEoSN1MqGwenH0dcywQ9U6/LcOlB5aQsXuPX1ZYfJ
`protect end_protected
