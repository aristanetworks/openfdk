--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
JAqsnBzK9SgBB2aQsnQzS4EGMcL91Xv4ZNbJIDnqrMeN3zbhlhkiwhS/JQe9vZSD/elgqpH80Ayy
Ikv2IkzSTGVuE609VQbe3VTrTBO+9OboCIv+np7wQwjd4nphk7Ilwi3mHOHV/ll/InldOZ9erAaD
ek78qjT0mU9jatnf6BgcS0ZmztZE1PzbI1hutENl+UVSzb4MLBofd1ZlTQRgqquo2CZylC+eS4Ic
dH3C/HcROEjqEiNFi31EZrmGHab9xRu2KDuP083n/7xNE9mWV14o8CG81b3FOETqZiQYBeNg0xxR
ZrYKO7JMR8QqeMSyPP+hbpFL0OG5Kss2CCf8tg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="7a/YXDUafrclEWBXpo+ulkCzXirepEWhi4c+iqCS5sg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
Q7/RwI2HDHdK3VyGmiXphYiwMP1vdiNOEc2pkghnlrL/C2Wgo4FEzIdYv5Zq8KpjS8ZS2Ioxn6LJ
mcGjmiI/wK9AfRFd2Gthmmp1Qx9H9XUuCdGhanUq9e1GJ2lq9rQI27NQoom+Xf1DwajutxYRd+tO
RsgTsdGX+gVWDh8MV5Gf39n+r6ctox8/NIhvNaLzyWtwkh2NAZGjMRDzZNhkjPFl4vI+CA0AZqeJ
x7x72xr/arti+uWNrWaItTffdNVWP7feeKOBzgQUqpuhcWEHsUe9K6UqtLtPJr2dAmRSeik/EgLP
uPf5hWryI3TLEtkWhp5Z3IdS/keZYVgVD85VHw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="z5s9GmXSONKk0EZQLwpiHXwFouLFRTwrk7Lj+0FsTJQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4368)
`protect data_block
k3qWE/Bb/uazBWQoFDGP1PERliuJFAtHIXnTMUmjYhFyFepz76tS9TKCdr7OkYLw10ctn3oBHIS8
kShpD0m7pzC7cFwO0RgcrkGxuwRZMROR8XwbFlhIq+porZ/6vFeTJGodWWD1gpKZUa3h4sgJ66SD
3DiDECe+epMLFVcOYO8sJMSDtpuOfjVeytwSOF7ea+r7MIWZJWe1ncZsS9iCFxVfurLSyZSIsQ3I
DfPPS+3hCL7PkYmD1VXIaYGnpIfhqIMFxqScIacQQc+MAwevc13yMruYkZAwULeYEHEF4jataYBL
s7JGczsoXqTub9THxD5OAasmK0JtXhc6vBdqK/R5xTEYfwPUETbxDAFrHVB0OkOIEMHi8zHNTERx
5biVVk23d6Ui2rYwsVG6xUTNYuRUoihZFH1KO5JASquirH8yPKOl5L9LUaHnvaiiebzpKam2yvk0
/4XjWN6K/D+DHQ+m3XUfld6CM6Uf94455dKsiJUa6NltG88/MEu1y2upSf2XAmQfTxYVeRSonz4b
vH7WCzgbLrUtL2hUkWmh7ew/WIdCsOoKcJr6qpTpTB1cRKIbYmsY9ye7w9IwQLRqUNfUK1bd98mG
VwfZam5bzt2jWr0dLGCAMp17OPA7bD9ldi1AD4a5aJnt5R7zKc+VtzqErVDN3jeOPrm1+MJIyqHl
MdTQVBtERKSfqUXAeE7TDzAR3VQGdaU8Yc2f3nfc2yUq6Yd7govUqv8evSYUp00AC+5pagG0N95e
bDmeVXYzUfKUOE52CcinIYGhcM+8wftaaERVjn1AE6oCbaBtXzzvSXht7KWsnwQQorBHBvqrc9vM
aZoreeI9H6t+ne8wDbS1SfjuaTxIuJNokTaXjf6Ei+lWtSTY1K65L1R71DbJ3qztSUvYTL3wePiS
eYycQU50+KbAwn6YqnLXLaUJ8wPdPZM+YJe2xh24K3S0pyCbISMYjPRlKiN1CjgaFEudS4O3XoA+
XAV4M89WkHgPvfAG8IyLuIy2fW9zoxUJ1q5cGVmEtl+FzaaFHFu8yTVCRW9SalaNH/BzcPW47XDA
7QLMyWBLS6dYqjSRNre7nlmTQFJQoc5KWm6PVMOm6Cy4bIsFs/eNzrTSFoHOsH2y7s0w4RzFKPU/
VHcauHY+9qD2lbAfgz9F7Qu0a/Ko76RA8xzn0ZEw7i2vxyDLn02vqvLE/P+yn5pAZSynXFfm3Sz3
X+WJPryDJxkXur1cffCf5LqgrVgLCtkhGUcZ+glSeRlxrBqIw63Fv5niRsFtbUoWX+t/pCw4UnPC
SBH+UwY9YAbMxgdnMELX5FqbgjZ1pzvO23tkoSVy/4d2wKX6/mNzVFLkqOeUbFZN3u0OXaAxxTuE
C4Smdq3ad5o7kMdhf4RRvpAIeX7lGV+y3bN9oqP6KOJgbA5mA3cT/a5HicKhj0v4v6WjdTjkNqMG
pDUENouNHNK7vgA7D/EJNSdowYl47+KemyhNeBrD1xsqwKDVQL7TXobppERYTTJKYhWNbX8VlaCW
0mTZliplmJoJwiYRjM7vWgYcurROPgRp4MHBQyYCHfuNRknv4FWa923zRo6XjEP6fgwoq4k1Ln4K
s01PMbsY0g0YnqA7WpUngpKM3XJJzYNy5xzxF6s0v8zyHoxHhumKxP3k4RopJGgzryYZsjGxT8Yj
6hP9TjsbTv79onVk/CVu6v9qHvS8mxeAnnmT/x2izQvcBbA/Swaoyi1y70R1E0xAyQqBnVKd4Ab1
RZn450l5UrY1+U+k1P+E/8Zmr6dqJMNjCnjVzlSPWWU93gnwL8b5Uypb3J0kiYt9BOAZwGm9khs+
SGHA/k9avRZW4cV6ozv7fOMhCFNd+mhSAPC/MTxlIXbAdEjlzBbbUfU1m7qWo8EoSbOdy/HtDBMk
ocs92q6THMZta9RMLKmacqw8nYjJtWorjblTFdNJ3Vpp9CDAzKtjaJuxvjawky7d3KWPRPS+kkqQ
VrDPwkKHm32yPjOkfZQUE94FX41kP07syEoZ0IjKH8+iVh6EuaXdLroU05rn3EBFrDSSGX8G4MpK
WpTrGsXMiL2uBEKiXDJ0hqYatJsUnFpLvPkHmpXMOHsKhE3hU0WGK8Y6gwjXNzUuBmTfedPUxdIv
tZqrZgoCbOFN3XzMQjeiGgVFFO45IodOX8v23XFkn7iBsqWRJ3FcLiihbrmtb/67tPslYdPC3LNm
Xp8GdC4CdPXtA8WHYzX+bmu/XrJ5WCJHcxzdPgKmgmkvvotq1nJ5QEu5jXwcKoLSrQ5+h9KEKvG8
Rj30BMOWNlDSNVtw7OZitek6CMRnDq02odHxHL/h+zWyt/dfb7lQanQ3NVMmr3dfotQCo4W6XiIS
TGycnIPFjotqD2ZmF/9EIoCaAtR9udUc3lLgRUbSoxJI7a1Z1GsMwLvghke65HAdlcV1llKEz5US
JtX4dLhC3KX7ZGRVQrmnUfqbkd52PhuEOoyhSTxFloJwiqoROnXg1DpeMfXYHIWzJk+Zwy6YoamK
U48t8AyYXgUPERz8FKdBzL6bh3Tm230HH5evkkHcP0Fky7pRdUGzhrEBlhxooUuFpyOefiVDhNJ0
a9rduOg259x23R02nJ4Bb7tVSHHSfZryGP2G21ufsB8oKwiwb0cdkYqzkgRJXmLRFajxlDine3iO
IzlyEge9t1BNE2e0xSe0NHZI5qY5Ed4I5YPnN6Bq+oXKsMIf+7Llm+2gCX9SJEIxm9ASbNEiEnl/
V15jRwc0Ks6OntPEkxwpeVT9bouo4dtpxmnIYFmii74niFXSRpsXNYGjcpPkSgjcBD6A6ZabYmRN
2k1eKCdN0hzhPbiKxrGZUK9BC6qVDr8qruQSo2jONFhKU4yziI1aaPzsPJjdVhrFj9LadYglQ8rN
kEFjdGOO2VMQKh1u04aRVKWrUTouH/TmvxZW9Nk5XxGeH4TNl66IZafWsQtD+Xx1JfIu8IiI0D1S
Oqs+vjbAvI+phCFzonWy9/NJvWqhrErfPH1ofLpju8nUmjoRGdTK1+ZId3AF4adQn9x+YVAj+gvR
eGlo+dRBpXLB16ArD92UX6wwVK1pW5rM8+XpCp9O6aFnO3/zAZsoz8d8zN5mD6fKvtSOPPFf82bn
3S26Iyy5aK8Gz+JW+7LL87Ui3fXzw3wSqISHT+cSVBMe9sCgy0WMRKfm/ioqY1jKE/CLx3WQ/4lr
VLjQesYFFqfS12YkmGpnGX6mriVAR0eCbC8huZpKkHEf8b+7RU7PZ9+VI+Mx17ORAiqPffDuaGLP
/kIBzZqHBYUB4BOzf7CqrVst/Rm2i3Jlf/fjfHKn3tAwUxNW23HF8z7HFeyEPamKcXtKZO3hgCQn
NpV9IJH9NvFewMvxs+r7Z/GeDjAVzhvmL57Qn7UKHfJ/8cLoAEWR+FC+xIlF/+4tkbWClvlnVD3f
QPikUcX6JdUf5ZuYqO8ZASYv81AV85CYkwI7RJ3VLJ7KOfwwpGUQYU0UKFgceg0NdUWMYsa3Ia8G
1i9qmsa6fYJPwx+O683+ZMuNaiz23xP3ZtRpnIzNS4HrnL04hrWhAF1j84KL56w8wyR9OQPo1OE9
GEgWoiRpKBt1WhpbOY334UEiR+whJop2Mjd9g0Kvrag+c4oGLdCALHq4jil25FdOc1WwlxXj9Xmx
v2SbMr6LYtHuoBDOa3IRL8Cfb3F4egxgyomhQ8R9Oqi5dBwSi8ux9RDc3bAs+lumnlAkpWLwmMo4
Nn7G3KDvNrYABywv08FNJjp8W1EQiXn6D6WPCnrx9hWV5FK7zBFEUHgpQp17IxrxpyYXaiodW9Gd
peDFKTqb4P90smY6PQoAMKg1kHblXaO5eA34BON+QQETsmEse/WVZAuT9fPCFGELTOZH14kgjsw6
2xoRzB9gAZMmSihRAsWJPKByiSmXu1e4YGTVSG6RTPnQsCoyeWHRLbgT6PbJDy9a99wAyr/Ms089
h3tOCyYzq/FIPWxFLoQE4Q8TtlRK+eKcmSEkgs6S4BR5i/8YJ1JKMYql9y/Fwo90ojl7rumEt+EW
y+F3fz1tTzHMttL4WGNa1dES1wNBW/aStKqaalpBpAwLMfEp/xU79H4ys4ctX5eQXo2YYxFp0XtR
Qf2O9y1CNoS+OsfzrNCJfW0DDUnP9bXjtsX1LKmBByQy2kxb8zpqJXoGGjtHOBju+NxKHUPsjxSs
tz1oH8Qxh1MUhAC+pkTEeMPMfbcQZQdrS9LTu4FUqJOPeJFyoYAxB+CD+QvaT9hKTs61MJYn7lHm
TCSNrgEOqXt28FRITem98zp+JyoMzIm8wOPkFbe922xozcTpbxxs5XSfdJU4rGnxMfLN+pzasP+4
hHsm4pusEs13yDg3ULJ2tOZDxytALSIkdlVS30yjJnglIemiCm5OLQ/flt8esG1Rj7XUsGdfStlr
gTjVKNdTXRm8KM9wsx7L+cPb7Zx7bB/Qv8bGpfRY07k0cHs41y2qtud78FHnAPiQThinXP5Flte/
Yfwf+wyotrPkWePFAUmp8CBJP4XvSqFiQoZSEURq6eoUQOZmP7cvRENFZEdKXvhT1enrfMkElQCH
WL1sRot+EuHelvGFcaAZT7jAeJGE5FQEU9HnoszLATo7vBd1iLRti8f+yQsjitSqwTFJJ+xqEtGe
+LCsysugXn78LhXNofqeJGbZ512XtCw2kUt2kdmHu6EKinKbUcskCaCGBQjjIKBwOn50KTq/++0Z
EQJbXGn7Ovwtn9cWhiCgaENlCQR+lLK6cDYMOvjJFOZEZ7GydEUmqUpi+W/DjLXhDgtZSxDDn++f
asH+cQNhhdFoedQYyGnBHUxsa69yBnjeXWgXE3ulV6SLkTCpfK4JnqTCgoN86hTBnWoJ3YuNqkGG
sHC9ssXMk85BxFfDuFezWCSOL1q448Cge5Jp2fcHwgcr38+ddeY7LS7dy5f7sC6N8H/cn5IxhBmt
b5PV9qbh+OLd/2A3n1GMDi70GKuhJiY1ZDO3E5Xe6nMGrkNVp41gmO46/WDaugjXoqclc1hToLCs
sVmJ38TMuyu8WwOVYoygYx9FwRCz0OTurBtAoeTgOuEScFoyoAjdG80wj3dFkw87016L+sbm9TFF
2uwSvdP7MXo+15hX6y7p24j4lk3oq7+cRC7gW8aPnc6BpYs8dbu9sjKGhXCcxcNmJT0SmPQiPh+a
R8SUdCLIEev+MBbUjXyiWG3MU8M/ViOc/e1oybrv1i87cB2MhRO+ZEEe4yAQu98sDgFVFh6F32uY
Z4/5DK+vL2TIeqUXLl9zYA1uENgen/yqwuspDJeD86m4EtrtuN+5jeOWiarb39Q7LtTLpOe8FpUj
4/Bm0KrLEznAH/Tq4pjn6crckVe0K7phtKgrRrdeOvcxltrZBiOJIlV4CqvxE8s6dTmOWnwFTYxR
uhQ9Dhsxkj9dy12nNOafB3HQfRy2TgZ5L+jZuRMlJY2YzvmWZYW9qqrdWZAe9nwTdR5MIcW6etei
xbBWasZ1cRK8cz6TuoZpxkBNDxeR6AhosRCEaolY2mipufImbT7/eaSIHAA6u0g4xXBQa/MmWPpr
gkvNSUF81jpK7hXr2tNCp5M+I1ft6/ZCR9nn/8HRbP7une9UUyHkaDRxcQyHEezsXs159ftqp5Tm
dxzlEC9VAE5xIS4u50dpdweePYEETB8bC68OwBcQmSmlNBIbT1E7CXFokBu+OTV/ciTPTWmr/hZD
NUlp4EsfbZbmfGnnpQXQ+PLN+I0zWh+8BX3tUMraLnfUJp0oAJLFtTrLULbQQbpKA7SBgGitK3qo
Ah/ASQLlUlf9zbAvLSwLc7GEO54nYe67eUjBDy29d6K5mNMx
`protect end_protected
