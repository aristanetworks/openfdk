--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
SKuK4ujb11eORxYyIFKjkXnrSlXKM2gaXq6Boe4VVQML4cvAXH3qKwtT6EJoq7eN3HOyoCyfXKqu
sOucmlucNnb9strdxKpVRdUFghkiVbKK5lc+JU3fo3sx5eXDOKdIiM060LpJSyjnSAzHdv2JUzCJ
RI+dNvu5MQSz6H3F8kZC8jyzlqv7SmqEGPhSUMdhEQruA+ZZe2WZSPt0n5t6M3FkJVWW8kGvIivI
OzgZyqJ/knSN96HhichZzm36w8p9JbiGq3wa7rV9g8KMAIn1RYbUf/ARPxPYhMlWv5500noNpB6T
xw3KaO+qRRP5SaeSfTbwWqmT1nI2pSVujGjDfA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="To0TdVe1Sev7UXRzaznz/c7ARC/O7CR2iwwP9dhI6cA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
FZLTvuT4iibPQ0Q0ATKAYYNXftG6Xrht2iwvH3UdffOnu3seDgFeO7wdnwK7/JJVk+l9zjy/SXLr
eibO0ySKMh+gYnaZf83XX4mIVbxEaXlNnTiIHCTBHEtKmZBhMpgpt++voI07qdwcpoKftx++0teE
Qg7ip33fB4praoToHzhmfbf70vBsJub2YLWDAOm5bl01ZM8r+nUw6RbJe8eIVqAA9w4hWuxeJSAg
5XDPinY3luJK3MJR1qGpTPCf/KlWVI8pBFqINkLt5bEX2ATqdqMhyR0MvVvbANHyfSmajboQxrC4
rI8AdCmatYUP+zOIupmlFlFkpTSicrtwnpqYgA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="QyZ4ZKAxPSDkPl7PJxAI3vxcd/ewGLMG+rHUv6uq3/0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3888)
`protect data_block
lBSmnuxhvlx8lyvQlFEMF+sLUbUHo51CdiIGU3NAe0SY+FKxmjnsQIDy3K2apvYz90N1L0nwv8X9
e+sirerRpAT/nrr18TEGlcnZgFSHYqgU/DRkYFWXra/PVJR/tVXuClD3Quza00wZqd21mSkJTROG
DVuDg4SZje9e0PrMOoSRIf0tU7WyKYnAEVENAuOka1t77SfoNM+CJoJZ3RAwE27/7Ycl2UckJ6Vg
atwMS/TXlM4WWvAHAlmGv2PhXS+3G09I/1BLEUyMIs+zAmgC/y+I+/lIIjpXeFgVDepTGdl3UdSa
ADjq6956s8cPY5+O97mECQDtLfYagw9p95k8mPJFpapDXBtZZkbFJckva3CRUjH2KdDZwDKGujQT
bbTkN7DV8biNWaPrpSjqPAaz9Zu5Hp+efXCx4JVFvIRLhvFXocBUdaBbY60ojEenk1yKvVjnQ+x1
jDXnJIChwWGd7qG2o0kdZeAk3FYtKdxIdrR5NshKws1+2LLNbAGUamZeqqObytBozNpT4R6g/TrU
dw+R3cBEvO1Y10FtU99INEUhLc8yDgpJ5FwOQz4jdlU0QSG0PgPUna9xvHyCOMQ9IdoWAJq6plCC
FrUKeuRDT37tFG4e9rOM957TxdkXw7XJn2iQ7zHT3/83UYjw4WriE6Of1+q4c8P85ddSY/Nj58Iq
4k9Zdxn2vL/NoRO1jZnV/RbDIvxWleXbVTDk9cSIyOdAH6Oud7NZdv6BTHJsvvyAK+2eOlsGg2m5
ys3wpZ985o0gAJocsa6AXk2dcKniWxiL9b8kMjuXeHWmMbogyt5jwt7hHBvTMgIafIm0ndlRRNWq
Hwwu5LZauf2IZisGbZ3gG2Fs2K0uPOZJowa6vXmqhIZli70pImrytZSGuVjkXpWHRjsm7sZdmf87
7vtN2ACBv2eKT0x6h7ctHnvK4VEGtuDHj5kUtYGqsEmGcux08jD/GGMCvfVFXwhaKh1+IjtJQBW1
KmvxqQDcPswm6paTJNZaPWFvy4HaVm0q42kXFm0P5xz+S/naQcTF2YDiCAHzKDnqjyu84+EaFNE3
KlFWj3oUB/hgwQEJ8VmHyzgHp4uZMP3ET9bUJojImAn7YG7PnoHjGh8AfMR13STZqqxuznD50eq1
dYJjz/6XEKjF2h/hALbo36s2TnT1xKWigCLql2rAt3/kWDSoDKj9GIrNuB3d0tXOlD41uRm29dJ1
dhDQVyD/M42cI9ze5D94wxA8pjkeFtEDl084i/xM2I5xjtnJbjvVlTKJubU88Jqmh1caoUa/sWy7
KEvovSVgMZQroho4/Fcyx/2OXAFKYhnQeBipXmJ7s6/muNewLpSoDYw7gE67jPK2B4FHqNKnCcLS
2mANPnNFy00x1He8juCGS05CLJg1k8oZUtokLZlbvBk8zwz6DWruTpYk8ukrwpZwFeALHuKePNg9
nhQOmQYNzQ7BdhR3Ldld0wIABByAgQukVKVfHXXfaqRgjmaRGEc7kQbUAR56TGaeNeeaN3g9pdK7
QanRuIZTWCM0d3ZfT5MAfQc8L5TV0VRmb7Prf4Fx0hfXOvVCDY0YtYGUxkNXbswcgKtz2Wh/sEgp
WGDA7aDxzfQCo3JCCROh3xcstwTxN5XtxtVRujEPdG/CUCH1DWAbfDmD1b/uiNaIfNmIveB2+eD/
i+uSHRHPEK1O0DTm0bkDMDk+gUMJ4PWn3e9wUwHHueBTKS0ZTRVEIm+xk8M43rQoHg13R6atZosY
lLhbDR49WZw1MIFapmq+mCmWtcmSCfJx0pv58dviBQ4SVXVq1nB2uAQjCrZVR97fG5yCrMIXJI9q
c+IPsyNDYPdzlygw0KIPWXCkAwt9mwAnxHbf6obamDmhfvhbdcnpu1qHnZI/+nOwHzkVmg7XDla9
y+/k2iXMZF4Jpa6D+BrTbbjcouBgBDo9s/uJjN/YSgKWzRG/LqkjLwB6eDeE1aEMa3q3ONi9K9le
WqtqeF0MEX0aGIB7kiU66G5ju63b4Zypy0yGSObmIm8R5eRncrWdGXtFPJjGVKVi8xclZj31EaBt
iLE9RMIji0QnOk+O52uNEo+oDVwIbyP8hMvI6KebBRtKVk6S3KwV/ZXHZBTl55V7ZIPk4B0Jilg3
ZU6E7DeaPkcJWzv5GiDVrrKToDCPqKTga5NRFpTRpqa+5frgz0DsLRAG1LLCQO/EmxlwiNFRJYsR
FxJKYafixHBG+F2htUKgPb8ITmauZ1qRyGtKQz7yu2zJmnmNyX8JPxw0EdQFnVcoCXa7sAuuw0vN
87z9bCwq1RXLV5ypC80Z+/9d4pPxbWvelwHzdeG+zKuID8YfUzggcw+JWe+5R/tNVIp9Mup1fabo
IksWdBX5BPaqun3c006HHf5yKyp7r/kgFuHcHRsrr+zVaNnWegaKFM/R1+KnsA6aIWDtd5/Zr4mz
p//2vU6CEDPMArpFt0VsZ0RHJua6ZoEvZ0DSpZw4oASzB1sqn43phaD6KjrOlf1WC2LOnQVC0BpS
Q9STf9pV7mAXWTyEWyjCR9/jUrWmj0hQVHAIeVgivE//LmsOHBEZm8ff1ORWtMjjVEpCNz80Eq/L
PZ+gvDvB+uduQ25cS+4WCqsepoB54a1i1fvYYVU2t2haVllsxhfi2g1oEpHEGLooIp6s7/bALgUQ
6VUulWr10LXeK5DzCsps68gJ3do/0RDao+Qrf9BnsvBLMaZSX9xWalNbwrpk70z0ZAoXwO5jShus
EMDHKuWE9yoQwIMheU/QuNoe4gxruQg1x7JwXabVanBA64TE2SOVJdFQoJ5xgeBUdrvbs38umpFj
ZnYF608G6qlEi+6Ws76fqQ/OwtvyhJDwbK0aZ22NXjsYDMLRG1HYyAIt4wTLJuw9xiqhptDwQdaT
h0n2yJ52JXN0ilAW2LZ8k8O1oSRH70E68LWI7z9nNB/Wa94FiSmIqxEGYGEdMMCbRcOVaBCZrsQJ
VnTbsugeULJQIHKCy8X6D4rYFxa28QO5BRQkYH8f9AgJh1vHOBhdOQ9fQKPYhVG/gxv9T7Anw0OV
umJXnXLkJaGawX7Oee3uoSGw5YDVFp+AGp/GiBzx7NaAtpOGCEPtr1GuE9qRcmoitH+QmEwTOMEp
J7LI4db1G4t1lp79U2h4ny+Ijd5yG2AsVvOCkh8zYW+GdDAOcWyLhY7RdcE3h/EGNPuRdkHJc9GI
LRXJuc9Dm+AMWuMYsIvJU1bBzVQz+DXsqZw56va75W+sA5rqRKjwvXuXb2fqJaDgZ+eBEaCXPF1H
6C7VWiVY1C6+zFVFTHKS088chakcyf0CQK/imLcgt6+oYd4Wrtoj/P0yw7kFsF33rqUs+fkBLxQG
9yqDKb4iAwThw5AnS3cR1ErSULgqQiwJjpifQJdX9bvJKr5ZRcC5N0GuyGRGredLymC+onpd/dYn
9/174Ln2MMK2mchCd8O2bxdhWS7ojikHmGXZRncQ25sSc+N6+C+Gw9bfE2Angpo4zygicAhQ3H1J
5O6OjeR2uNJxg/+MIRIL3LQudNux4eIopageHInKD+kl808HcBJmCc0FMjbNBTUTUQcuVXSfCl4i
7ZDWxWraGVG7SNR+cI/Q2lDO5mDP/MYXZ+li4revKsiicxRauEOSRamwnBsp4qe4u8ePqI7OArbc
O/oZZrdQvJgSHVbd/Z4DRywRO0KXlkchBCILcP68FQcX1JcfvQwe17PRMRfNuQMw6J/poFHpUl/B
IYgSXzVxRNNoT4SQhgwczXQai5oxCmq/OF/Tqxfg4GJgK7PN4L5dN2ysCtWCQpDp+uIOjzLBp2aN
fZrX073Kcl4SGKcOKaqMlNx2dn1fO1VlKN7M8e2Bdb+f5VF2pJhARMmlrLUVFFI0cZPrkdrLKmv7
1t3QhVhz8FEiVMRH1lrvdXg/94zw7VWLgGUAtM3ecrXyNQS1FlacNO6p0ygMnmX4UPzV29BoTsgm
rieKwQ/1QUPURHwSCaH5n6XZ/kkZaMqTdApDABYMdmRwkPMOAEYv/NRMzi/0Z7LneaFrHHfqJhur
CD0KPfVM7LIloo9EP6ceQHJNw4jCDIG819Zo/KWhBpW5aF7PDWzFZQYSX8O1YO3iwaO1ZB7oIkB7
HFR53kGHgoDwAsHEFcLDUH17rjfk1CHHFK1bMJ9Jtkf3MatQroBlp5Wm7w86oYZEvUR7dVtvy2vn
Ff68pPMv9+iF2sLK01eAeq3iVAM+WdIo9kzVC0i8xYCJQVuqZz9S5H4hm5MqLJVX5KLsyhDyuWpE
Y4Kzvc8+ESIRRQ8skBd+4uBTDZWOJavSn88Xim8k0DrJ+NC/nIrCrcmjTEDhI5l8KzmXIn26yVIb
mqZJBeCr38cPGOj7Y6ubdAY7i266yoYJgxGW0MB3Ad9laGsFxWCvmKwgpFkKa+pEqeDhBMwuNwRi
N/CSmKauZNAuU1/OUz2bjZae0jbEWd6NJNf+9McUHb0uXfxKyUQq0XKOE9XUxcU5HRDjQL5Rpdi0
AXIoT7rbGlVqNV4CUz5Y9cLpNgYBR8eAFokMGVF6j41r57At0byht/x/xZ1KBuR7ZLurZJDNHk2d
QE2TCmvg2jFktdgy/WeOIwiIdE7oM4tUV0UQfelhEdO6rdKRMTzrGanUuoqMk8GcjHWPp4YAys1R
GIHhqJ1Z11/P+hxrUZ1Q6pbVeiM5fuKANmL5Q2gM/JA579Y3BDgk4xkSZzeu8YIDyWweKKo/Wwut
BsmAiBwzVCLlQtqMwTHbtVfcNlbatBDn5lrHfclM6uFCLKBVq4TrAGQrBZve0KR5knTKpmgxkFZu
UtyHOOjIVLkg9NGnZcSCecPruf38eQyQszkFpPs6r+QPXoo8wOf0sV1rStbhiGhNTp68Hc+KBdJX
fi3JIBLk/LB2sEhfa2HJBCNtYT3MoKC2w0Jk4wWI+5A4DYP1CM+oN9OWj+85ONWgzqYni6THIkKQ
Y/CJdL7WuZt+IDBKRm5leN2oN/qI2LZzqwtOMuuoTCTrfTg4WbQ7ABpOuvCu0u6msOkCNcJZeaNI
QVustFk/QnOfrMToOhNj0mHku/SuhiTMcFaRDlgKqIPsEkenIX13hLFsLfNaK7tg1KU4FhM8dP7U
M9n4AcyIlb+q7tX4fqyfFkj1dDlgnFbTD+r3Yyu5f7NQEql83UO2TtZSlmkiM3tAKt98rIr/QOI8
ZHRrWW+WCEJd99ze
`protect end_protected
