--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
fTkF2oIZaVPhlbNlj7dlrtr027/OPCqSRH0DZ965t+JLbSWwoJxE5Cat9HQ0vpsYFTOnkBGF+dfF
Fh8jsr15XjRy2UNs5bNyl90BG0Ux8D6q7uwYC1EuEdJYGo1gpKcJwbnFtyFeXMwyRO5WyXidikw1
pvGnv3cmQtEid0URlRMyMRNGSq5h8hL8nYDJDrm48q74dl7hA6mbAGM69urypiclcV2MP4K8HoWZ
d36Y3Xdl3KEZ2a4Y5NktpV77ENsqrDv37IRx4G/nDGcE13owrLJ3du6v6VJ8ZwHQjXQptwdxTG6I
SYOF5SrXgIzxuWcPCRiNVUner8JZgBIJmDZbKA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="hfXKsPz6eSVVNbEOIWEn4MxIHatoB0j9cmtxv5laS3k="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
PI+5n6bieSDX/eKHppY8YGzwOAyi8u40sRHBSBl8J1yRg1DRN9U9xxQ5bxOd0U9W4es6cDYZiNwA
MhMX/tTxul9bAb3XgiHnO5hDvp5v7gQbfe4KXqCkddUDcrF7TgwPkKqtJ5wq76GPb5T+BbJ7nie3
gjoNZhZt8kxRPa6945wOolXsjbrk86OWGF5AGda+ic7D4MRpoC4qkXDz7NsJ+iBVG+OuKxZa3q2r
1lHVF7F07jvXDIV6I7wLyWwmDUDF8tLvUwsq47hzqvkwBO+K+eRN3WPRM90FGJ7pV84jZ07FwxYu
e7iZ6ND9yVnBG49IwRcX4o1Na0LheFrl0HdVIg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="+GPbkwCRYzdSVyGv/6gJelqvf98LbvihH9eAJqzrsRo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 61728)
`protect data_block
tS1BiqTyJ3kH1Bzh6R5pimftrBiIkz6xRjbObd7YuiMjOr37ZmKHceC8ekjrJ6iHvMsBKY8CI1gq
maGx1hJsMyk2EJRrDJPPGJ0B9h1dUThGSfPWm+Ku4Jp3/QvT/Q7v5qwPgglxsLjRbhtGIIFSZZ+t
rlFMN1YOcPWzRsPuDrQE4EJjCXI01+ku+7WodyrZkABGwmDImlBKg4sTsgcJ43t8g7pCRLwEG5yd
4gbz43WWgIOrSnjNR8g07KW5YzLZvrpVJeYTRmspEDryE+4e/5eU2GA+6Pb4uwWI484hIEBf97nN
QE43YTHolVVo1SzUB7n2nZ2cxYN1Kt1YDSFLteL4BMBI2wwX8R7UpcCJbRlIH0i4hWbvq+0cdqdv
8Khywbsn38FH07U8UnJgMZukSjZgt8jEHrAgsC3OA4NaJnkMJWxdpXYQdjIj2XFfeG99oTR4Oe18
QW4P8abcDevhD25RBf+kMofLYBU6/SGP8bFmCOz3kcR5ZSiYgEFhOf6/ygoK34/kMVmlBL6DJXEz
3nwxNyK2wJu4arQyCfRCoY5GwmZ/aXAFB+v5M3Ozpq0F/oHoCnD54Y5VRYbapMRhlImvHfNWXQiE
w71ZkKwur8z4fDqubD79MgoN3ZtCD2ZWrf8CDiWEFbjS+zjLYmRthsPUx4Y3wd6x1HmXKKfnHMPE
MXGac3swBFX55CtKock3WFSVDpd3tJBrIAlsAAN02d/Nf631//OrU+0/temMrFT1vugvnkKT2Llb
HCDOxIfSgdTcDN0ufkCBOn3jb5qqeHBz+aI374+YCqHhsZQ3G6p0Ahq0z56RxUyEvrteCHpos6bD
oQdWkUprZk/mkA8j0rEb2qOrgFQhkGZq3jqXfp67CWoHH87GvFOb6KqjIPue6PTVqROiWSrw0dQz
jFy8xrUL8vO06VH/jzlaEy4kbwEZNVot1I9cpcpTxQZroz7lqZ0/aK6kkgVb8gJXOIV2sKW+DVeC
FEabRxo190cov3xjhHObWfCnrSlCe3rF0MqTnZqkqUgbArKcnhmm6WqN7KmfYiiqWr7V4A6IUy2D
Nus0Bo7EuZV9F1SiZjmwaiO7AUUvWYkYMJpcnD6mwoUVFd7mGga4araAGF/8D6IeKLgDQfu+7rI9
EJrVCxmc08ILmBw/uWJM53p73XI826hq6EyZUAtjiU2/jdzcD/2BxB0RXd76fsbp/Fvem1UM+bmh
GqIlcJYLGSgVQ/D90jM3wZv061fnV/PIYfOjnFMQJVrcEI0pvO6JzSOoCw6bbrAgqES2UZM/I/fk
OUKFKpKqqD3TookLQbJEmjj9jDc/J1gG0SSKyqsPrzaGGHXVmGevfNspMQtbtc+gzXnVN093FDMF
gRlDiA0lprvRh0ymrAjgAnsGA5xPQp6IkEM7ROjBTbRO7ctYP1fmBoMYxMnH8mOK2Ev5CdD8roXB
sfL4hXmauy+MkI09jXSxLXwbWassbzX0ZLZOwvS9dkSNUc6mi9LhCKs67IPz4mvj1r0cpJci1/Me
qz160qk7+nMfI3/0KfI1WMLbZuiR+me72Bj8AZpVIoQMqi55LZyumdafAfbu6aiBFbUqgllT8rCf
eCizFjrza1inVpLGxZ6iVwIfsbiRZrqZlqo1S2cPn1UXZccqRYTIp8sLYyiMv7m8rH/dt1wTb1dO
9nsJnqhNQiKv5QeC4ziT8vvpmw+vGnPs4lyutfhTMfMCMmMhf2G9S0v20ikatnCZBhThLAZ5Qqtw
TMVHTwcrSFnuS6bZNoUIs53wa0/wnTt8khaHHkx3Bscj2YvRPK1TFpLc3VtJ4pVBUGFsYIsNb/6i
DxeHPWi2Un0PAJh03Tgzl8zvz+Lab2UYf9wS7AhzxcyViNVoc9kDOwNw4upav2U+oqsyb+A4NWaC
8oOkFxEomMOoPgGEWeSF8nBSLXXnM6rHLYV2MGMwoviUnnmm2DmyYA5QRICRhtKgIMyi78ftULp7
1ujXn6YozXjywjKfHFDZm4JwmaAO9GMDwbHvhatUL3YrCK0rrv8LoD47EFyxBh6DXFae4kkY/IMh
KUS1zbfW2Xlk5TL4ip6qKpIZfHNC8t5xRm++h33NwvvP7xw/nrpxpYu7NPvfU9RAR5KBie2zvBOY
+u2KoX/RrC2tznUPaU2kFVgbMSxVJ1535Aq8ug6nQwtgKrme1XmFeb5eaJm9c3VqcdgcRCX0mnEI
TN87iJ1Tw/TpqvvLZ561/ho5fr4fGNoQti5rk7ijg27HHqyC0R2GF1bl4MQd5+sJrq9U3BMpxLf3
1aoCXbUGJ6c6xWfwTZqkmBAJaqaRhf1AUzirQaf8oxWCcjFtzvT1DyoBVwLKEKnK70RR6sSESh/Q
We31NL0itMgL2yfUstgu5o9sQOAIVBPaoyxbMUr3F3tdQNeyGX/8iLaGuFM3x9KHhVAifoz80pDB
6ChJeB68/hrlkdU51Nx40z55FWyJqqlbQqhOwxhHSiA8jbMyBRIXPHE74MduMbv3ARDngOVqZl/K
q6uKQ6C45dk/21YcJ2sjMXevpP/Yx7qdsI1MG4AZgPuklRVVGOF2wP2TTj9sBZaieUHPBFJo6w/K
/K0rqlGtN026U40whGSNSQ6pYsYrwasjD2P15hcdJE4MKX25TrEGFgZzhPkvyoaGqkZUAv8fFRdw
Y4ZHBFBrOSYqgcu2AGzTE4+HDourJSAGylTyYty0nTKpYpT+rAZMcei6rDNiBcYHGeVIn2cgsx8v
ZA2EB1jAkdUuOTz00XJIh7lJgR0Tpp6frGWv+oQXnY5sk2cH4kHS2fffu3t69cRmJXdeadGCNCS5
cxAIdky+5zlDNQnAxDcb0nYZXI2ObnwaRN2fTJuj6m0XXS11nIpqKJ6Sgh/qAKUsqpmw4+rx1Av0
rIrqgVRcOg3wgHPAjbvpKcZdCDsluFpw1Euf0IT74rOqGJ4Q6GlajyhlFj5EV+xB+WrifuwO6Jcq
MHhYYgaEoMWwLKSJZwUxPQsivWJb4Gd58y4xFfna/NRAKgMLuqfRbu19cEHusbIAFOFv6RgfAN/T
i0ryQI7MfYoHnPzG1w1ch5hUl5/KZtmgPvylD/uSNWDdfbGoZOJsQyrUPXq4E3TSg5nsAFOVyx4E
AXQGGC2/WPCbWXWdZ0DW7CSE9VbULQah6Sv+/pLJXNwVlx/bhFYxelbNJu4dVQ7NhWms+fUOsdS6
UfrCVfQoqwaaOxrw8fypVmV+Ft4xxMQeCTvSfGTH/6B4Ge0rmy1NPORFOQoFCB/nleLuuu90xbz/
y0EcF7r3nHI/p2V3xTO+kwIshvXGgxAZioc/4OWEKYdYxRwSehXpLFcQJrcrlmlUhdeXlaSDdr36
P6la3OFaQXdSV5oZU1H618hy585TNrx7vg1iCbua2u7DIzFp73/RludF9cg6JHzgPuflxJGi3rvG
qIdaJodIDBxRIeHO9EJYu5E6EKMU6uuypgaFPVEXIfKcZ82jhEYPNuB4Q78pBjw5QVxCIYBBfFmB
VRP+KaY1Hp8QZmaI1q8xOALX4S9/B+gbcDXZcTPfIsbZlTH6e8hg7rFDiPy/hkT23l0VOm1W7hev
LYom6FWO4GfeseaEyjS5b/1khbCk4O6bwmPYLA1XVYnrj8EbPOOnY7TRNLlHiTEpTANlkIwW0Rmb
KmP0s3GWc/D6sTH9D5wztzr2dFfJ+W/Sz39+swPMv2siWNDeE17xyhStKipH8rjuur/lZrW2tcTW
WR1arxX3jzat3oU2VJOflov350dqPJWWmVHsptfAjQyndlxmhNFdsZjTU8JXSpyFY+UfmB1fWBq1
3d98oV2TJKhkklNr+Kzo2bq/tal1jBoDWZ3ZI85gU/ehdSnQ0GEdMpIIZ2iOw8q42Hp052L+x+8a
kGwbaTWCxkYBFxLtNtb8sgPjUpG3WdO6BbNwDDkudo5Xzv09260zfq3StAGUmczDQqTo6iCGEfDj
rU3afCXmNbG8pVPOHQarXKPlY2lamChj7s9ijG39fcWhjFVHg6N1yfnIV1wZ9Wx4vN5fUZhC3686
Lj5/rxPfhwjbkjxUoQKbi2e/4JvQA/xkFIt5BZ5wZ+blzHG+r+mhkrSUpSASUdxpC8Ch21D2lp7o
SFtyza7GAb8SjLsrx87+kMn34tKvMBzceyOr4khYS001Vf4zVnW9P6NqRFNWbC7O7qL6/ZB/lgNi
x/uZCfhXwvCxm48oWrCyTh1f39maLyS7V2Y2Cv/zCtG9nInmFWSbQ6sQS+8PpuQQwnewpIVyZR9X
1RJ5h7fQE3sjPnTab90CZupMFMfaATF8GEi8mwwRONJUFFuhtQ3UEQqoaUUwiJwVcCd16x1cZACR
D4T+MLnNy1nB73lZr4lAzoPDFlPNKQLXhOrmBenHnFn0T2CBH77PqefdzOydJSVFVfp6kMrFvf0Z
oBjzOvO6Fw9h/h5+GOTS5dEqNPHCfx3E4Y/2SIM51tyceXUSGAgTttsgtKiAAgHXFV5GYz5AZeB9
JTZnwp4KjDv+pSot2Xqo651bNJTpSr+TnZNlN5KcLs+eDlz7PALp3qtRcFfwxPodTJKYLcWtM7GW
6LrISz/wLYZDVhDp8HDPEe3w8DSX5cw7u682eXRmQgQoZicgrE+tXzr9IQMChLv9jnYmsAsAbgx1
/NzFrxuQ5w7Ffy5vA5tLkzHp1bvay2A62eTlPSy6Ucxn3ss8gwQZCrLqeCe1y4P8vnFxxLKCFln+
AVY/3SoAwudEupbUGiMXEN1GCELZTAoS3qcCV9+bLld0PPqiXbKCJJTR83REJfBnsT62f7JRpzja
4XHn7FOwgXm+HbzAW6voCOOD93Ho2Qxi8zIjuEuBmM5tvkQymGBCOHCgYsgBByaou7TLxGhCGU0w
aRHz3ojzTbajmh9CMpnT2wdNlHRsS1XubzPXpB+Rkc64kIQTJ8ZcBe0DFcy3LAjPL80WIRb/+sIA
ksRrKHyyX4tXCJFpmja7mmoVeowZ57egYGTphO53ksfFr90gLhjWungUbcjIYo4o+/Zllf0ElaY/
a5ONWJ+m2WKnfXhc10aFeP/hlzmA7M1xNz9FkLSE2sBjIUX89jLWcfs6awoV7EW61ceaIyCVQ4WZ
b/tBtJwnUdQUdFgQK2F8mChaP33x7WHiy+QAlcaDx3w9Yko7HDb+ZuIrO0XHCXNGSj5b2al4MXEr
7K6qYg+xPLdS78ek5U8GUEk48tL6ZVyxMAJcYHpvuTfYiC84t16T3gvqKJZysEKo5tbklTyFvuvT
xU1vpZSLNz/TF/+LH+/qPbax/rkl+fkfl+dc6J10R77oN7fWlQwf2ruyp0sjfUNarHmC30v0QVpT
zUjdruh0a/u8tuu5WL1JXkYFGOohNsSGVWA2eEXUUNBc3CHK01vt7+IgEJp+Wtc5RjO4Sdu3aiVi
ScdVGBna1X65C01UFH3MDHRRF0Ajl55xDfnoW6qdbXnVYIQqZk31KFzsoh/MSZNihhKuOLmIyTD4
qncTcjPyPFo3LhVDaKq1ltleEmQcHcDD1ZYRKr3ghGmfzyc72/ffWZPSOeDQYuyehwQA19V+ksHE
suX9yvs7b/cdNA7s5dRI8h90yxsfJ4O3Fy3k7yF16xIChH36NIOgx0u3/wl4JWfhIlK2kevOLvMy
EhsJ07duu9XPNKO9mwFtcm/NYezyCkIm9+46GO4VE+Wlshf0jis79S0bSmGPNWZGEgcioKz/p3e+
C8/dilY9BCPAfcoM1H5o+JdpCoEWSWX0P0dAiBm06anPP/OJS088F/ak9msHFSn8h3b9mRoypVuk
DZkfZpo0CT2uRcOFYtf60XpjxnqP6j3vkt2B99N6DSwi5ZV/FLba4yEXu27W4dTLYe0upt/WUwZh
XyJnXj739tbCUN+hDDc31q37GYJ5jSLY+NLjNB9Ot/d3t9e1TlBW1N9p8gJ97HQeBsvyOYophoRL
+LmzcDPcjZMIjUMlijE2t/trX2kiYX+CAdd2clwWlvHyGtt1Ynt3bLpAzrUaWYi2m18Kr1qH0fUG
WFXrI907vEA9GcvXBDkUVaAMj5DaL2+hOPcHyJ9G3l3E9xkFRYTHpqbzIFut4FgNSW/IeT4iT9II
YZ1f6Yy00qOy6W44RUk7JHD/I4I34zJ5C1WzGRUAiwWEnm9QDTfOR7bi89AzrvUqKyrzWqMWqVKD
pgIVpdkIYBRKkdfDXPcaXkAJbr5rmQaT72Y+UCMuYUlqFM6L+roOo5Mfi34aI1zzMH8sfTMbBtrf
TccKszRtw8AKoR+U2JL+8ws9y1m5SU7Y2PkLcmRa14R8c4ZRYedaaOaFDKQpbm6WyqUUlw7cOlK/
pHCc0XroL7AQIkW3w0uweKMJSNBoElZxuNhAEPHzswcmXMmp2c/xCYMdglOVA/BbqTwkrgXFeJxd
XetoTgYnlgimQeSpQ6H7JSrbjNd464sZRRQSTxB6KFmliWxvp8iisMHZRJWZbUCYjGgufzVEPOMF
WwB/gM2NX372H5/gJ+rb0pxrKTEe0SKhFMUJp3pnQK+WVX8KJqjnbquK5IePVeeuI0dPXCTrUV8e
o7iIPT2Hn5RnRmoLKmCvbIchYXvB5SBTqOvSwcx8t+ESWlmobG67z0WUwfKf64YzU/IA3GEzd7lZ
SYyV4dtpI4ZcYl5+0tpyqDLW2bdEyIBn7Byrj/L+CkdhIr2FjSEdcv110JduTiw3gGt8EcrG1rfV
PpHPq/i+NQ5x7k1REyBS3X1Zl2AwKkqbd5a6YG1mYWmHGtsyYE/fyPeorVQOBCtwlo3SE/cY2+i2
7qHODCO7mH4BxheeZSHcmMM8kAplwFJca5xpueCfsWSmAsJIxzrUMOvlchOPzMwyO/gST6iEKdTO
r2iYNAtS0HVM4cYNhmuPcQ8LOvbveDuoSjXdqicxuoKrPKFn8Ym6EKIQtTd7PZmE0fJLcpvtEq7Y
s7X1K+3YWFuvf0YUksXboutacbwxoAf9NrBCsg2rWttn32UaWCdkT1vF7TE/o9gfufXDFEGWFgKN
hAEckWQgqfOQtPQE3+Z0oDIvtXRdtU7R13bRI8fZ1jTgdpN8vKbhyTS1lhN8MOy4C8fnICPcZ0be
Ifa3Bhr1+I7WAGn0UgVY7sB9x1IES6+JAlIJRRXZEfMcX4f/+mPh1AhuScAORR4ovvd/M78Rkj7n
nZ5GK5d0Rf09CKr/XYYJmu0jOTptPYhuDJvdnrzYVcJ2K2yYf6ZQqBUZbDc4WhR3rJ5aLoXwAJIA
AwhsbmOX+D8H/e66hPjMSD57Af5Wcgs/Bawa46CpYqg5ps7+a0PrQCz9dO2Fvu0Ef29zqTCvuHzm
uCPQSk0fqdqywI4ymKgFxSsr9/UWYOJ5L75TpOF5Vq0pCj9B+/KC10m76Scarw/jVmfg2ViG4BH3
FAAXUo41R47dneszpqyyBJPidVw8G9j3aFfWmaygkOt3dXW4SKnoVuK4DHQSO4LBs+XHEAHOc9B+
0bogXGGuP8fS8ofefQUpC+70JH/ytPrfxwgXNx1zAp5VthroYyb9YL/FyLc5DF/qI3qp032ecEdD
P7HZlZX+isVjnBoVhE8TlYMMmKgr916iJuthVE4X7sbKaLdHaARJfnuJV14Ou8SG6tbOstGc3/sf
StYnMBRsgogNL134g/D6bf+JEHSabMOkL4yJv2uYufwtFCbb9WzoY+L4ypQO7LEaL6P5Xg/zLhOx
EmN2XGTbGmr8BKe3Bt21cj6A2e46F/PzUHelM6xYVNQngzOMNcRhPQnLehcrIlKvX/CPdVTr/llJ
6DUPilyYKMBM2qM5l7ac1AwxoWNPGWrnrIx+Tqv7HcJiOxzbC3G+n21iD4hn+xtMAEw8pSSZIB48
dRHqT0h0twkTMKE5UTxpShbJnKSTiJufGrNe8YE0GoIvZtRQ3EknCmfzolx6gW5/lfFjyQDQ0IzL
cA7y0aEtdYMH0Iyx5NWc0mbP654QSFC3/8eYkvZQkNMICtJ+fem8bIO5ThsKzJgXyWLYQkVa1i8A
ty9dRpQC68rMXCdwaSAri+hiTg4vPQiP9zzTF6PnXapyOVT7VfsLCqcAIWjIHto01V4vHYzukcY5
W0mM7rd6SA0xmRhxB4WOUt9J/UYonDoHX5C3Kmg1kfyO2iWZ6M01Wh651Z6PmzSH0mxyB30fGazn
ib+HSmTJSMlOxrfKycsNJVR175WC30owHR1RwkEbkJ34Wi6S3EUX93FR66+0AB2Y8KpMkIKIrkD2
myo1PAC52/NyuQ8UkH9p8b50ZAV6cfSHNugA2zO+NCwFR41pECjXuAua4zDp9l1yz3+zK9L+4RQV
WhNfS4/J6xUBUKjtTA5/OSril0C90HpLAsQHWH4/TH13CMZyF0ry+lfAAUajP9BIP3MmpfBgFq/A
WTV8pMBn2Q4edxCurbTEOEDjGwkC6Ly5wbRzwtkg1lAMMmAhP7CSEGwN1iR6MI6AXT8XgoPGirZP
Vz8d6E1nO/cQJU3Nn1cNbEeRqxgcvBtK+8f1vfwHs1EkizNWuKuC7p5aj1iBmIgOgtM40AQpKKHl
IMszEBoMNlnI4F0xGetTowELXoQIEokHALGfeQ9spYoqAI5uFlpy1lqNqiA6qWunNlybcNTmmE0N
kdA5FcT+Oj9PPTW6ZoGzwNZYSi3BbaJa+CgEIFnr2d0jsgaz2bPEZVikS8dBNDJCJ74/Qd3BKJzF
bL3CNT1faL1agCJF37B5VAx1xYsxtBtPLKtzsUoTLPZIMQyzlX6IXCDkfoi3bT0S9Z6FFa9d6uhx
cuqh84GQLliKj45iGNQOzTvGy1HOaG56Rsjf9/06CObCs57Y+jcvWAMZQ+NBVg1lmt4XHv/RRe0r
pJXaP+uijoM6zDq6i7GQCwiPHgTtljfeHze99BD3YnwZyXukMe2MYmY0B9PS7wXf/i5oqI3Lwj/0
tg7nsDzKFk+LWtlXy+0XuEEGkfI24QmQ2gKu/gI3VF4GhB7ed11CXF2n26wWtIswBpjR9UQVGNrE
0zpbo/HU2URKliEC77dEVhJ4kGWSYGMnA+DXXN8WA/fETQfYzMsIiP02r7LTYZf/nQAz7sOirNQJ
FimQVorFCc4XwwDFG/RZVNG+ASl28fhoF59g4WUCJ7dkLpcjA8IN568dmpp+0qN+hmMsSY+qu4rB
2b86iD1RXwh/naIKkcjMoJDcv3UmCFxjYZNVuOL0anLvuAA7mWiGHqxWDSMKPpd1xTBPdXHx8LWN
o7jXEVXU7yOMRQYtis5oOvMk+eIGVQTjCKEVPEJzD92d7b2VElxVMwL2Pl20BtECzhHzE9lPV56S
Ocuu2Wo+h20GWmrj3rzO739izV/5PbdSfw1Z9B0P2R+J/bwMliXzzyX24bk8ZJkTDQSFzrRR76CW
Veb8SizBTI3gnhXoYp+AviSg/IK27Q0ixdVQAV9DSRpnXtMIeEwU0qqHc2znlyumxyPiI0Y7sNqB
SKvTKJw4qGa7AIgV4M+a7iLJ176XorNURxuRt7Zvnj7awEuz7eB+2ZrzlKHc2wwpdeJpPcBxzBgG
+oE8znjVH4OwM5tSd5H5bn9M4m/jBzeHrXYQ8JrhrJ6mqtyIq8BqZNQgl6rUuQid6L6QrdCxYHcL
TKT57yRfCueXw+N4SAtDT5Gq16LD4BduufzUMCGiCrGsB0AJwg3uiiMh8rpnakVb05qgg7zG4Y76
6Jh2rxfhxQ+pmsqAnS035cPlWQCWvzHKQunbNprtL0ecd+7+5MHK4M5AIFt55xtVFSHCYxc1b8JK
8IyG9A8Tls/JBYG55MTr+ZUMel03ZydGo2kBDtKa4bnHwkGOSb5sXw/W5uohieRqnPW7W4R9Kq97
6BfRP7cieEin/yES8pgusnOn3koT+Rz1NPR2TyiDls6Vn+4Wwj6CbdWpKaZuEtWRaOEyYKxmabQ8
/XHjShUo14FXyN/KnLLd9frrOQGnXv9bV11Uqu8lnse+/qDRmJAlaF6HZlWCQbQyWNO0erNQqWrP
akO0SN3ZyBEiYnH8+UTP86oVXuq2krMonM+1llObcc2hBQlSm+eikTvSShTLcD5aHP2aceP31XT0
4Yt6CC118R3KSkWCkeWUcOrx2OfxnVjkCvIpvDX6Jo3JSWmeHykwQMKu7FLKzzbAzPb46xRZuchz
F0DdXqxKGbcIyfvoLlF4jv+EZ0k9a9s7a8s5MlNM+3+hBpZg0u59j3y56yZ0+m9RUpwE47HwEhgt
Yqs8EACN79ACGYPM7Ta/GpIXDFhI//resWuQcvYBHaSOAyJ0iK5aKBWfkWUlZcSHjHq6MkEz4BxW
k9xaSou3OwOfO2BgcAOr2tTREItmUGNnH3fdxOMsnLEepVEN8X6mxdt6F6eeyjIZ6VeNciT5i9eV
9AzgFTWzDztv3x6NeN8dfqNAYIiXeMTHffUoxJPUF5/f2Mn4YLBDuDpT14Ko+p9syYGKu5s9J73X
p82BRUzzyqApqgYuP51MeF3DojbNmPRqjsjZVLNBAkNibpUK8y4YIZNARTII3jZE374zUPgi3Z6m
gA8D2n5N1m6R6KL0/ycbXBuH5PU8XnHNHVHS2PxJF6WaHoXKb5aYguXnV5vs8IsdnzENS3HF+NNk
Q0QKE+ieljAVI8Kjkvb3toWLG7JBwBqnp3nyIMiij02eqJfdsej10rYkt2zJqDD6FuaJrUzKCL0J
XhUM3kqYkHOU+YqJn/e0SMXeSUwbCGmu1kBdH+FS8r9CYoC9nyfNi+NMY93vKuNZ82ukIZmJfi/A
DSn5qEZuVGC6PQlZ5iS7Jz7MfyMid623uyGBWMIDTteKc9cdYHeoJCBCQodXEhmCuX7mMbZ0kjMG
iDM6dbZ8uhzAcWyBh7c6Vi8pI4bYAbI1OYgz7NsfGJQENBqoJUENablqGzXouJyYxiN7JDsE/INc
sMAGLvfWGNM5GGkOvlBlYyf4fof7liecnZAH/5xaw1UOKFkEzkyv+2zZQAAN6FexsP0L4aMj9h5A
x7Q2DlbstxKbIUg/Okg9rKfM3Zncqkaf+X0kLHSzghoOv7gT/QX7c3Qz38b+9VDB16jg7NN6WboG
EjKb/VxA3ZkUG5+6623rwITU/9xh3Q81OrdXK+C/Qw7XH2KUJLuALt1Km+dEdic/dyWQ8mUA0D7U
otTNMWe0TBk5Y1l0isGsII5EEg6eDRqt+j4TAiMZYlOxs2hp5ba7fqYbQpGSPkm7S3vxHEUPO2Se
GWf5QBeuczYuvqDkJjaA+DfFsD8Ub0P/38tICV2A1a7izBJf8GLtX3948USi5vlRLpnp3E4P3xbI
j4rWdQJV+oP8YWmHHEQThXCKgVhFDF7xI6pbke04V3bWjMSb+DQZn2/y7RkMMLAZjEN7LYRg6cND
IP0XQJuBgxzw0kz9yVZIen5B2tkFWMqnbFb/hE4YJDzevaElwrnSppnuARYHBlIjtMzNp6kcYO1C
Qsq6jB6H+rQtrDxMX26FwvmpCPUeTCOpgH2ehMJoEpKwZnTMddsZufDEoWTO11khXRfBl/qsST4G
byQX6+TKrTFpqjAyoGOiNUl8EXR0cAYGjWF9eMT1MKYbmhl/n/KiN7KDMbxccdwI/rKb8fq+tExW
1fSC3QCbOmaU8GsuZ5BIKcM10ZLcrUfAg7HNYU1TrQN/5JQ4tbTMY3ADn9MvhIt65xXOh7njyfra
m89j61j5ECVOn8Fjw2ertOJA1ZL+F4l8FWTr9jamD50pKt23rQh4h9s58sPlLBCyP8VjCPIhXgZA
qq1mWPBSyYxlSnyRQablASlNdv0L6zrb//WNo+AtfIXjxCYHPh/78K2zeRAFWMO0SQpi8V3gfUfK
93vGyCcr24Cn4bNDODxDecyki9WwHTdp2DllrSvcGmhGB2rIIVbX75inyz8vZohkO0OwnpTYUEWw
CMVZt0UMIVIVwakLVvnPpa1UHG8GAWUqp4030IBWzDt/N4GI8LTi9vshcculXsCFAzEq3WeyELkD
9+qRVRfhR9Zadv176oyVr1cGkhHbWW//OY4rMmet7jy6YD4dNmntFV49JDJeKijFBCnPyGXcGUcN
5+HTa0qSaCvbhRWQZUGW9tVs02wBsUt4I+1tKZbNxi/DcAv7Yt2++cH/Jj01/nslYxKDxDyBYyqh
M487pcdUNR9+buQ8vcqW731uTdgEK53lrJY/+g2xhwwRUUfKarwxLWwBE3YoEC/hg0vecmOdmVl7
UvSWwG9kEhirPpVL8qNMg2uRxl/UgyyUQknq73LDRcQCJtVzaXsmeLGHF2aAjadIjrMjti7sqjCK
IBnkZpLkgKzcMnk/UDNIX2+DzXiJL5QdCLbo5tyy57v9Gax4Q/alP5tw1Pl+XOgeC9yo4N0flwoZ
oz1pJed635Vz8J4yziJWm5SGCYg7y5gFw/2fUi1ZsWTMBGcqecA3McA4PRSq1fqRSOpNzWnZJ7qX
zvirBTrmhROvke3+Eu7fMeRBzeYf2qlKWKqbeeDjlLzkAnh1qgP5Jo7hZpsCO3umjZ8Dpi3KXBBg
cfHzwDvyya40DLyVDjcYxas7bgQUVzYxSDnn8giLb6yhCneEl5d5uAQGjh9HF2b4ye8tSHYyMwZe
N+ePFYMvZaeEr349rth3i/9WycHkxsdfY+uqhvy8dJ2WYlzm3vA0t7RF4/ZdsQHQAZ/PRIK/Dwzc
IIr2Gaizkrwmu/oGsk6C76Nl+leC4D1e5dSfKndqwj7ZSBCVNE2haiK/ekPYVZRlUilX0K/TDQx0
egOGlRMU1u1uKix8HCsZ8l2LslTm0GUh7nvl2uFoIi3Z+TDGlFVi7flGmPodIxswS/IVlQCI2cud
vUlnYXId+sFEca8KUAO5NWQmN+0yjlb1FYdFo0lgauAVJ8fcvcEiDlPVJjXip7RUFyG4eEzrqH9l
5YKiC52YWK3V6bIA71iczmqTeEpqw6yIyVgiWneMV/YiqolTwRKm1oFZgGlpUqh2NP8lFxGZ2EMR
cAQn/Wk1UMyfJihdUv9llmpt5PxQYZJn5HrzDZI4rwjqQQkQM3J9HVZKsbU/AbTORR+xEzc6oWBs
qnY+XxHVSdkTqQsUh3rhKyMh/P7fSQBOikRbpLz3+UepJZkq9KBOznvoik1ganiextFz3c9KnPLl
auQU1rdtGBOlmisha/yWSReVkDWqgtPhMFevrC16HFnzmAlaZ9FDTZiheS9614cCHAm8fHptWNAh
RNMg2vNo1C2vYDAMkuExjrZipl6jPD5Ak2D1Jj8h00tFn87FogiqnWKeCNEVKbBRdlIrDQ6k7emW
PcmLlSD3fAosPjFdg26jlrRDRD89UnttQtJPlLChyIWHqJ+qj0QGkj+5sn/2GihPZmu/hyhTeVrd
psZyWKiulMd2AXSuKNDSTlZf4esTLI/CXgJiCJbmahI8tlHIuGa+K7IhlsYGWJ8aq61Ycao9kT52
TGHOxYN0ti+BpPUFCW+QkuWHuG9WRU/Kf76ZosWnljB76O1IL24arjYqeOwFxYITDbL73tUgi9ww
arti1HXxxQ0kBgieHqZ1eqcDGCmsWXE4W7ZmKx/LSIYipuLkAXo5Hmj1zsu0jgyIsffL6QNlJSX5
gLVvn75Vt2fEzj6+tX/y1myvOMoL0JxwC0OdWFne82MC8z0DKIduS91RV4yF59clqTonb1DQTnHE
NbznE8pmmlOz2kp7akYdSUE6GbDxpLrsp3RhI78KlXKozxL5xWEoA64j359+JypZLoWWBvvBvPbB
3VQZx9Yb4tjjfhd/i98qjghVcPIVAGr1ymklUuGbpLkOZWnUBLa0ld3CrEhQtRNNLnaewuAPwb+/
7MeoaQRj5ovrmwPmur1qI6+YlPaEkOaCTc+ag9on/rnOQoO2jl9KCopVqUjQuJ6ImKZSy7qulcbh
zifYMCuyQqRRm7xI+xDSxtc0PvwUz3qiyL9X3rXyKWjhqSOjEp6/SJWyV3/7xicGervaoVqVSAZn
i2FwLrZt41j8P9jdtEmid7kxEDPPvGkNzmDMTtJCWqAct5/xHrdZRLrITX5jafHrzC6IL5kCx4ZG
qUN6OIhS/11EqhunA8rAsPk/HCFMzRRzOCm1aBqpgYHmLjEl/5jz6pyqCuMhTjHRX1uniX5QE0Mg
ICYJC2hZbTcvgZRLkAz+NlXwOtfwiA4T9ZZsNRgtcxOTRHebLrQ6roUmpaf+zKETRF/kfiQ//Ndp
feMxgG3iYSinf00wtF/1uVi8hES1/PjjkCx/Vlc4WrP6rZexu61xXXY62bg/BhWAUw1Oeu5U8BbB
U2UUOh7O1eE+uHuoRwSR/OvfJYhhK2/ahvyFoHwt8n8ukX6D9KJb8CK6FMEn4l7wSHTinA6eqSO2
6W/L9+gvd7XoWog9afmjRDquvugRfLQoA8s8nW6WQLWDfDZZ3BFcmY32CMq1oV/VzoeZuHqMDvkl
PEWn1T+hXsETNtkFuYxMoa9QKvLKcf8ZhGICtKeoseGY1O2/ppRSQ1H0nYYuXUCOjP8XDnTmIDsx
oVlWQFYEOwbIc1F5EayrOX17J2bTGeZHBTONpFH6SQH0g8MZ/1f4S9qOJKl/kPk29lC9sxmVTIpB
aTPQ+WLXNdaYF3g7SJ6gaIJlxw/K9r4hMk5N4AkqTNtepZE4YZdAmVPwZE3tMneDYetqaWC1lAeR
Iw77vhquQZHoZ5MNbp4qDcQYNTblzpcg9kgNi3H4LlPUuYTDqvDAWNYmpZep2Zb4Hn3dS9zIi559
lmnAl+O0Ym+DbCgJJeW/X94chVkOWRpeFhpFNWanLScJq7lHvca51fGrqgWbST7Vy/S3am5Z1iW8
GR84ND9QnnwsaHdWMBJ1+5ZjTPXmUOfjd+PaA82uJZFF2MfwiizhSRKKZ8kzfx3aP5QCCTwn6Egz
vMouWL3WlQsDC00CyEkPZc7Xwu5EekHmWG0a0iv76kzsBs/xr/AcLLXodJ8hLMXe+yLG2BEU9iW3
AGuaC7o4C+gKacfkB7Bdh8DKhycbsPxkdACp0SHaJmsaAhrZML2DHo3k8JUZdzSCIvI44pEZU5qA
DWm5OSDWrdYR0kB9hMtZcV7Oij1aqIdT4A857mZm/+onDVlQOljGnl/9h4GBhSWbwDmiTs8F4huG
wLNfBBT5q55trhTKmWqzKV5TRMxOT4O/q/u35QuxnljtG/cctUrIYRIX56zbY/xeW1W9QpQdf178
5lmEkXpEMaNUR/WYznR6lc1C+DsimWjbR5keDgKVgfsC50CVMQ92AQD1oPzmg4CnJbg0uQzZhiyb
JkRzzkJBEyqFx3CtTgEJn8TZvedeOw1hnoXjBa76D/1eUrN9ae87tWswEl6rJc43Wtr6QLUT0esD
CHJ2qucs1Yek3trHo0hT8J7Z2YOYgNx6B5R+qDgD1/ezFIWjRMc1RPofamBwBTxDAkeDgQSiBNHu
FZXQ4ghypYmTi7p+vygn/4CbNv25qqcrenGI5dZMzQowCetiAm/o34PUbNxJLrFgmY1+aNSLGGw0
rDyfWAX6Uf1f1+qEURls74S7P3DJpKPaS43O7AuxXBdN76yb3iPCWLs60zxqhHchoHlEGoELI0rh
STL0xxaZvLhPsgGnGxHymnFTR3lJNiIaxZ5nolvWnjNqTe17IC6eG45dAFH8c1gEz/OtoYyMSHXD
9x/4fDaoYA2xa+3UAJWhLmpRd6LhGPyQR4lSRp1qljiocmDKK9f0IU9mDXQrhaLO7912arcjkFFz
c9xDFN8V7jltdj3zz7sk7r7WLa9IKRQoSIIAetxKgR90hoSzHzbjt64wVrU9eehL3m+ifZtlQbsa
d/1A/bzbq/Why72NSlcqFkOIP8Epbpup2LD1im0hac2QQT8hTYlKoPdgD7ltQws5EITebk703oo9
qX5RFjcHFH9Zn8176EkCVq5EpS7o7LhqhlXObaVKBU4OcpDRrW71m3wO22ixgmS8GqWHlhzmD0mN
IZyLuO9GNNySrw9UxNfOXo7xN+a0OKyZEofYnxZtOGEd9m7z5OanbqD68IkP0a4CsEYqvi2Bt4U8
Sz0G6+3sSz1f45RTklf7DEgzT9CYE/AIBTl/5KDikswWoLozjUT5mNod0CTjfaNrEU+UlY65E8hE
Dvq8joMhAEUIoUo6HrcOxK0mR1sBtysN8aAAnz4sSKs0uPqL7u0Se2b9fN61TKrf5r0ICEOIf7OX
/Toh3eg8/PDkqUjh/TstbmdudFLNodl3lXNNWG7Yh0ObrFylYiEFDcj6EmEAA2a+FtaIJRojC+nj
MDnDiW7v/NuvhoO9OvlcvyHHITS8s2QRf4Ud4cSmpxdo+dkqQ6dcnsVnSqyuMDDQFk+sg0jfNajQ
WxkkblHQHBY6zGe2zARuQ/0cjhp5ki6cu9pCCgGNHKIs6QtmRv95w0/gu6cdEK8+xRB14Jzle6O4
f5F12ADUsKyEjAjnhLdBtjAgAvXP4lo+KWNQRsD1ZVWemFnram8nLxDPQM9uNSO+0H/Pv969FQSl
30zzeg8w1fRDusjma4suYxoWSMAuW+ePo5F9HGhNcCCRjBza6Nmg+SF4uwtEXVZ4zxS5i9FvXG1n
WjE/uU8aTZzvdCNv/Z0RWfld4pRPcIG03vV5xCOFNtnchlEcX4Zlr7dcrAB8r5ddf3MkJ3f+OuE5
39ffYWZHn1haoEiHBIa2yQ1kQay33OkbHcmGbyTSxGbu5KYHF96fzKGZ2lqhmygYbrGikMQHJm86
eL+aSqF2oWe7r7ONIQTvdJ+NRQ2OctiDs0QSK8u4oW1HWHNXuZLv66PmFMRH442Zfy7uuCoMo0i0
BAw9IH+nF/k2DdsoazxakMHkSFmvcXebXUWVGUCiij0YAl82vZ6yHwrkcCWiuMSqI/HvAajPZTnn
CY0rOs1sGRkPnY1uC/YyetaJu053nUmrFy5uERYyVW5emIDwBoTZVrJml3Qq7ZJzkwiqdikTz2SH
gkltLPaLLRT5sfiO5W1Wgbj/SOb5iQ8fStg22ZQYtFbebTsf3vwSGJPhgxotCptnVFWIowIbao3W
Fy26dejSe9gea2Rr54O+kqqmQXxE6sQ6S4gdeDOnOKtNe6iLZvXERx2/ig0R4jUPkqoVKCZQ5zUq
BBX3NHw7degWo+2Jmol6Bu8Kh5wwI58Jwx6m3tffdSLiC0lVYkvgMX3NM0zsxqAHczYfgLpgDYop
hXxavYTUKEK1vUSK+a5QaOrs1Wj+v1s2YvwHeHoexy6CWFIBjwDgEGhQMVjwdwjFdcKnT7obcHS+
N+5DJdazkpyTn4rAbC2pi88fH31iR9SjH8zteCE8xMM85EteIdXeIAJLl6aBlCd4ZjB59iBhr2gJ
r48OeoYMNYq4iSmN7KdTZzMkemfcYrx7PBOOKzFjMl75aW/fCgKUuaBXWPVLOZiPT8kYA9IbZnAc
ax4ZAZIQfF9BgqeXk0hiETEcyb6KaxDs8WlzE6oy8oV9R/tJTsak8brcCZMO2Z9cmg+oidESTS1T
67qXgjq0/nvFjm4hUHXVdausrgkpVs+jtijz6/5Pdczv1eKWM2qEIbh8zpKo9I47GojWUsuyBEro
EDt7bbUL7nTTWAE3t+Jg+B4RSiEoB+uS7sDdvrCuDAlX2XY6+zr/gaqzOt52HIHKSU2nkcE+Ampe
kixr1tU5AZ6usg7NcI90Vr19hxgE44iRQIY8WB/nCz87anODWbLt/M9XlbZxQGxiJ9Fhi8uDiAsE
No1iqIFgK19uwiEH3X0A2GFgmSRigaCw01DOF7DL3HyGd1z3pTIqhsHmKyUeo6zjr2xsvMEpm1tI
TP4SxoWRgUF1oDrpMgFr+snerKkXt7kbd9wXjJ2G1uGZ2HCMJ7zo7KmeYKcwyL8QCCT4Wg/JiBgr
uxOvWLX9TZbDbIWljn2nCkm+/AEcqppKBQfApW+yFqIo1hpd/zCQ3Ye4kHidarwEbh5UDBEFVR4I
uu+AHRol69W3edPBxt4qWvZWrLWfI5ON0zVJU8VNYBqzZLDll+ANgkyJ8R2/VEntIvb8jCVNaFbe
PL0jEZ1jhnAuYH9FyOMIPVwiCVviV6yXdFVBjDjJbWjC2JgQLHwMVhJlSPiACw7BKznfeFcwgEY4
7wx+kAo4zB5t9+2A7Rd7O61JRawwXso1jZgikRzZcmOXo2MWaFouJ7qsYUjO7imAtXU03bsAwVj+
p7Q3lJu8hvTdMUKMbuKOxYA5EHoPpdQu5Fg3PxyQ5+hS5pNaDYTO7jL5xP6B1oVe0o5q7jYJKThq
rPELh8UC7GD8raS1Hzsdx15k/eynBlf9XR9lO0Wwc6Yq/qIPlI1si/86HHDBa5VdbPAL2MhWNDCT
IL4nxyF253QBPVFz+1XAje+LmYsVf34E/ENWNtsyhrTsYpluvA0g826GcvwW4Q06xkYYAbwY9aFA
Phe9mJbj1yb7ps0eVAemJbUqMA5pR/dBrtbyt7pR0fGv1xCb8bwBgpBXMlvKUVytoQOVDnje2bAh
daYMD3e0XikLkoDUPk5QDrkOLR9etybOsUfPAZ9fUFVjk3sPuUtU0NfSArmBzWxdMTjw/gU5IQBT
eHmyWX0th+AR+JxjL5F0o6DKpfrKxJ9WT6Che1IhBDPQB9vmXjuYtbFjFlurzeiR4pDDkVpoVQAh
SFZU5M1rBF8a7wlKbgjaeAOLQQT6gAYSSW/mSiD6oyIOl4bATbgOvxIDvrxedPm/DKSFybpWQaRs
4hut9VjJWQhm7y9LTvYSYkb+9eXg7cW+DkBb8ZuMvTx+Y91Zx9yXVlZjaxLEtd/jjFIXCy+B3fvW
NLiyGL58TVy14T5gxlsIP2RW8UJlY9HfEs1/cbrYgnIDiBsCCHbB4aTooqSOhpbZ+fA3wAJH8v33
M9xT6AD1ns8TCCrwF13BBTkqealhrxIIiA9M94lAGMlFBCIhejClgLQwu2dpGkqoFNRS/teNEv4n
/iWq67eOLaA0KlemHZVHqLFTlnDdO5mWaFQvhbWKqczFJQFDi71Gb958lTQaKMrNRlhvI+Hctkd9
T7kPfRbJRABX550AUN6yuzUG8UK2JwyxSAxANG2P6ZZIZ8CUgEgU/CHAbjv/VQsBMVo8xGzKKzMQ
wgJt39Q3d3gXhXTUg/ef1kKyd/E69+Mc2pqeok2qkmBJnfrXSvoF5JpiOyM0cu0d+McHiCZrCr1w
qxAF2lk9iO1rJIvnbyHiyqw5rHemIaM+CVLz2gD9VoI65mqGpV00mjo6rBI5O99ou9rOofIdcVFi
ptpTcWUzdsSbzEJtoLoGfVgN9gGnrQP4wWiL6UwkskNaPhebSeNl2iL/amfSXg5XVnDp8yX0mrTY
HmPl6Yqxp/ruSTtd6hJaG7MZKPnZ6PnksAhRIbmtUsa1pmWttYGU5urIjmwW5Ea011tpEPWEhVkh
LiovWguhL8+5rHBwnUTu+k9vWg7KKM5jlV6yJxZAVO+D2UvM+fNTAxBx6lcSxtTXvXiv6yexhoZB
ynWjoez2ap3Jw7/cFfSgyrr0PsloO45TkyvrOQsS28s5Ym54ERugVdlOd8h87tiXaJBYuKVbHyQw
s2jq9o8tCmu3JXgL0/WTCQWCon4XcGdqLhGrpSE6t6IxtSGvdDsdKmuY/09UMTVPkPVjM9Tc6gZ9
DGbLLoLX/7fUbl707bwT+AbdDpkHkvrEoQo5rvRmLdv9/QN6YHrf2CSXYE2ee2f5kQDAwjxkR78G
BgeJA9KMzrocRGZSRRXOZbw9PIMdcP/hbFBc1a1jNMMWW1l951ZVIirwv0zc1XSkbh8DirTxh64n
Ue3SHx+isRqT6zkisCMsqOsfltdPo5AjTBQ7R3D6VvpdyZPCPxoKmycXIlfC8jDe+7lAbhjUl9/i
s8m5AfFFGNf4ohe2ilwcQMMRUTpKG2vsnj5pSxgkAOvsRzX1r6TL98ET98WuCWJe20XuQlPFJexH
Z0vkMXEseN7UdUrZIoGfj5iY86nPdbONV8HLnNl9eB+cQd/ZnBkSw44G64lKdSuSPSoX9rVi6JlW
UGTXVn4iHCdbact3QKzJ6cyYwcM243wBfAdp9ZsZQ2wqUwUbXWkgLxdUzYmok135p+Zk29catIpD
VCjZ/L6KPyKzqkDRroxUoqdyLvcoxpDTqc64PzHGDEhoE5r6sEFIKlzlGrcCN/iPiHLIHk2CqOYv
pB7HBl3L3iNAqah/39BidNriaNtzFddGbPFGhiYbXMfG3Xul2mYvBiJzpU/jRB9OqKsrqWTx1Zfw
mvcbegzr1iO9H5PlIg1ThjacaB5VVVHoIqIsti8W+QREpgd8DoeJQOIibpUs8rHboDt/Y7OgSc2B
z+SW6gmItxYzqh7I/58pAmv7pIIp1YrePEBR8WTOhpZXvoqNQdaYteJB2dVXNpBFmXrAp4w8Sd4S
deULKaNYqUdSVcRchUc/W8L3ckrsvmxv/PqQtEpbuG8/1WS0ul/i3BGFGsjbMd7GHBn5Y/QLke0G
qOnjANOtKrlmottTmU8H5Vy3JAn6LVSk393bN6bP9BEoVaR2QrKan5TxhHn3yiMU4sEfutju8ImT
o+UMQxkhFmO4BGTQ8OfAKEaWQ7Pug9AHJU9bBj+7gomN+/qzAGfWOIX1ek8vVUg4mJH7S6rmv0Yr
7xm6Cp7mxH+P2t5JtB5JZ88YagEzNsyy4xd1JzF1mCQG28M+sQb65QXk2s7nMp7B+ox6Lcgqv74U
10tQtg6JW7xNukamnA8cdvL1j/i/8OznKOKC2WrptMpP2k7l1rGBV3w8XmTA2v0b6RhH9jKfEU0w
AVWlPQB2aqe5xGJLiS5YBSFAuxvhaBrlIiWUJFD15BIz32TJWeTkHFalIEKOvW3nW48q2/JCzlb5
zkKcuzkBpnvUg6f3qBs9HhtqD2LGilfvEF/0oGkfhh5KPVjxe9Fb+j7DUMISvNybxn3rhkZZ65Lm
YRAbiFIdc0I+nAAdG5Fyza9Y6uPg1Pm1lf4XIin9ehIQk8tnSYeMxNXRu6hbm6q8aCtU0KRmuj4g
5hJ0IBHfvW9EpEV+X8kcXZ8mNcG6GR7pSkXElFtex2IRoTSx3hdlvaFuG6vfXeSCmAKQVL39Gf47
qGT6HbiBjDwDM+wLbD93dDRSdA3iggp+X9GVRneVfNfFEnm1mC0Cckndh7wVrUVzT4Ub1TNcZacU
tFRZHPAd9f2NphZ74oGgnE55u1stTKNzrQ5u2iRAMJQI4n/k20y66F/c0DoRyzTV7nt2JMus0IeA
K8f25aQ0JCrUCXUABV0+U0W3yaX6mlZ7QMgq8EqqSNlV+thlQAwVyT8fClwFRNdf6wpwlOlQ52Cf
OPyCTt+Gu2MHnqX4uXzYDPoSD6mQSelmN1lDvImrz5sPEuOGc3XMtyraaJB9CjT2WP8Qqq48+KPS
i4nHFIXpL7zwNGugdDBJgUHicIgBq0tsdlPnaC9hgynrCbDM+q9gQ6vKkVRRisxWCt2V3a74uspm
S/xVSd4Q22KHcSIlARnCQWtVKQiqOzbu9/QMrDEy9MIechEKiHHzqplL8n+BT4S75jz/oEtWzeZ1
kz30Ou/g/B823+U9N0AdljiB8TTub8Bo0XWdPwYOuXu7DFTfmg30KnunGPKdJiiPfKXniossiF4R
PgTrD7xMfn27+VPoQQ2gz6zfWuUBy6sdKlLUmBrLFmYzJanoPcRvuXPibuXhUk6wE5OQRYiKyev6
kTeTMWnTGS9TK/XZLGeP0VBN0B+Ko6sIRGQDnZj0CcBz2rGKnrWq4CyTWqY4B4mydd7j1fIR1+1i
PuF8iUoHF4Z4t3mUD2ae37/kfmkPJreG/dkyN1zBhKn1su64wqq+5at77SS6FWVNOi4YW+ttE2/4
1okVnmITJJdZRLnHbQ1epzo0D7bbCUBbVS8i2Xq12Wk+hZR+BH7zS//PgCbnrA7G9QTaZUHKCRbY
Ya9uSRikO2AyVUB6s61VbfT080PqfH0RzQ/GuE6V73kYQ0s9979SU78mqxLoscvRX50NIQ0yvFsT
sp6rUEP9/KHtobeivh5XeH9SvXC9FbyuAnCpJEpxa3GIl0mZdfxuwo/cAsRRS+DXiCfrqnD8S0p6
pU0IkOZV2bszaHVYC6E0GDSaQcpn7y9V81HR6ikG0kwzhfanv5es+DYELFk6g/VMtUgeMq4AJGtO
k85gjNG1oakP68uat5oGjHo2+FGLnWSplWMKJGpRpJvqn+wBgOpZY3xXu2FNEC3CcJV1CAcOGobe
cUu/D8Lkrve0lJSbAFEQlPTZqWiYBwTANZRKs78fj1iKs/JMCKOkyyJpIIaAJbtE1vFK/f0w4hAB
HqFW1a0xQfsSMv1P3AFgoPDKgbrQS/0FDERkqMF8bqSTpqJuQu7S0pAmjn8WCzu/9oFjbRMbN24A
LY9+9MVH7XUZ1HDhAENYs3rhDh1kwMwN2OMh/t8Qdhu2d1xwFcuDqd/VPu4+N41KZKwRu2dV58b8
64SFj+vUDg4G7KlEvDVISFDy03i7GZOWK12j0k3tGRHP7LNH7qCzVg9g4lz+4AeTYncK+m/DbWII
zOv0evjlEBOkQdx71Van3QJdjL1jmS2DFC4bIPK4xp6wCk9lxLWiBOX6OUoqV9yZfZO7VYxgmmdR
Rx+Nl/WtUoO1790OIdTHREZ01EGBBcEKLNMPb0N5JrCvjd4Mac2e8Yc1ZDMtlXUVj2TOo7TGH3qM
5CUjr/rgIIqxe+g4WZTDdUyfuu68o49SdbzmYe8xkX+cXfL9ILH5XAidi2km58CPuZ44i63M8waT
OwrDh4yr2+3fpLjB95e+HtpEl+RiDprYwLuU+1qWlhrJc9fwn0pWgK+HrDbcoYPUD0DIWHt9IKlZ
Ilg/C44yck8qasXezJ1InR5/MES0DCSzdwiK2v/OLlRlAZEw+0415hcEi4CqVF0i5Ta3wM1sObGO
zp/BXgmhiwS3kPkP3ZJLM0hkh6KV4RDoBwta2NIUyAKmOQNO7gy/y292TQX79a/epAI/b4v0rxRX
UUXwF0dnw0zxmLFSsa0eW+gkxpKrCAEm7Q4O5CIshIBVKJgLztI2mkRHnBHgY+As/UqR4vaguSeY
87+9oksu9KcOTNTFAECbv8IGhVJFnbkQFiEfh5bx0FHzjp4+vTe3AScWl8fvfnvq5AC7bG9n1PO6
FoFpuR9dfVnOji/T7PeBNHPdep1JEfmGPwIQGsS//19GmhyKV1WGS9+vCjkM7G8CzUlfdkmsM2s0
VaT80XfJQvD+n8JcXW2O+1oTmXinsB5TKc/3HB0DPfnrSGq3QOqQbAWu6JKi3WVjszNnAJSpOb1j
AlJQ6rIYUsY8qhDsrYw0WyB3QTgqJQS9AMfTx1fqTUFMq0gweIM5vxzFQb7LAjMQX21wofUiFvLv
lFUiANvJO3qnkh6OSPEeCL7ZXR113CdWSGZKXmnCB09OOGEGL8Bd54Qi0RU4AqgU1GD7D0kHZ8mN
z54MHuU20w7ek0rLgDLBoOEvJgCLdpHlkSy5eGvA7yzbxjSFleFpXZLirxIK5+IVvlrbeMq3eNys
tZ8SC5wQ6MOClBTI7yloI/d88XcEPO5LA6l5G5/7NQSMBeE6hBY8phCIBkb2fmefAhKVTwNL56MG
1tUCm4C2yZ8MLgbqru9HkA1BU1+EZeT1/hhrNqD1f2mauHWL4PO3wy6RTYNejR2mv+pqAcUtFS/l
vPcX2hC5MXGRsl2DWYwKGWpHTZ8krnWjYjl3/9XdPj6whRYVIxm8REnMKIUOpNZayjzVi4YGzckE
bvGClgIMc1AIkEZADWLBJHUBziV0BCxwxUIc9i/4oH44Ce/cVpBu2CEr7qIuNVw27et+KDhJcNML
g7tQ4oYqo8eJddpm4+Ksvpr3ev67EcvVrEdGLnKXnAdpQhD2vianL3YeG7EJ5cnSG4Cwm5nBrnUT
nk+kOxQO9qzS/6rdqrCPGC4sHIwn5CvnDc/lMx0hdEfT2IMYau0D4Yr61K7KnxAP6dhUKi5ruDGP
BSdb4NJGAvwKEVdHtc9OUA5h1tfd+8kJeQBssHdHJn/p9aDuZodu08U1jsai9NBaR3r24xfZN8IQ
aXx8sYuIbgOzYqDOARMvH1DQuU/ktL7faEpT6mRnSBgNTCP9d2jeBSg7E9bIUEFfQfcY+PmRiHg9
HNHfwfGgR+CIS1SATEhw38SOdu6wUPpC7dABqRMLMtZBvWb549P4Tx71MPeAjrTkTphtggJ3q4bu
dPdtx1wUfXHvcoWInWUrpLcwQ998kEX8xmcvytJYzowoKf9lOjdMcU3gdhCyYAx2OMGGc1Sw/gem
JEsOQzEECacjJ4ZpiGUkU6lelDUFTmmP79UhTefM+ZttEm1wIoFTRN0rzfJphVr0bGNk/aqOcrYR
/zAU8c9KXeO3ju+Np+GwmZFqVSRWQOclBXDE97kxLTcy4nnBGCG1WYTgigzqzUTUTyQBDsjrDXbF
kk9+/4ZPFdSw5jTT6iwEB3k5a4W6rLXO5gzAvH0YRhjR60/t8El5iYshZw7NkuoDlTPnS3wr2/bR
v16imgwJrr56aAj4CoI85bwD5YTUb4+VEojMK61nojjy1/bfPARQ2pDo/UN4hSwC6qFRVNDj1O84
2vKk22gj0AZEqosOdc7YShRDHged1gr0MIclUXvjbyPfqn0jTXaxtC9p+Uygpbo9BNsJgYaf8F3N
sXHseGPhxq1KhpAEqAnNjNurwozZEEpzcWQakfz5TAr1e/lZgkv8uSdf5DlizXxauEPX7VqrMhFQ
nNF5dvls90Fjaru6ThT9FqB3dE7N0PfiEIGBTukAvENo1dUPtlG4d06mFX0EGLw4zC/pXl9TGZ9f
3x9j+iEJJQhnLw+5O2X7k3BecGtKVWJec7NMmOLUr50w6T7OyXIahg7w7RmfBUdlfh3ZdjtHSBN2
I1xCp4s7q1lsWBdL+JdEcc67yyEusL1trj4dFJSeOyVpV9W5VjBbV8zoiDTyaQQ6pDqS6LZczfyK
C/o6H/PEiDVOknqbuQkDUARcG+ANzvmLwsbS1ta3iH/hkPZUOMkPeM/71pPOZFHtkk6lgu/cwewh
7hIiKsCkdaK+L6S/M908pfPox8y6j5ULEVJdG/UMIextnEHQAB+ZmYtrL9RDR4OhrO9HE5RQa+id
DXuMwTtF0JcVUU7q3cvsy+Sj4cTm8Hnc3JKFmpHu4tDlJvLqHtm8kN8+jljC4q/RMUWG6lnA+VHH
SylYamL9c/jD/t77w63A+jgQjHlT3BEtqTEli4Ek6W/AXD/FadpRLnzM/hCKEPdIE71o1+dPGSeb
kYv9D4sEn7SfpfNEVyKkliDw1BGboZl1adEjlTYziLdxVrpPVMT3wGBaQqrnhmXFXdy/aimNxw+7
Gn7NuFbQ6hCvecj2s0BoUSgpULOHAo2z2urQyW2V18jd9PVRc2u7rzbLxJQSPd20n/V9go/pGluR
b9KX6OZArhkntl6qVkdP2RJliKeyuvbRfkLLuwOEERFFVVsM3pDIIqAUZnTga9z+rdTYhJ1tnvzX
0FGycqBytNXoqwqTkjlI5hjbDb4yFBhU1nmFACJCBF8VD3aV8zXZ0IZZvuhCBHmnKSY5Q0Mm+Ra2
zhNdcuSTSgR4U8WOtdoCd9i+LSaraWFCM6rwpgwGOxE+lhhh+zAc7RLFjC1n07Zfjn6e7vfuRKtR
KHGwnjdQQWtAk57QpCUC0r7LPrFG2RVEUIBkF3G89FwVNn0t05hhjVsZT5MVZxwh+/YYvh6//Z4H
cb9SZHfWWwucLzUj8PagjMQc9qxC195fiL6Aj2ieBvGgtpvjuFTsMCRiDAeSbAUuE1VWss2OjHki
9OdNoQFo2buIzgSeyJGsZW8fmoLI4Hv8omiFYwq05gzczULbTEvelr1Zi3flOkuSUpPeEzGtaKnp
5OdS+7Zx4XAOSbGiPvNXpvsJxzJM7LyOO3HWQgzSIRtVqKlYHu7/Q/v0/OGFPgLKCNA6igm//P8d
OXy6sKUAVSi1bQDWSgXaqsI5CjiaaQRHtDioUzLNwZcsh1nQrnJoaZ2eAN/0CykEUw9wFwkOiyT4
7j0oJ3i4CqkbSQMXZxrv/RiwJ0dajXYFUr8Q8fB3rKCbZ77qHm5FobGmrpygqruU+6KstG3r9kJb
tCeCny/n0f+jOfZ+W5C4lfI1sj8wSqlT4kU5GVFpvPqCehjz8BFh1Z7nxSnYNT8VrIy6SWx53Xdz
RZF21QPtZzqVt0lAa28voPLA3dA0dtGD1BPYfhGkgq6cky9TZuq+yVr8G5i4dH8/BBJmlEAQlePB
eKWeTQUJOVNnYo2vfY/DW48kQrhra4b43W7Jm9lEZvpI87chlWK82pvxoCpqXQO1IDZ9q3WRsVKX
AV/0V+00XueqmSv92n+WEJ3amRAfU5nuQ4XOPoABWEQb3Yr+wgHri5PCfRIEDXsaMD9f6+kAqXXf
ZL2jeKJRO3RO2cln/6z6vX5oJ9nVsUImLNOrMqLnYkls9zlLm6sRgCC+O26zBlsSFAtc9xggL67m
0p9EoXJGRANCimlSYhpuhlsxopFxyHG76ZViWi2knS0lsnlUOBHGuDq3lWr6FiOQxGjOtdr2IaJC
4Yb/CrifZU5LdEHaastNRkCzOvfkeQgZ+e5TItyys/j91cN86mFOslezR3rZMAaG3KlEXT5BWFhm
mmAsd2J85pZCRlSFETw8gaTKIyNaj/jnS6arJ1dZY23tHBFroxZRj8aG++UvoK753gcmYZAjZLoo
x2MZ/HHdk1FgBg+yERx8Lp6uPmTwR7IROV6Q9ZrXB7WZlbf9AosQLSLDOmH0X7I4shAHBH9FOE3F
jjAyGy69UsRTT1vN3UK7tCbKz49eiBHQHSBEfTRCCwh6zkupwxus0hacj/KzqLOVK/lS59M07Zfj
GiT+POyf//cqHU+Q8Ov7ElAKSzNEPfMIXfqXkditSTz+y56E+FCU0l47dE4hDRpDKD0OGoccJMLJ
iqJJAm0znr/786YyoWl2Q2temKsTCru5qAJtBy41XZK2RZv8KxI+QHchhM7OzMavEFiHFay96r2T
7TxwHUfAxvnpcyBNL8Daxci65RKVLeXd+1hZaXkhFNsF6sr8vNnHrUyX24G6mAzRhZSnYt1KCmr0
nh7JIodK5Ag0BK+igt2UKrLU4+lPkMOZ92J5AP6jQiX3Phv/3My1A38tGM83HWmG9QLiCZEvjl6u
Ve0lhgz8W0MpALmQpPuIlVRqt5opE+0jKP1QdOdrUECnfgaz9+KHPCO1Rt0bc0S9ljNdWYQ6ugX4
pvX1RPkRQSYyYWDpc9dnGoy1MLBzr6DziYEOM5dRRwbWvhfQv7AsksS/a7wBaQdx14RHGuzKYdl1
tQGes/AmLxr6GQU4WDs4Or3RQ1teGEHviglZaanSixqtgB/C2mraO3yBzbwgdMlCdPRroQeT1Xir
X+3ydec3J1mw5lEJv1DeDS1/VlTac/2z5i4zkuhJOlBHvnIjwFaOZqSCNHVIf941oFmpuYOoL97k
aBGq9V90pZg/+3uGtsRcA4n4ldo8nQvUZq4mg3oClItTxffgRGGgjJJuADyVz6Ge6uVXTrQRy8BN
pEhTIkphlyVNR3zjYmuRUO9745vKLjtbOOCYvMAtGCf5PQDwqfFp8unZVrgeFG26wzBj/SiYl4Aj
VAEWBny9MzsT59c6K4oo2vuXIIHPu4s2yY6i8BW3Cs5mwDD0BAC0m1L2dTeMPiYM13LyYGpWyhCu
ekblp8HSAHTj9+DrIPv5LZ2dR0GZxqoizqELjkxSFwzlpnT63wi0iH1YYgc7U+JRwe2ioVk/asrJ
vIwYzOYOFiPRHzreqBwK0Zt65IUVpySgQLWXEmHt7BzkgpAfzvqXM+4fmcnjS15+xPWTLwRZy2JT
AMkj8rsAKZAUF7VI9juCgi2YCjzxeUdIvRtCi13ggkUgDKlOLcCV9fHtYyXJDjPm3C+J//sShH7G
0Tf7ISVQQMd2jq2wHrXorRhMxGi2JTZGho8WhJt2J2QKzHYhvWS9c3WTdOp3mD1igxa9ojhX4bW1
YgKG4gXI6hTfB6NRvbmqsQk1FvRODlTCAyOet6cl4WY97YNioqI4zyVGBmocxmyu+7eghLiWSwNN
Riyopl/+SEkZBkOAjC96HiGhUaNq1iFY8/e9aDqWykrwZe/2yK2NtrhwxFe72S9/HGHmzisznGC5
95PjUmOZnvqwA4uIuKE81spHTizZuPzBTvwHOP0soL0AtmAI78dZOhPw+LDDLLJ2p0Pbe9pklNcK
yItZsfVYoQcJgNKuVV1ypxnubhYYqlAoqpNamSFRQ8NFjcZdAglpiHJYQN9n2s6A8p4Svz1lMWCO
Y5CnaegMdH5XgfUUJeMs9yzTQHyi7KzYPy5VC8MdcF7AMJ269Ly5vBGzJ1GyaWCke9XtjKGCz7wB
P81OUqWEngnmhAtl/s+tKI75wAjle7/xC232kSUZXPe97K9nrNT/R7xxj13EVNitk8O3C6KskVW8
H2jAQSNYJ5j8lOSbUPqY6KbJ40I2YVrC14AmOu4bWsFvf3p22J8v4MNQCif975/Ooxtk0AmXJQUF
L2JXYJC567Ri0X06O2s+MF+5GMmxeaLfNvtoGtD25+yD2AGA90ilalx+PvZEff3K50jVYFZSRz1N
aCFmwNXLRLyOPH6Yvuv+mScY7sA2gBtkJyEx6j6TcUOt5upEMc7axGfEN4M2W/KV/XoHV6680W9N
X59jpx1CZNxpRqCtKqSr7bUC7D6g+WrkVTsGY6QQREsmpi66i9/CsAakj1r85eprNs3Cp2ETCOX0
CbaOtMr9B2qzILbbyBGp7y0rz330FrhuEySSND5rd93IvI60fKG/2guFi0w0tS8qay1UwkCs2YIv
6dnpj/9vuMtkqnia+nUTFw0w5n6jrNMqOubu9eo/GeUwbWCM4Q8+81Sbt1eAcQbdpjvaKwHFxhfH
H04kxG1RYHhDh+9VMv9/RBTQD7QQoiF8ouioxlxbdACo2nz5Yx8E/ANs1dogJwqhxNkZuAKEwEyr
9iraodOENQW08zbEosyNyGnv/6PoYCd3Kw1EKb1EJ4nYTbTU1eokqw3BL9S8yic1gFum+nklzOXa
76REuk3orhL0lBzPvWiBw3pv5A7bJ1bsa4xCc3VMWLi2qixUn9/bA1y6oZxg4YPonaBdem2Xbe+U
+TzD+X81vJFzy1bTezgTqxCuoAuOO4E1D/ojfILvh4ziooEDksS1XjBBl+GBZHpDFyYbY/glbPPt
tPGAwwqjPnJafqLjnegtqPQ/6UOq/KwIK2rvH4jnyoKKROCNtRfswQOamKESMvDhT8PZ+eo4a8ON
T2EG47t/yEB6N09tiU+BpK53GMO4XwY+6d9l5AwO9cGSS7nQx6tUAoeBQSnbzdyQcoV5u+UN6wEJ
eUXZb9NKmEnuQS5BOfVm6Tpe1FOtZSHBAbbC8LnO3vzXyd0SCXgC3gjO7+kh4BETtVN0KsjOrJ7D
Idi3n0yq+/2MHkJRVO+OvEFArGD+53igMejFgzO7OOcoa3OpA9aQx+9C3cA0cFSsQ74AReLqiXlI
061ExnF7QDt6ox8a9fkqhfhIUXeSHgM44PLavs5sjzLF7ZGHeSrxg9GXf0TcukR3QgWlfRHwJgTl
4MA5gz5VVZL98ammtOnDzR8kQkYpDw7N6f4MULEweYzvGs5Iqj79EumbiGV2aMPPFFYXSs9BsJrd
QqEimAkouHcHLAI4cdeuNJZQH+XmhNU8u24rnRRNX6eT/LwC3+aheGX7HMwri9R4O9Px7d+X99Ha
/jLZvAoD6hbWckpGbKx5kyL3IRoneGufUQmlSmfbwjxcno7hK1QJyZ2tnQfQWVNg5Zg92ogMaByK
8PgOVkKtiNotxkJiLD2JD/zuTlqKC30SjvC7Fn0MqfW8N5Y72WZ02nEcHVRLzBrGgL7+fVjDiANo
tyixnOKXxHryf5an4ygN4A8Y/4PT/CBQmnBXV05jdTd53E3Pi8wivwwvYT9jZ6E+QHewTtvo3AW1
vNmzQovOjGb+MWZdIn7I/Vi2gRlfbJ21g/b3kZ0PyhB7J2BDthF9NfjtvDHRfMesgRD9UOM/gy5N
7zVla0c01mB63VjlaOKfuOhLPyYm45R8JRN/AL9HvbLRaGwixN2IPkUUUF45E9Egwc9DDoCCLH72
UTIB5pgshXQ8JpnVPvVBuhJg9H3wSxxBedLzp8iB8dzqVc++iF9HiwB7TbcXrbKYVjoIn4oyJlCY
A2BWvtVZ8pFmh20hNl5ruhT9mIu/mnEJFk5TstNasTl03M5DmEbKs6+fagWIF1kExK56zdTzPTEH
0geSMW6uR1m80rrTpq3NEF90L3PMa1xLvq6fHePYR8OtaKwLwOA50ono+GPVDneFN1gUYXCyTtb8
6yEt+FEuQbQzzdQtQtUYj+LXkOVehG1zLTPf1LH8zoCus55nVT8ic0hFxlHb+eLEMl9voLw+/ytK
walIq0YN7JKCXrVwJfBmDD038FSSd0gfLoGHEwA8qVrDwX0ZOZ2bl9XdXX4dosnqZxZxHF/AfE4E
rSfQ5HJcQwkr1Cru4HIve3OdnxbZv4nFEy1JChoPA91BdxzmBSPmOZPwppBQ0i0z/iM9Vkxuii5b
Wnr+XMu/kGbz0aOc+b69Fiv1217XBfb6oiTSKFDfFRa0B2Qf9nHLMU+T4Mc6CSuSyrMhCxitvz4D
pa7rkeWxo1ItXSMzDMUh8+gwICSj2NGG0OZiNYEvNXkc0Ea0T6nzZMwbQEp3vEEPdVuVtD3koO4v
eYMzwyd7GMa6PpxwC0PFt8mGvbuPjQ4pKqteIIz4hND4p12DiEyNCVFr6DEFTNjkhgj0wF4pX/C5
mIX12yiCyFUgDf9Ro02QZEtgy1iB2bzB/Sfmywn4U6FVr/NA4F5F9GQEi76ao0uc3WFR33cbxdhE
U84y3KMf1r7jgm3pUXBRcXzFZA7viHTcXduAIEO/7KV19+3UAvgiKqctkCFzCopSr04AaSinjzDF
A/Upf1A1uqqATqxqUH+wNaQjd1bfo8ex74+aYZb9WUMijOZjV2rZZYR5nDkgKWI96uQNnJLILozd
39P+ERTfCo/iTEBi1b3qcU1ZtTmhrBeK4A0VsNiVvpH0+EfmL7Dh+2CCNeKBmWjMnk3UfRpDsyHl
BgMtmjEstaLVw7tu2irI8kb6jURYhMApEDL5DQ1km+r67/nkxJG3I7oRYZeUac6tVLSKAir95H8T
gIAHYH+mXIJLt0ro49SgYQDHdBx5uXz0L4QtbpVuz9xUw0vU/hiHgpq3CKlYle8rFCmX+GS9Ue4N
Nsh0FM1XcQjYJeZstrApkIUIk/xFL/nmFtyhlUcWa4GuqTu18oYEOWwOSIwDGp+CB0TUVtM3dVFl
YWtsuvHP+GAybrCojlHHnQ8SVt5xD664CNH8yltWh+9b6YP+4GL64ADS6enmHNaf2u9aSkMImiM2
ZCKSfctxzz4+l2WvqJE79DM55JZ7aH9BUSR+nP2dPRwwlhAWDtutLQJcHpsYNJpeoHgoNLyNFdhX
5hkGw8AVNWzF8jOYCHBZl2jgyL9YYWkS6YDPvGWwtnoipaAqzydKENg9Dl2NnifC5W3hBJszzMDB
AILr31R7RE8VPkAfUpMmbaVs83dUaRn+BzvbdeEhmcW0D4QplYJ+Qq4B/5VymeELJKZH/oKPc30r
LHd8mBaAaIXel4lsJEcTdRK4Gnlf1gmrov1aaLWQ3ZYi6zj7Etgy9paGIM2fcWxJy30yXsmsQ9iF
dJh95gRLvQry8R5jKQFpeXrOV9UyfN5UjVkFtzz0hx0PVxtIIgaUEceba4paPOn/g0cqNsEnehkk
Ccg93i+zoDQu3XIZF4eJmmSt+yR/scyfcFWFMS8Tn20Ity/pZqX8Yd/VazY1eyF5LgKHcytArMsQ
JbYxcdeBDqvo8nj3rLA4+ZD+px8amy0tqd7Z8hglsjghb1gnMcdDSv3HS0+kTTRhW1YQyHndS7vH
C2a6k4QNVRYPF9DGQY5H2pJqeuwM+DAkS6mXplzeoQK7mhHtXvGHqRYQTmlsBkwHbKIKt0UASQAv
yYaUeKJVaEvnIlSCnV+eCnG/OjfRfsV+cMCXMYeuN0TPtnlyj2o7/1BKXK5UEsSXe0wE3NCdZFAB
MdDcic7c9hsn/LIh1vbwFE6HM4Y1gwryUhcFAK+cOBwWNuXAbIhKXAGWzHWC5PXW0i+SE2K5p7ny
NOjSsFK4Vw258ABSNdBAlW+G9JyWS12GyCPZSFL086FIDWGu1jrLy8P038rYcFq27U76Li4G2w55
DVPGYAdd4SDdIEmsE+5xJO2xquKC1wnpH6/9gXIypEJqRDxqQ5W4cKBzP2ic+ygTWKTwIhWjBRCD
stX6ajPk1Yb9or1Vr3vk0vEkchpmZMGC25//nYtoTtg4U2vfZWMCXgKJaFvRtcO3lqMXHGsTlQZl
5B/GkL1NVXS1+GSJzBLToAkKkQtDYwRbj7kfXH0IsLIbt41CWk5X8abVWPiaNRt5QfJZYkYbikhR
RW2g3gF0HRdCQSMuZMHuh7IBY5ntKnRq+VENE0YhWDk26APs50o5XtcK3n807GtzxeRj/ljfVxQK
M53cw0TUQHSOcWVGib9BGD6bB/VMcIvdf3Sx6HBBMUWJOpiWD2s7rhPIAxniKrRWkVY5eSEMWm9r
dQJIxBOqHrOSgUC7WoIGmRuk4s//Wr7JZbToFkU4XM1RqiBm97LfEEzkWGUx9/PgUFpWp931bwPG
20r6fUchWQY/JJ+6cUA4rs0XABhPcnUE3iMHSsZshZV7XEc8rlFKxHO+0dni+2BSf9pllzjXdMJ+
nDMhSaucmCl81sZZcpKX+ZgP/oU2wfFEE+ZF3EzvixS0/rvO/fBwgNL2w9yTCLM+R08SatV7+0U3
0jbdGoKl32WWt7RbFQ8UMP33UoUyOoLEi6C4r2/lkNvuF4ethjjjhL1x4WuRjjxxQDfTuACj8Aje
JmfguWTy7zYMeM+1WowGoQLpfmCScxj99/7R0o7DHfjcCE/eTIq3frs7cYIYJx4kOi8y4VwMN65V
VIVkGTRB8GDJfS2Q2ZOj1G4Agr9YsuMiV2TRtLOuhR2/6GdcCjCPS40e4UPuLoBNmIKAAEC27AhR
+Sp8GwBr0YJndyUf/N2JFKLLatuDCMPtsbXXZeGjOV5J1h3IkCbwQRnK/wYYaRRKPy3+ADfrnWVk
fANvUmANbNYodZQRuPxHjWZv0he85YGSrDgwys2P6od54PItCepJTqWMwq+t3XUC7sWJJ6htOF9L
f6Dpu5dRs6XGGlyIWWs2PxuPRn0oq6jBAst373Htaf9nvktNKEs0d0SBaFz1ZYkXphppTf66dQ9r
8r+xnVygu4dsxgBidJMulAlcInAPAOsQzf4z91he8T+HJLPPQ0Uc6BDVU4WTnI15X+w6ijXPZt0C
DIO50BPMYKSHCcl4CtTO59jSkl7CqSbHjyCJXollg0OHekti7MzpzvTORdLwFeCk2wmrl1eVvmMW
zyxLgfowvwum0d+WrQBbgOyWFv5IWWi/DlF7tA4TpYgikjavPnKAo4XU82SRskwGWPTLZYboC6rI
dVbbq+aJyV1QxreEYfYipOHjcl+aTEPxJIXtHmBQE28wACkT31eSdHTSyayVrQDoVj6oFzGT8u52
OMPCX/lcexB39EgHVAEmgo7YypXOG0CNaeBHmE1XturqxVtlZP7vKIOmktpzwChm2zmQAPUb3IiR
b8CGq7lr8hDbu7k1AaZIrmCb7dj9JSY1jd8eiNN6DeCJz3vU4IV4OgzkFTp1STWRP+0y+YyOY7pJ
21eqwi2CDzYA1G/2qBfUi7qQN3RhqLM9bGpnx3vZk/j7p+Ra8+0smviYOF6oj13N+xGnK+STAUVe
vxbLMt+p2YXaJccatBFljLLSe6DAMYdhJbtQFn9JmX7fu7XIuf9kSNNM6mb0yFsZZkXmR4Bogic6
lWSoHgEtFudtZV6szxkt6DjDW7BeYteM2YsXerUUdazClGdBCvLqjpcOVb64apRa+Zsgia3WWH3g
zYnwWNMVpFWb1gGG/V/G+t+vyu9aAePpLpzbYj59VAepfTS8zA2iFcyEeBFv4t13ySWwXYvtjD8u
1hI4CjzURF/dHm3I0ZnjxGgni+Vpw1GBFV+UcS6Cg41O9oIfqsP2hwhOB7zmH/D5qZ2C883pspAk
KvkbHyWAT1sYEmKuhtqTPo1nbQZlaWherHqikxXsvrJH3IHyFtmmniqGmMlzcMFGCKfrOHaqeVik
YLC9jj1hXq6kZnLga0aprIfTD7zbpJ9lq4mPv87PabXZmlxqskYxLCBqZcg8/lr9XvJMikglLoz4
+A3xVubjn4NWahzQt196IFE/nXwoVMLJ5UeUjPIPUVnfEVYsKFAJ9Fsk272RI5o8BEHhnYz6HNkW
MQM7zqeu/j7tS2I39xHzr79wKPZNV3MqKOjRgZvRA37UA+1DuWzJ7065XAUgguErSaY9Gifmb3Qf
rVPuxUkNoxTo1rYRe42ulzT6wY8ElBTenyPlXc5rFmwRSAemi0kfymShm+l58yoyaCo5Vxn5/M60
XJwCDurA/Mv4rU5HMYqaeNgptuSTAw95M0v3YCQsj17q9X4CTemEeWBxehF9tg25QeKd19wtAvJ+
TqXFp//ot5XXhLQWLJYy/ecKR5eWpUXen2oWo3L+VNHTytm/GpZqrw86NiBC7Iy6yBzlbV2vg/XZ
VA0HzyjJSyU8O20wPWuUkHTwa+0Vm7HG3Kud2jQ8WbqIXXhlVFBPaJg6S6i9b/f4M1sVF91PgYTd
ZI9G94/aD1iiNEY+hUv/hgUxb/w3Pq074503WhEYofGlPWXLvryLZeBSlCMfjH/eIIkmnsZxMOT3
XnbvDUFvoFktVWJXgm1EAcoWXR+YLPOlDsOqC5fTYvegkpxK+W1BEaBTIyfWwaEm3fMWeDZr02qz
iLKxBrhgGLcW2Sg5bGn7Ng6xNZxrWxeuxktiP20N8DzCVzFbNsjH2sa4tgTOPWfliurp4OKjwY0a
XRWLsLY/JuT8hkr+i8PDcXyqanKAtqcRrN2plRcYqqdGk7JJaNtZ7WptmdKYG294GMtIQJu4W6W0
4qB5pVbrEq3QMlZvjLBCZpBzb/UIDgJAnpuTdgsfjLdTlpjNobVI9CjwZF/I6tyCktDkcuYcuCus
mUqsrZsQmpLaFzBmQ6RDwPSIDhfSCEUxUzzaWhPKhms2XO6pYUI/Kx8ZY+vpzT6t6st5SV41VmOa
6llyQdVdVq4s0tyRs8PXZ3P/MdG4ndaSAb2DtDaz5NCfNCYlxzUu2NSggJnosijAHrqgpEkFdsEE
OLYahNgII7gU7aXv/580HXjyaZ8SBSae9VC7gHGb1CIJGEyq2tLX7cRrfMh4EdYgBahGrGviEgML
CvaSz18kmCpndcjUdyAQl9KzcQQPWNqUgjCivD4H6tBSP7F9GWvHGttPf1lDFPy01WBStxZqGcC2
Ruuzzd/pgqVIW9pmd3k6kURkE3a8BA5tM0AP7bmUNtR3ZXIP6wklyzhuK8qvfIGV6GJHVEAQHjWT
OAm+jn3X2AOSOEEAjRgCkD+HOhZnCgqLjC4RAASxWDXiqwSxV4V6Pin3tfWPfcvpwlhxfZf1ti8N
rfzgtieqtmcm71RchG47txkaLjeAcn1tFuG2mz7xA9uOLporysy8fzg2yxFUziyqyHtEY2Vix2Mp
aW1NNuunF+5vZtRIXys7EZPlsDX79go52sr/ODidObBbJJJwzYIvRh71ewxX6OChODfCuuD5uyr+
qRSGS1QdEuokj+VacAPTessZe1YPW7pGG7yyK24AnGGJX580aZ2Ct/8zSR7Lgp35xPRHn4yrwZF4
bv1Z/paSToyqn+kAL/0TxAjIQfrb87I1k17q/tcHtFXATpOID+1cXLOiO+B9FGTbj/LrtKUOyk7B
cAIyFCA+PsbL/Lu/WuPdXQPWONXrYsr8lpptmdoKwJmknnAsDSk2twZ0jEhIzLMrBOp6/2L9CfxS
3RiscGbBhMsdMeu+8tzXAyt9WhM33Zp3Mbbx3utFl46zixJZhtpgT5DKhMPN0q6jty1Kkf1sRXd0
XpddQo+fFN01XL2DM8Qjfb/qMiEQY/FowlhIpKhqfkPBXMuWL397T7PT1wcEN3uZ58G530KvR8nD
huLIrC9J6YU4Nnc1DNfrVnZSDi2d/NXlWZUZN+C47tJJufaihcQyOJ+RlHiGq6CNffxn6/VtkDy2
hN7kNuPBD93Bm4UOnexnIlFUymx0fz4KNHoQObEOgudP/XV+TnVm2s64R4vBlZROmj0HkflTovWd
JuoWfrKt1vD0Er8PaAvRgZFDSlIWhzbrpRxapfILZftpJF7Gz/eYOUFjxUQqpdepXMVV5DGvwdtH
9wVikCQIsaWVNTb1x+jBHoJEkpoedgqcZflDKS5sjcFR4B1hHNJ65OQ9W8l5C4y7yqiFdQiOmGP5
KBsWRsrWkO24k2k4Hc/OZY21sTaiJ+2e0xwiixoFjVWYn3NCQ/U9iZZA8uRIvyq8aQWqtF7C+YgX
PyLkgFjKG4GRfMMF03jp03En5wnC2P0MYMIDbSugLy49WutVYhp4slE1Oh61+7C6VH6g+Ue5nyHo
Ok+rnn3riGkY1dtCRwRnouTsR4rhemSzc83uAyvz20wXwZvu5H45MlCFFAusR18LxkoMdHArc2ce
u1eGjVtFb/qDn+tfsTm8dDMaW3bgTdZPPC/PgIc5Nw7vzDGXfZvMgWzwXx2LNro3888CRGq3/mFl
nB1Nol/3VlJaLwYs0reTyK1RSffqlF/St3SyE4AK/TMfbOou9wgnNptCUYKQk5lC4qidhriLAzrT
hlUO0hqdcieVo0DBmO8D6K6jglTnWO9PKYHBkfShD/zrfaPRrB4GaY/mY2+AdftJFVBSPjYsfQ6t
YTUzX37JJk1vIIVgh3zAR54KSrwWB1J8LQfqwk0FGWQe/D3+7BSqDKRsVLg/xLAJhPC+5Pqf4s4u
t+3tTrFfbnMTuwuciGDKF6jrXPuOnCTMnxY5Y1OwgkVl7obEik5uy6e5+L1MEO6YSst3HOeMBvyd
xZlkrWdNtALGwCEQqqoJXlwbN5uUACEmzJRTB2OI0X/pFyTRoR9uy2TThZk7L4VvAIxaEImaMrPR
K+ItyrW1zuY3Ne5P+onH5WfOUAjlV542QF3HgtocODqc7E1bsLIc53xvJFHluGDAuZ1ReTOszY4Q
XiZjdpCp4Zpa7ZbigKh1BmwCvD8SM0A7P54I4luxl2Q2K9Wgbzv13SrNkA2MDs8CHFaezoZ/j3TY
4fbsw+bupdJrAExn+47sxfiyOwCOo6yUSqEpY1rt2wUSyHGFUW0bavz/cqHiedtvtN8TzJ4B/+CO
qsmPj7ULjMwx9hSXpMmCv18RaocaVQrIDjJQlFKhq2vqq6R+vFkfV+l7t1eLEf8Tb6AmitcC/mRe
AvoTeUhQdwOnTr+nXBDDZGSVGanSTAv16v1OFkSUIFkg7CLkjxGSAbPBA7ndaRT2wBIfdL+lWYpy
tewi0JaMrMJcqzZLMmxdhMsFJerh7F+plPbk2oYzQ+cWPQXxLqyad6Wt2csVhnN8+/ojDEqsnuet
OEvs1w7nj3QZEv6pIJu51f1QV9SNqmt3hP7iXw7vkhwYTMdh299P9P42eX2Mytq/Ps8rj6842wd8
pV9gPSqnL/tMgsROMV4u2NjCkoJFiMJMm+hvVLhGojvT6yjZD7juKq0mQLk3/Rw5x9N9KCd0nHtU
W6E8okb+d+oY7yXKDZXCX91W9IffXBHDELyxwuiQ7U3+SsSZMxQcOQhCcfXPA5mkANKL4HrjIA/y
86dyzn7kJGLyrDKk9K6vXqoD+GqDqyoBcg80tKaLgPrvpTxZJxsp65MikT+/rUYSGNtsN8ODV21s
QQ96PrRuP9LZilIivyzbQyfOSHQsUPmsLdbw+Sm3EXQu0pVM7Bi6eEDYcYUq3dmcLBSIM7ieBGyJ
Tgr3K1qXYTWJ/gxlWsQ16n65uHKvNbRLi9biESbp2BwUhcBAj9t8Eof95F+0lmmDEGGAiT3kM1sf
nWxBztCvuIlE/zJIOWj3cS+rU5iIa6MF/u9BpIAP+TJETjtxG+LMo2PUSQXcBgz+PR1LEK5bcycg
Jl7zHCWxD+KK4dFz2fohF/iXaT9x3cDs28KSIg9mPitdQ9iVJD/MDmEV67fhY2B0H+RSvIcvDdSf
LWstglIPlcsWdoxr1fXmbVPNfJ52lj6a7dtTKNjGxUVejgbpIupR99dPgNrPY86U1DOiV3+LnyiH
3OrVJnqX6Z875GF1P6lTP05Cqj2ryYbFjlj1WFlw8jaCZvuDIoOPZj1ODkwGjPf7fXWlXCrRnMUL
BLxBeh08+701DrWKQOg6h20A0hQRDsrqTjxDUN34FODEfq8o2r0QoB7a1n26tc6wOXJMsIfFodut
9jnicHwy8xICHw1bM/SCFGUBRy5J4HbPtnAiFXrKlHdHnoxrq0vLESsUl0zasj4KlBQUiOaVSFTG
6h7G3FXE1ZGgaiOhciIBBqcAu/fqFVDnkTbGp6Mgh1bSrv7ZceKmYsYSAV1f1/JVbUif68Mz2h3D
jXXNlITYGjkqjll1wcI3PDYevTNE91uUFvdG/Fk1wYqus8TLrUftfD4R06hke1ySLGlm+H9aLzMk
elTfmwy4sF5V+8D9rs8KgcTXhvnU8o7UP5hQmRkeus0jr9GAvT+hL8Gsp1RTv/EcB8QrYvM+2+HA
/rsqsxGUBK9Z9YCkNCyJAYfIxNhXeD+/kBbDreNOYV9OJGhbLE91QOL7gNVaoZrSfZqCcKmkuKCk
9GKXZ8UUqqX138S9G0heIlhuKCHjyt3sl7G8pghYw7kKswaoi5ve0oLR1tp5HEGhhij4BR/0cDxk
2X7D0stLOjxHkwsseFwfaQb3ZW7VOHBrmrzdYsNIe/bbOKfxtpfX+DDCpEkypaY4A49uQuDn68Z3
6aGlqOE1VVpq2mqU37t6rU4ZSYZa5BGf1DCAN9wjMeLKo1V1lPQHoUV+5yLdtALtrX6kMtTSFQ4S
f9c8VJVkoM/z7c8MhkWuKsgBIlyFH8MvgUvtxCxv9XYNbfzjAzJET7ouEy+6k0MO//7tbYzIUM4P
VK8sl+xbG4Yx9RzBfT+9fnClaqFwosDFMJaDO69oHZpyoRK7YJ1ov1QHaRyK+RsffxqsZZsj81ri
dyyjv+kpPafoibx3gx+hKcfzGYV29ipxg01mYfBQpD2UMaKvQzQ6q75NznMSI5dMq/XLip9F59/n
LZ+yYwXVkIdgJhR6QEcaCQPDi80RatnMvtu+/dhmzxBQrDIURzQUPIjteObcRIrn1WvxaIL0ZXxK
/Dw9AIPWpx+4XRpFiPHPYOII9jOnfaVRcUgrdX6W0NM8P2Y4PWSTAEdg6NhE5npBEQBYX0Sqoojn
wybNHdYSdIu/Rs/AxZGGr2RGdBCTbu4BJDgN103zdHp7BDM2yOQjplF9hiZBIYDW2OZTGp1y0gaO
GN7R9W5U3ePBS1jOLj2yqrnbUFxegL7JfNfHowY0+qEsRb/xs030qo7fefXCjh+nWj443U6+VRzt
tYCKp/rWdy5RIkZIrx1VnmDgQbld/e6pjb5SkPNm6eo4pVs7zVyivQ1jE9FYoVVL+KNqVpiisp6E
DdqDwpVRdRF+31WhE6jz2+bIj/Efk8szi0J2FY9hpcNVdG8BmlHdjfTNOG0j/W7yKTSR4CQBBAkL
+Ho/vej3bl3rkMFZ5C9H1AyTDgFvIcdVSRXA8ViT/tbu/xUgYkUUyqXN3pBAbNnOLIA/H2BIV/py
WLx7AcDVQMII3Jse/mqt3ZXW1w+KSTgUY9KiFlZqdc3kjhtyWbDmpKQVzEEXnlTPRmtMR9zOw++O
0fiag5Bhu6kUJ1tk6UVbAWZLN14qVxffjE5rn8p+U/9BYMpyJvxXssPPEGHA3AmnnFa7XLkzNHH5
ixbCfCOk/gxhaHnRNdL+QQR8+x2srdjDpaSBl+4za7W3+di2ssxefZaujWu0otU1rtgfOlNn/LBn
R5WIRJNCkOD7z15Ve+hdy9rS/9q31/EqGy1MoTp5NZHuY+pfP/vdwlLXx3B4raHss2Ww4/+Fj6Do
SbaXzYmAym7imRDACFQFXg6KFHMwK7lZYYOIh/S5FhPt3Em+hgO/d73z/kqlwW7ITJHW3r8kAYgl
pg7ktLd4/Ne2RyKdmGkkLNMOy13QGulcdiMJ3YF0kcg/ef3JbDGjcmwYQYOSi4ZzN8D63lPc7Iy2
ZBEFVTiYwkkSU9j6llfKev6jFmzzhvt1g/RhozW/cEj5jicyBPTCulJcrvEOVkrbbNf4yELZIC7z
y0mJnTp2aHJspYZVUa8uCJWoOlUiNKhVSZvXXFI/j/AXuGM2LuXLf+NZObc89F7nolMp0+I4Hxeu
xPNQrhVszsp8R5pH0H4t0NmsTDQbH6zhNQxlCI2jPPX88DD3s8GWL+WW5Xdjr0zrs51yZNK8cafy
70F3THdiH3JPbjW7brRhtxZhAyCMY6WCfIE0fAM+3KLcdKUx4ow4BJCAiMh1/GsHbCyEuIkUbzfs
o+y7e8J8CK5fkSVoMxzR9ruNxmUC2O4HRG2WEsuKFczWV2HS5JnV/k84909yGmODSSBLTysXyhgG
BU0XOUzHDhc5ZwdKlZP4K7BaQbRK7I9REmwGK4jHlRFcAfIEXUv7r7+JxhHpDg9wuIUC0lR81aq6
sAa+//H7f1ky76DQfSmKj6T9QJO20H7SOhu/2Ur54qgwCEfC8JMRAeCydVF5OKvvAvCB6CyaEhCh
wp6XOjqfszSzjBZMPtzS3XxLVt+I6XFAOwA6F171j/NT+t5pKcWQAyvX6Hp7WsimI+ENDctuac/C
tpCH+NA+LQjKRHqJ6CRZdt7tNAFmB9ziPlMMUD6iOwHSkG36v6RiCZfIf+KujR+sFoETypBMVC0Y
FXrGxtj21crt50XvIVEwuElRHEcbQsCBFHjwzQSKZRls8sQmtx9tWdhXY50odfR6wt1wki8sM3e8
sPmLBcumlGxj2SqaObQ6mgx5g0RaZzHAonfPNMWA/brtB3JhqUvCUY+WDNnMEdRM79WyLcWDVHPh
BzNkWYo7oYG6e5AGt79xdDG5w/VD+z04t6JRqzQEEGPABu4ynXUytcnbYfG0dL31kaE3hkt6nEO5
cPuOERKHSdz5bIDrysI9xQlI3VSJ+5X+M3GvO5sT6XVUGkPLunZGGB2leWa2jjNvE4JT1OTKx8lo
ElAEnVEgTWFmncnI6KH3n37dX7jBybB6HcofvUADTyyg0qUG7LPt6Ep5PVS5LdZWZ0K0Jqpj2bNs
tBs/Wkpn604fpjUTmnsFRcBouVlbjB4UfAFqRXS23Es62HwZMqUe1t5bMe4wG710AquKcrp9W1vg
/sp+7znC86XZa0Wdc/icuQY0aP/itrApebjZGoJMlzOaGxWRvlXL26lNFuCxXK+7IZ0/93axYPrQ
dyRm7VxzSaL3izm7LqJ7XTgMoJKofHcXPfFhiaKXokPBmE//aYYZveeZ3h3/y48Cu29yWeKl/XzY
pt8pEzq4KQHMK/TebDIDuqZ/KQpAnMviGcew5TTmolsD7iVdgHvjjm3JG81K1wOdCZi8bdmn1hCC
OQNSD4JKIJfh8qQBTdI+a2L54axXcsa5JYhMLFzY8M6TMayvOLGQqPRjfQZ9C3jhSMi37TWpQQQc
V6dtHtx9ybS8Qc5QG0A4Eh6KmRjun3WrLHUb3emdRjT4ftcbuxsduZDfBDdRiESQsR3LX3zhbbMQ
0FoJUVDgOH9DrEQY2dsl1L9tGHtlJq+C+WU5tKI8ixPU9QDgPVBg71wyWiLN6ChnuI3+lvnsm65x
AaIjrsFltA7EUmkCdBAj/VFnDKZqjuBTr9v2zvcnjaf2EGWpQPelYfVSXrPAw+jIAvBDvl7gp398
DeZ7tX7khDqCmutodzLS09mu/U/MJR9MWK5aAACmSVdYebRmrJsvvIwIRzVhSoO/bzSsVz51cVIg
/OFINLtYDAks5AfVMd8vczdJPu4PLggIAywAzxz1KQbaezEn5yr81nC/G8UuudHCeQOWavwlrd/a
bSoE0555TQRjb79GFWpv8cGHXLtai4/Ga8rg4NA9dNfu2UVxWlxh0S02eNzS42dREspOg8nVWf2T
ZrDnbfNoiFAxRmBo7DEt1D1op/IgH6YRuyM+9ptQmFQ0Sl/L21FQSUMR4Qoj9CPv8JPFvv5X5Qhz
hv03ub6nm9JYT0GaMi257quq28ZUn9+nMvI1UooAejztAyQhsnGFoCSctFL3QvH8OegAifMHzV0W
d7sPnGZIGOugBfxOjA5Rndo48gv9SIAqHT/0dWVpZ8lEzwsAz81Rgzs/js2B69AtSvA/Y6WxLSqb
FZMItV6/InzhxHx5aCdDgu5bY4JfTkpKn4NUczG1bpFTgDn0QfgIvG1EJ/9Cd9vN2t/L9gATCmCy
0ioykFsCDMWc2T9oCeKWZIG3knTI/oa5qT4pGlVrbfL/oUmlBQAc0f5ETLoFqVU8hm3FyPKHSOHk
fWU+pkWYCqDVuoA12e74JdMon5TPqnKfMDp4XRK/k6zbcId37K+7Op13AX5eWJlOyfsIoj7KR4/5
QooEJlSstq4dQ21n6CliUCslE5XRbnqxu/MA3o0pW1pwrgET2xt9965ZZRn8Nfh3zgQmPed4mBLl
5FFz+hzbsXjF/P/2TlT0bWGpr+TkH0OKbmFuuyS0LXrZeU63jvVLgrXZPus79uaGvpyMuVWPvP3M
gruHP//i9zkvZ7kzjNphG1W+znt15Bg8pz9mZJmJqnGFs40llq+c3600bkbqPG/ZwnFksaF7KC+l
jpRy1SKwJ2zYducb7CkP5O5MKjF/oh6Ti1Cqmq8TmBDLY7TbT17080v2FHMagQ8MjAWeiMPiSCQd
0Em1EQfxVF+A1PN0LHV0/fGmoJhJa3k+J2WKpSQpIdfYJXSYb/6VcF0R1Xg4KiFf64xaSR9YaFVb
CTSkLwnA2hurifqBUapVbidPQXGfdPqBXy3n5CfhdhVraDoa8YiLGYWQcKgUxqM1XVN6l9sWFs+g
i1enV1qguUhNdHu7AhnK1Wk9EtmiLHlbksYoc0czFBWq5pdOJ7JLcQVLxnMzqfz+sDmNxNenDoiC
PH46rv8VqWwZ48THgZSaATiUQD/cBX7nfHr0TV6gX/Hw86jDNQuaKzf7sGQPMnA6wUjnrXwC/bob
4zd02CgA7047WmCgLy3cs8cwXxtBWF1dNCbJ4VosGZoF6X/x3jcAziIQcBTp+F+BomJXWV8bTa+g
5VjjU1cVlCgtLQ+6eY70xqjd05+MPemIwX1MFxIBdF9APthU4IX7bBuPi9sVIur2llpSi2SHeOAR
lR/trCi2PzdLmbYDirdYRyU/w23QHpnqhvlEUAY2RAZ5twoqHdzE8jVDuTMNnUPBPSIxkS48wwln
67LSxucAtmu6UdQbY9G7g8/d9i1e+3Hy+UzWtNfLPqDeM2NJdXXSarQkOwvtwjeVyaNQiM4rPChw
ZqJSm/bT6/I8lWOXn22/VoOTGBePAxXhF1l4eeQhkWB4ei9VcwTQKLQig0SVU8JxjLV40VRtwVad
neOSgW/pCDwoozjon4GpYqPWBn0//PZjPBvu221cWgWZaDkY1CsINjxLZeJ5+/6iAY8SgGiGrWbp
B6DXxJP0iMuD4xX63K8rf8ItsxKQeO8jFD8bmtcpzesZp8vYfLJ/AeZakshKvUdbAjBDkjBa4bDb
fai030QKfE/ZlsmrPOSwM9UpVgWpQmQG6DiISufnKML7ZXZMiN4+TxZEvnj8+RnH8dg2/wQYEl3n
vuE5I9X90CIFsatvUMNfulcmAKxYtbzzyO/CBr9UELHAq9FY0QV+5nxNrjG6rfDHrbaeywc3Z5Y1
B1d6CO8kXH6PfGxC/0F90NX1p6eadspGPyH4GWU/h/rmhKg4O6IlGj/w4YtAmpLNj7gGrOThGdqn
2F4Zp0o5Yd3Zb82V9gPhehQE/+2ubOb6lA/80fKQgjIQb4/a9Frp+al1zyIbD1guud09+7wWs228
QMjp94T29JYK+OLuefVZf6zFa5xJdGqfdVm5aP5P30f/L8kzr7XOeGLbxzLltv1kSbHSv7jx+Cuq
shiAQsIsnj8BL69bkHRuPudpdM2yS1ZMa34QTdrIzfnSfocPtVHQwegJSmhKkXWCV6b9E8zO9Tte
p7hZT5PmZjTYTvpX1EUFR/yxtfdffISJ895el083alPOKWOw5QSgeMY2iR4ukLc9tvK00MpkLzP0
L6FjGzx2u6FpquOuVB7bIA0dJ35tBdiradXmLT4r+IHMH55SQspPnoEi42kA6RQkyAItSewRkNrw
rH6wD73fwrasAmhkC0A2QsAK1YUl0+G/QsPFWTIxCHvbhEFoFZCkOc9JJQmHIgKOA4xSiOV416u5
ZxcMtmZ20lxgNMQlc2LhB0uRg5xg10Eo1ThE8NHQVxOw3fSiPqEbwFYfDSV1IWpid3Bjw8IxW3OA
Ty2Vu7Z33OmA2M5qrK2MvWZGTYJ/XnwRonturMVCX+AyXFUkA1B5zL4FfOkGRcP8/y8ZYCBxI0Pj
Zn9yUzVKIY0EiZxehtuUPENGDPpXKE5jezYHXFyGqKk7M4KlNuF9k7PFyJAaAMG+jzVmwKGlaVaL
pOlMWcHiCyDy+gPXWBS9ga51IJjXdqUwmle2D0KIWeVmZNwOdbPAGsR2tsfZTcWb/qXGv6pjgwmD
bwo006leL0hocotIhxDpBhhoeg8P5t2IPRjwjDBeogSsXoGGx8/r5WOKLSnf8tWClIitkiLvvvyA
gp3+PmqsrZJ3b40CCPwV9sJhkntEv6EgnRTgMETVUkgTlkCBAxKkDoFI6+V1sFrQlFCKvXhWzmWE
mrknwxKzgLWHAcT0xGEG1rbxFszGDfeUksGLamHju7UlpnDryXIn7fA9Trcubawv58uzk7KpABS7
c01VsN2RYsSk2IHwbnmXaSnY4V51ZlEBZQuDpU4WPQ1QEa820QTwSx/V0OPM2ijFxY4LbGsLa7za
oFbWaouwRgrCh+cRW3magnV0647hQWkEQOhWJ87XQBZmj4LOc6ycOYf/AVP+mzi65iJFYUTWHzhI
uvp2QC78S7pd7t6aHEQjrgWwh74VoT5xLsU1hzwiTFdR0zYAHldVKKxVWxy/KQa5dtXd2BXlBKwE
eZKOTCpvID3zCI8qsPxXdct710MkQ+9U568pPMPXY93jRjXrAL1/a9BKTvfPpKVs6JtGP/pydjSX
t+Nf+wNL9oibp2+QtH9+xzkSZhzJhdp4desmqb/1mM1JwZP+hGwuncEO+LhCQxPADbOxU72YmStv
iz4gNR2T0kaDQPMD98bEsq9ogtSe35in/6RplyX5NHTWf0LRcaO7V1SfbCGo3HZH0L5WWPFdJ5L1
k6pFarsrMYpR4g51O8xiDAc2iqXpaWWfghycNraTR9LIpCrEOf2BldbW/yoKohkqjpDHK/L3rfAH
4Bf0uqszmdosb+CQEaHKt4Zh6OGJVxz6BeBPe0bQfRNVvUlNVH1xzEoMFZa4+KtXSWb2xCQuBYWF
n8tf3uDuP3I1/KQHS9QbY/58o2QltxFny+95KttJ7pT6ppHoYOPll3oDZ3TvI0RNkQ3pjCW5k6E8
Qfk26UlxffoRhut/UG0aZ+WrtdhvF6r4M0KQ80OA7B8IL9kkcDVCVNZ9E/gIPXDGxh3Fuj58e+c/
g6G/H4bsLQwgQDzH3AALk/wrtORwY3HPgMG8itTcAdEh1UejQpybDyPj6QkhjsHqem4Abg+gC3+R
2NzLnN6SOgRts0b1QQwrN9I59drBm4NlnjOP09Ft7fu6Zz1gbSt9O/7D74qLkH2RWeUnGmxJjlEO
tqlpH0zMOjBtMAMbiGD3Ek8vh11gaDY9fZ/M2wMRBGMf8k4l78AprcC9mBjK7xZ6T13qOvq8tE82
LxYONkFLS2FrMyotzfyYsCxNgMNNCFjpTbV9vfDFd8VF/Iy4d4spwACl+JgvwiTq0CT3mQ0qtrLt
G6QUdKp2FX4Nb2xo++3sk4i1IVDCmMiWElSm63wCNFNErG4RbWB2annCMNwWiExBPjL3MzDMQRVT
tQVmc27TrU01aua5aMi0R1hIDkJN+DM0FBjM+9aRhfqg7wXo7Gh1GRr5LdzvbSbmKBywlUJRRfZb
/B+R1xMWdzsoxIMFUv8q6JAvycPDRsvISCrzKD7gR9CKbpG38pA8DGxKJkl5yhguDNu9BqZLGMhn
Qppfd6+qtRZdqBs1iqyUlJAg9BtL3cBlC3RDWX6FhKwwa1gXGqdFyMykChXdJqdznx/sAEcqxFiB
4JYs2erHKT1nzbdD/Lf28dX6wmgIgxxGw1xV70p8vT+z/caeu8EIsssHB7YsIpkHphyrQLSomjF9
bDF0PocDBifQAZ65pTafH37+OSsGPIrNSO+mrRuIppBk39IlB7T2xGOqFXZxXnMI+r2Px+OC50sE
Vb2JCVwJ71x4pK3t59jXoAMeohCFPrW0ME6P6zhwbP7hJO+f9oukgtTyWucq9mDC5JBdLnODgYWl
FjHmPKIjHfA4fEe1nMSFIamJUqluVBtSwGOQk31geOzr9IF6mNf2VPFxa5C9wErrmfsl5wXewSdp
ZNAgIjnfAq+Qe1ebvT8q4VLIBmdywpJ/30I+GTIzSFXEMjLT0E7ojzToB6a4DvtvdGNwfw6kNYa7
n+TvnQkpGGs+ZtVqnJ1duQZC4SRvT8s5rBqEOZVbK4sonDltsoTZ+bY+WLZPlEsYCLLZmVlo7Mlw
hfiGXSIQM42s1KWYe6mOFV3fbhxWR/rFLZk9c5Ungyz0A58Pbek05sRvZZQxRo0mzYN1+UOGIru+
CFjG6OURa9IbYaIdm/5GBUxxuXk+2tZbAxI7ibaRMsKedU/cp54vTJNMEkRQfENP6vjEM5NmNAgd
2y9VJWX9cVVwM9BCclKn0tRbiPpb9CBPoRsRc5R/C6NBZ14vfdwFb7aGp6ZalA2orpYMm98RfrPJ
4h5xUCA8Z/6RLhSwy+Cnk6I3K168ZbI6J3pMHV75NaNPtoxTc5fY+Fn2slCeT1sZfd3byg6u34U7
VGypHhANCmN2cSs9Hu6E1IHEu6DcIco4z8ZtXQ13IcpWIoTU3N03vSVJYmOSToLM/9LWx37a3jzz
Au/HIzpe1+bVpDsB+IgX9DlGdQeTCxFdbJxLgg09PaUeuC1k00sbTQSzGyitbpKk77YBVMcaC8yR
oQ/wpte/WKKGHgYiiGcs1OJgj5EFG5sKImeBbPWxniWA8hB9HWkt6u26YjjaPdqultZ3Phw5X70S
EHPgV81JmoC+7rJsD9NRpIssYslBBMbHb0+pm60WjkfB4AXvxcvupqrFGRU6cN0dN5/dMnbIjKWT
j3FdRZbaKh0LB94iOTDod165uEqp0GYpF//J79G5GjTe7hknotj5tGYpHT1lL+bS5KOo4FpzVMlw
nlSwKnEKzAV+jBh7kMH8AsWZJTIpLnQp7GhfXlIUCQfSigTn89uD/613jAVVelcsJCdNVE1YvQt5
l7P/AFOaxdbot65W21wItK9hTYQcSQHNXnEUydUxcXl/HHN2H+1Z7TkQ15zk2UadNt60LFOEC0NE
R2929SfcpjL+Hl8SCz1WnMqnVcOgPr0X43WKlGiz8FVKIhJoJo7kmqUsNuGpMoHXKiqFGPAK8vRk
z5u4z+GuvJvvSXehT/wqRpLQWnEmbHv1q7yy4PujEU8lDOj5KCfMBJhtBIJY0uKNSNvrcO7lC4Ci
wuPKK74hMCXRc/Q5+FachbY/HCSKnOiiftGZ0q2Fg97Ijqdq2aN5yp0vF7FHJoCfIKN1E5B9yprj
/L5L1P7XBlWy9XPMPUM4mwSz/FWiqXXsKUk5+3ewW4Q3chnKkyNceTn5iLRuSioJWLJFFMog7d+5
UI4BsAj5lYN2tYjmlYYvAYTnK6qbnJZEf4SJCW7DwMA6tqG5QyeNdaSuWATOcNZdDSPo9j196jMs
XkRGI8e7FcHqUWCByMqFoWATbwq7lns2mOcZ5Jej4EnoQMTpIlZtKgL5Lr2Fxq+Yy6N4dNAFm/rz
gbscyh5cRNXKxZDw5nY95t/E4hiUKlNQi53n0LPeZbUtcCQmz7E4nPrx85kx68RVYOl1FNMmwMZE
8V19UEyPdCLUcuWLPko3x8mk2UqZExmZEXMBfJfnIKiwBof6TDGgpxH98ZpDNR//tP7wTP5+UY8o
aOYPMF7sTokbSJvGkC/2lmWEf+W8aUQDqi5VPuqi/Qm2XCSFKl0fqP5z08ro3bld3oiqIZUojYQ9
OTNkBwGn1P/9bhLaCQJS2ydV/KAUzFnU/qCUUahZ8kxdW/1u6HJB5u6QPoda5Jslh2HpqWAns22M
Dwa48Kr4vIt+wj2DkCq6ooFqesMoKEuVI5ItC+IbWnzTp8M3hg6Pq9L1zrjJSf0xVJj0NHlK9e8t
fFXLu0q0XIIjeNVgK64gqwNrfB6Y42z3QDX4BJOkO+BIR2NBD03ryP034cSgL+hH7k4/wQGkkwCJ
9Nv5lG/zZTCvIAjj5qz7iVjKOEVOxoUyMu3VYuibf231I/Y4XjZMpngfN8WamaHQrx62ZqCzDbiT
sxiD6Qyrev0X3JCG0Uhc3BL87bV2q8sTtbsXskla4lnm2k8F13gaADtza4WZxlfwbiRE3GwRYwlA
KouRBdIckBbxsczZQ7SGaUDNK7ekIrjT3DHoC3CKOmAq5rLc5NKQTHHHqpJ9U2+pVkPSNehaAqMD
2J7O00hWxaMc6bu4ezkRwDLeNb3w04sg2N7SZ9KX641mxYOLaP9ujZinbvWrjA7PZocl/WDDX2zP
3Rd/6xekU/Lai4rWDthmEWuDWSgM/lqkdGTG89odd0i9vFC1JKs7gAtfD7d7VRrBBGM4TlScVmhb
8DYHF7pp3CI6nst/3dFCIlc3FNUtCyJrDgOzs9eqadgis2pziVtx3k3j0KJRLOXgr3c8fFKJyz6y
BqpY9QeQK1fNl74vYlJKc1OJQhZAXUH3FXMRxBdSu/0c8JtcFd0jeXip96921BTS5HHZ/lZqrkZw
YOwXMxr7ngCeyw5ui5HzooBr3uChlvQepBrcGvNfkbH3hdhzMUMIAYpAzY9U5akIfvH5/p3h3jY4
RKwI2XavjPTTdrZ40ysSvK0wWvffJcVwcW0JmvZCU8foFhg8zR3EBjnaMGJfeaDU+1KjfUNGizh5
7rH0XFavx0ppHlpqXtpQouy7FOU+Gwt77gvtgKzXpJp8uWBwoTi9iduEH6+c5imqNstaUzwniXcr
/6ZF8VnB2pC9gVrmu0B1f7N2gElFs1LmS42RttwrLQ1ESOS4HjWI1W1/yI2urEdMfMyI3CuS7DxE
hNMJxg/OTHotQ4UxW14VYXD98wXMgpQBd7kROxkwxJyi6WRWL3LBS2omPCCfyV36h6/uiSknar7A
Pc+oNsBnlkDyeUBkMvI2cPlSu3UM4A/5u7XXO5sLcdjz2zQwgNkZo5OX3E/LtXKLqlXB9sMR6ibT
TDZrCF3Ij/1TynAnQroL+DU2vlGKN6BqpM5oPj5Gepp8MHbX2GSvnE0fOEaMFHwiiouZ6ubkTwwb
7FcaPnhZIUZQqmv3YV39hlkot2bYwW8u7HU7qtUONMEQpMYWGDjl2x2vcaHA9qGNeu1nDOp87j/c
sKde9fnRz33BlZQ7tmx5KTiAjkmE7TLmcEVm+523bIhtcZoTCKLJfU+Tx1BPXZkNY7V78SM5zQjU
nMErYweeni4v3FK3u4uYtjOMMPVMsk3+UPMSy2XbQMe0hejqlEorI7aGMmulsfXoRY4iyL3+CfbM
FWQINhYeIwL5vW4t28XXW6CZi+XgHrlRKr3bfGX/iApryejkRPl0xeFawin302nLiMqmXamCjSfu
oGEilNbhSQVv5hQtWK+6+en6a7ybl1+j0zgUK4namw1mGjE4tgjknJ3Zt1Rx3hKEXeWJHoT0LQqe
zN0rhVw8htrAnXsdjqzkS/4NqZ7B82d8cR8VPgxBKoFy5nNwVks8XE2h1x+ie4lcTrQ3aH0SCdVt
4+0BQyWaNvML/mkv0PpC66V7a8mchR2OC0+Dau4zQeZ+oql+TZDdSqHSFzPZsOQrQErGUlgeJsal
RQ063hKk7z2e2MpFbjVa7yihovlXj2EFSQmytl0uBoBOzVluf0OzfXUgxb3SdHoNoermZ2jsDyCn
EV9E2GgANFt22iP0lorgzZ3FXPo8iNAdFEPP6Qe/KQX5P+TL8QE7DLyw4tX7HzrE4P6a71pVjxSf
+Z5eyfs6FNvy6aC6KSn4WzaPC2x12fJoAG0N+BSL+ud3u+WblnW8r1iXhF/BBEOdqBEL52GwfTO4
tnqe8wxBXwaxuu24GrElILR00DE3KxbQUN5uoLg12NDpKLgQ957E+iJ6xLd0Ja0UbKgcAskG7SSL
xer4LESjb4f72jaHekjhwLSkGFR0uBrnmv3Pu3L8XOqDH4i8qYAR9ALpJjKMgXJEsZmcbKCcz3pO
jHTA+0KNR60jb4Pr1/8DxsCEEqPod8Qyhr6iccGWeUXMSA4XdxB/3W+vEE2mqlvnnbS/gd58tR6F
sINeFnQxAPJFSZfyguv+uw4wFOMEQVglGKomaDexaXm0HFnjdLRelDcvKuP9ZBe0+2KyLVKcCLD9
ehp4UkeZaRSWa2tDzwL3CeRBZDq5irIvRHHeT/umrDO8AtsrNL6STi099/W6oMWZB6pHj4wRbw4a
eHFS2kiPc5pP/+eF29voaQ8NRdA6q7ey6vyfojYsD4CEiQ8tkElTpdPZYrvjU6TCSOzgZkU1Yl4j
yJvF2IQp0gR9heXxjgHCYg9011siFihC5/L4AR58m326JtVnd/v2pzXJlzk0mZSF8zOUGBcdJ6vb
zxlTDo0tm+6NOYxTCx30/j8C43cZe7MP0fQCA0vwv3avqznMYG0QqvfP0CKBpX/uHBBNGFLMeVaM
kscpYrKt59aJLY5/aI/KYlWaNbo/FdcCKxKEaWfWkcgoQUSA4GCAbtlPJFOTjewKfEcTd5FSOr+i
Y5nShVdtbSDwTcsNZbYzU8t5qfaZL9GcDhMPVqABPKZNIro75NyYwlbx3JG1zFyglSGe7QE+e8Ni
UIkKGNRTpkacct5TU6rSxkHYQ/zRAFZN6pbQ5wrvHxmgEwmFUAS0oZLuFnSraocK5PTEq472t+7T
YAsNcRZp50EtGbcK2UHkgYhqQ+aPF8i+VYyg5smEXE+tDUO0BwWicQR3h1K0WEYIwRGrV7hddd1k
/YIdb2lcZZccXIhEjX39oH1SiULUBJJPIdAMkCjLRnMQgUyf2TP+weEMgxx78i8EPjddJLcGCXay
8s9ME2XFR986/zCaWIEPw14FTsnG0HejN+5WERrA0Yy6O9hGSF3YNIDPNFYttiBUuzJruR2C3Pnt
bI3BjVuT5Cv622lVDbHV0wvOdMbyrUoSLNDnnZTiF/dnIegKQy3z/0l7T4Ca1wDStE3OfesD7Tod
lKHdGiFUXtgN6KzjYIc9ID1MtEFLRjmWuifHTjdClfZNwi3DN4iZMZmZa7j4lIK0S05QtCG3cOrA
1CWz1zWzzAmNJIaTZVSn9yqXEs9fgUZKgvObQ63l5ZhWBzp1ghRHHv48JUGI1sRkDm2YP5JgNpsa
bjXR6qwwaBBRW6Ws5hkQwoOLbVbZQH2qDEUkHmbePGGHu+ShV3THiJe0ivTEc7AUyNliDhUfkhl6
/g7eLj/CEw6CmT4gebpipjnTFSo8gnW9mwfTJf8KAZIPC/CCTWhLC5BmGIyy1v+SyOfwkKsQ1j/d
Z3EX+rRkEYUsdj6uIsLcsVt78eKh1dVAUzHJAo6I7qSM0V9TkwXQpG0OXW4783yuv5AVTExT9yK+
GcyujD/J+X20AZJIr7bJjbSIazaA65bO0loXiTGygVhtCL5cJunuO31oPR4cl/TCIhpG5KA+yWkd
iUgP5/khTQ/dX3a287OnDo5XxlYt9NCZDPdxFY2XUG7Jxqyr5xxVyewkbMDfYoCKHQV4BA7Ma9Db
l7EZ0NTK7mHwF+NqJlsZ4BIjyfB0nPakCx1M18kDYCGy1XhcYFwQXLDeIP1LsgjTpDFuSb/esLMM
/MdTWFQqXO03Pfnn39GCQQubULyJG93+cK2XBuy7TE6iGVQUIXUordQFaaCi/FQoSg8Jsa4OocuK
G6cYkCZn1vdDp+JV+YChkEzkK9X+q1YZTrMIiwDol+KM2d0RpTII17tseGkjGGhyeeETWvewEaAN
PiAUDUEcQRCboZKr47YtCkg9c4q+ZoOExyTg4gR0aZHFgONiiqTV61igJ9KQThq5WpZ4f3G8iVrO
SItk4XgTMbjTjnT0ZCR1U+EeIC7Y9Vnj6XPFgl4bgvB8NHLbIoqIUFPSiVz1IEUI1au9x7US/OW1
g4+KouQoxxi512nfrwCE+ozIrSrVY+E4neC/jlJwJ75HD/JMoh5N8QT7UrbENBKl0bMQpkYh0uq/
jt2Es7tf1mPx82Xh7xP/cIWWXBWu71Cp9A5322lhFxHsRppN3ByIltdCLXDmhvKtcZuUKyNvVlrK
shrt9ehol1pijzRwjQ0LBwlPmePkJsNbwPS1gtG2CMNvE9LB154tW8te25oGSLn/Eiu00/barU57
K54rACvCDblKIXS64X+Royj9E7PKfGE09HNANkgdnV083VB1cY4ZtlEXf433meU8ExuYw7YAfz8D
XZ/gIcs469NvGWQb7KKmqok4gIzF281TTw1Dc8BtfBHDykQRgegQy2Hh9CTYJ3SfbifcQXeIeSoh
/foWnIe/R19m3H7fvAh7MmDHNDY4uodFFyeJG/Dti0gmJDv11EcvGzow8aklpD9HrykNWTmxnZEb
c9k7RFUSnNshoIzGZrXhpOQZ1KTTovdHfYQYVZSk203C5kmWnO9V+xQVTvYvOp284Ef1Agqyj99l
kVSGdlmsq9G2O4Q5V3XGipua7iLEyqegqqH7+B+ASMAZeQzAmlgg3IAqWCHIw+pQcXzXvbgQwNan
6RiSZQIDefxfMmdPbTsKJETR4o9DjRN3UA9YHjuLx/M1/TRtT/ZlLgNP6Cj7W9juVj3XCz58Fb0Q
LIUmuiqKSdXLn0zobUC1DSoq+HKRbQdFwa5F33mtNAdsvGtKfcjHoZjjfqptUOcdDn8N134Rkxrv
ZQlhkBgC6hAReb83M3NvzTOwcDNHMAsWSFreaZ9u2bXeIVv6DyjQAiaDmKDzphjHaVRtp63Lg8s9
RxvdqWUDGm2X20Vxiiot/f24vNnTLNpkufEyvg2cIfKK9i6KoZOPK1oMM3gbcutKn9idhNF8DSsK
71t1AjV+g86GwZ7OqwcRhJ9agIwjHheBXH3bPuo0foJpDUz0cxorGg8ta/Ezdq1LhUAQ+fU+c2ub
irwsmi7C8WqQNxqwZ7OlVmdPqfxKN3BfASko2TXqbFpz67dCJjT9Asgu3rsuIOlfJPX5VD/XGg/6
9DS2LpJa0CwCLCqIOHTIKqtIoxp5McIYZwJfrDxjM+TDu88MRFWYm486TRpZr+CAVaq6U04QMngY
OuuyK/o/Bc1wE1jVfcTsMRBimWYOMHEl07PsAtIfBSpGeBvjZxvyTHnNJYmcm+jSJ3F2AKo2E5+5
2f+C+qEtKzucyqnhxukTkzcn73ATN5kz1/noFpJWMEH8/OG5tv16KCEZQKhQ4blfMHLVPjuxJ4R6
8jcHXQyhGpHAOIYvqTl/dlOHRoURCRW1MDtH3yLxtAo0sXKG+oSYxaC5LK8yv3s7HCKbMqm3fSvy
pdi3UNWbIjumIO9E3QJIhb/SvzebppCDqiI9dKe5IYyHVWsUR52A2IN2xO89TYaVBNsJFNq6SiBU
DFhSZQxmWDiWVtXxm5Xk2Zs9I8Guj81dUtz2UyfnXqISDR7T2R9UlCzLxOUQz9TphjxI0xOUciSK
V+4+vvROYv3R4uU6TxRgCMm+YV3Ty6TSjpjcN3r3RUhKoqGHrJebZ63/uMfXvmmXOjnC4x8lcF5n
++GqfeKs3TzTH2MG2LEaWCdwJG004L3J0gr9hUrsWVNH8PI2h1dS2MOenAuJy7BFEt53hkRRTIh+
GVpExgBdZsYI7TZ7QSbNhFVgb+lGs6tNpA/BcNS9KCp6T4K88q7IYCIhKkmRv6SapbbVciTFu0/n
3GkkRKR2vffjLgq3EWckEdAVI0oiF5EKbb+0bSbfYb1GaNYNWScuDEGQLg/HXAw3zA+XE3keEVhj
JSX24f73MS3ghZNoK7oWzN36Lm9yImT04OUos+iUQKivm47i2AH03DUBUrkdi2RaFSrN07CjFrXd
RpTsFicw0HSTv7V9dO5olaKLz2FFgc99XtfNqsQ7a7cTFeUwH0oFupfPVjyqzepucM18tKcrM4QG
rZZHDP9ltUqHWTacX2Yf57n4G4XvRBSaXXZnw85SxetCyn/3B8StCyo6aTRd7qhDttgcfUqskrQS
gijC3V86bCF/gdVRoy7WMSJamHPGJ9jhVqApjOJpuvUYN1nwirD1zsEjSq/j/+PJxj1DycqiMYTw
5ZzoXypvz8ddrl9QtwxqTAohbCID2nPC6FsjfOWeQI9N4MUq5lpTA+jp/GPQt0aKXGXuQHjarajf
l+IxJRCZJBbCriyjr1fmcdx5kciqBto+kWjBhkTGHwYpWRcA1zZU+Gb/Eeo4cquQLZjrtwY/039Z
eJ8syzagABpjR0SaHRujjnAk1fixwj7vblGE3FSwEpHtwSS9Tv/itSjlzlueilQB/MwMxcNTs2Rk
5/bwIYpTBJkqpVmNVg2legZj5uHQq/PtHdGnJqXlKA22s7x4mNPpmWVgGhlFm79wLmMur7jh/dOV
M5ZTLUoZ/7P3AHk7U+PFN2uaDpW7wQ5qlLbjDaHMaWIT9wJlOApBL6aztnSXGmCR7iRs7Dkmx0uU
n4N+NcJDVQM6Np/WphCMQTHCG9teRe3gtxsX5ICiJwDnce7PbathSb4AiMKxhpRWG3IYsclt2Olj
1psIV/01gpjZ7nkt7WRXj3MrWxQYOpbbKmuHbc+jCKRQecWEepXr4/fnvvKr+Vd1MDnfRRLBLoEd
D+JMUKXAAMhkPJaGXb5wFU0vIfh/i3WXmPWcDMs/aEus86ax9q+S+jPaCaDsGCKMKeTbTzQ96UwQ
d544K+w/qcJKOTNfohy4UUP+GUecJmcMTCcrZR27UxM2e0XrkLkWPjMagiJRyG+M+wIZhImaZjhx
l0pL1V12gQbP3vxiK/a3uGVX/9jp8BaopS8GPidEHk9BFindsyqvGsFEMM8WB51l5j23MMxrhpqn
+rGfO9ZqnmGPLseAtNT2hY+GpCpGLnR9/YG3mdseOxOhmKRNjjmU5E0MEkfcXpcWNYgA5/N/bp0j
2yWPM8kQY7dUpY53z1c0TPwea4jf6Fp30TibaqPaQxs+hhHfWKiMUlBgMiwFwqsqwTE2hjsFL+/k
1YQcx9mekMwZx+qB+W6cilA8E5w5O4rxT0+P9QM2pnf76fgkoBK39phCuMWkgIRQ0kEuU34M+s8b
qmHM4HeNibs60cNEV6HAyQ1UDHY2QzoxrSzfYJ0H7nRzhH0m+XZDLyY65K6ex+9VJWFxs/O3APAf
3tiRzRkeDldmAH9lmQH3r29Q2be3P5E5x4dratB70i96IsQZZSI+dYXWfZw8Q6PvuRPB2/iPh3wj
LwobW1cokPEqt1X/zw21zeg0Ds+az3knrpZQoSKEXlVBVt1i9dyQ1b1J4qAZO/11TlzPbkVEI18R
CYmNIQoBd6gTqqi5W2gMBc7zVpadgl3metpObc2O1zr7hXwXwOJX7ZDCZa/UeENXj7hgjbDDBtzQ
O0VdEq15HodfrLGoCt5EyPzP1UKhmbwzSKYOFtOKSFCzOPz6JI1ZDyIcCNQ55PXzelwNA4xaHkAP
uPid/tRcNeE06HxIyQ3wXP/xN9COrubwGcDP++l7cWaBJ+3sl/UTzpb8/eLi/HFrh9yqjf0cBKGJ
rjpqYn5SnGmS9xZ+q17wbD8nvfN120zgMXgnFXD3HokNh4P6ZE1z31mUfaIAN43I1caLkmew6blv
S5Qvi+JQjP9w3WifYOEjGyG4LFR47teVzrvokqFu0twbv4yYheyB+MsgpPdWOpum63eMWbp1tTbH
H1cCWNJaaiSnfs4/VuvzRQCzsucIbr2EbM7oDBJzSE2KI4wTJZU0VEkAWrUHppuw4yJJ4TvUfr0I
SnvqVbKPlO3gKFW+t8S8i/JvimATDenRUIxzlsEB+8OL9qoXz7lsrgRovtYySBNHA3ZhfPzprfHu
ubNueOxrPZJhCHFksQ0n9gXFig429HtndDeKIAVCtF9dAeiCEVcsQJnrtndTWPmEZI6zYKt5cAHZ
+DB19nlmY5KtSkgke0LOqtlYhplQQ7VD35ql2YJInVDvs28yBqpCoMgj6YKTWigpvfNsTdxmACD4
ZYgyNbS1rTL1d8CO73lTM3HDr9x0IiHuifD2eqR1YHhpVQRt0PtqDbsk7bIwzd0MxP0ZiOuDKmdy
XLvJn9FuGeiSA0oqSOd/9mOhJGqM7PbzdlF0EMxN/gzv/VmEJTAw0GCuFFObb0ePGi8e7da4Gi3m
Q+5sNtVAWIzPHcyJB72OYuQDI820b+Y6BnBWgArtXU2T++WemIIBywUohQ2OunSZKzQlH+0tVMPu
VWy+AA+QrUiCYOcrDypgfbiELcDkqMLfLN5JpvtQ6sSxIjh7w+VE9HBJRLfL5UwFv7o4++sgfv2+
GLBEJND+altp64YW6GStMsUscT8Vx9J9e4bra5kivhOnFPFI6meeE6Eh8Id3G4n0B4ZYB+txodKw
y1CqdYDrdgBjtmZjYDD4jYsTH84WasshPiqwVE9SquuZbq5ZsiakkQU40b8ak3dCUtIEHYq454wh
vLy1uVS8Xjkzmx7S0GVci5Vzs8hRe715bCJstJUIymq8pskg83f4HNJSdUc4SUPBphY7mvTWvswo
L6zvqQmNVZpQNNvB1a1F+PDGLN0QLgjR3peT9/upYvtz9CEBK2jxposurH/kafM4Svzo0ANQm5Me
HvBmR+brZVKc92NM+fSUB5KjfFgZoN3Mx21HoBvjLN1tiwR1hO7A245hmrlmXmSncXbNkC/3kb+g
1vSUUl00uQhzV1Pkji7ukTXnj3ANavlazK265hogtRggJTKlr6X0sHbq6NsmuM8L6eB2TDGDIGx7
m5mtf9/9H04X0S2ihwQOIF5vE3N8u+aDNEQbHJmAFenWPwcqKCu0FSbh+0ou6E5xoo5m4nALCfZl
bjGhvsG6CBReBciZgz2RnebxiSSr6hYJKFdMzZ06y0hYG728QnPD0um4umLcoc2k0w/8zd4aM2fX
4qtope8x48zl4LJP9eqA9icMp6Dx1YfVINtHHgfIbvuli/orDearPphYoo86Lx78E12atPTry5uK
9uD8WY5S9fZMqLxhWNeMG0/1lnnOSgc9s+6m+muG0MjgreXCh/fWKVLYE9hgJSVHvEcel+xJl0yf
BoJlOSVY8Kh4RAX7vjEaXS4VWeSq3E1zcg5mlbMq8nNi9EzJ4L4poOoLEcwmwNi5xlI0Ppl8K6qB
rD9OYkiOY/vXJ3gbChtS72+naibmL1c4NiOH3LkZb7ki6/BB4lRHPtIu7uTG1pQ+R1A9i3kfAaje
qMYGT6nnXtg7fa4Ejen+C/6S+Fn4PX8pNFggn6wztuVMjzv6lDs4crHln54J7ipBCqS832pLGggC
WSxPFJe4I+xRjoPg89Ygi0zwbNAL0Nhd6+hEoqbL3Ai8TeLAZ+Lf+B70BfzYM2sxFF4Sj1G3M8sP
FQsyaJRDulf9pl+aJFPJonDs44NKInz9zd4n0O15HtBn4h4wugfB4TkWLcpBH8WkEQOMaGgzuWbv
k5VVn/vIo3Vt6dnHZaJIZ/Zq9BkZPcc/zxew7i3uxh10PJelP9YSu61lCLqyVr+wQuDsatD1vrZn
Sg0l1/WcywlrVghuowtRLdLtsQ9+HmwcEEw7+dVOI/BYA66aBKkfpMIlexJQ/QPG7zM4P9BlsDXU
QWlRVP29YtC4UL+L82afg/L9cEATBLYjmB+UCCSbKDoS6tZTL7igHFWIfCI2B/vacIWwTK/EwO/2
V7XFShiLwjQf5M3H65h3/HYeqwdmw9AnTrYetuKVViv5apnrCK0qUsU+GI0iwHDjRkF4LRvg/4NW
mAJAHpE3bAX3BBauO5RmphsP9hwxCEnYBCPBrT0qk5j3eyIfix0zD0Xk9p3YWq2hws+tRkazcPGq
oAi/7/RFEbvN/qbKWPeBJx74zNh2RkpRcmXt/ir1nppnnyBS8HtLa09RUk7WGjezD135yghYQO9x
+skxPjWy6Z/RwQGoTLtFPYKyYtKWONNwyRXRHlIbsuGKG/8F0v69hiPXnSC2w0AnsiILixn0mjbK
AwDnrKUNuSHY++Z76XBJquhEaJsG2VHdq1P3GXDJSZC5NcgdjsnLwvu8OTHfNRMFfmpiTEfUgavj
JFP4yh3iOY+1xBh5NYhxdTG+bpjwbVSs77UEZgX/9O4cf4KWm7pdQR/Txe4TWI/cWqU/vb/Z3FUu
B4M4RqRFZ2uWpOgJjlcP1++yyrwiXMzyxkda+ud6gct39bXXHjW1KWFyJk3P/Owp4vZ2u2qG3+ph
eduq/aRWi5FVd2n5l4RKJx8JI+PrOtS5zQ7Wc03S3nDmSpSFQZcMsMz5inN5CPzX4scLz4mMyDpj
FSPhb0UfEn+Qb6OmQIGb8vNcSqpOpRUlPYMqKx3y+rlcmItCEM0k0kgD0flyXUP+JMBX421SMFty
6Kkd0YIWwi6IAZjCwm09RH0OCsIyrppAEMpp1ln9rFcPTkynwxYKoTy6Mt0btaXGkrVQmqk6Nq3c
sjS7MUZQCs2e9R9s/5F/oknXcsQ4RKpuQP2tPtRKOamACLmrL8QTWxleuSsqGhsot3L+ffqHpZ86
98zECSlIfNldK5D2HMnjyMYokbv7EqYw6MYeMU7h+QTBvdT/4c7+lylKDD42pBl2kJVtU9sB6Sx7
Spgdva1UlwcNhvAX4cexMg9vaElsz/+ThuWx89peFQpFJn5Tof8E5j+DEZBPO96cu8r/Pcb31K99
dY4zsJlXchSQc7hn4fJ+pUzfRzd/7PaKMVUoWSqK/On/7l8vdrHCH+34SV3WcAdCV1MCwxnEgSvX
mrhPA9bJmV5A3T3WMrAd+2TiglClSV83esvd673x22e3qtANooNIYdYuT9UcxluJXb+b4RiJ12rl
1/dZt0c+ZMkDCBYLtMs2PDu4BMhRQH8VZ1MajTfqIpX6hXAOvuxSLloHAxdRCsDd0Mmj+hLv7ZwN
BELQTSSm4QTkCp5dtZYgrsaHTLkndNV6N7RCXWE9/AL6fISdqvCAQdynJ/ZXsubg/LLOiW5P8T1F
HH7PPiJ2JHcHgyMVDoYP5YohVt0T0APh7qSZbC0te30wWMA66s2Vguq4ypqgXFO3x8ZfOk1Qq15h
HTyLzb/KVBAyQEFwZLSZGeHr225dV6077gikt4QuEPZPjbgrbVhEPsbuIrmiIQvkN6SR/GjFYZNr
CR2SbDWUF0eYgiCeOJc6IEs4wNPllQMx9EqX/+IXn5OQEohqNldetO5UYp3vx+Bp5JWwba06hAAo
1haYlfoiF5RMM7b+g7Iez3VLs5qmDS5MuT2DH1uw9BDlBTPO0/O+nl8gPwvgmFdyk0toZ4xFt7a7
xNfq6iR8g9WcBaNjmX7zi4Xf10KES3/YNOCIaUGVxPah0uGg7ROlPgEUYxIJiMFxqwTHek6II8uv
XB3qA/yFdJEFUXWLa7jMzzc5cK7zUwV89EXERihTh45F1Xo1sf2TFMoJ1Y46SHZVgHqodu4In8Rq
9VwX5GqgN8qMdrstjZvIyp8JucWsiLoET3aknJ8vZGFdgZRzpv3W3kEs1kZvfnXsaK86jKnH69Mc
Xw5EwV+TPrsd0aRsQoOO+vKuklJQFAnUqAFIQXPC1AXfn473KabljJVf4ArKj+EEArVs0B2J1wnL
XxV7OZ+8BYYzty+tOJG6X0nRs3r2zYEH7KfFh4NZN/cRa/ozsnd/dUIehIP+hVxjxNjCdhEFHSlf
EtYvqH8pKFLGGIhl66EGf+YZSKGgOoDIald+hF1WNZUhY5LoPkstAfnRiF9Ik96VrsgHjfPe59sm
3HlBhXTlDo0JszYBH3DAx0lyW4feOopZZHGUHepBjZrXXrEB3h+7Mdo0rOjQLV/1x7tZPlM03uXI
a5g0FqSXEkngt/QE/H5n4DnxFUdVMIXjirdmxyRFfnlef6eEpL500fPfriUEBZldO/IvPO6LOO5w
WYtm1JF5QfGtEmls1AOBijyeAezvhNSWpF79FRJU35jD934i+F2zixr8ZbdKLOAkBG+NtJto2H4Q
2IQYEDdZPtY21hneKXpVw3j5w3Phx8liysnzLOrB/tftXvH+uXkLqvSXD4L1mHXlU2fet1nHYGYf
4TAC3MuZCQN6OqT0mignJLAZAvw2K805HceL1y/yIm5yCNJM8Yr+GvSAllaCIE30YNrM0E5LE4hj
GYaakEAC19bf/VsKK0VS2+ZSm5CenAsphsQJDk/5it65sPk/Pov78NN1iPgRpRORqlT6c8ezADbv
h6JulmC32TB7iyJQJQ+FsQ4vFw0RIZKtb+KE8fPugtmn0Dm1saMM16oAdNsR4aGjolzMax6gGiID
RNBZxtR8juNW54Kw9KtVZPUF5tagS7m2UOOOiMNSdZr40Yjx+As2Ch7gyekj/lrBXxLkZThq4y5/
0OnVv9MBt9nb1fm6IZm+beb6RLzA77Ru8wpVE0BcLaiqMoJ5VxtQbLoUjI9YldLXTLWWiEKMbUZ+
SLRE82igXh7QsZOnYgb0dk8tnUmK1lW+fLe0OP2ViprcKSv11EoZRrS8xpOjWlbe2pDueY362rAb
mZSOcuColoaYCWf4g8n4mpw01QObhonskWIB6R20fGVUoE7Asht2S4x4Es2+Om0FFRm+M2A5kDjM
SHnNgHjbS+aKvI8IweiNESX+RnVqRUBwjFcM4wEpgnuaewJYaScmPvYk4IbhxH6LDmxp09J6OafB
lO2zU/WmnjEZZP7l1V17sIYUkmBBfziGjMeVlJ21KnRypIcc88+RPSzGt+8LUyuk2rBhr0rlcr3l
uFiVmqaKOZH8fEmTM+jzKLEWgAlZD3yTgZ1/TXSqsNbQNroqnjEbNvelt1WwHDcF6vaOc9ThZZyF
pGJs0kfixPhCUl4mmRKhtgQaplz23rjwUDQp2G/6PbSktmo8FBOMp2Qw19Coz9VA4Wx/Tvq+nYCS
JLA1vldQ/CyLJQrukKlNRkpmUn2rl7vRkE8EvJSSnjeZllcQMUi0WnPpSzXlg3LbrW7VTZr27uJE
NHgRyKPVK+BJFYYII0uO7NVHNy/diAlvEuFr+Sb/LIhcXbgNBsj5nQt6pV/Ka86bvvpdsjUKCTaK
iHcbcTyZEFzxcJYB9PgwOx9yUosGUQ9NvB9HTjBHiZL8bj1LoU5BrGmIr7VmhOVr5uaVtFrc9ljh
dIX2xRvDYhBDFScK/gY6eFsoO8CEGfVutKt1flp/3zYuyGed0glJ/JPNLEbAJ5t/XhFNMGxYmYO4
FL2iKezNJ2+MDpIrXkZAjG0RabTdqyrwZAp6nCi5c8ZUKjyE2gAvi09zUG28/qbeALVJ3CGW+BSs
Xv10qS7in/lcPizgCmsrZveUpRd0L6+OVeS3/tx7hqm3WLe9XcVidIXM8CTysjYp0poWGRaVHXKb
fPVPkSwFzYKQVX/FfPi+fz3bUDQorfqOqWSZwd2vmFLIY7nfPdQ7odzihObB/8E2X4feid1FwHB5
9wipp+2gnQsT55L8rplGSjSSshua2UGEmZSk54DAb6/2ng4WTL63TJXYMwvRMFSHut31fN9QeZYd
7BMzkK2ZeHgMXEN2PkK1roNndT7H6edXPwO1g9Mqw1OgtYoehQbTa6SPyGGHfHK0WOQ5sZEB7Ysa
qzi0kBCv34oXsAHY/HKbtVHJIiNBwr5RETCDGMJ4gIudaKpHLxze9EopIT4VnY2cdx5z7KD7rHPO
MWNMOQP2bxdzSSYq7Cm5JaQrsf/CzIwVHCbTjmKrD5oWxbqI+PxC6eCY2DTb9WnsImyA2SCRU8MU
g8VDTq/9JCvEXNa/+mpXpQRUr0z5dzuu57WOykDsl+8SeeHZk9QavxojHdNucI6PPQAImyzRZgmn
VjzKF9X2sj9qjTmEnOUq84KyylPzNJxj6aWld5RinA6Hi9CXAY2dAiY3zq0s2y7Cv+2vgixzr99c
PHzUjcPsk3FdV1n5Rd9eCbbGLROAtfki1b8Dfucg8I1Su5Egh1CHAzrOD6BOKwIICPLq3VCeLtoF
M4rjjdg//85BwozBPsd+Q+jdZGg3Bo3pWMOfjasWhESjiH0Y4cmY/gM3wSJUHBUo4n5bVpS8Uvho
3oCS6HRqLnvobBuIwQs1OPoQSl0hHjGWlP03pWaMru5wxOpJFkyaFZcwDqqpcjjC32vX9QD/8Tv4
lJzrZ5WE/gekk4TWR7OpH9+48h5872gKURN1zEo0bSI+DiFKoiSPo7LGFV+6plZhiIu9uE5aYnxO
vZF1QYtCxQqJhOF8BL7DV2sr5uURWKXom4J3amsW6AhZ+UMUO/joJJECc45K4uAlT+Zidz4z/Gps
bSZTAt0QbTonqEASNGnp/zllsbruFIx77vUxMJp1bjiSJ/Rq9uZgQ13Ax627ThyPe33KEAv9lkJ7
bsoRJrOseY3/HDZ+wetNf6eNWVsEJR/n9WVPOUA4b5WFSY7BETW8ryykq7C+5vky6mXiV2B+fUCB
sQvFtaorU4GShWwmfV7b65YBUASJj6oCN2HbLTnet5hB9HPH1qsoAm0VU33tl0BH5CTSUUgBqN+p
HoHOTlHzmweX5aNhrA+KP6jDvAk9gD1hM0d6EUoj08GFwOjcdTWIXCqyn/CUfyE6qNcxuV0XMr2u
jwENO2huY06lh6aKvY0wAQHc+E4Uy8Tum0qdUBeYG0JQzJ81U6TEaoLDXy120HoQgToVQYQ4uYYD
2sgjnrbAOq1YxVhIp9lI93b1VGjHQyf/STXIG/ri/E1rtS3D71mVerxn8DHiOCYGcyAzXgLadaLZ
CO8eDuEWV38uX4gUXVtKdFERyHXqFMpYx5C/+gQlaG7BqxitptYhDuwHx1VjdPrGVYGRkaS0YK/9
kUiE6oSIIrPty5EI4JWBBACF0XoxZ8WvrCrIY6a69YjvpO4ET7Jqa/o2lBTGssjektQs/YMXftEv
3x3mKC7sjPtTefatesq4tWqak2n02LH64Q7ohgV9T/7NY9BWg9q3mUMdBwmzXBjfgFcBOg2nHHa2
ejm3a+o0pu18l/Z8e4aliHLlVB2OOWPtw1Tvr8/ygQ9DgDifFE/eqekaHS0cCHPK3MFZzdYQegoA
looTtbrnhWUMsctkcUJSRBklxaWQ6VPysYgT5D0NpOiX5I+OEBazh3N1H0nPm3WPTkeRtc9nX7Fs
SK0UpN6liC0H6bBDH3cw6VJ15mnLdy6+cWmmC8dOlPJ2aUmKWZrDxukIXCS9bCT/F6mcRVSbxv9C
Z5U2dskldV/1gGh+4KL8mfXx/LHYWrRs9E1mV0rFV72KW9fYxlCest4Z4yRTPHdgX6pht75a26Wn
dVjaoAQvVtQl2dGa9I/spikhVYvOYFmi7AZAy8dejPXVR+GVxfjj+JS/o8OvHhlZQUeezFZADI3W
jP5cfa1CuRmrPs2FVMOS34mKA5MZ3TfkLlXJgjERrJVbExsTr5VyRK357vvb2fh9EB8ggYH/Wjlp
OtXweujhAavz1Sk7S3VgDtfu/4PJnhfR29CfgPTMX8rBaZWrEwKKGuXLy7FwjVpBj+IA4meFoOn5
nbxh4xuC5nrLDR8AcjUaLYDK8MaA+yQxmr8c4RRcTJDDo1ZIuSn33IL1GILPeOG66pDjpJPwCj6M
q4wN7eK1IOpORijRt/7neeIGoMQqLSmYk1izPZ5m5Y2TqHzBCnKu4zyuK49e6296n9x3S27ZcoKv
YI8JhX93S78wTIk05peniElTUKkuBAjXJlR4oVvbnPqg0ylDZeAM+IpUrwPVPjAinLc74bNDpBph
2mGlZE0ps0UruhYPvMu4Gt5xsAo4gqkQhFTCq1HKoA/ht9pVaIA5MNL/GMr8y62+en4ZcyxjdRau
e3xDvGT9n+7XgI+6mjQZJnaSRhYwzQNSc466SwX7k+GZmcpzQblIxlbd3hV/qd5ewlgehQIhY7Qq
HxvIwbSNrAIs2KU4lwfdYvTY/h55oJi4hMWJcp43ariSwcnoYIRy3DEMvt7KnvTNil1tgLiFceEG
wT8Wv/xkuCrJJ69ExbhTgehF4b2/I2Zq118EJgE/tICMXWeJem1fOpOhGblVLf/pCsPn02IRxFFj
2dBMfiSS1J5U4wEuWT0WivmMbVY/dSHoJEG5fEKMhmNs9yF1TYSwhfnK3JovmH+00Zu3cguh4y4T
g61jHBSezikXNV8GD/AATE4vG9PpR87+rVSpVE0C3jrY2DZZ22tzouXYUg8NfczcyYViNatstveo
Vfa0IRGwIgJ/hvBsM7ggM2uSGpmPuI77hXgLOFy6Rt516ybWRX8TNw3Txmz99sYdoI342vwL1Yg+
PmVi190TpqD1iYEDmC9Pzm/UWI+rUwElpl7NgPmmFYugjvtmUhAPJdWJdQ9hpSzUPN9KbK4oCzoQ
iWJ6kLRO6QEHlNUk2W996qu6IUILnI+OLrmWvuijSj8sVzuzrH5NevFNI960mpRhFK8NV8lfK7JZ
gdsHf+Meuif+sm7lO0p4DR8cXNtrF2XIFcYw9gk4yaYeQJUe/P8wOCg7++cUJfkIyiMSbRArJn12
NrR8OFbRAe4sq9LafoxE5cXh6lQClGkBDXvFQjQVLLzF4AGKWlr144yrzW/B5jfqgsIikI7lbYr4
ovcqu2RuB76OMeUyC0YkKsUTnm6i2qOaKtmZ62hMfeE816Tx0QrA8RQVExGpY29WmdkCaoARg0ZM
qGDzgaJC2EX8PNEp1O1XzKVeXJDoyGw/hGEjp8o5J52jOUOVDpkRUZcJzJQ2KyA89iX9fwKdwSbt
cc4bewtu7g9BINgzDQ/6h2OwqI/KQbT3UcqPAZBJ42yNkvqtaAP5EYyCrLyfel8aMvcB9Acg68Sb
fAnoEkkwDFV2Qt5I6nbDqusCv+2iVX7+5P90onxi0RZMLrVxGN19vglydbgCK9/m7aC/hu2ccMLB
XXnQwm3mI6qYV/1itnUvZBJ602Y0q1Ned72C6Q6CUyaA89z9AX8q4mrtSPb8jiqos6ZGPR7KFsYQ
/KL3WRXI6LqI3E68AzDufu8qDUIegPwF0MxNJZQmk51vOpl0tvz+bVnS6v0BhY9eTR9bO0L7iqLw
sFrxEIPXuzhwCjvHl1OmWHB4tG90Ejg0xvb+uzSsUTBdlxxxXdPPZEGOP8vzmOcDae3E1HhUac8d
r+4ZM2tvUyoe9NOpordlyGHTOrekyRJ3jqKuqULvuslcAN2spc1Knlyky7hc4RyAFsADKqEYAPgD
SGhXyDeqGG73pJ60q4ikrIPcwETSOjkFjATg319KWS6JenszIc+1xZ8KB6Ms6+a8sI213+Aqet7t
A+YAsusSvnG1uVWW6hx1rwEvWp9oQSeDs6HETdFx/KlO6s6jEidBMVNuvVkrclSu53oU1qsx/N5H
4m4yJHqd6FjEg/7S674VPHRXSYlZgVa+WkbWk1locdbvF3Ss8cOGmKUMxwIq3WAdzICYhsYP5Hjv
RdSQ7Ai3SFL4wz4yAekM61oiFEZZn/uamfM1s6eW7qgmBaSG/Ymx9gpLQ79aLZNWBuLVksr7CSoW
AMYQMeAwWNvRzsecvOKhV3cujXC4i8SKbDBwiNDAIXhYSBIbPmBZ2fZsu/ZLdFwk9Y/jZdSH+ARu
MwIuyix36MXnpd+eeD3eJWSV9ZQB/ukINKjlKbrrh9vLKr4UljtMxGcnyMcNYf32wsiMrIdt/Qxv
kuFj+tCWaJMqDSAeu3ygnIdQqRYugbXC26MRDOBMM3VKZWUHZZZs0+g/EtAVrdYY2dP6icJQj39W
98FuwzC6wHlXcEaolJ6YjhZhw0HI+/Q7cuhRXH8CR+Zg7GvbJeHllL03fqfaZRql6n05g2cLODx3
vn6RKohzwuBm2RhvIuvj7S0vHR5Vx8M70vJMAy6UtrjLYPPRnctj01Q/+SOTOH+1uTpQPPJnr/xM
PJiPzIpVua+6c27TpJWW+UFNaUO/4ULJOhNFr/mMpuoLWyziEliPqEweaCfV1ahG+1V3+EJKmScD
J0e3sqBblMP7AkAbKUNL0yQNApPWQ/msqsQxwAWpQKaDZIZ6f5zrm466s2LqbUGxMXbmV0s0VJ6X
zhGO9SaO8TMs9eulB3WB60r5/P42WFCUcNER3tYCb4GR/n0jQs/H239P7Ga7rkqx6SHL4DL4CUl5
w1GsKUmRbMcyhhPaHNH5INtPFqWf6HUljqEkBlXpgkFq61ks6NYBHvO6mb7n8KtXMf70MFO9uCTN
VV0t2Hilx4/yuD7uBoKpuMsMzkGTzTr8ipje781km1a1B1sxfhymAOIkKLugjHW6122sEtTu9OJw
xE6FGxLFpT3OexHFgA99nHQ/i66iovpU5VxOzMO/FapxqAi8FsOJgkxJ6psqDa+4Lf23ftSeGAWQ
aOWVO9FPnmE5mcBdX5qbpSWsmHmhhx+VMPOCiViBty2wBUKE32Qtw4mdbgjDkFPeJhjhjYEGxsGH
yIybYqCuJTR29Za1FO226ZfkcuE/6qMCwwac91heC+5DLcHZ1aNg58F8ygVRYhTjfe486E+LenOR
ZvBhMrjSihxu8kYsivfZ7rkPu4WARabNs6WX43SpQ82OtwL13LYyZfAdb857S03HuuIiOy6FDpjD
JIotycWZ088jB6vZEC1bsNPuHdIsYxiNYd3RtzJR8tW89AJTHsj97kpmwaZmJ7lIgoo409g6HqGq
Bbf9HlCE3scpVu+aVPmf7P6SprMth+rM6QPdc95OMwcqf98cUFxU/4VWWMYeC6djzJdqsEiEZye8
YYIYEtZkJwKN/HLNteVV87rin0jNXINa9P7IDJWgz2PjlQaCCp9veKEiZYykYMrwHmMrcdDUvV58
C0C4/4XgYO41Qw8HJvwKmL+CnZilmc/iFGJ+XO0lqm8cu2y33xvPSJ4u+cWoc0HB/PkEvA25U4lZ
6oed8Atu19+xqkj3EMbJuPETegPSFv6yZCSnjVxAAQ9FnwViCGxI2RjnpfOHYn7FRntLL/h6Tv/9
jdpxkSLXBJ4NbYSts9dyjVxXrtml9XqxoWh3/0hTmBxw2gWgwTtC3LEfpl8GShlQjndtB/SDrhtK
pr07e37CAlgQNpGsyqlPxhayqVmNpe0rIPHBk5dMqpIzQ+sNQ42eHTl0eDrgU2CjVmSqPQd4gbOm
Q70ZhpglgGjG2Wy+i2kwApqg6KJVstOSz1XExmlTDgbCfsSF5OmBy4zQhmEkl3Jmt6XzdnPKfT2D
0nz1BD02Adq00Zi8t8cRgEZpOn/i30OqE65x+sbMUPT2Ka3W4Tteqymu98HVx2l86pVy5zT/yMXF
p0S+/a99lwbbCnFIbZfgscFHBQOAYAcr8XtuTCo8jHAEhk+OW0+avaR+YMRJYhm2KT6oy0LJfI2x
pfasM78bdvKt/OojpQBFfMIu/6x3hqyKISRfqWnGoxG8eAggeMKHuQ456E6SZ1kPeCsjiNWy+wt6
LuaS0aHd0yCvdVst5JXGxchhaKZlq6tMFE/4NdmG0CkA7KU3iyStnBnYf8Q4Ts9Uas2BszCdSSJR
cuWSwV6P0n4Q5DwB9lg21Xq6UWWo1flQ4KPk0+5PnAstMiw54YiQKuYNGyuYt/p7jl0nll6PNjvy
93SVHvROsWjkjXaVScUG34Yvk2TgWLY5jPEkE9A/yUqHMd6tBqoeHHZhGMJxd1O/B8RHmw0JpjDs
G8vk4TgzhaLqdgL+8hta/737FhLAvgAta/SoaDhNl1rh/E7kz4GqrociA/fGQgdGk8u7zC23n0OS
oZq3uPv92qgXwxxC4a5U6McbIomQD4iqyBcGcHSi4kXKPNbTrVMroWzJjNJf/L7Kr4Gi0x0+NDSa
Cg9GHJPmEk0w2IF3wgxOhNRRyklIEDXcKOMgy7mT7kVSbXjiR9A872dB2FY8ZIz8uWX2XV0m3vRC
s5eAIg41+5kapVr3t2aFz5qXNfIuyNfG8PnKLgFBoW3QWQAcdcEt8ai9iMlaZcx7RyIgxGEm5VRI
QghOLBVRTHETP/L0s2WIOqlu5WTK+hc0PHx/Fa2dGiebJmku8jmx0+cHnZQI/91UZ9gWi+VkWZHq
OCVjIoGyIZgW8xvWN2pc/+lazqGAMcQHWBsQMHKxPcyrpNlIw2eE2LHboa2JnjZ5n4gNlGMWc7JD
Vz+g3PvONQrwcryltl9OmqNKaA2Fg8TXX69tWJNeSePo5YGmsh1Ur9SWWh5JeWBtuAaCuKu1FMxW
jm+czFMgf+dgdTXa2dqxt6Yg09V4mTIBIx1hDUirKTdxOpVTZLR6JeyoW56ZRic8oDR41kzja56t
25gxwy1jr7c96Nn9JAsHNII7teMUOqSeonzPXqp7VWelVXW8q7bAyilGdYbSDz08I8Ep9cbjn/K4
qNrqGSM3rEeZXIQSyp6v6WyZbU6k96U95G23MBIeXsCAzPNv2pdbkkUUeeCucIAmDI0dS5/ski/W
ZJdD2p5fRQ2IJswcWA8c7vbQQqFTykTg80fhzmLohNqvyhCnejorAa7zN/bw30oh2AV4vpO0UD9F
Pg6OwZLOr4LbxCQBhaajcNgi1zPRCnDC13+S6WN9oKGAudIR3oBzBuebVQ4CcvwfPApP/iVbDUxU
6dD734BK1oJZiD7ux/Lftw9+hjdAuJqrHaZrpeTKv1Jf6JfxkvsqKlrjrgmY2IPSkWHXNaJZqByz
iIuOd3SfeLq0rIuH7Yw4bLtnu6DGjU4rj2HUWW6dycKZjW+BD1kU7mWftkKuyRTn1WOSh4B/Be13
yUTsXL72zzN1OZlYo1thnJYAsH2zbZVbGHDo84C9RpwcisVLrVF80lJ2cAVmJHAYL1F0cVTWx9e1
WQR46Q1Lyz1MNxSOCxrCm+PODoTBosn3cIVcOlXRBfdOJT7WnviqmV2uFKLTxEp8Rp/NjC42Djvi
YYv//Wdpg9Mjj3j7yPDAm9JxWg/JvnXIupgNX467leDstoJrpt5Lt8qgaCdiO/72y07fkvV1LO/b
fiq5qgnrM1sKW+FDodb9v5EAIh8rOiDhlAyUfoXbOkKj+qETpm4+DpPyZTCG92KzgiCtbDhalDvt
RcOi232p8GEu0DJh2dXB+AuYIL7xgNdTOFz5JxRn89C1mEppCi64WyQwovglSm9yEH+hB0Yv9O9i
lqO56GLc1n2M9bgJHrBmt1TuuIkUjcdEUaE9/Ztfa7zUSHpqHL+elnK4VBJDaWge8McDHJmZ+l6f
i4Ss0AccSIsUXYqAc118dRLasOPaykT1k2IcV9IJG4xNmqvpMUGI733fiMbRYnBHK1sGDIifW3Zg
vLlwk4cStVOvKUT6wynlP+wL+e4LgFZN1/rHU65fiEFYmux8sLqEUyoQD4tLd0X1SSt8P1b0tk9F
TRTiMMARs1mjBZdKL/qsDoye8pHhZN2k5lswyVJXptWdwWNEwQOPaHzQf392I2i5xd+ZKEI7+i81
ZbKdE9Alg4lgntjcXWzmt6zsYwotfTwCcTUuQyi661PlspbQlF5YOh/9Y0Y/b9a4TBWrXj6TPHGk
vnFAmHmQqe8jYmN76O7HEVZRcQSe4Zi3iyi35F45JrT9djiqLXNAgkIdWXIy5uiUbpqO84JUctGH
KsuHqi97yHe+r70nA8uFm3nZp7N4kukXbeUhSMTpWVSP1argLktttDOlo+xX880NGKHKtJcHwhgG
zufg9scK0pHcZ97yst+KonmZ5xGjSIfchGnnthj5w5WY4Fku9NCixtv89W1Xu6+afrn6Bia1o4KI
DTGF9NDMK8jlzETB9cbyUkmH/XmKOJ5aG0cCx3Xh+t9J/qxg39SMgtGSBrjvA7e9Zn1R0e7LdS1D
loAuOdEo/SO1Tk35zCv13guNV1L/pGldden9o3jlS0fRVufPiqO61xkq2V5SXb1vXtbFGXJXKYfO
h85M881v92rqWDZHJRpqhSXsPXgcZMfj9YoR/u52DB4sYfKUuWw/GVTp2/4rDa3HVH48zjCg9QUS
bOvYPEXQAXlutoQq2KN/ublLIIopG5dfyOh1kk4xMN+YiKeOk63cNmyPa8p8d2h4YMVplLRAPpdM
+i+J9E24t1znG7jG3DULnZ9XOK6Cz4hfd0/GPBJ+uJLG/3gvpynw205cMxCWIIDKsAy5I77Z1tBh
7GIzE9p8ivWD2SaNUTzrZNAdKUJVd6MLbSsWE1GSHTIhkjk3xFyzE+xTS0J4iW5p9UXIxUk1qgIw
rR2rwDzNDY85i59SQYWrDS7AXoNvAMihJMLsqvWe9qDebaPSl3Z+rbMl7m+jR2LsW5lKm5Qr9ZbA
VhODJv9buzY7rDeTM7gqMo1xSxQtw09Xv7lyw4QzdTHltOFqr7wNl5IAePQGp7nAZzN/eBpazkOV
OCjErfwF1V1D7pxdCA4RGrpldjOg6oOdBG+aTD6Au+m+YyJlzF7Tp57cRgz+Eh+Y09T2vo7H7OMa
K0rDPHox+0dp2wXDN3uGq/Y8O+b2s14uC3LG0Y4CICoOE4tXJgEalQrItBi6xm8Ytv2UM9cFfGFe
V+FPEasq8jWA9PfEx03W34kPhG2tBma9u5Ql+nJzUIq2PDnhsdVS6yh3Jzen31yVJI5yO94P/j9b
O+L21RHZBT5wHvpghnQDz4DIgQ1Blj252pE2k+9l2IG2qJ+btite0ESDq7Ng3+n6FreV2CXMQIqX
hXr2auEiIeIPQizYD8rRuNQX0hLYCpGTawbE1N1tI5QNQK9g+Ag1ZAFePFUsY7pkleYPeuzv2NOV
42u+G0aQGqafg2ZUBmoFvEX7PiQtrCBtPRUi2xuUwaxkffpvN2tKfS5uH0B/EghbnZoB3lX4VdUs
NauL9A4K5a6sTbwXG0JRAVP+er21mfmIn//obX9xR8j8QXpjmQIB4rBCVqOv0IZDoIwl4n+bojv9
gI1Fd12ECP85VPUo4T45KTutVJAM9WFOKfBUaG2duyKOZW0/Kp8LGhJoh5ArLc6ybn7TX3LXR+us
sQH40MtmSkOp/9oILvK8IIZ80Z+j7n8WgwUDJA1P8j9Ov9XL4bSPsSvAaNQfFx+uRY8S+tPyXRfh
xo286B1S4UEBG4Tc0dROeqPNGWGIqlRoqYdMLcxJrAerK3TxzLfqDuVa7rcyGhcjoaO/KDdwula2
rFWdSfBxzIFKRAkxzfRNnJQ6ncploCslxzcwIzo5F/L9tOwBudWHh1YqQdc2yUOk27wevNucn4Nw
LWyfGEo0rTbt6hf/4ks9vTM6tVVY0NslKfxLWq9LzzIXQ3T3AJybo5fnb4G03S/bGd4Xv+YLTcEt
hDlR6KBShAm+CseIq0vIYMlEo9GHcB2Ii9g6F0dzfDaVQqakvw9RTkKBXD0RWE0G0w0wYmN5zwN0
mlTzLk/y+ivv2Snf7FC0mgjXnEWiXUag+LzVJtAHOGGCR+CAbRCjPEaQGgTeVtDYQTVYQGFicVZw
nW9ZUSXa6wJ6EZ99s0SOuL1iMiselujrVq9I0e17+S6Z93TZjJTmS175VUbs0GX1TDB1FRaK96Zv
0icoSgm3Dp2y74C+DOdvNGQGneBS+3RqDU5jQZlFV8tOwLnXlWonnToGPX5if+xV/modWsyaw3qU
c1eRogk7fWsHUaWbyH4wF7eCo6cK3WKWCvpFadNWpHfoNpzcWaukrQts+BfZb7ChTTH7giddBmdG
9Qou7TUvQDq4CY+DM5hIWnvN9LUe63moZgHFT+pTgx8fjnnsdO2J1f0MKsz8udS2TbOdxYIM6l05
rREjinJJjpYMvxSZ6kA6G5PcQAHaEVNWBhfMIWmYQkBAlJsneFdttooYJjs4XbRQu9juNOA3JpPt
c9JKRQUGarrzdRUNpsZO5aTmHZXSI/L845CMmnMJi6d4R1eGXLgF1kp6obrrRFtKjNnqbEpVArUJ
S6ze9GimmUk/+UWs04us2BaWTGlMxHOqEYhVQxzk2XSEQ1bzAtNPJrNFfz/abhhzD8fm6O5JRXLM
iekPQmxLR2NBw71MVk3KfSG6umtyVPMs9v6nYdyMWhJdCGIEJwezVFUKaTdwqRvCCekmDHTdSkbQ
6lJaOz6ZvLTTzE9YcyLOmYii3XjGroGh2uYtKVXorehqkL2BIEwuvMd+moN3aZggrJVDhcbawr9B
sFPnTpxrosx9XpzqVFmJnpiRdKxdk/mY+PoHPbWZpkSYpPcw5DhDlrYvMQDfu6O3mi8dHhvZjGda
ymhNloX0RizZrKA8Pkln69bTDst8l3g8B2dCkJPTqin+ljleSD5IIwHWwMFaEYVAzW0cyRwcv92c
xehjHq4POPmwTb2eTSuJytkxa2Qd3CcqqHuJ3I+B+GsWldf4s9Sgw3kt0ZDBsrqi9NjYf2EYVTDl
uRGyOI/FMXndZfXimHulzI0tLti/5IN/KJw5L2soL2b9sa/Iw4Fz4XpNqN6EVm8q58dOnIp0MRr4
w2DTdd4IKybJTJMPwqlC75gMHlRoAbp+X9lsAA3F8Nw1sx5YU4pqdwFMrID0eNZhRHgm0Ux+/ftC
QEfy+zlVkZJZOwfGpCM8sorCTKc+HkgqqVmy9vakybC4squ1k7nhAlsye8KXVFOuDF8Wgg6VZ9EE
olwSpNmymdNvOi0Q/eXTGWZ0ByVv9aJXEIEcDdEyvQeA6/CfHvOnyIZnQ1/dNA2AI/ZzjVgUauy7
8FrbaEIT4/MAyYFevy9nYd4QWOK7XJUqKYdF1SZ7fGFlr7UQl2VIUKf6AU3Am6hYsKjg6bEd9ajK
NJtwMQOYFHI6B3DKnNk1N5labKu6Qi0PXU2pX0g7++SGU09ePSCwVvcPEqsRolhqPOdnZHo7JqU/
q9JA68OMrsETi+38ixIRJ5U2OqVlNyBmMhqIFUH1z4RGuTE4kWeBDcXhpuaRTgs6vvUP9IAOj+KG
xzBsSNfExPYHZhJIz0eWLKC7Glq2vR08UuvRs6e7aEoZLPAfz3/UuwhIB++4FHBeend41tx0rAuk
J3kbRUTB0Ia7ZDTmx9yUvNFFExdL1TufadG72MrhOTMX5asorPyb5O5l1f11De9GfZ+pKqGPIuRa
zgmBbnLjST6kL/4H2ysYwnI3rJFvKYMwwUO9/h57s3rQ9t64CzqyMNBsexpj5D9Mnp/G/vkGHQOG
INj9WslDVAmACUGtwIFMwCWoGtxg2eMv9Ha4SmcFJ7T4azNsRRdo9Q9e9viTjB/dcZ+/mW6F6gHe
gvWUl8Ee6V1hNwOFNcvF3TNNxL2AN/EHRnQd1Toieu1wJeIxh5ilzGsIlPecMS0nQ+JHXY4ICGbQ
JdqS92JKZkY6m5wePl9N3eo3eQzfSkaNb47TBNciIb3x3szPurtxJEa64M9JWZhsuRusasxljvae
q7V7cpDRmKjv07t4F5j5vlYokiLXWlu4XWLMIlWvuCCpnfSL6ZHfJEUxr+6BFJ9zgwyHnXeK+rVQ
hAQD5eQk4fKSZDkDLnBaKLpZ51d/FkucOeZnLz8DkaFGmLOWBzFyTUqbo8YLmtWASwvgJupBf0Ed
8LE4MjLNuD48O2pJAQ4Mu9cZ4oTRaxgAjRl051+323GqiJaa4xsYmEMvq84/GfECzCgCf8CUflt3
CkLVmYJxi9uEnUX9446rUoJAT/W4tmvWA8ZV2oWpI8J4wzYB0kApSI/wzpsrUeQu4hAQ55BpEcG7
4ARPwAtcTdBamTMaqkhUwTSe8gyfnLVplISTTrIDrXfs0oiYnkykGeGRUp/SazlQ7RfSi8NRjCok
POehf8NBw5r7spfutgrwi0g+SmdIF7h5jq/PXedkENYUX77+k9XqKJESZK4zIfdrzEYBgjy7iVuj
oLMqlz7RO3PN4DolJFpoEbBqauiiGafWNKKZ0EX4PyxasCqkS0OwrdG802lQD58Wb3hWe8BSvZqH
KzqW/6kphv/mhc7CaYLpIOUGwO4l8G9nJzL8vCiuP2HVe4VM2WJUVBf2GlR30vrbOOY1DBvga+Jr
eb7KHjbMwxB54CKg+l3xwUrrpw8shaVFDWP7bZdIeZmSoObq1DZInD1Tye5PucWrHxnvbDkz4JQd
KL5Yf3Zlqav9CnjelNtYjheZhTDbiVbZSsjpIQYoxq02FB9xbKuuXc2qeJijzgibhGmwMep+hxqh
8ceLZQjrF9AIOzCjezw13aFJtLhSV87WXTJ5iqyPYQrMjRCp0zWgkt7e4t/LhnXhqfZH+ybJ3sjQ
niTci54Ofhv286Vv68uJTx3luHYqIZrCFGQbNhJoCQex6GhoaP6GtFQhS45YgoiYDL3sJWbulRN7
PHxWf1h3nLANXsEqo1aj0hMo4We7aWgIUQzry46tyaCAOvlQnqdvrbabQGGzGTJDIvcIi4cf7enD
YcJxXvT2U0vbx4O2SlCFtG44tEbb3VaCkIodn/5MhVfd6/4N9GaUZp5gr8xWi/hIwSd1quZvy4Gu
LSaOTvNeDYPCUJqrqs3ugmZrgKzawS4MVGMGIC6RRw4Qn6dTByJEQCKjWv1QD7RTwh8OrfPndloN
Ul/8GwkOzcJcSdHTkULO90jKTq94FWfK8yWl2/ho7k6kQv9Qd+JlNgoWHzUyWigBopKdYAutLIUQ
6/pJBsoVZpOihxaiuHTfF+1txxhPfGG0BaR1w+X7r8x7h0MkCd4l2SFWpVJ0zX5SY8iNGaxttOCy
Vv/Nb7qYzYuU54uwvcWVzInfsZgNYiXP3YtzuDGJyVIAb1665yhVxvKfD+alCSFQ59wYayHR3Q0M
nMI1GL9I5pny4J247yKbsBSbu1UBVksTIeyNKc0eIrMBEXq+qiUSjitk20kV9RhU9/oHcFQnjnJk
NCa7xY3B7nFGhSS19fygk7o1DiPD26BLTm4I1e/XdOx20XzbGRlJ4bLTmq69XJLzSed2gwWpl3yl
FhHyyvPZHFG7ICCQ+3UDlVcze+Y3w6kQXgKtlT2odZqsa3KIyLcodrAqwun+Zbk7QMZ7JtaTLHJS
wkqwbveYhsnLMXILm8NAWeCAM6Ykpg8ZpURVas+meKrHD+rN5wOQPvdx75AqLtjtwuwcIjqjBWR0
5b58i3AkldYkEQ5ni1EoDbUXKwUirovmLt2m/jSOzzIOXBFzBCq4wfq1bruS0+SOJgAOcljaW1+b
u1oRGpsNyGrYswh59nqqVQBj/P6og38UtDF6VOjP8IrZh8/Ka3OATF9yHfM0FImTDY63+chzTTtI
Z89casPSk5qLO8tCpT2jOyiPW9w96ciwnDn798wx3cnYOBMY4J/W2TzPUh7o7h1f0QbID8eVJITC
z6yMiJjOZ9r50xLjjZ1AKO5miHHAyeH+tS21zYJi+Tp2StT2n0ua4hSFycSPNZ732e56Ce2L1nnQ
0nvElsryog2mcwGQgKJKt8I1bz2MH+xRreDgABBrqIWObwPGNyG1X6a2AkEkK+Y2QFRm1dTTSWd9
EIlFd9KkudgL7hHDaYWUOV3SjVgCUFjO/DT7ZkjcQ60yKytIkEwBWbEzTvWW4KDtxq6+IQl4zSz4
BHiMqijU8Qwm7uyTbYurGiqpxR/tK7mQ9PRCkH0NKNF1jJ2XPIx+kk1PL7X9sLiuG5+iuwCar74R
xezOW8bNqzOum97zib0d7K+zT9ERsMYLP6eiLq71h/KrSXhxzIIsVRUyuqnCnIM8kIwHA+KWLrrF
xGssLyjdo255xs9ZjZqWUXNPYPmmE/lQrnYRWiVuTQEWWujtYpd8H2fSBTj5Oie0IHGz6j1kjP9x
KF9v3CrOKJfrYAdKVfUvDMAgCG71jZumGBBr+R2jdaRNl/kIMx5lE60WWRrPezAhfkL+yL3GBwKn
fR3sE/xRgEEhtstD1MR8JATRqJJ6qe07pw4688yBpvBlBFUUd0KceuLxvZLafURQYjrJo+Xxp2qV
N+M7+VU/Fx5RaEx5BlQTRnN6Amu+qRFu5RXcgJGqOM/FoVVHRi+wJDT5hj1pyL9wxmQ0gg9zR6Ir
O687pY5lmF3VGj7z0G3oMPz0DFWE7+4MTOZGp+g6dXDiDU4v4nZB3xynCaSVlw2bRCrnF2Fcdd6M
EK4/y4iWchjkgbnc55sHQgU1o2XFj4NIVnqDbDnOe+hi4sASGNyf5uHF9Mk6v3o/QiQoH1D9g/dm
fuH+XYHJyKqohEBmuVsAeNKFWZrViwdWC9QS2y1HlOEs6YpJfLl21S8Hc91UPAeN2G2fYwF2utwg
QU/A/q7l1r4L5VkBqRvIkdYsGjnZvf/EYGNtqCFuMGosgVtCFGka3x5erprZwnm4zZhbb0RbMUaE
ZeJMqQDxWMrSUGw/rcxfyXUnYl9/fH8V764a4BC0E4vu5myr6DGL1ddRWkMVPdRW/mS0yOGtn5JE
WbrSABsnGz/y007lHGHAmPN6XCNNAu8QpH/ny7/JhjiCGKoAMzpuGrUA8BBmzwutioNW8CtNSdMy
aXB10OnalKvCjjXwIQO4A2Q+b/FyuOcVdr8J4RJxk0pNvjicxDeQsElrTYOz6EwbauR2cwDa0MG0
pMy2rWS7aeEOGKl+d5r8f+lUrcGkxv89xB+Ov6C/JXReGbUXAOByOnU25JzgRVJnQIRIa8w7ycQ1
lohUE1JQOkfK0bSBC5RoubVOCGdon0UdcnDl8hOMXTSVFrj1DKMGhERjdTnAWEx5W1NNLlNYXD21
hFbvAhYxCfb6lElgWiLYtSUna8UfNcf/bHCzgzYC/ai/PtKBAOFjwq9qlnCtnOPdiSB2qYXewcb8
2JpqA9l+0BmoYn2sADaVT0jD1C836CuCRtfP9kcRAFRmtm0ZU3O1iM8ZPWxEkW5OsIxGOi9hZCua
F8q69pXFQQfoMeWrzty9de5iG554A+yuaiKTY+33/inLFFbC6orJFcBpFEKW4K8faO9EbqeSarjB
D7J49m5Wq46oftE2r5LBJWn69IUQOWZwQ2EiBiJKGhZkrxaVV+KcCX7TcV3IPABocHOPi0Wy8SmK
VL9ZQ7TBOMUuI93bxGMWzt91jKNwBcn7nzr3m//xbA+RYXIC2mcDawTeFwwWUmAi3aLSjM9pbNdv
p+4uEHH4MOWQEFyVIAbC39ZB+gUnAfgMDxItNIszSNFLQLqYCHy9QvMHE+kX3126b5uyRoMNdti1
iPU358kBnsxJlXCBmrMeQOsi4VwhetdK9YBzYFyZVeQZfEoy0Q20amxN0gTk/Z20394CPXA7HZfI
z063HHf5tujau+gkv9aZwJ+bneT6w8vTsyWsIhdvOX7ccAqkoEtiqeUX2b2u+OnJnQ5u29FzxLB3
qzWfyEb8aD5c0eGXvtcxOTekFnZaVHONM+ZYKW0RF9LFporfAHJl0kMZlkpOJjUcgcZYKolLFOpF
FsWLx1Acc2WQkUO80TwaW9WAILnqWCWpx/bV9NyhLjeFCbgkVSjctwJRwmJzk3jE6M0XS4+DvQYh
eO4FzDoym7Ik38PT60UmMIOFZCkcbPvbAgupl/L0NvLq7DdtsK1pPZcosmkd30ED6eFlCAikbLhi
Bs9h2WaRTTTSMY3c+ah+lcXPzV9CogWkQFedRQStJUNQaHoFAUu/ztnM26K5b/fyOj4YLfULcnoW
cG6sljEeNsHYmBUWt7RmJ+IbcDAD+5aJQYg9bOqVUdxTA17kMruVaKA3rSXaMJMIDpOlmQGqe2Up
J5OP2QdZUDeA2hbrDamgFF05Et+lM2DRBb3yTD1Fuowfti+tKow4T7YXpMjjd5PyHtNn6a3I5zjs
LMcfcZ+KDFcjBUQbInU5hE5tpX+1RAee4JpLQsJ43MABI63Twroet6bExdGc63HqMrY/9X6c4NTD
N6ReycZ1xVZ4ZnbyzHzsnQanmz95HeKcjDSbGeaSnIYDCeV8LJgJf2kyPdY4TnO4nfGj/lP5hpXn
Uv4Yp++uKKjhUtRpQp5dtqu65f4PeS7T4MLZuXPlb0FZFniDvipj3tUMD+H6AlFfNGT+4bYZsSpV
yCWX+iCdp7lyqWr/k0QmKI4PW6cZIfwQyDPYbJn4foMd44VAq2B1DAI7qfmr1S5Bzq6MnxDEeajd
C5rtTu86Bua4eK3BT973ZE88GDdRy0F7TwPTdPKtVN3/87UFpw9I7xPJRthpRLjJMgXiag4J40XK
6WQA70xtjIei2IIovbfJrsn/1bPgjYf63kzdbSkcTuX9fp2xsaQ6JjF60U7DXj5ae35YJxxMmZXk
CiO2gA0EM7c2fkyfnULSyi0rr7xh/Bf2heR5FN31Dyj8qfxC/kthc4p3Dw00AQTvC7lzXLdjL4s1
ZtCykyymj04NcfWgxQ8pd+zbp4OgUOxX+iGkbZsU4H11dlBMfSdEN+PTxDSV7so1P+K7yeowzffo
Dt/JP3IPcNYTTP09Q3MZv+Ucpkvy44Oyv0OfjB8SQbBzYutbor4B5Xswwb8T8IjY6H+FwnB0jOAd
fLcW8kK40lt2VCO6BBd8OXy9Smiy1PKqBbdEzSaPBf63hAa+8qDY6jNrpG5CRus6VFpcZnN6FJ9J
1BXlx2JfmcYyhGpqgc0HPhiENpy2uSUIKRaY5BV+rufKvhvTtfiM+YITPtObNBO1lMvTglqeBy50
08V1zJdLW0EYayOjkMge7pB/luAgMnIw+R8YlT82SGMzXWKftVpQvhxQW1z60KwW1VDv+/4sapJp
dEU2LbbXgVCR22fKsQ04SCBCPOu/cwwnxcnjHBhjOY7buwiGl1h9rlES9wk97rIMAZOyfujMroz9
0sY3JfUDACTzHqCpYZ4IEI8iyg/5lCJSrJotGdHnelj+kWWG8f35NOI67QZXTmuDUre6J65x3aWu
5iK6KNZ0Y43yQ6XOLpaudd7ikm83QxmvrEvhRlkbjzGfvM2/B4mXx/WBt5D/m9enR3Y/z0/NTJDC
SWWiOLcwgHo9G1WqeFe6o+I7h2qv04+xGKcN/qPwcxSfVCPEeVi3cEzvcc+azMcOxwfw8fKh3g1Y
hrkPpLlIKpsmMrPbqIk6B/VdEpuEtqEb2OV43vuuPHSNyeDy2FZIAANM1oRSHIB8TPLhKCav1C0/
nVarFIXHiLYIwFQsi3rfe8+iw+iGwXHtgpI4B6MdVdNweVWuz2wOxxsUNbjmCYQgGrOL19uL305/
9lbagWTzz1qi2Iae09pzh1f6hwpoW71bLHGRnQqLJXY+4mvyN6VGfa+MPAdrXpIjCl7Jw7e9vLZ9
mws+P4LLFhMIntA461+U1vJLjRNj3H/uYP+Ox/5mj4D0rRunJPCSfQI1RC8AiCwxzDNzygLOVRlI
Pom0yM1a4IwwG46wQtcU3HN+NsQBlt4N7pWl5bK1YoVEtZ8cwud2qm7Fi8wJs1zPBIHw7JMrOBuo
9UO3teqcMi+mAaeC8Qr8EhFml1FApUU881LLtWILz5BnvfUHbo5pkCTd41DKW5vfCABL/jcmQtH3
UClt+xAsdURgaCiRzMdcQv42VrrMGGrAvmAvn78SsZ27EP+qTvyO9//GXhmID0V8E7t/9EhdA8r7
Pgt8yl+g9afcWAsjRQJWWX6VimT3PKPdmzCsTe0dJKQAmizavvMBaLOHDhGWE0cfZSyXwASMHcz5
kg2xkqH/KoDkZsIxJwzYKF3AtC3tvgN83RVA0roxWsHchfTERP1YDNpu6qzkInDw8LJnTkE+zzuP
ihZCIomQRQeyrIm3OMwcLRIuvfCkFIlIt4DnB7M+hCbARdM/ESwHWFi1DNAWhHfEMCFJTICRnp/u
4GJcP2YBBPm1v2RH8+Opi6CW2yzRyPVuCCZVC6wBbiuWv1rlfArnRfLyTn9fkY/jnD0U3ukDxAjb
+lx59N+qnQE5fY1feShmpF7AheMnAoTQrYUehBBoCViT8iWBuUYr60BsbOmGnoa9c6D49vs3/sH/
/wEK5wJ1t03lk/pqyAJgWQw219GxmxfVrP6sWlRwISuT9TIbOjHgMSoYYvid6WtN1m8ICHBK5IaO
APhBVI60eB6B5KtFLZ4i6RqZdtVs9VyXwRdmnJQLX9keWfsuBjFMVPY9A8bnwQl3JEAcAEH+UdyB
zGw5578beH1CMSrxbMWFZTL1XcazMaDH6OhR/F3m2chQVkCnHFCt7Z7MnQ/DofddXNCg3fWqeW24
A9eF/easdPxehXUS5THxrxQYOIOr0TJwea/6qfYSSJLTcD3BN8jmhmZT4rtXZ6fpadCjbjlrzxLt
lcWtnHgfuKHueuBtl7JVCuZDZYNtADgdcUyvbdm+GwTWboz1i/i/ZxuFC5uBF2QMEiqEObsppwRi
3nZ3VAOeJ/8Dh/bHa0I9HUymzi3hyPgv6LESIhXaP8FLNMu8WsJQfG5GIjThf+xWiqMlnUOY0TxQ
hmVnThB8KDghSD1wQKDNcyjj8dUbLMEzMG8i0Te/9TxhdhpdekrehNtxfURQ372i0iXCiY8MpOMm
nUiY62Uaq/BuER/8Fx4uWu9mYu9IW85Xn1hBhYQsqdqqfNbxmgOUuJLQ531WQITDS5l9IqtsfbDI
8KNao3UMtqrDxwerYPBoccQwyRoP8jNScLyIZGgDSYLBYvuclAcN8ne1guIIEftS95qCUBerpm7z
6XYTvKAo6efJqRZyE+zf1OMY8jPkrxqxeUCr1aDwdEPl0+Dy6b2pe/MjUc1dSJZHIY24jVgfnb5W
n61VxKIdX5kF/g4PKfHtU8pAY74OGxdCEyFJxeBjRqah9VWboqj0e7rcaR53Sqt92g5fOnAn/Xlf
MDgtkHjrpYqwG4pVwmS/v6nv9IHRNHxwFkeOLh5j89gVtcG+VWJS7aIR2MS8m01hcbfNfXOmZGIj
jhPTzNBm+5lIp137dOWnL43MEBknm+QJZAY0ZBPVOcqpSkjH3RQjHa9pYW63kKSNCus1SKrh3zol
ZtB/wL7GpLEHt3i0VJ6JqSc4Yf6WtR5p1DiO8nBeSRDJIezIW9SQa8E/E+tDkD5xPVfH8eWfgFt3
AS/hkQoAmiiuE7FBKbyZudZZ4t0hV6369q66tZGZE2Z1R24OOXLKy98R5EbaylfGhKjIP5bzuOzP
3DII8ItUnwF1WD3E/U8vOXvH1yMlKcgoE7eipVoqzF0Cs/fKfWWEGsMN1m8Hy7NvsM5V+W6+fUBf
Nnp54EJD9lanESwuEJ4gJuClwApZp59JqMw8VFq5bRnhr9XnBxCNM1oTVqV8kPIauq/Dn+WxLNTa
nIchJjBI+hoLnsEVR8zQwZXdszeZ+RF3KGDlsizmI4LNaG43kRoaD2D3B1ASlcyfndVxL8OHyMbc
JcqBxp24p260aWMyaBEa/WQ0Q27cr+WoSol2htX52JgIjgfqw1++qyeiLprwzACx6Yq8U4ChNMOm
R+Y9+S1Wv2H9vCD/PR2/veehyK1ha4PDxuJRJl8boogvR962JLMrThokjsuUcp8OkR+E4FQDSbwu
JYacpjBOABvaY8uYSQ0f4RV6bfbAa0U4XP8C58r7LQIOozyTDoM+pJGerdTJ/q0Z0l7R2b9Et9sp
Zb2c+FWi4gLANJQx55+cD52tcV782GSFqWQ/s784OckQCrF9LDjz0pPThefN7hsWrvntAXrSBnqy
TtyMycwzBeFaEyA5NJMMF3nbP7yPw6j4AqrHkn8Y/YpBLUqtBfdPXBA9vF/fZDSCN+G0UU2Btw8Y
hX6iHSLMVlbEydXhD8txCDWI8t1n6Ybpb6YpZjpOJbM9QIQmKK7TH+X9KqT8eHovc6ML/xJRmIqJ
GsmGNZNd+PeLTbGbaQou32ITkVwxf4NpiYE1nfp/VAhFdKFqxU7gJkgjsGTSqe53+SGyXJ79v0uk
7gC2rZq1ccLXe0zhnaGYVejACQIdUsXmPsRTuuGfiY9L5qrR2YLQxQX9aFzoKVYhYmV9BRnSUZsb
LTKSeTkExljH9WWvLCnRR5uzKXeUVLk8aPgBl8aamq+ogbcPpOVBzsZIk/qujNPIdpFkoeKE2ali
D059wqZpzOrOgsH4Uet1uMsDy8Z3eIHIAMhwmHglFp1mI0VpXWkXfyjoQZcS3UXCYj9TPri/1QR4
0Uz2s5JUiFs3NJ3Mr0LxuXmxq+uVxsnRBZP6b8AKjRRpd5sxz8ZGH9luB8y74tCf51l+A+zNZTV7
BSu0tqoKBVgqcBbr8CzefSpNvsnF0hWpg5GCk6u4YpY1vssTJp/E6JYYZafeGJG7BANNwYGJ3jvp
x1JaqJTDZd2VhMgiZiXqc5e0biCtxyjLDldzBtlDaPHYrrCJ3NhNUdGvBCep+rAc470Oi+3m
`protect end_protected
