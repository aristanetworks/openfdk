--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
dk1nLNEdHApdpIKi8hZBHd6sg5Wo7XfeseLqYDBfZ+Ad/VN3ULQj12DHoAawqRVA9jE2hXEbQefj
t/QKE8mjJo14fbWgyJmDXjtPVGk/JyVzklqPwkOVgs47Z0O2+o6pDPYBTO8IS2ptaFEV8Ppgwqtg
cZg800EFJg15TCZjYMiQuzTVXrxo0e1z5a8TInNihsQFp+VzSP6oNz81/UJ7+E4rSA6kfj6FWK1m
1mD2pBMFCmOOCNRRiegAZe5nJfuF0/VGVp8yrwTZ6ZdGA0246hQMSXDsx42BN7enXmHVhfzpUPME
cUgtyh04Ttg0CKzBejLNGtj7/0+WoQh/c1nLAQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="xtuaNMqFeNZ9DlXHi20seu7d4Y7NiSRaWuLkXhetcjA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
DuAksg3LKF3eh2pRSCrtkktSKJ8j90xqgzk5SDCo9yJ37mqO2Z2JiZyxH/E5jFz17Py6L1tAiREl
VmMyGaiE0JhR2szGTzviNoWRO9KY/YQ+FFgjtZDID97J40tr/nHAaBMlMjjwkn9zvorEOICgOPK9
/6XFx3oaXsMgCOULvXzRDKhSHTimXlWCZibYe5bzJDJGwAuUrVeYat59q57ZbJcPJqimW0ZxeWIR
o9APXUbNikkro+0lP19MZIhxa6zhj72r5cb0L+J9HHadYmrn+90TQTcMV1/t/yYVfhK4OALxMz4b
8Z0JJpP+NVwWsuOe9oqaPAlC+RVrB4lBmIKnjg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="UrZo1L/cme1mGFP8s7PVguVTCCBOo5qBc/IgLpxEd6I="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10592)
`protect data_block
TyjEwOiacPNHkwMFPaFW9DalQ8fCEylDbg0Ont9ReGEAvAEnrxS8CZWEM4vRE8zDRJ6w43FvlD9M
B4XsMW5G/umXYELC/gPrHW0uBDeKcVsjsMKkPJ23T7zA+zVfRJXMj3svhiudB0M5Plx2qjpyXF+l
jGQzjITPo4HS0b2gNmn9uhhwwW06a22rnZtwg3KMpJl9JRT/m27e7MfmP3zbHeNQKgyQB+0v6zTk
j13wFfABYbM/Vc1aOjI+ByiUR+rG7afGgdc2hhmQWG7IiaHaX6kX4XfCAO64hP9wJVaHPZAylKR/
E37zELC0KF6JfgJjQEwF7pG1mPQ2ZWeW3XKltXjmXpn2t/1QOgE2Ar9KoAcU1JTTCVta9hQJp+vO
DlMgncwVfi2hO2XcuBrEP2H10YLIRZBO8HPptPYDuGtugwSQjkxhKdLbAKdY0cDTCXrB0wfC2DL8
tGLcJSQVKUxDXDvCw6FnSk30Ul7stgTS5KchGBwkugqZrrGl3MzrI7i2UFVhP2oxJQsvmrCJW+5c
whtU7pmIn4BJtZ2YZdirhdddHOjkUSqOiVq3goaRN4yzYy9U/pAOYQi/Hhpz0UcxDsblPb7LU7jr
6Y/YuE005g9/cTufSoNptMg/tZD0eiqqIAsqPXupeUD0Re0zt+p0oDFP4sI2sE16YE7En38B1/ME
6UPlb4n97n2vn9VGPZZc6XRoDLuInQXlfWCtC8zCnLANlQNuFINNds5/SgeIvAkTrWb4rb3Driue
oziU7vYcdOTpDJcAwUwa4TYSbq+JB8EA1OCtVGBLo/GUndi2GfEn32QYODci40t7V5i6f8wtB9Ye
lEVq9oAjHp1bBOEFwZ0VFa5QkYifVYghPulyZzhuMoI6GZVxodLZyOM3f/4fzvRJ1OxXGoOM7tg1
hnd4M16deZlTaMbdWp5SjNyhTdlCMn5eedK4pVoNdkmrL5dTzyfSBbV+riRDsuvJRq9Z/6GQ6Lom
u4RxeLcN5UJH8SpeSZl99cQRBE7oSX3lVTsW/+EXQJIFamFiHS+KwJ3dHg9aZB8Blcy4vwUkaFJ6
lbgvbeeRrIAhWEzUfMSVImjCKk1z/s0P6FEkm+HH/kstyb4igQG5A1SVb1bbWI/nIegUic3TQJdC
6hHVMlWpn6J2h3dlb6Rk7emOPgLtB16RAYnitQ2F6a+8/ntinL+Y9kV+SlU00AYlBZaKWlBe1y3/
L1cuNXcDCmvN0Dmn2Qtaag4yuwB45SFC/eQcinUvYAgTQ3ncMwRQpeeBT5IASBSF+Gsp2FMcmvbX
HAW8VqSTaDCCOSx9Qt/PVxmNBF3xwXnZXjU8XiSVQ2dIEnSiWufhoJXXwDQo/kbWOy80Dcugr9nA
C7I3meq09w1DILb0P7wrtZFqD4hNA5bK6q6cVPD7UjlBwvqaMo/puQ8npUo+WaktiX/FEcY4q8li
txjbq+4ZIbpgu2sYhm2GrrDWS8s1B4AQKU2RbzYDqRt1/9yjeyf9oQFy92Wp2RYCZypYPEuwvDuD
vgDrJFT84niozGi9m0fZqqoCAnLLjZrGweQfj6ZN+nDTfu4ZGScNuUeivYTdoo9d750cVdXCkOU3
22LAqMCyhJqbmSlNqc/BPnvB5WrRbC/9T5fpQCtPvrvxbmzMnYLg9+3zIeqQK5OQA01PO+H9nEgM
JNAEvwllr6j2Vu0oKH4WvKCKi70a62JOyusvSENULjBASejMbbsuaFg+5uIcbYsmSM8FRbAASX3G
SwkgSBjIOcZlp5kY5Fysq252GrAfS578G6fOCa9Nm9qPUMZafwub7z/RT8Y9UBetnKPWD7hpL2o/
afPTQTxMU1fDOOzkp9UVlJ15H5+FJEe5U3esYmo/orcZ6fFCFnsmIxo9rVy9dCRaQSfIAhcPTDjM
Lwt53jse/xw0Wck2yGLbI+BwxgT/fS796NKRbDpvdjjrttnN6LZGWaPZrPOonH/H0c0zr4KlLGvN
sGIp5b8fuzeJ3sCG9BxsmTp5s/TJo3j7TeO0lPhsc7uWLZjnfl+6rwpClHFgjwlml5qtycMTG/aT
8Y7f88C1KZQkpd7a4ZcEWcaynwhVwqwsjhr7ApLtUmh8+wJurMO8T6VBlyy3ksPHC46QeERrfyh1
yt+y7oF6vMt7fmHmegKoZF8T+xwotOrh/XIeumYUjWUCkLXn/GftnugUP30ry0BF5OqZl6OEz514
Z+k571usjKQNUsqgAve/usKiM/8BAKNeiKvB30CrPIwFtu+x8usI9pKXA6ZYuiUbLhlWHOWs6TWa
PVJ1nxT6k3tHkbIcuKICjglcKFa5MZSjC5TUhZYy6a6bSoytcUJ5FXMYXorP5FFOm6fkwvRIDByK
P2GT6ud8z3KpjefayaGzqmKffz5unzy9wqaRDhVAMzUhNYeS+fWlpWrAp5eHSxa/q3GzlJ0zt7q2
qUpAVwWqnCWrz60OIenesRQgXFTJOWPJXANkNBVcfBhwVt4BsN2QYzhE/Cdnsi6w1gu4g9GUg3hS
5zp4Ncoz33nEg46k5pxRuC+2MXwoR1bqr/DHQRh/JEM0nHz6eoU7ZSIDZ9ZZ0nRhat41dgJ0D06H
VmxuprRadE5F+qtr5qCGfWFLpgswb2g3pw3c/oiE+U2fOLXqmtnSYwGUH8fd7pedTNph68t/tIbv
HhSPZZkLzi7uXr156WQkMmTQUZJKZ6FIjv2bv6x3ZBwKjZMt8aGWHhnzu2fV4l5AmxCo9p4ZhBDj
0KDK3tougifikD5SCG/XY87+tp8C1xr2RFW8TjpVO8J8OxqqhJde0k5fvCjVzGS03zTmoI4NW8P+
3o8jf+Wejo+lsQdZOnwYzIzFMUiXWhrI/giOmYSHVTp7q1U6lotUSTKMhjjRMShloiZNH2/tyY0e
tEsGvgOgYHygKP4Ja4xC5JG1m1OzczkDZ2WZFSRxmf1SC6w+vaIzINK8kKEmSY+ytmitQLEwgf9h
+VwzNVTYVkw3acYiPz0mHwHQsWwJ5s0YF6bGRGySwphRgzI7CK5q1NQgtCaVyi3xL65rnFPCSy6B
IYeE7thloAu4tUqCStQPp5LpQb/2kjzcUkBnbEFU7o/9IZtIMJdMzlQ+prxoq/IzzWphqmJ27i/x
LKrU8SZ0Vj/HrgfgLSdNm6rRdwz9K3VidOj6f61JA7oA7+ZPShYh7cRfKJZjkk88b5dKf3m0mjpT
ntZEz3SL8lZpjeuOS1I8yFmCAhtzramCJfK5igPs9nkbRwVC3FyIzh7aK96puFerzIM6W8/NHSA+
XXwaaWSFO49CJL6iRiebaNelK/odX26Q3S4m2F/pdiuy2jSj/gQNzNNK266NkiSImQDsX7FoMiB1
oNWYEX84fWPT5w6x+0k1s774yZgEXr4SwD2NjaQf4OolA27ymocYnx4nGQuH4isnvnmOPOaixBiE
eFd80Zk3OLnqher0wiBnhzr73RIWdOlXCn5o/x1ChErRa81eyt/1b55o15dLMMOIx1YzZolF4k35
qt7ggn01jPMmAjSIHtVROnRvJXYyTz5UKAeenQKvtD3LqpHClSp9w178haK+vHo0s7jMmUVGM2q2
QWAvZXu83m5y/xcRE8LeaSsioLLDosqGeryE+In8QhUubrlN2+Clxiinux9vudpXb6lQOFNDlwYL
LcrBWsUkmXkINVlABOQ2cQj0pcPC3TcSQ5Uud+PfgeDRnVHjPxkbLr9n/KAqGrXVaFNRP5LG6P2g
wmfyTkIKxhsO4GJmrlAdYrN4HNGn5Rzxvk5CR9bDktcyMDuBelOE1kcHOHkRXdiWBCV0am2awB5w
UIK3Klsma/uh1UC0blocaV1LlXyz7rP7ivqZ6DDt5+IfcZZ8La0+a92Bzz1tscuKntwiwl7knlnA
F0TEyNP5MMbT2/0rPsVFSKw9iGg+zn83WTJrVbmerDECqi2Ghcmc1C1HOBwTVsuKIGgzRx4CDQQe
gy/v+GB3BARKTUrDkNnBBSvpJlweyXzHBs1FxEqo7DYrLQqxw9dtpVpklvJofniSE44a1ouNg3dp
AbMcfvjwg+u5DIufzDENha4JOvdpDhg/YPpJO20+Os7hjzS+RCBPKXhA99r+nfCaoaFdbz0SoQPd
e1tOVH0Rxv1oMfnqHaO0Qh1EN7I7x+YQDy40vlAZlzGNDqIz8hW+69TuvOOxPC8rLJXHxhkF+zwT
RYHdGhSprfeS4asXiA+T58uaiJY32glm0lvUzBvRgsSYIMxsxUrJUdbae2YW71xCG/J0hSQz+MwO
RssvHKoi3MzoMz1M3PPXaPJ1J7cqGrfCzV3knv4So1wmUcT6nRpyFYltxEYRkgVLfWePysjFTUrz
XnxLkECThVnRdFVSv7QYgkpdzM/Tg0ZrOqIrro32ZHORy5UWyAeIgNwe5xjClLYDzeCzknMV20FS
uFkj7ubejLlDuxKeHcbD56dEzld22KgDLtzwDYX2fx1gzPNCRF4+JbmLacY91mOua9SlSAlyyDR4
e844JvhZ+WG+Y/Hcpo2+04Z9gzJKrrvSIIs+bZWpYOxfqmwNZ+qlIdXd5Llh9OnbFvgiONuxYHFm
JAMN//Sz5LHN9F6fE+DieWbduwTT5krkNhS4Eburjn936qo0A+WRixpGfBYwNL6upBR7K7m/fXlz
gOBtVi6+SdXffj8B7rQ/lwJY9qUzpKLZ/y9TUP9rJgNipMHtY+zOjX5paNCwqDXw3OiA8RccUTht
q57kmeiBJOIVHAB18qofyeLvh4xMdHbzPBKeXOxqMJit74ekKuYU08lnrkXmHkKgf7cEu6Tf025P
jTO4iMYkPFSkua6DORQ1AgXCGhPJSdHclkRjTSuCh6ND0cmXjZy0+YNvotNEiF8joOtADVydyVhH
bbMOzIlCLpZWCUCDGUFJkh7HF5+sVyjFYycK2M8aAOc/IrhKB7v4LjaXewFcxGTuHRWJC/y/EQEn
vbhsUpG9OUNhLiaFCrOjfJ+OFAog1P9yrd+uT2fPYk/EW7aeZIMq9d3ie5qdMFbdLFokDJ7c8c9H
UyvmmurjwS9SENUWONYrczrFNUdHmmZmVMhyVwMCDL1kI85FnJMKpv0Duy8+bJ3MsPdqBoRD3o4X
k3EkaOgLeslgFo7yhCwuhB4M+7KtaBhIay5lAGL7YYrDNMToeF0cx6w13h14HE++w+yG7ZgAoemg
TZzUUxBD94uLfw0YcoOEjx1RYuTFJJ+oBG16Rwvpjf+TksNHfPh7pjhX6jAOB/B12UzKlkWjaSJn
8J4w6o4K1u9Sh6vpwn3k/qD3qBae9i7PwvPb+QeR+CYM17cVy+8NFGnnkZnbkbQXRXknhPNYOnYs
Pis9PmFy/WODvbkEJJE9ahbszwbU75CsZ0tTMmNyFXxWE9ZOs3jUFgXozlS8zubRP0AVHAeid3+P
5Vy/g+aMQc+J8Q+990sgXsE/V2458Hj2FnTb5Qx/PCuI+HgO0+d7oyXyLOso5xFPXDGcS37lNt29
FKJ/YbYfmXH/ZuE0emyWuE6Cdg8iu5ibU0iJCgbv/wJaoBgdG+RTto1cIwEnPPivdtK/AwiTBkYN
QMafeSchY3ZFkemf+nBJ/7cd5iJ0i93qqE8qZf0L+yLkysuEl4YE0c0+QZuCqbMDsv/11ONIgZmN
IITqvzC+k1nqoXSpjUpPZiTt2SDxvbD7/a5GfeLawtI9EvIva7kfcT7VNz8/LujLBvCbF/JjIJlq
+XUeYGnLzQpQR181SDOq+cWjcpCqWoPT51y9VTGPHQzb1gsTdc6CLSyBPnzHcOeyTtNzkWzxbWHE
HsU2NofIu4ShoXuccv3As0zJy8YFK1ZkPiVsHcJw52sE+UOHh7Sovkjtt0VsByk9cXkLVlkyCoj/
5aiUmrBAVoONbDDDIKE9hXax45YhdVu0c73WygsYB0s+BaIb/c9uVh632rBY/M0RGPGlr9HJPYz5
VYzvLQ5NF7ratXatX+DmkP3Iv5a/UddAj2aISJ2ClZnFUHOAFIGzNIO/G3JPM+R6jXYDg5o+Cj1H
PUhhHUyf4s347PmVSivgxzW5XY6gGoWXjvO3Pcq0ngI3z097tbFKN18irh+H1zHX0RSq0vorwxpW
JVJaKf8vnEMCqETVTbVTEKMX76cN/IOWM2jc55qQYUsBfgKCAiaUYu634uI8jtSgFXh21+Jqn8g1
Og/HgSp/wq+rB7gtqp8EgHv33dZlX+GQRl1OsJ2xTN1OYSh2zdbjFKlua3qbrm26j5I1pgDJrKD3
oonkCZ6sMuppvlYCYLED7d++LDN5L4J9AM1O8rLwhEQ9Z7nDyP+K7Qum/A3+WWljm8MhgxoLOaeg
SpxW5rTWGVS1k2uSW9xQAdvwwsPTBjlrCzMajsAQ8d2IbfjAq6XAn6niOj2j4qKRRzJTtQqcafas
R4rzTFYpna2DkRGIuQfckJ8fscdUWeSQB9jME4lKQcO7u3Q71lXH4FFlgqxNEtWX7KmRz5lCEzaO
CttM5K0bHwQyf6S5I72JyoIjlCjICb7BJsI2ZUust2RiYaKmCo/yKuC7+2Mw703+DX9iSymEvVji
9LpaH3uhKhlqvgWvrnNqcn8Aq3wIjW46h8wcQDLHArBgaY0Fsv0IT93bdnuYosw3aHJETBEqu3wQ
xE82qcu5R8wuF3wAtAPRwX8P0BCt45bVugO2ssZK6slRuZIP/RTcJX0QNSY+d5ZECLxXdf0RuiCQ
Ln20onYU0cYY5zzAz6ao6x6E0VmKxOMYSAhW0pMCR7Dzl8Gm9Bcc8sWLiqWXX/76lnFkG3ZR8jOy
f90YnLRwbuzI/CrBpQrOMSktSRVqeXVkpCS8zzeOx3tCtSG7YuOmo7UaBzJuk4Hnz65AzaAKOfxB
1G4B7fcZjQn/fJ9VM6eR0JhlJzkJn252vYShKvuyQ542E5nYBXkjX13E4ZtLXrPvT544e78KDwq3
uqUv7MfoILwNjl/CDCqvwoEQHPNirr6GiWoNUJHFnuayg+0E/pczL6VaeSf5MlNRGzmWMETjsor7
e3l232LdEC11mFrKAXNWecdq4bXlnFy6FRmmFFkQTl+VKF2ooqmeheJ82x9fAtlXgoJJblR9ZgrG
h4ucJL1mS0TicddqOTVvkyowJysaPernfQTajjwW7nAMK96Ih+XgZqymMH6dws+Mt9fEDR5/wHue
Nz4w0TEJunDPtAY8StUNcOMmkXF3rniFfc/QvN5UCRYBpAc8pZDCuNHLLg9qCSsv5Z6uzfvrBM66
KhrvwMaQep7MViwDa0w1P6F3V79Wp9Ts/eUJqdgh0hZtIyA080+SVipYguvF6zXNEdCcACsSJ6/Z
lL2wIuNDCSysUszVc73TO7nDkx4723DGA4o4jrNYzHlMfAB2PPwAtHJyx4lFcqJcTJh0DaDPaJZ0
DVbkmwyk3uUTjsHCXJZxJ+i4/rfnyfaD1zsf2GFwyi/sPHNE0ymAnV0Y4+c9Z9RKTQoXCoFecMIB
PwXJx9LkI3YT5q8VamCJVukkCWYMEgu5Gt/V4sVlhMFSeAqMw3jInXJeEhRJtzkEWFSMrG0cz6Ce
bX21B+gggPW+P2O9/pXt+qH1DcsEQzNP4tm+rQCZukxTXUKvHHUhlbLR2jVv54ZI/8JQGDK7PcO5
brO/dobXL13KuR9IXpfogeFHB+ZhUxRSjCEBOBMlfyt8Wuex7PYMx9RsPcx06inEPRJIZQQrqOHd
/ue4iAYW6d3cXa6dorZn00VeGSEj3KPm4hO8Punnb2Rk56yHR9erG8EgnueXoG65wy61+/8ahEoX
dWKB6GzA250J2S7vxELxrL4aYIjVqzq4DjEIyM3egS1nrAcQlccUezO8a9DExLUV2wwPGKCmigcp
bqadD33UeWyS+wFaMGBmw8DDqJWajJCro5vz8OVVDqZ2u4aiv5nk8EYfsqSpeAqQGeJqQb2sBpEL
oK2f+etHYmBzIGYfM+gagyMqHBCa1lhMhVUGlMRHNTVRYKEc6KjsI8oA3oYC5jh8QvnxMjFXPq4F
0v4EYCCVas9KpCaI05zRSo28QnmibPKq9fT6VjpdEyNGSVVwpYMkk+wqdgy9mlQOHkl4tsXaXfEe
udFfSkHqpBA06hCqY/iPzgnOaEAcpqfONfwGfcPVPLgAMeJmj0NI8uoUsK6lm0JzYcuJzgfrjd7H
w/NWAsYQ9z81dn3dIjSKjL/xpmPyRHdDGMXsXpQShI7U/kuHE41WC+grDMivRn0f1wykmSkftT3M
WhsWh8FCegriWFpdF+ubrpqsEjIhIhcqBbnLGnoEBG4dhG/617Xfjyap9OuJ9pJbouHkCEKuqOkx
6+2l5HJmocu8O1dpyqYHcq/CoVfLS0e8QGtSu83jiSpU68oP1/BkUImUb7Xgt9QgDDHNpdGr7fq5
zUq8lkva9SpRPS7PfDkk8+rPrEM0I1vOgEFnY/rByNKQHmYpljQgMmxzUucLkAAkkRxjA9tSYIyU
IsgZhqRqr5YxAJsfxRBctfZrk4nwb8KpPvncHTA9WtcTit5FOHXOREjGI7Y2AfRERwS5wpW/y6Re
Zv5mH3s4GRHCJELmUI5rBQNii9gQaW3nsAgJfKiJZTEdQH9tuTnx2hcZYHweFsZ+4DnHFx4hG10K
0+sWxvprD7MSjv1zMyZeaM4UtATfqSqzZps4RsXw4Vi4dP2kW8RvSFthhZa+NojRZJsDtdfWyIeW
32Pj+V4oXotYbb8M57e5TIxv7rmwJhaLM73cnZad+JbLYq1X9zD0ESwVhELZEBBatzWN4x6/xGVb
rZf+GE57bVTFoHQxQEPLhWP63VDoHIY7NUig7oBpDdZquOjdGSVhT5mbY1UKjfLoHH6Fv/h4waZg
Q8ohwdBrluTxo4UYExocT0EBlXKIWgZLf+VKIPzJmz0mJSKHLUW552I1qTV7k8JizU5fNwi06AIp
a9bOHuOuan18dg89la+ZnXeAOtUwco8invBCsXkoUH849xj6RRn/mV3Iy90R7GLQaHw6Qzzn/+cV
bvjmflzvJOCMpxcHffSGFEqy+wLsOs9EkuBCwmHQir/LmeFMx9xfrqghyyjg+r2UESXIqY02CEOK
RgIoCcoPRrgFMGAaHoB7h2ipIGALa/rNClrQy9m+3Xakb8y+qLwrJgBxZ599NxpCuUoFCCHVnAHk
oRnq5GqZEqeP/+sqCBIzGr/YCaE+Fa7mn9mmrQs5cdeD7ZMl/dlAEOVJaoC4BzTlwHQQ1BW5Mlm+
z5aeRj8Z/JoCtF0MipSmTL0Egeqvjnls5VKeP8OXU1a8T47blXtFTkE8vQAqKGUO+V/RFAH5uAnd
McZIVzW/EZsb9usSi42gvxICgkA/VIVGXvhcEyJaBOra/vqNWWbUuYn9QHPIZV7rqp3CA94t0SUt
6lWD4eYTlnRMP53xvEiSH5bcqk5uEn13UyYkvr/MUoG92w/r1TIors1rSjLP7afGQV0smKUGjRjo
uL9DtqdoTTGfDmEtzHIIgU5Pxlr76BN7zo/CRCnjj+/QdoKJLq+MGQSjHxSjj7bLAur4Kx2VBwf1
ZAVnZoZ8RaINSiogKkWKkdFfJUpICB8cfxW+PBMSEvSNFSezYC62K5dzx+BCMa2Jg1S65BqBTQDe
Wl/wP5ZZujfI6wEBzRft5wygfAYNRBQyNVVkljhaIItIu7BQ99ry/ngZoguGXNsugJWtMzMlZSJ5
EMxxWx1/4nprO9J/OkXC0hYgTL9/A7MF4QlSMt5dD8CbzGv304N3CEdryIfOc2VGHgMtB4DO25Cx
V8EWdP5kWmq/4xP3Ougsudu6aWmHA54iq0ty0nL5B19Tfs38hlCutQTM91hbzblScWNXfwF+0tof
9wwYD83aD5vWCCMC2iDl0PxwoRZpxV5jtBOJslRXuOJTjvD3Cg4Teiu+iyF0xIYmZKSzedeJnhKi
Y0vhm1xUDxT478hfEHyma7b7p/dg8Pw1nGnaE+pWFF53oOyfGmkblC22SQPN13oOfjbr2OsuobIm
84563q6uZ4B36M27WniSk69DvLe1holDHRNJr5zTB+mmgyomF0PF/EpmAGlasp4A5EZBt/iPsMSa
6Ld+VlHbr1PSINAa6yVfySQlAEkyQtXzB8d+tuRBnId0ur/YyBE6hceobstLhThqvyMXDu5cyrDL
AdCnTXHJ+ZrcEm8utaQgH1d2hFxZP6VzPH8eqEWzFa/rfEYUKznTbwsGq/Yah0cy3if63FhfCUi0
lsjVjB7YKFETR7oqx+2OaqJXPVv/BZgU1iZvKdLHLuwg2RvGZztIGNr1yj4xFQ9xvKBTXeoH/e3E
N/X5m4iCrQQys7ZYK6OtMKPkJwfCaI9Po7O67VminGfUL/iVHOiPtnC1UKzMb7Ly6u5VIvQCzWNM
vHB7FyOrsAu54qkM/0jyfkJfxi5k+aQGTYU5s2Ch8TL/XjmTljbPDVNvpFMZQBEDEGy6jzy/ON1j
Bgb3WEI/SyWB1zkfZlKwMW85w6EPGMhlRyV31ZepIMZlZSIdCOpaaYx0uylorzH78AK63E+zIqsI
dAOamN1L7eh1KwEjuROP22hjpL8hyjJoSLwTkcvlSvBMSYM8J/DL9OoDunctZ44HVbitNLNh1Y+W
2oODZiHj+qW+XtSXKFcES1ir3wElT9eRLkLqBqi/WCcE3hfhKJF74NlQSb6phl6rDdfjlHfifAFu
hQ6A8pDmeix839UzGqb51Ci7Azi7BBJnALKBgBFWhMxhRGmXlcyg9afrqdlK+1LgSNZz6FwiBmsd
leRqYpHoChozCUBw/5C3WDntnTGZbik4W28Zhl+qQa7oGyi16T+wuTxpDgBXrZdK/IbBq9ShluPj
VVNKPvSpdVbsA7Qn3jhZNEAYY339r3lUsVs6sR1qOqK0o8nJHAYgORO8JapbRjETTIHYhQf6v38r
fcJ/bfM5CuCo5xs+KKqmRyKmVil8RU+f/2jjXq2gZ2mdyyHbZfLZJOWAmjFnqz1buc78WsUw8FI4
cVLcpSWWYd0SOPajMHoksTaYdmETWXBlUED0QEYH4BEBGI9YIJQkLIlUu+vUCbdr5ZhzB5u2pWeI
xn2pW2Pm/71DBjrPiJJ5/62R2GFurJd9eXNjqNM21I+6cNkLPqOqGZzegfH/naWOVv35ekm0X7Oa
s4bwvHfd/AlJG/rtxD14KkUjEEf4+KaGqherTXkoYmplt99XftxAeGdgUnOQsCmvkf0sScjyGGJH
VVFexRExoiW/ZB0EmAQfz2rrTG5y1ISZQwL/v4sF+MxaLdCcGhnJgntZO1sXlKRkuqU5kTkTPSxV
0Ygr3FfNTvM84rnAFmhZaC2rJLdYuYq0eyj9lkZ43Iu8WI30tzSKX43OB8Z/wYNwjiwXT8W4j5Jj
AXS6Zhf+yd4vlpJRd7gxMRpIuiaoEwQpwQ/+Sh/Mbp1HAjGX70XYzmkeOKerM3AjBr5DX8MGRPNS
v4vCWMhvBrsRBBI+f+9zgkR43H8GlrUdYCZ0J0AkfFpqRPUfqis4psNLpphLcr9Bqm0ovThQRzcS
+/rhYT/bljHqcItFd+TbcNbKrwo0w0MaY7H1OV2ZzGs1e5rt0ovSAdgW4VSmPqIQzEhSs+n0SNYS
Fz//lkWW01cDoptwSH1PmeGtI4vjxqloaFPAmaqyggWWapODQcHA6EdXhirVkTwo7bfkZ6KJkGp7
dfK5pysSHhXhpdq75EBKFRzT00AzNiD/O7ji4DxBIHluHnf6v0csVEf4CUCZQ5dgWkQl9+SVktfM
1shkzSxz1uRnvCrVNUOM/xR/rYruV9oqy/hyHPiVDFWUQP4+ukwIcGgThVsT8fwAtHln2a7FKFqb
sbWysaRYTe7TA68o4Tw1F1ZoPSIVhrjhM3TfEa/J9IvywiDsvXTZ7w+8wQ5nOA9BEvu+U06y7cay
miv3OBGDugE/C9lC3vNi+dSgnJg5OArTypgd+vlHkaTB1DXueUwDT19fPrQeLncFvzw3THiNQ1FT
t8XIIGTBXE9p5zPnYSfG5wPQfSMaUdS08oeUHeLge3aCuateTBr1Ks0Va8fq/qa1jmHqWCtbFQYV
BBVFfavJGzuoqBD8Dml/77HmH7o/IqDXB/qkilEf4iv2FMqxmCrBMTagqQdhCFG9Npf1Ud00QXvK
DPFqUIDuaQ3nt1AcI0UhBbZOHPcJ+HY4MGFFfiVncPDDvOA0GV1N8hZqrV7+aYuVAGCTO+DLjEZ0
4JWCAXgbjveCt5cEUaZZTm1t98VVcv6cAvPXq9WKaZlHCqbEIG4ocLb0bFDx4nTM8Let7/Rn/CIM
fo6Vf9SWBjJW3q1WqgReHbcQ/wMIIPzwCqBc1W59wBDZiDRB0jhZe9z+i9H1I8wA3BR6SDE15D7o
XF9F/1LoDN+rrErQGquqBQ96lkF6sAcUR9BrY3ayoXYvIjCYxne88Gee81MXJgas6/mZwxcvHy9b
TM7mtbvt1xcrDTKhyQZzFrQC0Igv80NLcOjyA7iUQ1ThC3bQYQQsF585wQ9BYlfhFr6tBsGd4+TO
8v3jwnAMVGww9AcfFum6cH4qATHk486I5zUeBK67tCcP6XZR3nriJMl1xlsijJPkc7FRCtmXdxC8
ze7ZkbOhuHOXwCA07CLRqlk//S/kCzCtC/b6OTifClZwMtK/mRy6gI0CwIEWByfkMgsAt0Bud6Bc
jR6CeF+aZ6cmTepAXMEBPAne+x0dozcKu84zJpoliAhC4EdoprL58UaoWLKWFiQa3aNyHqfL+p8J
lZBnEI7rgaYSWlZLPkUURtEz55/lqR2m4F2Z+KiMDRcejcop0QvFmu7CN0HcXAG73ZYHs8kWIp8W
selINQ9BNnrgDN6cWnRxAkYFrz8JiIGO1LgZzNBSbrxeJ1yXbk19I2yOIUpRyYEKE1pVDvV4u8jJ
pltpJu5LXW9LXdMmDyYJn0f9Qtks7ZNCec5jv88iy5YWl43slwmRGyLrXAPH9uZolEgr1uBSwaLj
YdbSice4UOhvNrPIrc0z9o16jcRJ8rwVYnbgIdkxhn/vImzUQFWAwUJ6qVZkn8DpZxLd9D61sYcN
Cwm4lMo/P4KRtkOfM7cEQ/r7oVEWrLDnqxGTG8hEhiCJtYB/CYk+2S3+lWsEx63HgPvnPGdT4rmW
v8Nm9+TlMlTkT3XRUy6Q+j7/dph1tOYZ87n2FL9cWCGYhaccIa3HoqIRXYBajnQ8N4/nyu0rDtN3
FFR0T+/0B1ttuKmTTIU045ECHg8MQ0EvfRc1WLPGmNfQ1ufdj+Co9hNpLvUWkkO7zvHqchfiDaAG
cmh7TTlY54ccOP1nQl3AfJ7nFixaS96REFnQnZt0v6cwA+bocKgg//vzWNFvWHOkk/CaVolfPmHT
tM1dJ/oS+snyZgk8RSAIhOydcCxP9o+uRWgzpWN2F/oqI1GcRRoOurKuW1AW/GT2EVjHnj3CNtiy
N3MX4u97Cx6uaCHySS8LsOsVZyS4nirhvU3Rmrv0ob6fO1rkpXGZdj6HGxb1CKVOQYVKoJKHjESe
z3ZqCj/cuppRzHMgZT7WMi1r56bq8NH8nCyPTnSXBdcwxHiuqR3TQU252GaSpceuO4sZIu0VNcya
9+kdXuJ+DGIP2PnwaH1nxCy6Se4AzowtCc06Td9uIyzho9FDtwHghRiyxt9vBBoa5HHmM8rgkCBA
TrIadwE6wU/CDtP7hY+JGUMHkT+Ug02L289koB5XeD8Q8mxu4iAxgChUsIZrPzi0WtkZEBjPDW9I
t9SsmONY13+2dJvTVPIp57qKP7vXqgn9YK6ouNTj4Zake491DhTfDJwhCtWqKrT5K3qOiXeKYS1l
kA8sIJV4yAnauffOQV+U8P7pMNuxc6IFr4J2ihyAcOI6iGTU5F6goW+yWDE1hQKrEQBEOLKbaFtO
NLXp6FUJHZjW15Vl+JKLsR30+tUVSDsjqn8id+VgOquZihwRnfyAbmNWPJDHUO3iWgHUbnZZh+Bm
MSZQ1ZGJR7iapXMUViFVpk/za/wd4LttWFGpnPdaOA2jDFGzII8BaAOOdYUAy54yZU6lcB81BGjk
nx1pzcnmHM849IYv7DRIFfBzMBCmrqyItAKho6/codkXFZkOUVEcZTBIWH341jlvMibT7cSAHRfr
d5b6V/1dl6rX3jyiOjV9WcGCl6Ha6gA1dtxj9MIyuAjF4tWu4sXrwUc0oF+RH5I=
`protect end_protected
