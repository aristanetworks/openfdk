--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
IHgNB45RC4IPcgCBsP7wnR9h8I5kZ7AnSHxI9Sed5mCf9GFgtY5/SqJOaofh/Djz+MZNna0FPJCL
5kiBUSvkUJu7Z/lwvr2XcDCsyQY5Ssi0ql47zTTmv2De8291gp+strANSLeZK4glNyQOdilsBF3G
XnNPaLrNaVREvtzrMhcQ4zOoxstAoU7otuVldYxPjm7Xb7LKBZAZ9L7THplhApPWEyowp3+zinSa
We+8tNv1cA9G4iwwbRYfvvwHEq7GBDWLmaY9yUhe10kfBXzZxdsLc7/o3ZsHgOlEM+O5obwz/RA9
KdvFFfcOUi+h2LHdnjDAAU6pS/ZP6XheO1yaJw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="itn84wUh+5tlDzadIkkyATKJVPRMcEqLedbLr3z1kDc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
EWOcK6+eFNMen1JRZortqlQSF3Gmx98YS4skhEnsp0Axw4d3gMAJfI4JAXsNcTB9tUMXZM9tnlCR
H90Q0SztcbKrHLWb57jmCR9QW6I1Qj5pM0vIVQ3d3Osm5MF5FckQY7e/irSyVDMKJZ5CMvpOrlRE
ZKpEU8F4J3/wD6YYzyfsSkN1veFwepXZIwZdvwMpDwuhfxo1X+++RyMpvSOU84PItEdUDTfB6noE
qdjQ1oIo//g4EwhboU1bA9NpuFkY7NAuRqOaDyoGCi4kAuVrQlgoymqBrD9JRcW1WapO/+460Uc4
vM8+6BIAHepdeJwrsFEjVtPdo2gQNJnXGF5urw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="deFhqHhWoygMouJTDeG+/Ncn1TAnskd35/bvSw4SSwg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2896)
`protect data_block
AzrFy+dhdVKyH1iMHg9ofCEpPuHizdPZJ59dl/gi9dOPu7Gcg6FBSE9w2ZgZj9zZyzKgDde5OdJZ
jli0spNSKYGA91D6Hh/hX1MT1Ulq3IiiIfxLb8PMESo6qTpVoUmUZiX2euPcETRZ6fUKGAvbTnmj
SJq3iou79bdnJH4zSzrF5AQjzIv0Q/tXkeksZQTX88hra//P4wMLulMa827hEIIG9iYH47bBOzVf
AmiFY57B5s72VAdhUXPA+Hgmq/nFMgWuWcvxruhVIocs+JlJ4A6DSHK5qIPnM3pZvD5qWu3KJsEs
3UDWj3WjAcFBZK4L1oNtO4A9mDHnfqxoj/HOpY6Bja89RxmLPGc1CncAxbghDZLIE30ywrirS1UE
bDMi6FY+Ir//a4Cp/8DQcJRuY5lr2Sf5La38weB3lWYwH+Bbyot/nzKLXOCJB56QzV2JoDod9GpM
ZS9COVzMjMY6sP6toEyYlx5Dy2/C7CJNnW5tYHIrVGr36N0F4CoancB5HB9BVaN8ZrWrlZbrcK83
VB4fRZops8c75ST6loww0xdePzxjOxqu9iJ3el/602/vQamd9eJoOUbSL9OBgfaLn9/Nzs5yEAwG
9J1q04IIEU/ZZnOGx38jRx/LM3OKKbK0uhlmGw7Qp9orZ6eH7ytsgMJl2tpqUUtJt5JOUz8oJk8g
DLO092BX3Y0Wu3Lywh6XyvITQFFeNiXVuMd5zSwhIgIB7FWCfDfnwupslU8PV9G2l2sS6VWGxlse
qo8qnhpMg/nBjzwd9NQDXT2M6ICAf/YZnnUjN6UsC+B7ggGqBebtvJ2QclQz8PfVYayaV06Jyvod
EVdQ8eGARKIVY4qdab+fNBVPWQGuFWKJqSL5JW/rLoxaIg/82Q1Kip2JmAoF8pQoUiyCc9oBv02R
aVA+JLr7zyvJkUf0SOiMLYDICdblpR03pbos9GuCsGf/h2SirSh0pr4KU75qqT9dMBarIWNlyVYg
E0Dix1SK1pOCndDx0r12e1zLrvDTk5TLSmJil/tOfiPD14m11wqFbByLGQovR2MIn8xPTWVvn0sC
lrWEFUo78wDA2HoFbRUnsGeMQZVoWkiOLKeZyAyKKd/dyAutZkYJPtAgJfreeXnxt4JE/TwR7h2Q
mQdfzeQNx2w617hMvZZMT1irNWDbaDL1lwGQudSHCrAKHfocsLLTcDVBb7ypyQ7BAfjbi/BDzJKG
t015xviprzjhfSGTSx+FKYfDYHtGxxIS2LD6yAcU2uHnROWitDFrZqZHmSpUUd8spndgPQHuq3JF
x/a04QJvYKPWoGZgvt8DjBnIYeoJC+qQrwjncBjF5lI77pduIzkMUm2uO5pHz+HZeAT0waZPUUuh
v4ALlFlWdSjwUJ5CozAGtLJU8i7371ALbYcz4NH6kMWuLBrFYdg5Ln7xNrJ8GG5psZQczZ8EDbke
L09jvQIOoIkh+nsnNtX21F7HdePtpQ5iuErMHCY69w1GyBLmRA54Ew8KmNIMVxhsOMiPHR0koG9R
3E2tISo/1KV6YLJarcVZWl7l0aVc2rwgLq6/twUH++VgHPzTk2wENBQFx1Jfoy97mhYcyGcVmh4Q
Q9WOxfoo+gtLIdn6SHf6K28sU0hpyS8xVKsbGQzO2RJb/SoJgSTOlUT1SJhi8Cp4ztwiK8o0Tv+2
WZkrjtr29DXHcmgybbRN+AT6M4z3oktYbPvbi9sstiJ0g3aoByRuk0E24yYxCYRIVVHnne/B74Wk
OHk43pnU5xQ2jmQEWAYCrMz0ml8Aea7AHCCFw1DBfxEnzqLbPOv2WDURetUsmQEvITAF0rgUEtJM
zO82uRKJh58gqyprUML0J3Byc+wGdn9u8WAo46VnmoazpyD5xNMRNEdSOnJjAx2e/Sg/OLHwqlfv
I3wHBpmfbflMHTkm5GQr8pQRGlXIXEzGrFqyeyn+qc8ICMsdEtus1N35TpegZB4wHwo7HsyiTt8d
fryQsewuu6YoJAPd8rjzZVCt6j4HkmnPvVJWzNLrCsDzx8ioAmwyFmU5AYnJ59dnwl1lGxZw3bkD
FLGMGDE3eem7zn/RA9ZA49d6FXdFQ71RTMDFE2jLmUxjKppPpDzr0F1VJ4hYaDJ44T0tJWTtuKnM
a45yAY47UZWyV9tRYBP0iydDsj7Vfchd9Ay43EllyiiNEDs1at3nOe5YuoPmSlzF31gtLg+fUEEp
SuszrZ5Jh5El+SV66pw1KS9CN9fPfmBilPbuiEIL25BOYfQpu/MoF7po3xqPQKxfBJqIrJL0Kw+z
AggNtazJd+ADykCCxISlcpJAue5Cfs5k4aQWcXA3HQ7ogtCkgiTfX2Sh6J4WqWaK7EwyX11Rf6S8
U/rq1aNjDVNeSPxD7xmLczv2z5bDy2mvsBTXjSPRQ8vkcOgwkxBHkD/h4L5PbtwufpqmXGxIIqe7
cVbVPXMgzsPAiuCW2VikDtaRKkYJjmGqawzbbLLmv6ypezVxvsbduDfD9Qo/Lccrv/ybBieUV0mP
u8jv+WP9iorvEmppuOuwdhGFH7A4lQ1k+Tf/+dtK58QWms+r5/autSO/gyb7p7rvmmiQNY4dYXal
J7S9YWz4Ay0JBQ/LvwzoYfPqzawwzXBz2WG8ss+84fsDEn13javsAS3/2bnp2dwFlNUkcir9IuFt
b3WFQLttiHOjdX5VGykoVKIIeXNPo7AncUGjnigspODtat7ZRSslRgTyFxrq5AwoGl4G/Tb+NmxT
wiMCG86Y3aEMp552wCeli5IbPb3E990SapxhANWWS/MxnCaEYKIeOYETSfZyc0NQ/OL3rL+w+79U
XW1zLuokRA8aHMkVtpTRxJPOyy0pJBtcM27dYKiUV42s5E3WMvWRMOQNXAc/O15gMqPNri0rdSN0
6X2JzkX8OtO/ugZVd7WhTpMoy5HqmXe4kKcyfbCS33cuzcnQgkmSy0IgvHhGdvd0kCxKz/R+tswj
dOPpj1CKByFL6PvPJw6djupIQQOfTd8+xj+ZO/LD7yybXbF2Sg9+oS4ItLUEfCyktGa585QiyCWL
tUUmA0FHbpGbQLFnx0E5NbP79k7FFITUlXX/jacPORgBaHA6M/wAqGIaiXgzQrzful9AxJWvVJVg
/FZfaFSsrd41JOwQtxKpUlKnutbew6x40+l5SpF4AKqurfJl1Yy+FsNZYxlLB9zvC2b6Nl2+HsbM
AFtnWYOGkxqSI1PHB9n9iN3VI1z9kbVUWm0Y0CKrfCoLxHKT97LZKD/Ksw/uAq/JA2Zr5Enka1aD
e3AKpVeXMA7A7HzC3gd2ywIbHJSCHELYnHyRuXNGOOkNBwTFZihHoj9VykCDDmyR+nImdf6PiCjw
Flmt99/JH/UXYggngyAZGJxaSu27IWRGCYeEzAZCEe86+vlUGI14+OVJ27mIOOHfEd7etjlsqmnX
T+3C90mbbLIb3kK/0wCxtWG/InKIAFsu8DDj3t62j/WTkbJThR1ukzmOAVREMYNx1o3dKYEuSMpr
3EZHH9AFgBFaCkE6rJqvHzO5x2MNIjZeItrTTdUGQppLIvZ4lCix6LJINyqwWq7/NXtJbJXGNca5
3v5htRnQylu88JSLCLKrvz7dqA4f0rm6TzS7QxUF+p7ZqrUw7FRumEtmM8LkWoDt/k8YjG8iWOdy
91zfQkzHKI5g2vMC66qKOzsmblAlI92cUcGLz4bcLDRJiCPYdquR8HR7RbNgmfaPCfX+Q+VPulj6
fFJ2hPb8pWKBxfObWuQcl3BLg3ZUTnwBCcHZTdTKiVNaA7Oc0j8mvdgchXzhE/JLVSk2CB21JwIw
apuMR/LyYoRctTtoPYipxkPdjM8hfeO6GcfIVHhu2eiIyneMeaitzBTJts87OQ==
`protect end_protected
