--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
n2UibME/DryCt/1WOTkQoEQAawRlx/IXLKqrRQ95Sg7FpNsmQVCdGUKtkmxmJ6FA9OlBdx3tUR94
0F1lodqu5R5fL+z0ER3N6qLBdW3avScYNl81z3MZ1HJ0qQwaRGT1mhfBzSo+7kB0Rgc6EA4sjjvS
dXT5LODc5EOuWu2FNL9KH5AF0GK7VitI7qiStE/kbIowl2T/tnnoEZAPiKO1O+KznfTBw5/g/wpY
EPVmOu9buyPQhmF/5eHdi545w0hz+gG9SP1zMkv7Fn7zVfwIecsZEewuYd9KXUHSUuX5MfG2EhwB
7xSKJ5lY9f6htJDdRR/H9kZ/4SWn0DMZX8VOZg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="UDd6BdZCgIzgrLdGOq4t7M2E01Bjwc7LvUqon27b7qg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
o1I52vKca0zflOstXxckFkl4yS+4wpw/yVHo4xzbJSRmasTcJPVVdPSjmn5DzmQCZmCJQSm6QQKk
rfVPQB5nx4Ixmn+GcoqN+Yk4e9AVYcmrKd048l2/wBFMpS8vaE9QgTW3XhIiax9ZJ9NRglI48keT
hRHOcJvf2r+cVP0bR2cTJK/4UZoVUQMURl4XcQYQqRGlEU0oEQfdI31AYSiCP9UbV6aKyz7RYwER
MsobdzTUthte+t/SYmAn6ZK7xL12IzYtPSVUB3WgiYAy7Vmd6IdZBXShzfmba08HgnZ7T+6AGSIb
uZhqJ/WusgW/vLsfpuiRjplDzI18kNQIXdX+Nw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="em5ksAg18IxNmcTtN82uxpUEEnSFPk0ZhjWX/kGqsAI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34672)
`protect data_block
Kn7XjzPjQ5X04Z1NOM0gN7IFeDRR85rZ8vhjJk4a78a214x2mBo1cj1fAvmMW17VgvfQGmFIge6W
Eq2rjbgfPsykdcOo1MuZT/9JWrUWGeZ8zB5fJdackCJYgVsnj604ecj3OMCfCNDvqOJKwWgKmYsu
ZHxDFxrGP7HHvrbUJqeYr2aGx3rsfjrcFT/M7jhDya1XTLn4zZVdF+2VTMJ0sOh05piAtVtYOJp5
JqoD7C2pzES/Q6Jkj8Zox6/Ciqs7BJy/BlVgdEgyobExOvKabCJBntaDGT2x6TVRWu6LSoCabwIT
YJrN4WrmjK7p6ru9YNvZx+BP7UGeL5G60/jboct0aVFCXf9mToIVvPFuk1iVtMG2AE8k+h1TX6b4
bsbnHGQPtVd1A1kG57Hfr5MgINK7NcTCxOH8HeN0LrpYSHIg0b/oFXmNYK63DaqSck971XCAceOJ
LOfEbvNRYnPnwiLyZXkPYgoG553gsYaz+2DBiWGho/HPbtX6HLCg01FH8l23wZhKkkAF4RXpmLnu
lD05sXpoEsMnOtRymwg/EwiST24090sx9go8yyWMAckoPk2D7tmKd4EXEAy7N9W6GeRZgKbr5K0w
d7SlRZ9OO83Z3UjgfNEsqkD6XihoaNqvwaSbW1VdWw6iqZCoV1vK6OcltwGLVjh6EHuPpEadS+e9
TU1sloPasKX06XbsL0AzpPnYWhlV6EHOSoT9QNHJuhTBM8KaWp6IMSH/6kwNNnNnhVuE9wO0Ejkh
UhILm4VobKJwjb0f7C1GFkEAll6H0A9Z7IrbZ/1lAD+OCBrvScNiciIUqjir+ZhiPy/m3pTvpMIP
JRwpAiPKlfIiH4n/Ory0pCWwrXGNyQQ3txMjLasScA/64xNacOsLwZS24RT3Z/kvXuesjej+5KRH
ppmdbyKBDgKC/8XuHDX7IgjgQeE6uQQvCdEDLTIuNA0oIvfMCausnFWU0TskSPQNbk5amc7e+Bi7
gf7WUflGexfBwMw0OTZGJmvL3tCUVYO3UTfQN9hEcd3UTxrFFO/cDHi8/Es4ddjMB0rKuswVC3xZ
5Uwkxo8PWqqzXQGJ6+5hS01UQGGqfq68tNUZyz2ynhPXG7BzvDR3f7CaTQD/kDXIp0xWuJEMA5ZW
caEobWEUjIqt+Rst5sAbXyecZQv98ARzVzE7rM6IvL3e4Mopu7XORh6HGsuARAVh0kVnjzHtTtW4
42dpjAX/sRvlE6dqjumPSgs6nXM9xadCs/h9iGO7wc8mLDB0XXaFPNas7CHzrN6AUPejMYeL8rft
mAFhR2kExsyQcdGkDA5NqOcN8NnVM8feym8F5vuaaCSFbzJ14fDEv+00zv8v399UeulknCEhBsB2
0fEEQStNpGMx90YvC2BHp4qZhcA74KLamGe3plDT6HyDsDpBN4DJ8Ct/AB6afmfhrHArcRxnLDch
tYT9WsxpiZxEd5AmFHYzhJvhfFQdGbca8Ld0Hiwq01y655alht8zCkqWKXyVxPwS4putLqLGtDRd
LTnR/K9by61Pd6OBNhdFHYPIsFQ/tJoP1DTllhIeewB2ncUD4NlS3JIrdjC9vOWQae0T9odQCpRv
uN3Q0mr/kQNIstc9XSAyxaqes17GQblgkfR/4m6i3HRo9aSmeqSHk9QJZU/lWIiVeCSO1c5BuGPc
CizCXz1snEMEAycqQuB0Qj2kbtRRkdJFA66/6L1S8S0brgt2eY8y+lHG0Dz3m1qCDZ5BZ3KuRyzS
duIwC+X73jusB5BPFYnKiMcoRiswR2i4o8wKIy7POQJgh7p8X8JEDIhnGb5j2xd8sf/v7c/0BEMk
yxp8oGurEwZqsXotTtbZ+qNRkB7IbGiA4M6aeT8X2ypd1zV6vgYOV43+lGmDmi0rZuN2duRdN5U2
/SBGdDihF8hFW10vcftmljgWOb8TTbL2yEG/w2pgC/pdrbVNvls1Cws9KbBcaYk7zT7ZhWPIAABI
HYgZP3TWzC4ckrm8SRVraHH6RqssNhnEXN1tekN70EvcP33oByNK5vbWqZWPzq4ays6+qb+pWStX
mD8QU2V2L5Ug7+Y2PARcWZE3nZq5cS9uLtebbhH6X51KgzkQumrNj586bqqcKyhhfLp54ujqoV5m
xru7HxV6+Mhe52uJ8FxLiKvTn+H799JWaNrBjSAKjOpeChex3zGE1mqirmjtI3bw2AZ4l0GpzpCm
tB7UEpmYhnGMutWORj01RWw7H6IU+tPGSn/RL+HIhjON2K9Pn+f/SxVtlX0nkEor3fHZKRgfVVad
3Fz4cPGCdEJslMdzZvFmYZoEnQt13jT1FTEXg9YQm+ZtbF4o06zK5vuQtDcmCKc1FI42UrgwzR+c
Bt8NdiEqAvoU/DG/NQiFXlLMzhiroh8If7v6W9eCeoEnto9TYQ5rW1h/Bwen6bcgiPZPNtHGwykC
7kPWpsKszw0F21DKdVgkDLv0OWqMJbkGP6dPQUlHpNUgx39ptidE58eUziKJnjonSU0vBEtwClih
0UHOKxABShJpMmYcFZDJYDCyA2NFEJ0Fz4xzy5qRNC4+W7jq2yMuZv/5zPogrxw84aFdaWXiu7ND
ZD1BQwX32qmvuZuHGxk/geK/Wh8JfVDKoA23zRmUOqdZFhnYN0WApHOfaanshd41ZcJqeh1JEt/7
HvDtzQnyzJw4yEBcQYvHjmHbGLMlG9xnnIUcsz4SDSGv86dWp1cPRiNL8nM7j/zk61zMUDj4jL//
Wf7OIDA/Mj8U85X9oWMhC+dJGqrWh1w8nmcee/dkDHfMejO067NAExqW9xkGr+565VgOier4kTVe
BeboEoocg/5cCeUuos0dnpezZG9k392JVARmYAsc4sf8gsNm8cXffAASrWjxO9hMDGLVBiY2OvsC
8bpZg1QXRZrVGfeS/NGRNbj6x4TBygMoOy5SUcitnSUQOBR0vFCy+1asSjZCLtC4NBNdEPPNBdkR
/r9YX+y2dj4CUAKDFeVfI7xDVYvJLisTlSWn1m9i9K+MDrPc8bl+cirLWJfwTtN8xt6Fp+VndYGV
ITvIMFte4pBYu7ETV6PtzUIN8SP1a75Z+Mb3xNrwiHiZOJDQ2w3/PyHK81HReAcnrpd7to/DXIPP
DOZgW+VDdFTF15aRaiSFG7SDX/omm7pWMksvFlpUv7D8wUReh4S5UqdQ7Oi89luisOKFTHkZvNU7
vtXkDfTQr7NdjrcVLMVG1nZgSBv5zEtszbj5kGRvmVmu9vGRGknTRJzk8UEULWiV4J701OJCyqKk
l38Wg4JLKF3pBRK9evMCp+ixZaO7NgRy60C3Cz0+5w+apbFtsN3w25DEPhvm2eOzvFmEnyyTul+5
cM7x4724rGIh52ejq5X9H1Riwou5mvWZ3sKpUaXm67z/if54CoJayyQdXGqtktShJLsGYZlj82bK
6PLJZqqxsahScpIia4KZPVkBhSU4VPO7kD1T2qQlRKmpH2wF5cavXvSCkPRzmMMLx7KH9igKl86F
HBycF0MoJxyuPdvse2eiNjKjChpaA/96r0wVtWt1bAjXp0rEEj7VeUAhghaz7A62GhUevGkTeMnI
T6ZY+Ehg5szlN6tMLweBs8bzvG2mUjVH4jW11w91Rsr+5fpCst57EhTlwRrhgt+EL72fflLtdxrV
l/d9j8qmYr586MAHnvn5Fa3xmJyBrlbXS5pbu766vhwcxGQP1c6AigKx6pSLv269KUo67TINLNzT
R3GLSHSgtIIlSYB3kqgYec3vJeoKsZhxWEfEcnzbwwGUGuqQhR7ZDrOOcwDFyOXHdTtkeu2qgmj3
yayJvHhupb6LKiMlfPh9fGVlkmw3scHFdD+zLDGwXMe/hG2bpg7N7TZJ69gUC+P/pJ2mSEo3uciQ
y505Vv/NEXk5eHVgoEsFqYeabCwPsOzSfVEBOKIVbARLjqs4v22JS6pnWKgneJZ29jY13ehNrrVx
ZxcXRGpyWl7jdYYmYga1Cgo+CmvcedvPSi5Xu2P0tghEcvX2zTcLPpT2mrvlNjql0Gl7F8cvqHwy
8eGS4gWDRGmF5R7CGvLmiPWYCJUyKGQZLYmMmvx+ZJe9Q7YMw70raPC20j2kjppwVNhKfHsfQxNH
VbF7a9xwsNCugLvjgiyGoHN0Zvw/cpoEEMp41sYY2BqKero8C498CB1wPVpx1xc5sI6e0Wi63S1l
RAOZlvmvdv8wH/Sz4i9nWbo9whr1CUHITIpZH+VJOp+f6BHCxbaU0DVqARtgzj3JQq6yLJo322Vr
hIyjCbo4WOq8ITLiKPrSvnxB7qRco1tFJFHIfKfez/xJF5OF5Phv6mnnz/7f+Z5/VZFmGSsw0fCx
+sqWnEQjZw9i3AHq1LSxRVEbkAbPIACjNM3TP6NotEp+OB3a3iLrDCl4WJwdSyg9R45pILt8Z9W2
QdzFr0SoOtbpfpY+extIJXO74Vue9xQq0sK2Jgiy6Y6+Mdp8jjtecJlFMg3HlM5r9jNwuBfw0zPS
1MqZBA8cBwD3OI6GVIXbm5aDFyXtTxOwY95QZx8Xeesad4xaMhOta+KjP4v5qqXoJaK+mUFXknft
ne3eSIGFvG/SbgTp9i/pVT/tx5SSaa+8xbzmFDGGZQRbdXsAkVhJGVuODwURK/T/ywFdEl8IXnQt
FepwbjIZ/AlwURCpvYtugzhyFI16yJRnynn41EFCAzXcOD/57BTMIx7bbWkCOpRbw0HiPbPqghY/
D5HPsOzOyh2AztuieYyfEwxE7wHpwq1ILFJG32abKxcU7e5/zr9GtWJvwyS+irhpmCT2/PLqNGNM
QM5NCDU3lqHNRI/lmkkVJ9+z2dLf6PxkwAY/kt+TJRdb8PjAvz7GmZzWRZK6uDuoJRNV7DJRWDq+
CdEUNrWGrZfescAO/X01jN23KX3Dz6dChOoPgfR09LBHwnzLNaI3Kr8ZeeSZAsIBze3q9GFu+bK6
lz6rBuki665h2h135U/+1pqfOrSWe1OENMOcfZMjlZacsnM1GbO+9Qmif9WHw6sbKfQQmDyGb5Fj
23/m3mm5uEzeG8SGY+D7XI8kHJ4oPBi1g30o/BxYW+3C95HSb8jokPMC3BdNWBHEEH323SWKe5SX
S9L6A9TYqYsmfvZAcficm2Iz7eINKW1v4duf+Yms5E58utqOrRIWE70RQkLL+z5UtGeyXstzIs60
FVflxyc3VJHRlu6QfYN4sMuqVVrCX7eQyhG6V7YFgwOUkJMVTgfrYY1no8KDbEybc7Iqs6gFmEA2
E/ajA7ktMkfRLmBTumSKVh0ixJIM3MUcY/hbYrTbj9OHch+2ZZw5gL83mlT7v09B+Q7OBJ0VdP+b
I0y/eOCnLf3H54mBzdjnWz6TN0xUwLNmTt/O4HemmN8j8NRGKH0K3i3su2XeoofjZNHSajPm5p98
AVqCCqMal8lMXhMPAKx3j4CZgNS2TqTDLThC2oAq4cKDZF1a9pU3BaEZ4A6QKkR9F/mig/JLU9l3
WNZKV+PMglZ7/KYgL51lWBWblRsBVXHY419dtRFIK5mdLCcefgfVpUfyllUFV6zUd/+o+1pXFupz
bi4XlrBXGTBwYSTD4OkVZSn3969EV96JPnbUgA4iNxgVJAy1RiL8LrlIWlc8fJio9F+gdRRTzuLH
1ll3mLKi5jTFXOmVO95gI4BSQDd7x0wLc1xEB2ZxzyEXG7gWa9yyYDP+17tQ6HL6xxHqHPP02MMg
0c1/zFaGUNUJ3DsWIvhOSKExoblMafLxLxyz4kZrYwBBMS1qL77CDQROjVQS3c8Wzz7EVNBQp3kR
6KRMADrLTZf5rWG9i8S2vVtSgP69579KJOcAshljUrWPnhZxUU6lFoPnTPewjfKP8MyOO79R5wh0
vGzY1hIwz8zlJmeoJH6D+eR9yHE5PDjdaJFEknWEC16aNS3K4hu8e391FVHnJgKblYBaUTcX0jw2
J3XkCIOmWtWQqYznsSJibmwYS2sFQ+W9fxspx+VRGjGupMCWArso3bytLLd/AYkHrzYvDhIOdeuL
NupRZSffFUCGcDN3c8/M3lIUocduFBjkFo0vttnX3ecz+ow5hwE1qwRFy4Umw5Yk2b3qg9IMZXQ2
pUOaxBBsiUkhKH9shbd+P83rHiAc8TUk/f9myxIMKdCgOwkzw+im43fKVdP8XRuHW4TN7lBjea7V
rmwRC4Jn5ydWDhIoOwXyqf8J6EF6DbeKlbg6jokUAWsZClW1p9nZxhnhZuWBp873/9Qrkbmdsh23
GVRfzOlVzBzs629s1BGTSmoNZZtEyxjbMVpy7VSM2V9/h+48x5DeMRIeSMmswGrC+i3ILYkP5nw6
sRD8ZqiKkgHHxCzs8lM2IwKEJHDmhb7SB7ctA9V7KyiaKMlYJ9cEaQ4cjRIqcTC9Hq/WnjlgSw21
blEUJtPN/fi200XFEBxT56PgzGG2+GedXTmDwAwwS7XUzgyF4Ih2HNm+uJFN0KkahNzZRkQgwIeE
TcW4NBlXnRvACbS48N5cU/ilV0kkO7qst3EaXSNpTGiZWgWTJjydYZZLNH0MXcogCFjYoMXyiZRn
hJRpy7SEyhpReT43My45SwYxENJH33aeA+Ank3Jg+Y90jZTad6zMIBTLT07KWiaOsiHxLPVPl8qb
8S3Oy7U6JzlJ6gxsEC5C2qJEb5KBY114IjJdrWt2rM6mucGAAuFXo6TRo20r2FtTnlynLHnoQ4Sj
L/dENwOX9YzlGeVZ9BQYebG2WFq+7chZWOtGOSmllGjV1AlIZvhiG22NVUqHxHL5rgyHHiLCaCC5
S0aH1FWUUyoq+t24su+wYlWnbJk7meYIeMITEurmpAPh1WcBAv2mVTXaN7GYr47uUY+cjpNhZb5P
ZoH24sGDWwBUXqCHxm25LROIBP5QfXTXHCcVgYMsdGc9usfi/zgeYB069+KnxoRfEolbCLySdvXq
jlxNJ/1v3Ldmj/76TCuKpCJmUhr9jFVGuS5jA4R/pILNiflUmrloYwqJQ0KgQl9VaCXwbIOYBB25
9U8D3zFCi0ubBTSNS1OfofETPj5BdIOnorPZMQJsI+d1Uctx60qZp5xEEqjZ/1D04FHnOGjaCDgA
LjEqL71P+hwjfG957h7fLw/Rhwa9oLnLV2D5u2mzW7eAeBW8qMOTs4I9iM/y0EivBQFubrs0pcxd
eno52YBim6UDYEUvU8RtX02SM0hRLdivR40hKHrbkdAVElzUOmjugL7wNIz47OiZ+tSuAcpdvv4+
gXMmBJPy8cqXp/E5PhoYwlu2YX4jXVjGDzLWM+HI5dkM6MUDf2L9rstOgdXEUgDRhfleNcA3rS74
TttTnBd7PlgttWjl6qk9iMDYhulSklN9cL0z/sJ1yJAXo0XqYrKKXvEEXbRCzF+SqQSS/Qxl3/Q/
9fzeFmi6bgo8W7AmrEXsr5tTRc6junCe3ohPchlWDJg/P3upLfdUMwy2VTPjaHy/63D06TitFIir
042nS4P5qCUSYYt+yTyJIWgyn6NjZlElRgxn+7mC578wTdIfPCrS41Emzk4GBdTUUzRPEqFBVulC
7v7I/aF2+BJu5sBlLZizeHJ7mPmK+aE/WtVSWh+/KQiBpYFsw0DtltossLF8BOuU0Nm+Jm+jCIjF
XLr5fFzQZYFjL55Ashn0IeGsZzvpXWvVDu4cghd6v1jFaPA5Eakk25W99HBoelXAyK6d2bG+zy/b
8QJrgT/wpiNYonxsACJ9XDQGU+xbq4hIann5N1og2MmbFPM28XtM7+hEVbUaoPdu/oW918ugifSN
FUWCI/lQF+UQyoE2LG4yjZ6faTPuB89zQqK4+idNHt/FLAEZYjEEz2bOA42glhfvkWojSi/SMjRT
2ZA/U6UcqI32lpMlTgDiwblaQGvy1FzUQZsh52su5amYISrA7b2QAWsBY7NPM3uwvW7FqBPzDYlx
l2GkJjZqB9idq/rlxDr3P8YIAmigY6R1AJ4bh6/s8s88t/S/BLS97TROITHBzhGK3lkj328hcquS
ZyUD8ubew3cSAgrS9dkoZkjShtH53WVW+rE7sE5yyMFs00IFXAv4NvAcskDFNBkjW1c0+mQUuU27
uSlhnHNfaemdizJ7Kse+g3sUaxrgFc7xvzOgyyuuUVrKRKIaF/kET2fODsp+WfAS0ybJ5JC+Vhqf
SZVSUn6tWWmrPoNINCnB72DHqYj8U2tOBriD/IavBmMx4fgxMBdVicNSJg+c2RLyWOxtzxjDSW1w
GrpILrpMM2lfIsU1brWW8NPNa13RIf51si3jRGqTth6vpsr7QxVKilu4yLM0P6qp0gSj2VDHKZE7
1yVW0mvSzuuYvkV4cSBsJ5ZrNL6IVwDrZnEiOWIH9EJUprhg+jwP6jCva22reTbX6LladeyCPnYw
fl15vGxXNA/T072See3cjYWhnIwjQ7L+zYipAn+JkMr+4u+33MiFD3xgR4Yq6il2Ep/iumHqpjJb
hV9/7kr03NY/3FBHT8NTH/SMOYQKqMisk6UKLh26/GE1EzplnocwGv/xZn14AEvU7ZB4baiNWXNm
0pSdoGKTKWs5+uuELbJENtzymHoxy+gnTf/93SNBz5SpLjBGDA/hMTP/1+RUIW7nXR1r7O4DL3nx
FIS5NL0GuWmVGYi0dOSmHvJBVGBUWYYOHQ7wGFS8gT5uUp5kXnYrVd+OZ3FGANrdQN6RxPTuPT7v
QbyVUQUBqT4QhTz7i5CCnNsdi2DISaHJoiruZvKzG8JLnP7iIN/Z9XwKrjgRhrmgT3i26th4XEqj
X1vyUm0D2srLGa206yzUYU9ia0SibzE67Nn+ZPf70Mk+RW3k8kWhfk8EKtl8Y6MBtvc21tqEF7gy
8N03DMRt7bGO84zzOtUv1z05FDNs59MdPjyKm1+3IwVHi3EmctQO69SyKfDOXu5xqpJNyqRFr9ZQ
t3m4vuuxSKz6BHrHcsRhk0JK0j15JVhKtFUk7ldNbF/5gi4ST0qY8P337PWTpdNvTUk9+rUSGQoB
VOvtr6LTQrupxQ0leNTB5gByMHzuWNpzwfuJYearIz9t56cBETWM6V7oe/2LElAJa0C8s7vjr9fl
XwRsDYLEU4shYwhsPWguA4tw6HBMQghJfZNt3irLhahHrw3FRAK8Xg68J2829s51ykLLDi9+SoqQ
eS1lSGmS9dDByGKkb1DsTzQEcyOqwv5GRvXj3WOPGAS1PjP0JRUH793BL3AAo9Tw4OSGdxockQ0W
TmC9/EvNSPHF4/HU82zlvkfHGd+R16DRWPIF3z07fKMw8LsSV1F6VgDQY6XJDs8AIggY4aUPUnE1
CjKW+Icpyv9+G7776WnZzG6MJe3MpSXwYaHH12qiWfqyFu0Q6ok6wm00AYtOBc06T25FSt0CjNlC
4WLDJT446rErX+f6gsnUawKGpGEu5h1KizmbrK2RTcsaILwhE8D/oRLjWxBq3DdXoB5L0Phsqx+6
IQeQ452ZTZgdSUwbAYtjnZAF3M31xDLT5UXxZeOWqGUgqawq0vJ8c/FnPm4w423L2jU0rxx6nP4V
6v7GtwBXnECyKJPR9hMZ42snCB/HTW/CB64NVnpEpwd5p3QBJ5ouXeqWS6T9aGNA/Pr4TMQnXorY
7RvNwInaRECvlM7YU4gyYNkYb75JvGseBgEhL+PgRUc/GIiOX3mj3BEjKw4sCW3aLJaaTlYpPYpX
RctKjSlqrvUGGx1JwHcyiwjgYcF1cExmkdc4A0h1IithdXXVoJ4jNdX2x191na3S12M5h/LUQjAo
kBkE9CbS/pdx6eqoxfRkyy2Uc52XGa1+gaZwAERwkZ3zuemHT0BFdztzDM/0iT32H0NmxdKFAiJq
UE2f7azSbtlqo5RKDrj6FATZOcAQEj1H6dgOjE0OYCTMVdT+eviAO5/d7LdFfsn9XWaYUPS3k5/V
FKG+V9NHvO8JlzwzuH28HQ9xzUHStUElT1F+Hra+BT5zO2UECjy1rg22CF/5o8+5PAiO0x+Thjr8
LBX6k+LrfBtFA92ixwjBWzMz7q3enx9z5QrzIpZV95zdvohsnvDVE0huy9J/+BFT3VytpB/m3sxV
8U8ObBYcyGbhyXoTJ+5b0gs9YYtUR9dUSOLyR4D+E6WR9sHP7CoGSzugy22VGZxG6+N2sXUH69W7
OByry32GYjtT+yJ7+pVKzm6iMe00o43TnYNmbfmcVTDmrMoRDNQZfowLCv3Byz1cWG/HkzsIWZDe
7OoGC8jn4RiUivXehPvQQHUsPnGp1tPiHGt6VqQ3HrVvxOV+2eb6XMgeNrJN6dtQM0nxEImFF4rr
q65JEl4g2I4DFeJproO2NhNEAUtbV4Gy6zLsi8NjKf1Teuhhzt4MAJm/T4oKrMMs2eI8D3wcuewQ
mjlUqJl3F6k8hx+THwXiNM53cWzkSBZaS9JnbMjVk2Kav/V+Dp77SzYxeR/JQKVZMf3j6vMW6qm6
J9pp7lwwZUQ6XvpeYGyC502rwSR1hoSTBXZHoLbmEBB1QepecE05JAVIeBacD2Pat2NIWIHcOiR3
uvBIiyRQ6Wn5WuvcTsqKZ/Uc/J7ZgOyEDP348j1kGAWok7yB65MKJwrIclk0M68XwSUaRYb79dXc
YKLRnWGxUHWBWVf0zO09nB1Qu2F8kPDV+cr6+dGsejnr8u34oOfF9irV0k9G9uT+80dap7C40JUc
EoTur/LTuD4aKRXUAfqraen66ssr1fOvlxP5cbFYEYcTQgqWLGPfSqnvBDUxBlgSR9ujgn36EisD
fnu1aAIAmGP2PYrOV1/wEIi0eoV7mzD3nA2yecS3RHAHkOH9ENE9zgGmtBPzS88hT3ptFL8IDSeU
2KHB7LgQ2ssJLbrszbm57ANJZPZIncR0nbkCX7cK8rnu/lajv2Cnq4vSoc4NRqothBpE7FRixsUG
20mpE+kYWn5CFe9lki/wTCsCD52fasm1QR5P8hp4WRfybiMB63j5YkdpJmZ32z/bZKERB9WeL7jU
X2NIdR1/BEj/NhcWW2G1u1mAI9LWYsPAYh95GQTQG31F/nwp8XSiQRIce8MnXsjqPgczN2PpyBla
vcsdp7GbJSgLqtN7Dvz2kYV2pPKUHWjFdINW5odpW7taFfc34sFTFLatY4/Ahk+armTkKFTkmVGU
F7jfGCS0yx3bVjHtvCVrAbN8RDx1UW5zcsXWIvOkp7Bv5Vf9cNeDA3ILRyknu5uHocjDQ5tTMqLL
lMNHpdtxp4jYtmtCxKwnpUMsN1Fpo1HtS1jZyjl8MLFY4qluzQ7Y3V2UYymqTmrmBc23inu+pQiU
tgVUKm4DMPWYZZvd93HF+YUPookAvd213RwiUaPgy/5P/mk0qIi6g1AJoKs2Gwreww1yI+ylqJJg
zdFfrW10d1kdrozlrkEN5cijwzbgwb0LFVeZTiSOZxGeEAMH57MviD2Yp/CS/SkBI7T6WsQ4Ai1w
J0zsh6MSq+r+CbFN6Jzpwu8srMyJjZ6bz6srobY/5/EJQEkk5t4DLu2e5jVF9hKY1W6dK8HPRwRY
gPaDKQyWJlPsz/EBa2YWXun6EM6AihfSrUpUGa0fJiak3ZNbzxvYSjlnQYQZFNJzq9IUAD1QwZFw
V6S2qp7dOd1zwaUnvf78JqAveK0Vamm1p7iCc92+AUYb2Ll7EKWpTz01zIye7vPdTur5d/JwITqf
SQUZulz0vuOI1NGQdJpzVIt+a7dYqdqgN48AYrNesS7CbUENseshrQsmBLLU3I/QV8j9Z3HnGJUp
anPf7N0YP1y7twGvuemVnyoxaGAcub1iNZfOWP85/4UxdM0DREXUiFGzCXrO1LTGycL2IDMGCMmj
/fBLhy2DmAIsdJ5jirUW0zpzzKgmZ/Sh21iocGuAuWGLe/RyM398wieuq64uEpYrN3QbKFwHsq13
q+74xpWjq2mBM4b1HfwjO0ZVKfvW8pLbn70wOXnwKGcq9x2ilEmZ1rHEJcJJTWpxTUpV4nYOQpFN
z1ty0yDUZUAU+C7s2NB6ZPME/nPQ6HvOhVtRxSvr1VXanPuNwQECvwEPubOoVG02RHr0If7zRuJz
z/1cVVR+4iEeLqBDhnIhm67LgknOqtpeJID2WuvCjv/UgwSPPUDdoUQcA3asS+3LZ58YR761E6WK
hjkD2BPVXLLa6+P8kNTQLZx1kJ1CwUj+RiwzXiVWViqqPvDjjEOo6h40+GTgv1kPp/Lw9ykzxBVT
/xal4kPH1sE+Am2fqgMVdmGucMS1VzECT/UnxS49C2Cs2Gbu5qGFqzA1Zqzz9aggR+DYOt07poJG
A+LfEecJ7xTXAt1Vll9C7lAwFDaLrn9S+klYmBZcOaIsblOGKHMB6y6Mu4NOfe2m4stBrBCr/s7k
I7YSrP4Jt9iDWvKzM+dWqFzSYxb2vkvi1u8imVfzJw9fif6GAQZEoQsewFOxvO1+XhS3Ylc3+VW+
b95fpO6BOH3SfMeq3eMVIaO/znOu9neXonR/wrItfyqpfXFZSX9zaFLmzpv8blVmMelV5slW8ENa
TXqJR/h8Q6+SE1R+46Lzss4Jkzcpnxf8/IY4y4zRHb/m3tiSwZc8ZGpLK1brOSHWL+RAWIxhM2w3
6ODdl99muPf5lJnlFN6epoSQOepRdf/qxvY5Za9youTTcw+L95YxjyNEbPxoDXjsuSF829nDI3jT
q+2AoO6ktzNXAUpnB7YSWoPrJRPjuU78zXGV82ZvmFSFdIE1eaB4tKnPWUPZMpcBh3aLeENvMZN4
zRlzRAVtS4bV6adSghv1hWY+M6KQZebS68T0VScpgXUQ0i8QEcyDhngJ5PELQPtaGVjundfdqxNN
IxDlALpMHzsh1sSclcVbeQzswqkpCgQ6aAmE1DUirkDBUAjJKbPIoULpxXKJ/agkXxwb6lO29GP3
NqwojWh0jD1GcAqLVbhkXnjHbR/yI3PmYbqtiftHVY2OdFisl1OaYbxWX5HBunLLdcS7KdqTtNUW
XfpF/Gey8hsnsVtVBRznxJbs6gwIMZ2P3RCDVeSlhapuGEt8/VtbgtbZQWinlbyhKxlDAOwqIsCB
f2ijH7VAtzGprzp/6SXyUkRImQ8nFzGWgVmqk9QyNqJBtRQKjn2BFdkmPj/VUUImT7clkXrz1HNF
ITpP78aRW37SSWP8v+clca3RcqHOHzeVOjs/dT5mb73UXGlN7LJQman5CGzsWmxZliu+oYrv/9ZK
TlB91vbwMawqgsLHWkzs7Q+K7SZfIxkFodEqoA0KueDq1iFX1ahJwPIh5/ikPJPlYE8yTBN5GN5D
m2+q1SCdBd4lJ2hzRASyrfR+mzMoj45FfbiGj3xpS3P8yUIkg9HgUYwEJR1s4Z4oTciMShw61eZV
hnCnl82pXO18ZsZ8Sov2MQ0wcqnHGYwOdlrx8sNJ621jTzgS8UvlC1DaGGCfO4lazpp6QtKU5rAF
y91R6skorp0TR9nkX1xPyCDIcU+MRw8tjNIrR7Jqx6Jwi7d9dSdxhXPBHs/W/6bHrGxvrSNGpr45
51tpr4VBdahFNh6z/KAwPTfA8qUtn16igH7XjuLuAVcKbpPSZmLYfP1T2vAJqWn7ymhfy+YOtaMx
cygwbSJy0EMCxJT1Kzbo9ou7PNd9PiNUWqU++7qVjJ9t6+Uu9z1/Bgk1gm57sqiW32ehZWmFf2zv
NqH4hzBsEaw9jOjIeULZkbhybckVHkVnBnJ9oqgCiauptjlSdMOFlr1RjIpgkLL555T4K06zXfff
54yeGrM8dFdxRWd4z+yYxZFijDy0VyNY7mZOfODzJstx34sG3BrsJEGejj+YgaidvAqOGP9jL75C
LKb7CtRgGMCJLlIy7glmgLt268OpxWdsB2CiB0Ql0lOFViZ3TTL11M/H4hbZQOjxO3g61oIamhb2
awnYy9z64ZUTgnuIic3XIPiIxAMgA5tIfPh1MZNgzV5jaW9ezHdi5emSIb9ny6eZHDlB8QCcgDdY
eB04ahOi/kPhco1l7QZseX7CGp+y+1diwOYoxuENiEynG0yCeESyDQNWxWpCXi7MuI6OAKxMzziK
CtLU/3UMSdCawDjAgW7fC8JfELBI7nMtvOUfg13Uy0CKBDg3cMPIZCrnfJfDNorQ9xk9rXVTcLk/
hfzy461xqhZYRrgW0fbBbyomYiipQ9sM7sXmZoLIeKRsqnHMS/6EAJ/cIa7xB2+7yyQvye/BZUSf
hf4rmyRkiQyK1dcuDb4zErMx7vFSl30+V+6Zdmtod3BP2Ludo9f/Ep20kuRtv4lkdnWXd/xhZYR1
OP+9Aflh5FABpWPVHaf3uViCN8e3sXRiTsIylV8koZ09GEmPTylcKoxtsKmVr09FqYOoZ/YqwTTt
nPmrXHMiKllesrprOaThnwMcZxJnE7U0Wj3DPnESLuibhpE2zSo+kHbMdYW+3lfgD192nytNTjtp
gSLbPqcJvzZFh0acV/RLomrSzpErX76tm6kyKcc+GVTOcIY5DJlM/SLLyP7BCcZgeG07Qq9jUOKg
Yt7VvqQa9f9OG/2u2sL2RjY6OpFzo1oYhok0Hu4JbwClJnQhjWW9IEIV4tV55ZHiOFFlvPfcLfjR
JhvnX9Ycteuc2g2OeOCQClIUdgI4LXVbCYuTtZaOJIxHKygVH/FkdnmSOiWv0GvqKETC2KoEb3pC
v44r7GsJuo0We4Imzu/jozReITixDucJKW7d898dTc4DLDHc6TS1yRhI5dH6xxfx4q/G0I9FWUt+
Cws0fVXM1PI1aloSpwWj8BrfDyMnukcvvuvSoZU4QGtHjImGDhltsWT6A2icUw0kKIR+kkktaHzW
TdXoSF6Ci/XYMjj7o9r57rC92KVIA75yAW7VRHbab1izCuNM9Z0Q/ynK/FsYFmrhEYkrqbUhpUtD
H80NAkkcD6jYZgNtOy49GvbFk9Bjd9KAISXLA0x7Pn2jnwAPWGVJgvsjI1WMBSQli4pGy5qdHimK
BDyuzGWihiIm8tVvbznYBg5BJd6Pcv6MxnTXG0PHYykjaOltqsdR0sLbWeSRTPJrhOCOOeMQKhVS
0NGQUegqkUXHC44XXTQbL+BHppJRsdZsb9VBBVFtE3sz0LaZb07fzCHoJr210VJ38vujdApgATC/
CXeDvHXrny+Bedr8erxcme0DzIqA3ElCl7+pwvQ2B/eWxz0xUGHfo2ayhJgKRJ3qHai8/jH2P8lv
Qqw9zQUGCkVW47BsocLb7CHQzxJDg3ibrVni5XkAdOfciU0GqTL1YZjcJPStVg3GFiCDifZhI1Q4
cZuLb/WWa4Sw+RtAm1egpB+equM5z8N3VR8b6ida6H3yd+ID3t1GLW93ZM1jTeexYL/jx//LeIbJ
BEfoPKtjGhZkWcsbf/H2A+UbyXjpdhAP4W7H2NMPhXFrpDe9aPVZdmCSXnxlf/Czg4XQF2tLFFag
LKr6RsXNrwjr2VFj/0vIzaqFIhivNx+/ZvLUobu8dZOsNS2aLJPU+hg0y+3/zv9Mn7xulyS3WYoi
+2uWBuc/oe5W3p9b99SLUQEs/gsKXvGiB97XlsWVs/u9/wsZAdOYMB+aZZUMg+JD3GnVVM+RGzpy
xcfT9+I9gnpZU6fU2IWqtxBx+WDUwCHvo1IJGkgHJOzC7D3srmw0NpgLCo8iHRHZCLOQRoqYGO2x
HxX9T+whkyLd8lOKN5FeF077DUT7Ycx+xiXpU1+c4I/BDhX7bhODdIdWMBKGQiDsLfEWVPFrdgff
V0BbwU29J71i3IvJIiUsMyxqpeilxu4N2dubro7hArkefbFihe1pd1j6JU/5IH3TbAe6vM0BMPNQ
5q6QSYz78t/WUtbZapOzsG1XAdStOPw4M29ZIkFcl4nQ0kktZcDZRc8crQpx//E+x43w7K1Skos3
oh3a7l2jziQh01mzVh7dfO0sKK71RP/vWZe378depzKxuJ8Db0fbcmO9MGKZ+LoJne1YxG7Jd3cY
vnXf78nm7AeNdDDTK07u+pBELAQTbBlg+PbwjVVIGofhzNE7Tt0Rtl0zDOaSfgAq2x4NqoeuDYeH
/HugFjDpbciyr60WffHA/hE66MzL7y8BpLX935uJ6HhOSP/uAbvUOtu14paD7CIh7Mg4Q4RmHkix
wSA2c+ic3f41qBc8zoXWss0jQbKAKiXJQrFkYANt+CyHlFmh2ko4lOfXPsOINujEvg7sTRYym/Rj
KjYXPWl0vUzSa0dym28YdaUCVj2zMknhpJUTVEjs3ioQFVh7r16PRLaKjgMWNvcPp9e0EYe+BOcJ
T0VvyCYRytWHMQTdfIDGO1KdSDJLN4gSG/RfFFpWjFNDYoHy5gshc0lHicaGwsgqL+1rgcaIwan6
OyXuFPkuroxZhOFXe7H3QWy551OcfgQd7VbZkfisDeEgTkSawELj7/ZWZJ9rWDdP7djTg1VZwKwq
zc/KhUAXSMXlBY6aSzbtqiyJUZc+5sXc8iy/vSOAcFH2hV2URchfm6lpJgYq3Aa7NOJSCgB74Q/c
Lq6pg/Zto4feo3mKaO70G9FBmkhrFMFcb5Of4g0qmM96dQPr6JBxAhSTKVOT6oFNjbTJFeQiV69H
qabOwnl6ryHPaaZYcgX+wo0H2674/DZBuhjipAFx6gHpJhwDlG32LZxwJqeLG7qhELEVSFsEaIkd
DKPW8I9yaLb/ImXdd+Lwu2heUodF7oTCorwAIlkyeVYYSTu0cITAE1SPaNs9s7rhTuVl+EU8Pp01
MLiR8j2Kmq1gTqW4twYVvfKMG3u5qWHPj6F3YRb5D9szVPmlAzPZ4G0+GW5f5GDx/BR+7N6aqFEz
Ji3o5NPIXCDyJCSn9vu3TKwOfJAob/+raVVWKQ30wlTF3X0QbhrHlQgyRrgcZEkC0gTq/QR4sLKC
BnrXxCKlXMIT4SxaJPGY7R7abkk4elWDOadslY1s6VMAGZ5hnjrMLhMEMX+2Y6ulRHZlrssE/E6D
uZEiFwArARbnoodBgwZW03E3P6oZ8ByzDt7SLTgyenVUt6tCvtQk+YIxtsBtXBS+n+kuvxL3dAU3
8eqgCWF2X1f55nFfFNfpDUhH6N6D+A7tUNAApbMDu6/mDKcfojM4f/XeKrx8GywBZXZZLfB6I9KE
mVrZ7u8BFDKROgH7fgcT8hcz0BMkMtHeVqIX/0u23LG1boZ45cV0FwnodTF50QvKo1FWMaWenHjc
RwMJrjszIHkDmIpGVMYUGpufoZ2/iIHAtbRo+rBVOkjD1MR9ZTdN1557L/f/3pRDgIOqHczCSf8k
4f9BJM6E24e9pUEsnL5TRv/P9gG+JVncYuExqGb6G36j/00sGjf7g3wyPy0+1Tpz5AWqMC37V52U
UbDCLkCLouQBP/IHQs0UbIeYF7Je26u2yY/HsQWdx6lLllgh8/H+ZD5c0CsRoBTqbD4TyVZ2YDQz
O7xr3K0wkT2NJ1eOLaheshsQhyhOr3aH1O7MAi0PMpmO57hc1GknUkHKAMPop3e3V9vSFjqrMTOe
3ePSzperHoLhc/Ay8k51KwzJJr+3ovqNpF/9Bb0O+TiDAoFNRWgMcfqb9DpN2YAhOIZ4Nrb4CtbA
xSSZ2Dl1ybHv1dftQudpYEn17qDK7TtJnDqjtw2e+lL93PRKW5eE8dt9om/vIQMDr7mEWWoMFERy
g4ClrDEUv6u3EOyaBFN3qyiizozFlM9Bd//U7HVXHyvGFob8+lufMoEEbVeW/aQJDawGq/LSwowx
sHwH9Q+83La60s9wQN1b0gUgUI1YkXwJe/sX49FaUo9l9P9RfufnDcCZ1QBhLcRP+Y136vk3DzPN
x8Ni+QkXZvA8PPJ8sQr3cn1BXBnGSEJUA4TjS4+VjrPc478RupyKZJxP8H8MBXwt6dMYcsvW6K0g
Ape5hwsPZkxjlsvNbAnOQ7KpAWMK5X35bSy1lVrO9M3Vovx6eme+HFefDPxBa1k6jP7a44VBzEQi
5ihCpRsCU769rrQtG/JMEJewGFGn7IBVMacRvZnv54BJQ2XQaN4GLwDr3iat3zOk1kgOX2HQ21RQ
qxLjruaYZjwsNqqPrzOljPgLnjTg6RphHlgys3NHVHF4JaRnmdiVVPq4Pt9bkf6Y786haQpVbGJX
mgzjc7TO8EC1856q7QwEo80o7clDjJX8BEEnF2ssI26fFwcVWamDXyTpkc4n7WjP1CKt/E4/cLUq
KVLxZPHtj+H9EdgxjcOhGBoA4aUV/YFurMizxe92IVGM+UyQa0u58c1Gb3Iobbpfa8q8YRDgrU8y
WltSXw0e+BoMz5Dh3YzDvFFgYf+om3rGY2/nm/vtiNGOGiGXD573di6sK/EhgbhXz10nlijg5GV0
xyB9WfMdEtvIGdcogtejlIOhZQamSJAOGRLk+fT1J8UIqHN7hLP5efRHoL8+d2p4W1mJBc167mzq
2f4oagVCrmEBV9+8BZ6vR0TVrD8DFZqQgxOrX9cttKaisJZcDE4JG1heg9Gu/mQrtjC/dRDARi/f
CjxzAWJ3FLBMdk0d6JFIIe+hm07p5FE5S1R/LlZ4+cIz7TJtXuOWFdsJet2ZCjc/V2krGQ9vG3+E
oqNYitCuXer8wACC55zJUX5SiaO9SK7cHgbt63tcct5Gd7oJRByxoAKkb52Rj1PU9nz6RBB5TiUQ
8e578YxHHZ++dnekktACmGIrmFQoUuTyVRkYE6lHDZS65pw/Ynrii6yNqUbk2TXce8+9QDacUSnf
ap1NhKNccxU2yVS81P/WdnBjV6tOvAPEf3wKP3jYpa040FMmzNoWInYcmRGTgnGdL4ohfrSxijhL
/xwZpirUq9MBuqc+OGsKUYBLe2dmsoQHAiJWc/9rP989vEblXavWc/Gv9buPZNXz5yTfi6NhpQ71
m4c3L3vULEl4n5Vp4fdQWUA3JgdvdCOm44smyon2BJkcuDvbEh3N0noMlhK4ek3KH9vrtLMRk403
O1FjmllzCxyKwh6dUKH/CroJS+P2aauD8N01t7u5t4CKjVgDAYE90QYP7712ev6bAhuB/C8NiKOc
Z1nUDVnT7fzgny2FRacNiZq/uBqtU9XFP9RYh0IUYPdveG2mjZgwzJViK+260nhekyD1C1V3RznN
ZEMcGDzJyOyKNUeb97zi+W2/XnGVEqEBdWdEq5OflXBmAb06amX8cpZzTEdH0vBoP+C9y+p+J/CH
tZao0Ql9d2SSkj+Dhb9wVkaDPoJrIpKfTj9nIl+04HgXHP2p1CwycqDBdl+AkSH6oyuXvAQz2/aD
AFr1XnT8mWwGYQlFuxMpVri8Q+VbetGEIstAlGDe1hhbj9jbN7s7/tLzPEhMkhBwf/DtpOfeoHGb
jWmWN6QCtDUVXDWxk/+HV/c/TTXi4DPUQP6CL9pVbBaSOvSWixRiD+tnlR90kaRRPyAjnJEQKUoM
seEaidfPI89Z4ToVHOcT/VM19+79XD8C7Cu9X65bZ+akng77Ft/QkakUiatRYyWx9IDOmQo0lAnR
vPSJhBHwIV4Ttx7P2nFykz6W/vtDwtpR4sXhCxw9FKNyT0N6qE/cGKwJegV0v/WH9Kj6LdK9mSxR
WGC31dGwZNnNXHHPXpRujjPt+f0c8SD8+0p4jk3okjbIYCCRXiVTDRECfcPFk1IsrjmZex4qM2or
1f36X+wgDexR+GEf8+4bwwjYErOEpceosA5LVp3KTbTFXHtFfYTQs3K0fYdMNdF7uKCGAQUggDAJ
FGUWVwjdJJ0r2+6XHIYXQVFJmGJ6T2fAL68Qj26WNvnW+8atVv8MPynzbF9HE63nQEik2IyYMvfk
GL82iFm2qKUG0yjzUmQZulYAU8eDHyb7EuuJtXG7bMyg4Hb6xJUormIQY1w8rmWuwgHh9KbwV4e2
8NuHPiuma3Pu/kKVDa7nbij2oMw9uTg8yfRg3XZaRTF/a6FBw/qT0FI2HP7oRZiOiZ3VeUBrKmVe
O+dxP+MENIXTXc2PcVNWalzjouA/jgkusPcMvLAX7kyWBF2beWd5U3iVEEXBK7ehRM7mMtSbfXzu
4RnUVoEGU4L5laOSjaNZUQBPpaSAzecfYvP3lzDGiz2TPyvCjn33xCKildpVzPTs6XFhpOT4Xh0o
l/9islYcy2yejzb1KfL5xPKj3B1Hu99z9wVz43bJy7SLHD/7xCJrYGbwObE3DoMdCfTQ9R2USJb6
su4AdldRCX7f92s6EU3p/PKbJfuo1TLqdsl2oK75bIblfcg+lu+VRCvo2usDcCOhZuTLgk7srvTu
CvtVLosUnv+5ADMOO38pYUsU73Smje2zr+o4jjtX+6Z8fadgrCtbptk/EChOYlFgOqbG3thI4w8C
N1Pc1YXGdB782YKp+sTxxgB4EZWKL+cxLpJXNDgIG3wNvHsqwLk9BUaB2lFcL68vm1vTHvHJDgHD
fvxB+nSloZUCH32FR4XGpZU5oCP4uGP9jn5aXSslNoXI+04AgcYevttk4n8Q+Ggjny9qJeqNM7q3
aptH7/m0aV/q2/+qf9i7pDgqz6l8OejZAlT3vn/Jb7bJvPFrMGLK50SXu9AUJYuH44n7aX1LeaKC
ym/jH31xilbpnncH7f+5+f8Xfc5ST84senUfCF820IXuFQmiQS0lAPwWzPGjisIf22/nxx2UTfSQ
/ASdrhGlwxVZDAPOAOsqhUOVqHMLm6fWuslAfmmnoHfrrFXB5VWaF6E6auw0J6oalqkYhKNzuml4
zVfwJICa3+HQUp2IYonV14sJ3snKxyks35QDHRUxOdecX+Pv1d6mQz3J5HbIPb8ko4Lz7LMwtGHG
xUJ5V0M7i6pqIX/STfzJ8WWPWU8hE7Ze6bNp0gO9IieJ0HOC6V9xr6KscpIzv3Ku/dfB1BAzkINI
3HhI+brmQK9euKkqARBMIgjhRvWROxX8pD3uodI90q83La9BOfQmncnfWY+fAReYDu0xzBExL/0w
bVBDSD4zSuKiba5+Tv3DmeSUCTeLEwm/DgOndm1RTvau/260oXSmHq8H6Xa/TWojqacUzq7M/vcn
HlrKIzKv/JEwloA3XTGhgB5TSSm7uK+m+e+RwgGyUzOhD+JTheXa6ClIExntFE1kH05IL0vvGeF2
7Ll9GWd/m2VN3w6X7GQ7gq26ze4IIxezM6t1dOXaniPw02Jn9u6q/2oXqIzSPEZ1zW3wY4iaC/VS
L0wABDAvdrHXNoAlMP1RiZAAqI16BHEonTQ2Im8RAlyV6GWayYy6LiKZ11YWpNgMrSpyuCPxs8Hy
mS6xbug0WB4PKy/3TqYcGmBS4HNyYhZCiSa7Xh2ZTbJKJh5st77WpNph0zeX+BU0f1T2GxB5yi3J
FVoBO/NdFHeujAWB6Aq5bhh8DPcFh3JIYreJLfNpXHDCJgZ6twvH8NN7mDMssSN1PrnwqHTSE3ho
uRG1hkeTFNdscvtQs8QFUu1fxXJNblY8CH6ynJFkauT17almA4NbPRhJ9C2wU+B94ZDjqzudH4ze
7AVVbrwwth9/QTGBwicoh7QD+4NJlCnUd4cLToV+paCbDx2tAzkk8CMuK101EHP2p5NN4gpnci9i
MvqClOjQKa8CXRrYwLgxfL30nSGqwi55Mrl6Y1dp/G6VtWqwWzOHP4gR4L3z2KSd61IbnzRv61+o
X/s5xXGOV7oaS+K+RwFpR8AZGrdo1mEuQ+dxHs/1F5fWjlHjvAEf2gr01uDGjBqXXsllfHh08qf0
TlYq+DOSdyUcW7kdA5efekZPGFU65jzzTVpn/k5aVCN24MRccnqPBPVTg0n7SSuu97KLrg4oevmq
B3nGWbwtYHl4ksiKxafMxO2t0jt+uXzn4UX8JYb9C1U9AdD3elxR5TWrl6vTUwOsvg/tTwhPKwBG
rzzhj9nySq51n7+ikI7xRT8XIcUCO1ITv4A0N2gjS2VKnWbaAj82jl/EAYhrqLkxfAwRz13PAdzs
+LTg+CVzQlNNrlCuUoihtH8WvPIlF3v7Qlzr6o9b0P3kdkTxSBzQnSQbKGzXI0W6pf208Dzizj8p
Ah21PH4bxXHGtzYBJ6Jp+0c/glocA8b/WrM51Eri78xPuEjldsxTPw7Nwhmn1GEVt0NjhnuqCkYI
46tGvKLx+eKEqkt/VcxQ48+RNHxrxni9WKYs+Vn7Exa5cODJaMf8P3q9wTDiPrLaBURwuoBC1iys
M2078gslahAdxkB+LjwCPUWKraTrz+Xu6dDNOYHzW/+VVJOn3k1Rb0xQGtte65FCPnSICH+ehFPS
8ONVq6Dlu0xnOuz7scyKunrrkXP88dGznL4No3q5nWoG20dpDDB8nBIQcL/kynMEryccdcBmpyyQ
qVylbdy6sheN02d6ylj1HPWusGLdeZ3sO2g88Ocle7EodevuSF1oQ5pgALxldbtEj9MPcg5UMQOq
wPYAkMd4RRVLXhtSO5zPx3ICA3sWX/ObLt9tat5CD5+N8UOD8p8vXu7BiHEPKlty3foAQ1/FDABQ
ge5iTnQhAOjThXgYrRp34P/4hxu7ji1vXALipF+eoBVviIyF7+eSO6CIhj8pU63dUGQvvmOGosGv
KTh49IcRydsEnEeVLbeaWFGifJCe3AuTFo18VQ9mEpwtD+a5/DhmC9FoeOWc6YiZM++faf4DrWgk
1ESBqks5hbiCWnpjX3jQV+Tk0MiIJixHhSB+4QzX5kC9o6XbMGeUpVRwU0ohDhQolRDN0HwREwgM
Eo9V/qJU+bsE6dZLieZOmo5ILFA9sBGglkf8TVLojCLOtIeV8L9NqlpDv5qleXJVlrv2AhofBPUP
Mla6X45A3CU5odObSuiVyCp8faMaViIOTJAVbFPceRdar4Kz4RSeWoRaOS59YqWB6v2wx+myDRs1
NrvWoIMu60w0Eymam/J/1I4WO3srVicEcRx8lC/xr3KATN+Mf4nh86Z9IS6LKlBd2XH7IFJjdM8F
HtnyDACvfwYJZzTr0cObVTQGeqFuiKqMDsMibIX41UoDBR4mVfpNtHWXY4m5vNCAQX3qbe/vOlWP
5xXZk36WUskZdvlScJQCX0od/pK27qatjb79Q1Q1UUrhIEYANm3Vxs3fX2bNQJNriwaOtYbr+XCn
rizT6Yn34Gs3qTqZAFkY6xD1B2vCVYK67216uQgpGQQ4vu7JTvQfbGO2M0sxAMDo0UTTvHWG2Hy0
IH5xegxmFTlSOBl2xirPEcBva+W4ix9R+bw3h/VkfF5RbkssfsQxy3J4JpT0KnCRM2a0zJIzvfZm
LWTHbrajgz5ruMNJAfnvftdyEbIgT8zDVaKL+oOHH2Fge2FQc/VuHmnYtejlE7aqJMheljIx0BIy
3816nj2Xs0CFJ3HnuDGBlhRx76HTSU1m/rrHIP4XeXR1dcPOXQicsENslOgRQc/6pzF2cU7HvGd/
I4pAvRJv7lAtZyC3itXH99D1Qzl7R075HPJtIV8ah4Eu9bmr1TGdpKCKlCyLd+kk39sUYT1EmlxQ
zd0Uv1W7GoEIduwYaMy703jUE97MH/f4hKjNKFuA4e+bp+45r/eUVwxuOcmrJ5TjxZ4ebM2Y28+o
vX82vuhg7g/zociKumea9vLSAj7frLKMkMHOGF2s3IIUET3+XG2tsg3czu3b6e0Gv9Zvnx89W6uz
cBxq6y5GKMoUMzpmL5b82LrrOQBXq9D0Qm8yULdX4CutJGs9uxGBviIjGh0tLMbdHreWVZb1S3ra
aYsRM7GnvBFPdJF1NtsbDNpVKgkhfDQ8EMCx1gaqOOur4qO/zy9+DBorxmsiXAHdEPg74srvvt4j
ksi/1+6mHuNEkKOyetcYvU1Q7hWKGxJsmVqkuTEH9tvCBWup1SX+8Coj7rcZ4XrqqxiUF/rUK/Jm
5RPBoCbcIJngpavYhd6fyZZEiBeEDSktwe0r024ZvZa2UKYx6xIHCt17W9u0paprQeUidLcen5/y
qbZGJo8QAQBS7FCw1b5b0NQiudepFD9yGgpTFWe4dcu08tFdWYIPRvPqBlquNpBW+qZXBT49oVy9
APzcNKoIfVZimaXfB60p15WbBaiR1V3mxuXpBeOms5AXmxpsVIcdL+1g1MSsOETpSJVrO3IBGvec
cNBGe0cV+SQw4TGWKqr3SzcSFWTfLpR3ZX9juRguzzQ92AY3FZoi37OI3D/hncwU3wCOuaQJ3ka2
LTv6cC/OZeiRqEp8tYHnjuN1qFKU8EVPkvAm56ZawxvlNEaZZgfy9JM3HvRiXh0V4rtdQaLfzue8
ch1xyA+fMfpChUIGV+yb83ztqpODCzz+P6X2ta6DOtL8KVqobdYOT2ajJlvul+prJtBO8VFYRv57
t9EZejyWfQXX1m6TfUEIzd5p8ncjnNyE+RA85aoB7laRMLC6eSPoFC57Y2+IrievSypHpN+HE+jL
LwYI0XAatWURWsMBtfsLjtnRO348pP7ZumimpUe6riORjR25Ho2K9tv6WsIM6DwE3S5ey+C9srdH
m1rzMlJKHdlSaR9Y2gMmXReV79iwL/onQ80wNlnmX4SnH7jkHdOi22nskUrHsFDp2HElpkYJuvTr
WxouA2a3SgwqqtiekV3GeomM4aOORAauBPPAUWEPAxxnLt5Zr3jazpIu+T2EJUlfc7WfsSOID9fs
TwbaoGoPNZMCEY/Rj1RhfUratYOk5c9J27+wv5QZyB6LqGIbJFUC59zBp1lSG9E8VXe/yG5A+UN8
rbns+JQ8QJD8Nbs506QWmvFEuPGSrNmusz2QKnHIaOUdZkJ++GxrFncT5TvR7zLbDrBgOpjB1jaC
VeLgEdxgjQrFDf/BZdMZqqsL3fQDvI8uzFCagjtRhcGFJ5+0R38+57/FV/jgrTl/cSZhYIE6lIdg
4TRMX9S2VKYBvdrpgA04F7wQ6qBK1098VNa0Zy5YzgIFQvmi9EOcyNg49EoLK6ICTJ0XTg5SK3ff
+AhNJRWsXwrdkTP9hmLKDzY7WnRL6VaJm7mY5Jvpan+WsR5CaZyUg47h6sdKBZSr5n6oHe4M8gmn
9W1eNFyaQp6Nh7biHeY3x3tau5XrroESHyy/gpKJXTgIafXGBnkZgks+eyyAXe/aczGCvCLpxO/m
HlPGL1J+HWArLYK4/nc3Xkgr+6wFrtG9hUR4AoAkvEmSriScNDEKuU3iFeSoYvf24HozStMNsXg/
P5cawsUcAFpMs+i56/22RFTRlNfjQX5Bd2wmBKRWfMxOYV30mcdeAiqD/8LzZdxbdFsoNo5/zxIs
w5XUeGQQatmlsEQBLbCpF3L6rJyZVBv7GdQycdVoFB7xtcFirBNJVaZWus4g+gbsn/s4M9IJQWqm
14Um0BVCVOhKKMmf+iNvR2rMrs7nLbPxPwNcId4DkdgU1aELlJhCD2jLVWFcz6e513BjMs9p5OGQ
3bRPaecUel9s0t8vKjew17F35OyTwg8bf5XV0C8353OVTYqJaTkxtXTQ6ji0lrWC3ljPhmpQlIsd
11uqnNaBpinYPMndjfKv1f7Jj3F+Zi4uRgQP1NbvPAtMtM3Yx0/J4fnuTojV5oJwYfq3bBwDgJ0M
KOPDU0rm61n2Wuhueqv7jtFxsCW7ZDS/ykfzWBc/23UKO+cqJQqvgzZHY+0hyB3vL14fkCda0AWH
J1mkJ55cKCK5dQXKD9zpnJlfxEdQak31jMZrCDUK18HWfIMtGApMrh8lLMbCYqJR6Et3ZzsfqAKk
+oqLgd7FLfyl0pL1p7L6ihP3Ia7d95nPR/CWTd2W1NCQP0UGHMO9uqrU46/Lfb9zSThfdS9Sn3r2
nDRfgGwUKA0jLWpZBq7CyWDvTZyXGaS5iSAnLIHhzNuInx6/uXfu+0DN9UPQ1Lfb1qdXy85XeMrR
HuiLyQn84ccMpgLhClgztypLFsUYUmN4T5b4JvuJQngVzSuK7yWNquYrPTW5imouYxkRYLt5Szdl
RfHPknEdCOmLpl3k//FC7VolphzsC8Ug32dOI1D0Zh2SH2BtKFvJ3XmONjUAWSAc8JOwQYQr5teN
cMTVZFwkWKWyycxOJWbNMCq+uIAyid0gIDDsZFCbEVBfyh15ax3mlWC2ZKbsuvex0JwQF2DqyNN9
RXLSMFNzPcnbjYEaT6FZe0wGo/9pXJHGsM69RSz41ZfTa4/5u7u3o+kS7aBTaERSiZcm0L/tiX0c
86ZUdQEArORNWQFUD/7d4rgO4ONO/keLFnHcCAWoesPRIa3Mjl2Up/HEDnCpb/ly3BX3TiKxNJjS
E/Gykahjz4FFI3NyccHbIgp2WUbUGUTfyxEyZn3iaigeKv/uvvDR/PY7SUozE9qU+M8+Czze2OXR
apqbT9Y7Aw40CXzic8CUwuLpgSYHgtY+WopIab56c3e3BN3wMuBlO3BtaQYxxilJLBEPAqerg3L2
k0Ez7815FffjUT5B274w3fWTPSYEf5U2jncACXTEz4CAGY0fpEnJH3MG01JPTtnOz2ycGWz/J027
pKHOaIPgPj8x2IFW4ptjlfeehQZKJ5UBGRZUopbcUBoNMlumS05TZpTf0yJANBuaYMLFalTy4dB6
NYWjN+6J9l/po/+eqqsiBqTQiPmAV4iAZYLGwKJ9Vqfcgwnl/uLvwjCu24dvwZMhMHia4Hl5cPdJ
Px4TDa+7PO7gvJyp7rYX8oj/mbjOTUuTfUBoeVZtprXFVvRyqVJojz5FW+7TYzSyrTFBs8QBViWa
fbIYPajo9dq1vlEEaSXUh0TO7yjTtE1/esZd4biPBp2EHEeis3R2y+OsCd7wcCSBh4ulU1pKHNSn
nB4RS6YD0vXCDXWf6TuCt/S41yghFNFVRRwJH7HkKTGZ10h2ys6/MyDMby69nidyFFzK4JNXQsuu
IIoBVLs2t5wkrOGSg0WRdoqovi5PgHf/cUC6cUuiz9N6YNN+pc7rizeC2E4y4FmSO7ZAqrMhG2QM
W10X6OUrieSH4G00ME+C2Rj54bs8wJ77ub0nLYO5zzt+IBERm/D3I3l7RV/tUHMGg5DC1rrjFRUq
Ws2IHYe5USRgATz5e7KRuGb+3ka+NyiKgKG302sb8d6Ujp5pMUsyu7raqUEN1rZG2JOyohJPQnNF
JMTcMDY7+w58Ms+E+BpmFEgPtuWff1JuDNtsPpUNpYDqoxBN6vQdOj6vpWuZQBklaT8v2IMr+5+J
TyDIjSxpr9NncBSvQZ+GTE38X6Wm5GW1yFPNIu6WEUvRoDwLj43rMqzUJaO96dM3cPb9twSC95eD
RI355GeFd8vuqi/0eGo95KoCklEmcoJQNAdKsyB0jHHbsoNYC3prt5oNbD8En2eteP1VVSJioBEL
PtS00v3kZPwESCW7I52/u8vC5uaSkNhAW8zAs+uUrQGh0i5Y99EdCn3dy0OY5TRTp3WMM5KmlPKG
I2ZFfzomyylk025262Q9+ZSsum1gVVxAU5rRUhuVr3WN6km5QT9aYC5pnbeXZqWHzGRDIVHMzr5C
PLO9h4CLk66hTXY3bC6WYI7qHhj9XlcKGBuEDIFHON8tKzSdHpSZLH9hv/CAS2Zl010b+tj584Nz
Ad8z2mlQFoQ551R9VOspecQKJ6H17bXjSs5l2QnncvAGd+y34wNTkt53tzLcneIabc5QMpsCAW0k
Mjhuqqg0bXPeMV87MjaFASuesAPlUM+xwqQAraTI/AH9Nn26xUnunVjod3JdTFeHkn7YbxEo31eM
t8SJRMIYeHq0YInvO6kpPAGOMqZYlPvS+J393xIM6FCnEzuCvpaINHYVnOuhJr5LMVLv9VNsOkju
/VB44Hoh1f7hhk6nz9OygKc04vkT88xE3hw82PUyqal8i8EOtRhqMFV8DYcor/quXB17xKykoESC
HeH8krv/X69EznSpPfvcXPcLOB2K8zOyuTQdS1LAvjd1RPXUctLmyUc7jctoRmIjPHNjThRyKbDw
cEUCoHBtErraI7iT8lLu07xRh8vDeU9bXxy8E5wKAKZU463+xxq72711xBndwl215lg9l4kAyuCN
LFKCzY/2xXLbjxnSJyR2lOm1yWo409O/LadtrFo2Wip916XHJfSnPdUM0gjmnMLDY+U6oT8YI6LL
TlQuuMkjV/81k+nY/+MkzX1Wu54QvXtJQH2SL064OWXDBei/reE0PjNyWihY0eIlpWqIsRAZBXqZ
qt1FjKmps83HzLMzvHZ4ORtAdi2U+QArSUei9Uy/lPrRUVx3NOr7tbJdZLMVjnwro3+OXg/4RNPB
wvpAeieiEmehT7OYlC/0HOtroMFPXAHNiqF4D/O48BifDAcxCWvF5odK9TKXI7QfiQnIhjoepDqw
0khF0sEdU1ltpgX4GwDQBXnTB4oO2T6+/+DuXBmYDTNxNJhPyKXd6iPvn/StrzPYCFfrvxAeWsfD
F8g1ktZ8sflTHoPS1XjNY8O1T/wj5Z7I28F9+iT0ZARCaH3mpEnDzSj2y1LOqcdRAuM6Ev94UO44
6CsQXBH5d/GPCtTCRwkgYOvVvSyIMYb6FXicVpmovLhClsk3qkg8Klcn4ufoVekPPsrVu9OSZrrJ
oIfkfAiRZWMOOfCyOhKghAwYsgn8B9I3inKk7IftMuTkJomZ+4nB97SLVCWyCBnyxtxeYesYC+EH
gYY9im+jzCWlyvVK4yaueu5CLm/6FCjo+rBSfDjC6Mq01SkDDSbzxcMtBVU7VrB7I2NOlwpSqpnN
d5N+tHsQTPix84HrFW+NATpd3hFz9+Z9KLluhm5SYYJZCd8izTm+tGFC80nlM4A4G11EjCOZwOJ9
chTf8AOaCpnXNondtnURNoiFCucZatmKn9/uxu4wgQR9vKsmwx2+XlKJJ9HlXqpAFWNHG8thuKrY
8LHDsn/zkNhVXwlvWsKQmIQM4XHE57Pxz9civywNfqsFRxbYbu+wZjLSEEegolOHoAx3VqPSy84i
cN4GnVFXKqXpoSejMQyaSDQet90rb9RiCAgKlM01j3qudBIgHEnKVEUwkrBOn+owMfNN7aUs78u4
+n5t/00/pnKc0UIjdJHgpXBlG+ZOdExjZKdOrBU9UCf6+LyOdLa7m1Z+waml0hq8nlT5JboSJtnD
zYzu0Nysc1aNmX116ILqEVhuSOxzxAhADmjOVcnglcRdZiyN2H6m/qV7Jo+CenRsd12PS+IlwScz
z5KFe02qr6pdQkT8/d6j+/EvRjEdJIdr7LEO9/y9HpPVSGrhGBfgUS4f82zsh/yh3OX1tuvy10DG
GD2TImHMTkIY6DnkzCDWebhGnpagK7kWTy4qsQfGKuWj++Kp9ustNdHeS0H5ucwiTKozjIRvyAWK
yhT1HDR89USgJIvZhjfE7p3RlRvmHM49TVHILYUUVaZ+4Efcud732V7rKamgYZa2u/QWVFSKk7vD
YRYeXrcPQvA41oizw1fR9H2CN16cNoj4iDXLyLAenZS3tpfid5jxR89h6IjIWH2XY2R1N6PAnsQk
dR67ijOT+OhSBVfX55uD7RuCMOEWf+pJEy1GTFgsiM95+JK4OQeFVvg5dMsamna9JJnuRrV6H79k
3th0W2fslpH5QOlyBFwBNzIWaTwNrttPTz+CzYqw86N2hcPpP/3nXmmc9ac6CV9bxK1iU7/eYt0B
9fFRLchbjcUT1pxZOxaWqvo0Xc4wR+4L3yoxAMPugmCgCAA7xigScN4YdrtZc7cOX7Lo+AUEPlWh
cSAy9voNSKt47tHbohkmB04+e2ghFXP1lGY1II80n6npz9/DvRENBwit8pVxHusOQzb7JjiB0MSU
kLwu8RWrXPX+5Xjc8xbQTq/IvsTWybX1fgS2ox6XMHGFttWymU0AA9qWs6ZtrIdJpIRUJp+vD0uI
dCsHDsdfvgqATohM7RP6sJQdrBlGbfOXHsNUhK8Z0h5TGvGE9umElY5NGkqyhZJwPNOq+uyoGwo5
225XsnTXeSvBrtWYJD2xpyZhx4s4pd0+2qNsId+qb3KAXr3/RUQUXvH5Q4HOOOGiEMbPNB/OhNrw
guaKXQx+s+s4WcIVDC0c4a2fU1YJbV9cTbEAADg8tj2dCOe6iRkkL6RfjhkUgMBO6BxjSnuOD6oa
iuCLU/i8nlslX9afRbQHqdFEB5V6fPl3B+H/zIzNhgxRiAJ9kzRp91Nkw5I7Tdinj9rTpnDzmRQp
qFr4zKgVQUKGYZhJtJF/6ATF+j3alqOCd62owb8wXPPHP1lTBEfMy0hTko0Nt39JY0SFtsKmW1nh
OBggkcKC4cRGMK3hiE+fZuaG7VWwcXnUrussOQm9EmHRZc8q0UPJPBVv5ovq4vs5/fzZagq0Pqy7
nIZ4UaqYJPtcVPlOnLw0ikWT8Dh4JzBpSLiR5W/Nb9iml8g3tL4ULVuDpochSPuy39dyxryVMtOn
AQ6VGJM+pTlSQh4ghOa5xhPUXmqaVainCX70VQ/O+LaToRFfmXLw/Cf3OwWxXTz/QJ6Pi3D725z6
7ze9tIMisrxtwpFH6sFkSz7PDwSwyXYB9OfT7HzSOyXf8CBJTIE4Y/GT+U8F4QZp5SAlXPhlqsmK
Sd0KfKiJEd3OOTpLl9lqNOSF+Qb1YUgKPTR40E4QyoGiMr+ybzGMGhII1ShtmHSp4+N17fAjZbFG
KLM/FUdVSB6eYwrXWpF5TSM80WSkTomjgtI6NTYtW/Jo+ZbDo/b23Ks8+nmdJEyeC67IeoQNSyoP
W4PBQRRAHr7aiesERkXse1L0DypCnc+9nqX150zD6SV2WCJIXS95EzcIRaBSDjXAkItXuHkSTgp9
zGq+ndZk/dDui2wtn0ieNj9yWQqyNqX4vyPfexVdmXZ2Os5JVqkbKF2c+hKtBbNPerSciRLu+qDK
fi6USODkklF9hId18KqT2gZd23PFH2/0RGHUOYGov9JqKbI7BCm7d6H9BkyFDKhb6nMF3uWwxN+q
UOEzXicUAjOXfLTW/0y4v8K4uxHx6WDT1P+lWz97gXnA/HNGU3q8poEeZ6ZjtFP6N2Vr3mePkyAg
12kaL3c0UyZzW89ftveFlvkFN9B7kJkfRCflCthV8FQ20GUbHcAsNxZms/vgMzvLX09vF/XEwNJF
8qyE/ijFLxv65G7T+kII6y6FjqW+uDAXXKcDIz6Q8VHM7kNyxtjj6aOucTLC8BWwpxeIaSqbVpBb
Ebm7JIYbF70kiqphRx41SzWz6lOivsrlR2pHoH9IYMbAzbsgSsxi5rpAKdBieHXskTUYToqiKjg5
zNyFg8DzWA3w8uwJE8ye8EaHnYDUdlkPeNVzwTGdvYSXOVqjRU6uRNFADBZFuAAODXzvpz97WgNr
o2CLTXllVuMx2gvkCdLT6FMU+TEPC0HPgAd9DccyglXXjaBWzwyhJRoESbp5cYH9cr540dBi/9RE
9Q5usVjpQ+v/yz6/ogX/PupM8+hW5yoejc4Z7Wf4U0Y1J3bZEtpW4lC/SZaGjjQVGcTvL/dIepT3
LcO8EKQeqULcYEGG1VL+isLphWCx+x51mXE1pmpDfQCt1QTxMsC3uJerQ5LRVuO0Y30+rymQW/5t
n5OJBy97Y5va8yPFm84Kj/jvHsB26KY8paVSLrsmriVhAp9EJ1CKTzP4EPeFsytO6tOY6ntWAhsy
c92P214EG0Q1IjAdIIFq5Do4Avhs8H7dfoTKpQx4wGedfI5s+lgI52WZ6/jGa5k0JVk5VPl3k9OC
WBcVOoG4GKUnQdVsFFDx3Rwex31M12SA7qtYUZ2rNpI9p9vjaX1TPDWqjCfEPRVA2PcbCvSnCbBn
gPJWjk/a5M2tG/Plm+wFo6AY7dP022gaDFhEdrIk35PcwJQSiSE5Tghawyk5s/wWuWfFLnlhq9Zd
PH1fPQSvOgGVKe6XH7TJ+pIT1w9tIs2IifitYG+csfdBNF71xx4R7xqDbGcnFonwrfaH58+y4wOO
5gg909NTXxaHzUGk19KR/5jge0HMNTPeqw+MhlqtnsDg5+RKNB/t38h4SVhWnjkJJnjJanM71Ln5
1MUzzF6Jt1oLeZpEs6HLGawG+E+nWmzytqtGMVVGfC3+tR5bRLHG1yN+YZZOB9fi+vIZPWfG8UlB
7FDW4rCb564BI/dXQmxCPP1M1UBWyewNla0/sYJoU8VKRoiOptYpOdpimNnHE500p3NYUE+8eccF
vvMagfKiNXU7yviFDS9fHwOhuzncoPjQ5f+DXnQM8n/X0eiawLqHg+WtuX4Qk2G+OMUdTdClgpL6
Eme283pDF+pk0JogMTS3h7/T5g8z7yQCCihWGFRKVOcjlPaOkCZIJ/Sw3au0HS5mcBLJ90u4iGOp
BQTAqDwvTMeesAiQVPe9YOrfenRT2NXaam+uY4opOdMCnysXxyoR079Ij+yCFiitXPZHsgtRt54g
5JM+AUYODOATF3aDW+DQik+PCzPb9m/uagcXvyNuZhIdnv5c2ozEmcIv3p81kxN3VRSk6so9mUrS
Sl6/TdpxMZOM1w3hA55IojQw2eEDpzR+O2B+UeO0lyj5pnjbeKoDLdXOFR3lQTfsY3ExjzRy5Ij1
4Pzph/3YA5Wm43Ok3TbwfHIaWUwKir7mz8v3UWOgTatHquMi9uzj6CGCX4RE6a25nUhsg6hJewgw
1wIp5sRGjrS2Vk8pOqgTkgqv8ZC78qviYnHmyYGXkYh+TYEWdGF791d4NF4nB1FeppvZn23dRWQI
lqhvAkCfJFaU1tpsKpNkL8QAZuxd9UmyvfOgrq1ZZcZt9ule1X6r7v5J4BV3Vuw4lWxk4AdUpJPq
4c43ugWxFgr04ZcQkJEtZx3c9qEhTi5q+k6QCwusyRTQkMPvqGBI0Fjdbc0q+M5IndgMk0Fpt6XS
ruNx7xYlH7uga7Ucf0j8H9wtYhKUxg5Z1pk1a4HUz0Sh22mRSAt0OAuj4Y2QAm+91nxax4EG+eEE
J3bP/WK8h4aYkEa96soYxTsChc4wW80jv3LfAd+MEqNRFRNi5nrV8d2eavQMucLUkcdrOI8wCL1/
3oMF9sA0y+Osi1P+L/VtKxJNujg+Acln8EWUXD2Oh54wfbG8W/QW3gwoAJcKwDUnj0JP3LWU+gwG
zXchPwZ/wXd26alKwGJ2ISKHITgP+K7moFmUH5EPqyOFtseZd6ku/wZqTDUQh6/uBOlg/S6WKbQB
+V9nLhpZLA5yoZXIwfGNq7cgmnZFQMHzLUeukQwZujP3Me2cZG8MULcYUk5CCoKD6fBgtAlUn6vx
CQFteODew5u1k1plvCdTo0UPnxcaooVxuZAORe5NXgWRc+FwNtbgaJnrR/pPZruyuNGXfHPUmV2j
ubBQlyJwmK0UuCYPtUQhUMPKvQD/bYGJd9OOxKoMhLT0WjitjwunWIPhhjks86pvxMcmM/m2wGcQ
qmUYqfsv9lDDQQpF2gH3d+82dq8/frb1I5kqriJsNsQrYFPU+qLRFEPgse1eT5C1T5lsMdy1W8Bd
6GHHcpmtbRD6MDlZ7buUL64eqKUr8Nbe5xhB7ZmRawXstZg4RlycZcoLCqO/MXN8wcbazHwC/4QQ
LuVV42nRbpmUNGmaQz0qADhNjSNv9G/wK2EpDMwOax7Zl3sDvxkrICzE5XfJGgRAPGdy2/u6F9tH
2Ns91+fJvuwRKft9bRgXDmqs95FfzlNoZc4UCpDDJpzJdXLQA7zmeScQcxvweKNbI9sjxAOKyokJ
fx5Wmuh9iRuZ3IhaTyKFLVHueICMWMwIaLxu/phmMWzA4u6gqGUYLblzXlWNGR+CMCnsQaFeKMhT
ct/8tVe12orJDJpuIBn3OnUsUM3Wl4fQN0BIw+R4/Kpkw9UOfsVXHGTc61npu6dLn/pwAaijSOM4
8/Rvrjz+J6XqWMb4WIBJoC9jq3XViytOIPuGCqaf3L1ALEGGG9VsTvxRlK1tUIhlu+j/bIg9HOZO
GDwmpcVpEzUhTkTwasOPwZWdcvxzXtlg+oFpLg8T/BNrEkZdu1I4ucZu93pl0qrUpeqau01hxsdE
nwv+1wCRolU+ewDLg+TRNz7uvL+qn+RBP6LzMhKGxp+wwx/RqI4WTFAx0fNTd1Gpjq5dhy6yp0JV
42+1NpU85707DSSmoKhukKWKWuc0jwuduB8HRKzgegpPV1GRo88M2nbMwjiIVQi6o8SJiitVXbw1
x/hBCQ8W9oH6Vy4ITm2vUGmyFA59ZVSL1bS5jfPLS7ApvZd58CSg3/BaUBgwP8A/xsssKV6qF8zg
n8E3CIk7adFmq9JCRgkrk6ShawRCTWe3jICxz1RojiEPkyOUCofmuW+jh8qYrYoJG42DyDAdw8fF
2Ekz9TdCQNVLK7kzatEC+Nah7g3Ts11rRad9GyP5WYGcx0f9wqOoOwrTmRxICrPMh8gTD+qzVg+/
bIn50Htzxn3IJ60PVApniKaLp/WnZzlbVzuhr1m26qGP1g1CSp0DpwHLPxZrNxd00J39tcUVU27e
DtUFkrq/Q9SlUq0phXqeuvbn8+f2O7f/n2Mn1fMaSCfM59nEU9NBq7sNbIsyqqPCXEuKGt1yaBMY
9GoDLHxI6Fxj1SC8IQHcN9/hP8qG/l25QBkKHzT629uFKO8BLBKEAMHj154GChDRD2uRbWIOuqLL
qpr+URyODeGOctnrncqXJWBht852z+7OD65mY32FMXnkl/iVSKXdpqI7XS/nLa1IcMDopIZ/hwsH
SE6WMet00BpD/Tq0d1hv1UF6XbyMHt6i9DEPemvL8XEbG/GQwg0CmrrrtamZhee8UKlNmivkrfE2
5cqxB8IoRsiB4frFyrYluZhThQRYc5lDsCYO1F6be1vkVSc7/gyVJZV4+ovNCJBHP93dOE3+WKgl
059z1XiBzQR7lEDSWsnPILOyntGgvKmGR/yAUmKYBpRDLE0Hr7TgzsGRXC1JzwWEgs24ccvJ2fsW
3rxZd7puixx2x8mhObnxIUGfUIQycQom/vIzEUtpLFnLLfVc/OYHw3vK/OLiEINcNbSsjOJe0XqH
GtQEu7EkHAUWYdRF7aD1D1CEYlbjhvbB4AauLb84gJoXpCl/aONwSkNmVUPHg4AQFGhHWiM3lVpa
iXgGHzItzh6C2IP3DJ5VpNpd5qxtBARqPh7S9PwLg6rq9JhvwAnv+m0MZDyZu2v6keZTYm4ojDfz
m99CJAzJ0n0wX7QiB/n6xcwneu8rSrcX5XkfRoKcjxzzHgzjUZAhMsTIevzCblZ7ApDX2rpfd2nI
QQKoI8txmkXxU9kkbbec1KwrsDm+akCzjBSjYnk2Ox+R2Pmor44iX7hTVbVJZyfS9gHlIDMiO5dP
PPBoxwXYkCDGRXSE1fd7h1ZSBjP8noGJT4vbf3QxepdAoPBTHEQ7xQ1lXUl4/0bTepxYUS512a5m
BcIT/Sa2yjGQx1K4ZyW3iDcu9+/Bj0C5v0HyV3egoe4LMHk3m8bQBLVIOyHxTUl5DUFcCfl2BptA
BPHAdsnCcj3dH75Eh9aZrtVJ97SGSJyqkXgXV9jO2z9Hlyfvx1UfeCaQm4W0JaAqHnLRw0e+dUoA
PScb4lYD/ddim8x2CxwIR7pEEedamEZlt9kAodRe2YWAG5LclRawhNjf5NiHWqoIGlpVKrZvF0Um
v7Px6c8Mf0LE2q8vUZIQFq8Gvl4z5JL3/fRpA+8Crl5kn+EdPwHF7yrd9/4OgQulQlSvxG01rYpn
p7c1P+20DZOa6PBpt+JkZDU0kcgTUUX0BwzLxbldzUYOA990t33RHI+bb90qYckU0KdiV79Q7Z2q
SXqtPhv5k+UYShcIHy03AAIquy+JLrmL4vLrFMohMF5P99TLcn7SSV2mKhTcATqSPdWeoPY3qtAi
dlME4smBkkqtvoXV/BzNzWl19p/SwUdom4thZIH2aPwvRErwH3Wh9Y4x50O0ZP2Q9fg2MPqP/81X
hpzidG0x8mZoYni39Cd6sU6JMpmG4Y/MsGSz32naB1Cdui3AuncZRLFmHuv5allNNoTU38uIeNNy
g/F03LcObo5waYDZYdQMTulNLjhLahJy/kMNzkts75+4PhT2RwqIDoZDqLQ4jlh+/fSxJRJsAaB/
Y0U4HYPJYe6mePyTFm7AbzOszq8aKPlPVXHMoaqC+pdTyTDeuTOFiqXn8Er/GthRjSKFRPrpTsqc
qWQFctPtwXgPZrJuhBkFAxrwXEdo0BwreHtkPoyU2TLxlEiiXc74XN/Sd46UBpP/hxqQgMK43tvb
mLciWc4KwK4FFRur4X4hXIVzpBBpFZuwJEuxjQ89iBStXYiljyfDqG4IWGj+abDcsz+8ud5qmarX
sW9vMU+kG+t2xfZksKpXSaxS6aesXg7zZODVohPSXRG+yIVgTkAf0sUky72UnCRYU3utSGRyEurM
xfsSqDZQf0se8sx91I7L20YQkhv2X4yihAUVGW3yAm2a4oPF7j1vCEkzwMRyrCNwJ9UcbQGpVfky
moyL18IB5BdsgH+26dSMGKHrv8haoSri6P7ebWarD5Qrdf1spy2g2Mnpnur2jESabWQ9CvjzYLN7
r7bh2E32A7KvJOJwdU1P5neG/AEJZLMwd3Qobg2rrYiYywr4lfdQZiWvf/5rRXgpz+RVWjzF6oqf
kxmzMypaqfzMUzdB9HzIXnVEf2cX/kYF2nqe5YIQBZS5ZsZfAEZxgLfEDBoo8EzzE6a5Iv4txZsb
Kd/VoYGdqtZkKylFw6a3mu+Ba45hnxOcigokv6jQklnVznv6OV1hSbF5vXQ1e0jLhBrtRTgHsRdg
FAzXBdarauJK7QLMQRkxvzHKL3mq5b1b94Zrv5vK1Xxagr0ms+pvDQ9eBMnp0PMR7A6nNG7cQd/F
prgszsKURRZEnGCGyKX3pE5vR6FpSHkHDu7wXIkzRy123AKcllEJg20FhXJ4OUBScTzuivh64uUU
u9sLXaVXY3IlG9lrlFG50G1JfqOegS59gJnD7w4JINekdz+hFEAyBgHpJc6LQTWVQz/lqZkZWI52
079G3FKTNDg+DYijAkviuf0st37OXzOFYmTPeAVGw/v4jCxjq57DNGUjuehIegAHabrUm3kwfG0o
bBqCfuz+TpB+HDEc6PB0zKmgpMvXPZFcvp9z3X+3oZMc1fwZcNQ1iNG00eoaqiLGCDq22JucX/JS
H6dieXwY1UgnxDOuBs1Pp2vniAYDIiKXl+UIJLS2KFvMGHpIKC5oWzFp4V222y21ibyJm445zQwa
Ps81u2M2K5vUUPSqzaWSW9EES3v7NQsywhsTlIPZV3nXIa3IMpf7I2LUaZMA5119GFnrgPwzulxy
UaZ2zQT/Phz+v7BxE/jOT3D26a44WnYk1hgBslqiOH4t6+2CkbYGqnze3EtIP5xhfI5ukOBaUvBH
+ooT8C1cXy2CGn59TbqaRkCbKbdr4bhC00vhCW/Ti+DUmvOc5MJ1yK9HiBU5KLNKdQ9Ntk79hmYG
9C0WRe9XK3r3XFv3rOGJFh3786xqPIDo5t9JifySKakUwxwL2uCZRd3cCVESeCOr54id+IHc7wyx
96UYqN8z159sG//Lp5pXpBdFFC5s35+ySsbMjDFd/qi782tkZ+DQkwftJeW+9aNdenXEi3sZfBrQ
CxE82TXoRCBCwOhh0EmYMwErPomO5nlQQ5BtIosOpcrbOCfes2tAWwISr4BeYz0MuOPmgdPzEpnR
BqEKVBB3QW6dB0pyP2p9nyA1BZLG0sr5yIBFDkOHKUIaEfuyhEB83OilmJkOm6OW8ogx+96+Ekki
AzzVpP1vSTMqABR+yrQn2P5xFvHPM+lgSIqjfYPB3bvyhr1IpxHN5m+8VFtgL7UovxqhMymlByRd
IItvlNA7KOm2+yY85i+JU+0n2BWK2YXvhInGksSew2fMu/3BPvgDnBUQ3/CDbxrdZd4eSc/IcAFi
rb6KnisesIKyqhaqZZYnLmwCcFJaOinar0mo16yxWgIst5g5NAeHOxIbzgtEK/cRQ+J8atX4Ggh9
gPNdIau3/QmTolc1Pxfjgo6lkn7bZBcH1KmJrOJdtDb64XT8xtIlY/nbCVVh95la6eeBLQb7V1ZO
MxkjdIxJAMZZThjnXIgddwDQZZVyG8PuUr73hHqf5xRF4vAjDCuj3rgbaR4Hd+52KUPmT+2W+rQs
DQkN13KL92mVpo6Gtmfpl35mpGFAatbcG7iLGI92EmmX+hTLkFy9jA1d8I+EBSI9Wt/Y/FaFHpU9
rXLKiTBU93stMqxRJp7C2I31vK6JZAs7VMeBiNM3wTMQErlicAreMxN3vfAeSWe72XGUxaTrptJK
m13EsSrwJNPivnJeh3w5xOc9EOqdOaRdnc0amMPNQ6i3rG8/XTokUW3nzofFn5hThoWxhA2RNhuz
lOCCDmY2QOv7zgnFvwDZAShzTt6SXOkFXWNpKhIicClX8vjs3SImGnzwLW2a/vkUcEYMw9kRwg17
q+dLYMiNYQoRCSIvcoSza6uSh4ZDAdEN3Q23t/iSM7E5STUvHZ+U6IMKvaHKj6Kzk72a2C9YeLxm
bli0a9vA8HsLrQYvbXFeWZSyz9d9Z3yIIn0ATEuHLytrjDPejOFEDKy//MPhjFHZfsjqOOoLKyhD
OvHcuLNTXxbPWrs64Iyg2A6UU2plYPFJUf9K+HdSGBkmQQpMXxXCk0o5iAvYh45/HhU5dxkWmAIl
DoPg9aTW3zasmMlbRyeNBEX6ewoNjjjXvOx/Vxej3I9kqZgxqZct6HecKebEYT77NqaFLs8o8K7n
IUlqwyAYEQiR0kpCb+XQPTs6a8/CB5vNkoCMHgwMS1HmV7O9q08Ia/CqxtfwhJ21JWr9WMVJpnpn
tM0zvSnTJcOKVFwg5JeHNJhc/oJCGsOQV3HV7GXN43OR2WwCA+gaXR2flFF6lY6vtJsHfpEbiu/d
sK5e0sq1G5ledc1HqJklphjSJg85WvXI6kBwp5hFU536QynDoKgnhrjuxPkXVpol0u+bQBIJjgLx
g3PNMqGwaDMs4pyEWXsenoQfH987FcrZ0fivxTWtE8/pQ4wkIsMtLycBCIYI+dkgI/AQ3zTNXIkv
BzmoYYBvd7ZMBpw4jadG5SV0qtXbixkD/qJwY8Mj1d4fNse0ciDXXzNOJES8iisNVTE8artSg3ZC
I6YDLlWb7l2YpZmIpkXTut+y561T4cH0dT/ZdOZYRW5sk07+fHrYosOF7I4cnQY5Z+g8hSE8tlgZ
Pc67981zpi6GFi5LB2Q4dyzC+g8vBGXZAaWtnpRRJztPDzuXiS+WgXusqXcGCLiSM+WYMZkNE606
sAUG+IgFFT2m30EEIeVSZyIKOpDSPpyP6L3RsXBzJEGbRgo9Da55LVG9OYLLS4+Nc7uexX4aJ9EH
Ay97MZV7cLw2y2yFy28jtfApKBxzZ8goiQaKOd6oW6luzPJ42iuxcB8US+/21Xk905XuyyIPXf6W
Pv4e3CJVnGZlQHIbwShzU7CtI9Y4PWJw29ijZ0B5J+TkzWWI3xXGO9BcfFj8YAltYNAvwEDRP+xE
x4HJIsFxGy6O9bL+6fgVqY00XuDOxbet4G1bNR4pVXi5VhEAyijw0LixRY7tXcL8KLTnbUWd7VLy
ShAxwF8YgMTDjvRROO7TX1zy2nuSCWjSyUHqCZqNBCx05x2fj55hYhlLcUDeURK692Y+F3atT36Z
Kb561UoQLO1gUj+Nk8oDCEAsQq+Hq4QX/fuCkQO4uOwuXhic6FaHoUDDs2VehlrhBck5tSYXw7wF
rebdDkNB8lLEeu/4WtoLGB2Pi1xhlOpewMVZFZWFpxBiOEO6UNRClJEKlsAuZVlvzmpjmmeFap08
2YiAOcD0Zy/L+STMvfUtH+Fz2YePCcM/WgybqAp8BtV+seUTVwkUVn7CgbYCmna+/ownmUkVRPNc
VKxyP28Ot/uBokJHaOFPPOYgs9/wTYdsHbbtN++7BnkNtsEyPcNOjSdBiYTQEpYOueLYwyGnlCis
IK11QEkY5DFXt65L5Df8XzhHF+ytKUt1x3+/dckCe5CzXDRJ0exHircE5ukElU503IOlhvWA3Ml/
f1sfwxzKl+yAnKdjmab89yfo+iPwNKYG4i8jiRpgYrDhG5uOGPEx/MbG4FW88Edm5YSveq1vPOfo
mTNQu71gX/91QkJmUyy/zYXwjc/0IZJyj6Q8g2MmL3mgBpX78LkvwCqFg/LMc6PO4IxCXtFaE24M
DOlYYXbFHcvOTPIVlsFISUDG/+CkvZ8pZG83TjwodjT/6x79dEJ01uprb2bAgLshUH+26Fm3bsXG
Biks6lY+bcuJK6sIE1UCvjz556nTUMEHlEqaj3ZhcJQ5Y03+BPMjEM+rYIcUWcrFkD3LAAcYQHzc
ZaDxcehNTR6CLDmXu5BvxEsPNHy9SzFJE/uv96EvU5qLOedq0BoyJXehwdnnlZmH9WFj2bRpE4hK
Ry5SEsJlXOYtihiDWOc2pWu/paKGDZDEVt+3qHAG+r65oc5ERbVjGejS1Xm8v1tk6T9yBxGc7+cI
QHK7Vd2enp8/DPbFFi13t9LvDSuyiV6g3tCCdh1tLJemrnHjHW6wWbgOFlarkriVpic4FHOlLWtl
CC5cr6igrN7MT9V6y2Qxm+duqz2a5Y8Fnoi2aTERUta+ckXAAkXsvQgDt2cRPzR83D73bnl9TOcN
vuI9eav7vtu5ct7jc2FqM5gqETkAd+PXyFOtxYkoOaHY7L0BB1GvbpRwDQTgFgN+X5rpZxgE9mKx
yOjYNlabOG161l7KVn2cqrAs10znrKmLa9GhxKBcGayHResBz3BkD2E+E3YS8AAGBoU8NcvjEFuA
PXdnfpM054RcLZfc4YkoBTwjC/wZjGA6TH3bEVg6sO0mOanTixn003eKaCM3fQKA5mx7WUYojy+0
5F7lOZZljsdWzxTwNIxEgcbKBhX4KAkCmulLYEh/jgEVd62G6hoH38FvJE13zO0BCVy8ZNnR708v
7EKnUWe6o10WVhCzeDOf7iz1xJpaLTdw7XoBXR01wor4Eg8tIhqp5/x03EvJ3FYquL/NjD/Hdlul
HLH7UnIpCs2pD3pAcrCnvF6F8NAyqgA9SdSLJAHvdoBQ/Ee/z+pLkemJ7GVQ9IPGgMkyOQCBBoTI
3a/Wa8RzcD+O510oh3WI+VuRy7iGH0BJkVoJwUK6WRqqPJmbFL4D+zogoIMxIVRcdzuWg6mycPdz
Rn2l0C2ldT/C5/9KCWcOpVLo2Yc0HsWIcD2bS3DN8smeV6t7lhAzwYNJL6fM1LF4RHiezoeJf33i
LW8j9H5+0orcWYYmX6/Mf2bH6BROYzdP3kZYehF+ROrGxWftYWEQsvDlsO0oH8cyV815XX8yY9uD
sdwrNSHtTq/ukocTUi7T+0tMrZGOaL4LmXd/4pcIlvcvKKY1HsNIHL7NuPICOsO92ZbuYczQHU9h
K/TjexajLCX56NeCNr8Lj7DyD0HiLlwykwzUGdK7CAV1jwIPMShDfyLVPgUGAtPwyLaIAlZuuvEd
+bKsxw6gUo9w9BLT3ioRvTLBh9s8VvnVN9iFG8+2fmyPabHM1CYDw6qdxRl48kMO96xu8UjGlLdV
YXwOZBNvNgWnwVKlD0PskSklXhyLzeTMSSw6sP/8qoPCD2Lq0bYs24j+ytbc1yU6WHTbCAks4XEm
Ebb11XSOpBBGDPOey1nu42dYPpQcSy5bYIJ8tfTt3230DOH0Fdo6MXrgGK26Dy8D8HOihBewAhSg
0IupkL5xcOuzEP8BDPkfHNvkntDuVFkiZ7QU/0Ol+opnIEFpBk1zyENeFtjHcaTVWhJ30SRYUrQ3
MX0Ny3Lg2I1hME7cahdpAkVlg3TDvU/wjQqEs8hMl5dFsEY0afRW9FylUTto6Va2Hv/wToz0spT0
NubscSG5k5/ILfmMDg67aaJVAAJnO8xS3lZI4TQEpfDn7Kou+yIDWi5rXMYesAZnUBLJ/np4CXp7
zVrNTHt1cmt6QyYx/tLI3fSz0mp3zjJHM7GY54c2KBMaFOrsWxcqvSWwn2CsfTCPP6eI7Szyt4Ua
tOIUA+t4CJ6KPTHfWUBHPUk7NbHkI+cb7cCdrVFLteKEYGKGIMGiBSnyv8pW/nPj1AtVp+VF7yZX
mGNU32U9oRibBctcLdJKMo5c+wO8jrv6LDuOzaTkVsl5tdytC8gcACDPNnnQjRvaGefS1BlEhmJS
UVpo9gvtU0EiEl5oRn4kcEWIQZ6Y8IgcPTXTDU5NzzhM1rjqd1d61Ldu1kGdF6UoEpgP78ZCMbdB
bBTKELjK9vJBEKKor5DNYuy4guRlitcgCdC07IXj4XXfDD6FB/8UPedTIzF+MuzCdMppg9dms5Ko
knz/8OTG3FTYdALEN0JwvwKb+qBTYxhef3ZBbqahu/7G8AJiWST51txpDecq7cWKDpPKVTpxIkAm
89NxHmYGUExV4yHdGvfKEBOP21KL7apJ4JrhTyKbMDlDabBWtUp2lxrKANxOyUgl7HrF/e1Zmh13
vWWIUDI56M4GWO0RQlONOaeeBuAfKKLg0+PNOrB5fe8qKoDp1WzExMPAPbbNvoEWEXwC5lvdL2bN
35aKgIyjBXI6Phx0gUOmESbL0LuiA7mRhzWY0Yrikf45B8ytDbiebvRyK/4Gl6DKthcTvmBK6pk0
tXBWHqxC757Y6VYSO+d6q5yH/TvZfPFqHad5rTBNIn3rQypmoldcBYc30YT+u3SdYZI2KuZJcPUw
OPmYoD5Amcd2GbTP+kvYws4id6B7geRlXIejGrrJSSeMkSJZdzLQ1tRb44DJefeA8YlDwcuDzYH+
92g361BLF5OBMECbyZtRpO+sWopsRQb26Kbe8CYuf8Tdk+W1GnRCm3b7M1ycjQIfQhYgvKXB4snu
lfo9H4PaUvrK7NDFBzsbiWzmh0fhP1y4aI+jOGJYo6zP3MjlrHhAm8SvBZI6xK9LMOyTaZo7Zr+1
yLeqIBLINJA6i/ySCW6T7r7kSRIgUiX5vaXYt0x1qStE35jQsQEpGpOtyaJ7QhwgO/jI5l0E8sq6
pa63B1SjDdHQjkfhVoiViQtCJIJQfUsl1R1+QYNwvqxKJRxRv3+t9Bm+VJa3ixeu0lggpSUnKfYA
Cc2UiMBP8+DOQxIG6gWgrynZSp6gwQA72gmguLEP8vyiQ1J+IabeeqelbTDvMEAb8r/dd00xMNPM
2QRDvmmh0/npNImbxALdnCH/8+LjNvcYcMfYhG/tgNgQsZhO2rb4uo6LIRJ3P/q+PpQ/f3PQXnSW
mDCiXR7HSjUoY2A/1CWrdGiU+oHp/LZhZuXppAan1VYHP4G0KZ+WzJigaJTsjH3i4n3PpqDnI81A
8U3XRW32+UVLF3En/Qu6o6n04arsI4omgSXkFb0h9r6J8mOCn3a3RdE9eUHoZ2WxbJq51ukgag8r
8v1WNgxg0GhX17Pi4Xwk2zj4WCG89t2UBxheVYmgUXYYD7DnVGaqL4I5vqaLlW0ros44V8PPz82d
kAjaZTtPFJ8vGIkGazzva1lvZ512k3Hh3Dtf82PIshq7iaJluDIIGS5sfsoq0Akys6eqeCRYK9Ig
AvaSgOLYpVK0eiw9VERkH/THB/dTmyyakJicJPD6KMaG5vpbivQ9UoKaw/Ys8cJhlbphtyBMuxEc
WPtz/6MPIbcZUdC938j1othii6UPaH17aWWXS/cPIiVTBtin6O2gNzQJJGKKr/4XtJK+y2DUZ0No
ERC7NmaQ+xGdNOF7R6YRdfNcQT7TP8EM+/sBOxuEdiIdQffbaKNpCdc4vAA63O4QsurjQWci1tbd
BdoT0BsLOOchbiH5/4vRuWK0H6ZS57ovV6UlGqYGuBs84dNdvGw5sHan4dySGYYGZo3xcWw/zbYv
VCJmMAY2FtEaaW4j5rZdEKzdBOk2DbI/uGufyc22QEAeQe1cO4TZW37St1cfMvKHzdFlfrX4lSIE
w7wVL0Ai8sBo6x+EoEJqx/Rtj52sMRBc6EBQeuiPZSpfvPZmFth96tkP+2djn07Rm/AQZNkqWe7H
IN5veszIuMD3vuuj3CfrXYBQLdWYRtkJ1kuIYunMCFYA0HW30tJqK+G+NxtG9tJ9qjkvMvJjOKmh
duODm5j7U97myfRCP5lSDlgbhrhbwxLC3hDCCSLeBJG9pxLqR2kZjdjBHoVkHCl7gW8rtT9W/IRD
rpvHnhTGi1HlRmFHu/UHcJbV6wmXyYFYz9ADvNSW6hH+eHO+SvJd5q3het1q+HgStNFlBlpqQ90G
eHgUtx/P2qhjvcgwYMl5oD5aIPlE9h0JFTfNIaN9vn5DU0wRNxOYWev/BzSYFcNVcYQwljiee+MH
m1zPL6LXO+ek6p8cqVjhUYvdQNoQ7GCopeJVDftzUaNO4mLVgwyNwqAk0bekAWoJn/SwXToITiXm
cH3XYqmmM+gkzxjT7zD+J8zL1xm80Z9AAqd+UuaB6mrIQ7gE87UghVgdHWhIJ+oGC5xOTAgb2vwR
r5k7DFQgQCx5S7MZUbbkFifPQktrnTFMQHdB6G2avMhypO7svVKdfnjX4iT5m39UhMCf6qmxA6at
9O/MTjjqyk0U5UxiqFlBpgpa1KDv2v6mv2BxF7OX+z/xDW6Y/6Gjt5VGg06d3Kr5mBEujOASKojq
RKEXvDQ0eVVKMAzd3vNb29J6wUnCGGvIMB6IQ2zZz0pxar379hLoX5m9DnrvomoPuqJUZ/dO5CTp
A4UiuBXuU/Ft/iasjfGIq+29JAWw2if4TxrQ566Vql6h/dlIIrOFyQH7i1k9xvJ10ZWnZTR07Ml5
0AO2bEqzSV38uaSiWndaO/wapqvpqz8kxFpe3NlRU22bR5XLWNmFC3MELqIzaSNjm8nzwDQVBTeR
W+dYRtxziQ4I1OSu9jLshn+WDdatECeIdV39BR5cPdjC4gTOXsaXnrMMLRiFvN6H6A/tXsoUJ2+E
vgMYUV7GbBargO8Pm5CylNwLwlIQOTPXRXIf+HHWBmHdYv/zA8DHIqCUDh/1P5KgXDOaJ7yJ+9zD
H1QyVgOcfI+2THt8RqQiChGHkYvvQaP0Im1hiHov2auEYdJEX/TIijkn1ct4g5x+QzDKSckl1vym
V/LrZ5suAPTZmQ5631StqDL2mbG57aT9Fkmgq7sjCYWJ1Gnuk6VM9uJNyrDpuT0NO3/eGDxGFBIU
3G2C5vDZ4EOwBrUjuSXuCYqDp1v8ZdYCFmbZD9u6JiDqo0p2ymLjYSuh0sZiuuVnK7uXmML+6TmM
Rd1GrGBDda6vPGPCnV/rxCb8lsjZT+bOITRA9yt012Ue3qYjVBmDKhT0//StFRLnWSXicr1gKETQ
/6jpz7CLYq4E22+E48ZVueV8cwpNWeORFRgb71k+DD1k0qTRQdMxYIHlfxnZZxrYDqc2ioysC9+L
8yK7b8Ju64JfiPEho48SxrI1q8BoJ7829cICELi+ld39DUbmse2mBN5hCjVdfnb+THmJFkhqRiRy
IA9ozRzlRvImwUKursMDZAnAVay5yYx+GQ4sBwHJIp0vwMsEX3x7VotphQ9Wx7Us3Dw/S6kLP1GC
6jNJfiRdQUM3WsZwe48QPxONWd/1g0vfEZ56353XzwDjy8TQggjp/RO0mQyKQp69wvDpZnMtwVeC
9GY2iwHo66fmcZ291zEMvfTjBn8jo7SQeI8NUZos33gtZPjqOHZ7lpkk6gDSepoA9iojxTrjLyKn
J6h/w0eTgCf9X+dTSDsgwrg1/pMjv0Bx/ucbwrMRP0IrodqfKD/GPN2NRJSd0raex6rIgu4iz3IE
tl0uEEinGA2w9+NU1Hycbvn7MXiG2WwKCBVxBOGI+z/CFo7COMNouBuTRO0bpd7SxCX5zhoLEYPT
m848RvN0SYPcp6JcQBcYvhfKmE97GYWsrZFOZ0w7LhDp/ZEvpGGwN2yMNZf0Ecjj2+YgfqI5z/k3
296kWb5kO4WlDLptEiSuatkDFEb5Fz2Hsq8s2lUGyfUhSTaQebrYTg6rLdZTpyZvs9ormu3vbLgU
g+3v3daZkccoy6Rr37Fj2GsUXs+9kaPKDFu7xbgl5Dp3t+ldyaxIALlzsUamtT7W2fhTXEeWb2ss
mM29fF/xtWe6GLnO4+wl93JGpvlcCLRTIjlgOzZhpfOFWpvqiv7dOMvIW8NheHiRbLCvzZ8Mx8YV
7kP2HTNxXjmbZguJM7xqsV1uMmU44hSdVQuLXcd0FXmr7wV6g+stTPz3q4ugPQQxuYtCUiMfsVx8
7hX1x0neCNfAGFYPXXxO8vjil1Xlg3KVn4IF8H2Mghr0lhE0WD54N/Zo9Ybc6WeubKVCz8kraFg2
ib9sWd/jSqbPBHOZSQN30RaKO0YKPdF1G5/cyU3KjehuRLtYr0PpDT4lATwrnSYrA5ZKqoFCFd5O
PBgcGYMTebVBg0b9bMS464KPzDT6eHZpL0KNRBmfm5joiPTVN1N+DuH55g47p9zVGEpAGuLxFB2G
qEYof4loAFfqO/Wa/fr8yKuxMlKmilAKT/iB58gO9kXdAnBLsr+SYRtIAk3wBm1q3FsivNXtBiir
ogCBr5+L4mDX3F6tpeDe7w==
`protect end_protected
