--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
GUrC1l/a+PmqMtsNSytI2ohfSWuHL6GfEj8cO3yktQd6GQuWtu4hU8jyHbtMKnpQLIyfzWd8N3Je
yJh2DPkJrK0DZxQRxBiKlDCu1tWcO5NSp9yNkqqx6K0UP2YgcULuCf4rnDXK26VfkcW+WR8q3Ks4
70nGOk8cFtABcr+VOQXkc2/Ldkwf+o8FbWFAwz4VBwZ3953wJtVdh+o7xLXmER9dyZ1WJzjwUYvh
alhJVOykSyEQ+lfpkQI0tyI6j7570nzHhjfCDdttWE3vUHT9Iupv/o1MxDnwYP9ePTpk5u+Lkfxc
66Oop+zkBzin+Y9QsT59ZNzzdCLPCt+qV5ppFA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="azkouSewRgx1yxBDabAnZKK+GrGULjGcqDgEqHbljCE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
GAhrmmMzH6QOwaTItS2Yy+Fe7wEcfmD1nKyx7usyqo6lCyxqvanEyxS5VypAgPz2gcnX9E5euAdG
kRGlnP00JCg07C6rNpuQHMYSzgZMVVLnfmcZEAKcptd9RsiBFM2yHmMQhlLDiMJYeaWpW8M2o6ET
mKNTk0TK2dJvVnn+SyMd6eGpy1Pqw647JfARP6YC12FnIbswt2B3ANFq//po5tlZSDmdQSvzp1OO
W8YU6JWQsQty+CeLeuWHvhGedCi8gkLFOqFNALdUk9SyCg8SfVSACBoSSiR/ssnfTwlwRxZtNaqH
FQ3MEsiB6F/WC4ZGB5W895sMf4SUogYCrUqTGg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="wv2ZlmzOUs0v+VRo7ZBxNHbchRNIGHLjRETa/b7SVZI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4208)
`protect data_block
+PfriXD5woC+SXBWAB5VAhLDRc51yQgrawW/n8re4K8kNBrMq+SLXcbEV6rvHgjYGMN/CY+2u9Mt
DUlpQ1RLZBUNoK8MdDYi5e7ZZ1gyALLr/uTnzjWZE8j5pCfKC9oMte9Dnym/40NhoSmulYOFYPsF
5HMJ4o2+Sg73/DJ+DXy4HXsDc/ssRi7QQHynMJe/EBZoVVVG4HLIoRcssAvECKtEs5y6UvP6Y9oA
GenxygyWz0QF/5ySiUgSACjUQQYW/uGk7xLkB2l1ymzxlCNwKFIvucMI4oGeVVCR8cSNg2X0dynI
qZqfkP9T1d8K/JQLgoQfcQMretuCtjPmWcDJIysZ1g5XA4rzp7Cf8B9NxaiNGrUsi8uZ+8FGrLHh
+vUfWp3Uz0Ur23g3T5UHusota3Ls4+pAgfkjFEx1DxBOzUl+unZOyItaNXIgvvFOwHnyXepk2tKa
gPh9DsJDF45IQ+IoRHsVD0j+Se0tQZSE5+sYQN7pQWFPLscEMopeT4wpL/+4HGcc3VLnNggj8/+g
AD80Tnd3V2Pquh2JN1DCFWNdtYzHTbgXr6nzljIB1xAXuNFUe/u2pdTE0pGKrcO1BQPTCCw+CyBT
OCcEBjNWLaIzFPKHlCJ1GuLQYekRcpM7EfpV8dj4+MntN2XPOiLBErcCJM16IMPwgjbah74Ca0az
sTjo3QYzzivfU9khObnHUzhKUgpRuyscF91/GBYu3qnE4iJIzyp9cV+ZkaRIpj6hxsoo9dYs1Xz5
lanc4KZE6YBgAjKkVHY+MCaEaJmTNYkoq7mz7Ofntd3l8UPEZl5sHTW3JT+GFGEPVFbIeMaOBiaQ
CyqXz3jUIokH0CFzzQxncQzsBTo6PAHtLOsw4eGW0JvEM0nl7wAiI4mdFOAcMWKCvdqFPXMOO5e+
J2vpRvKd3hBrVRQv6nlOtd5EzhEF267NMzKreC6Keqhrk4mHjj82UdBhm79xttGN8KG59lAykHI4
RH3pAIgs9gzZwZf2wcJ5G4Jva9zI296iGHPNRFAMUuTxfuClI/RuR7ZRv85q9mA6U292verGn7z5
NKAvaDDb3n/pQTaLwJ5jFzAOU5rcyc/57ud5Xh1pWIRsG3CbTt7AmAWLnSRz3jiyhzHc5r2vObR5
hxJkQw+sRWy6PfeXyR0JyRiKvSGMPtknaXI3mFm0eI/r1Ax1vPO28av9SwQyOhXM31wrTOp7w2ET
P09t5sd/XCtg+NiYb76D3Rn6RC2RXrRNTSCUO2IMydIiM+O/3aeARm6M+Z8UABysdkWdYsUb9u4m
Rdh9WS8DPOJ6R2bEQvTGx5OtZIrDcmR9iPbkJs+N/llvBfqtfn8jkXKoXMlGMX+2ViXwtJyUnb82
VdaK43qq4/IPjGQZkxvJiDA1uexC4MkeuLnJCGcneYMraDt8lQR6qUUHaQSn1foJv5i5tZZsDFDI
vICVNi0UrVaf4v5tMgDhCafilEKgrlIrlpwzF/jKisqwu1MOsvwqLvxzIbGsyxe5wCL0okphbgfP
3IjZ+xD05Def2sg/K76+Ro7omRt5kTBnLX4ApFwIuz8tBr5PeoVjnvQYU3kTl8HMyCgQgP4MhYuh
EzfWmrSoZJLyPYacQhNtfO/8W7eq46EB+U26Y7/UpLXlm+DsoYsh8jnWEdyS4iy/Frw1uWmPJAy4
W97hFQsDwEl/jmLirkNPmoGUQi0417D3fg2oDnmPnNZGzML73mBwX5eXqYRl+K/QqZnKRpBjromm
bJdK+IUNgOUhwiggVtAPdcWTkZ0X5Z/Nb3mu1ogB/xroJl4yoaSPkFla7VucxM+d6yu2uj01s2wP
SXYhjMfvEZZXTJg+gZdbyCg8V75h8QbFoK4K2cbaxAkf9soArJD77GZq0pUZ5QA3HL0AEebwIEzb
VOArYf5Dmnag53Ww5Z2c8YO/BKtlzIya0+J6PqVWS9At5vHpZa4+eb4v8Ap6jMz2hk+r/LJm9rXu
rkOUGcIox5fifBAXOL6BqIGTfGKMI69v2KMy3z91CHITY3dXuDs8nDP4cSTE/hSZ2hS4ur6Uu1ZN
I7AeO2vgakEk1yxXxPSLzUj51Xt3OYoTI11IfA4qrhx01lyPJqF8XbR0mle8V7ao2rjJiHC2a9IR
aqTKMQ9wl3zb8ZIG4CSi+5alC3vsZ8vS7BvCleiy0CKCWaR3l1conC/z0gpGqKxfljwnGTQb3f8O
zQ+owHjZKVv/hxD8WEWJ2XeQPbUR7MsyDd3Nhzb4jJlYgrdVxrxv27cucSzG55x7F9Ypod8s2Lq6
K+Whd5mkoivv0FdrajnFkOdFr4lPPeiwf3mKFM5DTwZQo4Cg+nwFOvU2+u0RR8qNOISZ0PjdiYt3
riVFGSJLTOl0X0iEuPJwqXJD5rPSf1ULdHV0Vud5LUjrbPOmiCA2RoqxVNtuDYYK2UXPD5olJb7K
dQWt4PCGn1qpfoeuTwUsp/Un3F4XZcC7UUJsGV60I3SykYv5ah6JB4ibUTVqSVdFx0jGAugW6JyO
HLDXCk2nuUO3qOagG0MsLBioOiH1/qVhYHvmttdpa2KmBhUX3iPi82ETieeQQcP+EXcE4y3ln9Ap
xUVFBR8V9e3Ora7o6VUaItPRtEPIgV61h6zbP079s9zZI/NfRpRK7zFjk5Qa2mlNBOS+o4/B2322
TIkVXm3JFQUaUisFgGNNSOoBsaU1tvjDCFLR9xSLtd/kP8WfVPEDggbC3hdWk3RYXiJ13qQtr3ZZ
yUelynb6pgzPiUbktbwoUjuKBopz9NdGrBlvqJBI2fwGvvtZY/kBZfNQeY5T1rkVLDgkq48hdAZ9
vVJ9gsw9z10ldnWOJptvSXj6qaCtbvAAqYxBrwEVpOOI3ebbPUItYGtW4oxfQArHDluMKUIZOYd5
IGQVQNPiGcAh8CdrCg9PTKi+hhtGWj/R4bZCMNOapqgQ6Ud8SH7CayiGoyo6WKiFywgmPmglK1aG
qRk5nsMTytnxw4nzdYsB140hd/xjANUulApccQ86IbnZKM9ZdrstQLE2QxWFpwZioawfVp7EASlP
e+9Chp5+DuydbAp8u3A0Li8LJitKXdtzs6cElZA+N0V4jXGgC1Ds8SeL35oEQSwsXHCUX2bPDZFd
USRf4qP6BM6l2sofQH3UP6/6o6c/9jsUIsJXS0HAe2crSeHXqW1HOjYB+DZkko/QYkfL0CANNRcY
aNVfcPqTuloZp4IIftH7G3pnIK5kJDjAqvMJTxPnSndcyZsbqZf7VavAJcKz5W0i/Al+zpPfZODK
3UhN2T0/g/xx2W+jt6MKzysLYiW7kd8VXY0xkyLi9KJuWbZ0Ujh0cZ2JCh9zhMlskwoEpdxJtzTo
/ABxUExPECvepMeGa8Hv13CSvoqON552zaxNxeSTR4+7aY9gp4iZPxnuFb8ueAHzNL5oxjgx/Dk/
a7SLP0TcD8OK00So3/rV3/sTx+p581EWQoXa50cYgKTO4zlBavsdCHY+mI6/c6lU1iwZQMpt7yrU
e+ppW888rNVViFr6Cwe0LQ0Bwm7HPJHd/oLl5xiDwhOhhSDHh+OJmFJ1MiGZ0ZKDjcyIyBIzr8Bb
D1OK54Evq0UjNDw6wPa/ermDNo3j4gchcOzsvBAodvk3dPUGWTccu1E3jDtSsBOzkOx2MuLSadac
ansfFCRs4EZNlkpQP0YSi8SDiFKpIgf66+tw3gRcGvVddCUhDWB1pPM0TkdEFlPUlRn2Ose5j4T2
jsrdpLH5RD+0MbzXaFwZXOD/viqGgmkCSKfA6sAnta/Los076lEvE4H13sbyn4hJtaKIapiB+iVo
HCsrPeMmQYqCpd8Y8beCO9nwVWpDrQ+lU+pwgwF9nzp0RNslo7GX55/qAevBDWMDctdpxGRghpq8
63N04ZZuuMvTxK5p98xTSZc4F00szenWpCKRzzutIYmoCCx19Sc73Y2a+X+dF8iWNM2Gl7A7RQ4I
q5yHd6mEzqb6ria8Jc5bihna5MUOeLXu48Rvt+dA/l7rKm26BSEI/lr5L0tsT0CZ73HNiQe2b8aO
qhApHLHy06gQKPK5KiibKuHunlYexcYz0odzvBpUOmfPYayOd4WClJCgH5lf5Y9igOLu4NWC6BaJ
kVCiDykqh+DVStZRy0GVRiwwW0o7E6ANuesu4OpY3K6WOjlZcQLMq+j3+oXwM3P0LwNE375F72KD
M5DJ6w4mIa5CNeqpcmR5KX+M03e7lMSRhIAWHjqWea2N6wM6D0MxYkEFmoujAMk4KSHYGzHxxckU
/CnlfxiHBpDucq10vipoeqS6PxqlZJwjdgXGPnJke6yttxknG6KGwtb96hD68NA6gXCw93gJn0NC
XKeRMYXuAIDye5cr5QkHb4QVx7V3xymIMdxfYJg3R6cpwp5vwbRmXS+nZD3a0lfP0ZgSlZC8e68S
hJbWgFB5HceHyexMWckweO92dS8D9hZBaOUWF0kiqO9AQKvJ2H9u/gPefgTkcCbp3kHES8Io1vW7
Fs1lNm2g8lwIn3Tqn1XnhJzJdmC2rmiEtUhHDQhMXjN72eG2RCU/nosdxBqdPVJ1isaSWMovjRYV
Yb7ZXj9F/+Ce4IFj3hBoYIHyvApbcNxvuT4+7oevB/7xMU9eEeGtho99o9lK0yTVzJI+XOOHgBkZ
n1CTdLPtzDHd26jxZ6iiCzV6lSnlEHFQak64fDfpmk3mpVwkFmNiyyFLPZumtdtZmCiKwCgZgkvK
adHRmHL9/s37dDGl22WkS4hl2Ckql0xJ5qu+S00DUsvHd6NSx37ueQaVyVgQ5nktf+yjfCBPffjt
IoQC0JGXo6Yj7GWPvNENLgQl86fI4lNBN8ZDhnIjkX498WvCE/RUr0iSSiqM7p3HPrlsOyC3u9bO
lhrcTcesFhEB4r8u6QqFv0dHv6QAo+7ToLx02ybLrAuD0JvKC07oSHyLvHtpcqMqLR6ZGxp3YOwL
1I9w/09z/fL0RqFqzzFwPUkoQKey60CKYMFCF3BFKA7h4kuvkPob6ssR3Duoq2C/kvMoVDCImN8v
pHnmLd+j5WYyGyP7c1p8BaBdDRDy4IcsRPWBfcBktGQGJTdkikBy078M5G/0ucvfS/UoXaEhzPEa
RqVZN6g9u8+xEpqtWpMn/UdsPgKH4AEURHmCOa6/Rn654kXRGhThw7DvT+omRVIPHNV4ec3jMkOm
D7n5K0jU7eK3N5Bedbmfd7iz5WOsHuCT0oWJs6Q53p4LVrbWhU+1Us1FO9sqE9RkjVNbEuKyzLq2
dpSIOk+NdJX0fa+oMwHWO0jXXMsfXJoczAX7XSG6i6Ze6pVUgFlHG04JtEOTzlvVvxXXcLAc437i
4vfs6vSFErjMc5kjJOskxqIFodbirUcMQrq9fyOhRKcekLbEdx6vO9jPIgnOl15jIO1zipzAGseV
BMX6xmzvJ0ldWoOSM1KML1yr1Kg/KjkvYi0FMlo7miAQ5iRuU46QwKQnvxnPoOi2huGHZhNgEdgx
cWvFX+vJ/fsDNnxl7RKtZfL9tPPnp1RVy/8vOR6+vLdwD1fXk5RtaGtritAj+BtlEFCaaYQoi/Cc
VYhYqWCHNAC1ZrmcN3i18VxUzl4PyELNKMKCmpsiW5YoebQkF/u8YDcIFcoGflE=
`protect end_protected
