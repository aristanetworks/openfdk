--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
UY9DKXmL/BZfYANPt/EDxDJ6q7Bv5yJral8mpMgVNpa3//CZhwQkGnrjeU/cGP2HkhOYHOAfHEsZ
03TzE1BJc8kpSsgEVV35v5ZJTNMSoDD4BvOePIQyFg9XrW3j95LT1UDZkP/4ReeJqvy/7Pj5xG+k
ZZGpomKdMnSa4n73gUXS9L/4eS1xKOkU7DJxPxgflK5w9z083sNH7hnTJIWmSuOqS4OUp/v5kj6X
wesXc8KjRb8T8+oNqXhdTRyHO2cLS+zK5u1/3MM1lCwHT/DGPny0lE7tRpJAc50Dp8A8tAJeUOWF
8SkWNsXL1UOKC66jK/LpVMMQj1gDO3YgQoNQxw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="ED6ol6HdPoxmnge0eA1s+Wr89BsP/dD8GAAYJ4G8zrE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
oafaE/Or6LT7kNJmAEby70N189t9WFVjlXzMdFiWI/RstA7xLz6/sfSF8O3FUGtFMkr2otOQ5Q1v
iO1/DlEbrtwIPOmHaGB12YdDaDO1cIVaEP/CqyyxeWIiUtaRHL01KhCdMzH2Q5HdE0ozIVmodgm6
OHp1t5qaQB3gjw87IPgVLWYPh3ThwHH5DtvD6BJiH8edFSHX8GDr2tkfPoCR9JTSIbZL9VGDCTcf
VP8kA2bGdA4MuUZsM8SaTOubugBwPcNcsUPkgMvxo1D3u/Gt9n4j8qMXbBpciS9s3fJEik+xE809
9EfPmdw862gcS9JVEUGNlR5K5d8Y7Oto3NI50Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="BGo9H9bKepWl0I+o4lpworqQ0sYttVntecxFfCtnn2U="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2080)
`protect data_block
MbnrXEdseR2Tz2cMWjW3bzulaMQSwduTz+PtpZpzmWtvow2cd54ZkF93xaqjAG0tikzk+T1ac8ck
JyTpv404fVQyciV4ExqMcy5FmXNUaWwkoQgIbeCkATI0VMrjzxyEJLxuGPcRlSr9zImq37K6D72S
ECMo/5TU+8hHSrupe/Oh055mv8F7RgIRtidk0hpvT7bEoLYL+eCVU8C180FclnoThiP/e1OxagdM
wPSteIHU4Vfq8pUdzUqAJGWp2/UfSrYPaYOAOyHAxj7fl8w9PU3oQrc1g+pmWZ58x6QnWS7SpH11
ezkIn10he+btmXne0me/wf6Vz69DrXuKznCyuykmhfQTVpCIagze9QAla8Bcpx/gkdXrqELfm+83
tjVT11f41AmEmvjIrGgjj0J1LoFW+FvMbc0lgl673XpkMMWBS1Kc1NYaejTF5WsmVOF8Cf7B66A5
G4Tm3d1U3HX4rVg82mhL7ANVXZiW5hgNxgZCuwNFA1pINH0nNZ8e4cTlL2uxbci2KXAfpVBWzyx1
KtqQ9309rym7ybxXYvqpLWzmWn3KRz2EMA6WQcftl4JdjyRgbvVjVHAuG3YWvIIOjXNGCH0iVFNc
e2KG+ED+qyc36/74p76E0WpjmUF/qWPf+Cv7fAUk7xNKEtoKj0H6kMrifr2gr08lXi+ylHrTpbDX
/CspluvjkHnPtwUUbjispsEfflmqaTxFvlOUlktrsp2/fuUYAqzZBi3xti2O8NIPCvT7HFS2k2Uc
EEsHv/PbeDoFJN2+PlvKL1Npum8DKFDIn/nO1ZnEPQjig6CheweUWHMrVj6y7o2HCzk6+W+8HHow
ivPB9c7UxbbsMGPYa5ifFhD1bFZjaELMrrWgae9OjvdtOfpVgUIM3rM283ETkAqtqJz0x/1A2dFJ
hxgINQaU0gUze+sgrbISsv5lDXg0g1cI/MMRgRMwb/aAVWn8kiKVopHVB70CrgD6IgJw2jCl+H1+
0qefh6prGpm1lZ9NZJAVGyNkrodzGu2NnIagRRu55C2aX0arpYypITVXIFHfwUOUtJzliU+35iO2
yFwP7frnW8ksJnDOENAQU3CCXymCns6r9xbi092QmTKnOlpAckPeQgaRuT2u3zOmdeyZ+F3oNFlA
OP6ZHqLKyu6AsPqjRPdSHwEWS3+enUw3pOeFm+XpRJHPuoi9s1TNqpjsDCK6XAHGJbXwy7FJFT66
mCqsG384y4doWGM5sZOt4l9nQDBMoZN6kWGfsHbcS0JCL+Gkl5KCb0GNwNF3mACFt5w+uUY/+LoS
v5xiRuTgZOZtCot0KRuhlrXOTKJGYsK59TqZcQvIhvwC7XmG8WOXU4n1zliZBH1ctzQiCbQjT5HI
ifeDkqlVNxaacA/pmJz638MGBCPcs0L80QAo/+pbx7Vu3JhIE31rr2O3Bls7csLQS2MC7Zrkwuyt
eoKrN1LZ3/sJ0csb7YVB0fJ9tNMayDhAcrV1h66QTxWXM1zBhYYxcTUr6De92PCL+PatVSaTFOGa
Ecqc2DjVbKBjQbYVrETM9lpEFhNEfKTRkUKeT5zuLmyG1NPU5hzUfHw/NhlMBngCkt1oXCTUXQJk
XhX5c8YSFiSoBez0SYY5XyIGj+YRrP26hKXrAG6py2a/pTQnHfThs8xdu5QWVxddmYEq5SqkUTxo
/Zg6e0Dl0WS6gf98vJUup5FC+JxoXj6fLpHCM6JLcRJhrxdg47TjHiH/QaeAtAmuGJ/sN3HgtCAp
WGp1A4mq+PlIgWtelxvPuOHrs1Pgg34jo5MtfcYq3ff67ZQ0MiTqMQM0jxICb+4jWYMMEnDIJL8Z
iVd2qizFnaagT6NMBd9vfl2+corFNXdN4SAVCAj4zZcD9W84avWqGSmDM+pulo2oymi92BX3egBQ
1RWrrOM40NCP8NwJkAbnpwfE3pVIG37MMFDKHz+aBIgLAX7v0Miv0/15Q/G71diUvNUXJv5pJ326
HeMr4uCVh2/6H/AwTTjnI9RFzEsHxFYSZJvfgexDZSWXAv/hG4DSYwUYRAL8UkjEpH0uQkzo4rdI
uAyg8mXB3ufsMGEP1HClw2v+UxdwSFBxxspx37CPqhfp0BXn6EEEDPSmWd3ued1qrfHr+sW9urrx
mkcpsjzrBvPaEcy/xX99p12dcl+WWgHmduntRY4lFHtbtEjxEGpO0YU5iczpTUj5QGt9C0w0b+Na
op1I5otpkSLmRWg1IVOr93Y9AeZsBxc7qAdj9jdvRUKgTAUkz8Kmog7Lao4cwkx8drgs7judq1p3
dK7ZeO4WxH6mATCjV8ri9dsMKnSbFZriYaS6BMC+X2XR5g362hzoRaCZxXVndH9Fi0ScSatTnwaa
JWcRUbmJhPSNweSGFo3vfq70x9lBhc3xDjosTt/5gtg6Kf3nF5MXY6dhcjNsiLHTDOoz1/wFVJ0T
s99oYpKRI3Lyj/4PJWEKfRXCnCy8evEty7xFcD1nEfNVIwNTyAwRCz5jBfCqSuZDaruoNG1AUnDq
rYgLxzV+4g2B4P9ymjxwzPZ89BbtMwwGPaVZDmmGk8kgRVoYKbcFMMjIPSMokA+YzL0pBDxzP9t2
gBFtT7v1kTplJdfCZ+MbWtQuoWiraMhrliyJgn0uOadTc546nwXQ84HLsoLGnb7JJl7JlzqFGQna
8ctGoPwBPVnKyPBfUgTjrHhAFXzeoNlBGCaT0XCFcWWsG7FxvuXRpFI2HnSNnnZCp1Do0z1AY5OS
c9I8RqfDqqKjqhVgxvZaGxhv9X2f6TNQgiZY8Q==
`protect end_protected
