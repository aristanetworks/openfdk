--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
UdL5FldFe/wEIua9QEquYeQnCoKbWnv23MFVvpJSAKuXU1DDKYPgVpFwkHNiZp2NxA051lMy3JW2
/iP7QKC+K0+xNALx2jyQ8hWHhmylep7LqK+xhMAQKMIJtXiVDdb7w1sIg1tXaJ+q9sj2YInHE5uE
m68yHl59iqqPG03Smbao+4ltixDdEGAH7zpc29ch/8VT/1vTeIwY87zVuCilU/eMlHfHVR3aO9a/
UfFi725qzAAz6M6hjfspSgzFdO/0pe2iLcf6MZ94YmUOIQ5kZCTUGWYGwJbIBpDQGuosFNnCMzz+
piFa9Q2CQFyeNXY5QcHQps+DJ0uy6EMNtXGiCw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="/78uUBueRT/3P8cEnH4hqaAplsm+vkz2387W8veJNkg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
bZmnltjkbAFoWMPG6VoQ5MCe3mAmrQ1+IO1OWwpnM6x73j2cCJqUEAon7oDpSEcwwVXj5JFEn4To
7dq/B7xAfAKKgFAvNp5m8fxvHW1H1B7DZTMK0iltyH3cuXk+q63RcLg9Z2gD4YiYj58g8jRyKsGt
EvcxLtKt90JICX30UKuiFFts5hWsJB1DdZsB0iY4RRyESH7YwI1OUkUXxDG2M/tYVkTMpC83//k0
jtQQquZI4XQL7vwpsG8SPxpq48h1ae1t+tBvFYNU3VczaVwp+xQ/OJLt5vg/e7PVtnx5moKW95DU
J/BvPyYDn32BWZ1Zp0ahQu24qSZHiLrRxV6bNA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="y8F0v680Mkd/QN8jVs1YujaS6pnPS30bbCLSU9sSGp4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22288)
`protect data_block
2/d0AlWvuQ88QwhUz3x/nP4GlEebxM5S1y0reuBReZ1Qjx7zucY1OkywG1W3+e3OebBi5kJZOSMs
3n3quiWqkvQubyXOi0SsYyRj9NwDmewzFOCQ15GVsc1pqes5pAoyXtvxK8UrsY4KHb6eusbi2Qda
ccdnK1kzea/ygmjuDkTTr/mBfn18AlQFUFAfidnAYM08dnqwVD//K9BfAidd2vdZM7Ye6ADQfuvE
m+aoysIdWALN+EA4YCSe3Ywk2ABnuEMQEyoQw5tJiwWCuF29CLsGYLjDmKt8Fxdt0nCZV7/wu17g
BBarwtqPZYchCd1dXQZEmFJrbRNKzqJNdWn3OCARTlt0NExX3JuNs+6mHos4AsXzsG3zO8iLpm8Y
5KI4IUKHlO9t7KwnV3ZzUyiu42p0yls9ZjKFbV0O9Nx3lZ/1Vedf+XBCftfYYJKTcxam/MFCnqGl
fWLnqlgaJYgqtCNk0VPZ1KnRBM0c9dBPcMlGHy7yB9wo+G+yUGUdDLQ1w+wntALDfFFSo3iO4j3Y
ucc/8wtStrcUBDS3s4Aph0CgrlGa8XfVICJcUgO/6d2Vdk8MoQKmU4ZYTyPOgkYsDB9lBTlATwFH
dRQUkJPVfXTIM/SY52pdINY8vpgaZOgLGQuq6d0LiOY5MYBNqf9e2W7RNIPM98Unte5b4JcaK852
a3rr+H/UzE/uQW+EfVtK77pJ62oCYCC9LaNhLUOSxih7wIjUIoMVipBIUGdzUf++7Oo6KaixqtKg
3+wOwZEMTWucjnRnGj7WtzY52opRHgvlGUFhlgzErlMMBxine5sTRaruVOlr2+vSWCeRkseUIpYn
HfuIA/eZhI2pAtpx+5jtGnJ5O3UIiFQf5AltlqJwX1NSsKHuO70MekqMV7CHXSj9989ZeVs5/KUp
xDGPkqB+mw2cmj/KA8KgM48RWFjLqkCpMZhFth0mvFPdvfLAfg3KlC6H/2FB8HC0A7jkYn4B07lE
7Vr9YQ9n1iHjwdOuEJSPzic1EM/TRqI6tqqGF33sJ+UMdxljj1cacsWLmK6l4SYz1+k7vzoyCUzP
0tWM92eYfyxJKNM8e/U/V817T1CzejewBp/DeszAMPpq+ca5v5OqdUDTeKoFsgRl7KL0BBk8vdU9
LS5q923/ZHrABzl17vVv3wJxlwrwzXp5Au1U3AnULTU0dMH0AV+XUWrOYxOVilepSpg1aLQm9DmA
c8nuX5u6VF9/vs9wAv9rREw16iSCWHrjyle3ydwkXikoYkprGuOUM5NlYcE4SNttJFPZYqXB42We
t9J2wqX41Sb1QGav13zPeaOCqAE7S3NHdibxhda2Nb4SUvu+v1ZH6QWCjfuRgdLz+VU1Dl2+XEac
1H8Mn+d1xWal+37NsTepUw3/0BXI0/HAOclhaKGswFO9HAXEN3aO/Je1/t/y8AwAwvK5zsNwlbVa
1ashyzkwv92qB4SFoo9QKw2ZwOr5zjv+P1gHjbxSYMP/rv3qorAyBw6m9kb3P8P4NKQWjzm3PTCx
ngla3ZIP4zfhU65JbY5q8ndc9Optl7bqxDEIQrgtXB03CCsmkzwPnUa/xe/nkPT1Lfh9+dH0hw/y
uDEJl+r6k03rdyNkICvNpZebj/8N4LDZ9uJv7/GW+Dk8LH2b8R69plwLLqXzhzHwu4DbKYk3VFzD
h80T9AcRki2Q6vcKieTgcOcYQF7TVA3Y0OFAVcwOyK32jSNm5oWevKT2lk3Ylv+KB4KhxdwoJlvU
tKvDyjYwsqHJdTESZLV2ftG0IiIkVKiyyn9VkaSzJMKNJNmvlXW57A4bnNK115a5+bHN2ZBDVTDN
SV6sN9cqacTjGQeUBULep9NIxFRzBoUGg4YIz/Fh7ClMPgidePN2x+G/GUiY1KBXaByP9Oa9I6LY
SJfjg8S7PXK/lwCnBBoW3+xx2gi+3Bx11DnSwyJ2UCRCP/NmVAYPDt3nKYXCXko0Si6Hi+bQh9VF
l1bNXKtrsSIoYyK1L01tNczhoSuVSnucqEK5RR0DnWUE3DtNeldAuQnTLNa2UHy432OghMMiNmL6
VzabS19tqykkg4qcUE6+lagllxoI353YeBZWzOVD2D95pqwEljNjwBuhgHmkSoSFyzq9gruvV8+p
hA9aVw5+GK15BHBLhg9zf8nYfegn0DG1UYWPSwmClvgXI08RzZXS20Xd461M8ssp9BMaSV4pb4Ae
wH2iATrEI0o8PDqM7SHy8en18Jk3ewhbkOwYv8lbtSkk3+39wapaTTeepcZ6FjhDaB9nWguOXVR1
wBkyT/KlmKjwMZR++HkM2+t5pmLkvl6CCor6lnCJtkG7MLmCJCc+N12Q/Hg+qmN5I9fVl8eKazGf
3GYnfJaL+bUEc9jKvgJowtQmSd0qgfOegKQpJt01P7Z8DmFyFjk9Pjfyyv9pdkZfv1RxSA+Aoiru
X34zJAvRvK1ixoAQE5fqYKDiwBmAd/5p02z6cwSEHLqewd+6JxXy6A/5ANcS2q9RgYER27b7bhyR
p34g+w1awFeRyYhGXvKd1bX5M9tQ28v+VoguHg8jtwklycT7AznvVwH8LTnZ/zBILChrUR9PQ2WD
iE7sVVAD2KU4hll1YRVeBbm4iQmValQIjNzkI91/1vsBwaGmIRo5CYO1t/PkXpjj8Lr+tiElwA07
sX7KTygbjHjD1hXFRk3MBGpcOfsKhd2KvkcvuGJTPD06LspyyZWmGehs0kYQe9mF9k9mxxvU0SUT
ztthCmfpg277O3pPzq5fxO6F3DjmRRvUDbWmQIM9mcHI1CeI+N3q0SmkKuIzcMnL/bEqhrBvowVb
/i5ATyKvUDU0Xx0C3uBq5PMbzWJBiHubBuRMRufRYlf8DruepzWKWKUooQsrjdiAoGCiGQPqm12Q
OA2+Xz1j39RgiT2O5u6f6Dzrb0VW/JE6J9UG00mKfkgJxRtyW64WWdfwRIFZjZ6a6L2OIS/JREOr
8ZEsJr5ELVZVxMNB3kqDF1bhQxTdkAlW6MiibZRfUuMT62kLgjqkN9XZgSMFhNpu8nZcbI6a5v3Y
wA1T9aE2ieBblK8W47/pKzJWK7ML/hnn8igOTZjfOeiR3iTBHBgh9BYm7m7tKagP/A1K5brG1/8K
GjD7NQdO59kmTDS8cCpuv9i5jEtv8yYrE4yi/v8J1tlsCZNJsF/xx6HN6fvhU1r5uLVcmaRxR4TY
dWTxkhMyNWh4fgM2SPHUXxAsJCA9M/Xk25A6kzo2UNfpw8t6/PJe/khv4n9yDmcpW9DjAbqCFl4I
H4KUg9ty25fh8YB7CJfo4/ZR+xuJ7XAXXY14v4r4453W5Y8XDZzJQVyJp6XA235Oab2/pugV1bZl
zfwwj+v+ykjg33KmtFxg8om7w1NAWBJKaI08qsBhvA3SPE6Wuq5FNsCPAv6kynMAzYQokejlnWQF
DvgXpDB7cmerJcuZm8k7KiAyzWfgq49JfA5Mihj3TjSyA9i7RSwvjIebrwZy1/TwvoRuUAM3GFRW
Wx5pky/EXl44RAhDysafvA9sq3LT6uzkd9ImRIeYueE8zwL4iayFPqcPtQ/WmUBGIHlkCX3jqKU1
KqbMfJHAn4XJeipQEH863amIo1YhCldxQ+KvYf0A9srgWg1ZkgobdoHpebWSNdtWHGW1m9KACAlr
7pB5UL5G53rFGNTPK7uqNhm02AgEv+cjDr1+DcZAQrisf6sEZnG/nu6INsHIoT4Z+Xfg4yOXLtyA
zguvVcqMgAvHsSuRPSs3vGKiCAb8CsrZzHw60XdOKgKZSN6tQ3Bx7aFgkP/15oiWUu03m0LNlsNI
iX5EZg+Uo9YiSwiTCqQZTpgvANShmc81GlDCDLYi6eqCLhl45keOrUZrQnpYUFG/LbOdEWfqZrax
6OMmM+pt18uOo3r56wsrBcm3bQl5tEfpGmDmUINSSq7Tcvy6OIEsNWxOf94Se29lVa5ZflvZsu1Q
aIAkYOSAZfxspJ19fU1THzPFcUmjW1vi5FnJ/RH/oq0X2CwJ/VnuLChmqhGchgpqcbP8Syac2wzX
PmTIREgX3VBS2qH/cZ5+oIKsWvDwxfpyUKm4O1tIU+Hog5wEQ+KQpZh773THc2XZJcN+E2djFHC5
IlzhXOxB3gaRUwRtEiGboOo6RC4wXbHte83gyt2r/nDvyl/cyt75lRs615GCtYYM202RoEBWRTm0
tbst70k/oejo5mEfZUW517mI/93iM4zLASd1xD2LpykS7j7mE4wEMN6kD1JviV2JictnmPmwhQeO
w6ArGbm8aemfJIP+ImnsJUksErV5eFE7c1oGZwKr2kupvAq8ait9oASXByGs8Pwa6PEmNarU5AuB
41eQXEeddAWepTKnbLcFFcb6xAjJ46PMto013ocui8DtvIDTgMv9VTcydOCv4Cknvlr1lFHntne5
brtAsaMOycryXOcWHs9VdkDUN0U4O0y79DARenFY/NT2zvxgUqcW2JPqqPNcYpU8SgK43pjqDIuu
P/ZgNsQgdgVBB2f0BxGAboqkbi9czGsDfAJVRvgXPm+c12+2mh9ceoNc7JExhbbZywhasN6KyF0A
IpWdMP7BNR955BFJa4t/ADDfqA0B9WwwcrI44ac1Dm2Z887tKryWrfYExdH3rQa5UiOJLZkP/h/6
w8GtPMZHnQs8QY0PoNkA96ye4F9kIf40ATt8ZzMOppGQVE09s8aBJ423bnMFE4u7/T5WkzNv5AAb
9eqQ8NmM3qm+YDRkhuCXTdWt90/nKpRcw/WDuCtDN2NLlmJDcR2ez+9woKX2NGAkTYc7UJlIapQm
4D9u2xlxDS+3ZI1CXc9SYxpFjDeu7lkSx+ZmxOl5WMIxVanJqPkWexUBrZKlRcoDrDIg9eKKV+ZH
qHyzHH+8urECjFAeBcEnySrd0GPa/n9/lGHORxrXgnQnNhp4YMmLXSjTmHkPAEi/MGuZg2ulWqDx
LQhwUjwTAaIUyEazTuYhW6BDH6vhOBcgJSjxn5YfDY+K+a6USiqfG9KVsLS24SjHwFfZkRAo6yJL
6vJMRjdoEWc2BAYtrUxD2/5oeOkGre4x1mnIbpKejsCMGkp6bQRbw2DBXCQDQcaLBzLELEGeBAFK
ZfV6aU5YFH2WA296TdjZ9J+9R9KfIKT0B+YDDpEFlgJek0tfrtt1CnV6FuwujBgXWln/cLLEpVMw
Ohk0HEO2of/3OCEZesIY3RYgngDOo3RngwRIffQPKHPx9i9lY1u4OgYoiqXDK9tnleQNapCX9vuK
ukFJYw6WM9IEAawM+MQXLlevCTuYUkuPAsOprzbSKXuToZBmLW8Dw61Myv9M3vTsCxFtrLMk0ox/
3g+/eEs9dQJsKC8QiecNPRBlYygLznBM46Wm3tdW/DkbxePSW9/IU48ZlltXoxh5mF8IBiHCWOfO
dkaK+zHaUE/U7DgIUvsExU2karaH5IbgbJxXHI2wtS4Dj0mdZ354SqQkfKmT8pVkq+Ny7ggZkvjN
uDe27BqypKO3GFNrsfwMCyEbKaaHogMMFQM4ctlO5ilJePTyMUoVWYG8ddyfhbZ4IwyUmXFvIvk+
tLHprgC58EJS78EjD95+gw6GpmRD7+tKPisfIk+SPdTw+Bcp6lln83prleZgYskx1pANBQ/GfzBS
Fzj4cNhZqVWOrwavIcJRY07XJM0eGHALQVIwnzGcIh3SbW15CwHEe+N/E6n81SSrEa+lMObDJUjU
/jM9ns/hXW1MzSjf01O20pgBvOM6mDMZ2iM+5ioThAvHrv5LbqOeY7Y14y2Qg1IB9/lW7rQbdKuR
6S+GPIO/SeABaZtWEeQORmOcVo7zfvveaa26EQ160hjp1OyvMUdSaTSlb5eozezXVPkWq59Myein
Hdh0kzorewnSnbP/xkAsS+wo381Ifkct7QcV8igH1meyMuZMkRSrWT5X9lHYT4Be/4RTG+TsOFZN
SM/WIaiUow+HRcE2DyIpTTyziMdyJT1hIsjjHUsYCfRh3u0QzKEVjMGIliXUcXeh7dj+9s/XVsgC
tl+KoMNUQd+5cqUG9qStLJ67Ov0n+6fBxcN8vHbgeAixqbZUeRYvGc5Gt/dOzOTFC6RFkdFxqrGD
4HIj6lwbTMebxeXH6U6XOo+dE+SnkPaE8vFRtX3A/Xy6khFqyjzOUW9tVlNye8xro9dSEt4n2Y1i
kgCEan6OGGYyHB8KZk/kTZMOptVaNsOFnuK/0uRI42PGeUE3v4EBLdarEbiu+e5eckB1a4VwDajL
5UWaisJT2t8qhpcbyO9E3KN+1vXWdhX+frh0xlBsif2fqfkMx/qNUkCkDJbqzArezBpOZMtuO/FU
u/Q1odArB9OP+WJo/zIGcAjk2k5FY+jmQ2unR3l1MAET0+GSmHl5eWo8i2jh2eLwZPGbKEnIwVvJ
yoRSJN9p+WpTHXirgaKTyITaUQdUjBGJIlLjyWlLsQI4Vh03ca1RFTUAIZKj0HlOb70bt7bnV4qi
z6PCX498XfURrqbO9020EWcKM3HrIOoN3SCEVxsaxasm3bJDS+xnaXzw+dJn9TPG19OP+dv/1O1c
96wYaUlaMb3LuCW1TgfOG/XXMx6qqh8085P3HRvBDeNX4Euo1dzeeM7GvWz1eIR0ubT1B+OJo/8V
/j4LPlBaGciHXFRYr9yJUXLp7PfeZT5ArCfhda5AwMVO6N/hwB7YiKnT85uvLhv4cEyE02E/WDpT
FueATcRIYaQpG4lkCQnB9OV0MG2KdWFNzhGtbxSBWsEHQh8TncuLBIYITIwuU7GxvJz1lLCzxwGy
8IqS6uLypPpkzvWerlQgX8/ARoeSFyHUUmy0TZEFhcgrdtevQdCFCRE1lbGOVoGXE9J4UkYY5Xeo
BANZa/TqqDEKNPPNxWRUngM8rFoa7Om6lN35qr4coJjdIFfK46/M4WN474i7HlolLAUWJU2x8rUE
tU2lIMMRTy9A4YnPp6aVY2++BrJGzN0eEdB2hqLL1ZsFBX5TGjTlzoOMJwmOTzErJ40SNyf2z1zT
9iuyYcsL9w6wyzzWEddVhhYcDEi64Fm9GEQ7NNlz0jNArk/UzV5DSbr/FKHG9EcpjJHopLpuHWwZ
xV7UzUkaeaDc2NalzCOEU6jpRsn8QkzfXp3DZ1Sybe8YY3sT1wx/sEbOglxua92ryuS2kI8iuWgq
W7/qoG8MbSkkzXjJQpqsfFtPi3xD4QXGdqyVd3o2qsPDUCYz0RGxE6qfH1BWtpC0uu9RtUkxLbdS
fXE+aL0Hdho1Dzd19kRD3ToSPZ/TVcRAgDjjspKsueKBW6UXobrB3nZKW0bxzlkt2e5BIV8RKwi5
1hEs9fjy5CnkdwgDJ2jTKGvG5XApP4cXNKkqFHK/31b4vScMZyIbCq5RUUzCZCtaq+Hy6P06WxAi
liffrTeeXtMnW23EO7TZrYGU0VQED42LvHJbH64rkHOfxyhom6zj+FJUHKCCrRUxSz7gcs/sDEM6
YAfCxDsJP3Azsl/eAZPgnhkCQ4ul/ObaylvePNSGDkkvam8TOKdoz16yk3q7dVCsOJaF6gCp6MHx
28k9hOLdNakDp2c67+9lB0WTSbzr0eno3dVBZpBfCK8PIQ08OjevzmnZJunXtXH74MYcuSEHnXDp
18G4TF6FWj5nWkcgVXAAPgmSt3IDBlFoAP8FddvCPNHNiaH7bncD1TsIFchrh8/8MJOidraSpkjE
nbk5NnXcvk6isLiG4aQlGLj8Kc+2LHvWvg/XYlvoHMQHEWFOJq1QJWa2eHYogk119n+yqXO9vgZN
EL0gep1KUuIlFOPNUP4AnAHp3KhmaMf18Zn5elY86QdSxQ8ah+kAp/S1848+ibZ+T64duyYg+7Lm
uxLtEEI1HIs2+MkB4bU8MBplAZz1X4QQqIFKuyntgpQTHNHx8RylpGPFUThUOkQ4O9seEcOfvNPK
yktFSPygynfd2tY77poH24YoO3Rj9oWCpqqDRz4cvpleZx60wNAlqgBPNeyraotrQsgkEBsDNBaE
NiPofvHk/9qE8gNJ8AwCHgB/44vzimFIv6Gus7wRsaxwgOK2/AZvXzDtBMa7i7iuBh66tIHhQvVz
dt3XTkDV87LKEKUFrufwkwgSBB+n1iScT76WY4eCyS+BZNPOgtBpGmF7XfER6rBjXt/NIGFe61+D
bOOnSExx6w3akZ/aweoOhUI7XiRGzazYL91HiurQfS/HjAWtItWmY0U9CcyQuWQ8bcjjrTeN0Cvl
/qNUmh3dh9cPH7MauMEvJEgWoUrGkqmyrVUPTY89VOHEWcYyOc8wWQPVH1PZcPTN0QOXX5pitEqz
/jiAgptWIs2UwKXk/Y1W/2YCOohJDe59MKXyDQ7eyAt6Y9Cb89BF8RLP9CbYL8BQRejQUIq7TCQ6
d5S9oxfopy/7YIcEPDXh6J4pRusLZdomtZu3vrPdKDC8hEfyBKep4ITXS9fOWD2h8Rk4akWIOcHb
M500LZeFFdmyNSsHy5tPg29nWuumcLbzVBSdO1bEEWp9mALlmmUrE1H6xXcapVa4C7Xyhi0k/nH8
WgsTIjyA1gKAZxHYAwdHQwlNORZ8IiQuRN6mY4LCVYJqRhmWLobh1/OwWGk8X/iynndzS0iehWgK
5rbBHGDSdxXaSLVEtDiWEU/j/abRuCWNoEymtKF95YhS3CDz26AqqX5pDHS5aylA0DJ9iymOQu0/
oKEP0d08ZQiznmXFiP5WUwXMsm/eOVAgPsyedZ2DrTqPGVppC0RG+3lcNi+kuItgUh9bNT7LrcDW
hz2P7Uib4Tj1Ma1c+g78aBhYQV20a2qz83PWHTJFtl97AX1oFlf1wUSkmAZrL2BbSC+EjjVwrei5
+cA7LqLyS+ZTsjp2ev4oinK59wHqkXlSyoxK5ShrkKxSp9YEHBJ4ctdiHkTBdCpsDoXLfV68ZG0r
RCdNr+P0k65wXTX1HAshgDqKYVU9vAG0HKJD2YWEHL/Uws4XxQTlN8M7V7kN/pyBbRMS+890NZZj
xiOLIyeXtdeqcWqA1lRKtQBvjfBNMGgRo2y+ZZd/2djAkPwMFS35mUqN/InyMWCQW3RbKGm+eJYx
opZtc0S/MfcRAwXD1ZdcSBlaeLy48x2UHrh178AI+rP8rx00U1aNXb+dnxeW/cQs7dm9iaDeHU3c
WFE5weYqOdfs6pMt1+Zih/tSZ4H9oW1OEO2CV+7btWUkjxp8p+60DDXL5RQrCwON17zwJQ5jltDe
7UMcXDrejybN0SJ/JML9eIxjJm+k5NwUxtpd/xO/P+CVblZo1LANSSQTpun6YavK1y+bgqqo8RjR
uyrim0vKW6c4sasOrW+1wGxcKaceq7QchMLrFdN1I0bWl3HkFfbAw5SkzqoSud1VKr8p/B50q9ry
TS+T1XJEr9pBjFKWMHDe0d4WA1++CgzkesBhxm0ChEF+BQjx5nZnv5UNtAukO43GjzdKKt4vBXyr
6FvD/LhKIp9f4zarPiLgR3LEkDt/0HdpO2hfOJ/4iTLDc+zBxmQ79klXSLBdD/CXaCiIuco86c7t
6E6IVwxpnw0J62P6o2zQyacuf8zU0518wzabhxjlLwhPR6Qf2eH2A1z2sUQQ2RdzVwWPKFQyPGMZ
zhYHmTA0ieDokXCLADzYRsRTZVhcUxjFpGHczcO07pPJ2oi8hE/4I9nlbfOoWjwBgmA1Vjm+i9pa
uvTCJkGDOQAvk2i0PCZ4df2a3jqilIKyTeXRNvC1WbOCstbShkk2fOa7epVLfMc3CstMKG22/S9B
aumY4foQRDp4/Tlh9LzER8n7YU/hz/lEZlM3F9DTutp3SdMe81L/T6j3kZ6DEVyIVAFOLg9GdWGW
G+PddpPBp6Il5L1gGm7zerxK9nsyfJfRh8Oeb89w5iE6b7xiRYhpxophGnp4bUUy37RkVFsNAO0/
MGsB4rhMJiskp4YAl4NHPV+tXADfZqOu2vDlyIgRBMVZ8qgtBSOzkN5px4HkPiW5/X5CIo6lrKj+
nuICwV7+MIP8d9c5yGMrCwVAc/vswW2ki68UTjgP4Hy6nF9cpWu3hH64/mizncWKKpSQhmoe2ZFM
13dGHEOwWEGVDmDcVC9KD0cr3EuExvLV4XTsnpCC+m8ebTP/bavLR64/bPJMz0Pg8fhMIfMReUUh
UtiITa7U85RwBQPQgz3qCCbwBkQJs1x5nf4LCp1WZMLbJZk4tKGLGbMoH7h9fdOsWzUpZCcLuASG
KY/zCwP/LwkyFTtWtpluyQetX/23tdsVVOjLRgbRio3eWpBE3EzJ3Xrygrj4BR37Z90qiDinS0Zo
nyj8wE/E7yolhTr1run4c3Cirrhcoj3dIZ9nbhkCQiUNnQpB8lm2/ZWn6x8V/GQzt+uTG0PWU3Xr
mHveKt3knQeUkk7KN3LYtYbmicuKjn6bHQ96nb/9dvaDXdg2Y40+KuQ6dWIpHsk/6hQTtdJn1Vf0
FQxmYJVp95U6GnlmLXHMu+NpaatIWkNIqiW7ubsxaxr1T0bdwVTcL3AFuCF7/NzWZDG7IxiOFc6i
Hj6PQXUycrv2koq4hMselI1u7KvfF9WXWpav/Rrlv5J7dnfUSf/3Cnjb/pAsusGESBgTjv1HYOM7
kQ7AzDplz6vT38awf6Bdb6tYuTb4+p5blfq2zeRQew4fvidTuh2DzVftpAeFhph462zVX7IA2QoS
Rm00ZQw+W71SEeuxGXCouKHpC8yx9MQYO8ptm+NIG9SBPsromnuraKLAeE5oyjeccbWaacBKhRkw
sbJr2RIDZ108BHEKdziqqZj/AI3EAzdAp2Gq6aWyAsVqbWNN3spNekvaV6WbVOFuGPb20CMMSwly
dUKKlwssaRsIn3J8W8QZFtEpMits22IWshNvyscw43vwzfDWuQjfHA4V7RgXL0T4KRVuWJSCHENN
ypKXWtx5FUU3+MLBUFuQykcFV296qDHX7OhvcSaO1jXpIrVUIy0krZLP8KC/fbuaeIoY7DzGz4+a
d7jFfKukaz1DDJkEkSq74BWO9nXME0ZXyqPA3Cnu6XINaGH1khZGtXn8SmAAoaoZg092nB/UbQda
Y2xWZZBFDjyub+hiReK8PJn9nS3Z0BEs3bnhf/mDA+Dpy/f45mQY8G7RBA+ZoNH0mJSFHXgeuKTQ
6wW1RIyTV9n8vLEPiPdBWWU/HbTaW1LWrWcxz7CxphyoJYziIxzDNjStg98/HOsa6q1rXsFIgMEl
JxWDGgc9eju2RlA2xU+xWU9RBR/UvQpD62jfs6TGgJ+VwntnGwAdcRlnKo/QbtOpi1RWr31mRs4e
2a0BEl/hX34qogG2JLGSMO8LorPFSwrkzwqoCAcYrJ7Ttj15iBgfvRkqsHeAcEprGWrd5mYtdBPG
pJCcVrWZG1BmlFDZ7/gVIyLRonWundmmc8xbdqeIcSkKc6o0xpk6bQhQ5is7qIdCEa8m7PkHrVl7
O4OhjDvnjrtyVufbtOnhj3xOfBza1PCCMJ8KRW1VZcUY4OFSLLohrTm3MxrsmcKxVAClGX9odk0q
G7HaFdgRaYBZt/AdANwQw+0feznegdYct40Sc8nGohtddRUsn8G22JnHLot6MpmzUjTAV4qAb8WY
ZDCNd/s94+OGbNXFPxTyNwEO1LbDqkC8rPTQFtgvx1D8rdDJ+3Hxri9qGlmHHru9b3aRDd6+dAN7
j/PJCPiuU5eMBNmYP4tQD0zOn8AOFLcjQkJKrUsLmVwhikpQNBR3Xz2kcN9gRJchdMAxVxra/jUy
cSea2gBQWaQwZ6XsT4IE0A4Yrn5jyahCWtHzrup3DqJv74OvHdZUf+NVJSUwCT9mg0kIZPdigliG
1VKuo3+Bf9PCRScHdBtVmRyaB20llvQHLLCF4XpZKUD9VQcbCBql08eWVBoy+Igqev86R3opbyQv
7u7CRc6MIRo91TPFactk5bxecqjiCQUOvzFgOejKRwjxGM/TyxJ5t4a4Ary3AqVN8joOH7sYuU2z
C2NxQ8JXQMKvnKaNGJJJhfWrzRYnHEDua+fhNlDmiS4bXGcG/nK1ubVUEKpHUbj0NA9dbTL/N/O9
l1nQGpwf4dfsX5yyolBJnL/cYMWOI15J7BYP8NaJSy7mGOlxUDA4FoTC23nrVMYliYLKtMwC0w0f
N6oWg7jfWPWaaKo05JiSUxV0KQBdk7c9sqyyOXeqlF0CXmU0OJ8qzAOXLkruL8tkyN+z4fDh0Hlh
b9Yt5aU05QrOi72F1V7G932g5DgGDHVUMwqnn3+haGT4eTkZQUBtiA93ExdvbuBqEXg+tvmFSdus
eP0AQnPhPEaIMQHYOG2wByNYfSHSAo46smvCCDviA7PCoHb3bx2HWQ42qUlPRYj8Y5Zou+fcno5m
3ZlnVDbFX1S+w0yHanXS2r0/Y2Q4kcej2Qdk10+pfZ8WKUAB4toyKCOX2FSXMYhcuEH4I45eNzy5
NCGqT/2Hlqh7vtXe1E8WQLggNtt9kQRJxuY4WuYugeNQHFIYL+Z0SAC34xPyoco3wM0yw3fx385M
FE/7mjoko0sEL9VudELm8eILfNvqlQZcjrx8c3ap5sZgZjUUnlJ0NrfOjMzmIHMjmhfcNdB9Uv08
/oIZJF1kZsivrVjK7RS85kWaKzjPCua7uvNYnZg/XrPHxd+L9JOn3VxOj0Jg2o924zwjl0131yYS
Elkn6h9XcJDZr51Otu8qiDFU3ZzVV8DeSHRf/0cnbMeBioAnpwd5xjXfat+Kc1oeN3WUZF2CPU8X
82u6W5vKVu2Oej5EB57+nRmhIAo4z0vtRl6w0d55nk2vBfMEIf+0mipZog8RSUAIZQH5TqZEZ4Pp
TK6o6ZWIS7TcUdayagn/2WWcSl0Gq1bs1z+Y1HE1x/JqtAnY/0p5pUMrKf5j2ReaPO1JgE0BjH8o
5jFZ1K4TReXEAss1s9C8TGvYMLJEXV4Ze05uofOdnIkbjv3XefsnJ72yZLZwmeHLZId22yBmZtmp
96ugUbM6DP3vNdvQIaFo2nQa7jNNiQ+rhEQhVmN5H6P238wmuLChBYNzdF1WBMY3JaUfCBfk8oNJ
9zLcPwryk8nSNlLz9awqZ8hOUXnkbrctAng2v9L3p2aQdVjkYoZxR2d5EPSVeltr5lIjppcPUbHP
eAtonJGsoZ9ffHSawokaG24nN/pMbtCAm4Aqc+Vq0f55CBYbuZ15owvNfTw3/JQYyf0PEX1PuCtw
WadGBW3hdAfgV2Wo4WxhXjLBXpGrhGeT8l9WxYCHxEsoolLwlUDFOivnuHAAKXzSv0C1G/5bzBm0
vJ7aior8UIfw9Po3ZoNFu2iS+IYLQA9fXSx6IDWZo2x6e1tStgYRFEQQwxVIGK1fcMva5dGVnVE4
nzXZXEwf5ecUm+OtyRx5aofiXD8YXAS3c6joFi5KrvM6N9pJSyPuju/VAvFKlU9tZtATlF9x1vLM
CpLYr92mmg/rbCZEn3rkcU+MCrV20k/aggs1MXQnKzzA9eKrqxjhjmiZvSMhIVVZuTQJfNv6sR5A
B7fCt5uMwWOIuQLee+dRULaWMrovkpJ0VTPZ+XJYBkQjK4kOaSoxVTaFhrFJgT0rhFrCNoWpvWG4
1I2oDjcMNL9ixdPvIrqWvXOnv6AfFxKQmF4L30oXHrdBo7L4dnMSf/awIpC+d/Gziy/9COAsVy3E
GWsagwLQj02sWf7kofEYAHk7mVEnLgcfN+VjJMpfZbzNeopNIy6DZJXWZsuJ+1E6WMkdSSOOERQU
6LC/PQShNGFNK2P1F5kAnsi8bAiSwTh7btCN/1HrAO05/5u7ycxIa3XE5mbiZ3zk75UW//NdyOhS
G3T4JCVz5z/62kF3UGUe2b35On7nT3X2F6VsJqGH4gEyKLIK3CPalE3FD0FO5QANv/M3ieek+sep
X2MRrft8ubsZ8ltcmJdCOVq2WdradUU4NChcj2G5v1MFwF6CaSRTnE/cZi0pqbEVXWeiHZlLWddm
fBSJxaQo4bi06VrhV0xaAEU5kiiDg7Gj8KnZvaUbOi9QyrLF1oXnS5DPQBLZp44l3cn/2sjNolFz
ikTNHNodtAbwAupzVqAC2mjnBmT3lLyqvGETP4WAn4Z5ENeui5+hUQ25hIO7TiNda0Es704qneXl
4ln3EGI4hNQBclzJd/8aZi1ExL0vB3U4ECksiq+kzh2Qz4DRA1iQFz1dr2Jz9eZUI+XFMXhmU56Q
amYg0rhmDG20oa/kjc6q3BGskZcDwisRjNIEXIppi5XpWsfEj4Hqklhi9oLcVeG9DJfO2MWF/Jva
MTDUIuXL6L6qI60DdoFJvpMVs1BAvEr0jM0VfNILdZyjZ8McA5A6JXB83GOk6afZqYLn4+LacqOb
FTY3wD5EPYv1DyiKXQGeq2x+UjjY9WSWmhW3hOGofLj9e51OsOUM/h/eJR7bAzAK1WaaU5SiEvUd
QQiaxV6ifaN28Ueu4tz+luxFyxA2VaZacgtnFEBnyJZo8GdolT2fznxwVE0ST9wDS3zwLYIT0TnE
Kjyk48uXT+hk8Q22rt1PZZ79v8aChjP6++UJGjmXYqxRuboy7CID8PRsLvB7r96IJ85oB0LBgIZW
54gkrhHM+LlHTBRp6+XMRvZ9VEyfmy2wYNxsI+Ba0k8G23OFXOnQZQQu4hCeOQPf1hevWMHxF5c3
AhasArUmt79h24Qz8vgJFqMDHRTB6GhkdWV2ZX07sg+rnb3kH/K9kBLQpyVlQvI8NX4/thkzDQTC
oRBHahL6zc1SLEUbu09UQgQP9MvW3LthkTaKtaNJmX8umGWQw3qInzw9BPQfcHEk+5LhjcUjC0kW
ODaJV3Iutqw2h+CtslsmeaL6XnLnaiR7QSUmoMjlV4SclWkEhIfVIYVpuWrukQ6Hqf9xKxOmkYn1
z7CnoAZVkkOEuW037/TDFBxL0bTw+4UuPtrV1GoDd2TJ8WERacABSKMFHrR6C+MFnO/p38puUCUI
F/xsXCAlDZKTSITumis0hV3thHBgAnERL0be5dP9apuIqbWSijmX2nQ0OUd24HKopVUnPzIvAkjh
F0z/EjwoPtX/Vm7mUrGK1Uu8kNfznzFfajfX+aZFWgqfeeDFPC5a5gJAdqrH3K/9sIB0oEodNtbJ
f0LQT2lngJC4D756DbmmrwxyDda+EYK/vBuzNvrw7goM8oHHpmCT7QwYKymIPtmNWN6B/oPgdIyG
pSuEdNVi32uVB4nlHYeZ7EH8Skiqp9VdZAgZB0XWOGV8XnBx+TjkoY5++zWLnqgIsHW4G0tP8dpv
Ou3x9YLV6xB0liWAr7VTZXA8d8103TLrvPs8oSgi+94/6M2RtGBRkGRvWxw8/T69ApMK9aL+eWzu
req8acw0nlyv5sJ3klMe9aoGVxy4waOHY2xtU0S81Gnwt3q9B0O+XDlwBjncCI8kNAzPWo/LazCw
ViChjOypUsv1IVu1h+V3SG9ravSNHzprRNbvnRtd77mlVQ3JT19AiuJtTpeOs+AsH1idV99UJWVD
rNX4O81/MtsNC3CrZXIBjOAL70Pg/SXRYrqTAhRVSKQbFDQxkFmjZDwvLoaJ1t8Vk4Vsdh30PM0e
IGbD6+AVIP5ulsW9Sq2Fcgjac0lFY7YNhIuCEkeqaPEZj5Ax25AKqq566UN6K3ySPm7+TGPqn36J
jpc6vBAhEO1lod+Xf7g0k8ZnK+k4DEKrPHDuTdyRDWVHO7DX15uvQtZXrd0E1U00CI3s8oryQE47
IwDCr94t3us4/6uQ5fgxTP9E4RX8cP1Ek19BvAOTc21Yp8gRSQ/cPtgojYsZ6tQsmCJBva+KNxA1
l1xXcy7DD23erNBZMpZ/ZuSBfCP4VI1GTT7iXlmjcv1GgkLDDUvKbpfepYzNLuBg/G5DDOSrgBAg
+WSeQrWTcu5ekkjHgQ8nZbauu3Q5VZEiSEBgffu9fU0JsnGy1HErx0K7pH43Peqw5UzIIgHKejKg
4lHDzbR4cyUCz9eoPbArlCm5X6QNF0CR/bEfb/9VCja0MlV1dPQsmBASxe0IMMGz+Ji+g1Me9Fbo
QE9hWugC52GdDD4JFYgasiYNzBKmGTuTVXJEPgmhH9ItE5R2izjsEUTX+Y0sSd+nbEwMiME3wrSy
r+VB+ND47E8GEE8c0YY0XcYDvK6u/3CpIaDXlPQkVy66ZxqDnxO8vIaGpFqBpa22xB+8pmChtxWM
vbjRhS7KIabzekp/fFzPVQhv+048THv91f1ac7/6nbSMAKE844Es6111kAVvMdnJjHlnIOTkf4MS
8k734SfC06zx6OjXfCXlQkBho7bSd5L/VhmQQ8qbg7Bo8nUHU045VaJOgXvjX8xAPcHpremH/Ua4
pLQeJAzuHPkHo7zzSzhflrOI8LwarnuKI3UHyv3F2J6liC+zumYy7RiNjBdn9W9sfZu6/ZcN2FXJ
vz3Qeq/f0iWMno3Yqh6f8p3uRhf/aS9cA5O7vOyxgs0rcu8l0X7W9xt7k90KmRZ8WrYd3GGB/86e
QIL6lHfQu5uHtXuQaPTlZhS74guJmAyU09SQrwRPTdGilVOR27KDvO7ET9fSaGcQBeW4J9m2A3qB
ovNb46Q9b507lx+WVzG0amKJcw3JNnxU3oU0yRrbOqjb5qNgeATCricdYn+eSkByhc7IpPaN/bJg
eQJMmNL1Lzg7ON07461wHPAR/xHwjj9Na76U4bcRtklffq0LqpWGWr7SxC4ayix/YTVncQJq9grj
J/2sGy1hrnIIeD3LjdweJMWt7wK6VeUq/PBBiudx3QRrzetr3BNRSWTPzg45O7/ktCUVH7EW0L7H
Fq4PvcT0hIoidfXraiNHa9M+OanUTJ5IHuE92WZgLJuoSMg0hPmF03h42cyeS5JbCpkldcYZGgcD
xyf/4soSFDCihSAZPtlspE2i3btyxXLYYz1Ps/woBTdAcSNhLjGlCKnRnzvrjOyh9G2/a7u+zxkQ
3eneuWfRpm6oqg96Qfeyx8Ij7Mxj+/PP1F8Zamt/wdbKLdeIxStWWE45vYZIVx5YEh2LlyQ3ZFHM
Mu4bu4PorfCjUBx0jchzebZlEdqufwofSKsoR6x3PBsALpN8eltFVAXPlexpIREpC01ydJQ3XHxP
6juvhJJcVVYMZACblVsmGndFpw7JssVgo45XmDeVHsUMYiuYZIHjyM9LAyfOhF63hr1qVdWSyeE3
FfDZLuOk3dFpQwTnUjc71uBCpvqML/ihEZFjoiG5coSRcz4/6Z0WCC7BUGUH5sU6o6qmJLMoT2Q3
j7VvNau9ujlEcTo0FCDa0MOyu4IaoCzj9QDQBla/AM5ala63gN2lJwLgEsjImLEEbYJ1zzgwOxkj
6lQLgZK+6SYOtrQtk0hUdwP+iKH9vuQx/zI1Ffrm816LwnjG4ceKFVNjXv49uI00mZUv1oMU8mdy
txLRLcxLxYlUMon8fJtqDZ+Vb4qpgoB13k7F4p2wFdLeCmwpfGI2C+THFUMuR3sEcKsJLEjTeaUJ
GTp8n0XjHryLDzfrg7SxK3vdOYb2jqmTXuFe7NsbdiYz+9VH3KsayZTrqH93wmcowP4b5XI4U3MH
8JgBQt25nsnLVSn9zAAraH/aYrUUWpOASaWmlMx24GYNBY/Y/TJ8YcZhxUOWQ4rcZiF5pf6oJEKK
QPWNt/EeYcmwx3O1TgucGZQIQgl/Mz3FckS1O/6miUL9dWhKUN0/J9tGAXDJ8Hz1vSdiOUKtEdsQ
gR7eGAJPqDvSN2L4eQK/QXYc2AX5de8UDS7J3uohSimcF+BaDxIuil0qjwBOlZnyP9cJVEyZP4Lh
lZ0lMKDPnJK/IjV4QyWMoIW03cZtj0HdSneca1X1u+I95/b74rYgGXW/GVXH3ptzPQ6wNnGZB46T
aqECG2RTp8oVhVAkNpLP0hbH0YFVeJCptL/hgkpGSDgAVQxMqDnnWy6ljKYUNmgSwPHyFlNzzRyw
z6wykl79OjH2beSiXvfNvTtilaacBNfUX1Z5as20AGF5nqoEnxhAcKBXDk5WDICZiW0+DqhwhUZM
EGTffztOyWeP96wzURp5Llx1L0BIy5p+k8zENVjydHPC1fbYCuqnF+cr5EfrTxFi15GQNqTBSjjk
Nk8pKpD/eg8s0Y0R37iNwT7jFwN2uC5yVgissYBKyKRIJvWGTpWOH+ekfdjf2GBuGyZn72T/LtKw
qCzAds3DhW7lNKEqrO757MUGRq7m8UyXhvPofLZEqMPxxFunngIhJMzoWRVZFZLn7kRdkXkYZN54
sh2Nebq6jOKcpelSh7GPec+WVPU78QgGpmkABm7rUpFatF3kqniseJOCNrML5NfqINY5/vx0IBIv
HFu1t2vz41SyYdELH5FZSA+qNLvM6snbS6/bxmMZtLyPUMKM529C2Bd9H2GXGi2svIr0DX7Ghhab
8nrhPgAKUOqObza1S0pDznDkFB58TczaG1o2YrHNk/QTN/MzQn20MqPatLB19qXM7uCWPBeh3iYa
GnuVKe6ZhbzLFf2FV8zvMBH1RzNPWFc5Eu+2QhOfG5FkZAgSoPf9nU3ocMMwombpW6afrI+m+9QT
NqEGZzsuQJ8rneXJZxCvl7/aeCav+Q3CYkw0mH8RChGQWOO1h3lRiWOfX2NwcgQNvVu9wI9ZAURH
kj633y++br4XN+thHlwo7CO0C/OOT19iJ9B+CZEomMxILRMgCKhTUZaVz3M45gzfZXBfLOD1EK4t
wyXcE3CCzGf7EN2VDNvsCptcLTepJ5+BqNiGVsmb1YGlLqWVIWNawtaZzRtPinyXBpu9/EQUIW3u
8LQh1vmQFGRyn+Bpp5zIaCGS4k8kPdt3hVxBqip+2BTl9wjAoHRj4YrKGybtI8uvPoFgwUXDUfBl
2rBsaWDAkc9rLvvwOgL7h5mIulbjPermNpPezkLaEQ+SKF8B6ZQ3/LUXe2COo38yDc1frRQ7It3A
KxvcGgcSLmxTfIVqGs8OUxPzonHOqzO8irsgZ+RZ2Yx72moUML0w3lnIr5Bo8cjoh/VatLYj/rH5
cRCenNGpw3j2/ppsVy7NXaaCuP3B06IDhe4OWYRw+NS2Hhn+tM6Y/pHyb1JpCf5EYOnv8AMxHfDv
bI0d9UZ+cD1+QLtLyB23plq+j2pLWQRfJJVl+9JmkA/OXvjZUJsI9wJndM/8fI0s0a3gbJX9cQlP
37A9E9UNpSf05Ed+CWr7LEmcLDGqEWx03JYcTTsTa0vDY2BUNLaV5nvpUGyasm1w407K/AwDRVEs
fgYJuqP5ZWIQFc4dmWPmHZQVZvz7KbLcZcyruiZwRuMjWez/EOK55AbljgTrJpZ6L7uq2sBGzn4d
SZONqWlJ0AnevPH0Felt0UM0erK9115fztXT7j0SIT5cotXr0PM113NOSrrquNBrjt+pthjFvQII
NoY266DTpeREH2asbRPcIOYNI9U0XGgUUlG5KBhSTfF48i90OC5EKbqii1luVCh8Lcq/CbO71s0n
8PxQ+9clWN36hvu2HoyuxuhGRZlD8mMVo3o8SSiHO++WYBHDNRQTTfhl5n4qjzQRKTT5DraB/8lP
+VU7p2EURcv5bt3IF9hXBFYfNzDP4sYp7wSB0knjAl4bHJ0LkphccJQYUG7j5IUVCv6bRWm3BwTF
506fttd+/D2tqptvMOKELckp6yxmyNKON3e5LQtSr/RuliEWLb8CLBMR7mJml9RZTWXOJdsO5dE5
jgOC+zT+ZXOZQT4K2m/AfWyyY1kb8iYTt8pTJIxwf9koxGFhpEINN2pIDpEeDE+DH8wMTWMucnrS
ybqqV+EMPnYuPQ71mTcFtqM7ucfru7PkfFudvkux0Te/lzOA8aOEYCcGmCSTQVnZwv+RoM1Vzc8a
IQeX4TFjahHCGcNPOTeP5EBqdj5QTaqhacI5rsp4nKU9f/mvBT8W6Kez8cNITZlkZJSaDTCEXzI4
oAm7nUBRdGNIAomY9h/gXRmEWL982/JOMfEUFBSd61ZNvFFIYohaflY1AdEowbxdK4o+yJZj7gL5
80Y7YuMoGICz1HvggE8YCa8xWYa7C/y+rTD7xWmak7WW0vdDClfI+drA7RU1fmtRCsGtJnQT4F+m
XoLovcRVplRKnIRZitQ7LLn7EoYN112aUtNxydOYFRL4FRakaz+UtjSfvpQeneTPPsYUgHB37pQ0
wURx3XNNgFmTMZ7DFlgtNmpoq0BV/pOditnOECYdsNZDWvWABYMUzWw2bGRrPM7AxXa+VLzOAOyz
/A5sYhcTzof1uhtHju7GRabh9Ivfo92oIrSCbkpFmvyGcKJY/mOg0HcrlArlpRa9ytFYrqUg3HgR
9H8QQeDPSKZYmRtEddmBeZdnIOrzH0h5JnVtxaAcmEAM9mn4QyjCEXwFuFKXl3YUw4CY64QTrQOH
3V2k5huwzawtJ+4RPvpUVYXYiCpVOIsEFj2z3J4HFQSvzm7ec7GdNREZ5Eb8z4L9FenxQJYAvX8b
Eu9/5TLBrbAStS+7yk+oc7nRu32QRlxIMCl8LELCJz2hWUbwbDZF3GcRPZUoGVGTfQHlg6qGwFTr
r/KRIXlc+Ovb5/5WKeqVRwUwmyTy/lgDXYUL5tGRULIW7kmZ8dmkLZbNPWQ47945s6Dve+rvlrnU
0p98Euh83ZtB3nQtkU1Cks4/N47mx6O4Yq/arowq13Gmlu7sCXwDi5Ir0EOHZz7aKZcvEu46gxrF
KpZGIph83DLKcptIkTzn01iLqizx3GvitxFUD86vbv51jMbVI+EoBf1gqlhg5O2aoPlOlEiXbApK
Vsy9Q2MaVPpvlTHFHIzo6rkgvIC3wcgvzpzkrGRDMI8wbObr5sWC3FEZEjcX8mpsFCnI5n0KSEXo
UKHqtKx7NdtDZjdd7CkXf2e90lhAQpz3FNzpqlv9+IXRZozXUI0UEksQt7Qdv06SR3XU11FA37ti
AbCMin9gA6+SbmxmaS8MKVfVlaHnJYDpmx1R8sqglBNz7zK/Z4czu3/qQ52XpjeofZVrt4HcmjGF
NX03PYhBX8BE87rdTgcdpYt8bILHlf9sJk96hYSa7yM6REr9BZ788LU45pccmC1k8R7OiH8my+tL
WhUFh/pdzjcaCR9JhW/B906WNGNTfdLeIJIbE3dX/XWOwU5VXYK/Opqkis1exlvXsOXSwu4PSwbt
EVZECg4643A1AT8opvZ3VCu9f/epODpvIZc60/S/YGZhbWzQdAZXZMv3e1q5J5fcbr3VI3pyU9D4
SXCmif1e0zxSfwsoyjBQwt8nrZ1SoBVpUqDiEYnMH8W0Jk95ntFmljB1l5cehiSV4FmUoWfK/Xpd
j5a8Br9RcGftcUpCYg7xv+Qx/3E4KibaZwYyUVNEk8Y+3+GP8UxzTQYwsYj4aj/1whwlZFypm154
SsqREjMbl2Plet38S6imPRZDKwSF2gO8PWf73iJerp3R/dSJml3ugl9PAfh6xWRZ9jAY1JDUkfcG
viCLVh//7IQTunODMrPpGoZp1QlS/duY01DINAYkFe/UeTut/ds3hMmLbX+/M2OQuMlgpoZUqdmg
p0TXBsqC56IlW4HL0lL738FtmEtEsGLXjntEaGYYhlEYI3qutWdj8xhfXaDeOC/vAQgrMfk6Nz9V
d11lM9aT2MNDYhKcC/k/DhDf9ZoKQx8xeWO5XLKewqjODPXzJYb3/CNnGIUhUHgNmaYIn8/NhlXD
z43iNX/0DnUUQHbTJbib+pKEBTD9cG1KXT2UTDEEPsLUR2Wq/HPMWEPW3JHkkePa3mQtU8M9R0Ex
AjkHWqmMHkS5d7qBMolbgmBaH8WrNefSK6ju/CQCHNGBYoets0JT8QqinqK6M1eZiCo9xs/+w3yD
zsJxm1T5CgL97YoQ/H+QTZ/deX3oYpUQZAk2MfbxgBTxh86lz43w92+BOQ3Ji0n5LDw9jEYsrt1W
8kuSc0qRRMYj1d9RUAE+OIkPtmqxerriBIubkdq+xZgbYeiVGmma3QbWa96YjUKPWcr7C0COsATA
gpvanZ3EDjx8Ien3Cf86ZjOWpNPwCgYc2GVE3kBMfAFqf9VX0xkN9pettam/tSeIjg1/28TMBKeA
N5Ka4V/T0a8JJCHtaJYYXCCHYDHJdZjMyo//dYxqsyHUmmYBrOBvBIKrjV0VESH4ON/gOYnhKc4t
HnLOe2pUHLxSVsBHls7lR31Py3MzzajI6XRwAnw0bGfoT2z1dso5dA1hVETuiLrg2/8lCJUO78+g
Hkwi1MoCz9d3jXVu6t8Z2fkxYZTqY2nofpqmdZEkSOon5LD1uFaq3aEqrOXLXSeq9MPbjDgx+pK0
NUs/USpEoe7eBTpxXD5n09tvjbAjwTSWAFhhBOm4vaLHfsnyFPnTtsDTQVkR+UAZCpIA3sqH1MiZ
dfF+0kZMdMH2vmIel454YcRQBshyTqHrrHdsujpLRzoNgh1TU+5UlTaeCeLR4OChBkll8lN7dwY4
JSfcq/jKGBH5JYp4McxHXn3LWZqv/lZIZix48jiFgaFJ+J2vDc9sjEeZEQ+dCS+jdD2PPmz7q1pf
hsfRhfjY5vjMzFyLL00WZ6Hg310nGYaRYFdSRciLwfEupHeLTHOeM9QFw/QMesyNt43NNSLS/4eI
kN/RZ+iwHx/9c3lPI4TaXFqtVCrPgwqdlY5QN0qmVzxJRvuFVADNsUUENzeIpmIAGoFB0PJQWfii
/Uh45v+1ZZdDxIJZ7gFUU0fDK19nG1hdY27xxAjMkMfVLd/aoBSLd2Z8WZNp/Iiwghf0dYiAPVj5
cLofxpgFtbeptge+wkxvP0G3htQ7tjY73yLJYD10cZnjjMnciLNlHiBSSoJK+k2s1+JpcEx2E2RC
LduU/KWFDJKUi9exT9f0xvuIkPPR+EIVsgaeaW//BYj5KHrtZ95ARqUHrCU1TII0noupRL+PJZQS
OpswdXJooOF8iuRRHV4pZT6x4okTZORj+JPcxUARkXn1IxkM+GViKkSKuIFCXTN0Y+DZtAvNNU9r
suMhOERZxkj4B+RLhye9xmeoAzvxw7CPBqg8lbXjHy4w/S9bYNgRd/nXY8iffQLUOd8vxFkqyB4g
FSk7R9M2lrZQbgPl/ORLi34kscCfXW9abnDBnuulnGNge/TXO6Wm6E3GwzUF2O4w2THZ7riyB/2A
pBrZJNO+8D87CDw5iNA7ROxALm0PkUC7MMjQBC/fxANYt4USkW7pECNNQHI2L4SrloFlcwGwdAow
4iHIfJr4ElXHKFI9Y6nL/M63QwH3SJe+mpl8m6dtM7iTB2Bne46+j213Y6Qmu9zK3EvLbjPQHlcw
aqZaELQbp2Ezmeokflac/TdkgpPN44+v0xS9/TUXf6Gvmv4TYkjERlhqACnLXc/sOgCpMGpQ2GrB
T8TH+nVpVplM3sAXdR4xZyYj/zh7igE6FMgoKU6iQlYnVEfJNGF4LQ1SGWN3iPrjfAlOqMHsreJW
/x5dl/XckXI63ZglMdGwAXmGMXylFyWg1YpkM8kULIJETuMwlheBCdpB/H9A8q+/mCW9ue743796
tgevF7rfkSAZm6loehGN/Frvhm4NXPvJ2whpNxp3AikDKkDP1bSZnwqSKtOBS7EjsEVtECGl25QS
ugH+xK+pRsf62F1O8YTQDtFWINuETPxyv9klZab5WrILTsS8+YyKOn2+TKVX65rCal6OlFIzhkHb
9KolKycAwd1/F2d+Vm0OGvohvsqM9/GuJU6oGw68hQo5z8tvDDCGUZxbjNaBr07tyY/c4uL2XFt1
fvGdqggkWgwsgU52+AzaOxseo3pyI1TaJxE0iWwPpZEVnTBqCm+gmGnxPTVLA/1G+cm7LVDcc2Aj
NVdpPjXVnSIEP9yQNyNjt+ijlz4aMv2miLOTuOcnVbXc5veinK1NaJmNsqlXCy+Mml8SjA/xqPau
CYZEKruHUif1N39KGElsIt4PSmTFuI/84ZUPIvsj32dUTFijOmSIbr6UKzn7nq5gvbYlmaQTQIls
KqM+vbE6MQASZw6FzsuhYEial37APcS7IYzoYljIqg2cUXMyPr+awMULFSOETXl1zun1z/4vYPWk
BFWv40ZSuZsgdAEnkdbDwVQ8UzQNkeALvKyaXQf0T0+2WwuU5HHHwi/k9JSDUX5Hl6NREKaEDuKl
9dtSvejyitZdP1/vJoQ7j/Rupl0TTa2hdXBLhM48m7DXN93Cfa0yVdluj81h76lqRP04NN3wC7ae
ovWGYxTgZ+/RDkpLLx0LPfp0yL+zRk6sYw1QNpzWFWoqnvgjJPap+9sY4g1Z3zNe+gU8TWXtDX1q
mL38Es9/IMhSdbvA3uuH513jfz96oACDnvtcDIrn1XPXWBmAcfinySRESzXD4+uXjBqbjHeuKf7h
OA3Ve78CE9IC6p3WTeZuDnqftBI9ZFaJBdw4DCCzAupnPK1fCy38IqtnJgkhDviaNF0x+5h2UeMo
RNjHi4T6PUlmC1wu+RPzRSXxm5K4zKzgl87oLdyob93fGKyeqgMalhAqElx1L3Cx6u7EzUtZc/3x
fIBWZS1CxsprbN2+PInlsapOaE8nz/J+1qB0jySQ+adcTY/VnmsVVgJGQ8vcYyIbIKbpfsn/DDxO
iMtNdhmyd49LO+EOrAQxGzdeU8/qGWf+CaDd6FPPff2YUCeN3UDHuFB18l/IVnNfE6f4pIHb7Iix
NFKJoRippWtlTiQouv/umObux9SlDs33BaAqYn8Wh4SlCaD2D/gI64ARSTNyJQwvnVf/0RYAKeot
dE7oW8Zr94P1nGCgbY8Yx3RZyIA7uTebgziC1+LH6cQmEl4BFBbZtjJFEHkc5+8mFHN6uHNahIs8
LP0SBNKD/EEjLe9TfSfI315C+fG8yvYXRXAbO2NiNdXvYaYE4hNwO5PFRg9E9r7a+Auq7IJ8eKGz
laNfQ/Iia4xv6aB0fpnUFZrIe4VadPMu13ObyVaQlM7lV0iLdzGy9Unr1pagmDkBjMd0UpRdFcew
+cSGH/TOC5OC/2qkvcEEiHBg5b+JDKUjea8RT57LHM2OydW3wlFEhPXuK2EHO/dN0ypUk0y5f0bx
Q5+UXOWXdy7Vkc5Gmg17rpOLeb1vshQ7bCdoZS2aXGPCMo7GLR9W1z+peywoN/qYI1IBSnRsKP3v
376o5wseGUAct5ZbCGodrATnr6WBnATPsJeZAmZ25/qhQzV5Wjsxz2IF0wPOmtn8GBPg0u/d07y0
TpdLpQZMdROqNWaaIKbA95AwRU9n47Wc4XZSKCOFQjEeA9jET5Syqz7mW+otdoEFgl7Yk8KOEbQt
IUdiWFOpq3xEvc0yTb3LdzUKGY/MNTQXANpiFT1OiYk+tN6cHynWu0yuu8GdDyGHa/nEG4q0Je7x
1PX7XMPMmno1TtcH0Ru2Hzvy0cdO9ygHI6kpELR+VOS6vzeowJS/P/714bbIBy4Z+yt6X+NPJBUG
mLs7dY8HlCZvmD9VJiTEsysw9Whmk+KXwdFk1ahOINqm1hSZ8zI1XYYW1/+/6SIDAeSYI54/6fy4
gmN+y3BWLz4eUWYB90bI3sCn6EB1SS+Ttvl33TcqX9F4hjxj83UfR3fdhap5yibMBRqhrmeH7Dok
LdiA4nuKivLjD/gDEjNSOee8wo3h75N7RQmdlqN0wPs2BCtgiWVcXBHw7TO14dUZJTglXLi/lLvb
h6kWRCr45mi7A1aqKnBeY1P2MBe5qav3MZXHIKNXXy4HFFNego3od8LCo6Te5KKYpf5cNjd7DlVk
7PzUPc+1bLRHq/hKujoDuw1let4jDURe0cSN/eTH80Eg8fyBVAl08wZwJCyVbYw+aHDA7wDStGnG
ZBFH4wgSoydaNBisRqbVAxH130+u3RhEpUXzPgoapt/B0vz8jYi3MayW2yauNeIFCkgMTE/3iP9u
ovZ4f01me9F/gbZ8seNGRB9w6nlsxJqGzvaYIcqffutmRL4D7CofTCyfrJ920ZPu1JXU7+KSu2F7
YJNjn4XzRttCqChRhUl43kSAdli08RZN6bDeMBGxUxJQ44mGzUQK+KUwqu5z35udb7WeBeFKNG6m
h7xdXSXiHRgcGk/f0r/RY6oNo5rtuavE8Nbq6BpDK+FKdhcNkwc9WxjJ+U/27unXmucafX+AzD5U
ufSghKBdXMRgEfS/rZjCrAIrNOyE9HhRyUKL6q5S16kA0BI13jG9I8HyJ4g8zCqUgPXwWUvcApE8
ZGwwRJiMtQRNiF6qv1fw3KZnPqM2ak3sRAydx8aQ6zdHjagEHiG7vZcJleRQ7wZOp21+PGmhK1Xa
kYjXTahQ5ijJbvYLqu4xlqk0zAY+oxpTMovsZTjJvTpLBXussACGEhvqm3U0d9MDc+3IUBQufwPe
bWD6hrjQD2n2HsgVn8F2QEgY25UW0AEKPiNzPVOdXwj1BkDNB/x4NaT6v5loGI5ytE7ybN/KQ3VJ
WE53TpeJRqeoM7X8/Mm8101IdrfbY2PxOeLaL1t9njWA3GV/1IWayNLPZISdNtedXVkFcvlCb2Fg
zb1Z4v95wTXpHCPzniZn20NPeRGoua+c5oTlg9ig/jJ4AucbwWoU9yrOatfhEbcVMcrVk/IgW/ey
uRinEItAkazPK/V8ID9f57b7LGse+/pYhTCpoybdlpGqnEaGCXcFOYnyNQj6fMvGQgsVheVugu9h
4TMGTnjOcoawoxthF0m53AekdvAtaaHDXjnEmfI0haHKnFXvVFxi94KkBflwjJuIHlE2dfzyh0th
sFwDYO3hcbV9cVUnONfKbjqoYZI2ufO01GYDY5zn8ywmm58wPKDAGm9SSqZH6X4QVpUcqGGfaXgC
viLQkQThMCDPbLk75d47akfm5xVCLot10XfJXA9Xm/Rlq0JoYJw9tqUuDlB472j+ZLQlvV6xZztH
VPsrrtxRMO02lhB3fF8qVfKlgSUDyA2Ud0AFQWU/UYKdXZG993Y9PfzfdrxGNJTdT0iIvhn8S2W4
WU98p4b6kONVqJRO/Ka+GsnEtvC9sLhC4Hx7FU4eJBIVNuw71XnKTpW/3QETp+n6xnTF8nN6xyDl
LFg0YunV0WJpuxRJsgEhBrBBnYNXIntkBY6YoF9JKI9w4vkq3MMPglXLpNE7AxHgPEp4J3P0/vnn
oQyShXK7J/swqgXjHgStKWC8wwmxPpyDTVM909BsdZbUbYRkc/vKWjyC+r+DYar6v+gdUhweenzU
vvf9Br3c2ZU/1bAvEchqkFuNkyeoNzAYOcv6UUAkcd2M6fNXmPulXMBYAsJqS1CALk8CGGHUK8FW
G3QYHQ7Y7zWJed03zgJax6G4mVh6lKBMwKNjdgdZsktdHD2f9GN0kLjVJhl4dTeGgtzMNY8wsJQp
K6Hs5JKARLmc+q3gLbO5d8TiBRo1Mtg9SuabEuTABDALPX6TO7LRMLIr3V/j4HvEWolPNCbjoSXd
13E0AjO8tm1o0FHaXC5Q6jvIyYr6r1pLzwrruRpRqh4SAMToV1erQS7NbRXq3Y8H7xHJkyCTGSb0
W2wKA91en2cA851rYnIQXoEErpngcvEscxxM0X4JDnikXKXM1YCdo/wosVuAqAdc3+D1WcxBuEJZ
tyX3HSbCmTsa60wOg3F0yG/8K2RskvZDmGtreSaj+ZTfSf1JxbvkQ8me4sYTw/aFQp3Sn7ocsbiS
JSo2V+MYRKsg+yEaCtKyySfvSmRAgbaN8hNzlVxQIEwUv4+sBrjeGD+Ic6hZ9GOn0WGpOcuX7OlJ
RIbILYYbIo8fGF9N9g9ASm5rMK7RAS40rphXPP0I8QYyxeUxZ45e0fu6AT4NZ5/aCktyPf/jVp1M
OYIx9T+63hRV7WarwyaNr83Jp5kb1qvfC78VbWoQwIqo7Trzq77jTkXIsCSsVQxsTKnQN8WuoH8n
XB6FfP6pOxHHLH8fQsjZeeBJo7gtz+HWjBmrdh4edODdOEcUA4qoKybG4Um9P6ADObHjxZ3QshLj
SeJkMlQo0ZPUyyBW3NPeFDe4MyYc+9gWycGbK4/1+7PRzY+zwamS+BW30Ja5MR9VvUh7ekTgtHDZ
Uyjx9z3RWTfydEvxEzWtBNM0EPqjhIq1hNA1+TlnVeRf1iQsb2d9E7QDN3I/flV6xdKP1RMuY3Ak
vCpobkZDOAWkv9WGjw70jSTKqVkDV7wRGdYVefN36wq9/fzkY16Ungy+JKb0jKK6UQB3z99G9kl7
SVzdILs7rceoCffzn0HcoVxF7g4vhlPqW7FXXc15ELhqqqK2XyOupPNEzY/VnJEcdXqZieFrABPg
lLzxMFD7vZGU+Cbujjl/L8EEsL0O2D4MzlV7g7YsIhwkeSCbiTRqcob3fR8BAdCoei+U5jglyaDd
HhczEUWTPKa9kyCTTmbfGLzupUGtO4bANPZqUzf5QXdxd1wZKORDRgF94gR3IFkreRdO6PrrRBEJ
bUghdCXz9mPot0n9ikx3Bq2lRrVXbNJStN7V2KizmF9PD9Sbw9bRpYP8JOEoIsAsPhK+G2pJp8aH
2+dOdTrV1kY7Gpe0ds8xWAlw9vV2f7j2aPqYvvV3+pOg9bcO/ebB5QL3NCZk1Hh+AgdymwsvytQW
77P23fcyj1JuO+AckjASVgXMhmya4cfcvG6pPf1s8yjmg32VtMsSOAC3N9jP9L8Rf7fpSkC3HTxa
kFoxHKwPuIWW5Q8PjApgs06t+JpONq3TAVZG9AnxzEUp4jIFANyvy5kgm9/WZRvyQ5tzCrcVWKXo
8hFccPJnjN1ZW4d6xTw3dCNZFB4n//hf56wTNSXCO3LHpWplM6GYJxPbmvbNFfOFCCUrda3ch3yE
33atGdRo5R6GYvHk8xI2rKPrYmIiS62qPZCx7wUj2EF7rTQDJTehlhlJ/QM59nBh6Zy4xOvs9TTY
BeMRwWW2yxsMMqNsLHcDytjEyml6CoQGHDu3dRDVIxzs+jbnhdCr4h3noeVXz0obGzgkfwMdt2Cl
N8vvW2Iolt42FBSwZTuS6TzklAL3rzJ1XkNSBqDy4SrXoGYKMzFGXYMFE7uFxu6dj+D8ulUdbO2Q
1udfrKouK4QX/Xkz5RDviyOUn8z4YQWYPlx3yKE7Wb8oV5phD0feB5Qb7zQ6Wpvmyk5ksSRne+1I
FWdhYTUa51JegC1b7QykloigUwhicb6GKTNKA+1tO+X2fltQloKpk0pGAhS/jGYikXflMiRhjunT
NeanwjKBIAXlNah0w/lQGGu9t5AjjB3pKP98ztV8fGFnDvDKCPRhK4fyDs416V7lL0ynrfTF/kFp
z3TKJxJn9WL7R/MiRnczYNWo0s41JsJybG/DRmn3xGuFaCx3sb4X6EtRte0saYGpSXtqjgdGddeo
WxRZmWCt15zgreOGasjmsd/aoZKqUvrwmz1EapdRNd35aDQvSyJ6UzstzPqXXIRZXt4HDsbcDJ7T
olfe9Pmm7ms38PuT8NlAw5WcyzD0yc8WI/gGk7iel4OcF0gnw9K0yI8KMYZNyUGk5Mq5MfhUqvxR
5wC9XnJITz7AjZ+XjFQcXczKilM++BBGysOki5uVqQ92wenlryke0r0MPrydbzXsNx6r2xAvxY9H
9EbZtfxiBL1ZTWFizS5CfXzbgz5PGFKD9sYVib012/M1jRlZnfo/UuHPdMaGpNrLnkvVVISGc1rO
em9aXXphjFP8gugaEEFCzmFwwexlSNrrFK+JpCFP3Z+u0zYUX1U+3gDTbYRx5EK3uBDRokmKRukT
e/JMIqgHbxORMqrTNVJhuRlH/SMEknnh6jIM9KjMtWGdoJLZWCptHYeTm5/UNFtzC22omx93YsDs
RGY+t9qVsH/pQbg6lThze+k0MfAKK8lexF0gZ689Kn0nzI0Rk2ItqjsOjw5BlV9jfQSQkGd1ahxl
gA==
`protect end_protected
