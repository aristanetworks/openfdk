--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
m6ezz0n2ASmBQOB+Wep5qI6J71xYNCx37SZ1vhWOrGYz0e/2Y2/yPH7izluEVAT2z0bSKwP+XKWg
t7Gydbmy6hwFsMdAwMfh2hOyd1whNCYXZSrliiFIxOk26hRHXofwfmRionofjewGs6y7IObO4BpC
hDpyltOD4pD9yC+d7LgiNa3n3I8xUa6/Sc0cecr1NYJMWB7ZyLkK/rCcnGe4A16I49mLzN9TyrV2
reXm9+KromiJUNWD+2OK81QxMjxNHZUmeDzOe4jwmI/ahyklYv+0jIEdWOHJ0RWRQi1jiXTczOb0
uJx9KO01IFz6rGQFipAmJfNrN4KTaxsWL543Gw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="M/TgImOBcgFNZPWq6UvPnVdCyjpIHukTrI1MheuKxnU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
liYsDrt0xuFeHteZCec5xKdhMheDUAn2PhpyPg2soCPk4WXeRvxrjVN6YWw0IvCWQ031q90kp2HS
LYNx3xXqCkrIxbgGcBc34iTEcPmlqkrcNzY23Rzo+RhWYfQxBdR48WiRb7x4ZKJJyLES1H8C9XM2
bdTQUVaGe4hGXJiqBt6s2nCITmjlsNp/teaH+0U+WyxNeGpZdpZzorVl68N4gqusslvxyNifnI06
JaeRDOvZEMBg3BFDSXJizVtgK/J5OU1+drFXMX3LYP7GlHzzl34Sdtc59p76tXgJ/quoHlF5UtxM
gkp9MBR9ojfl07m5J/67Azx0TZX+popdxbqsWQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="nYlljZ9cOdyO7wdRdZJY3olhlrgcmVYUFenCLcUrvro="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19584)
`protect data_block
+cRSZtE0eN3rj+DnQ4DOOvWGv+f1LzCyxHVf9ngliPvmtzjbW2/YmacQGMfhxia2DLIaiNFEAyBn
Ux/X7q/e4oqPr/BWwQ3bOHCA2SPpcd8V6eCHKt+CgYevexLpnnbk6mariRvW6dlXUzab2flZuZPG
bMqkGhvuWHuIS56kCQVD+vB2aS4dgZmct4P1VldAdyBd2MdEJQPKM3b5OucPzt7NbrFqeBBuZaVQ
/CgnZsy5yGcKu9+1cPtdQcniiudIqtliUwzoEoyxmFUboOtXXBYHrHfZWVXrIgqDYAE3V9TpphgR
M4o+eEWUblQsEgOM94Ocxg/efyIMHumMkgdlWi9jEnvv0zSxg1VgkFXvBnfKInsUhLkkp22x77a4
pcreKQlgp18Wqj/mFs2n+JrIpD1VUckuWJQ1qa1R6IuSvuv0sqFZ7ryJ2vWbao4znFAsxz2tHybw
zJFzmt3ZBLLeooYGS8hRvPdW+Q1+lqR3wW1Jq9b6vYblmYEapLbiju2FQqnaenPcmD4WPoRRGZui
Kv5orRYB5b3GRadyA7im6WZWMAkArfCWKFdrAbTi7UJ/7/EGIFp4qZcpVDgOeDEcqp+rvv98p95n
9qPMTpCUyU+kuyMkrW1gtFCeIroLvRphlxoPuFWN7i82TaeTbpbJKVWsTnxnxNaP5b860Lx04PEL
KkP0Ore4GVKmK2niwSEcZDLb2SFLeRA5N6QEBM7v2/QM7LnD4OaDockvhVK4dWBts+wtDJ9PvvSt
vFycOId79pqZxmEBES1mKdZSR+oj0lwLHwCgxcGlT29NuMVO8VUVNUNXiJH4l/XFYyKvIZXyWV3L
kvt+VeYgC22UgXlXLM7fQa8oN2qMux7XbWZejVv1EXqNLVKhcDL6r7UdxQ6feVx+bywDPuckGdFb
5UebiaKDpGiwtbXdVEai5awxoCXgfPRz+CCm0Mg3tYTVavRjr5sUdsjl0ZKlv8qi2qmZNBmIh02z
EmE7DQphY51IHRXMZQ5dI+2JkB0gr3XQgKtemVFrtnnOdy50vYZJJhFX3FESp7sAcLz42+dWGm96
CBGwMtGaEW4/5XX1eEF7uRjg4fgempBHOGEECz3xc1nAEu28nTmEGemkOpDhMaxgn01tEqth1twc
/46R7U23QvB+Qz8PCCxrAWUIGvtfLurExyh4y8TR4AytA3mX4b79pcnabi9wKsbjsoAsagpk4zpP
7L4eCB6iKFw14lncyv7/KsscGDEasxf3X0fFoMwOgqvEBCchXc1ivZXZbgfJ/NMhf2/eQhZ5PT3H
c3maRreSMwOyOxwZFqipHj47qcBXC4qPXfbpdpxG1rci/2b+3ra7dThL1pUdV13iG4ttJ+0LVZNo
KDpu93DVDEtP1cTCFBrPO61lornWWffaHtfbCh4IzBsmLN+Ykdit24//kE59YQrzNir1eLbCMaj3
3X686heJDdUExJpRDx5zFtBxebOUbpENgsBU3lkSX6u+YZOEzscGF6Eh5dX5hTEyJAhRKIHDcPN8
3KxYPBkSWG8lyjSUEFCNCLQqrXutXCjtqEIIVEB12epBpELItQjBFwLRFsYGQuGq0oX9TXhw+MJr
Qv/DaLNimJqVyG+zWMKhKaDJFepMgmr6cV3XOGNusA/t0NUctbR7o332BcsB2coSnwHHRp85b0RC
L+2vxLHZMeKouM9AHGYf8jHaSe8f6WcbcUlvYvnRYnqxlEO+nwk/AvZaA4STUrq1iNB/Y+ij32Cc
rmqjp+1UsfjdZwf0S9W27+ZykvLlrapG+WmpBSTQTFrVg0YFREwIgSX9vua7LMnimTxNO67cvB42
H+V3pVb0rae9hdmYAArjAjljyuK4/JtjAGW5hly0vxmPAZtHzPyUdp+uNNZa8Booj75vwZqIPCwh
Leym1j40fAw9QDfW1r2dVHuJ8pmJAJ8FZ52O7+T1Bcfihnx+9Ym/zDQyg92mD38Jwjve1SuiNtpA
0GE4qigKxYhs0i8pJrl27pigi1TNd9mYVHtkDyfI0lPy+B6xbFgzak7DNgEaFF0Px0aNMAkQlb5L
DJC59kIihC73p+VTpOOPJEI4hfIPLaTYnD96P3Wj/2iCl5YyM7uDIQfWfUq8pfQqf43Tvj0a4A8n
9CFC6F3aWOrCFpyYY9oH2Yvft63ZK/bBb9JfegOewWgaTyqgapARhZufQn6aMEagSWvCBX2IagKs
UJC/7/xbMHSS5tsks62W3OTZnkgeaKiMtHPXCsRP+sQhkdyOuc+6hN6nP5Dy+GLVak6gUV/zWCfP
wvSVyhI8h64lgm1nlv5gwWIRJ75SOyYqNyceN2EzifJga1gPn5jKYosPBRm6EhgyHD5y8lswRQR+
tHwSu6ZT6pEZAf0AHsPrNGLPGYIBqJTRifaKj2ZoXuMX627QFEpymIeVnFjCFRyvbKRJ1Jua9Q0l
uXEy6jjwhlI267ZTm7lVlr/TZAaUAdtPEMtiDzQhDRFUavHMISCFQzF+5a/onl4hLshFbMCLP0WR
VARvgUfbk9LiOCNlrX5G3khRoZpFYmNkqTPoy8/d3Sv8ZY6WOLYT/pG39uXSEFOnAyR9phDYAtbt
gm3gf0VJAP744NACPBKDREKtW2hUzle9anCCHYRkAhYJshJxQufgSwPz11dRBSUtFRJkr4oZ5Dwh
Zml56pDOQjYEurDC5k5fDGf6usc5kJev+nFoFWu/iITFD5mptgQgMZeOjaV3G6d+UNqu9iNfkzIh
6ulvWVRx+u6ruFSppwqlFoxHLfrZQgNGo1xjXI31EGpcIpY6X0KgoEU+V7EBSmaieN2FAEmlndZi
I8RoyV40OdKabeGCFA56KYo7KslDViX2rbZBkRPD0NidlBxAbV3rIDAPyvDNL7c9951Ig/I4nqVQ
En8EOy+9WgP1U+XF0qC+Plk74cf1jUXWhb4FzUtP2WijhDrOU6Juwos9M6AP6qlZTFNrOsQtLYiP
YgtXaqmq9YM95Tzbz59YlVnyfOf7S/r3ccozq8gDq2FwAddBwPeNDLL2X6iVmTDr5BLKyrK4EPze
wVGhc9zRCCJXY/Pq8F9KSiuvoabK7wb7kclAvQnq9TChZbMqAcv2FX/TmtagIcg6ZowOCMpUbvcW
JOSc79A2BiixWWCtN93+T0lx3itEmPda+TFT23TS24DBC6FKNVBVIgEHTPjxKjGB3ZovRG4cuqO3
Y5HKJbyC85OZQem9lXvl1XLj9sADYWUEhG16jDHgBVcE6F45sc2Y5zwzM8hprYqhNrCe0goTDlM9
Qi6OHgGHsQFz00MXSjZjApKqxWUTqCHfQagONM6Da1y5ehtbKfMOxzIUdYPlo4o11/D/gCwoSuDZ
UJ4Sb7IjdupoNeWBMuo3Fp3a/haVitOW5ZlPYFxzAIXeP1Bg/4TYYOMkFpsK+9yDw6pNf1HJFPm8
qRDRpGPLYSUR8e1qwwiNBeVxYyPfz1dDzyQ4xjJwBmcpyAPNDCd+Lxu6tiAgaia8fG3kqaTaxCPH
4MkUegQJalkR19pgvy9i1E7Vyz8USX+/WAlufUpzTh1XLQ18eZ3EtX/3ldDYEbBFiVdTEJM5P1Hq
mqrqokcjq/M74RREVfh7fDney2+4ypYl6sJ5qwTXd0M0cL0EFqy0SIEoBEYRJTLp95tPZcWDMCfs
7M2C0FzvkTWAqkqOCvcLGDGP2AobdUyRLpekUP0Zr+x707zuMSQ5XpG5vT/l2kw/KdhcNN9u//AW
dYnOKuEm+80DJrFnHR0rPzDbeodKpaFenLNajuqDrfBZUIXdTpiEKzexr10gxlJhjjIZebXOzut+
hiBeyniPyDGgeY/5Ub8jUj56InJxQGB9q60g97FfFuNapSkrdoPfDI/tBM44BnMm4TqE9K1nyyZK
nKLVWUCDwwL2ZidMS+KuFBW38I85nf10IjbxjvK3ZccgRUR/MOoZ+VvdaHuiKdDaDszsKkOk/tCO
nsYXQJFBDaNangcCFXdgzu3j1uaGyiUNhVTwN9nCIeicoIlaFwCIPpR5cExZ2tM2a+xIOWHLqiyG
HHVLKlA/mfYQsGjpsbdVIeTZRxHgNx2ASmUjMxDhezLjMaKOe3ecT6YMXPAeOGWs21ySDJDdxDYB
y/vZmU1AKRZf24cwokRVkmf2K+MLVoxKz+78ZRM51HvrWmNu98c9E/7CWP+QxahRuwYzznrFjd2g
zq6y3A/IKlbSwo1e/y6ixppoJvZnP0beIfnGjnLBNN7u8UZOITPPNR5TXhl5isFYCqqlsBJjaxzQ
K1hQtHEkzxc0ODDb3XVIS9eS8S1EePm/bbVyPF4doJKFMATc/r+wd7GQGw78d4bYz6X4bRZ25zRC
k6ydJaEfJNrkspD6KWy6M6Xc5VrSSIw9DgfMtJyOpIgz8Gp5EsAFvAL80aVB9Jwr6jP3iTuTZUX3
OImFSjttvxIpSPBpZFgsHdPw/YmUxcOUPKDfYS5wMO1cJspGAKunzShdIKzG8ylzl6SezUSm4SKf
1ZlyxtNsMv1/n4iobTngN/DhV8HRbtuKf+CiUlqF46CJpOizat0RwnRmVshxZTz67O3Ht/AU+0RP
cd5JhfX6Y3xmBWyg8WbhN8iQc8sx52+tkxO2Cva8xcYSj8Lpsuzhvn2tsThxi6w5jMtzn3opPSex
HBkLqdyY0iW+jIOTJ+vBL8T/d4Gg71gDmMZcfFnpiMNjlpP4KMxn4SIIunMD/tFl6mBnoAaDPpkd
klH10ypocxsJji4NGfnGYnfz1bFFS9qbE/hF5phM9D8YxIAj/hd4wQoeMg5545/lWr95fKiXzD7x
EPc73HmlgXv/N0H7vnMaVgBHg2UUHAAupxzTBJ2rr5yGKhZz+E+IJcpE15tw/3A1P/MnsJIcT/pc
T3hC2d7f4qMo09p1R3V1kSp+7SSjcud5MwTvg72uzmHu/u0tlVAyzXRJk82KVt11deWK5GMMe7Cf
xJg85bF3tMdFUYDAEjVStpfmJHZzaDtxSrTVpQwl7EW346p1K57IfYb1tMGVN2TZ2EEAl3TznTZ5
lG3DZZl6ib+b2D9dzyS6V4gSrq9CGZnPoCPafGr43c0MXiu73iBcXLXxDrn4cVzj3UzgCOWF28VU
ymIhsehRlr5mg+aj2yQOjbeOQduyih+NIW7YoUbBekCbbzeN/Fx3edUP6h6UoLrJVcD7IlRnavik
REyZU1AxBZnw8yjtGVxfTJNhs1RxsEa/TaXRttiM2m97x6cDZAlo0kPEZEEIkESr5Rvm271Z4Pt/
5/6kKu5GiXCKSw1ahxs6YOpFAbLRRvVcdlZM3LEwbQAlJaOgmMuoQHCCsc4CZ/0nRmZIxYSI7RmD
EcACaPrUMABfZpVIDO6yVxs+H9I8FeXG7dsfhoRuvRwDycyRjg/LQE8T1IJk9KG8p5AMQ++lV1CI
BwYDQZldLfBFKJsoNuBeh7EW2L6NosBzwLdW0hUy2jStUhv0BD/Z0mxUL86GqUm2w56T8Qxkn+4b
wgPvZBoGSxfH6e45xOglema3IOilKkUBmPkA5t1FUiTvrbXc6HuZ/TRBx7fhq3czUWSGhiZelii3
/NZz4xYBsZAV9vQRQA1736pzWGTOIY28cdB3wGai7JW1VvlEPCx/fdU08nU2wpa5jWvarR3u2LG5
3eUppj4m13e03AqpyxdqxIv4CpxxW30L8GU/xhwFvVvAa2C1w9ACH5WvKTVaRtCbMs7SlhVzVzw4
xnjAsjv8G7SRAkkQOcwWhSm2RKuzlbmxFxpJT4F2Ybwa4pt3iAYRn4hJh/s/cRaLT8HakNqByqO/
oHI/Lcv8LUNSjFunhhK3gg+2WvA1zBgSo6+0trRdk+vbVstKkru+DXTaw3sCyRKB8FMM1F6YMv8E
iiuut8kBUPQ9/amTq00oqb95CpR8jQlLzCmH+vqy1UDq38ms+bD9JT1+atEO4+sCCQHmFOHfGmTd
wCKbvyhBQkQnTlLAYM0Bi6PWJEEQ8RRhu6lb0vt21tU4EwVgDWERV8KGs79wZ6qBpKrNWvFjTbuq
a9G+FUj4dnoQRBXcO5wqZvds78sKAV5t3KKwCQeknSbGyj4VBnP2uMW2x7L4tbE8HFUq+NegWneI
jew0+a6eOFuBZRuUDHAWEdreKL8ScvyKnsziX1iCaFlUHwGl5Mzouuz52/A8B5QC6wBKsQQyFQfE
XO/KiOprw80fV/cug/KtIUKgbJ+nHw5DU+KccsouB3zo454hDeUx6ZHTT9S0bjuIxqYOp20iVR4R
bFXpB/yE6IlEDq0IuC+THYNlsAhnkyDC8HzDwLVXGYdimyv2dPJl1VzRummAXokXFmaR64PS3rn4
2kPI02LQQhGhzsuD+STgKSGjEtZqIHTACOt6pF5d1iBKY1SARXItZ0nF3iYya4uPOzzKNbACH6Ac
eepDhxUi9RuZdHb2BXHDKgVCUui0PRhpaLQ0y7g6V2bvzeJGkfsbpHwXQNSO7BAu63orK8U1570l
j10/ag3TRT5k57z+uRfGPEnv20o1tzW0So3TA40GIiyYuhd4w8B6siikCn/uz/eLdi4g6JSNIekS
YyhKniz3hvnF0T4vqpXc4tfH+D/pYAlkhuVab+tpi+KWcIpfr344N59qv4PkSXkYgj0I1MaluSmB
mPHXJogz/3ToCGVetTHehcP7182eOb/tau0k/lcUcJvNNsI/htkG1tD2+JKs1b7g1duIqj06jqlb
8mz9JulY7Pnqc8nLGCmHOw4oKccWMXR/prktV7g6gM5hoV/YKIUmRa6QFDoavs6nsF/6LvBcKVdU
LHJoyfprlALcUx9/91TdRjy5kvyJ6iw0cB0Ir9Hx1ZbHHzRumd/I3ffZHSavlX8qImcjHp87A092
CYpTgOqvLflGkWU6G+Tjxqe4ks4gMftKtUpy68padKvNGfZ7ymJw1cUxUp1PpXbXCWQW40a7B292
96UBUMZ09SOknXXoTcttfCqfnYt+ISqQDgZxf+sjl05u8vaUbQVdK7JCpk28VdL5IaxZfj6c179W
kzYM/ghJbG0W9/5oNNpQdMRviLTF7mjd9y+oiFM72of9eFG+5OgzLCMk/QkfL8eLLElEq3iAkDal
4jc8FjFmgRV79MHoSrf6WG7qm7O2ifppG3BiWlWuFHfhGAumf5P7ufUqETqIYz7qBLxdERlXWrJ7
cjVFj9CUU/tWm8LcgjJhz/6lVTtd/NdoDBBdw2mTYns2M/oIK5e6IJaZjDKGNBjKYQLnWEuXP5Dy
zNufd/Qs194VqlUTqT4OLF2IWCLJi0MZp+2BcPBEXn26prh4zxDV+L83igL5bSmxntnwMJb0PLmP
2yBuyHk8pi+ioMPLAU5hfDpzZvXBq33XcnWMyYbK9SweiYNxPbUz9RJmJJfXbX/IVhRkVbgLwzQi
YSYoAKlp7Lt4DK97CgHvDeEix2G9HZL/Zp5I+PrYSq7rOgJIJHYbGKBHQfzwgNMb0VHHUaq1v6IC
rMQsmHDZKXMILyfMr1CK3AeB6IaMWXoc1rZvxlKR2/knd/SOgM8C1iakdGRf7qpHaLZ3pTXpSb1J
oaQ88leXghwBHoflRYyMaBxJbH4z7qEeg9F1zdgM0lXqUJecD6HJCDUvZxu9sA3MrqSOQFA+amSs
MOpQfkt3/NKjBx50AuH8fc82J2Y0U3l2oMHpYEQuCL2mU1V/UQWGtBkzvcV1jGZ0vQExIJJUUvkV
2I48u48VaAanKvjGi5ylQzsni4qL/sedLkCnQG4TLCB0k4ttYeVkwEQ9+BWZDgZvL764Ci8BKhoa
sCkpC7LjWoUZQHQQu1jhF/Eqa3SiHmT64pQbES98Mktc2dcvqZlKK7q18fH1+KaLy935ORymHRui
AlIliLyAaiDKmTRqo2SfUzcy8W3jaqagxW7bK0JQaC+nC8W8gENXwEUmOg9rwHnm+mGww+sLaBxf
vUOQpiMaZu7i3CyPA10Xd/oL3xX7AneSpPiCgrxwrPYCPtHD57ksIpCKGDZZH1vNIYY/ZT6zzyAE
pfN4Qsccelm7nnlqAMvjv38l1LHcare8IgWvUaYm55kRKKcM2LTgpxk398TFZZzmaGly7SD0sR7k
/WT+fhI52vMAXMYatAVH0LGOzpAkk+aHnNcPuW6Zkc/PgjmmpkDFEd7P7Xcxz6FY58vpMzqU0fr/
AMrOi1kXKuqFPPtNxUNt3OSwhBgg1bJy1ICGmmnlQzC8M28QNMcIkwEM39kANN6lOkVs/jRb0CoD
rmtiTFXOOrtlsM/OECYM8g7guzXxOv/8DOWeL1raqccXhC1OEU8GWt71p93H6C2n1qhH+dOXjOjN
5XMmqQ2J01/G+1UsZqMkm4GH3/ydUU+dU9Fjypdw2O/QLmAkHZgZJ5S01XBL00MLYtOfcgQ38JUr
vnViymmSqtzlUsfHcRXpxXuCpIa2EoIbRrbFV3dRNYZhvS93xl9z+QWB+zzsLsy+kzG5Z1n0Rky7
H7Rj7L2cCyYheUitPbavVN0rNb0O19EV0fZJ5OuJS0rvi03061V8dLoZL92LkyAowa9inxH0v1oj
MRor2M9YeF2OmslMFDm1w2B1w1vPvAajsXmdKHJoceMLPu9Rzjfp+VRL/15KtuFutw9zM61650TM
q04UOqMslvRb/3DlukoBdOzURVCFPghNgQEjinKcIr9sO/OsmRcIPHi0ZVdFSElCL4ioJQNf8agc
9V0s0Ut2ZZpILR2pCBOmsQjOAamXSVLEULpHOjLzusdTBesmXvYOnc34OABu2mZF5wKNCvycXtB8
ZcO4O0WMKUeDSnigYLAeFhXwpsD39UZ/7HML7Ej4CeC6hRVQ6Fy6wbZkJWSDa0jUDpoDk/FC9Boz
fUOM8lu8Xd4T5aizLKJJzFV7Cx6jQKkme9ITQ+NuNY/I5+oM+f0q1r3HEwUQN8Be2SBhFfgkevyI
IXXT0mC7l4LaR4DEl5XO90Lh6CAGnkIeK5bsDOL7GBC6Kz1A6+1JYefAYLwqXGXGWlrUz11AgnWM
be7qA2XcJgs6GLyHxwAZoMR9mUlPt8p5u7r4CJiUK0mD2mmF7qVl8YUBCnCT7sl2DlLvT8oExZU5
eoIFd+F+fDLvlNbShZyjs2MuTsbALzRpCwlq8apDaPNoaT8D9+TPx1LaxnjitmqowA2HZCgq0eWE
xt5y4xyLWRXevE+6xK3Vmv+qYar4vrF6gvlChJMXC0i962/05Yj1RxlIdwiiiBW6w1oH7mT94G/5
8OjiaSZN5mjcZgtuKVWmwmEo9ulvbjnZXQ9ISbfNe6YZGikf8O/n3plsW1tvV0JtmQsdb2yAtgD9
GIw/lDQpntyJE9knP9ft1/60s7sGG8hPTBFpJNj9/EWlIerIBYZXDx/3+l1C3Ay3zexAgBIJi/0M
u597mG6SM12UEVvw8tgVBkot2K1PbhSP4QqUDKGX+jUCbKwYJ7rSQorRr9XrqMvqFGk0wTQkLV2B
mrbfVaa/tpj1l3q5/IrjpvC/Nus+DbXd5+qqCLLtqbrjTSgAnc8KCNnqMUhDCjV6Xq0+7mSpjTaU
Gkx8Y/NuQQLDt2xy+vWiIRAcXd6D0hIpNKV770t/DBtcbN+8kx7tZXDb6QZyAdpfMPj0LAGMACYZ
3uGcwddQKoBe5plIn30zk1OSDpgXssvn48JMyXTNbG9PKHMYDkzbpZyHSmc/oMDLPKN27o4safR8
YVyYWY5FdMhq9RW9XHbxoQukAx9rl6WIsp+PiHRf2FP1a4oxRlNbeUmv5Nmo6pnVm1dWxO1fOUqH
M7ej0vpCyAxzftIE71tG/GjIq/Mp0zlUNpOJhzBkg5ABm6GGVSt/G1HneT7dsXpEaQOe168QtIY3
aflY7jgClULgp7tYGBjfyXXPQsRmFqWMe105P5esRs+XrMStwaSu9dCKCx6rkiEYUW5c0059mVP3
rhLAhSyLLLqnBBbMGBvAInHY1xCCBEfmMRRZR3ZdvqIUgX0VvWYyA9p0WAxfWuYm6gObgvdKdn/N
SmJj4hCmoZcPjAqFDcmqFgeMlkcKZ+OibEh6RMQjK8VfdwqbPdwX95iafQn4xBKELc3d8gDqaPGv
1dhdM6ZWFMlOpoagsg5R9tXQfPWb6kbVhIu20liWqtjQD+mCp0vnXBkPEQuDEIqFgkPcOPcaybx6
wxZko23x9XynL8ELYiB1pIndVu5jAIvfZ8kvOPLo5Gck9hf4ptjeR15ZXx5QQA5TiZkSR0OTweFc
HtBe7SkZZKv18pqDeRKPvrDV+5/ilUdZEWmNg9uvmPlvtSXnjPnp7FizKqo63tlnjHrOfIWDsGfR
0lB0WhI0EwUgjFqAFLFUe136YnPPXOWd+m/CtII0u2uSija/RQttMocfYtRxbOdfr0WK/ExmHEYI
JrqKzM8/IKtRnbuOa/qoG/oa9pFLj6E3xU04FXxdvPQBy1kKgY4+8PvkRge6Stz0InhJcmnAIdPc
+WuWZADvq8Fg/zIOCdkjGXpxugNkEQTZ0PXcriaLUw2RBDlL8vQq1ZGxswg4nT4aDiXy48SF9t9S
rwK4E8oM8MfMzv3oU+d1JpNb13zguQgsVgntHgNa3xolvuCbtnf0qWZ5uONZUs53sPx/Ixxy5AIw
YLlyAjQpEkhfNhH71bFLuptkPfsJYWJP51VvnBLWyzemSC9pc5XpjZs0axROVlFLZcMGToxB1RKJ
g56ag8gFz9Zo000O/hnusXbpFhK/ScTelcbJmo3R9lAOYdWzKFqWAH+010+CkVALeAyNOaXTngjp
yduqogHRdF4EfO259bM+XfV/94CKaZIMYuFxNbSvUJEpj868DEkomnAlrbb3yYYf4YfZzbVmkF9y
YLL5XdeWYJvVcXSraOnIJoKJxtLzZw+Uy/SAmNGRjN7xK2+3Z6/UPYihwwe2gsLpLI0rVW+G3SNl
2mV7ZhCHB2Bq2IlKJYUc32Q+S21Q8g/MMdx/VcDtZrk0l2gtVwc2DUHfYmzGO2WN4jaIcbBja0k/
QCtXqoG+X9BEe/jspVFfu5QkSg+ps4lxrh3dLk1+oCCNYtm/h/6pM7/bFBCLHNcrWOunXwowKE1T
1oDKbJHSycJh9eLShM2PYJx7+qzzp+cOM+ARiNYEQlSb6eWdv7rtlh/LS5OSOJpvsLY05cymsf3+
pmouu4ZuVQYvMvac6uSpKaM5Euip4Co76wRwlp391ojNZYR2GQRrFc1AtQctzebE4aTbwkfnStkn
zbSuHoK9gud1uLbu9W/j9hJTAT1H8enFJU21g3fMg3jwMYhKzx68NlOEgr5V+h+s3MsB/X2qb2Z2
Y8GAE1+TPE6e1TdgCYogGLjBq6GoBXWEZvVKlaWmZWjUJ1CDE5dWuwIwHVoP7KGyshRZDPOuWMuT
rdBHKw8V1GBNV1t+eAvSIXZd21yr4Upfp2/916h6SI4lerQ+6rfVD4hEwJeKwJlt0QoQSCi8lDfL
g1ciC3dp+39WY91EedJupKQcVW22twH389M0bOlyW72lyOY+lYZ0aBFWJtDZGT0Bjy/UP4Lw86eO
4Ggo1+OehY1ia7AL5VpR8CHXiFn2AunDe0qgJEiryGbXy8oE923O4/Po8uKqPLhwsE8x1yQae9uI
/GPegrpbIB3R63AlCCKYWnBcOs1OgDtHklYSvw1rVORrnuFxJD7WIfF1ysQaRoxO+xTWZtaiCpr/
+wpUbgLEfmskJfT181Ye3Top6rYAssJVQFuYNLZ4D9ZAQw5o0QNpogCCkFQpmi0gGVW3sBQJCXmW
H9oaR38hmjDB5HwsuTGztaR8yrnWDDNgU+0Mw7TQ2Nsun/Md/2CpL8QuHV4Jdx4gwwukLd85Y9D3
9kOV7j3NCQRuK7axaMun/Yu/74zNCO4kVvVJgimH82w+NLorRV1fJURqirbywST9KnVXYxtKU5/E
HBSiC/j2z0sHYwd+MTIUzhbP9nNFEudZeNSstYMVdG0EaNzb9X9ohh5y6j03h7KuB55bxpR5RQgW
5wWAUROFsJpex64GrJeWWADhMd+OqfSJTRHlr95EIMxSlXaZe94EKrbuJPA1zeff2XhAwOk9dZ8L
oIdpLeKF7Qb1G6rcMiTZE04/K9Uoza76Itf7iU1GwjqB0ODdnu6rByW0ls246BndZrxTiaky1xAJ
YvamJVULN4jOzx66+GA8GL9vsYZtXhXkKnr82JU/0MYQz5GGXsS0cWVVW7qVxfhPGEgjHvFqsLXv
fCMelKRncsfnv+A+iIuQkkrUTixotVDLZcdP0v9dj60n5wRZJJDXxxMf4beKsV9oZzN/AyT0PLlB
3RAKqEzd/yut1hBejoLAaNDnFQzmqFa1tid+fzAolpYoQqk1oRsrjhYGjKpBJcEP4zQf/cbblm40
CdHANh6F75FJ9yI0AdTgUoxff3WFZ+UFfIrvAXJSxXktXoBHtQlVAqeWeyBUnonmyWPGsXTWR/r3
4FFy8hAQYx6x6hOJjbJkhUp8JtL3RpCKAhnu8RB4h8Yv+LxZnSqaoLpLrRppfibgSDq1oLQUHEHC
4rf8sl/zn751Xlgt6qca6BNjHybISIBxuVqHSDLQ6MwA2hPV7nh0p7e8XexxezhuG4D5dR7FVpDo
2ZaPWqTpbYOIGPm6nlDdFistuHemtutVNWxIjG2g5KtPW3AX6ppFWt77jq0p7m2JIzGn6krddHt4
29JCH1JndEbcrIPdULwtW4KT0XfinKv5+nnNZfP+9mwpMxcYIG5a9c7KKZn03XfN503ya8KaKHGu
BLLcTMjya6PojtornHi0/dKyV8XyDNcjjJdddxqi9J0vx+aBF1oS6ydHS+mal0vDV3TOTqsPvCV6
oHfXu2ur075lKqPAffCnKm8INgKzfS8dVMzKg+tkkZkDlnWrnugNqcN9j9AY2qVQI8MW39yIKxf3
8y9qZYT2L1k545FZvbEns99EachXDY7Hi7LiJSMRq67rd7Wy22KF9jum3q5pEWR13Hs/LFCgC7r7
peGvmHg/yC4KgmrHcQBAwbQi6iN43HEJSYYfB0Hia7ZjW623al30C7r5uXt1PeXMMEyN8aA8n8lC
A9HHCGStr/ayFDyXfOLxGB7rsCNK2+8RQf8j/3lqQE0V+jaZ+XDwdo5SJU3pVs8/YoliAXmdbTBJ
bdUHKh0+bKbZyKfO0gaCZ09pVnlf+sCtHG42kKue1JuVQg+Jf78b8pP5Q2QHkB8pVWirzccUcFjQ
DowbxJJXC/KI5JIRwojuIeRpyuNTvii3ez2CnBsfBzQLML74pwrHWRelFIFM1zIVbosvDELgzJVM
qA93MNBPU1USZjM6cQ+sTb93qfW+IQgN6S6gZWnJWu7N+FTT4xmgB45mvNjEW7rmDmayfpnYaOd/
k6+Wf23eQz6f6WyCotCYvtXnhtRN0r+U34lI/J7HmQHxak32dBpmR4P8Mra6JFuNEY6ox6lEkTw8
V8ERxzc1WSJocqWDCsn1pxzaDKg2acd6uCCFL2tHOAtkoEiUs32C+ukVGYUkuIQJuVst38wNw5M0
wRr5gOtKTBUmQRecUXfyZ3urH6XunnMD5nS7W5pBusQZHNTVSn0TKC5jN8jIrsbACxRy7SoHHqnx
w+8n1XKhcb4TDJMbkoNtUGFQMswdLTC4aXMBsACjWUd5boqTbxbQEJkVmt339ggnw38+YepeKDMf
+JEpLQlzUaGna366J/iJxK2kXJ8VwtzfEwXsxNtKU4jzZeEZ8m4GO59m+q0TxYwpurAiFVTwbpCQ
jYmQ0SxkU6BxGJnW3bNPoS4XIAjR27d/Fi0jYxYK6/OhORZ5+kdSguz6/jXpOyrZ45T3N1TJO8Kx
V+X/+51hjTIxtfBqdPhJjE4BN2/KFw3rLA2DRNPNrpHGmZMOmqNcORdQf4l+pie7UfTmZAAeqklt
LkArWYaeBTESvpgJcAcp+3B2BOs+3xpSHvXy5MvxS/gJ+a4crz3L7bt4VzY3k2PPMQuHwmdF2y7R
j26kNN05sd7jRKfU4FqkvJWzJu+H4JRP39KkYt2Kvrn0TpFqk/HhhHXm7WmXVNrbeGHdN6ieqjO3
lhbDg4TuLPcysROpfRKeiDKs19/TLq2c2iz8LAnOTNngj4doKZmQBrnT7U3Uq15E3r0fG86SR7AC
uHpHdgqc7ZsemseNByeiRXQr+J425uuKA4BoxPiAp/gRZyh4K1fGY7Ekrd1q3pAR8Ly8+3Ggsnls
VvIR9OOB40Tso04K8DICx473IbphPu+vhNKKwffs908mVZNOJxUbd+o0tMpkEyoZxg7IDGmlCZqo
0J64168xl4I83LyVCtlINCgKAvmsHkUfETLVWnBbOfB+aKtZUDBuQPF0bl+1J8pmiX7N9M6TBDl2
Bu+m4zoUHIBmyr2yaZUBBFRMc6ETXPcqT+26HSIdjdXOmBAXOXylyjpTyBvm6pv55ilsjqw7Gd+n
DFLDl5EEffXii97YtO0dkJOPmFlhvcKAgsHWGb5YwYGrVxbCaS48hrH/ck2c2/5ObyW1+lGB8sbZ
MfPWI1bLalgFTfzp/z/bxzx+pbYtRfBJDUp2W/omw5nbS4nOP63ayaXh1J5kqK2BuxxoFgDrW2Gc
INGOOuJzLimZEtfdVmTyaCx1JCf3omNpHiG0g9isRwqZw8NCjkn0ohgNBpiXcNI9faAzpROpGtsL
WKDTVUQ7sr7fbHCQ1TXb1QGH3/cwQJu15D+bQc+4ux6fFQnmZDZ40UzfxsOHT5yzXGZwJ/RvxXRS
GUwheEN0w/m+UB7YeVGBf+umPO+GKnTlCcW+CuynUrwXFM+ILauswCKy8ryFrFn5aUBD4ZCuz8Uf
8CfEWvTS9oRNpDRi4PDVbGTdk5CZglJY1FXEhFIBWcDtsvxd00HNoaDgH9HBe9597pEhYVXINrAh
7sogUtYzA5wdMgjbZSTo2vrGX5mo2douauSph2hbz6LcQSIlZyZ/JUBjJ++sjR+CFu1wvIl7Rzko
tbxN8Vmh9TgnVxOj4xlRYvDWY3Jhkw8SivhYpf5GhIfY7lGNdm3fWGkLbdClxwHt2zZKmgCr1T7G
ak8LM9EtCO11tHP2KgUSQIEAQ1h6YoWP3V6lmckpDjV1ZBqQ7EcH/OeVyfgXmeNZKkTloAw01A6s
Y0RHZKchIq7j8TTafBSy5dWYvu8pAdlRxmSXiMDcgnbzjBCTDjX/lY5son3fyq3Sep8I0sPff8pt
G0P8aJdadsXJ6bcP3Q91DUpGAH6J/whVRQG93W3sZgLV9JDkctpz25m1ySKWtXqbeDS8AOczgPA0
fXdfN3P+kJXxFgxW8wfhMjRQLgbA4jh2YVpTqZUbGsr4stVwy8VVLvQZky7a120VYHctrEhCPddK
kywO98wiHWOq0kcAG30aASIROasLu2p/ri30fpy6k14ZogxfAdTjuw576kvlleI5g/TaYAJcBnc/
+AljQ/AaA/nuR4td7N/zvb6P1FMSgxS6Q2ID1UajqFekc+klhXlqVM4KyoDb/4Is5ouaFld4zvgn
P7SwR9jz4aT/escwuQNm1A5s6zUFQQTrw+PEEloEgLCGhqoTmPT27FjQZ6D6hog2+WBDbKDq7eg7
NKp7YUcE/bgTRUqqtbTcIzTzQzZaB9tdgJI06+QG07rsPWihMiHM3ywgQgEVd2XtkdUvXLs5WLyq
t268D/W1y5b5uN+UeE88170CpD+7c8Y3hLCt+9l3B7dhaJLTPZB2B+T8+9BJKv1sFrG9/9RmpIin
DH67+lv4nKR4vzm935WJPYl1NjK6m8B7qYODsrWsZwwGtciilbgkBjnDAmkD1+mOGVwBcOghMhui
MXQRsSB+2fRrjzMwdX8v8u8LxMM7lf/Zc4FP8M2xgteKiNxGqk6N3U0NAXerWEtfcwt9hNoKqX+F
Oa0dLAFHikPOEkWCH+hqjSqyrZCsTpX2hPC3r2EZUpGMqI1QbboFbCgpqZF/ZCrS4iTpoovtz75y
UqEWv2BGCJ0QNKw9sMuAfVcBE+hmPT/BKOiwsGepUWFIHTpaowNpl3BOQe3hhIQut5Dns3zB912/
+b8t3cWzhk3Yy4Lrs4nijPm8SGrZeKjS5yMSkUciyHGHX9kYXoAZq+ouB4eUjvYJrinoOvr7mex2
rdy4LyDBt3VODoNOFPSlzwVrNFcXsKf+Zjnuv3nEDapdmDGNHlsnxgmflAUN0giHmTbRYKxOtYSn
i5U7kbp89zR2raL1sZFHh2NhhQci2AL3APqA79PKQyqu62e0xH7oUymYz/zBjGacdsGIKWOSkhhO
lZ8Vc3D4uves1OybfnMsP4Qa2i8RtLALTFzZdJcwltKXCZjj0TkOsp9/JvwHEmrEUVdYRAqU70h4
4VMkiIrtd+DWQQk8OZnw1Drbgqh/a9l+mgl6bVZLNtfufEIGjQDh+Fn7G+V1+tWmhkRDwu6EjvBs
n9RJLE69HGXWTWqwokWJxJ8g4Yt+7wti2bCOq/4wIkPFn6A2gh0l1qpMYFh9j/OWa4AxzAhXCUOF
NnVZJSRvFxnsI16OQ7Kyw8wfirWONzK6CNINz5H8X77EqXhNNxvRlTHjObiZHAqDmUsy7gYdf9a1
ZHYAaY/G4ZD8VEPUwtJ2mHiLGCq9zMivPFJzzuyfaOTeM7EBr+izIGzdo25GwLSCAuiFO17Ij0Vj
n6YOaV817f6/NUbVpIN7WFIQpV/j4W06I/YoJvOKpqjvnCgSNH9i+yUvlt3ZeCtMx58ttekSbc4i
5l/IPceQvi280P/gC8v7+io4KZrjpSdczVHHXDAJeHUpu9mDvIl4hecohrkfJmn/cm/tlnXkvBi8
8PZLt48vHgrby3kQ7QsBY+LQkJrHZ3bdDKVSUuI+6Ikpirul+O5k7Wj/vUHyMPEWvlhaGWKMUdAF
HuBQBuOsHL5xwj4/BFfSI7BUUjjU24AgoZ+2CmthUjcj5qPC4I9FClGwjzIP5bGnvH5cZelsBGYk
xwYtyVXYSJlRfpMwvCqo1CVTvPVP8MtPmTnnxZOYFQGUC4fYck7f36QSzIXWWoOllUwQ/+F8XmND
cP0MTXAuFMhx/8RujdOM2FZOGMRa/x7vUhfJZoNcPvUHIfjpF1dtLSyWpP/VJ7dAzPRr8T77B1qj
x8WuNUzZLjjaUYVQrBxGk38PqTZR9rPFX3zXbBfnaMEsYidtOhDvNtV9vIC983VVgPZHtdpKKjXN
hnvG5uzrb391ppkc0Ea8aXYA4kl/RoadeuOVIC6mYJl+IQQTD0UILYtDgdYq9ebWNrm2QlLpm+zP
uuDs+jvojH+APyLmjt7ZPbp7lOLcfKT4WdZmbsCvDP6TPc/OMKi4Bo/+oqr0ucLyarvbzM8i4Hqd
faVYPWuHeMR8dZ36Iar1birE2LabbZB+9Gcw8TJzN79zOvMZ3va4tv4Od+8nwziNFPNFVjimTp6I
mJxoRDSuld/3H8myrWbL9qBMvrmBPazJpNvaX/6vwn1SIeb1jS7piqLQDO/sBOs0LjQKR9l4U8U9
O7PhwmhW4WBKevnPuLS4hqbfzdyfQBDrbIytWC6IypYDz+GvwK+1GA00p1A3FFi258n2EFQlJiCo
s60vHw5AxZoaH9Dnc7HjxCgmxRmBVD5/D3/8/Ad/qFFLLA5oQklqpvOGoaAwx9xDyAxvS9DRMhUo
Amo6+dWEfmf3Y2FM7qm+ZPfbaB/6DU8vwunJMVuO56E448Aa6pJgvYOS//UnGgohNt2zZTOF4199
n+poxyTKnh0L8hBHMB0D92xTxk5W1TeyXU0kZ5uYTJlT5F031mIAcr2Kau991wbm124ugSsXwmtK
B1X85vc8AFEJ32OoQ65EuWSUwdxOa8Xh3kNKPVI53p7qxY+R3Vdtb4AoCODLvdMa8q2H2pjHOmkO
5sz3cWMhNocfcBF32XSpoNxHh3Z6fn7ZRxWwMUaAGBtBPucnQe+8N4HBKdLQyvqWKpXaAE3ylDc2
+bZR/jcYylDf0sAHsaSa+dgfLPoreqyT7BAJtIwbGeSAwTL3/Tn7ps+v63s+U4f/HtU4LCcPwEf6
EB1Pv6lXnXZB20OWq7Qu5AFeZcYp5gqGFZ1u/GMtdvY5aMJLSRI5KwQ5OljyZ8LB6uXXBiF8KnLx
XzAwWzcxifQ06QtHHOEKt0Z8B4fGf5oo25cwkuCQd/XmGcu2o6fqqtjsAsOfx4TeBZRgf7h99VwJ
B3K6eu4Oq4t/hKrRxD/16DqvF4JhEMoPTF8hBvZYUZ+I2gkD1mQyOVQYXBtMWgGgvazjLqT/cCQs
GtZmqWmH7DL3R0gPlDg4f7nlCbQGXz9f14M+2aj8NQ+snih106/kXZBZOGGub+HPG94ntEs5+zbS
k7c32QLnCoCpQvARPHq2vbPF3Eyxm/XcPDJnRkObg9C02zmXKJEYvinjsZXyHMAn6oI6o+9/HH3r
Gv/QISRFL9L99r7qpqaRPklHsh3Tmef+GwLxGP79JXaevLwouP9fRfvQ4g7+HcDzemO0NigZAQzA
MA+Tl/ZeDgPW5E+nxs+Ppm7rUzCuxSvpaOLHyc5NFGxYFaiPl0sTwdNtjrPYTSr62oGcBhMXbY3g
2lhkMkCyJ+i26RyPq23XsKPIzEN7DgbcPEiQtZ/+LznOsuVAuu/m7iIX0KiwxP7z+xW3OqJO19JY
uMOaEWZOT5WydYIKzRnlucwIEGVl3ZjcI7Fmy7f28Pi2ei8yM7s1s62PRyW2axy0+2jeKgTXAEi/
gvz7e/s0/KCXroTQa3NgJhR9SHYwiGxASh1cWqeECWI2Ap2tjdteysahHN98EUg0qPuSrWhhcOlQ
UNJFunKki3SGXv4YBYy7KsLAa/46o9DoHfKGp5FAzUIIwDHV4+XylGk4gZPm1peFY/+tePe3tdcs
gkzxm44TEqSFVO7usr4Yh543TbI6VZq6glLEst1jHwe5iIZhiFJcFLRSTzORukMfBA2pCRgdsrJO
pHTjc8kFBoFxIYoxQvzy3myTvyFQEGgsBKOXoQsRujRxA8ugTDDMJoBKAJmKNwHVxblhJc6TO4fM
6smIxWy7sE3MBVy/cB3BjEQlsxNm+ti2E2w5U1pqK8AkhqZWMrcPCpW8gKmaNdnnXfOQoieowt/M
uw0OIJPql/0bWPo7MgWjgbjcY/3t6VU2Al2NS3p6IdY5V+khzFna16VKYpqAxf9WoqnpK4pEBGMT
1ibUJiRzRr7H7+41H5kudkuvKTdDk8a3t3AidNZhjBRbLRrNSJPQe6gFUGz20B094UmFMtkKOERF
+JR9fCrfl0a8kc7lM6S+amkPG++sPbWzglmqVL6FyawCYRklTeq520EMkFEo2QiLMnj3Ju3hJcq9
B03rAz9US/cIfbPnRvDFWEHOkkJx5kMTZRlDvsJKp9L3aF6CWjUmcUL4FSCN2Nnqjzh8kKet2No7
7MBhlviYW0WpyZ0rAzwEoW4VeAPE+G8Tc/b1t790uG6QFRSnaoknasartkgG+udfbK2cEyi1HkWb
vneQ4jtHfvMw6uC8cnJhvhtFkzljOKeaFwNU0wXOlvKEyu3lgCxoTaBiU6uPMtUWsgdfojFYlpbU
pU4nfMdUnP2X/MC4Iz/c9obu5XVNLF4/RIh0zl79KWojqhPZECzCvLK37jp0ScVDLXF63efMaF3n
/hr0TJ4O/3SXEyG4cpntEEOLsVBgAXLSPxSU0fyobG6zJLmBAHenJFXobr9r564p0gruVEwuOCXs
YCUlZHN00bSxHZ/H/WtT5V7X1/k2HBx9lyNlNnCeGEv/bxwSovje72STCkb5PQsYHC+l1ngZ4SoC
bonASRp67nRZDfz87SVUdFDRrxvExwVh5Ro06b3D50VqKYXaRQ26yoKqttcQcitpfdByjAUaIMYu
pTHWLFbNvGZER/FulkMEXbdd2w6R2tVX7qm6Ue9IiL6x4+pNyR/xuuE5L34jRPWBi8ceUCaPjeu9
OdzntI9XcARSd+dpOpS2IhnQuNp83VdorqueyxU4L8424tZoc2FC/hyuXU/wfo6SXMeqiM/uyu5X
EnavrKZbIMKwbxPdOZjjNWt1HwiTh92ECqqhIIY8lq35otSTxP/HxJNYC1bJaQOxZQvE43yIGGi1
lEXyfa5O7gjYWtSvXwOaTs71Auseudy5HpBbHSPLzOXcrpDai12src0CFGQdrEPjDESvBWsXc5gA
0fWksbCRyIEP40iNOyY9tPDxB9EZ4owsY1qwJn68neLZ5ynkF2/6K+QSuE6gu997y0Gt4fdELmP0
r2lWN7lio9HPhCSATswe2agUD4p4gySmYkvH+SOW9vB8TdLiZvfEuqBUL1l83sjGtyev9kH2Tu57
l8DSuwZuh/sIduzcfDCakBJ9V0yoCJiXmF0qzNAp5hxNTRnrq01pM35ifdGLPR+czS4C5b0WmgSu
QIpwK/dTkej/gC7A0PiwFraEkQ1fa4AuYNEOC2Gfxy8iJW1DwZhkTm3fOXOSXbR3QlCxLsXBNBIu
OzgtKdHZipoRr+5yMGYtq2iwPGuQWzUCdb0kEg2FBmCQyvWehPBDoPV073HqYHo2mbzMBRsF61TP
fhgR24SbEL9nLTZDZ5pRxt1KeB0izpvBtlBH5smVc8iVVqW2zHxPlEvdnLnCpjDZcEIoJx+7v6mI
hPriODZF+jlN0Pu4GxgRBlMcWj6Mgm1KR4Gak0dvDrIROCHjmv0nTFHOtzOosgLvjI7YI/nu/mgk
+2haFDLifuX/Hy00zx8+w/m/NPWHWrKo1HeMN8jTUBIw4VF4wgEfZw7M1635oVxvPdkeYkpCv4ge
yQ7Wo4DHJqag/sBCFtBXlnkewBcmKXUMpLz6UxK9Fjo+bDZZbTmNBYdO1dQoD3Z+VeEbYLe6zpFd
Ais74O7W0HJ0610DfHD6JbZmPHxYl+xyyc4NmrfL9wNVhaCifCsAu/Oe1FKUMOPePUcC9xHXR+ov
BLd33qN1TXzczr5N1ZpQiVzV6b/nyFSo8v1O3crTOKvRv4RLbIkKvzqKPBesX0PGI0zdjx0Gsuc5
uImDojh0Y9WpXxX/IDigSx90YEnodVmDCXG/wRklihQmEMCkb/g8a25Rb056UedkKchC0PJjuExw
2ezF6NA9Uiks96JELm19MNTxQLv04mMRvZT2pZnUFD6buAjL69KjMgwWsLAwqbOLGcoXaAe2q9EO
8Cp4JFGAfjfdx8fQm+W0MfzuSKBMXoMkPYEbtWckcsvoKAiIuTogdfQJjQN9MCf3+TM7gRpIl9ui
GHQjbJwvOjgy03G39cW8EQzCCNYED1h28tZeIrqNF7aXONIYP9xQgYCtWYyM+UXnYSvpKVjihDLD
ExEMKF+KMZBlBXQuPOxViAWt9u/wEV9Q/D0m3xGkWMnemlKXWcIRvlmgevrnbYOxG7DS8HixKu8p
TqA87Jy7InniRV+jLcA6Zf4fpmGPFcHci3eWAkxhnMmzsSpTXFCpzr/zG8fVNJhwRGJ8LqYbxpAs
gGbjdypdm9m+z+m2YKGHHRNqlFdmTw0fCp3pR1wXNOMudu2mkB/Mu3+1negw62jPnfU9vh0nk1tD
UOn9LHB7VNCK9ACxmghXj2Xzr3QjUWvuqzqN28UdCKERmkHP0sk6MpooUjgtvbR79REgRAwBoSBT
SZV9Jd7rDMnxPD2DrTa+4iUUtvbvKVdP0yj1azFDVBMX/P21nw9E4rQeSJWuZHYPGbRO/0Vixu41
5drpnWpcN4BQNzlV2GebTaJLaiBIEoOjwXauetZYFTxUsIGRebt93I0E8OxawkIW40V5Mavdadxw
h3gMPlqcfEg8j9ioajWZQdN9G/wjX2mX2Ychh+iGGG3Hzaf9L/pHoqUwEm1Hs7HgKqGIdtnsKdN4
A6SUMaVrcBTn3/3I9Q3lrB/LpuXB383O0Csjz62AgLoeXyPJ8J6/M9n9C9dU4RoQZukwgiklIPgE
SjAnS5XIf5n7l0XY9EjybMm6k6YxjoCwsYl+UePEx4wRyd8Sm9YuBwC6Q41kZqMOPqdkixF3GVhD
FfNv4Awf9JpezvR5B5q1xRrK4Zd6pPfHkrckqOMN72f07WD8f0mSYKxyvBLDcmwkmrG57VI06YdN
9xWYqL+/tmdskwgdNfDdD8DgW0KYkw47YUcOC49gTKEmZCu8gE6bQoumavpkN3lhmZB+hHfb1f6X
yv7p5MQyCapQQrxSL9zmpLuJiGp5GjW8qzoBPu9TheslfRMFxB/djfx6Y6V0yJjcsANiKnLIzj8N
4+Fnh5DRJ4oAxChbwFMBDnvajQqoRmB7wD2665WdeDyu6IdfgRRoD00dUzo8foeDtQFx8Rg25MWD
IKQ4KqzyP01V8llj4H7rED1/rq7m892DlUwfx/yqKLmFb0ju66BIUPUFykXmTbNAsIwEDh7md+6P
PeM2I7btoi1PcIGbgQWu6v53t0rK9YW3vb2jhJw3zP2oPHxC7tTiPxSnM2JTJw8zVOZyoszmQAHI
UDar5kYztEN7sfrYJEO6KZKY8RFAvKh69gFvSVxHR9hTRKaeDJzNrhT8A0sRD2FTpY6kHnQDbx5m
Z+cVjurqaD5IxWCIrguAMdKh4SwXSPkAhinQd1Mguq1S4/4Usu9ZDsf7kGA+QygVWXoD/kf2xlBQ
lkAeU5+/egiyGgLzTb5WMUfyi/PwfOouNd7t1SWpKrYOQMz2mVtZYv8yA9jEahz4LSVc0PKz4xZ3
gKUBsmiq2yxqWsgxDJIt36rt8nvQr7yxColjrejneuFXGztOP7DtQ3/PmoOhyxxHpEXPbWU7dJ/T
fpVaZ10wI6dIDX8x0HVaVsoMCizRLkv1Pa2aVKp4vxkppK5K1Sb4vZB8zPQ4IHGUPVEl6LJ2jrNR
6aH+sPAnAKb6vfMOJQxnHGNXzo7F8vicZtosgW0Hy4hV98VBzM1K8cVF4vlPUt9lddk+sZx7tF1X
+W8BPq6cPCuUdsw+Dzq7f0RxqbgGB5lr7HgzeWeFkZX3oZeSvWFh8aFuzF4O+JkUee/Z/t4ejz7B
qSjrostTTofPgXSZrVuRMLYR0MouNAnkfQvgnlImF2hAMNpd4F/fe1hGlQlvNoLKf9pXiPOTndPr
m5O5Z9MfOCGIyacOBS163hPpXn8EKqMWEVIHOQqCgCxqfN5/7q7aEv1scBDwOj731BDZ0ucjzE0P
TaJzp8rqHo7wvMlN0kjRp1Arefg1xZPpE/aYq3xw/2vWTL9wpa31OEFmP0PlRBfTRPRSXUx8Ykzj
gt3VFfN9oAAfZAHM9duRKAt7H1H3+SxOOPdR2hC2yz3papNb+o9yy6bDZCUPNY6d3tcZwq8hCL05
bpFMQJBEgPXrlIzUXH2fFfFwTJk1K1iu139sUIHDPCCbVg8JXnWb9TaTA75O9/oiEeNVEd2BDYxq
skUbfY5ZP5Hgstk492BUyFmgh5aEeRct23kn1B80AfuRKosBn9dbvz7Y5cu7H+kgwnHvkuX76fkc
KmHChr8ak6ekf+aXZfdSEJzxkwedYId9YfX/2Ws7h8GeVg5TukQJU1kyx6g6GzvUmpzllEIZFcnn
+jf/YvitwEjR/ctOxaZoaqulJo34suheJHwYIz/8PvPYszGhqHsF/8tE3mz4RGgyve8ZmAyjMC+s
M6P4JdaBKw5aYoOdVk6H3PyhwKxjniJGSBg1bqKF4PrbbdWElChVPjQgyTcpWUI8xdEr8AmDUpwA
KXMDreZda46sC2yJWj6FLIc5qbY/Vkip6A4S5IPYEiGhuD9aMw/76CelqXu+pk8cDJlTS6mqv90Y
qRg6EKkeb1JH9mnfE5g4lLzuMoGGySbdp1pgRpYtWg5WBj0l953g9NueaK5C5vBaFaI9I57mqAhJ
ZaxBV/s8QFZLU6LHiRq8Vbslri49nBIAOpaLQAIlLVk2EcNRYty6pBVPdlSxnLqtVdWzgNKi2JZY
mKJGfeYbLZ4NlokdkEHpkEQTVEmGAn80nqPcQOtUOObxiXgQASd+eFDzyTFA62nxtn8vhBEP7tGy
LZLFb7kto5F3W2iZNh8jpmW897/9W6CWbg0nZl4W9qPg43ZUomjUbLjWOmp+YJup0vBMdHDRN/z0
zq8ED//iIxl27RPhkztevZSOcbhigoB8XPBpURU6Vm3NxIkRP5ewDFz5+MXuJSXzt6GI8AbL1zLl
L3ndwCDR+EyAQKF5uXbIrR63EV7rMGIlirNJglUbSGqxLBy68GZb0ic/iyo4LVfrR8nhnOx0fTOv
rXvHFqx0WJI7VM/tWY89XKUfP0PaAZqzcVghbyq4ERdc9N/17LVKLuegP+xyBzCr4s5G4DJDWNTS
i6qWVn0dnzmDWUk/o6/3pS2fmM8D78LUI6v51WHANR7burGcAa2P8yDSxU/tfOUXErqJuSHhwmX9
inbijXuyCBY0iHMWhG3n/NNppojOa0eIAjwOwu4YrFoMEddSSGNSPSuoNyfW8h3lMKQiJyQbSqmu
1BDWd3Twew55lSq24cZ+x6HLnTnsvVCEP/GllstN+Il6quCPR2lBR0gHOwRnhOSZZhiZ33FtB9XB
kEv/qiaf0WBcxsf1FxgBaC3vvz0sMeWSKFAEfibrOlroREygQVw5cbX+GbV/lFkJJuHlNaDZ0uVR
aqocmMgqq3IVI1W/WQE6MNsJGtujD0mrwKNeV38smy4wGY4VWr7F1rOz+kSuz0pTP6Jr75+FB/xX
b5oXisQ2X5dS1ZSIrV9FdncH3pZ2UH4cxDp0pwC4ZJPttLw1SN9MNKsfJrHRBKkaTNbAsUn8JqvV
fgxB+e+cr+IHaT7tDpLN/Qnh07eEp2G5GbF/bvA/Nknxo1AvPt9Npe7rYcyNCNdfHLF98zCIFlkA
nuaXOlu3SnlDMkSXNIxBuGxGx2dUlPVg5Na3YmlZOEFjvwkh28LQ44YjBqsz1lRQSo5uuyRZwVAa
JJMJ5Kj8npk1xHiyIavNB4FMUdG1q5yrj1SXGHJQlCIKlomU1exHG4FRVr9k4NjvUENYAHnNCiMY
Kgv7s1rdGM48DKO+rtsROa0wT+aL0x0PJQdyPiU9/v5G/elRFDKPvxtuy4027H1g6YQOPCj96F2L
WbKkayyFLynx3p5+Eiee8V/VjRpXKBAd21fNpWkdtdr4vbvmHquB7sI53hBMMiTNcw/Y7BZMqaSt
OylgORIzTUTk6Hge7MbVHNOwA0kWk0gJW6Biq9ZgX3jn45Ltru/i12vDcivogJcKDb+/2SplwADa
dYXIIf8mS8koU/FioNyCf+yGLBfp0Iu9rVrgwQ82apTiKOX71E/P9SR9uKq+9ZQMUTVYBCDaBFkY
zhFIHMZMa2BZdHEogvuU30tYNW1XPtAk71mIpsFwMwmHqympXQ7XUKn0eyEaODeqJ8ryvNcMNK5T
oQYSU1YneAN74Eu7VoWA8aK1mrFSxDbLDEVhTrnm3pUzSx1DPI8n6Q019fqI265VDUtgp18SWdwc
siFfdUyvng+9+DrSjOyZ/axzorIkYQAGc3D7bM4A4kB/dV65cxqFrmKsFfFfc8RULM9rciHYos8K
VUwcKWC14TRKVpuBPV9/ceO8Vqe7weMujTyxCgGXJPrP2Zn/qVeA2i4brKB9pRRnrAk1+4F5oCo1
LmdQBpiMQPwRw7zi/WOOpbYCzstTjNekO3/jxJzynvGGTPLf7I49c7hYrbezNHcUe+wJIMfx56oA
Ksj4ReOUTjLuOupHtjlVaG9daKYAsZuZJqH4/jFmh+EjRL8DyLZ2RF+8N1xgSdpto6DHmanE6QyQ
+QBPAawG1/gHELv+IXY4jOJOkH2o+QR70ytWjNGy68nQyFnAalGZYHpyIvClqmMxctuYo/SnyiRt
zMQ5y9dsuAI4IS6wwB8pF1iogCloPxO6vmyN+gdWTrXeTe7nEzjfouiYywEWBx60mYafSx/wu1xY
r3J4G9gbuN4EPrLBhZiMofgXhff71jIrJubS7B/GmOCv5g3Sy82H0/8kcAbY39Enp3WsolupO80G
F2HaEGPW24Fu+fNCsIpwCoTsN29CpBOMjSO4Zx7PrlCNeXMZfty5XnQNkpTBhBPXTOrLczxPSQdm
n8Povz7NCRByl6XBgLUpAncf2bsQJQmZJOjtAEBq6RuXuaAdfN9xy8kivoYfO/9pkIwMfnFCmgyK
tMaSZKK1MBxb7W1sxr2MMv0mTGQWEEaqVqVgxmuHtz5hConwiSunORpB9OiuQu+nvry6pgZz8Kd2
MOrXt1Ko7s3olGdO3wPmrc1qXOKMqhsepGRrcuvnIwtB
`protect end_protected
