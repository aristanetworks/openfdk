--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
MBT5P7y4GdumBri/Kcdi4ihF5uz+uvmAsNJ4U7dWqN4eZefj4j4Lc4EXlHrbKBmrAQa2qjSd5rcg
R5i2+QVN62dG1A8DoKCM2qr48tML+8TgpvHMUuYq60tW1I8jUqV7NeLkuXsrRot19LisYdhFKUv3
pQbb17XI+VE3VskAzWct9oNzWP9UZC4Ml3QtWynOVogxMu8qZDZ4sPaKV0ZCiTzcSGmFxdo7NJPr
E4DVi308cT26l8TJSB3X9FmcyVWvJE/SisGn09XU3n8OpNkcvlfmnjkN3szMTBiDdjGAT2aoByXN
unCOHNsmOHylJkcKzrjtJ96bduV4awQdbQpR/g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="fDEIPwNt3+R7w9ogG/23zfCPZR89wjYlNN5NSdSRLM0="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
ZVeNfJOabsbN4pl0EsDnHP3huEjjSpKxqxHl8YRavaDrrXTqzkS/GLkkd09c+iWuUpyEBntvm192
wcsbV+xp8KaIGvi7ohl3JkFeY8+SgcIfSOyF9NUQg9NUAR1BYOoioNUy+A2d/vhmomLoQyqQqddH
0oFOJx+DQrSxUgZQGSD8qqdVANq/SxN0bYJmSVGF9rBf1uQj0hKjX9nv5uNk+sMXkgGeGfLTcvez
ViTQfUB5WNZBsdleTXLdxMCSmVMfREmJXlw9VjEdPYbNrbbq33mrkX5wPnSICf6mLVEWgJFQl3x+
2ZrsIeyvxw5kfBRoia54NSXZAH7ioq7yXpPr3w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="ARmTnDxzzzqHLJpTt9Smvpo4NNp6D+Ufo6zSXfo5fTU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14560)
`protect data_block
ijcJQSkWRZV7TNoz+/AO2r9VyX1NICZCcHKzXivFLCROwM2I6cPLKGnRQVO0TYN55qkUlPUNRBq/
f1RUegHVrCX9hQPjVgdo5Nap9ruQGhgsyWqY186tlIJuv9TPOBgsWhZlIRtpdToDhax7JXQrXt5K
J7Mrvf8aWwKC3kEe+3ectgJ9RI7X0B8lxUGb6Wi8FIIvQtc+Pv4aOeBNSaRS/eE2uoY/revAPN0x
47R3+I4hV93Mp1DW8ISdBeNnTgPz7eY2R9xYNXgj89B9MKaXVPgxoWCATAcF1D13oIbKjNI4XqlL
Iey+DWSNv46n2yNd7grzEIxrYXu8L/rRA5g3Mpez9mASIO2z2UTsNN7W6Yb1YIX0C2tPApI9b9qT
0fgj0bD7ijKNJ4GjDsQcJyVoEN7f9CnkmcPma9ap9weCuHczYWNdDMisv7yK07nJL3/ey9e3jmnW
QuimHyedONnUsOS0jS5magSMMFB4YjR7KLZPdCs2JS2ugsr4kakxXzfZFL6FgUyKVxTa5VgBgPgm
pAYaT6E8WqXo9nOMmQPcHnXOIbSI6HHnN/oagNxdlUGuZ1RJDGOVUx/zbu+SRn4l/Goi7xF3QspQ
sGW6JWY3NLXQVj7Guopc07XKihfkN1EZRhMYeRRy/zEkXaR6irS8dwQyBShnq/M+bi59uAqBgIW1
tNcUkZeIluXuuYol36l2XynQWxweRGawA3rB2c+MkOu/AnLulADGfnJZljQBNIaezRvqA0URi0AC
xIJFMOYNWb8Mb6yWEVd2qBvg3Jwr0jTecq0HE+4C3T8FUqaRQ/eG35OeH2P/d0KcT1fa0cq1469c
DGhrfN0WiocW9ftCqbfF87YxEL/PZyr3HQ3/Imf7QCk1sktzJQyldz9ljNvxq2k0//F6CVRmJ+UE
2wm7GxbivuTbycb6dBM8X97kw/iwgamJuF7XE/K9w/SkhSPcnsLkRw8pjJr6LCcFumC1CI1jWDb7
kN74PFOC/p/AwfxfU8lZKej+R4q18m0Ug4lhenlFD9YsjSz42ahBLNuDopDkFDpKADu132kAupCn
TBRFXMjTy5gMCFuBkytj/+jSTEiv3tHhuucCQkGXV1EOXoBky3IMHAeJc4W71TjjPMX8A+8JbEoA
eFM2nYdF05BX/OGdJvQA6XxqXTAPBVW41yW8mxvke8RdmJ+ZbRuob3pYefDu0WYgkd8otJqWgFW1
J+f+nLwzqhSxCZRFQ38GJbadBYGkJQHaeZoTnKUY6pD6Y2YhPbO1kwkfwtwUp7HTyeketuuUS0EM
i3kb/CuNYe2Jcan+wnF60z4153OZTZMCK/1s1InYEE/mhZnyNxWq8lxne7pYLN9MyVViMmguF1KF
JQsuh2KEQzf+xQ1Kk/C0XNX7bIk86datOxnYIgCauvmWhm/WZ6q5zsvjfLLHnNIOjqlnWt5cA0yh
TndpN0P+ubqWyrrY0ZyIAMqLBBIUbyuAKjbW5Mug4lSqia/VJ07FGRXHIJVNtus+J7S955PPBsCN
F6L6iZnHVvOlcnC7X+AbskFZqaqc+3yv/pJXnLEw32iwoMxZFhj7B2+4pIAi/YDeR5pzq2e/MnC5
wd6ZDfxcV+QFmg8VepZcmt7I7cYCgGv/10PvyVjmhMItdFXWFiup/1fWGMCxsaZd8d8D6H7vIK8Q
pMmQN8SfqOvWB7zD8FESGrs3erl6mvEe87lOJgpzLDwf9diNgNh2bxo8b4mVX930PV02hRWG2UdP
x8oeF5JPa0VZUTtFHyHrP7vKyB2rPAh2jolpdrLNvSG3V52bwOS+7QUR2gcjxSG4SPFgORrNnWbR
LR4mx/FFSfyd9MWLrpYj2NrmwX5lQ2dC385YDZZ7+kq6NKZIAbKAL1Kd20+kjn8TEk/4hIb22oPi
FXJk8U4zMMj3XfgXw8BoISdzxs9uK701+9EN9VEJVLoeEvVv6R7FpkevWp3+N1ZHKtt4eYr4tQCq
rrZIZ+8You8tJXz1nbZA42CiNGFFlMsu+oRsedYxciMxCwc3wVIZ0wWGTk6mafHBntNfB9cU1kI0
akfMxpKyVuN+/oo8hukShEqJQ+of58id+Q13pJOFQYLdT+Ae7irK2792Xii1bFpFVkbqiThJ1A9O
Mx8YfpiS0MJWT61QiAq68cP79i+twIBkxtKJ6qJty+72fPp9E9EK0fTIl7P6jqQ+zDJug5wR175Z
6bwQRwmPdmGVpJDVNHmSsFvS2KiJiMzJQG1lKTmee2Q8rPiAugBh0DjKx7GsL6pUvdeWLSbk82Ue
YLuHiYA42gfYb5YQ2iDaR+OfeJrlAWTCysYHPqstAiGY1JxRWSs+Oj3Zmt6NvozwaUS6wLgU31BW
8Ml8dKjKcuwne5OJjWrHwf/a9OctJWwkjTkJ3zjRr1VDLOxrGLNPp9utk2JEfh6l1w4gcNE46vWs
i00ANDXxUTHpjmG4MUwOoWweL+drtA1praEdfUDeQEnniLhNiaY1XimJWO7knICg5PzZVzsdV/XZ
MT7AgwJ+pwudZJSTYSAXcrxyDMJVWFi9tPuyg9Ww0aXpkvXJZ9P7HYpUL4KQg9g7lXdAhcl7tP9+
iStDIaB5hpi5GIbcJqhRNllwHAbQeUcxTn1+tgNGvk4DvkrH+absM1J8loK4OQAf9cff6qagIST8
iGAhIu96MymxiDqJ7jDPU3kU4GZKZyYeWbwG62/HWXd6H2IHVCoK1fdGpvL+ghkYlw+002B407kC
XYs1XEh+lTYaW6y6F+bNmuHO1D6IyY9ax5aXORwGw8+7hxROpyO3wQYx54LcCAp28hGbdOmuDN7Q
CbbEZse0G1l1l0EJvRx+bq5wtYMJ7h3BA5NtsmShruLM6ECYCiEwomH3bZEZA/Ej6EU5WThvNfVm
EtwvlvDchJ/4ET7AZPS1Ck6ooP8/ZJapfviZ8pdyYgrvITQd42ixGMyirRA0z8QLshRRnXves2ZM
zKGpjls64jfz6sjw+EAQknmqtFVFUp+XNm7AUTzcrG/J6gLrAunp7yg1XchDBzKtwf4tzrahN+kl
BWXGebmEppxERow+f7dIJn5YNPGfIGCKXUBR7oXjpdbbAWO+3BOYZz7xJ/m1kMUgwBgUzq1a8DqH
NR82qNuXoKTmIR7gsRuVpZP5dbqdFPeKzGAJ0B+zh7gSL2cFUU5rv84XlPuqDDzjUA9K+dhpyGAp
Iur2HOcZ2pYwItVUSrZL/zvepNMGL+JYqWgE6UwyClPYamdnGwczkrcg/osF3fTf04ztRp5iCLVh
4oMRdHmIKk/8ppl0W8a9T4XZkIkq+DRwVgWWyNOofkaWKxqM+KWa8PS+ah5BcSPC7z7CcYrnV47f
T2E6iA/hYwCx8qh9utvq+CZHpbq7cdiX3pQXzQvkv8fSL8Tcx71yyuVLGDlPzUwaldv9Mz2Nb53u
mTpkMgYWz2IK8K6KoBdq5qfACVzN17Y+Hx/Hxq21gyhn9mNuTwP33mAPYXPP35b3czK1cOzAZwTy
VppwPDbzoiipwlyqk7/7lpquhhoelwCSwAs87MpLJ2tDj39j5q8nzqJOikv2ab8EnMgmvXnuJ8fe
L70/z4GpwZnrqR5lAlsRLookaHklCbxU2jkH51zETCqy9GpjoQAUFpK3tpbYpp/k9GXmPD293KJL
hmr7lbvrKA2vdUtHIflBV01pb1ZJ0GzGMUCrMxOQfSM5kosyY5Ojf4DWMfVLw875Bfd3D1AYEiCf
UCwfFgcb4CIAVJNhdiyZkS1WYor1+cvCHCCMPgUyOQuCoFI1eilxZZGllXOEWQTKz+sCGCo2EvCv
MVI/fYtnS5M2aW3DEJiA81HF7ivLaaTGZ4O7tmw6msjmWrmq1oUAz4vtdBxhUXNOITVWHkbtAK8V
CGJXeHYll5c00fY2bbkXmhAXjHTO3zwabJ6HYdEcX/XO11G8vOpZrcFZmgcz6E5SngpG1iS+pVNS
0Af8mQ5vSOt+n9Dw+YgtG/gxlGgCAoYVpD8DAwQIWSyyWkERrH2OiyfVZO8bcIwILHvyOj+8xY0T
Nh5dy5mzNF1taSZvbGuKbSvx0TSo5Il6MwkAZuovIfg1n+XClIZgZXCqgnhVOSw/3XjSfYsuiRXQ
oc0WxLFSg6h7MwkSV3qqkSBTbR0x9/cJ7+JIyLwdT2K7x2NOLKFVg0oDEKZPMAb/o8esIS3DeAmE
SD1dWxjlyfOufeEXFG9BW0HaaT596cynywWqiFconsDNxA3a8Lk52WOlSjf7QJcOSwUuqQ4wxOdJ
vBYExFwmka7jesCvPg9q686uy+dvaCIOu3/1ReGZqdxDinqlnn57K3b/FBvU+W5wP7IICnDGUEqQ
G2+sL4pY2A0S8C01aVQ8XbaQgBo+VFlFUXlOyCMWPEa9dmmrRLr8dDjTleMNS8c0pSqAJCddR4A9
S9ooec9VNMxQRpjQ4KPxeig/t1BVpIre5RCp2NS/lEbCDSnYcUHuv2O+ksWlsnDEjmnxY5ReXHMK
6jm1Mraj9jooxSh7IgxegjVAqLwSLXwZ4BFzNMMYJPdVoUKgpZq28E/NvKwgtD94bh75FG/GKt7F
UljArG1FOxOW8970d7vIevRu+qp4XpJijUQiEgsrHMmzlILexOualITsaPxMRskTrjzWvH7Krb+3
rOMuxReIYAR+AriWYFMVqZ2ZmWWD1t8rfXRuufg5lu8Ho1YW8g9An41xd40gk/1u6MPf9BIhS3iC
+dv1gntpRlXYTTVvkfCEBA21aUB0o53TMVaDHyB+NQcgI8OP+EtdcckiuUu9UDGcdFQlQKJcQ4Eq
v0PuSZq0jpMyoL2iY2tD7kuKNS7SETFav6CU2GBCLMtFKucElWy5QNFuscJK891PxC++ywmdfsB6
9GE5PIw0umoPmh0vU+8liaawTTj1KezwCrg6AKvTx9z+/FDcnqtG8JHIU+0kP9hBDY80NUlyLEO+
rDQpRbu+H1jsKGGDmqEEr5Yj50n5AjQVjruL15tx85iJ8ocOUSyhgpXBeYl2MvAF3jVv04AFqGmw
tRMohGeTyH0w7Nu1Z/SuTsX78X2RYVGFa5NVJnD04pbR5WfNcHzgyuVHCPNEbzx7Mj1EcIe6Py8M
qa4+x9+dJyXnEQAkxALWKMn1NP9uJMbzLryX+N7faiE8G332xRewt1euwu8uKjgHY3W6coMRIqgr
SfuUnztcYpqK1uLkn0a/lZgm8d8yRwPYNY3KSIN0Mnm4PteRhzu6d4OJhnMWdQ0kwHqvxB+1RySQ
j9RyGDC1DJrPp4jpyyK9JMjwfM5r+CJYhfITUmSexU9lBJCAH0n31ymFjlwuK32/IHBpCs6CMsQp
oE7Fbo41OzL/o42plp70f58zvNpL812cH2nAIlcvl/WjM+mEwaizPsScdBTKHMgyaBPwZKg4Hw+c
QYQM7zXhDyl8ZcdwAzqB+xzKMtsroqa/vghtKOaV5He3ZlX6TT6KZjVMGCZRIjsjh9VFumjYyfuR
YDYaA0QKNBytawyKDviqTA9GAYVDDGctj2Uf8wxe0PJf+1tXzAtOOKnuE8DSvVKtVjDdvaLDwhJi
tLaOTrueWllQaVAQkb75iT4hSEu/9DfSQjvxkkz2NNcYCgVV91d893r+vvpEFQHBgvC13jy5r3na
0e/Z4IIzo3ErxfJJD7eSdTNdeFD1rFEbV7dk3m3xs2vzSvQvOfB3LndYvl3511YV5Rjqg07WX5CB
L2EO3LYylcNSLOi8UD1c7VBnjRzfXZ5wSBfE7hLeexDIqX0TCDJskfOyWvTaglYTAeL+dU+eLXT8
bbb1iXzVgqUSGCYKkR8MwofsNE+dTyfN8sHyw35yLlf56/Kbkvtm3wnviRXtAK+Qi0NOr3Be8FVq
swsNWKLok54Zg/lezu9ktrOONlmwK3wsNkN9pRnlW2Cx5EhnO+9O9wJnilr8p6gLdYXnVcuf4tXD
7fnF+5gPmisBUcxInoIMHo8kaeuagr0cldcH70BkNVGZtwEHvtVV+WHF3w6NMm1eDFxhddMw7v0r
YI77k3/HKTjsG66FRdMxSJtXhOvgpS6Axbv+uKrkhzbS+A9obMwxFnGk+LXIObkeeqHvhTR5K2T+
0eddSZUFjC5S1o8RF5Z7KZTO7D9w5m6L4BdFX/2yA6D04G7TFXLo7LMMELBfiE25VpwpjwSK+ojb
OiN/r4m49mwIg/gRn1oSSpAw4Nmj3cb6lAHsJHuKXSYOEh8LNNOGWqsXdb9LdyCa6/GItrUqScUv
cP0XfNYn3HYDueeyfZ6v18VcddyPlCU/h+LT9c32yflLVcHXICaTPqNmGnXfHEo53W9eQcVYAs3n
5CzHnRDDWtzoGyttWDL48ZRtj/dsCG00iWef7/jkvC1PSmaD+xUVqEh68XOLyh6b5FsXxr+APAWP
U5Rv5LfAUr/UZu7gojEWNrLwFdIr3IhF7WNsugnoEWJoSYSZCJpsNAAw/MFQO/2gUtJGPokWeqZ1
RY7/dBOm5lZriWZT0MMYRFQ4bJyZ1Skkqc3v6/RTUO6CjGEq+tTWV/2CpxE7feMN0QyWmsiv0dni
s0hJdqIkiPTaOmF1mvDIwndcScK3n7u/aqbk5kTqlIS1+VD7KvA9Sqkq0Ts6pRX82I+fNAS5nij0
4y1gOMInw0XRrr5YS/wDFJ4KjCdnwVaFBhVTdK2tA5nPXj87pez1AL4tcCyL+7GeM6rP6z/3ye/a
XATBlY4QCBzZVBxh9q6cq6PdZVChPwRO0iykwrGljZAUim6UydGosIepJQM5lDOQupZvUPUCbg/u
2XbKhCEtqwGnYOKMTkkib7hewgfdMLBt78YiG3apVNnZzjA9IatTcpZvZHSvF4DapQqkbBzjWBcn
BYO+qLmWPvc9Z8ffscCzqpJ37wK/cIxgjg/z8mxWO4dYkQd6ERPuCu7AfgJqLebDChc41PRfe1Ee
/HayKUxo/ES5+Yls0k0HqSYC+lFxPZvDKScPxFobjtH3Z4X6szJO6zShmb6DuVW6qA4PmKY/QrvZ
CKhdjP8BaubqUy7/6yN/ga9cxZ8ogeCbmUKCgZy8H1SHFnfwLs1P39ubnKJlNl2alH67vdiFmhTu
odsZV9eNTBD1SvyohSX5j9p2qPje679DCYNnumeuQs1yDysDTpYYAV/PjQU07uLvjdyotbkH/7pj
PTm+YtktT+AQ8mBhSxR8czfgdsa5Fc/U+KQeqi9c8dXlFZZZvztgmTaFJ8Bft6HoB8W+hfJwtgI7
l8l8lpVhAATkg2ANnmNeYGcYIjqW41klWOiST3l+HzME36P7tzR58qLAoGltW6SuG8HpwGiWY/E2
OKR0hMu1MTeNp4rDROIjQddT4BlXZvpBDbz+wSq6gM+jotdngMlx6V8U0TMhoK2i2vv6flm29Ye4
QdKVoXi8ENCkgo0mIkU3TH38bOuJldDYM3rH6E0uU8dwqqiKtDGGv+kemsY0FYRQVHLNe780NpO3
qUh/+HNXCsUnuTzEB/ux/WA6zl6ppo7WrGDQChlpdGu0VR7q26UqfFVoERYJ/2bgk3f15nO7wKFs
e5SIl1rGvlV4d1oZg5KAI5O/j8yH8d6scuWSO9MAO6m8B9J3YKcMkUk+K3Qpc6OCHvSlzFVmwybr
+hNx8Bm/6BKFDnvWwbKvYyIXagrGhp2Kyl6oxBOfUgGr2ntwumM8CssMKmAC7d9zyzk+uRSfu+H3
PnNS628WfCoBgCPqBsWHByBJSedBedyhxvnFGTq2YaRufoVCPID5T/xNbJWehsyTdIYOxZ+HcJNt
57dQ5+XKXjirt0SXAi9yyonlUsehoGkyvNHxB/dSeIGZGZT4PWyHZnFo0ujuTFl278NaAGFS5v+A
W3caa4QlfSvclzotMhDoIKDZ4Sn5uaJ+ReRAfP2tPU/zyhGzYRsPrvSUZKyTLJLA2urVIUNDGQZx
SixnjH+6KcrTp/RyI2dEx2DA+AC8BN8C3T/zBlbwr2umwd9VaNUQNdAPVsnfY0ZD1v3IlkHN2g+V
WNg0zLom6GJ209fThnvN1CtN/BzedqNw0Xuy/bNt2wT6HyksCXti6SPzaqeqAZEhFgTi5uhPmx3o
Ca7BpeWv5/72ozUqR3WMBaubrsbC4ZyjaHntd+lgJ2sODOrFVJL5oIHhO6Mx8OTJGgX6ucWDqG0a
ftR57IjRamb3SX+uLl/AR6GBnOjdyaDwH8qKZMo8Tjrg803Nf2vMVwLKS04fMwHkU1KREPPqdChO
bf7hhXw8qUDNGaiZld5sWK5Q+RZSGlexLVewHf0kMgZLnpzsxqqDmUN1m8oe9FyDp/lRHkqGioQ2
8jxSZEme/WpWU1S4NVSlO2JO9ZuP+mVxBZYNk25zWf0Is7Dzyqd1bjvowPfhN3Xv1qRkrJCdsa/S
YB5wph3cvQ111NpeE5AxoOGSTbmMW1xzG2yLadXAOzVWEvoE4gHCDAZ6bJalG2BYiCMIBPG4iVvu
rNiMB94Ypd+oEP0MrzPXCCmaqjWN+ykVnXPqIB1kBYdyEote0Rsxh2tIE3IaawmAV/F3zORux7/Q
Q3xTeKnZuhZyEyuhabtuZrBkVLhByQgmQN6KjG/YkWCQGR287uS9R56BLJzEs10TtpzAXDZYIT/v
mEMxED1anX6THPQ6KwB2JPZWK+jJ56sFh6J5FKvydYABA497+0WYj0g0e4GxJDPcVTxZAM3UN0X4
gGaDB9JiyQtkYmp3cjpOQFtC4RsZ3jJcP0YNRC5R8lxwsFB3s7gDZO/lQNV6Yrb9WpdCMdM93r1h
eyjNdS+brRvThVRd4bybE6Z9ka5ouM+YAkxflLU62cGmlWjdc88HcOQzdObo4fY07Lq/1e5kvblQ
3io5CvudY+CZlGcee9dkoygYHpgBEkyqp1mBP1/cuHLWDLRhbuRoCGNAbaBfTunr0ffwyB3h1RcC
9BcwJKuOnKbQoXesiL9LDg2r3hEYXPmrnmm2kUGbtmuu/hXS4sgZch+yTR0mBbldgVeaLujW7e0S
JdaEUajo6YkhRq6EnpxYAhFI53cyddr0ifbmUmBAWFSZesqMWVnyIsme4YGb3+87PWu3MADFLlBe
K7c6XuhPMK5rIuuH6foee51KBLOeEMG1Hc0V/uMHjcke2DCU/enV2ptmYmLXSD6g7kd/P2cCejya
G57NHTd4zb++N5NJkrVwrUVaavbBXEILD0BCk0TxRChds9M0pXzgjqn9f+B5HfLoM12qND8XcfDq
URJWEAqZc6/ng8ulhxkO9fyIRe4vnvzbstBqRl0vKyAomqfll4YJojam0RoszEoS+xOj9oR81/0S
6eOZLAO5ApT/uvJWfxjROD6VtfdY5OEVTSqoIiCRt70f2TRNP9BSpR3l1Mw5Zyd4biLD4FkSe2xt
UjqdLaTQuhI2xqtzfVBv1Jrur0ElWCAi1mJcnR2diOAPInYE6J/5IoKSMpenRR+DouDUqfMvw6wu
LZ+m0k7pSOFtizzoIJ1NvY/iEl+jEuUNxwDja1ehGANXqkqRZe+N2AGrdgRbZ7k5hzvMFoX2EPTI
izkBW+RHIPx0e2DVS3pNpBkdJOiB4+eSdsJHPMy1ukvCh9LzccuV29vtIoDMjSrC+3Zlj67DSsLV
evuSzgJ8f03asQlYYXar31sVzoO4GzRsInbbbbW0lv4VJzrHBhTrVYza0ohp5fXXhvGJ0PJ8URSg
JK8UhH7oCPB2Vuzld6E0eNF1dwDJrgGzzD9H78vQNyjclOSUL8B2y6ut63jiQZgCWOFRTjbBIGD5
tTuGyaGyTiApdeB4aSU15Thxf7GGdNKfoIIPyfCoTeVTSx6FWA1Liga3A7KdgkBa+BNuNPLqSJCw
qQlo6X3S+rtKfur6WwyfzyG3X5goDCzXc0EZwme1Ai1vieoxeRyWPw+No0zif6bt0IpjthOislj2
ml7Z3mNrxYr7xS2xAenIF10i4sdGwBfsS4omFwDQ/q61blYoEE01HwopRoZQTXkY4uHP5dU43cvt
S+BMs4RJPrfCXF0ECqvGjT4o/g/xo1gcTYkqS8b4Cmc43cEOqfV2g39OAxY5BiB0/MCyX6ry9rF1
lHs66BQzsJYFXmAIHOmL0mrlU6S2bx7MWd0sDU+x7ExVwZwOL5wxrBYQBy0ufd6BzoW33wQ8GOgJ
Tmka7lExi5EfCZEGgn0sPpwvWBJq8vprcqWN3SXG/driTHIyJ6MIu1ii7OCGaz1fBO09kiatOzjX
lUvXPnqclPwS4JPjzMCbUGo1HvlgSCB+s+WaBVzuQbPQBjxFGsqTXPa+cA/2AvzaN05rVQ3onbQ5
4Y9qX5iFVgA8fR5iSpFv/1XhpbuYSce7mYqRNaurbBFGYvb8xU3nmlYASW2Cg7sRsiuQSMX3LtdR
tqAbRfUZsU17rd6ge9LgLe2dwW7VLJXVdRxTCLcjLd0l7xUJWe1WfGB7dek4I1VzaQqe1l+tU5XF
cTiYo/WNr9Xm6kpLJ0LjiF2O941PiCzWJ8sdq8AifXkqlJ2WegHVjjEqdwPBeFXil+35I/V3oWAG
Ytg9hMLqLcdnvdTCex/aYJJo88CN7TfNfm3qHTgK6G3lvs/Oi72kQ7nrB6O5DsZcDV11O7SI8N+L
j75bgBrKW43lfDKNnLtNN2aq7AIvzEwOqtm+oWLXQ2Tz0KVz5G91Xjo6tTEKHwohzWbNff2h6Z+9
lc7JH1SXnCF5z7DBL/dUEe38tpWM+eJGKEhRS1HrxPLle3+1ffMvLn7lkmbv3gR11b6LAChLNvFK
BPpko4VW3S6WUZPGWCXdIC7yYjCVMP5rW5mVxYFK3cCcIv0DFcLVrjL5fUXZNB366N79i7BX2Sbe
GJIj87aZTbV9EV0O3Dzyu3gty3olU+yOTP3Zc8OS12xdYRnAF2FaZyMvJ0zn5qsHou0w+cZZIRoV
07/aTCiv2FVz7lns6qeOHe/p+SjzBeFxuUQln9wn7YybT2npRgY2gTLgm2Ym9jyY7j26VNFXRYe1
v7fRmiKv7PdyxmGsqq7eKnvBYrvKGxHnzrnzvE/xjRD1PEvZokhCIQw8RIVQhtjOnD6Z3JmbiA+H
njoYXCxCq0FOllJu4+ANsqHt64zscLL37HFkBvA/uEFZzIunVJ+iOLjbAKmvYC6nfwuGbYcn0I9r
vZbXHYOTZppp3XdPHI+XyKho8hZM0FrK+QJuZL5o++O82eByQqPRtY7xiBYdOmNzeUpvVTViJoiq
4WUeqsBWOl67qayoYgwud+ICYXsrormMQ+pi+ommM69Yh20q60FkShUlXKQofukmoCL1+cfdRAV8
NYa06gIaPVrz+3b2tksCewPb0LEkrAgF9m+eUFbCalZUEbgxst7+MlsojtTSjPy+zLk7KpQCceqO
tS/PY5SYGLSYqdCAz2uuC4jO+90cRTHoxwYOLW6QfwwN4I3h4k87WPckZRsc7WaZrI4S5Fsazszk
6Wp4g9c4K1z1jqGQLHMU/fb7l+00DO8uiiqnJxl4tOrBeWEz0f9cuN7I35CQ1R9adBpwVdYuNGBt
O1g8sAegUerqIFjgWzrtVV4JuHiOpU5214aH9m43TaWyIbbw0nLv5/6kretqpsc+jOMdSp1oA6TS
zs6aZn8OJvTLW/ZdKyv1qRtzPLwJ95hlswDhlDO59PoUGun9lkVeVDKsRyhQ2y/Ec2fttog7ox2+
BRBFA3tEDXwjKvaY4bnxAifjDQHMaXHBC13ArZe8iqmM19p0STWWhlfN6Wdk7NTZlbnDpv3Kcx4Y
AG06PUY9zxi/4gnwTgrN/o1pb6wD1kucnhGIMk3cvrVS9Jjs75XgDXrZRNwbs94lno1WViB18Ea2
E+Vi2ubMi4Y2ALHIl1aw5tvUiVCWw/7Dc3J/+wLzPubaA/NKU5MoJ2ECJGf5jVTh6VAFfVcK+r7W
MIgNbTzSlyVVak92uXtpWVDDWCAgttJdw3y2MlhMKmuEa9qT/gbY2LLf2aDJPMpGg/GX5ec0b9vo
o2DOLDK+UawsUJZ5CCiDgMYvGGhFW/YSqBm1zL6plrq1MIpozsmRGZmj8ZLFhZ87TSeoZWlevcOw
vIIPJVIDJMkcpK/1DkECc4ODIw61N34/8wb0v6rjc+G3wWomgfK+9aowlCK7hx1qGDhC6Q7xfUvK
CXz3sm81ImQDlz7g4W1KV9GZW4jCoeiEuZQhRwIXbCUEz0zdNnaCPBmtbsc0WHkMongCDdULuxth
LKL5BsYpRSA1owdr8nDvG9VCMwpHCHNTdCNTEsKcG8OnEOj9Tg8TLwYdRob2b9KFUc+YnY1pP4aC
Lg9Ph8n8814H5RnNmuINElRiRKyKA0Hm89fzBU+D5+u49+e0S78z2m3rkinm8jxkxnDN4xarJr0Q
sY84yq4V6SaoEfKeBulF1CvT2BPppvXvYbiXBTM5xYdqFOrJSl+YYhbmZgnfp0tBlyEDN2kGUUHw
uN7NC9DjhjhFmzRHAg/ALJLR7oLwHLGPCgX1iALp7x15JUr7FnWYptdnOZ8ScuhucgGQ4cYlC01A
fQ9cDhm8BwrCshBDiRXaJB9tFF9vlwjrtLNO82EqC2ppmWMutowb20S0lH9aZ+aEJXYpK1UASyoT
Pu3HTAm9KrstpikMzY1RROZwK/3ZNIkX0B6QOZnMMW+rAtt+shdHbxUtJnhWHEoEsSdvSQmAgbpc
x3K6SMztWF2GX4sebzzXU+0bAYt/1CWgFpJywm9vClnsrmUuSmjfEM5jSsYpEfV22o6ZQg37PcQp
awSR+ZPIkvFWpG+Mgjd9ACA6QwnYkijppUEKsazK+aEV3rPWmXFFKi4w5+WdKdOcejgHh1/FOXb5
Gihs0iwUn37ogq78OhCCMgUHmL4Ibntlxmvv6yivcNVkEQGCgmrmLrq3zRmfb6pr2FS84hr1ltl0
PVhZ0tzcgCRaoxR9Yxd+PHFxiFwAAY8ETjDbqoiySXkDFqPMRXA75NiklDSaGmkZvSNJxqpVzQFd
F/aW6G/YrV4JIqEu6Ya4LbR8PV8v1l5SbcXCehnVzrFAKw/b7sXX+IqK9fYu+zRCbVIzW0B2rbF4
tGW2IhsGJ0AlSG23fBpuJUPgPwcWuI7UPwisrEuCwXCCv2+yS9R8H+0Der9MGuq1ENfn7vzR051v
/wEqGEaEwpz+n5uITcsoWOgdCKesLFmYmhciFm7S0KLxgO7IY81dT8OFMSGaoQMQ06H0omc+EvJH
eNEjWwPLE8qQVjXGR+8VWHsF4kgc0N+8Zpu15jm+1OQHU+FgDOatqOmzJBFtMm8UxwY/Oh3roA0A
CLrN1VCBtTi8MWsOxY4HFJ3yHBZlMTD8Roo/vBeqlw+sfwJfCSt+Ahi/rsFFVw+c5t6I3MijQ9+B
t2WRk6QxQQ7CbiLjRW7egtkLVJ0JVoVD4/R2OODZqs7TE21Ts9i6iokY6cASrwjnwVu59OHlfvVT
DMA+GcQmdm9x7gT1+paUASd5EMwP5C0ZwgBDkAZT/pboWClwmm48ual+HwHldyQMMP7dqv+2NNvK
LwsRehWxAAfay4/F5F5fomOi/RhZA7t8pWu70QFXdXcmbgoM+msneNAWKz+9bFZ8d+V/RMyUkNkr
wWamESEGFL6kk3zC66HaM0YRBeYWSRHnRutjqsTUOWIVrCIsFB9P2QeQUarW5nSbYBnBL9fjOPfp
09SaIjMBapqJ2LySgyfyo6Qki4Hra2WPgYFPfLXLeccO7VvOjAzZMndjsUhZJgQzyTjWoJnt1t10
l3qlifwgdpjZNgSHv7s//ecWHl8eN8hf/oJa9e5+GtgVQzYo+NvtqAm5EMsjpOfwnqK+5Ss7wLyo
VQ/rJZH+uGDr1iVhWJbISr7eRGNFdlQWw0YmzQX99oRy9PFJ9BnnGqto6mBe0mTmh3jWbp8G3cJx
ZL5B09pOSb9YwPgJopI9e6uO2C3XTBjHbK0QnEoBxBtaEk1JjruQuhawt70zxb1gtmHVdxoQdH5N
kGR5RYgcVaf4814tznF2naTNZQLZD755OT+7IGxs2i9y5QWRsfZU/2wUjKChg0hPnWXL/QcvprA1
ukSmyDvV65tg/TfLHOo5NomLXUQoP6cZ3uZrLNq0+QJKMWOpViHGaMXKOSNGirq/cBYSyI5yJ/7x
YcODL5JdhBSOOPYIV7lWI2dpQ2vyMI5/i3+BptI3HuNrxGwTTs707BE6WnGNDdlP+APeaV4ZWfLm
tRwlnscAhryBMl69kbxWmbySJ05048YLsVq5qQK4IPe387ouGWM1d5Nd6no4Tc8866LnLIANxdun
7tNNg2l8O6JQINsVz1hRC8gjvx+UQVJraAatZltT/tieJr7xZcgG9Kb7LkMZYvhykIkwRYot9wBi
fldABR2gCf5dTHbFmikm4CfMqkJMqxwF6jj82lyjyZajCu34IwG9gAPmNXQAAc7Y1AhjuKn7hVKh
3PFEhZtgj8cLwifXPWgSRBEsUsfse57RJBbh0/RH5xaSFK0CPBmF78yc4ABN/sy0uopHFc2a4eeE
L4ET+Bpz8g8Xb0VmR7lTpMirtp7LLz8fm845i+uW1qOLmDU9QMeSdyTbQ9DHPpqC0Ht5HailCpJx
58LZiorpRkXLKYae/+2pzmm0QG6mifVUtXVBSqi1jBQJGD7X1d0tBwQQvSX7HyBGUSoIQAaVIH30
YT3KjvL9kwTADPfZD7g1azQGcNC2tnoAxmu64E014jGygUYi8UdTovTylNJUNK8K7nQIvR3/1TRB
A6KbjvVc2djXPM9ejElXZvxlRidbwNuTHEm0SRmZEodYj96U/gWx7LSMBQLJddVDErS/ri66Xh6/
EihgbCP3AA1pd+Fu8JNggXICenh5yTISpZKGBusaYh5beMIFrXloqb7wPHa7Hk0zM5kRnIdHu2Ij
GKAHYmkng/7sFL3n4++WQBdtYkFIpAepeoEeMse/3KdjYrlxWAv1vcfqJJBnxvGGnQvLfN+dFgsN
iQzDddyHJdtmLWw3oL+gyytH5EWxcBhqkms6I0bIwTxuMkWVakzabCoQA9V/sxjrmpbBYKc58Y/h
EuKVcnk5fbE+q1cNdg3gNIWlMG/g6zOh5SD/1fMD5pPIKMSf2d6b+cuitCsJFHI+Bt7E+5kVIxU4
GeA9WV1E+JCzS2u5omsdWkz3UUt1pmc137WoqCTB9DOb7Lmng4Qd0uHdnHOCA0KuvN+WtoLv+Mlv
GxUewMG4j8XfyZeIk0y8Jw94lSHOhr7dxZLL1H00Hq5e03s4esbB/U61AjSaW0QEdE03/cGZDGpy
T2BDozqesdyM+2WjiM3uSqVB9y1b0dlRpKj0ykQAKTWT4Y9Laa5V7rU20ld8kUMO5Xrwjibl6uo5
PkfgpnEpZJjlQFlqaC7+CeVUq00JDAnSocBRKci7PwLKZl2Lg2wuNOURgjuKcTImgqciiXucieLz
cMrndsi3bNao/bfUw0jOZy81iqzqXI2BKveVK/acrncJzutBRUTlldQ81Oi61uzIxWTOvDjPB/kO
iZyNgrJhMoxD2NrcwmLWcIlqhhvrk9BpUcSLAvD5flMX7yMXcBsIr3FBNEwAWC/XEcvMGym66GG6
cKlLzZ2lFquXRFJJJT7AolraIzvC0Os1pfRcqACZpQ1+Yvq6HkRFF9F8qcbfhZJxGUREO9nxAE+T
8KCn1Ri7Snt6dBG/f4E4Xmphrv49W6ATHUg0Bwql02D7uoIvAf3U0Cc4NMJ0EjyqC+krhX4urj/F
2W7HNJaeAn/yS2/RjHou1e8jXXr4wRvc+Mg+xAquo1iMO5OAw+lLktj5h6UyLXX7NdpZ6V6J8BZ7
Fq7WvxQ+MBqrEDiTN8xROedqGSoF7eHPEfx5IYmDJDwA7+6BRY9MLhWDW8MlDllTCKIUx3ix/6Eg
QDFm83KM01B96/r1dcu8Z60NW0WvY93xJ57mvsC8FG4cKg4o4GDfrnUDUMysmGK6jigFU1r8y1bU
jF41wugnmYT3gwheCKboGc+h8A3beBzd1entzB1U7h/G2Fr8FnLVFpNxGYg8d8qi/V1V3bh23/CI
W4tBuxu31k+oGdz9NsD2CWceV+bG6TpoVpvJkta3NNEeOviAcze4HqmlxBb2MN+5FzjXStTvB264
Lz/IXQb2fIXjpaNNB8UaCU9juOf1u6Qm3jpQ85BF4kr6Y13ym3Ys5N4W8MK3FAIPUy8IrYTDPcVv
3HTvYIPXcP0pJaH2POrMAhF3fCt1DEEigo11pdiat0flr1GtN/8fLuWogKpUdXRihT8zHCJawiK+
Hi8JhfKroCJqBUnhq9bI6/G038odEP7dwlwedpElyoMI5UsSs2kmRytP0LCaPhKnZ8w9J1SKNbuP
iYR6ARgwvt0QoMPnuEgvZJ+YoFnBAA4+S6++ozAErJRVRbAgwhUojJ0OdFgLlzIFL2baKXDya7Ms
URbHe47a1SgmUWlQJ0C1bRtufLz4n1xfrkjf2EzLyvyxcLvC+vo4qzFr3cpplsFHC6cRtmGDdAho
iDIMXl6nofmjKXWhGAzjVHwjv70IZVCF0NDnpTG6viD42uDFl7bamBwnOe6YV6HG0Wzc/v4Eu2fE
mO4DIWPMne16Z+IireZ17du0NQDpgs/5/9wOjtKuAEJfb0UL4d/Yy5hQzRbNlzpQm3akX/WqiJHL
euDjQWt2qW/llwZn8+mP3Av1a6rSUQzEgfIvnLMgesAvB23PonC7nkrTR//mWWigkuT1UAucQiQo
ZigmzzqvU0gX27bh1MYmpLNGmqH/JlaO/6ExH60kpa0SNKWnX8IELm4zGurcnYRMKy4xDpWQADci
q67PCIwauUiun1JAo0yBsAJ+ZQe0g9pYmpx2jSXV6lF4gbBny0ycrLzZ2XhH7R8J1/+UKiAt3jU9
JQDa49uibjzcInFY47cUWcigvoiVbH+PlIMQ49bxcX86DEzBdcMnHucXBlftUuOCtmotJXPTw3En
BhNvtJe09KEvHMMCVx6Uj5VIY9yp5C5+Us2cGYJOmUsXpZgxgknnfv1b/e/z5N2KdHk1Y+0vcS+z
V3/5Nm64be2p9vjudI+jnZJiAcc4FaTUPxANQISu0oukrmnUkpuytZH1G2Z9JWcdCKAUDPoG0Cc2
oMdA6vD5qMM2+sQexLVzNMBNfxvrnrxZJo9+qhki/hBKSq3M+3O1s7LKKBJnPkwgbIb+nTLBvKq3
IKPGFS1nT3bR5ddHY6ZooagUGJ/YiDvvD/S/wsKotHBoUgy7CSqghRwBA8fzRtjyWwq2ZJEzn1d1
7apz02P5gHGXFPrUUR1P3gkHZvEXsLDqWXekQsfvfZ+Hpdo1w9eDggXhl5ObFX0AhhKXHkrmAsO5
/mxNZs4y4Ma77rD+APiAwBZxMwP2Bg/o55KuAqJpX43qFt4xGamcJWuSqCeRBF6tY52ti4wxdcQF
3VMdr2+Gk3oaMBvyLViiaNIqFRD3d/AQVwOYMJ1a603maNXnW03tQk2k0xRFNovR7M6wzMB595Wd
5FILlN2BPReH+yaS3JwiaOvvGM2HepZEYI+hMgqZCR34MUO6gyifI+xMZQrXJN3Yog5G/UVYlhJI
54/Y92GDATFL0FzMCr2igLTWuK13BEo+UvvE8kLneltyh2VHufxu5M0BN69Xdv4kO/V7QcSuC4Rj
Qo6Rc/FcfWz4sBLGQcsc6zMSPRFyYPyb4Hm1h4ifPBFGyPP1ZqaOwIYCzb67kTL1OdrxW8xdIrgu
3JA1b+lgPU8pLi5i0urxWY2RaIUpfhzsUaGP64WLuCvl5LROZNSrg5eaGjo+B241rQCkzGYlAlzF
lAPlzzEtmdfp8xjhmxZP9HXu3kIxZcxA5AYyLanxQrkme9er3jUKW2xUuoK12X8VTbBNaLPntX2L
TL0QoCJUB6ybRvX7AxEzr/WW7aS1UxGg6UhaEQLQ4zqBNe4s5Z0cHskFxpytv1RjVbheE5QZZHVG
Y2OamTkLc/j6pVYexW2QjYUZXqysVv8FYgYI39cgCFZJAxIqZvcwwK6pQvRdCJRRCFjYhzCkCOgN
Y53rljZT/8oSv6P5U6vfvt8d1rT4S39TTfxBEwXpb8aw7UiXZGcDm8K+0hAt1HEGuxbfRLzrtzt8
w5BS6RooEPGYJbnrpnGHc0d5P59PvXJjacgvycaJQjs7pEyf1iCxZJ9xKzdQdKWCVY/YtNW3yqpE
LdptmeSlxHCfeBuCKYbXm12lmERrVHqUx1KEeSZnsp7qKEJhXbbfGwyznHkxRduz4BuUk7Hpxs+U
bbrzw7Uyq5c/Hx/tu9JewUnXlEhK4Xy/lBeD0MPkaHIkVKHEnDa36nO+KHO8JI3YBkalcfPltDiy
q8DPabzCWWC5GITBTvPxfPAyUTwCL4OSIGrSkE4z5NNFF6tKpQbBb8l8cdsVNIggrTiGphzmzHIu
QGPhQ+2EXKT2/A83I5xinDhw8q+6wrXRKM4BGZoaf6wogOjp1MhhYd3x51XWKOZybXXRalkrsy25
GIw+5acwUHXMOk2utnpEMiVlLY/7Gg/a6HRc/nyBxt/UIVA6R56DEWZaqX2KnBF/Ytidykn//EOZ
FecZSOfOiTQVaQLB2gFM5HlwIF6QJmtG1mqo2P9A5tf0xUMo+yT/AGTZDgtfc0g86EFuqZYqWJri
Gmq44dURmAYgLvaE4516mnrvrxmERPQzWYw4TFhxWpGS9SinbgyY5vuA7xpY8/rT4BVhBKKBDt17
2sr7mWJil0D7MIPPC2+DyVxd1JInpSPxfsmJT+vkWDWVTfVqAXATXyu4iLJ1AAqdorg7f4wCfs3y
NJOHsAM63sFUeJdAUq89R/RKus/IWjjLh8/ukI4RMiwiu5GxPnURa0s1TA/g6cLKt+Zrf2WHP8WF
hUvaC75pebY7yyZGYvX6tZeFDWP0gb8Youpfo8TNRKa+MZXdMqTldovxDwJxFb7udv9cbKTRN7Vd
DK4A2YnDCKnpF/yERWRp0WrR0PQ0Xj6h0O1QRRRJbq1uU6g90ZKGnq7ihRpxMUVsH9uLQBq7sR9a
XevFi4l5hybKhBEFF1fPBS4dZnt8GUqPPw0J1C7jDc2v/uMUncTJH7MKO/eP54nBzlrnUBcsGpBs
Lm90oNDd6hmTzUCUN6UDM/Ff4D+zgIhiLu0TzIu7HdVf9fMDGLealL85D72/skRfZ8lf8MIdo5Fw
/ENX2SmkNNk3bEhRa4nPT6wnP5mmptU7kLRfXPSKYs6mK3JolLrTzR+b241unEchn7fQFmDHFQeI
IU260kiaOrxi18DQk0XpMZLbJuNESDxiD8kgMZkPxOH2Hi9aPy+rxzHCyMCiovIakQl7bJtOx6hP
4IEph01Tea3GC3YC4t8C3bwwFtRkf8Qt1BV+d7SHi5Q7b2y6sNhdKOIOJcmd6/HHM1ST+UxIlHZT
dwATVXWFmuP/sOHjIHZ7hxieJGua5hqWcM89LlwX2qlWOGqE0+pG6wd+7AiahZiNPidK65l/Um0H
V+W9OTalI4vEc/gGZRqpFiiQv2FjfFO0HA==
`protect end_protected
