--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
W5UXlPoLHfa5nsIUUkhbmSerZBM62Ts65ubcR20dCeIWZJsc06HbSFrnOvlIu/hD9aUWl0dynzw/
uJVQas/IVMSkp1md2thA4aH8eD/Wq6CtHMhLsBw4+al0LQHrt0XbLBziGNs747kK0va+nWAaCDEO
//jbASiaBSTqHD5LBBvtRAjWy5WzB0FWFirj1xyIU7ydHb3pypSCwOWWy64byZhXQ6EPjnSW7pf2
QzhCXBPdva2Gv/QsKez61aYEhA0eaao8FSU80HZ6MC7vgmOhMfFIChgLMHu/JYu/kxQe0TZ543vi
7eaR8c6iOPHWXA8QDH488Li+yWtO2P50MySn/Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="nTe8drqPqnIWFn0SuUEc+3o4mDBOKNN1hXSec87wmxQ="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
pMPd7vD3itgGNtLSbpQBN4AyJH9DS1u5Qwmcdh2DBIvG0tIOtrpXnMGivzX9FvL7EESXYkxynqOX
8cggtzRsOr65FZvh0veG19RimPb2YdjfK5gNfuTz5o0ogSqQ4e3FSBK9sGzPFBlnVnEGUBFi3vql
A7gd3lHlFX6AEyUeImtuyLlD+PqHXqcnbbTrOaNnmaRdjjvCJGXooyEUF+Tt3lgXjfU5F9/HBAIB
VExLKFAtr98jWtuG4HeavhnAv5BNIqXjHBsaIaPrzMH0MsagHeBomFOifC2vxdmerJmPjwNyzaSN
Vd+dBva7KVZPIVe79Cs+y6JKz2db0NskdZYvPQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="U+Fwu6wyuk7esD01KJoK5slo60hx7gIXybI0SE3sI7w="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10592)
`protect data_block
2Q5RVAvEdkdaWAzet63P80Lcl+STwPdUMTtKL+jSE2H/GyA/W5OKFf5128R+EUxH0UB2pW1ZCVmS
OuK22znhRV32e28i8oU1Y9c0zx42muChCQ7n2/13uwEhR2YrtdSovOxJKwF3SM2Yn+sfYnKRXSg7
qbUW+kxjyOECx/lo/ccSsg9J8SV0D2M+y0EHLYsze8QeqqIbE+KaFIpBnZebTdgCJdJzp7V041vy
j0HzAWbxP/qxtelHSvBaalUItT+8IdayKixQQTPckpA+4HUYPSz+IzbFtzmYkSSTXJ58cbp7M4cK
ab44RRZRFkhYYsVqD0jipuzoxqsYq3FbRKrqS9LsJHsERqqRMluN7UGtEq+IuEn6RiAfMryrJ6J3
oSQeOT5/o3ISBJFF8CoDo9Vjh0as9WNHQRtmij/mxBuVPAJicai4r0qbNs3SG9cICiMc4h6t8YOf
1a6tru9tBpfbI+h7vHccXTA6LR6oRTg+G8I0CIJbcXp+IbrTZb57gaSEC7oNCJxF2MOPK5xQV3QZ
LbZPkWRt6VO2AuCwBG2SPAn8H+16Ku4yfNpvinGGDUEPsqrpyD5GhTJX5OrGQS/qCsdZRsDaQ1Z9
PeQps7CECMQo6DJv2V5tBe7B8MQVbYlIu3Xx6kQ0dugfGu8WszF5LZ9Jn3JoQodJkVYEHmmkPqBc
7vEZ2wH3ST6SSWXzsP/X1otfYqdDF5dkdcjlUkFRVT6cWJPmpV7naeGSWwkL/YfLzQyCee1QcW9/
zCnuaKxrMTzO1kuyiJ27zrMuC4C16lyuKDH8Uo1t36+KLTvplrb6KyOg7yAmPz3dkBGkt+s3yDdP
sKlZGFm/DwfeDtL1Qjg8MgZtdRYRFycHUnVYKQbjs4zbsTXQrp0B45stZmxU6co0rEKYKZ15ffPO
UPG9A1Cufb0iNjSSVeceA2nM9JUzVs2dDQe5FfAzbBno+sOAaaBi404RNVqEP+PA2Qexqplw3+CO
wmSR/Z5V2ZjvG1pMdtxecUJjamRHBBeJu69Kg7C/c/yW2R0UwpZZx6eHXyp8+7N94JsNWU63N/bc
9oD7x0cqoKfKMyWPuKFam8oAs2dfqUaimnJ/6xglshS1SAPLy1mTeWtKll92OTF/bylia4Ap9//B
OyhOec8UI5zs/ilXkF4VUGDidMk1h8IXMMgXjInaSxPB9LgJjGl+/AfU2izNFGkSsFwofZMezdCp
kXe4l1fzCQ5pgpjgeH+mDOSXfOkOXQrxN8kMrCdrSfpHWX6BeQXlNFIlf70QlP6PN/3I5zHMWeCZ
qFPJFPNwlIev7ppg85+9ikv7oHy3M1DQ2tXjQJaOT/qIkmXO1nwLq8OGHyMDVkhC8IyX52AZLCU1
j2GghhFgUaxF7NCfHjcefhSZpjiJbnK+Cqofppu1SMAW+op5BQztX1uPI08g/5VP1bzKwYXglaWn
aT/wL6VYazWExlQqsEGbeHf8iq62w4BCsJGYWHsiKRYDh70dhenzht2glMm/wzNH/f1TuKvjiHAn
1x8ZTYAuRyVdGnMZjT7hfz+WV1NIZuHzcfdozbV1JgGFnYEG+KpUGjR1QyK21vTPOmh076EjyoqX
cnhCaD3XYUg1jAClVKq7QXWF3vPDi/ms0Y7PyQ99YuW/foEwtjGqgBvn9f9hpLtadjPf0+JoLrW0
5TmOApN/QG/rx+amYQ8dRb6BjfIhjmFzPxI08zz4jNB9zvC+PmU7OEZy8kpwRT38PBVDiotBqrWx
SUvzR+slMNduSBtFBtRy3pBjF3LTq+panBiRHd4FRbSm3jMOnqMMK1WIhax27umxNPJncuJuf3gG
IsMdQpRx6OnByGxT8rQvqCJAq5Z9MbQW1CFwcGlhpJTHqZkrqmYuS9wX3JZiOUhJh8dIuV4vrcnZ
i1yuSJOE/NaBpj94Z+iyL2+xi2ONQAyXfwHQCqhBpBQJ5uQvkRWpJY6OgKS8UP47LG+AsjWJ+QPq
UUhWmawuhYAXinW1cEIFuW00ZcuNVEKs/n8XjM5bFwYg4GIkqLR2MjhDqDfwgDMA6y8kNuK4kyTu
J7yowFcfFzGuZCTyyqUDEs03RZBIk2skzsVeEWPG1sI7yf0vPoXBVTKo2HC8XJG22R1+KvGp8Lz7
UoxoDb2qh47lqSSMBszDYS1zcNky2KqgyQL2Dl2Fv/2D/H5i+D5VgmRuGB3Hp+cEwhsaDv8KT/JV
XFoQytdwaTUEJDIdhUhllRDhh5LXU2uu8SOcouAzl3O/G147On88JcPkQESkyETvSZxukA2uFKCE
kmoPu+f/Gfszb4Wcw0pnzQj179gWASq2/mFAm2iU9E4hWtNQsG5Jbzb8n5JDbu5GQHCcar3ixlm4
HX7mzmJpLfiHGaCgdPJkJvrirpnvRK2+xBe5vFZn+rgeyGVuOAqe/nys34qMAOPIkAb5yc4N63gv
AmzoJrskZcX/qDefA9ItqVaBcHag+p+M6zodZkSfF//3AHWf2XQT8MMmjmqjbkR/zheQMAEaV4ot
wNvh8fdxn21GtixXZPV6P3TFeOO58+8sK006fFB1HZlTnyCWOyENqQEecgIRHTR5kTaqUzXuw2Ay
yWR+2xcJig6FzaEv33Ymz8hGHTKOZjOwIlqAocu+515GMs1T8m06de5OwkTGHxkMJLEzw9onzAjc
w88fHvk0JNGssCKhQfF1bmMv1mmkCr06lyB3E9ILEOC3NZH8BQB0U1FKyGgR78ASVl+210vO3ZB+
wsfI0eZwel3yGEOiQ83LAMovHeBn4XHW+TZaEZzE6JzAGT3v0EHTPCILT2+HtHNFletgNF2GWa9Y
47Rkw5QONnOdb2O4A12rXmv0PNPhjUcNMRFTiCutxenJxXHLYenpDe3qVHTT8U50KCoqXJUGUx/A
PqeprH+cRWgCt/0kLM54IAGKd4MEM2pa9qjBsLLw913qd+Zkx+DO2zxBwe35UpuyBvt4AqI3SdA5
pCM0NSxHD/pciKgIvOaEC490WKkbWC9BDMWGbmBr7hv14CLj3AYVIgWhQZJ8orVuJWN/YaSdhUnQ
O9rM1SDHDa0PHpNiKkQQ9pgqc7QwBz2b5KjyomIg+cN2FMnrWuuef45MKwAqBhDdyZV0wbEhdMbQ
zfq21qUGLdK7+gGLdBSuUC9gUj+mr/riJMVcXU1BVZbJPSszOgwJHLdC4w/dX/BB4zXGqCYeFdMC
+ySQUykIJobZfUJLvnXdYXpn+uKCN3rSfhJUI7Fji9d6CNkFIaAtjWH7TQjBHb7fwJ1ocZA6M/2t
fFtkwezpISjJqCCpndTm0LgpLD1y7hYlE8KT0A7q5P3MJTrxFNsyefsOyI5D7N0OY8b214d58MvP
73jpbIxQae1H2dKEhpXU5UhyhUgH+MIH7RlMB2O2zM11/t4VtOyvbp4kcf8WG8i8wGMhGl6+J8bY
RGnuOvfVY0s0RogMf17NV+Fe0qQ9xRzxjpK8u9bR6sLHuuc74ENTX088URep/ZXNX8U2I8t5ZY03
izmvktgPfZim6bAOAjKE9eA2fWtaP9NXB21awlVSKO4Q7PQFic8X8garhFLKN6xzsHu5QdAbqRer
ofCxX0b1kc9Z2PHHmdVp64HrIydvuo9DqLfC433I47CotojNTPiKYQaOPPnOZxav76ekyNA4c/5w
wlEd848N2ehL7u+w9BQSY3o6rhpGdFyR9WMsrSxh364XpPgTNuPrSkWP7xnD3ffbzwSgRTW4/rWn
rlBx4Id/zjoFk+B+kQ2T5047x9cucO/F4BNdXXF267UyZYpQZd/tdGYggyByg9kMmbuNP7KSZUuS
abjZCEoN69xdVeFKL78UT/PAZhHyWbVqP2S5YQtF+dEYsx7xTNV4jkh9I85hI39GA+27PQ7nfPSd
CjDxd/5zs59f+Yk9LhU3rtGXzsZsLrcaBxEDTmyG+Vpr6Fw8sIaW77OTBOrdTz/w5rbuRHvUxrgw
vm4r6mUKZ+lF6cvlCCJrahkZvj92pBdKGlf6Z9yQfesYoOLObFck8C/laPEkJyofbT6sq4+Ax6mg
JU07MAqPcA8lIkVeap+UG4OghCcPcVpzO2S7NhUdk9FehrDBJ5idar2hjtcvqF82YeWwB3DAJR08
1XATzBGLsX4YbbGjIQlH1FFCb+BybffQAXtBisfiOF95orPDD9SDIByyPCLsk90jkKMCZowQMMwm
CuHttMefZT3hcoHAVPyFToL5T0YQI12rlOJUba6jsKQTFs/j2vTcWEmr37ezHX7IK50oVL7QBHyy
reDnet+z9dOD2lHQSqPe6uTvGSrcq1FK6pgDaihupy/N79B16PrNCybzykF51A4zXFplfCK+ZNj2
eaDOti2hGlPlzenCtELybE2oHDNHaW6uh6NKMN5hGeHekHX10e3vnQx/CFMLPn44NyJoNdvf3z6/
rDOlTqidkMbKd2MNyedjSIzJAtmCdK+DaxWcJrRUFqgKu8r8kEiklZ0ZaRe2Q3yOwwFhVWPOYL0H
gSSHyrkhq0Me055AUHNu05g9O25d68rTnn1YEgVIWHPGplbBhs69gHmiq89sgtkBxmYXioGSv1r/
gmkdVm49d4esIax+GrpOKao4lwQ3+o878CwaR07lb16fYqULcoM9m1P8KBPv1fz7f0sSJehCl+dw
g0/QUisY3aniK2yD5dzxbt/KL0Honc4na60AWq7dcTkSCQR+VtM6Mie4sm+pU8fJ2cih/ehgRtBF
i+V/dtLhb0/BBjD9Ye2my8inigll++J6s3vNTi9l4TW26XhyPCo9K+6mpQocf445Co6NVNj5gSbQ
hlqe9nZ5CianeJiFwRIL6SX6/VTXnuqNHmKlWmkwV9r1jCoTLC3ERLT9h1hAs9EDHUi9MRtSye6P
TJx1cTmzkyXUD+YdcgLkxqZlrXCI1s3wl3hHRHaI4V62XxErZPylLfdsGXksuuf8v5HOC66jGMde
hpi2W5YUKg2e8XZ4viOPq5m+XcLd26WaD8NaBD9CGWvUiRkYpy8cmwSs37yt2y2aDIF84AjKXKfD
g3bLMvZS5bQjN8PwcAO745c+U+CXngkjv00epFutFJv5tk3C0sO4t8OTA7G2sbxVGKeYVyif3sLv
5DH40CGIxc2WionC/GURW9tBdpe5L7htjWMF21OOTOI614AeoeajMs4YdaQhtOgAFMMHFgS35wxw
j5XdP/tuFUzhd5LwDGJ+cj6qthhFBSSXnCyaHz1cTSpKDUdeYOoIx8J+G/SHLOP1CI6IUVdH8qwY
GDr2gJlq2yuvWkwBpgqh/7ARSqV90rD/TFJA2TnAgwIPScrPKgSxE6/uEHlRmTtGIKo4ULbVqDoF
KeFzGTrC8E4ESSCPDKBgQeyg9WPfMpVF7gH5jNLYzI4C20lgeeE9CFxFA3LTSTrX16JBhFIF3q8G
EmBC6DwS5WMAu19UF3nxpm8KwcstrAoFmxwiCHgQdAhPr9/9OlTAJzTEWpsvIYOGdnD4e42Bd9+u
WwqXaeIzZWLXnd7S3fHL14MtP3vA02hkAXUakCsJEo9Sd3he0IuJpgmfciG90bbWBKAHorwqB+pa
LK8cRLauiA5g0FNcXA32mE5BawBzJd4M3f4r0lcPaAx6xySAWgnj+GmF9GHHDq7/gPAdil1CVEMW
xTqVe1urn+ts6r6CXzIxxGJSnIyzkRSdgcYD6XWtdYlZ+5I9Vig+WsGcSa7KYgoVESxxfcwYZJBx
eHayAGBqIpZAEK+aiPznc5oKVAnkTi+j96V0iDyLCXEiVmoc1H8CsU9TSgeU3hkzYJeTKEdlLTIY
bWY+6VLLJIBVdMWS2fkLQB1VAN76wZCFj1hs9NPU22zDrBsdwBGU2hXzmZ1jTvldJ7Pd0XMjLPj/
yTIiV7Q2hQvBMvYNa6Ci139GAxtB/pUGa/SchF9aiEUxCibV0Wqpv0m5Cr7wjr7SNhm5ITb4S6wZ
aQiNouPw0ThVcM6azFuXXL33YuZ6xwSpJwZSf5WAeuSew4Cfvn6lytRm/aL9KR4LFXIc0iGeQFlU
2cpm1tNnpqG/N+pKEh/m0KrQ8nr2/WfmBGnjofD693mOyPuTaIuDGhspRT9cfrhgAq90KXwl5CR5
6GFvfwd9NTNTbuGePsMnS4v6V0cTu692LvcJGmogyHRmDT9OpmlgGcfAH0eQ059082ep6eCAaSPi
BZ67k8rHDk21sjtbNF1t9mGOPyByl1hKR2ANpPZBt5YEslUbBuha7OCU6ueDy/JVz2Cf7JSJI1Tg
Q5KOl69Th4UY6ayoRGHbZgocvwBHZl144wfrZLcMvLv9hZKou9nK7t6tYqYzfuJUqEa/cTUBST1f
OLR2G1e1SNKlkn+ItMjTEIaY1c85ki6QLfHoNpT7KsAZohm9hgDA/YgISHtKNgrHd7tjPAuQZrFA
GoRCX8sZNXDZSurqK+/c3jgFFNvq5stem5SNriNbiEWNy+em9rdhXNNl/ZsR82zsvaiiHd/ky7Yj
DP+7qhWcg+Q6UyRFkC3vtwaLT6IFoTNq97Ctlr+3VtLCGJH3U6lX3VDyzeqVmmt7Ki0nER4Af7TT
MyLBqbMKnt6aL6iVMVDK4FQDnGv6R77oiqdlnfmxBs+kK6a3aL2+sX97cZN2DcBnlDScT/597MfU
popR95G+zVXkCc41ZqLVN+bydZkyYIV1Ar1oTkWwooPVXQfOawm8yUv4ncRNlbBCxtKI7HevTq+l
lwkpb6EwDTRYpNWIh7uYy0YpH17lZ1Ua5UUvDKAXxZBiWZLs/PSrvDRV6fuI8Nnq6EIXs5dvtZQf
IK7K5G8yJ2vTKI155sORby+wgokfVjcKJnipu1Kev+4D9grzG0nlOB6lhGKbC1PksWdBRekEUZFV
5cB6Nf4tmU0BkCiXsWxWS527YfNkvkK6jfFsvOtLtYw/bK7UuEI9qpxyoDdQ53tjlyvoIxN5lT3T
ZxcIiZfGulQWAg8SzrIf3ZWor6CLpZdyX0t2TVuLSCCYh2RrB918WGBXroNPaC3XNYg7H052aJP6
cuJ4K/VK/buprkP9kUmAlab9MbIkvirV/1ihnPpOYctELsb3miQhX7nJ5KEeNHv1NKQNwsS4kTto
c29C1+7EOnp0eUqYa0O6dUykqB2lAVX5iQTy65Rn7xbqyDva0orHR4mzF8ib+m6u2VCNPga3rApW
AdWSJy0d1PrF0giPEoNbJ2qG+1dmd6HJXyTmDgU2m8rrEAVq1pueSUE1WDXxkL41ylmY0V3drnm2
MwOz42Z78noK2HEJKy9hhYpBNiaoOHHy4WNkr606MPDD5Cgu3UIMxBaNzthtCmVElQ/e2nnRIk/D
G2V9y91C9OjgQ8QaL2v9uu+0AyE+zMaDVhAreLNfqtpJcjTHkg4kqWVqzJ8Q28hscmEmhS3EQwyL
TDGJ1E6SmXWms/TgBHLqG1pTx25iV8V34XGc8oFF7fDbKWxEehxbVATk4F/YYend3T31FIEqfLo5
JP4TuJHTAdyplMDnrtWTGSV4GgkUyYBVWxWXv3UYICIDSqTsrAAc/I9f9C7pF+ROWvu7VM6Z7mQ7
Re4y0501kpRaWKOzhvqurjUqBT/man0sLYmIcJOJd8ns5EDno3RUV/VGPLjlnLHpIZ0Qww04f55S
BszL6dDVwP1xv15XXud+Mhq7DM8Qz8MbD/0E4UW0x16YJa4xFFs3tGAYwVmf6Tm+ftje4iVrms/O
lg52J5IjeAgKmsan4O6aL72v4P3fW7OX7JeuVDFJlmcSd5mOZn3rUyXeFqpMBokjejG1VyqG65qD
Uk9EtZn8x6IKp3xh30ApBG2CjAhwmE8/ab0FtrCbAOHgynzMpORGzXdPhKUVlia4cf6G7Av+8hLi
UkuwWSA6m44XtOvaKu3gPj3Dp5wvrYE5k7Z2RTJ3iwCIgeDBGjJkar7qP8EjVi/8rNsBJKJu+10E
Gaeg84hAd72760S/LqCoJdgc8wCfaDAo1dHdd52Oz8PHKV0Tl4zoxhbALiNGVaW4lB7QsTKDj7HV
SwHyuphqvFbqKlWJDY6x4OauT/3LsaDynjd31+4rq5PbJXo/GyKuxqAetHEdr6AjYeeMoO495zj6
jI6c6y/fXt2BxM7KmuDnDUBT91T/5dlWy+AbNRZ5VxeY7XPX0/1r8uArks9Hf1WsY8eSbNGCxQjR
JJKd8712eo8ou1boMqqPesnwfwPVOqJQ+W+YNCTHfF2BDviPtfTNtKtOdJxS2JOMerMG4pLpZ4dT
/WmAxLgCzhnkSMtD04WWVNEHoPNZ23LZ3pXx13j0LUykpPFAwUeBdNQVzCs7qXDufLE3PdRGDu8B
81OpgDSKfUvkDBaRZMpVrrNDfyKpzwCeRLC7jEbNvxvuRhiLWxxwV42izdefZ0MV7BmyKByZKEgp
vvHjh6CxEFSf4khsUfkzcK/RG89r+hTm6/TX5aVbzYPsKqDGkRET10LD6FIMIaGczMBAOn1uVfex
M1MscipmgkLAqY/pWNbVriKfF1RWjawnN67okoPf/8N58ua1eWgbCYM6zkGbpPXyrqQacHmieM8c
wpK3h42PuuzqaUnCii/2WSvwDooXFZ7AWLwOB4Q1N3CZUlKu1+culG/YGxveY2JDef54sMNjxmGs
FxhG/nmJ1/CAorVUQGIK/AUL/3+tka+lSYnGB5pPqVkGDyAwM4meaqilQV9qKgmwauIzdr132OIW
p9b8WBM6JmDMbIoEzXEKilhSQD0hcuyPy1mNcJPnnTdoWKwV3XAb9Zhe4qosorUVq7L8QsZEEhfL
40Ewk1mpkRMka5mZDw4ty8tzsmFWiZ0e09qiyTv1xyzbnuTWwClrbdELavgRJOWCDgqUKsdckXiw
B8+bYuSEv2bqzG9UXu5DIT6G7RpQb6RWy20D0aOR10aIC3/j+EePQxVlz1LURGZtgGH+4K5Xv6+Y
2t1vcjl4+IMlM/2k4UqIc8Bx/6mfHbRKkijvBLQUUJZYXzHEbLEk5lSoOZpCdyLlNv3Myuo6px3S
+dUwamt+s/4Pifaw3/AZdfqNcj7E8nKl7LEBhVzpVEVJmeasMltrvdlsc3zneMAtGMiF+9xKpnyq
x3z3PyAeGki2AAEwBZl8AJwRIMITTnxvzhWSJO10ueY0eKhPLjE1ZvVhmi3I6t1RKpuvkSbgPODR
LaZz9nE9qNhTpWxzk8JGsOWQ4SQtXmjXarZLFdEn5ox1CIJlyOoBhz0Fqf127et3KPW97LFkBcqf
XIcRY8IQTbzPD1kUB9FTigiHqqFpqEIbWRoCvTZglVqQkLAMgkC8bOahwxegGUnHXJOv6wHLXGYn
8c4ev1Hqc3TmV/l0B+ZBlmGL815Q0P36fgfPLjkfoC1sr+/1LYAM/szyJ1x4QOIwzlmXJkke05Kt
NvMJ1X6Ty+TI1xsQ73jQfz6XrtxROKIHCphE/nr5p0NCOZ4npDgc8FaARQUwJGUR6GXKGUJjinBn
ZZ30nR1X28Z4sTgqK77d/lQiQC+rZxjgZiSRWGTyPmg/sZyp3T+LKmPdWEXAE1TnwuANbGooZYos
ukPq5PXJW3A367VZGy0rGaIpor19+iRV0ioL7Lg8gEb4WGIgZHJjnVuOe/82DE8zkIUx619pHv3d
5PbntUUdpJGXLxta1KOUsFIv06yFFfZCT2pOmlma9Eb5OcJwnqONnrHUlBbrhTTU75d2S968UiCB
Cs8yu+lp3RwAjDqvANCO6f+vr/KTFnPYwPnp16Afr9fHoY/EUqped8DnB+FDynCoX8V7+UMHAN6o
Gt6sDFFSEsUnnt2bHaK/xLuXk4pfGhEwuJdn4rTrlK9g/mKTQ+7vdhu2rt0t9kZhEEQFdZ39c5uh
HZ0V2TyLLjtjn2kjRVNdUaynRsw8COu62rjSpP/s+MQDdocr/YSisKzLihB0j0hyr0qGmenJWkuV
n9bUsDu5izp5DadL24IOzdF9S+IPuSN8Zcnk0seoCZRp+MMZKirnwCTEtPARFC6F0TH5EELcTF0R
7M8KYYTVpGse6CCIM+0mAqtX2Psnvr+I+PLan5zrkXxXJBEb4OKIhV2NAizesAtGbA+j6WUcGS1K
aNumJULPX0T4tzK3BFvhkJ1o6V1k6thSw3rd2JIw/Gt7duafoN2tBpAoiRc0/9pM/Npz7oZjYjza
JerhEPltUuEcV6MW55E7Lz9Ayhm6+l7WGnx0MzMrYd7pOMK5kVEHnVCF/xk/58YHaYekUNAxSvrJ
5ImzHYGzZ67ra18C0gpuveFASU0c80+8CMzxjRe6Y0a/IPaIF9FiSQvDnuUqD8XYmb6nYEHcW5Xw
kPHFwqP+X/FPBQU5dfwSjz28LnTd/qAjZeewM88y1lPYxWsgLIgZqzsMorvdpTiBDK3pL8nPbfzD
E2/7L926DgFJbRK9biPwzU9bww9Aw3yZWtIezQ/fT2rxhX9pdAAcuI+euH1uDhDb9bzXldz9F3km
TtrUIC0gvzhLV6bHYRUCgQDT9S2jihqaOLrBHQfbX16g3RvsAwUN3eAw4baFxRuAnEQ1uLyr5gA7
mK9ZqB4e/Bi3NGi6VDCk7QkbnWfNZdiLOxolba1zKMppA6G7zk1YYzgcnZ9aQ8UGyYRM5LN4HYvU
ek+zDtnWzQwqRosc/pQ9wApbiu9pbClNDwPTkafucSXUNK77volTF/9CKXqxEDJHzYczR52qR2eF
lXdQNT3TfzHJ6jqkBzAi31zDl0oMlNAh9fgX+XeWoCJWgzzxOXxVaIwbWo3UFVUe69+09Wh4sbrP
+EQPGuv286MClQyFTZhbvK08mD/4nwGp3yj0yi1jzrVEY9xcGHXIv3FXGdqhfBxLSXCZl2EEiedQ
vXAl4JQqS7viFBMpnV6NxWG4qIn+P/ajVGreNslY95MAyxYn/Lx0F/NrwbPt41qab7U9hFDiXrIr
c1I5pKRIQiO1B2w8W8gfG4S+Ztec4pqbB5ej9M5Yl6gnZ6haVjGzicucg8bJPPNcUzP45Y1yQ7y7
yzTZNI5CkjjaEQfdJD2FNNbZ77kbx7o1WYWciRCkg9NRZefkB1DwEIQJ15sMXxsS9OtnXQaLZjk5
7L7klDxZgRn4YpA0G1D4hS+2DwUJ8QwvMZKbeyEIFE3ASWgUyCdnTc2ze3VH144ZVQfggLASE2f8
AQiWn/uehUsxZ9nZ8QY5h/ypEgZE7MmJEEXnxkr2x2ns1d7sVPvIdUxGdNdtXqErN4JBTDZJZZJi
mKoDQnM91WXo3WqM9ZgSIkmjtbcLhqhFWwozejwjC9X+j2dweJ3O4+6Sz/bHipZO3aY8+WkPLtFD
H/R7MfOXkI6B8fcrc8uA83qAWLd6ftgq/o/iBnQSPL2lUd+5smMQW/RAvt8Im7wF9u6Rl73iA7fJ
+6GNHurRCYCAesRdy0JjHMzw9nMxfkRaepWZYztiyjEtSb5oxAaztrptIJnJZGTH05KCxHQDthk6
Ug7O7yhuDmP0IeLoXWXFYlKzEqalZMp9xESfwAp3+HnSCOJEyUt6sqaaZwnRqYhWyO+P4D4nptib
3x/h9IxD1bwKf4RgClPF7PZ2p9WHFH1Lgw9Wi0MxX+nlI9U1xv9iz5YlYuOjaWIkqP2qNmvyjhZA
sMbErCfj4/YGthNS/uP1D9HdlbjWwGqLgZWRA5FdbBONVfpOgQLL1OS+tgdatyNnjrddg4PEILHt
exk+Xqb7EII0THNpIXZ8ORWMITBK85C6Er5/p6IQCoca+neofQ9f0GBQLJonin2mfiPIO9LfOFSd
j6d2DWaq4SpMlOW9CnS+f5JnCaQqcrAQ7Lh87HgL9IBfOwgkzG6eIMGu8p0rxH1X3KbX39+kyRUc
XldYre+wDoYeXbZSabr1mo11ohf5qD8jq7oUQA0JbbGmsyLqHsMSpxTOYUZs/m5oK67NZQu0Tylp
+yf3HXh4Lz2N4zVSK9QUptb4vPnADT1j7dHW6I0udzW9Q6S2s3JCbNAMXL1B/8hA2v7WCclUM7AL
a+1SbFyOPDanRCl6rgjAvl/TW8Pr+K6x4apFDW+SxfSYVZk9rVVB/1TW5A2oxqDwEy++D3Mo2lMW
pBb23tjA3K7X/t7jVYr3TS5zD0oEFqrCpV/rGJ3NY2jtMazDUt3CpDqKnYAYkBljZRFxkYVPZIzP
1KDF48XYQzEay2xSWHH8V3l2EKEqXwOwfWvtXHEtU6YT9iJX2xghj6SD/u+uphgYTkIJvKK0AiZo
FL9dPyXq2vrzZ8HIAxariBLmWey4DCeQo1sHoQerZ0FEPsTqxZXlyPRsQYBLUfSCMwIuvM9BnkmZ
5JdNuL7KAFn/9YqZlWa3eQzjM1uUNKggFhEjbpD2KUGCOb/7uc7l5Dt6V2Q7jsKwMx+jrqGSAIWL
hFvAFozfwnfpprkfmekqij6cXWXTBaYgtJTUuTaUs6I30ELDgnfdDSxnsXQuQSj0kXn5ytApNGXI
lWb5jJK3DpKDjQuDeMjb57rvKwpXOWuR5R/Zh4yMbuFwQK/2On0mAOdpfCk+wjLnLy85Bh4Rs+q7
2znKY2GRtDkf8XpJfLL71ceiYetw6UmN9mGMXAE+nS8LX87qFXHj9vtL+hWCLQStES3u/ySCe172
RSKBSEHx+81MaeTY4a85X+yQ2lPQoYK1ajh/WJvEK1ee/FpPqCcmBzzCKe5ngSilMSTseeQDc3w+
24bIvzVlxXxe8pzviPsvFZwnsR1LnhfAzE9Nhw7yjCfQYOx4RYHhN8sJR4fZxBuVNaoIC3f9JuEw
NjzVu99aiwapYPwgcUFc9Ob5P7AsEX21bbT3X85jjcCQIXzF4IW2nBO3kugcHKAnPzhJK3Gt3g4b
FV5ph2ELAZAu7zhZLDDTchGpHc9ZQXJSARK0Kic/lY01eegSPWgZToX8JTriWk+DdZpn8O3xGIpl
b0bT9Ei9BJH9srUwFwS6NMgazns0e7NSOKQRxwX+Lw03BGPUAKg6AaITe7Y5FCaVh/axjHy5isdU
IqzPkqT9WJ6XUXg6hoP1L7DGnLVtvl02y7R/aDg+5UlQ+64Mim9jwh49iLuUEvk88tgyNv+0xdlk
CSOqZDradhXWCAwkLSaDg2YgUbc36agfvFSVK0NTHCAwWRwQUvfmZtOmbM9bfUs5hAKPDm01zceg
PNjiUXwYh2xaKFtgveO8KHyYh2fuLaVt5WFYDqlv46c+Wd5iUPFRNVFoF0cKibcpScXVH3pC2FKE
D2B2zDdYR/vKFsFw+aRCSVATiuqH7XYDpZeWyv0omv7r/cfTG9QQSZXHuVjIfBd9ag1y9Yy7ONyq
A2iOPepMw2ox8sdwHw6LI/TPD05lsECCP8DJ4SQYfRsIylyCUYUb2DDFePTAyjp2+uycFkcjxcFh
vf+qKtPGqhy4a32Rz2ns0Op+9G6JXGGAh5XxYTFBhnIyx09Fsupg0QD0WXlASAfHYjtqSPBJOKFW
S1xwkQGZ/Vo00ZXhM8aJ34yYhKi2+I+J+mk/F13ytaXqVkiDhzI2sociM0nZOlB/7LXTjYi6XgVb
HoKpbplbq1bbTkV+dLiP76HQf0S75H1oSFO/K3a1jsepBg9ipF5Np+wYPcw9SicmDMFNm6Seo+vX
xz/6lcMyTCnCyUlBH4ze9lfGV2e/Jc76bP14Me5tPZ9VOGiq/JZAkRB/qNaceh1CEXQYUuLLhnCN
8wUu4TJP0hztYavfPmECVnXhbwkk4987D0rilVJPlp/JklPZlX611am89dzlWF2cWSB5BRkRPEfR
DP9Q7H73zDACSKMU3nXrrjW883aurpq4p/tJyiLWmr4Ts3DPBps2iaUQMKjpDltH5NRl8d2CZVmW
KsYCyme9kGyl/7XdA7JXcZzWuFvfw4HFrbrkZGQKRvcxRy9Qg/dq1ZJc/zE8lLG+An891kC27/Ov
DZemGUuWC8wBtcA2U4no3T16cCm8x10odxvmiSTlpthhwBYW9lWKIWKYpuOPRG2aUldlhwg2VSGl
JMi0MPApIQqWey1UGYDDM5W2Ze80FAk9sgbmMs4OlEYkPwf5mKoP1K+DTaoe9rKc/iZn6BAlR3tV
AYXUENOV1eg2bZtgDR9wKumByifioYnhMt9LKb+sg778o8VAqjiugoZqXQ9pb4T7lA1KNhKSRvl7
2cuT2wptWbIqbF613LBNOD1cDDMR9nCL1/s3EX7ybQKsCHlx3CmKqSan+H0UzWg=
`protect end_protected
