--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
OlBULwfxdJTTD/3rzvj6QEiQBDYei/SDwj1qXVAEdVvkF37AEZXXNz97x3D+86jWLfI2VYQj19KD
rCKdh/bXFz2dVuuACLt+GsSG38T+Fs86M8IvP1QgI6WFWMo4Q15ITE5Cg66qDVx8+vNLAVFy1Qdn
vRPw6mORDycyfgtM8pmq9YI/96T1Yn/KJfyhiL8D6yr+2pFGvvSx4qVokcm1xiOJ2kRHerKcz/7N
CKEdOnGnLZg/uW3Vjy9vcV9OmNhDTJueWTznlLM97uIuFn6arHfMywOz9/0XrLMf0hI5aaLUnnww
mCwBA3/ypHaqphpbH3FbQXfoMxYIc6QBTUtpWQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Eq+iN9PD3kGramidB7B3cdEBID9S4a5ZxLNtvYasXw4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
p46eic59iNI/aekmKwmvM4b+q8oAS1169/7oUPNawg3T2g/ldnC+UPcOq0NIBNsknLc15mlkNxnb
CbrqTpIPDOyz1DJ+T9gL0LWTfrAvayDrPcqY7kO1citBQ7Fz/MlCs/iC/BlaewKB9qhz1Z83GzRj
um18mEgfHx9VcfbUYy11A+7A6GNprgEvJyWf0h/76JZqk7vPLjXJOuHwicAyXF/OJOICe8EMrXqb
BDv4haWFIROGinCeV91nQBNnJCpERPA62gUqcOwKQCPD1DrpX+Og+iyNG6G8/xELAWBCDZDGq2ts
dVvV+Xgn9utIsazD/6eGEY6vU4WWtBPwEywOBw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="TsvkekuEvKlZuuoW7CDTqwuQaTA4QEDIEyttVkCmHf0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12336)
`protect data_block
C96JtQdchmYLtokCYXI0Or/og5SZYQDnsvw86uoHSGOoMMUkLLhN0INBvrLCkDbSHsos1mordAuN
Of08G+ciTKbYjRUB7/WWqf6RMtR5YcfDEkW9h2IoYZPhZXXCHorj/5qYcBn02RkGhR4BIi5y4UJo
QgduOnaznlrwvu+wxZ13+D8JmHZ6VDKtyVU4zWH9SpqJVGiuMfhW6AQHZ8NXdtecCcOAeqvDoKe/
Uih3WcRV8Vpb7BJmkQWOxdFHUCZ45bWnXk1qTF6yztBaNb0dn5cd1+bjx5mseYhHj7a/nhT5QoF6
IKDgF6LV+3NIZnMqhZMtIhm02ApJ27MIfd095gXKLjARW/yie+DO+ljC1Bv8vQ/dzQ18pqcrAuLd
BeBwybQEizQBkd+JV7Jnc9Il67JPk9e8aHQBnBR1VL+JuoXnOfcC6nXvHJiEPL6cwGJ+ikJSqqXt
HnlLp//9r534cLgL6GsovAt/ohFEmE1y5Z+u3ic4dUyMnlDEW/IC5DZ3I97Ff2ocvw+b4qcT55qk
ExTcS17uVYrOqN3U0zESRKp13JeoJxcyxw4qo4BSFit8NnU3NCkMoGreval/Y4bfbhvuNmpack+u
Xd83swLKYsGnIZaq+Tdm8gB4USYHH153gXBWoythM7Nw+rcwwjxqFGRpasFO/fYA5LlRhkFj0ins
Ih9tSXucqVzRgEyGUPwUbPhai2ySQAUKy6gqPNxtudC+u7NToJmXdr/bfspQXx1XsR9WgKW0BwQG
8/XFnEvnXWkZ8w1z6n3pN+TatZtnTKx06TXrLgGW+T+hxHp0zezlRAoY1pNjD03iX2nfPYNralPC
rO8YbNBHy0rlzRXU7bo6vzxsRO/YuvTicDBAqiq8Qtba3rIcp7CTshpJdawgfAu9Mn4Dnan9Sb/n
0I3i8xOWUTZUxcXobPNnVuPgdyukUvTaLNxJOMoowCyOWWsZaUBGRMNUcLqBseEmEAFaLuNZ7FYB
V2AVBHIkcrhu6bqSvHyIIReCxdazBejZocI1FcWmYL+YDDCpZoiYq+lBCatbbzGKFt2Zwhkkimjn
unhp8PYPkfQ8Rm9DEooh/jwCQexz9jGH3huaSZZxbnpuxh93OC/8RT0EwzdJEbgayDCOF3I/aTeg
t2ORr5X5sAh1F0WFDmq007fBI1mpGl06QEw4jk6wH3eNdxk11KwzxaON6+lZ4lIsvbBaElFXRRJF
8JmFDuk2UsXNP5SLD64andJ7/GUABGuzmf+IwJjSjyYuShSpBL0rFkc7hR0Uim8DW7p0TuD9jQvO
fpbLLDDQsraFlkho3dsywCNnpYzVQhti0aV/edqD+cN+aWQFj1FjpCeUz2HEz2TV8JOE+/jC1IsO
5s2b1GAHVjOY4Q6eg0rkWnBvWbm5OaiWE0UEwLZw3Cde5IfeFFW8RpB8Muy4+Z16S5YFr+cNKVJL
IL8uMlVkp0OtbzR5t/S+kUpGn6cvxEZA+dxbdGkZn/PkcnRA7qQAhOja+xI1Go6UeKkMA4N7AhrN
637W5vqdKNgeWHAasZU0yH4yAF+a/Yiembcyv5DB+copDrL4Lha0dzbpOgOZvcUGb2HASu2QNEXB
tpPBuh36saMg7+OE60CQs58v6735bxP4hJ3+FyAcny4vvfOtEkgL6GeGuQBuuVsc4N9P9Y+3SWD/
wYuQ7ojCT3y3/3gFJLIj1Rsxip8Hq8W5AQdh1vFkam0WiC8+t1USvx6BCQ6e1O54Zp1+xE65CZoP
WyUXmzT8R9B7ioHArvZ13c3l+jLOJ9G0sNm0J5erSfy3R9uAsceKhfEy/megXinxyAu3T664UM/P
08Ma/1yMPzVOD5I1b6CReDVf87HynsqMpwWxyLrvU8/rOEh5R8Kqj2CWwKvTfaN+CGATU0MaMmzV
SIE82SptyjlAvwejOvZq5iCVK6dTef4n5ou0Gh1wptMr6HVhmX5warNJ+fpJy2WHpMkaNIibhfLj
Lo/eGlFBVGjU4B99yT5NfLkN4e5Uu37lcNxEYQHY2i49Y3PK6OmNs+pTpVXZEKwY+tXMxdE0r6yK
Ho8kL90E8grYvZ8DSYabyvrlYPvgP5NrH1VlSFzNx1yc8ZCdwbuqOSrItqRogNHYGq5jw0ryjZo7
D9qYz6tPtQLg6GZ3Zh1uHn3iBXu5nw4uLtijf9dAFEXsdvSnkuN0EsQ2C/z9WRh40LaNeJTssiDq
ulzwlvNzGE6f9pWZQSUG8A05X2ZyeaNIa4HiQlyy1AuJi6X/EkEOA6DnxkYiFeEH1IfxipTZLW9w
m7bLAp1FQQvsBWnXMOLDj4kBWTas4KhYGY7Y5kjcsXCyVw5ajMZxBvgqrSnI/oaaKXHvcW3UdH0e
+Nd8cwHIhKd36yRHGsvX4GZiLmleWWo4x27qSrUoDhyIK2aoZpX5mDmyeEZnp6toAUcIJ8Sw1iZ2
TANdRfz3aK+FkLqTHfVJhnHWMSADjQzsMycNVE5D9ZH516VOqSso7QzSpy2H0DTBsfgDHWQMj4kY
1tj6jFeplVM9XTjvlDLhJ/L9XIKXQ7BWo4ZEr5clrAvB8zGueWdIwAqMwnk4PrS7arKbCYgy5aft
t5Y93+fA0rt5y1fClRBrjjTBgcaq8oszKT/Q8hfy56W1lCXGh07g/LcX6GQ4dfKtXMdYvCvlVf+B
y80VLCARqysFItTrwJeo1HSknxXHUxZ+J1t8p2pkeHfdzjih8zK5PHLL5iZw6guY2VBrqt1mIxGr
QF24YiZA18y11Kw6Z3vXKgY+hVRcvLUdONNm5bap8IoJCT7xO0I3NvqT2LqzlXQpnKqOY5iDE/gh
5IB6YWd7ef3akKJkNiZC/7C1cr2lxd41iLwaySXVABUZ/+Noqb1wnbXAIcZ46/3sg8ba6T/1MA2c
zE9236sNtJgkScn7V/BbW4idJW8WxwbtMrrgbbS+vMJ+m45rAC01RvXnO0JTur0pRQ0PI+Dfb9d/
o+sC9k0kVOvZdcPV5jKSBezfQvGAuZS1gGnLvMp37txT+tmibcMvekjWYEXmfVlo4RQkGlVSKBWe
avtdxdnq4JHLjx6X6zO0eHF3xKOj655KeVmmb2ZBDbZI3/3fdlY3BTW9rOsfX17BNFXLhGF0pxWL
yVYlHHQitNWbLuId0tWF/a/0oHAlfmN6ll7aNAlmEzo4oFd1mh3iYgoF6DSw5EwSIzCMpDfidLIx
ijlTd7KArtkGW5vzdIMRBm6u864P5GHulq4s8eaiqOpBa1GXK52dn/eYmtRIt88wWKc/LCyZCj0g
EpGlH2a/H7rwp39JkNS4dDrvfRATuivFpPk06fkANjr2DxoiTONT/vymNJrpz469uthmKxKVLBh9
lKLrjpFYPGDF1uK/PikUQ8ckEiKwPA/ckzqoRgDj8hv3Be8AbObouCNiItULmezKVLPeL6PyGDvA
lfwzuHdfwKS+gE1ogR7JfVWIOkmvAd1XEZYXdaJOHTq05h81HHKli7jCpG2ZhXV1JQHhhB3KoWcf
g7jqb1UJThEkyTu2H7YovO7LckV6FAtQaBU45d96GJKjl4alrnqD+TVGhmBcyAcDc9gyNulvArHh
6apbJA+bmMXbe/TFMEVS5TP6UKF/+MYznv2SCrxChJzt/R5KIS9NnzzGJ+E/yIly7PeEnK8+ZFOd
ap8yb6vf5v7N9xuhMF4sd5AI6ttIzIQ5ZIfGADRnxFN5FXSLKrun3gC0TtXsj4OooHZig45w2pCh
AulZHXpxzg7LqT7yI046AAsuiX1TobRqPxxwtEnodT+ePuo1stISY7SqLwYt4R0rVq3uxzp4arIm
3mTMTM0z3mJwZpt2OjFPHckjPMEYOltShUaeb4BdLmCYpMHsrwd0zKA799ctY8wNNNwutsGKlY0E
eUliLM2FLYFRf3kiBRKKLmAp3p4qE5EJzncNn76qI2ROdivIj6tuNZqm3WYYjxSnZ3/wIv1hX7PV
guc2dsVEKZ0pXbdoubM/tO22xvT6mB9CcfoxUljfhkA+cqazXHq/2ejLAr3rrlfO579q13uq8l2K
b/ePIcNjczNhKATHKZ1OiWnrUj5mm6ubq3VzbWmuRog5eUzPAhau+kVMKD4J6ksXmmWUUYxGZb0k
Nij9u97vto6OUeZTci8I72k/Zj9oroy67tchsEXl+465+GAl8//kRIGikQrUh5hVqHWCkcoVufK0
S9begwsq+QPDr1LMdK57cZdGu3Kv6GXn5rJGrPoqHENru3fp5NJ7f6PitERX5HkE1ObEy39gz9DP
h3nyXOBfB6ZzZh6O6wO4ttVL/myo7piOXc9qpnezfBjm3bged4kwNPNjnwP6YwvbDR+HygBwBqjk
XdF2Qnol8luDoFheLqIYz2ShRfHCSth5SRY6jkL9umXyJBZNFBaRJ3GzT4EFiz5NPRV/+67tsjn2
wvVUQmLOrlPdI+CJ86C5MTWr7V1yv3rNl/DTStuybthiqYxI50RLLezKnJc2x8JN0WGA3avPVeia
bgRTeem5DuKckNIEXXsdfofGoxPQNLcnvutbTVukOLPRE5IhiDqtdTpuwfF8vkjg0EkiLpDHMZ+H
OnGPO692q++TPrVAqeJ2aY28XWJ9fTq/qlj+0AXC/OpDABRtMbLRsMdzkx5LpOHY/rC5Sh+Kafda
OTB8FzCv2KmEdMU1JzOM6JfpE7xcKO9FW/0F2KQF6wAARVx4breFywCaGR1T3VuHHOLIrtk1qW8C
CAjx61Kmf1kpw+f2F3Nnp6tN6t24c8lRMfsHeKpwnLjXGzsOaAylelU3izlOZIYs5hSfaTlHa2ss
jr6piWqeTYNS6Ex6eFV56GEpPTV2R3p4kHs6ZfK9aCfwbSIPSzU+DyyKuAYEVR8S3ghk5shWPugc
u9Vsww0rhH4MSxXEDR0DpVibm9b1TqApJbKS1C7XEIxgJQHveMP8oXQzIk26fE+nnmSG/YQHBZnE
BMQ8dJu5UtFdHsgVRJ+JKWgNL1mfdgYXJP7v/0f7uV3RVRGwbXwpFiFOEYYVry4drcIi8hgWnzqd
zbBfcpCnXlfA+A2VbtsVUEjjiREYU234qaqWUbHJ9Z6uxd5RWPeZTP8yCsykY9X4Gp8eei9nBII/
WrkCfqi+dTJCdJzYPbBdmZyEX1v939KlsUfxrgUYtqGgUD+0hi8EHtGxRv8McJeppkaDp3+VxH4/
uC8KO5cCV2cz7OkJIGJ+ginrV5g5J00RrjH6dLqqrDo0Izu+6K/kZPoaHmjzxSp46POWRqU+bIuN
88Tq6G/RGEfv2bRqiuxNO2ydyTTem7xScI8vuftpViupVp+WLOpXQFnDxBTlik04j174zD/JZD0+
vRBNPg8N29i8+gENpQn8Fvr+bV8kK5ew8JodzGP/RoWpAlD832k092h4nHOF58Gl/ADA2MeqfIlk
H7reHIFAjwBndl6QlIaKNQB5zBNzKfVHtD7aQCGhO/Uh6lHqAAHytg8NJd308ZuLTEoCUB/E6wKu
Io24IOyTg7xEcBHevKGmvGaHsxGDmC1nhaTgdJ4aEcGJ5Ew7vasbYdaZBsvIXqqY9vnex4Jn12zl
Jj1MODCBmRGHsKo0YCaXOxNlA/oKuI06eVn+WVoLVCzsqVCpYVLW8uRLjs+VrxWz5S5F4C2Q0jpd
v8oOjZO1zSagvaBs/nfSu2H60v0fxUEpjzonmKdTHlzLL+b/FGUu0i7PQJXfFZCvs95bKqLB455K
ShUJTZwrpfNq+wdFJ2b2EsE5hwzHv1gwC6SkGEaq0b2+NtOIx00VuW/1XIgX2JKWFEsvzN/7OaWl
Lm04A9YGOW9F0n1oxuqFbIPLE1GAdExLbOql1iwzn+F/iiG4ljV+IX6K1aFnHmGBEd+fBtQN0sjv
UsTIufcxj3NsUa5/q/MTw01z7Qh5Z1KwPQWHpHNDWw5rAcjq+n9+vLJvHzadFBswvgUxLnYIjoVQ
B4Vc49ZSaq4WejzepYeQ+/XaZfh/mQGqHeEUGQJjipK6U25Q3YT7F4VGbIZ8VoNu/pQwHk8y6A8K
JFfMIIChC8fBGAnCmI/UOQKrQSltFItxWiVoD7y4ZE1b/oEScY9qr9EgIHKDPwdQofWVAmdc8ScY
rZcmVA/L0Umlb3YNJKawnB5y0/HzqyKmMGsf3yj+7/G9+3lIMhDhBGHNYF6hDna1cfcvllwcN86T
iytXp/UXeKV8ZEl0uPRXWkZft+Y74/C0FOLpIWJwoga+AsfTyg2GmhEgBR4nuvX5xpteiRF0D4Pf
m/DXtXWgTD6tYtGeozqrq1yK8OeZnOGn8XDn1LVXFL13fGDUrT9LiXxB8dvASpYEhyiW6a8h/y5p
pjZIqnivcl93GGkq0KV+o+mNIGjqAhNLHUJSiCQ5Fh+L7Y7kwq7llbYZs8itiXSaOLP9fGmP7ymD
vVUmn/FmFF5cnMndxGkAIYwCgyu4yWhwqh4kLCga61GnlFia0BQBUb7tIB3BFc8FvJXbAE8HAOs+
PaPSCS/a1YuJXRXiVthyn996tydDwB3Mrk/Hsb6GDaAz/3mCIUGN81gECs/omyEQkfd5meTuHULg
Y+hhF7mwLIHct+MzDIgT03gEAnZMh4xbEsi9h2YXuq9RrvPH8qjjsM11TlAauZiVaZfNYxLFxbT/
5ZA2/7/4NEMuBJqDSzlVJ8U87yvlUOa7LEYVDt5izU//T1px9h16hM0tbJ0xpH5QZED/PdYKoS7K
URqGpy8+JfOSVGPfa37KYfNOfuQ+N59OsQ5ox1bwBIqEU3H3h9BzTXWeGXmLQ/t0Qxg9eLPH8zE0
FmJov5tNEozJyANCD5w4I+52sxYQfcOIQPARLfK2ZEyCxHxUrHNTkKxJq6qIXWg/RFd7v5RbewFr
ZZusX15R6+RVt2YD8l0S9dD5OPw1YgpCiUP3AyAiC3G8V68/uGisB6oxnCAPAUemTwuFgPqOHmQ+
inL/bYzfGhWhWBKWp3FpxoZz6Y6fF5eDNinOUamGu92z6g6wtphEKXoPwxjfXeuW5F72Nmnk5ExD
qjtE3TQeDtcpmKcyZ5a3AjAZgBFMiQzsh6aurNoMRrLE85QMMvpcQK56z3hl2kwY9bDQkpGROhZe
eUBVksT3xwklldrsMqXgUzoSlneTZjRweSdI32rxSpKutyNRVj/2/GjQZZ268EzuVXrM6NYYIYpA
s6Cp5NK6utLvjbzM4BRMNJKxsHMQBAgbM4AwtliOcavdIK9y807E32zhiGAsxhP6EmvRq7yWuUS0
Jc/pWbg/q7UmwEp9k3rAUxsXxLA6kGtq4+z2I9TfrionJTJ0bO+WXjTNvKR1UpSmg8xrCtwLy47o
gJ9eIbf0ayI2yEVI51I5odGmTw+I48HqNymkVmiu9a3ji9ztx3RYeDENzSZbgUgsl3opMJzGpMT6
JpfULv2ovIyobrzVtaorz+E8/HxsDz9TxnNOeSPwkG4cakN8tS3o+cYhs1Je8OPQe+l6wc12EZdu
XywX591ovi+rhf42kYRTfwZIh1wVvMJEMei+ENokB+u6ZeNNPKK7JJ4Ew2yNNM8vJjctxXF3GaPH
yMLV6pa/8sSvzrFdsrgPY8Rd7XPekSL255nxuB0HORrjRwaC1jamnPJopJlbgmWewSNBAb+ews3B
Zx9h7i+XCWcpD41DhVK4+Pzq/zI/yzrNcfyHAxUrQmlfYRT3abc0uRVBvpUVuPKHCS0KMUIAxXGa
lSJVSzF1+fjrQUwxJouE2kT1nOWCCip4+uM6xdjNUOxlI/MCLuHEzuOA1x8Nyt+hCjs95s7uZRMj
WQwHAk90Gs0tZben89SBEZPJfOUkuzphaI0y9RCgjI2rEJC8QiDsYe1X+UZf1PsG5fAYp12f20iI
DSR9ZhOB+xsvRP7YeDl2o88nPjaXVmCcULonKSPJcIXZJqMEUBsW2F/WgiFUaUUzDtSfObn9oJ9S
HqG3dRVqCcQqhBl0KcyLNQfgDfz+xpmmOTueUXLKg9KNFm0vamFXp/NUotFIUryjkHKDsLWbi8JH
L4MaXuqwuPAe8i3hg7gdYUi3sCj1y5OjhbNBpxhauqR10JlqnW4mWgbgyn7dqdnj93uFMJs2pUGA
KUmdX/05Yh7NNPFns72kASS6/PgzvRrTHUi0KPTO/kMJQveEbqi1K93WAZB5lQAjnFqOsOku4f7i
IobZebA5w3clZSfl/afGPvSSggwrSM7Ub0WYYaTyFKuH5E8chyGqHIsEWqEmGlAoRQYrfl+NOJDa
hTCY9zNfUloG5D9+SOWWMEHf8ijRCMDJRyBXs8NTsJo7KbkyBuRqkqCoNrU7LIXqZyt7zs+qUGZM
N8Puz7ZdrOdX4fxnjyQw3qpNkWAb2XPuMQr8xnLylqbNkDHldwIdM0mhZHUYV4PyK3gs7vJnFhSS
2aO3iNsozBAIUnolWwzRNvX7BMlr1X0MycikS/xjExDYFU66h7VjkmFf0iYKHkIrnJRW/hTbuwrx
TdvC/fOKnD2GetFPW37ZPv5wZFvq2XkQIVXZJibtIeOvEW1VMdI9nR7mNjHcmIye8vrXz58WwmRk
GoWQoZUoDldktJ8X1AlYusjEWM/MTRPPMSWt38ctlkuh///lig7x0YxW/mL7tvfw37UfsRfoyJYV
attBHIFwjF/h34h56K34He4ecVgAM96SYTqjkaKiEe3+V8zKjI+3Mk7Il0JorLJ5cDPi46XA2hw1
Gi2x4c4K6IibyBM8UQ/t9nQRVCL2fKnop0dWU3JdTWW7X2KeAwPJzBv9XDLoX7EaZJT4cV1KJofz
hgvJm9UhldSq2Fp3QCb9LOxRFfGcYasDpwq851m3oa+HZHR69x3S7D53vtdrU1TvLXieC750hnGV
5/GamtaYEAa5zlqKVXHLlUQ5W3jpe42VxuXkkP2Vr+fe7kEUysz6V5TJXwA1N+ZL3zoyH4kDCCMR
pdVAJaCcoRPKMIyMrHjx5Qvra8/SmnR5Q50U/bg9LOvV7QbPF88W7AWoF9hp+ithBJiV1VhRFyQT
B0Xaw6bKY4YuEOwXCAMORL8Z//BV6Mv9EEFITbLDkL0WUMi0AtsdQRXZXpFNThdg6SUNxHgd0W4v
486ttELz/3DdMamnNAv0+0DIyDFpjD72qv7btzLGVkBmggeBOUUhoqkcHGlgrVmWcwg1c+EgnUcZ
u0RkKwN437z/EHPUed/6dhIgtdAiBEEChVNGb+vccaQqEhYQDD9Xtz8nHwmoMDvkaqvl9LjZ4ed0
ErHUJWncB+vT4FjeOV2YNhwVz6lrKhESvs2HIRIfI8SSEwcx4KRPpzP19jRCL0r5ubxEYKIb8mo+
myuNhMfkksWtCJ18rapXQBMVAWXVEx85cnkmC/nY89fhJtIoR8gpKtdDhuM+TottlWzStnkyCJ6n
AnjFcK6ig6LBht3FrmGCOemn21BvoprySaVMpFAK7IqQ796xPUS/ruXVwuR+jR8ctt3IzzIb9gau
pnk+AqIx4LPax+cV0x6z2PuQ9fcrO7FWOJHpyJhaNXdOwoV36MIGKMhtiCIBjfLyRAJPdJUy9Fk7
8+Tvy0mo3XTeJey1CDbDh6hk7NAqu4iqIkgCnk49W0plCSInpm09Za7ZCdN/1KaCgOgI8hi21Col
GB8uvW4WjMoe0BnbUZGS3qtqkGOg3OlD+Q6BT5lMkT7Gr0MyQM65RQL1vxLyctEuUDC/VR38j9Ke
zRFxinfWIFVpFx28OlCQF40VrnR+kEpYcYzOwX1nqNJUiRWFAdlFhQYCtXMfDUsJmP7KdtWPa+cQ
wa7BAbx5T9Ec6RZB9/rNunc0NUTht9S2nnFo1Xf5zJuh2TCxdHPOjxm0AtelWHfHVROR+sq2gPQ8
WTp4ySdDRgMCLDfVbkQ675ktikVHH/dB99YLixbaPj2FnZu1Kz5uDIpcVX6b5MCh71SfauMOnJQY
bOu/yGuunQ8qvr9CmdqsIIMl+OB9s3k5GSQdBFb33D/+5qeHAV9wrTgHV0b8+A4JEeuBxZQ20asb
yrcIsxLSstUWhkQ+8GdpupeRL7zO/fmInIM/D8S9Eawh6ML8lCdwsaJ2L81NmBP4lfJpFQP99GNB
FTDbmywRiCb/CaF07rDO6skwQ8+0HQmmDLYwvNzARNZnX/59hEESN/h7OiH18j2MAAJDE3+IE41n
IGXA4d1N6wb+/SJa0bb+hrDGEqwYbJC7qxUwpqLKoZUDlsaoE/rrTUVcpguFxMce5skUeFTTWbKl
PTv60h4I2nltdlWwX9mdrQ19ugMRNV1iGs0bC48cJ6GnM/Po+oigWzE6GbfyQ5bowGx6BV/Xg+k7
2VGDqvMd1hFxCHzABXb5xDFIUW1COE9wgr3SuTK6UNFlYCY+EGSAeLqDykqbLkbqpfel3/lRd+oF
rcIBJ7WCxI+/QnQe7URe918NXrG2SqSlcWaXro3aKJAi9jiboXVKEF5xhw5yDVoxHj070hbZII5F
CzfgHbuKVH0IFrx3V2ATNSsg5CrxmaGZGnd9VEeAXfakWLDlO1f2y+EBvLE8OU7/g4lTJF3KJ191
Nyz+FM5ngOwgxO/kRjyXsZOsU3tlJxJEdYxhKbKaa3DThfd2YS1rT6eCA/3bDAUMnSqIyXb14gL/
2kx/FB1fJZEwosD2QKgTI5z4CUlnycs89RUCNs9YyE4NNfn2Kc5oU/T+MUsR+PEP3Komv5Dx3iGT
rZvs9kBgnCEH5cnMoEu1u4O8nEHMu9Kc7RuTW2Ta5uNdctGSIvaEpgRsgUTDil9TW27Cl7pS0aQo
KM2SVhUS54YjRXKcko4YFxeGNEJXBk4qrG593thFQ6ZQIn9SWydzgmcppjgR8IQ9H2p+2Ds5kkqb
x7Fzgoy62zp3A3WUFejcXPrDUVcxO9IEPslReOSwmmXHfQwwtcX9AUGWyW/HTtcoEMvFFviic6s0
/kv2yk+GfSSnVi+yKrr4vlRwzZ42BaVF6DOwVA7XBZcJBA4iAZ4DruQVpSwxIXLJDSHRvO1Z6jcb
gVSKP6Uux/ydMM7smGY56mJhgLGU3oczv6zi/Xe24Q7m09ICox/c/3nsjnDFp9dw0/jJ1tDdCv+5
s1Rs1/PaaxmxK4petM0VK0/9YjQdI14KQpi9+uhEzikDe3kV51wTchA2qsTy2E51WSw67b992n0X
8EvQinrdwEljvZmPps40/JATCK9QiUgyfzVznSOefXtfHJxSzZdaX+ljveZHTSmSMlLOrGT+jgEi
q0JZiH3Blw9AUX5yERQenwsgE2p3QYKLJxqBtl4vZucPzSHuEVDrS/nP7aQzvrdJBHyXZ9o8hP5i
LnL9xBznECNwwbFOn/Bak2em33CfMH9Iwf5pODWAu4NGg+elbK8SkLA06l4pTclRNNdW/UQgT7Eb
BHwN/H5fN7qVVHBo1r7ELFF7rIcBoUMa2Jg75SEQaVzf1tcV2Goizx5O5COXaAvvs1Die1QHJNgF
8SolqYMoWSn5cNeWCLHqeLbbEIAd+AqgrBjTeD3swVlp7Y6x+KNL0baLoF0JO/nSI331NxuEnEMN
h0YC+lqqjkQBxE2yQdTmj1LiHZMpUhJH9ESmECjxsBhIbBY3Yq+kkGG3GQVHs2ovJfA4SiMpI4mM
Wqhltuyk50uzvomF7npO5AzWftBvg+5Ts1qLvfk4lrFAiwRHNnCLu/j0QzJ5CmdIZwBnkbXFAZA5
Gk6egTzU6if50p140NVPxBPSUll7aUbc6CcnpwDF0+e/ZbSIACmW3NWQmX3J6mNjB9t7DeXJTSSx
+bf76hvf55kf9NXe6Np26/1ubLzBLDAExyrnSSOqdhhVSETygC6In4Qq3+LRBDg4czs50u7o/13c
ugljWEICHUWokWK91nVWfxExtZfDe7bIAOLq6zenbyixELdVqyFhhHauR2Ny1uCVQ4R2elp3jzqT
rc5vqB8cwOkQJZc2ZXUW+g/JNle4qHi0JvLcsRJVN3CfRajrIjxTcGpbkMDI9AeCvbiiVorf3bYA
r40RxYq5QcgwEt9eNC16op20GpH06urZwTNJvOdeMS1EDgjMEwGSnyUjJbSMg4b+slHHvLbCc1Kv
rD489H6td9qrq4rBiLoPB0dX2Ff5f+TBl+mztriLQeQN5PZD/YH68+Hogrj+mXJfVpbhxfBgbOof
s5pQz337vhZCOiUlLVfjdfAaJi7qWTv8vPpgh9do/nXv2ymOfZssFq+iTqOff9w9SXFPvQIjC1Km
1ZUuLGRB0vBnDIHXvhKopnk2mz1xZzqLsdrrMqVEZunoapNV43AmbEgeFfM+qrALjm9k62mZURag
b/LNwCZrOeiITRFLb+824inYXkWsx1gujh19vnWxrT8X9MdNmp00TmGhs3SQX/j6YsUxg+WYcXx4
+wS4dlSHvLOhmXwI4J4tAcLeh28fK7KZcwDmAr5BWBCq3pl/t9HQH8yB/jHC3NaWjQAJ0BiirfiN
hkVHPM22mJgb7OmuXEcUYETHUgXilkuUmungsxgqVDV6STEDs/Irn1jkH4MgzY9LJY+a/QVjvA1O
swAaLlh0CFDqQdw5d3J2V1KnUfmeQlb/rJ5pPDWz9GJ+1Qxmw6Vmkpg79TUj6rjvimotUkvnsq3C
ahA0Dr7zrn84jyUpq0BLf6U4NCnKbH198QyuTg5a6EFVySzqugx7EDMSygM4ReOMIRzpdX8BX/nc
zwX0z8IZyk+N+cKj/J8CBU00xhUa+ulvqgWTcSUDradm+ciQVGqFhOBD8cGldmha5QyKbe0Tkx43
i9OyeRK9GUhqDOZ2cagkt/PvKWJYHnHA/yxJyTlIcOm3qIDP+8Yjw1zEdKv2RktVM8eELVRzrvSe
t7WZE5dVKwjm5/ncXvP2VaVuZZFGeB9iWRITZwqWYyRN1v8m8rLmmJbsugcGX2/HoaO1RJgNJpO9
CBSBvOk9xy20WrNMfvOwmTs7Rqx5eFnq0nQhZ8L1oTZnw7jakkP6/r77EBvEOSdtf3a5OYFGt8VX
2O9YVNMgZXgu5X+UDnIamdsQ6w1ovwWyk/do6qOFJCv7SocDkui6wtgdjZzN9MeP4kZfOlmAHqDB
l0l1b0HRd615tWmrq3n3/UU4cyGdYNI4gZFYbGxQMdfUkT+9s+J+6TsWsBfD461ESoqKvvYKiMAt
mYAGn3VLY+lOQ2yui+sjdf83FMAe+tGsRMUYqLT/1gPfIEO/N7oIBkodLm4h/Zb5qOVwaAUdEPPU
4odhVM7s8do8oouXCdwZS2lnfn8sSuv1gPbnkzrHAsYegfaj0vxt3HCo3z1WmoaU+KXepEZG3+SH
P6i28mUxkedXSdQdYqcBNCNHGI7TXM6VrM0ySWj9UkGZGBLxDvWX6F4cwBsjKcBWpH+rb78h0u92
TSll80J4BcdmdOK4AC82ZMBabrmwUDhEt70OKFrHXCE9DLS2dYscSHehLZ4P45cFNvNfS4SdGyYj
tGnj8vIUagIAHAHbZZdO6i8X1jjrnDLeJjnjVbj2ziEduiABcRZ72MIoQt2b7H3eJ2dUmjedg2wI
9EgDdDoA/tBApFHZjwtWGYlOPQO4RmLmL9EuN/XjBeEp2kywEV9ZA4Uk4gI5l8bMcg7h6gc1RXHo
MUSgWZhh3QshR1Gt/ZFoFh3nXuOVm/f8XInEU6Mb6nBwruwgAFO2BNX1uZCW20yiqofcVEyuOsOp
VnxzXO/uUYotidVD/uSD+qanmRvtbQSQSJ9aTOij6YFmHGuuES+JlgF4vpFXo+xRwSr8hwC4VFIB
l4NJc6NI/w9KS6PhgAxZxIpg7olDGNByjbDmVWtg6z9fWgPDwcfFOs7JxNitPEg5Stmu/8zzVIS1
ngiXRWSe/iqYdEd0uuKhh/n9xx39hm0qzB/qu5ERuu7HnJhpBxSOtZGbOx5umpkx1uThNoekza7o
W8spj4+OohzG2EGJNuvXAEm4tKmKt9AeeQ2PrVZ5k+XVZJtoQPBUy5hrEBPDStdVmmtmK+ZKNm4G
Ceji5U6nDhNexto1RgZUpjE4Q1qh7xN2N0pkDsyfOKEqcf4DKNyxAefET8pLeAuKVqvAoOTGazPz
4xfsXjdFloBflYhUHbiP4M0IqqTGVHbFuLrRri/5fmZ9AKKSB/LwLfci0ogW9u6IjuI0VPv0QoYe
e6Vtxs/v/lOIL2hTETS1YMdr6uwitYQeL3cIOeTtnhOufl/qC57HcGMKvafpeN4CUz3LwDxG2Ojv
aoixGKiCbyUYl3D2nbxe3KeMu6vLMY7RU5dian1oaw9hsRq9uUAcCdt16RQj61gFFWocnTqq6V0r
4Us/NVCiG50aLaghC8SIHVzVNhYr/7F2AiGwCzBGjcZmsqgcOKdSr36SSjFintltDctIcS5M0HwY
FUA0nbW5Z0yvDf8g6cnanLNjIXNxfmd5Gq2P6bvebAQZJM2NgAvJYdr2x2fhZnhCiCRoLEs77la0
IMQ5IChxX/pMNN96Ko4H9bwy8ztsSB6S9/ltUwSikFd44HDKIo8KWTK4u7nlILtqvusSc4XZStpB
Rkf2zed/qN1XrO83zGbXW1q5rs3RFm98T47e9s98mWcGCZ9WCvbDjcuCe5VmHKG+lOE2ZnkIDTww
Bg2XeFg9Nxryq3XZ83i3hYFfIRiddLwWJbLKcr0BXCq9CNQSoDadzbIBUii+114vWrQunGvOkWUT
SBQVeWQCUD27/ZcWH64GcYWbHJuaVtHyyBRTwf+gRYk8F1oDYC0p+JvLBdWncszwDYuEylGe7K0B
2K1jwDwmQ5Pf9WsNyefULJCaY32Rbw1CNpxSfqevOqSxPbaNBu8n4O1tz/8/0UyBddsNewMZ/KmD
8dSxvY3DQjFKIaRecqFetJ0rOTxEQLo0wctpbvv5NFVHGMpi8eKsNRVJ5Wu6cvyDikm3I79bS3Le
SEulJI+Uo6uzSdaXtDee/AAZzJseWJ0T0m+yrwAmNtrn0wGZOCtddj7xAhcfiU6UEWSxeT8k7l3g
QUQByopASynGaofr7IZgS/TzzuDJS+IB2XGRHxf6vt2RdUWYq2sFm8nEdd5X3TD5lcD2tXQwpy59
iVSAQfh4atg3cK3f98/kCfq6XolXKVmAIydWfjGtFQsNtC3N08opuOJhMzJK+IdS1BwgjGPuCW1O
jkovr6l2s3Vzrk5gg/Em32mkhvP9ERqlFBYjxHGKD1OHctHkLZqijPgn0rninxo5iwJp2dmyTADw
S79RvRqFBrLTNvN2iwNL2p0q16/8wvq5kWwQq2lmyHzm7IX5AulyCFaVAM+DSEQOFRT9V5ZfUUE3
DeBdO4BKFL4j4K5QXwi7CqQEXTkmLYo4LqGoq/TtsNvaf4nch+e/4Zoa8W/aY1ToSlMlO8rvu7g0
5suy+zk0j18KjJM3OO7HBLoR7r1YsnarOc/OMEs6Iqh2ssqCSmax0UU/w22czmaKtirskTQcrww5
+5EgGJpX5wheXBCpCYejMasLk5DNhdfxYgucuixb3ROie1tgPHHDKHN6KqOAOz7zXsFBku3ihznD
2+BVFc4zl4Tps1x4a5YipFS5WwFoHMe6kX1II5C6gYa9fajqYvu09yJxWyGBjDKMbJMP3lKzZzFi
lJtzOmzhWt2ctyndlrSAHz5oyBP1rlrck3kizaG+f0jP57rdx/r8NlzmKYAD+VnBLZ8qDNW7opDq
x3rBU19kMFHmP2saZFSNMDgTenoyaZB9lkHdzaX0HrWOUhPC+OSBunaBNO5GC+50JF1Z1nj/Sw7M
w1AxI7FVDlv8sq3lyD4SOw/ss7hG2wU5vIt1bxx63kaF2Kzqt/3rWJc/Q8PxkbGh8hywIN3l2ZFT
5+Gcelox86HB6D+ofrA7GYCj2UjhgXf+QDM+bd1gHbLzXw8iY3JJSdfZym557wEfO2tJyP5tyqIW
ra/x370osljFLD3LDcmyIQQyftv+j0fpmn1Jkw29AKb/EPfaAhEgOnEFMEvFqmQkufi5n3SM70mS
gr3ygFDeWGpA9CUh1TYq4pgm1ptXPSM8iUx5PJCdn6Ml1k1R8oyQ3rVQnYnTkJZiURRn9iMBfGqA
ltRY75Jq+pRNkensKpaIN+2llSbBFNqdh+byYNHhZghECQkECykxvjO4M7ZERvSZRgBb01/8B5kc
aLcC9MKncFfVVvMoD2wgQ18lO5W5yzS1MYn7n7JAWxTgI+PJk33FS2eVKLZTglPbYkZr/0QNEkFZ
KLCmxirTTXA2P28AghVvkgZW6Wd6fg1775KnoMKVjH8r4YZNDsQSicWJdoqn9Zd2IsPNLGJ3FVi9
alVOG7+tPSoHa8FLKFEw4T0Xqe8xNEwXRy73UDlzoquY5YlZ+1Lp2UZigy18e2I7+EDr61F39/Sg
V5RHqwKyCmtObyh7C8wzofPbdTckrZne7KkamNVz7pgvVJvosm7TivV9Tv6CKuhyUlOL8WRcsjjI
+IRpP1PBHpAcq5TncbbmpE5NVZEVkoiYmSM0L98DP81tKHzuNtYbfCQO7d+MlhQTl2D3RFCwFJwf
VJSONfHOsZU/iAE8k9FVx6uTF3u6Svu9
`protect end_protected
