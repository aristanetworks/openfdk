--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
JyL1vP1RMjLvDDbIGaLLr9rKLz5ME8RvVDs6IwueNIdEdBxa9tlIR0gs9+H9PZkdsAh7wZoc0hWn
p9ugF6+7asHa0Qw2NXwsBl6QfygyaoxUqbbn5y+65Udl+P7SyTzuEhpAOLsqlh2VLLdW5ve7BBbs
K2yl4RYmvENgK0dgTtepmy8PzhAqmCIXYXla2sg4JqTznFmX0XaUy2RQRjY5BjrvtY/EuvdhjusJ
4E1U/ldvQhX1OeRdgZGH/vbWBOxp7z9CP9F/1ZboEPoRtB7S22j0I6BiEvlzC9DJUalHEAnYWiCL
ajPXNhgnUUlvqsuQ+u2f2nRexUNqfDZoOfTcVw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="eFmVf8DUetVQr4pfmipqC9SzzmjRLsYBci6X715zNR0="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
n8xapPQ1nQ1IJM09M6xvRTYFXllmHihXIApw37yAR0mMrw8v1If32OSnsSM4iurOjkmBoaAw3bWy
Jg4rr8qW1xWgarZfPiwBLpaPA9ojKrRONMnaBwAw9B1x6hNz4NUqxaLVG2r/4mgV7b5UnkQ4JxT1
i2dM3JynyQtAZdx8EKPwygPPBHpXF8KJDAItVVD4nIh3FjHfwFJ5sTxbFJjRHZ/jSNfCXya98wsz
+OqYy5sYIDizVNo3ECo0Yxg6DMoLPRpQOEc4RirUjTzV6YZphZewZp0iRD5rttLRMb0Hp/HpI/3S
HVMEvOQ+EZDLlnI5KRSuuRKIhIpRdPLJ4p4Y0Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="ib7O88uyEkWW2Xbb8SHRIItGWlGdLcV3sSXM8EAGu7U="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
LTMECtBJzRtT+Fv6rM97s/RzDDNRA3+IznNyNJJDDf1WzukLPxBHDWVWa9O0RxJbQhpdLLXqUhs8
oa9yYZ5ormUQvE26U9iyDeRVftMY2CkSZkulpAX7mi9UD80z4Xjp7XUT9fY5qGzQtUQBuGzgjWmC
aNUE05E/N9xmfZe518AeMip7wdpxTfLeaX1u27g+qN5g7xx+ZB+w1KrYgI2RqQwoCiyYPwlIKZGz
Je9VMmC/jUVHKP+n4YoTyQU8a51kburcjrtmDOoU582PZhfXEt7rapb2+WeijPgiUXIudq5PP2jJ
Qk1HsU2yU0oHB+HNBtLDT0OjaYUoCPDtFs74hGO5am+cyKWrb7NQDoVHfaTCRIgfSabsEfxK0uWb
WFqQ5026wQHeiLJdNLxTcqI9597lTBH1kwmdogSDRCfiVl3AQ8SuJmovm5EBH6245a4ctoRaIIlO
ALyltIcjF2/lvn1+UhgUMYLk/57+EaqYO+LAeQHzGRLfVlzq5dtn8afFNO76RS/kBvs6QIfn5vq6
HbWIBo7LhiD/kXG+ROl9wr9l5sPmmR94OsQx+kfbr9gpWIH4meRqD5zCJASythpZwftBJ39IAbUR
5vJYu2lkg5aBK9KylvQE7uRxpoBx+KyKN8zu0g980NYMpvxtVvCJYvPZ1P88XnfEKKKUa1kD3G/4
7iggTKfqa6pPsIl/HkDusdMoV0dkNpWru3O4pF6Q5rdG5VnFLI/4zLIwl2GIbet/sdvQhBbFSKby
nhBBgqvtHcuMCCMrLNO2b631F/NXC5OHdJaEIMSYPSQKTJEsOZOXcH6M7+68LnD60kpIJSeVObxY
hUZhhHJo71Nxj/IK0zoYCdPiB5F0nUjRgH3sD9rjHTgSgNcFEKbuDIXUFsmPU2u6HKZx7LCuGEdY
cXlYYsGWM3HCY5lj/skUgMK58hnR084do0fK2p1Y78ozyfU7pBnAmCWa24wUYRw58QCSp//GYW6B
77mOXNPeC38J3IZDDBG+e1q5pQXYkXVuRldww1zl0W0B6Hy7QfGOxJk8HYj3yTOrAR6xFbSq8lkQ
sHNcFPWpxa/mctjCU0l8vr2K4bZZNaxVMnNeFLxpZj3ablpCHdsKKpXTHXaiiy9Zj1a0QGD0xsXR
TneW+om/o3lLCBwnQSJi2H4xP1z/XaYWGmoViBowwz2rfj2dDWKVynXcAnnyNi5arA8yMlounkYP
cspWaOuPwgJztv1+2MlXR33RRoTwHB9+md5SvVtVW604WjVQCCYeEaR6zrit+HzFr4PIuGYrj6iF
yzWrmm2YmXTO8p9B2JxvQFboEcmlHUOpLYX+UuOXPDCEgqXULomuo7/72InsnENojKyeWcq4e04P
GhwAwAmgqA5MVXFNTRKcZbxg/HvNGZjXko6EdgR5DGVcogq/rS3zmZbv3nsSWNRVo8L5rhtfaxwv
DTQ4ZSj/QQCq8ZLbEzYmY1ig0iVS6rYlfeTcvPkBuNO/pRQdIL8QxmfzMG02tOlg5ctYzqbioy0D
advAi2HgXY0L2qC4gf74Pd3RaL7OtebVKle9pFID81f1iSSee6nHCI//7lrMHHtU6+DhHo9RB9Rr
n+2wYXpTjChWz+NwZVk8zKjxIJadAi/Axfwk1GLOTfKOTGbEiQQyaqirrThCbMewI8BENBcdhD6r
5Pf/dQKdBjKuRqsUtdi/tKYgHTYLiEJv5B90NjMP5GfUgtFBA5Fa13RPuQ9x1OZGNRK7h5kbmtBv
875R1uQIplqZW7pcYquxy9g9daHr3eEY66J0gwyRpg/IKx5pGr/5CrYRe0MtVv0DpiWvlEQSJNVB
ZWPTqsj8/P0zB5P38M9eY4G7s7mx15x25zI0aQgswFMzaEPPMu3aXdMNXz15u4bDlnqaV0OIDell
JZ+wdyduledrqO4hc8O48vozizIB/j/q2hAIB20w7yydCgHl1Ufh645OtvWfnMFWc7h4mOZQRyjm
2VMEQZNxYCyb+6Rm5TyiBHuxapLfuAghv8oo2veB2iFPO/VqTCqu67kxtyb51CJOtJq7KpOlFaNZ
HlP+xo2r4Bjy+XnnHwViD/2qrz+0M5+HTuJkbu/WfwG5NaLzp5gxtLe4ODyWC8k6Ifj83R0jhDuy
4EeABZdn9w49PZ/8XAvjhjHnbLi2zT/QFVpWIgVLRDbOC880jobjyqpBRTVROhLpAbftk+/u6y2A
3u/W9gu0HzyGS/HOV34i3U5SN51mKc6a61BPBgl+OW3XO+Eb8ZXH5I2ajb2Z6YsZ+zeReTre5yht
cX2r8Bw42fobnqgn8YZqOLnI0dytB1NBTTAdR5sVWWSkQYnJUuVW4CWGGw17gAALcjvfOTW85dJd
D1otwm/eU6gZP1PkIry6zXm0NIP62ZFa84Rd4gD4cMG99qs2NX3Wt+Z6aR7JJvSm6e0b2HU3ILX/
yBp21XD+DlhKVbpAuGMlmkGtLuTbisnmdZsqfoTQqyY4X9MtLZhcpAGaexM2UYUKs1e7f8LN0B3r
GxXquyO5UecRTPIe2Cb5HbH94GMYV3EOqIfo6l42h5sB7q1xWbbQw3B9SNJklnlSLkT6vOZXqsHE
KLkKzGlFULMnHEkqW3lq5GKi/1nzI2tPx0WCGx7DB3+rkSBeAMfBdVOVaFM83tta7B/zvdKGmwTP
wIpYe48jHZSXc52WKZvvzJZ+q7QXc9SnwR+WB7HBqngTfN/Ng3jHf77pGnyIJz1xq9kn8TKN6PAJ
GsTSMEPqh5GSe9FBwmhETEMnxwlQCL54Toj3M9eWBZ+0hJQhKubhTqbwcfVjIVnbhxi3Pwhqv1z2
nvADlPP731gkGnVu3vONlwi5D7VolrRzbTfpKcKHvOtBBP2G9sRb+IUbsccdecBlntZCOwN2MjKl
A1jLnfGvp9JrFqpGwIa7YIWh345tj+gLA84Ra+DNJr7izY4pDIjNHmT94m8osVfRMHjXsjLJGq5/
Rf2OSVirg0oGj/3wqhGdxqmlxxSfsTac0ZfwUDYgTMT36rjuAuQ70McV8rn1bcAhddnCtlCWENzR
pCEY7Vk/umrVSX9f0Xq+OpgwEtBEyGY7YBjDXoz3YZHGUtaAcaPo66ACVe8JndakgpxRnLLlhYmM
QxOKKoodAe6gV1Bx9v710v51AiG7nj3n1avRgKYVgtHhaWI+TDXh8qRQDjlQ4AEWT6dOHm9f7Slb
uhed4FCW+GKGqIpMp3lxKfHkzFg7vNEfxPW5e/JzMUgLxky0OQHZN7F7c/dKjncMFLVaZqqTdq5o
3XR2dO/8MleWav63dLACNEqWxKwaWEnwreUGzNcq9htFLtESp2E7Cba/w6YS8iYRjoOtLS33/liL
uGGrfZaX5FpJlpzk9XhEGZFnAc40ZflRtdiBF0SSvBNJCU8KPq7wIrNzgjXAXJRsseKT/W6kFW8C
4fWNnoNJBDY5cIGcpw8OnPs0rnc32NqnNmHRwQoGZyxF9LBnF/WAoSly+GKMEuXr9y75uiY3VTh/
w8YtHBjD0VrKhulGK6sH+3oY73kCJIZdzNjdE+4RMw6qaKi0mG9v7dcx+fpsx5n64FZzluBhFLLz
Kg1AMQAulXRuHpDYUsuwxhfBZdF6WORuvUoQhL8e0Urzgx3Mf0pdTqbaOH3iGJerlAbysChGUbON
9GbYBlGkxWVL9oJWtmDUIXCssL+jv+ac9HVsSqDSU8jFQujGh5TdonNkjQXMmLq5q3hf1QFZaEfK
nhok++IEE0hYceeAuAOL3GCwi9jDdM/Ciag4G9KtXkYTkyvTVGMFAOlnkCSAz+vBN0QlrzYvZS07
r283Gakqupx3HfXqufxWeu2YmnFcRF7wV05qQbAbdvaGsPs+89TwkppAGPYEEhMbGMBS0GItEqFm
xxVgZeLjDFdtIK7Cdr/nz75U9nvH/Hlh3M07aiQ9UMvCqd2fMrguM13EkKdUe2I9M8oqVFlzoR0v
31PT+unDZBP7EeQfantDeamzwE8OEbZTLCV08gpbBBFSwM6SPBUvGh/usqPbVEacycyOZxcEeCtY
9AWeszSA5uzpe43dnmxr0AP8tx2LW66rd/btV1aIEbT2Za/zadY+3bmx/AiOCAsuGcs39j1JKy78
P71Eh/VP7di3P8M935Oj+/Pp6JkNZhp8IINGbNEm/8N5gpQOpASTU1ty6P+aiRR4N0Q7r/hy1GsG
55nFDBQGHQqj8Cva0cRs0TX2mnHVO06kHaFAo+V4BaZTJxhwxz0RurBSTOUYBgMFtSJTGGU2ddd8
I8gWrJIhD9Vup6ydPzYku9T/CoPUHet3WIQIwXmQMfzPNCyMqgql6rBGWM3pWrlQcCckfFtTMsjH
fOCxbsB10YwzcF4VyhJYGFEqYz9IAEeNOJ1/ZJetJCnE4co3/U6VYnNDDCrfO9ePb0Sm4zzK8432
hk0DyYnEgUbT+meYLaBMbR54IksvyRxGEe7xM8cCyAZ3CE3Zb3sjzEJfZN3SS5K7c+Hk5SMpQnWp
gFJHMY9eTSl+ANAdFvd/SwGZ/ymfQHz1sVfCODLN5b2k8DyyWC4iG8Tr/2QX6shdXcQvy9CMsHxZ
diDgY07aAdVT9HWptP+9YeQXcL35iG4FwNdMdRpS5fWs1CsdvCPuQ9oRRMqcfaOOJnqTHbXqM7aY
MnWZKDtypf81UOk30a9paQcYhSuQHZVa5LJPClpCKL2MUkpHee12ETzDMloBI52r8BnbaNHBJQJc
GdiIyfDJMAsTchRvYT5rT5VefEcXsNIsXBYgp9q/fNkshOW5UCDg/z7KaZVJs2FJv4jBaDr4QQ7J
LxJxVsQVV8o+aOzgtw0HQMslC2M4Lm3zH5NYf4SVaDspXXzp28iNY6SxcqA17Tbn5cwMKtr1B1gf
XMNMQi1rjCBbfLuBbzA8QNQe7YtvlM6NScYRUUxgdEKyQHc7AAokNgb6P5LwDZbtRLrTvvH56agc
PPt380OIjhaX8eXXoTKzV0fEIkqc1FuY+3K8abFc0wKJGGZZrPmizadvUR1URZCIwkGQPLC0qAXb
efcuKdX/Go8ZWl+i9dqyTB/vimTuwLgdQDDfDNxD8hmVnSR6HNjqCRSs3JFxSgvvyCVa/5/nHsk8
Shsm6Iagin3JsOxJ6yGOZoEiaCW3KSZ/SeXcdrMXQaETiKK/ccu3dCkptmYHnHR6yzPuSQQouMZs
2fHomBfCA0HE5cGHAQCPWztBFYLdXOh5d6Sj6X3dN38eQwXZi2w8Aq2NdhELxnw3xLUnhATc8c9m
CZfwDqo0b8KMxZ3eHgPQktv16BRf1eQ9sMMYAc0gli7Cfe5U73v17pbFgDUdVxNUq+XRGmX/TiPf
kHtFewvFKAOX81Vo0Vu9rQ8h7glsz8kKzPr3JVYGij3Zus0Wh5OOwD3TNxi6e9Bcv9qxy6s2O8B5
Q+jyKYCaEWa90CLih5+xX8ra2BdqNFFHWyO5L334elzzz8VBkGGBdEqhpn7LchZvMZc8lzz2L6WP
A8w0/jBtzOm7e9KxyH6a5mgN43xfAxijx3ozl803J5G+JcE/BcjxJQ4SBWwT4aeO/NRYD4t6No/8
ySlNXtD1tfjrWBrlK/TepDGJCkHtaUByPyi+1nxPsIm4eq+gUQqjifvBY1vSx5e6eR2doazzD7q3
u46/QEiRrW0YXghXnmnlgi1PNjGLWNSJPdA9TT9QpTBJH2kZjFgz2LlasdqV7ctjZNuTQeHaBXol
KBF86CmjdPtiLy2mIFYf3YS/YiLp+1hIoRq50kzf2E4Z9HELPBfVFPnYyuzflvJr2dd3Cau5dho2
mC7vEhgUtmiEpL0x/H59Zhr/vRpRW2XZFlVhLew0bCvyleOBNpBrI+WDh4DJETVtMYgToFzopwKj
itqNvgNc14Z5Ki2i0b9mna0WoyOkuv1uqaqEzHdmiVzBS/fdQCC7Gt8WRKVjkZI6bPfnha9FD9rp
vf0b3W6z0HVn9WEZfQhiRFOvtwFpeuUGrjjmMRGYcsLR6V//+2PfxYWWdd/geV5rsOE3Fa57EY3V
3OGjS27LpnAr3x/WCUCrx4k+8srbJO4FTIej+uK9IBXrc+6ZdrZQh8BaeD6wBEx4KsfQTIbIM24z
KKolqBL6+pMThgRAsmgeEan5Ha71cIJITHaIVkhxnYnHKzJxeNoJr6bwiBqcSYBN50fqwDSdPbpo
qMwQtLb7is/d8HtdcRaPXaRdnWO71xnIJKTwCN1GoNG/n0pu28kuC/hHKpghsjhT3UYJ4HpHOE5m
TLQX76N5IURfgqzl+apOc3foZeNEg9xy/icKRpcHdtD0rgh74r+5rbI2p+UDHlw073Y9/UFeykVk
06Nesxxdv7fBP5iQENgO7pymEzS+BXuhQ900mfs/lDP2/oMt1dtaz/VqU64Z+7TPHm/dT43Fhq4k
MaCeb+6cmeten7MwZszxjrrDofiXDZAiCvdoD11/dVhsQKlf5eamKC2R6xlwaaj5IkAmHggJ3JRR
AZeCDW0gJ5I+JTzdf43/lDjB1Mk2tuvsxNkAJlA3OId1sRoBCzez8Yqs/xFjoWmZs/DcxEI8KWZL
f+kfa59nYl48xdXeoD8O36Q6/cWYOoCYG/4nb86yedoKalmq7iOJAnvW0HneFc+GwfbbRk+6CCRr
kKlcGvf60w5ITIvbyOtQi9AvKPPW0fWNtarqkwVNO0oiOfh27pqxwtQXML+JVT4b2+iPKKyWsLes
RL2UrifP/iB7R67ujYN4U1/63AqzxvHpVRHH3Kh6TX7IR4su7IgaGWQ5+LFkAtecYLFjp0lGlWCS
ir7NvNdEfAXZX5AHEhUuBPfKowg6f8o7q+vBLAAN+qaQ+f+6MplbRWFxcH17k3dlFuaEcu6F9X34
y3xvcXOyFwCOc4NZa7j7FUiDepnwzayuCuTgR3FiuyOa4nW2+u5EEXO4z0W6PcLfW80uYgPgoWR9
6r6JQ7HXsZRehnegzLgwzn3QREpw3g+P1UyUPL5ZYKM9qIjxVs34zLS3rsSjJmIp82htbOsKorp2
w1c+oshYIpB4WJ1SwdCfKOm0eiJ2Znuhj9JGEFToUd1m2aMVuszqY3taMsT0J6t/8EtzhbLHVJn9
yjEE3BjvjCPifT4=
`protect end_protected
