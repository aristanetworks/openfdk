--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
dJu5bqjS9AeOVf5VsXfWlOIkwcmgc2quvlKY6/R0jVycVNhN3yU4a5lritfSB84TScG1EGAN5anE
bvMXSJbNiEc/eh7xI9XS/uaskurMR1leSwat40AJhkB/5UQ+CV6yzeaGWWarJuaNz/n0LPm2OjEd
1XciXeFpayjX2UGJt3S51vnddCidEkvY/1DtuiMw7GYc2ZvNY4KdCtEcwGFp+Wo+WuIHIjkENUE2
xL6ZxxjR09CPU7mrK35C83KPyAghZ4Xo7AElhkeJFxJF4mf2GXGE8mo1bB3dC2TiHs0Ml9AtPdMz
bj731yV3AnR4yPtQUAfS3+5jkMR4dFH3oGQvEw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="QfGePeqn0MrIf0OAhj3Vpv//w8X3YwoD+k88Z4bDnLg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
UTDVVU4NMza9W3e4hiABHzIjqqi0aaubQFcl3HDwTX8LsUa5DnUN/39AtqTtKPT8t7ShlmEgTWDB
AK2UCNs37aDuYawhVhBCn2OM01fIgbB3v4r4nYJ+jwU6fANF94/efX4D0gerFLaEO1t4teC6Oj+K
zg/t+ZWOHRE6jXYDQMOwwjOBZD5wrwvyg407urpCpFnueCoXIBG13WhHS0uwy2jdVrQ11Pbus/UN
F0whyryaIJOsUsAGrb1SKIlN25MohHR4DmEiJkDm6TlPsg27P9QdsJzhHCJkmqsf2Cry6WAuyF27
FfwYvLmyRgmrTMw3kOdU9ngpAQIdJwZ2cDfKCQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="nEhfxYca3whjaIsEjh3r3Vc62Nvt3nPimko79f3QFjA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2608)
`protect data_block
ZbqVIuZe3f2rjpSww7rqFBH2+sVC7qJJW2e1mHdhd96NuvD1EtWyTgrQbUeGJhkznlePZdeDu1rQ
IwoL1wXU0Ej7z7ROhkE2raAKj6qT4ejjPaMxQPYq0FWkjcyYNjRQ86Vr7On3k2e7QJClPBMnbGGt
1YrAsCmo7a5KeSgk0JW3bWqncTY/xfYXR0e6ivbsfWylSUrHPbqEvJF5pCcdTlTiSudhN6uSia9h
vlCGsbm5kC1yoHJ6O4/f/TIAKkVyC3A3ErAJRMJ4ZWwRwYE7vH5kSKeS5QCTwW9gDwliAvOd6Rg6
Wwfbn3AxVOAnSPVQjXj82ICSFYDzi3I5xUkp1cJacaj49r6fCi7VApSyrT/ibUFQddq9wDD6TRL6
zMN5Y+0rDd2Vygr3eqavJCWTWd/V1b0FWduJpUjvcypOPsEK7aorBDUxADlyfv28jzpfdE6EfTtu
F/Qho5GbVhV61Et2+C9rpS91xItNsloLJzNpMrscIGKgWZxbhwXWuDefrgWYTU91ILr8mPsuW0J4
q1YeQ4INNGkPJTfRtacf/vw6AB1ddfkSKjqEgy2MTfdPIrsOBCJ3/7BeGXLAY0PoVky+RFiWfKZu
NYpFN3cIIQ2B119FW2dbKqAuYjPn9b6uObABvtfojkOHV7fIZQM8YgPLE5Rt4qCuqZ/L41MKLRf3
WysykeMO+96U8UX/Pphle33ieQdhNrbRb3jhd0Unh8HhSxqkEoVyEUpB8FsmwbdxXNfAgVLDjpfr
Bq3Q7IzUuQkCzUe1WryYHyIdrlzHWPYN0W/iAUIrxtrJyTPlbkK4XhIYSD7iGGCeAPNjRN86lR/u
SKadWOdC5x42l+N71jJft0b6iNWV3NNKZihVS8gPzGRhekwb8Mh1/vW6xX1cZsbXc6+8F1h/B0tO
/coZr+3vwvS1AoSdWFEvYl4+GSoIVMkNOWi2j6hJZwwR7oYFOQ4ywRC04Cq1U8l77b+f7+kAZJ/k
YJi50UzoxZdaJQLUlq0tWdPLRqH3utXPHiW1v+iRhJ33Ch4L+gAjo7bnGTqO5eIUpv8AG4nsawpQ
XE5+WD6/3ovL9bmv8CWePYYcFiij3RJGrF5OFZ7arT2Bzvm5/0aqdbDA4XKjqs3rk9tRmr3XvvEv
rHYc0obd2HJI20o0ZkSuCCml3wonTOqvbvPInFGeQBsXNf/12JpegHJqHTBN2NUisTzmZ7c1z2eV
9i/zvo78srUpkqKsxqGQfBOccBZEYWFyRHWxyv9y3DNrPR32UtxOisIqez5wOsxb9UKZOuaTSOPA
CVVAnTNRUuNiFBsZ2H79ts7uPk5UWXjRCN09MVWOgi0gtPSIjmV1FiFcaLj60i/ApHtX0vmNO1hP
pUhPy8qXguOf9W06tt2KG0DFh1ImA5xzc357K78/fP0mu7Mjf1L0lQHCuoaInUd0LbbRXP2Pb0gY
bgc87vULFWc0fAj5trK1s0Cp+SEckotc21uQvytdLyT/zRTTdZXKgummZ6MgS1fIGxZ8QLcIfzkL
vY+VAlz+F2QEsOY9K6TV7sW9JbFM6dJs7pHRPPG86Unil8GvDurMFRZ3ap0mZfWsYLsHJxzsdm/U
ikmdF/Lkb3iE5PEFq1e16dhr2dl55yvRr2yXCNlYLRVc/md9RNLyLFMX3O+UEjEZZGC/ZEzAsw7d
05iCPGUkeMQh0e6qwwsALk2IMu8FGcMIPUH1o09p0fVCUt3lT08cl/5U6yZ2ylPTHZ1/6r/akF7p
mvP/oF87R163TOGwGvoDKJoyg33htDoDZIqTs5vxxkuNsmWSSLO3DO4YnXnfJv3JPclOqTsWyZv3
8c7AD8IHuiU93BBq+7klzs+0K3AuuTVj0YjmGFcj7jlkPp/TzWGDfWfdKsVFPdWf7UjlLfBHJHX9
BJfiPjdk6+ld31qQDQfh6EDtmGS7dwe5JntRzwS+AcQCzuJCfkWm0qYmEevLKgyuF1dAAgY7o4cz
wqoWwmu4ltFSyFF/u1ZnqAWYV7AyxOT8V0kT7NaQ1++AV17SosUUWZNMJl0if2+CRRXkgUcD3wQQ
qxJLkvXtxRZyK6778MgBagowi6Ym8336dXTQrW2go6saT9JwDvfM+iA7xCuG9t4z9aKvkuj1DY7c
lVjw7kbFOKvJa9Ad0cvqu20H7sZDzSxRiUXtABXGpyi7WELlu77mgpYjovkhcEMczQTPjGooi2or
4FQzuX0heYfNVgeBvG+l+3rHncTHMsb/usRgPx2wXmVESG6piM4as0V+AInieP4BnggP1tzRQLfh
bkUaKYmmvl6FSPz9X4hH62pM5Y7EkFaPcw0mV2U5tPtct8jMAH5wQvYes9PSJIyl3aKzpUakv93g
RvkBLQ9Rzy2l0eHSmU53oyKsF+cOIyAyxYiyrFxm0LLkOIaITozq5Wum7IVix4uMZSHyIHDZGO89
irfgrYTauSy1kTntVpKjEGUA7pbYkCl2JVM4tDmHRXheguTlvt0UO1vMS0hy3Jp5tvUIABwUZ+S1
hnO2WCxEw7F9Cb2htCy60MEFc0xvOhyyCKvXrxpLbbqvyS9O4X1p63HEa2Vm8tWT7d2DbOoJYaSS
jm18O/F0UhQ5QiG15+jfswUWiEEgBMBEwcQXshEgeMF5QwYozri88Kq6NGR+fSwwIemkLuY9pfbv
kxCrD49gJqNYPvw/mpsCEgcT36KY/ScDjXCogOnXBkPWt0zYuqxWEXHUSmuE3MgLA49gAprZQjly
RcDu2LrC5aQydRnCPgHnJ9g47XfdSlF6QmIf19cnUYCNrktjshX3YREvmC1nYtutO4miuipN09ol
UvvUgy3txfo7gGNHvNluOcMiLifK7I2c+e7DgmqcA8cz6dK7WMX34YscQ+Tt16c1u7fdcW6rb5/9
nfwoWgeNjzmtWD04ZugTEVSkBA92y4WL9ZIQKGZM9ULPto4Mo/0rKwLvnfA6wcD1gbVBTe7UZgsX
2KrZ+/NceNi/yBzo/kufQZmZM7dIsjAqMmJ8KBUBLgejvu5+8PkvwncidRkuz+MXq/e79QVh57l2
Vde0zkvY11SgCPiZEHKrsGltHEuCvi1ALxfrGdLU6KV/w5ni2c+sqkWGXD2Ur8WJm0kVWkJ7Ukqa
EuagltFvUYFY4mTg0iQENrXZLAkuqX5hmro2YWILr/uJOssE3fH6Ythz8PUUZ1e8IOpajpduo5jf
4Vw5Dxe6Gv6mnDG/q0785+oJri4IEhFFztQPLa+c6bd/KXoxf/AdGH3yX2OHrnbTdpLyMuSNbj1k
ByQnW+DdxRC9MKRna0WywEfe//NaSole4n1aJNDLrYa+Tk+nXKTtsuKDg3zCPDI152InkNxke8JI
bolTdxlANCewIaycyUbzCZ2wW65qi+TFz+c06bvS9ecglRHbdlFTgb/q6JTkiv8om3puUnggihUH
Ihr8BSKx4lUnSvedtRLHhAgfkCt31u1yAwVFbqqsUZguAmSohnYwLIkpJg==
`protect end_protected
