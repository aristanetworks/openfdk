--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
QlXT0e5LDROmR6CeW7FrNntN8tz7cK0QGdcEnplPkVIPQKrudHZp6yDhrhKD+E7POUNndwk+vbxo
OxdIL1PeUlzHeJYmswsS7Pk9x7sf/IeeciM6Ww0RvhoEZivvTVYokRJ2r5EYgHdLaducpA4xDeTb
rda7H4oI1SHlNd3w37IovzN0aUfbim0feW9CLgpaxby40RidOosBEu1zS9rge6ITSKy6iAPYG9i/
DqoUqKWJbDml1eLa++tXn3EbIWKmHzm8kfTGY6th+IC0Xc3ElWhQ3nveWrk86tM5/v/RI0loOj3P
4ebBH1tCMVyDtfSNQoZ0YeXqjXueM8dBYiJZNg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="MBPgZocDS4cv5/haCe1oXCz59OqtRRdB0nUjykGpyko="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
WwP1/GArvvit3PBB1WZiFPf/+3pfVAFXskO6LC50J/o0WVSJca4LH7mH7XaTlf709zJj9ajKzWm6
WPQpliI7i8Lhz1Ojg9N9Tth6StXQ84olhz6n7lfXOJY5PRL7XDMaUacvy+n9Q0dhaWJUchF7Y/P1
4LOy21qmmMa+4hSiKF5WMRDjMFaUlZlhiz3pT5Pp/41xKCVuESXTJsifjcNUUdvUQwP3BCjYB68n
2Lwq5sqVfPSc6RWZTAoNKjSQ3+rBS6Q+CLdpHhY5GMrmxqz+8o5yvZSDv8y/ILKm5G7jAIh4UWh5
7fXNSSsTKcOPYPKWXpXK/yXvD51+CslYLreMLQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="ZaJPbfTu0b78rs38l1DbpOnjnYz6G3yhDTLtf8PdVDo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9440)
`protect data_block
/WWN8+3zwMu9PQHqVuWBhV6jEM8qAPzP4IQAeROKBN8dJXJJK50g5SQ+kI3gF1QD+yR34kY2zjCf
JovVQWnrWklYwBSIAxKvGhisWNnbyhKOS8Gd+4bZsmXIn8laDfXeKcdgVgoi0hurrB9IpdzU5FgF
tcFgZtBiVHr9+Qm5tgGG/EfigLg6wOSPTCTIMRqw+UsgO2MaP+dL/Wm/XYJYYmneXfa7hE/E2TtV
wjsmH58Nwef/unQ1QPwDNZY49tLnmawpt9j4jOB26wpKvfB1oT88f8HcTLycstoViWACoB5dWoIR
GNq4rOFbK0qwEhnbKCmsTdu+SNPDAlH/pavH6/4kgYBhookf0oG9U5IGgLtPVImysgt0nYWAJi1Z
GR4hR2mL85BrPqhfLBtHG9BVyLZO2LeLbGpf2OgDzbCID4pTQdrIp5jAduhSIqROnsJrtfrNNbmI
8ouoyieJGFWAfAPHIGqZpuqOCpY8cuilgHDhBmKEBnfGU7TI44/t9PziDHRCqOSlL8H107YuBkFt
vguxuRG2fNimrxHl9o4eXqzXGNprYMCpV4lmHDKYMbl7ciRj0gISnLRtoPZDBbQSR4yXCK8MCJAy
LiZ0OLfAXykS7q2dzU9c5maoNq8gXrh2F3S+vMdlvowcNtS5AB+kOigwPH9TzqHkyKC5+rWJxKWW
o/hufpCKnMQ9Kv+TtuAZYmz6CVifMMUlPOhTTHQJgQ3g5r6uaIQzuxwsR9kAwPNuxipP8GjbdVRO
8T0ozDS0CDclfvk4pbDiLxwvb0ARUhujytpTreWqtS5bZpUf9GaL+aWgFubsK+ZCqEECabX4FMTd
UgCJWjGji5jXgJwz6DlnwFkjerPI/Qzstyo0SCiZ7whZskpWZA6W6hZX7q3BJ1zfvUkGtrgRt6cM
SZCBogSdbkthvyOdEQYdOsn0qJUnNTlt5UFzsK52QcCwxhCOgrk01rYcLED6JATNP4HrwWb/miMX
J35zMn7xhQUhypqlyrL7rHCAAUC7KhK2JBCYqQ8EfPmA3EDsRnu4cxaXqGQdcsnLNh9+AqRF2ST2
gUoki4nySufx5a8SKsENU/X/Vc4aNu50Sego5LHX+sOgNamyPED9mWN+jNxLrwF6PWwpyo9nLwyN
E4Ljj4UBB9WfgsV8DrcFW0IJOXOi9paItyAXactkQGX5nBo/m/ow9kyPMhgQaOwYk0ITdcdMBxZy
VP+8xF+pFFM6GZDM/COWO/wOYQ1VClFz71oY6ckKRcIaozT5+ltIFH/or8za3gBUiYq1Z9vzeaeX
x/rKS0g0PMFy1bR3TJtpn35DL92tbGAzY25AbYo0eghAmI33MchmReiFMLYH/kPEJ1z10i041+v5
TpjTe/qIdUTgy7MDzQ4ppOC4dx8RAIf05l5aQhid6kyQ3EWCCyAli9A+oD7IkVdVgjjKvdzS1qyB
3Tsrdn3/heNCpphjf1iIWnfzsH3c6GArpM7SjpGpTajje6cYetiKVaBzK+0Btm0ue5VJvb06/8CX
k2ayS7MD2evzqSv1tXTBE3BzTYDY3gY2ShoR/BI2Xxk5fMhat5s4w+IpRExOUUTGKnIBE7yHwiN6
fd9RM+m3UmrBvsTfcO0+oQTKVPl8aebs+hvjEwLRGSJrEuC991FQ3ZG3Ag4O9gp+l6/aCPyBEbGe
qJUY0vCNyXlBLXO80ZtIrhMLS4DyaVztVAzlYAGQ81DnyOhiScZWkR3IpeVWtszEax2kYIlj7cFA
dyzn/YlgrFQRmghIJGZBgbROuoRn3j6Ng+E753m4qRtuq9i1Bl/aA6CbCyxhb47CrSMv6Stl0fdi
qkUfypO6HPVOjTZNpyfC/sPBw039sR0roNFzycq7j35a2UVnxnkyc2p8oxohrwlKGTNNZOT/zArO
RYCqx31mVqx8Ptzamn9fufVF5TOhCDWw/F0dmXILH0kk08X7J2fKmR9QiHET2gBWWdbN5iAEt2NQ
LTDzFB2gJIWkUDDudRAx69dM9CYltW4nSBjmtVIlljaHWfJZr06+amNOLyzbxbmBFCMXnSliKsTD
Yo2mwrIG7Q0MKnqbehV9h7T+Dp+cpqGAjIWzRW0U8wGcnejbvKHNqgju3McrnMNopRz4TgnwQZEG
QPuJbxmOv+Q8tIUoHRyUrlw8t4OhZ6hHBrcekv6rKp8vTJCNpvjNHJkpPCgUU+iZfH1PigYSvP2e
No5qd5BpfqUVupYIK2T2Ie1AdzxBR5KFQ3kauQTuYYYJ8jZtPdEpywFL/8gTNylm27g7AFPhy60+
QwiNv0hiugmFPosNlhB7skYrC7qEe5ZQeGb1RTRiP6XgKRUdpFJ9kZrYtfEaCkKebF/Wa1o3k6LO
pnGJBcdBz5kQmGCacpMhaPkGRAxZq8dcBbT0W65o+Vz1jNA5hBTufhPw2mWbeDjLRUC9lVbUC7h5
mZLYXXDgWdt8NSHz3z48fJk8Sv3ZQDm51Hmom2do9r/HtXQlah0j9ny2wFQSyUWRzCCDX0nE9H6U
ugZTWggMMqaYGaAfF9XE1W0xaCTN8H5gdfiqsMlXcylGZVKI85ETGHXEvvAhfDYrEuput6PNqSuD
Ghl6z0Lld13gHYqJxLOXJEHpimmvQk+vNvzwTDEjws4FhE2Gs5ICZLPIDYMe8Z3BDJJpbKUq7oE5
Sy8pn3sU+uSai7G5dU0CDtKpr1hfydSRccNIBRyHzgcMEEcZjsoTtmUF+JdzMNPVAsWeKJnWQ0g5
pDVTN3A9bIHO2TTxnQ2PC/xFHxthq0MMGTP2PmHORhv0J/9wBrIbGWtKvkRGsS+vCNbpwaRQo9FO
8KjbULIM1/rDtJMLmIxPk1fxgXjyyc9UgChTP0u1McZ6LANA7RCnvXJB9AQUi+N7D8HQ9sDvVNV4
7+4ss3PkJJtAok0H+o2DcaKeQSKQi9RzZR1Wl1a6MJrXkzpujC198lyljAfJKm40to+cslImLdCk
F0QCyc0wZJvLQDJIy6zqaRBqR5xNO5SWt/YpIvCDnMNECP3TaGbjlJsU/uE0O7l0ADXcB0eLNDfZ
fmSgcP1MCv1Gv2tWCNEFGw+Krz4+HGzjLMQKnhOc855zHuEqzMOsXhGfzcEgN1DoxDgQiaWOeyB9
6+Ub3eqgNvOsV9nYD6wlBk8AR/BA9QOWnktHs2qHbz6/9aYGYihSkoDFyltpcIkeb1uFF9bsfp4f
aptw4qsn/AYe4KrL0iRoEqAwM/K1OowlCxixoTt7FtGMefdWUUgV+BSdhs5ls4st5w+X1ozedfbA
PQf3/AUpoyCTFxfwl4HuwAp8W75Gbpfgc80zhFyGhLY7TJPtis7wE4zzDcgFzYWQAUI1h6t3dWjm
AirUhSpMvxigwDH/y9qctS21Ma4sOJKvvDv4+kz4aNANZOrJu/Aavk8+oSYaGstI3gIPAQDAKrKZ
2LxRoBWxIT0jFX+5aaTSaPi6tkzA8zcae99dKh1fmvnbDgQk0Xqf7/4zJuE52oVNuLGewRf2+0uy
dSg4Cnn3Da0KHdqYHr278vJ5M8HU+FuKt3caDvdEJnp1GUEqV0semMhwoEMttB7TyUVoD7cIkFt6
bijokP7U8YQnb+GIBFakHTYWWU1VE+Rla/K1m0vUR8u73RMX/+QmZdgH9s7zUIkI/sdLjmEoAf+J
I4lm1o3ivijtJvjByuUfAVO8UszkXZN/zX1gZ5XGsCziGb/V5DiJoSuSeSDzMkZkSbE+KdQvRuzY
zqiDRI8rwwlCzlnekGkk3YqKPaoMKxqKD35L8jd/JsHyibn40eaegEUzjViAaCZxk8LqMbnwhipY
iDC9VRBGYDMuQzusavJCKZTsD33G/ZGQlWedFjvyFq6lm/vLEdoVRzX2JfZc3qheZQ3eR6w6Ovhp
XxuXYGFXwK7l2+ldXbrBaYewEi9ujYvMvpqHkG5V7M+GcUK4kOaWH8pUpTcRaU7GE+x5Iqu8Vpg+
mMk7kpD8h81lWtJQULK9a2rftLoJ0j8MxTFW4IUROu9pCH6xZOPjiB05rTgAyb8Gp4CSvkWFQYHq
gIUuhRDQ6HEcjlJhonD1I9XpBz2B9KFlm4C0cxwk73ecbzMOFvgIdkTP2EBeLpsZzCIRd75xLM5M
5dW0dvoX6gvoZy4xRPk/fwznmwjxxwzM31LQqen2b02jYUi2/VRzlDF3Nenss0VBL6Kkj6rYfojd
w2jmNZ3PY4E612aWAsW3WUJDeNICNVeyDWcLwx8wqtz3UyxYtVJyxcYImvVUtwlMjr2G+9k3m+Ee
+RslEQ9WrBLAq14LppJF6i9OEyM5rd5FB3sW3PiwABzvrhoT+bXL3KIw5YaWZ1KhnpKrlVhioMEv
WoZNwBma+yQFA9HSERsWtQNbs+Dos4ENz7To3bQaK7CxaBmufVACWCEGRaVPykV7GaWqzwbam1nu
+Ykbe6NPmoPOWOubmNyuRm/mDlDkfUPNgF7HMQNocq/t6gYlGWuJ2x7OslK8tqlOKRmkaawjub5D
h4NlFUcJS2LD+Tr6SFd0GrxQLFstHSBLGyjGDZyfKzcqql3NGHaGSHnnptBtlD/qXb+TEpmtz4Im
bmyUj8e2wpb9Y/4myXdakCMJkP5PRqmkquMG2H/bRFLQMKzYrpAlgg59sCYW8AkWH6P0XTT56oqc
CTJIkGtxhqaiwiExqRaPpkmdMTcC7n8psrlyy+DsuedLMcFkBBmp6jJ0TU1/3mfLb9RZhElKmp2E
8ASq9n0oVvu4c67T5hthGUHspzx62/QU6qJZNt1df810fxx0cFqJd7fiwytAJovDXZEQb4sEkagH
a8pKDejAzPEB91wHOU0cN4qRvH7J2pd/PbHnqYrMxRhuLN/7mE7zyPk10q84kYym2plpVlfuWnhD
3LUbJHkoo0NOEWvtdlsFpB9n4JaaDxN+vANnpPUSIXWtlfTZKSWJyD6cUT5wECMLTA+4l7nUlciV
aAIdie9xjYbxIhf0EoS0NMt0u6bCltgR6wgobyFAN7Rj8fDdakABVxwhIZp5L5XAR5/uoFu4mTBq
v8bVePllXs3yf48RCnhhyJswdt5MCc4fHKBHgptLkR2nl3U37F8+mfzCK4WTgdQxZks6Y4FNIRVj
x7qHqQwjV9dD4IoFFeCeCIs9oECF3L0x6uneQdGK1ol9CN9SrBQQ/ODVk1B3O5Wgs7CnmkPGnf0b
IixyI4y7jvAWSm4OqwDSXsZdArht2ZzlUCEdI16Dts5RndRy0BnoRongBidoY1MrsBMyJlc6cmgG
xCbP35J2TqMG/rd/05PnHi9wWzKd0RuuyanBg+AHR9tTPgjDD2/fWHfBPCJJcT05jkYzTmShLic6
lpT6qAJfYK0jZ7qoMa0XzwFSCipeJBQjOX3royIs2MnY0H0Mzw2ktbrILklF02D4alnXmblY/c8P
kiOwitNZFbBuoSBvHNov4wSsmrzmLJaC6gXVAA2pLyE6kGjVMlwG0S0Ymi3FfDyv9SnHJfAl7r8Z
AsOrvksBYW3ahVXxF1FrqTx5AQUfljxvIRmXA/OMKv19YrlmYgjVtYpoec67q/brtVRBIzCUUKBt
OeaSYgnuZIJLiP7fuluOjOHvoKFR9oyIyFXxVIR/FIqcN807UTGe1vpGfM27pt0UX1Sb9lh5eQso
k8d0Cj+ylqBe0PK5QkmDiIT2Vyj9hjLcRdPxaBG+mD0YVjJ3p/s6Y1eWDLa3U+2eAQ8ZglRvS8P0
L/RACzXkRD9PP4pXsqS9MDWZNuaKXMbi8Zexeu50dNsoIIXkv/utggodFhGn0qj0mntCrvqT2gpk
lPVc93xywo7EqVS6Xf0/vUTyPp2ENgu3XQhdoZB5imBo1fSRFOFFVYzJHp7isB93cNujRDezhewr
MPhHbda3UWj64JTy+Wp/Sm6cJ7D2fXCEoV05McZEnwyeaAM9q/XWlSQ+boFadLTgewYZjZ1n+jxk
9xkAmn9Pz/YLuskeoboa3V/fGTH5edWsmIYLsyP2jkxMWaTAckv2yGGD9C5MKTSnV1j7rCZT2zVS
p5ShfgtCscPUdP/UJl0IeR9JqqETJ2HrN9Rjtpvm4XrGK1nOBQ997X43rfCb+BTytYN146GjBjUV
lCk204yAqaYaYbYi4Jx3gN9zzjBAp2sYEDfMaGUX2hb19CsFW1spp3g95IGiBX17ct3qeCkCkbhi
5dcbI1x0u817wRoTXN+RO6nYxch1VzeoR1hKSNWSSCW9HY2pQyArrQ9iuD7ZPcZHrxsXwysDx3ef
orCeYp/3lwWs5hs2xU6XE3BvZLppEMlUz+uiZ4VoquMM8wIvSK9SIwMwAugp9+Hax7/1mc8XSoh4
rRwi7o9rt3QrSdU3hnuXHO1SoB41DkfdAyajYmQWJnp9IWrMCBrazX/b6gTr8Cv1wT6DoSxtCU/0
tP1KIhZTmw6nV2zaTiu394ffiZgfYtQWd4J2T2HIbjBtQLtnwsQmNF8BI9jGL6VF5s4M1EGnial4
vBtKjX83AyhV8sy6FYIAjSdPiL8qgNOPPTl8CQn6eILIJ98RyKoqURJbi1EVeGTWP3ee9kuOfyT6
KJLWrKGRujeg+H8wA7PU/k6BxopMluf6Qp+Lx32OZrOq8zR5lUYiuyebKEtPcMjK6Rk0S3YILI4s
01MdJhRrXlgw/3cRyWxJ/mya+Dz/cIlqpK4NioSlc2fthQ7x9SWTBluhymi/VBeKOiENCPjD9gio
RL2DG2VsKbqAdeAm1L2dC8AlTj3xb6vmd/rrEFCMIg/14vP+4s83F43gNK76+KsQP5Cz5RFH2zOz
zEVUtQUeTnUtTQ4ZXwC8mK1eEZFwE9TlGQ+pBFt4b7G+yo6gWOd4whzCE8IX43InsYvtAYFrIS8k
uileyWssm4OVzkdxCnPU09qCjDdZW4q7GbvQLXpDC1Msdm0ADCBDpL+KwpGeA/ViccyyWMFJb3gR
oKavfbPGxWsW8gHdqHhcATLP2eFGhS61+GfdgjKFw6NfyiFw57Ga0bKIAucrgcbPEHXurHlT6xHs
lSstrbAiQwhR/grzMEotgHODLHls+ixBoHO1P9GARn4iRlxEc0u22gcpMdxjc7Xr7H4DqCcuPviV
dFRVVS5VM5j+010nJwiFd0ciMBqM84deD9SfdtLqRXBGVyQmcJOdj+KfExWxExANjbhuNwtunFA2
s7zRQc3ThRBcOA1fmGSnLoMaLtQGL/3UbC92RcHnkDUqwU6xey8tPcr72y5ls3gWDDAsdVKx8Hz6
5lp7UBwzMHjE6dVVr6abLnrhOBEoLWdM6EbkdfD9J53DJHq6I9OYsFj2Y9dhWZ6D74aIzUayUWHg
It6GZwU/67rqe37n5i0tx+xTQc+4UKPKbdEgK4NfCN7iWLWP9AU7PObQahBRLWjb1gOHyICDa2Y4
Qn4IM6o+w0XmYIUo5g3LkWc7zjAjPssalVodfOfZB0BDl9WY4ER0FqOZ3mmgMPvCDWRGfLPGpWi/
aIdiQGmz7cdxjD+1rR9gQkkW3UMtQeZ8nf1yShfouaKHWbiqwzqns/7SRrM6q4fbXhX0/N2siwRv
leIzozvSKjGqkGJF6z9T7U/riTwKl/iucrAKHb+P6QCbr9BB+vX/g0OViOTCmSJWrMdWPO6LCxWa
9pBTR9Hl8Jv/QJJqofGmmup756DPD5oj0WuQXy3qCpy6sHhKLB5mK09WupGXT/nKj7MPqTTVc88k
Vq2/J7uU5glAgWhpMYtGBAaLdmZMIPjCaILjpXXo2VEM/Q710SFJWJpoB6IbR2+0+7qFwE3pkYq0
fG+qzRd7hv/OAk6089A3hwN2ZVuQWbmtX7UuzERDWZfbQRWVsX3N80Oy+DeBxduGT1L6He7d6954
t/9MplH5X5c7XyDObA444+6mXAhlbcneSRVYwknx2mCwR7sjuOXKvzvMN0O478uOQU0qWZL9zcwR
UyROhyyEFi6SckEzPXXALNEYAcb8jOZhQ6bGDh1TA6T36/lJTqmi8H24kXvGjtQeWD0rMKHaXp9c
OdTnVMWBNwY6o0gponK6EN0rd50xzaNhzrwepcLTblQijCIl1W7dus/xlTIeCN+RtYePqcUKwlKx
oeGX5m9SszvVcTfDIwNGMH+KaxUD7T34G2rzcZi1yxjT06fRfw4G8laZqWPqFwL3l2iLEdTWtnM0
dzdqKbo9aZOEzNpykw/BtU1o0wM1QelbAJHe2fMyYB3xOQGf/PT88T0IHnZGsKSCDcIcc0sU9b3T
XoeVriQTDp2cbqzS+B2DH3UGw0OOHl0OshlNlg/d48quUtGG7+rEs17KX9Qt/onkgI+/KupYwnzt
JL73lgtWcUyBUzd4QRkFEtSr7NKhv/RWVgNK8b4p5r+5D3SN20r3N/ptDaC2ivMVJ4nijbPwuGsW
lcpLpzaE0npgJzFhVVBh/UK2k/GqEaX02INKd/g77ts3IKQsKo5WMH/XUat/8/IxR4f7l27jTxoS
SZYWhLkYIdR3anduJt3laivWNAmlf4XDTA+/RuoDRBIDkN2/7B/wD++1Zn5NBJDVKYVs6Wu0kksH
mNq+BA6G6wA+0KtHOwBifsCxVXgS4sD/dPuPIJTeaNbATVbAra4Efv8Gk+UEGz6y8KaN9IMjoBR+
gaqSLO8P25saBghhXrB6/v/0gXypwOyp3NA25w1iDGp1jBaPzaDtMjUDmkgPRvKZGp9BEmcd78oG
r7whR+uTT/l12anTnfXk/iU1UqwhZgX60EyydV39yHf8FPoZwVKnoc6lA+2Bgzi0enH5S7qGq7Vq
6SbJPE1nDzVuKBUPCx0leaD2ZxhD6arTO6xOAZ/WsFAjRRuq99/hEKlUyepHLU12/5JmqmsnYkSq
sd4qW1RxyVOGaJzlj6StfcL1F4cQAWSiUeqS/WXkijd+B0nL+7aPisexuNauZezG1c6SRvaxQ2Od
nc0pEmscxLeKpXN/KKatWwkvjLOzHA6/s4Cj7lhHkL9LCYWuFOICyJl5mrGNvOs8ZrlmJjRzFhV2
5IH2/YI8V00ufwjxnW8D8IRt8HEU68xvswcI6df9snZBwG4qho4VumBRgTjZ/Egr8O6NXK2UJDpt
GSRH4Nx0OMiPTadtJmVYshJ3pp03Nsndj2wRgEJg+i8afw42kJRTDKEwS05RqCYA2f2OCenqsrR6
HvF9MzqhW3VnjPCkBv8ezWwJutZ6VO8XOks16psus7f3mgy8tMtnyjijff9zwngICeggLcaIgSFo
4w5/s2XufFGpCiBWgUdNaBcukxgsVP73bqerlurOWDcwD1cdvN6vIXr2esMC3OfmUrQ3X0rRzwAK
0N3LXU4+CB9U3dAjRJjq5AcpJEZAl8dl6hKTKJuI9zWjf3ODBDqM2RPf6Kfvetf/v6BWVYgCwftL
dxX7SmMRKPI3vHqXWASXQMr9XDeLM2ylSoLZR/DK+dH8a/New8/R+tphDwJgT+MyZeP/oaeYi5IK
USNZDYMKC7aEjz1YQMNRg4wkYXnE8BjU7gepZ0cT/Y5LGbfC9KlvL9loFtmPJx3oMV6JBNeND08o
OEdtaqaYkuFOkFyB8P8Pbo9h3U4uXabButhBnvzaH6MO/vNrhOzfYvxsbmGw9wFN1KtzlMRg9VAN
fn+Eo/GZgOS6DE55+Mow5YXiJt/MkKHDTGScrm4HHk/fs7oiuEOKKPF5p8W8DL9AosfC6vs2y6BT
ud0RWYeVP9Xzfz+JbjIJeDZ/UCrl6HPCElKW2bPBPnY70qN43K/p8t+5GI05oIgp8/y3MKd87z/j
5Yr6tZJCeIvshPTduCMK4bfJoW0wNuYHDOEnylRw3saKEq77BVeA4RRb5bBd1FFmeNck9kFpdsOC
Z8q2mdZkOKz/vWND/Ek/C5CBa12Z3jnUP67s6hXb/Bs1ZnBfAecmf+w05bupW9Otx4rS+FheAt9l
JQVNURblJPnz6NPLuC1DlUj2z5DNIXe4bzNaFB1C7J1RSbQbRBXQvbi/Nilu9intmtNctmGWjgyn
C3aHJepAylD20kQjH8pz2tBctn5Z9CI8iFpYnwUvpquzQYhNkp0pBtFbdUG9VDarpTnk4u8mmhFp
OweK0orcKzq/wpBlhQLH48kPZ6iPu82eBS/HVFE28FfOkG4v4dNAGpb06RCuZKi8qEmK7/JfLDYm
k7z7DkI4olrsRDuLtw7Dm5/zc10r27f4nnk5JdClJi3dpHJbWStfdjbGOWO6+oMAv0X4gk2Xl2Bf
SIZLdLNzG4kJwRKulJc34ZtsMrnGhGAiV/7SnFQ0XyFpGVBnaQZhXhP6sk81Zvt4fAxxgeuK2nY4
8FerFZm06sPJBcdfbZxnKObZIVqUbqD3TqrShvnD8ewUDe8ZIJC2Bjvi4rEZPSrXd0+97Vq0mejW
HEXxYhATfSJMwxloluYzFGGTm4poD/Ydlevy/I+iukbDiinbIITgwM+xSegSNXLSwCMVa644+i2T
H5bLUtWkKoM2lAE6KsR//mpoVsLs9n88VKPa8Z3r15YltQfK5s/tHW7ujqXrnVhHqc9suaYNuhLG
xTYin9dn3gKjrEecQTejuc5EJeTur4rF/un5ca8L6hAeWkGZoxoXTULHM1ytin+YERI+aGyGXNsr
oxBhjZster2we7XqEZVY2Sxz7rMHCRjBufFtwZbL8VHGdLNAEBT373Pr+e5o3cnA/beQpeNa/9uj
fzqdGoQblkXOEz80rZFMoe8+b+DAzvHH7RjV+ieGmM4EiymuKfKzAL8fzlJfZx4fYV4mdMhtXvzT
pcNrJ3IFG+mHI9Kvc6aGgw3u8cbJwMwOks4mH0Dulaa6dILubKizDsVzD/Px/C4U2eaxIpLgZp1x
qydPupFdDuoADXcBzRigEHobD9ps2WiwKfUgYN/uES2t5pxqHsTwphESKNHgYZQIrCoZW5bVhJDR
fRzsVd9KgzetYubZ8cCH2Tzs2OYaGa302Yf4w7zgXb8tuFcOTvP4iCDOxuUngWXFbecJwm7A6Tnf
fED3QlBhq4F66Xlgu7yCpAKd2pXhxyvWqDbhv/dmn7lnqCHPTA0GpFZ1TNYcteC91Dq+O5vFO5FJ
bobYLYG41zJRWIoahsSigP9GQYQR4yWuGjsu3dFsFt2/RTg6ddsBSwNb0ZMA8q+1LJsuXlQhJM3q
o/I8mnkUnAd+6Bg6/btVtcPxdcnCa5KdYGUd4jJ0/BlJ3lJajFYQePDUOKJBE5zEq53uC4rBKGDB
4V7Iv+LAsCArSDRmfCaz0huOdppie21npNRqO6IaAPEURzSpD5ZpgY0ZRFHMrGXuvpd/czOCpEoI
+Mwzr41+Clkf+b3RTJXfPPTZosgCwo36ijUT3wP9Qs7CZOCW7EW8/kCR92m3GgY4z3bC4Y9tAspi
RCPWexZqJokIl6DqLXeLov8JoIvakUXUqAcVMY5ohSlvgQJel0Qg98yCsyb2y93uv7v3c5pRYZo6
segcQgsEWasXoK4H3IhisQRwH2SVfEyR437xxyEd7RfU8MWeYAhETsQ3PWCvJRilR6goaCHIB5Kf
VNZKF92UMWx6HZ7xggQ4jdJSQIcVBsbWpA31ZFMoXbYJ4B81hVIHZxJtgp3Cb73AkdrsQaGFIF7m
bo1wk1n6O1u38ixT+KN9O4jlrvufdIpHAd2P6mmYenzHd819zSpXhjDrfr84qw8iNrrxwQ/uGKWv
ErKtHCwmaU1rECh/oh3qiWfnQCGxQ03s99LY0i1pJvkAzbnHCPNjIXBwNCzPDW5OyspFWs9+BCPg
B2odN6iOiJNOGjbq0sW65jNbk8L/DZnWVqqaFX3nEDk7mapxjH6q4sSHoxFaofke9nol1kJWJ/er
95a5ssPqzlvqBEHZUXMF9ORNFWv4vIQaBvHjolMjTYX6d7Ssd36FBu+YDtaFajuHJhQtzsVVlOxq
HUjZcbAwKhI378zy/HoM4s7Cu2Rh8uZEo/3PYpHLwAYU7tF/ICbJLBF+f7JFKnl1TtpaJhm9OOSG
joaKHIfgxDWsfN5NdrytEIyQjCIJs/fKbCeZ4qeW5V9zR02GgSwEQF1HCB03CBYO+XjXxHYVA8ZW
yitG3mJ6iChsukOY0abdm4n/jddsBpd9AwTzrVBdmw11UmAX1LukJcGiyIpG9/iD3OxRla7C8V/9
iK0zLU3NPqi8lUpNE3WzOlXnDOCQI7z1CxwQ/A84g48EHze+uHJiMDmm2HOgQq1WoszNxwPNBM8O
4v3NHjyCPl7Wld4EhmvfE41zhyyBvvxo5M0mgwyRX6iPYjkJpHdlGFghUE0cHoMBQs/XQJKPusVO
qNege4RUOo494yJTsoVGIf411t13iqR08JqpqSKAe721VCNSmjnhoAETDcnJB3bFCVYV6tt724qI
nQsn9Lg1iOdobqn8TlFYkGsOx6UGQemUr4Kc6oGC9/TKTZmychd3CMPKoWi3yReVGA9pagQiodmq
NLk2W1LFXEpHW6in9UBBYX6bvduizQFrOc+/HGX8mxzwrjhFbQo/p3cjuXmZfyEnLozFgGGPEVcb
lNvxyuIjlPHrs7SGc6hByxMdkWttyFZMda3WjHuOl5/xxnW0B1gG3HbCD+++1yEykXGtOBRjRtMN
8qgVNMwhgWvHkflYzNMyUK1NkZqkn4bUDnKo6KpaK0ejjHA=
`protect end_protected
