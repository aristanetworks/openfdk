--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
HxvM5ewG8lSRV1/zF9hHi4ZGU3Me+JZJjQ53JtgPrIooMDa0ByDbv8eGeJAPybrzCBbFdxtP0pCg
edZRWYjnncFa15H3AbILiwgY1z2XhBTWm4qWHnpLnE4QMeL7jc38yM9UBLUEDB38Ym5TxHyjNH+1
qL1S5JPr9mCU4ZMrC4H5VcQWcJ5k71qwcysHoePon/33vdhwyHN9j9IxGi6V91svbQ8vHCWanK9c
LCHVeLhtkUkh6c+Q34GhBsRLQLdfPyjsrtZCe/7qaBGusyihr3AJmUfGB7/g37W101ZKIb+Bwj8H
tWV9Uymg1GWO4rjhyB3QY7bpiqmPYiO3ILCQ0Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="fJAnh3JSijoEdYp3lXlF+BJqrAcP15G0Cw4HVM49GLA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
GDvYwr3fOKIUbdPTbfQ1avOdEVON9xhO2aIpXLZg9VVBjx7Q7YWpaXWOSJ+T4piDDftHOUjJFsDj
XP+zlV1uuPod6oLQSpI0a0+n6N3cCVNUrAjGeeQ21R8m9g0evoqW5Sd6U4I2fUz2K3j09j3Hj8Sk
SugmT/CB8RrguwG37qHdNp4grMYakpJbbCDk+WK+nNqWBHl96QzYf5hzBUc3kepMwU7tkDV8zWuV
Y9KNDx4NgsiwkuITzqk6U9DX96AN8MFnayOZzA5f8uW2azjxKTlO1y8EvaM8HbdGjWJ51tyf2osu
ee6o4L0s+tfrFpWOC8a8vjDF8qSMVh7ZrVcGSg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="PT8kIYhKZ0N7uO/oS4SUVJMoE7kcPIE84ZWMc42oQlk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2912)
`protect data_block
MMg5uhbp9sx8UplhAMjsz/b/ivaQsT8A3tMaIINbwV1H+Pt73+bUqx7U4vggUGnYJiSMb+h/BM+b
Bp9CxEktBqFYGm6+CZpIHqvi6KZGDOlXR7cAfueqBonoqs6oKbR9tt6PzqHb4OgPe72Z84kI+DnR
dE71dAkI14zVN4vOjZxJqY9NKA1damrufhm+GuN4bxstBbPzrZBmfdO/WuUFLnGi5PuDxmNmKYyd
oUyti4NFmMajqasX8l7g+0K2VbNZgtuwo5BkSpEcnxTogSsk6TwAXFE1tcw8yeym6HONwuF0Ftv7
zUYZ2vK+xDWomHk977mbEYQgOVUoR8qB6TgHHPveQT/VjrNYi+46gFS7gxc8dlgotvodnm46P5q4
OFOvfLPmSem7KkUIKxnH4FIxGgChDfmuN+iSipUboNRP3+1W3dFbYDTHlnDHPSpm/KZ6sJQGxP+1
cttXTp9T66xIsWGnmQlMrd7N9hAJj74VxrcQVsb2x/quZRuz5CsbNWYe5dF+M0AvJMC7mMChid0g
+9sCj9UIcLbc7qqReo88+PTWfYM5limW/r/RGmB+xluafKKWkMIBXsIQj58toGklSy+6Ol+GGBPE
RGu/8G4u+9QsVp4GVWjoekOxMSuyoIZggUb7XaNk4KhqhEzoJSIIFev5NViFA0S8z5Nq0itk1cFC
iKZ5Vv6PT3tkACK7OpvJiY0LExfaNQTYxI1A96TSKuMGZ/8X/DKpWOb5V1dwIFYuUfC9ImnxU29P
1yRA9cJQ1YALHD1G6OiqZBTaX3e7ZdwCrUH/FCZQ6aV5wQ5eDmNpMFgk3ZtIMbDz49hwTkXXiN2w
5CRmjDxtYwP+54v59jl83tVhFM6T2npV61unN6R8mHG6zF4nXWU9gZVgSPcMBPx7/FiYZoE7GE8C
bS85esAAG7PFTGrN+jhIWRbbKdYjbeRvzDmGF34276zCpXMEzsw0zM8hAqB1Xze4tF3gJ2g6kTtT
Ogcc7KxyW12H6FWFQJDwNHQL6RZ6vxefdkiPWvZ4wtrNsI3Y52A686muCRYGfnBaVWKw2/rhiQqa
8s63Zl8IjmEssHZeRYHxzuL2a3F0Tq5DMwMtwbPrOMzzc/jZRkBBDMGtP/GBNLaUaWmwt3DI2D26
+p6R0mEuTaFMOIGCkW05Xq2SOr3SwrGAaWAIzlD3rsRr9wgjp6O2s9pUbN3xTV3DAGeCf6UfKs97
L8xleDmufTuEtN6ous6i0L7A4PeT3Q13aAaUTmEQctNmF9D/DR50+LrRIKtYUepAZApLeNwc3P0j
bOzAt6to2mfoZ/CzVd92sf0W0Zx1PeZQRfgcDwybu7hgOXk9+d7wACzeF3zoaklb9ghmKizeUgo7
6yTEU9nLFT65ZZD31dGXTDI1HnUT5nXCYosPIKRdp3BLR+CK6gc2lqo1gac3MHuI/FpnnVkKs8iH
sBCtU9w9pCxbSxmjjLTXsQ8uLhveO/YrTPvGyvgxLo4IBzC1vbded3ZDmkkWLI+hYudbHJzSy4V8
+Q+JRukfiXetn3qxKtK2JWr5tlQAkZSeNlQM6jTXZ35GpAW2nXW04XgQ6A4u/cah2/KFp3Oy6dgP
MsjklCh9FLq9U9wD3ps/AOAM3cuFFQixfcue1uC7UljS+8u2htScGy+X62XGeDTDm7Y+NVjAAgFo
W+VHYkHmLtNffiqAgA1ygscg8Cl2IxFxk99mCvX+mBzD8WdKbxFwxhlOfyvQUlTMtqrybgOEqNmo
jvyG1oiD5WGfIIG5ibR+cBluaXeMUFCzxmMYR10OiPgx724aNvsPXd7WQY+xLQQOW8qExiaNcuCr
dWbNzU02dql3pB2gSEIJ8kfY4eLHyi3KYbkhmpK60a8+8foO8IYQo8apqafb15vQR2M9fIFD1cuD
LoZdChF5mBb6jWG7hsgUtiE+7YZRdkp3NyCc5i2pbI2XBg6a0uLeyK9i7V9bEkaSSXKyqXj3lC9u
d5b64536Ov7vdiNmQhFqbMPHH+eyiLpQeO2Ov6Rm7lgKWXfJdJ1NIAuzbaTRunKJqtW0AR2yz2Pp
BdJV4N5dIacK8ss4ZCWsUPnNL3e/JcWvX/MoCrk2mZ2mEcnMRphEyIRTveQOBi/ADPbjQISL+ryh
JXhM1z+L4JSlyGRFMNwHqIkuUPVM47ljAUSfy5hjvjQ1trhsgV0RvnuGN5YSJjIhMWTVoKmtWsPu
DXtT0vqkp3KcMQkVfNrPhs5ewFu5NqNw1hGiEFJqf0qt3BfsP5a52mfzaGI8ee8OWfBfIPbBfbMI
uod4yaOootp+Arx0RdAZZfsEiIsEYRhPhX56KAvG0T3G751GJbk/O+WzOFZ8OCG/oMK1WBdRP2uh
T4FpE7/3r+Bg3AEroQdT0U/i4uaZo4/CuDUiozurPPeJysXUU531LVUmvt+GIONRNfcMLLWad1zq
gh7+0PQNO+po8Y1TsgoXqDqfPVkR8TcB5XNuFf6P6bTfvf2C4mjuCflr9fySG10lmPpPeAoGfega
9EZi3ea4nPlcQUiWI/zkTg/Rgt16P90N+7ZRsQldHQMArqZUuW6OsXC5io87/On9LPBaB5kuDXaj
emNiFKnc8L+CBjb+fOO/6Qo5r2mbTdWEYCN9OdOWU9tVGWKnc1lHov768fhKZ0DJ4Aga3v3O8aCB
9WLAStEpaQreClX+AQzHs5JudGPZVE6rq2gvKaN0kPo6bPiqb9hnWAPbkoejOlHJcnOGQPDStB3m
FOHXZWSy94AGpZueqeUE24Ei9AiBJdahoR+cCd0iNej6MhK1vCFoNVX9sPPtu51Y92fSO/8pDlEj
wKlKr2d1JAWwYAjGEVUDNj2v3LB7lxjzf2Nb/VmW8XJm+EzUWyDzVtrOPzHcVCweCQmkTctCgo2V
r4etLeuoIWX7LXp8+0kKrbaLBl1bzFysOk72rHPb48YYfciWKYY1+JdILLV7tatWetaE8ktUSxUj
1EHilSOuFEEGUUVyMDEM9CpmHQwKB/o/CYklo7CelOJf3k3fKBwQWbFrFDyvdynkiFAP2TEH7oKK
wni7ID4b/B+cBatA9B24kA5CrULkD1+f3XCvdQmjAamdd8k226eT2AZchZokXLKhsU+Fo5jvSd1S
NlAiCFvKXhjZTWOLeqYlXUwyJ0bcLk5K67Y2Me+aABKkCbNqQK9hrGBC9GguFzZSb7/KKoOgOlWO
3hbVthi8bFZH+/XuV1/VrE9R5d+GRxOEXc8H5q9rdooWK/fA8LJl2+3tDfzEubLXLk3uRlebCOC8
XToUri8w5SqbR2R4Re6K6dbLUAQy0k+5W9JBlOjFYpBbXrDHtHSfCJhcZueOCgSVPOb0hEBiWtDN
hCG5IVzbFhDidAqnfcmsy+wqU0886SgrqLzm538QXogJQLfUoF524qUEX0+GWVDeI2lPonxMoJT3
yyXeJ8qjjRB3BP5COw0FtC2ECHhg0YOh2ioTuRqy+D9/i0fldlbzOFZ6rHKiSyq9LatxNxhSEZNo
qwcdV9cKpQx0DKHc60HRtooHR9p5F36y8DfoTMEviQ97Pilb1S5laL9cyLQdxCJ47UGj362BTpIs
RqUCh0+69zmkkbBRed0huddGIOTKXiD6YNU/HSdYtuDW2b0g9pPRpcPEqkzcEQFC4tcv5Xpam/k2
I+jsCWXyi9E+7jyFSPmAItdtdC1cGK5FG9aIemutRxYY+U9RzsbX71jBzAjpexP4WBXJExJKGY5i
UEF+Ux/q8tZnhMgOGe7J0Od/C9rL/V3qaZQeDF5lFeORJignAbJpoVJXnuOL23jFoZSmqPdcq9Rv
9sWocbt5kCKYyVvZNTIHRzov/xqtFbxPbCxa6WgFFOWmUlRK22p5OYAh2fjxq39qRTPk7U/oXuQS
NDUVjOU=
`protect end_protected
