--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
RouO0yFSwz61TKFYxoc+wR4TRYbhuZwLlldJskrvj2g5y9YJhPOCS6aO4hHwbN3WJS8BPmMCc5h2
bs1wBKkUeEUjF3FshneVwcNCwlT/nRqPkBTngmgQLaazwKJTTHesIJ4+cBw5HV36SI94Cbj5wi3o
PzlR9DNwzKKhAOIS37tEnNPY4RrYwtToM7RGhjZZK2ZWTIXh1IdpULcq2dKXoJuwlffJ25jpVvTS
A8ptnrw1P/9+iT847Z21Svfb6DjFCZLi/FWCYq59vUGqNGjBExuRkubMo1Oqp2c5IB5Q2TTLlO+V
hdZdWHqA5NR2S56GNArDxn4o+jo86HHP8fYATA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="6iRlQ9RFB1AGp06f7uB0e+in7SREPL5PvealbCyv7Wo="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
GULwOo3avCjdXa8cywnj/K7TfxUHnt63PJke+wMPJ+nqWb5out7Udz2L08b7mWyL7cWVPKL3P0DS
juiCAXSLjPtBOgr9/w7k4u0LVsIG+AbIxhFruEDGegfU5ldmpEmneojWgA7EXOO/OkF/elxZaI3a
7Nl3SbEv0PcYvaGUMIfl36+yv6pW9BznyuGVDUOwEbZpCr3fJucPiKho7/r3IJMYL2T4Je8BxF8z
C/7nHrBni/cIYH0BHSBmX1yfeAfyjm9e+JNKL2bzOjjz8bQr0oNeV6pRp/yNbkms9H8B/es2CwMI
i9G0j4V0wG79/rWQi55RSKGkC5/tOLwGyM1JaQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="lUEkW/5+6KfXsaQAUEJvAANfoYreaeK5P1u4F8ZQmZ4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4480)
`protect data_block
MXXpWygjbyqVQ8HqGMhjB8cK3ThKm/wq+7Rjx0Iq4Y6bc70n2CB9pbKnsONT6kXvOWXopUzsnN5/
fnWfm02GVXUtTiDMuUSxe0MpQjdoJIhKlwPDmAr4fQKMqGtZjGFxjE82ttrv5jDrj/skeRVoMCXb
dcfVeP5C1AlPQNPrYbJNaicDHqxl60HM/rctfg5y2vmixXH6hfAUMQ6bx1hLhjZvsGf7YoalR5Oj
ALqSKzdxxlC5ZOpfLSlI1eA2uhC4AZvjGAtlc/b/HKKyMUsy2N8kTaaW3set88lOsylCqlHx3nnG
GzLqg8o4T5ndTWnn3qv0zrTQUgCZxH7v2ypg4xxFYCvBnTAOBPX6NuQBrHeuVSbXk3F/Tqr9fSPf
qBKvgGpNeBW0KfgWNfzMbpMy2XlAowuS3YO6rn7KN9/IhLtzuo6h1XMntz4ncScrHBSeruURtpvT
nyY1eiR40dFS9RGwJBQ0ZMpPhoWtSVJaoi/FU5jNC5gquDQvkSDbuu8j01W+s7Rlk7BAPYihQnh6
QQbUtVMp6qtsLH/xfniGQzxbgdEDwtV+oJfNPIg/AJiv0hdcMrzc1H00VHXLiSOXrATOzsczidoo
aezFTA0Hrh5yJS+HV34nkPOSUszJrWG+VN5Y5vbC5yZj5zjdUcvt9sl8fM5cDK2g7awhfsa43SOG
BnGA3oJRr/zqAIkAyZmKOsqpoAH3vwnHZIwiRYCHaROjSI2boM/fLrQo6zHJZ4xFNHcTXpvPjG6m
43dkGV9v7lL9b8YFnlHDnt6FiHEqH5DAptdHRvmwcp1M1K08TOaZvxQgdG9XYoYIkfz1PPUumn8q
M0bIcHStekoEhNvTNrUsR0mEo+aqMD+yr9Wzon2TUExjiW0gPVYs8tcF5Lf5fGGj9BRRinnGUP/N
TMF0WTf6kdc0foRxoOKYSopqdfb78hD8r6P2mS//m8Uhd96+PXV61h6dM4/NZkegO78axJQswCwh
fHD5o51IOWERhhA3cfAVhHo4KHqJd91YPuMc9ftNklHkP4RoHrZWx2JZ2l8P26Qjwt0bD6KKazR0
yWhY+0861g1BNcZ/dTjO9ifHQa197YSQrVTrGbJXBWBc4h0AwCXJW/uwAD4hR7Lvd9/bi8ralet0
OEOxASvNtMbTw1BbEL9nel0L3hsqocoI3FA6OxNdPifnFUN0QOZ+tSCXn/2JB/jukhJ6ya4J9Jja
NNLVAdgvafihRJWFSbE3EsxrgjRaI0JLQwqAQ18Ea3V069fwLjjSl7Fo0VdNZwO1rQomtBSPJ2iw
IGzqiVVF/q5p5+/UAGl0TMI3aoy/W5LzjcBmxPyXX+XTD7oJRm245/x1cnhB1BemXTuKDKY7oyvn
OWVcyUgLz1XTaAv0HGDKF8T8m9f9YUSOMrBmrTAi8YS4AZmXcIWCSqWwJJAYEK17CYmLni11nPQi
5DymnZyVDRtATzZTmAahcoH6jcPMFjVWXwBzad8atLJ+NTJjFEdtGCf+p6uHIDwF/tV01ULv2FCq
p781ljD1cRg7bsI4Agw+W2Y84gckP8icy/ADRVLpMpPTeoSFwF5cbEc+jvb+W/Po7QGJfK5VqhkA
uAFLmh8G3nAdspZyMkaZKLrfuESmFeoXyYFMZEYIwWtR7TnEFrQaQrMcFBc/2xiA/IQCur8coMp1
lU2MpI9igP3mBF+n+O2jGDZ+MeC9pq37Zhx5a3N8pPIKuDL9q2T7XHpJ+8AysKbXKFXPOr9GLHvY
RtsiYkwYCF3b7xjydQ3uVpTtIfHN7fv8xfmQs/8oDVNL7feH/1EuDQDKmX+C7+kU4u5RZuu4Z+Fq
S7oVLYkcO830PipXxl7ZhfTTSzFBEr0dVOcP0PCD/BrzS3sEumeU+jWYoAZ+Nwp5b5zB7h6N/WGo
l/jV+b+lm0tQmCwKfqEPyKBvkRP5O4xReewelil4bRRmdJwdgXPSG/j2O+6k9P2wQyvU814SgFao
MB7070Q9v+YpbYdR7R2ccpQpWX7bnS9D+XhLk1URGlACyWAcziwCsn4g8cEnyDj/HkLCgLKBbnmQ
TKrC+mfqCwKGWr4bmpLbvADPoOgkrxh7ysyHWC3UV0l/aKANG7lNBNU1xhQesymMXKO0SAljnKyX
w6a3fIC083ebm0UuV83Z2hZJNg86FXv7n243s/RGkR7QKBd6koXFb4IV67WsoECkB9BiY/Eyih6x
6zaOUe8wdKX+mGxFaev++MHHqltRZ8PAPtySr/NmX3HeomcyT9WREcyB72yzuhulJlw2Pagm8SxA
nR1QLOashTN34JGNnU6hwhlbSvn6QmUNxlnBpY7F+iFJiL02l8PzPv3R3lUCCx44Toq8bvosYh8O
rwNOtdZC/gdq2GagRk0sfIXh2pFcy9WufcPZNvi5BX1vxi6sV+CN8ltJuOD3bItzIv6mO3sABvrP
CbuNBWO2+Wym0OIUS/HHC5ctRJyGr04t+P+CIGVf29S0+RGhyhF5MudOPF9esZjgmkG2ibNgK10c
JS60etfKwMVT022NwGURsPiwo1I9F4b1ii0do5zHl9N/1BtpBP7Z5dPzfWd7FGMAisT0nCdc0xDP
0wk1JGIVuLOOTe9AYmJbxYp9fpG752fI9sMUDeAqJlQ2loMlvNX4rD2UbGShWXDJO8kVxbf718M/
XgtTTe06d+b5vpRYG5nsMvyx794tWqkmkUI4yk1M/wquEbBQlHmDJMboPNBVM76+92d4i2Qr7/ll
8nABVafd8gEXPIAinEkDtqXoVXHodNsn3UwDse3OmPdT36zJBFNlkeINUFra3plCv3IQyzLXM/8o
kL5fR6ZcypkEnq1OWlYan83URZohwo6gUdvy3+UL1e1pDgSpaWd9kku2qnvkEpR1HFI9vRuPN39e
Fk8zBQIG5KMzkR+N3+qEJB8naZ5pK5gm9CFBZxCTNmc9qKMNYboVYwMZOWwOsG5hgxPbOwl3wFbR
gEZN7zcNI6NGdyLgudcoJ4OPq4kjWjmkWtapGCbUjWjXRJE5N2+mTXvTQB/LQ5Yxg993OIGNevda
C/FUGnOCrLxyEKiwfdzMNpwnUYM55/+WhrvNr062wS9ocrYdkJdaK+ALz39g33H/1UUj9YRwMiMD
3GkTJcHBRIS8aetp7ys5uLZuIGx+C+ctY3pHOYAZtEyhNdCNRzs8cCMnBVs9Gb9XviOlV5x8Di/F
/Qyo0+e0xu+Ha88wsFp1RwjCiiDuDUqlCu6YRwFi1L0zqcN47cLnI9V+GWpJ5E2SaIINDL0Qsacf
7fXKc1JaPrCeeWFlkfa2takricaep6yWKOQqzt3qtd7nZ6pRpu1Vz4iWgrb4Hsy7KNlse78ouJLF
RgZbzOxrOmFgCGOMzh64OVm4ym+aZCZfd1UoFC6aIs8R3w44HeWLTcBuvIk9zLXGFuC/9XxOv2UD
EFk/57Lw0vyrbDit1ySoR3BYoEzdw6VXJqs4NFukQ4ZqMXRGHZqqQhRZrocw3AVOOOJwgQZvtRUt
0OHWSoaCG11M8isSf4W+m+7FPTMGwbkTc/a9gQnKUEtabbOuJzRmJaBp0X6P/BFLcl0dzZ+K3O0M
/ninFVd+IKojO7zjAgeLGAo+v7K4m9bX7xI5NgdXbDIEyr9nsXQ1H8ORnC0weqlLC87le/M8e72u
8I9956EzH770OqN/XXLBTnKhnDWuiJpXPQ1n6N+sDh2RcX+7PI/fjOkS0Ol+anDAgdPso6aqbwVN
7DVmc1LOk0ur9KDs/s8dYh3js6GtTLArqs8Z98crGmXVegl3s5rU9SOVWj4mf+HeX0cte4PP/bLk
6dgr1I34xbwwH0sBBn4w2CqjmoD9MuM16gMx895ynIYd5E5qUtH7vTg4qEWVB0HnXt6K54u66dHL
RJWsm7VBRV+GoiWKrqeRmw8GgBKYzULjN7KYfNnQLqvjpy8LuAZ78EDobWTjB41c9VA7+3Uh8QyK
Ivo5ot/jhYErJaPV17So3L+zXjfxrmV56BsSw2ZgzGXBZDDvICF3p/IJ4Xl83uZ6jPtwhd2MHHsN
LMV2tv4S+BtknvlnCpM6HxOqqzZdGWw6FvJ5lOVEYY6J2YsJYlsNli/yxjZDID/PcA5sKH/NiTc9
L/Ec59waX+uv+tvBcydAS3uv9x5GOMMSgYhoYQn/f2UdMoXSFbvafLMTtzS+7frtnxSYTw2cpyYt
AJeALaJ5dbm7FeP5lnli1gIB1wVf12pBOGez3njg91T9ZBTdPNCK0aydM9t9W1uakp7tCAMa201x
7l8nN1UXXrN25hpDLwqKuWkvisv63c2O/KcVKYyDgk5opaP7qc8miIYEcNKSk9kNZoEBrpkzuYzY
31LmJAeC7Fu4O++zvytclqHa9WXb0f9xsiQ84qoC660kOsh+zR2lrgRyL72xfYWXzUTrz26bWeys
3godgYrXhA9cvssp9Dg3gnjEko1K9dYFiCwqsVydMoIUynnzjGNvHb+qAu1zhb2WL11bBaTIYiwn
FYrxm03sUgQ9af21aalFuPjtBE6s1aV4ZIEGi7JUfeuNnuk8G89Wf/JhsbfG0AMexqC6gJ2M2lwR
fHUBQ71Tj53CR4zl2YDan7HHhkIPzAsgtMeRiWx8IAnneMBFbzcCQ6nvSeqix6TOwsYWniWx9zpd
LrKU0e/cyqwptAdji6hO8jpdsjmxjGf8ySsUnLlV+KHd0Y8eziGyguLxh/6khSYRBH8Vt9mP8mOH
nar7E+u7f1i0b8kuHF/epgYf1DFLeU+8+/gxahpNu1f4uo2SjajRndFGg+EAvq4NbhXcagNY6fFJ
1JiKMSvPlYJ2OgIoCFXc0Dv38HImzRGkJ3JXS9tWriwLujuf0v7Kn0+f/WByTsmbNalVKiUD3cF/
M+h/UUoLAqs6HkwHBXkMs/XvYGuhVW/AKMr6RJyNxtIdDD2gHjQRuZN7ZxR5qwMDv8wJJm+KRMxe
WECTASOdq++epwQAZ05sIn0ZtpkdDwL5hnWL/LOpDwtC+dkTonIxmoaC+CHDmQF/ACC+GmjOSYQC
l6pILo2SKsxxYyozddmV8VcjjhKVxIejiGj8ZBCc6K8r8JBhXYYSx7wSJaiK7e33RtoL3Wh3HsW1
m3VKUGEUiNeZvXB2k2Cq685PWaJBgrUI3jkAi25IVOn0TTNDHeAzKvJD2C1VpcVUmoic1EskXMug
jF1Wh6vLrqFLWI+Ze85i/caqGLwMQlE6VsRFzuo+htDtK8PqFoS0+qCRwsX7cDH4wLlo1gFLPz0/
T/TzYX+XNpb3cgPVikDipa7W/rVTzu28v7nhB/tYlWg6Y9N1UkTYNvKGIanI4TH79Ffv6tGfczTR
s6gWpY8Llw8v1c9ZM0lSKO5kw/9GpDO8/dZOQiuatyIdh5TycdYZsf9ShJvG7AUh9GhNR49cql0M
v0sE94bMg39v4AAA2v4pgXVn8bncv2I0yv2iq+UCGNGmpR3orylZAhsCG0+WYiAwR+2R+nzWuuyw
gyVogicKBoIIXPEqceeu+usIQZXXIJXUERxB9WjwqFjr4j9wrEAq8YHUXQg9a02u6/ZCR9l7cpSJ
FPH5evaz/UOfFoBGIxvW7Dtd9ugrmauJzFDQ9ErDvDPqGCwCAkXccUFUu03iacZsCmVZbBqN2H8E
AHri3ldJYXE9VR0z2itHrRdNMVA1l90yrn7+sfAAwzVsPA94dY3gy4z6z2vqabrFFPsA+UntePFl
5jppO/qCyClEDz7yk65kfbFKawGep70BICAsaI3KUUAchEDuVHCewSTo7St82Kn9FAywFFnyoNTU
fRdFSGMy7+Uo5W12Var16MV1KZr9gZuYAQ0LFNiTvRO+JHkQoF3WRy1mLrWmxMb40hWNQTQuq94G
ySFR9yP0EwQHDd5VC28D9O1byezID7D2HBv8QARw/EHi+K/YRKwcYOMICuMWaxJDH8La1v37lDi3
3x1xgP5C8qrZcz+QDxcWNhn602KHQCxVJ/9iGQOSl3zPRw==
`protect end_protected
