--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
DK3oHhAdB4V6hyGcgXlgaP+vvPm4ewAzRnoYCsoGTm4hPDEK/U4Wxp3KtNx/Y3RiXTrfboSxgTam
i6EfVITp8jISsjXP5xmneBLMj/eiMaO4ju6jwrGJSgzK0ujpSm9+ZIm5xFxGvj29NUbyb46wRqaf
ItsG16CMKEm5D2w5rNUP+D6wDiYy3an/B32TykSgnNKHFNCm+71HG0Qdp9G83826Vd3TUlsoFWcd
DfL+g+rcR4tny5NPJf3OLq5DjESsztc7I3NFzWG+otnT4o2uKKWJ4wLZUmTOgP0fWNdm38KksS8a
+VGfdCCWnao0vpC8RiKKHex0FZMDvcsnPUQdxg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="45CjT0UOD3Uf+Zr+ZYsjUpSDamKtDbOurm4VSV9g8ck="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
mEjjBNkUpnknowpwVTxHCGzVz4OBFmbvK7KNlG+SSTwAIMhY/R5HJrmkUClYp391KV6PDcHtZSdP
dWVM1Yb/lKIeAlQOohA0RVA+Syc/YxgjvsqmgxeMM3g9YoP+KshlYNVcRl0L/PDo+0nbS3u8xmFA
2Gf/xb3omfHnhAmLhOHqLanGNqCB2Ri3WcQNW6SjNx16rPgj836dkN4mzQNuuxyEQH+lZtJTYTFl
+xGLkzBxBIMJ6AGgmk+RnsZ1V1dn6kBf9JaMV16TUd5P8SLq+D3ud0GAlwE0I9OCF3xpv/hnIwuD
tESAqaSSYQZXB0dvXaIu/gMjaq1VD8mW2tNMEA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="ZEZYHejiY3a/+igJeBJMIdE6cs0jOP+a3e6vukUm0Mw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3968)
`protect data_block
IaKouwdiKhHNh9Rjh1dZHg0OOyk/jVb0upBDUoBqtHZytizwF2hV6fVdMnwGra+7Tmxyro1bt671
OJX5USP0GsCN2UpU1bu0jo5cDUmsPBAYdBekcO0Aez6WJ9r0OhN6BmYCPYlV7msE/lw6BxvPcEf2
E1jNSzoqxAkHmq2YHRSRjPL1rUFMAe3Re1dGzOs3wkaXI3NUr7tP+1WR8UCpDJGGEZx/0afdgZyP
hkhpSRVLCgxUQFpS3PdrlRqxY7mBQquFiI1/OHVlOEdFzU0DpAqG6whgMh03dChmUatqYvkRJCUo
d1d+NtIeSOj++5M6shKmQ4rWjJTlw0pTpPh99nwcAgDX7g+tlrqnaEb/UuhHahuwtcRE26WhVfx2
rBTbbseZEY4P1RwhdGbMPTXXjjyb7uYVTshetap40Cq0YFHIiB4FarMlwEtb7fJY/5elRwOTB+xb
wVrRn6guRdjwSBqHWDt1/V5X+QHy51Cx0cFzuPHvn8Q2uprXdTRrhzVKmpe6PBrLAAI/SGbnHYpu
4mBYXoPLvnWAZsUeyrn9fDwr0fr1jAFGyQIKaDRw/oK2B3+j0huyLdCbj22tsCVdjjSx2M11LQZV
gLyiTsZwhTXWSS9s0fLkU0VVGCP5SoTAHCTxtLPSuSE/5YueBoVlzyxyiT5/Cj/EnXuai3ovkBp4
pzkVYdj6me/d0GcE2Hq4KJt64mhFnQfzPLBcPTuGHApI8PLs9Td6/pvZOD/DMUTY9Poz7ApjfsRG
Af0Gx4VNymdgi+Wdj3IaL0U99jUPjUFTylhesVxWzeMXt4CsmGmerEhP7cNfKApwwJRMxnOXB71E
28NxKgA3FnjaAKzggXVu4eSfc2dqjwCRFQPAgylKnvi1zgTHYgPGhaNlS4f5/+UJz4ijZRM6OK/B
qdKtCC9y885uBbemu4W5RxQfpkgRYUfHBnIpwYPje81UHnbasnNKmnWPQleekYV9znZR1Ia4XyGX
ByKoVhhaylsdUFS+aZzdHkO6+G+T7LpTpBUVxs70l0COO9KM1+aao4ODl0Otpuz68hSu5C24kJ/9
ipcEy4FOHvD1loikDIDQ/229cMyo5qS95YhJpLY6z/37Fqxf44+C72dJJhWs+FmWV9HEeNJZxt/W
mjnKWtqWMhkB3VpSyq4/Na6Pxekb2QYfnYvroWPRUDFQnqbA6c0juGCmrA52tTk35MuFQ3URDjOt
9CReVgWgOXPVACijI5PFFine4GDnQY3+rKChcf7tccCi6xX2ODTBlzq1H93LywWXgeGdC0lGUTH9
/otlQA1UAV5n83lV60AU1LDsawi0qpytdF0Pl0dNMp52K+I8r8zAMtjapHNYgtUtqiFvcRIcMVoS
4tKJKbY8LTRIRkM4wbAIVdEseY6wsehATzPh2byjhsLiQ+TCaXpU1jowgNmdpdt0j9VpKfWzP7iX
lGYzMpTBbqF/9UkdRozKg0y0/ZvUhtvWDp5alBO0xcf3Wv8+wAuajxt43NCn98NK8stf89uO12vp
gaC96CeF94mPZpBfDkUM+WNQhEY2bzZ0gHJNul47ZLtqWY5bvvCXk3docemezPWQi+le40LFO5/+
Tl3uaqDS0nkNyawKoLczLEkImxXD+Knmdrcw0pWJqYJI10YKdBjg4pcS6WDZCV4OpWBdlwzKHfZZ
ZGKBPu3MYqt04HOVCAizUn3GEyt/GYhSoAW9OEvjPlknx+AZeLMWfekPkuu/87nHH9k8vFKyyJzr
ASDT4kVd1Mj2l0auqqC2djbdYr8CdBlKqJfNFDnhqpVaIgAA6cMwL99iSRSASYCEqw5tsvqPPUUU
C/tBfs/k0WdHhHxwBqCW4pFSLj7QhQiCs5qITw6rNDpJtp0rodnbt6tHjoxIK+oVZI8uVhP8w4ty
0wngxGIjguBDOKHuGbUhs273OdkgAgygyMuoyQS2fSb4S1KJ6ERWQADB0qsu/pLvYIlncGndvpvD
tp4SQQ7cQXIVcODKm3mU4Iu7xufCueuOIB1g92XIF8BsrE/DObKo9SHevFXggQkJD5qatIO/A/N5
mglX7tMwAaRwB6hcfVlgnoSZtBK/rovTGqFPiXoWPJ9+l7DwOxIeMw6qvpUZNkWTJgZ9m161qS0F
SjWaRw60O4kXMWPoPakP/KWh807oFa2NX0g+YOR+OTN3nGmsIAjc4Vb8wJk/iwwI4DCYksNISU6y
a/iunc0W7fsD9fd6JdyqM3RVj4rMGVlpiaXDHGfaT2x1UsF2R8lVAgi0mZqNhQzBHLFr26R1oU5k
xHcDUaZOSXRUPtgkMiOEb2g0y8Td21dv8kWpKsiG59O/htaUWidJmB4u7XGp6GRplHI1x+QIs9YA
coNXw0ObD4OchvJhsvRBe5sBesky1aBXmj5if9Mi88ccYDv271LvJ/rY90qrg4b4bA2AQ+PrXDov
29EpW0+GsHkPGNSHSoFWKyk/UdlasPB7D/91e3L0761DT/aFWXgGeQUd5Px3nUeURXuJ/O+68IRf
U2ASD9BCt4+VIO9B+5RhA2mySpcyxlgVs+hIlmhzRfz+JvhCaxwBWY8BGaiYKDvqaoUnj4DEAs3W
NLxBz48nfGciypzPGNn58nmWzZExWR8fautJ6Zga77MtmiEXHkybNQxe77g5LipRYgPv78BIezOo
S6GtlbGr9NEYrmP/rVaXjPvHWznBoBdl63mIeA3+IKTW+nR+rZua+H7n2DzeTjQBPIWsDCQt7+IN
XdSGDKRhPIxTUQQ3GFslMZqplZJfgr9H9CTj685mUoqixIH3dj4AOCddr0qoK4lUlXOO0whu5Ap8
lBRJxq0dL/gU5yp1GrRCyzMf8hzNTyzPoM9kSMDXFEwpacb/krFBEAG8nrCIezdD3pjhMeWHV0tF
fh399bHHtFPoUZc6AYIMpsfx4WP2TuSYzpAsVjQrqPKSrWhYss24ypGw5UvL5lpeF9HiP3EygKMq
I1FOKTFSenmfTTujeYDpHBUWV11Zu6yVG/N+R0oIbbEPt2/GxVTVZWyLffKq3X+kWSK7FmDUEix2
6TVeC2N8sW0DiX+ClUrcexL7vpPakDQUZAJSM4vPunmS4j5NPHCoZwHL3+ALay1eUyeRt7wqCgT3
lba3Tp1+ma9kzZGUrrKEyN8qMhamuv4uK4FjbUlzB5k75FSdqFs49WGJg4y/Vry8pl57iERcvQCi
XwGrnmyjZC6fRRFAaZD0YlKpnilEKcwc6qu9o1Trlc4OmDlRgkg1FjK6DDYGie0XADQpa+rns8tw
xun2ntzGww9vwDkyWyEcq4KhoTrhZC70TvrDkTvQ8CXfSi8C4ihs6TjxAFsnnMleHgl0XrQz1Okq
kMTgcqaL4ldQffuYotzuDpRlQfCSSpN8u4Ps3Tpjwbz+Cag0RKooyDlspQpat6Ze8D5JA/BFvdD5
KjiMaVfE4ASbjhZqXG5jVFsHsRWwsqUwg9W4g74C9VYRP3ucgO7yBDwIORjDl+RKYhsbQSD0A2Ji
vnmuyrWyTkTH24FYNZaFT5z8xVGz4kkul5LypxXl77tOKGal8P/0ji6AOmFQAIBf5TuYwh960n8k
IerGrqwjtfpNsQNZC+xBL82KWmlrs4nulRjafQD8m76pqFzaq4YU3nubJXQl62yfx5+g39Z8DK/c
ptG6Key1Y+kFh1eCgF4f06kmqTXQIQ1UCkYu7BsV2pXrKH4xkKV9PdpAn3/T+2W2iXOtu1w9hsEP
9ooFz6MVEkjpn9bZ/sM97C+zGrzRD3wvCCooaRVdpOpNwNNtghQwRufOE6XitrKO22E6MijNLhIv
Gxljbaa7ddg/px51ki5laaDQp5PANopTC9oKRt28jDobOQyJk5LISkIlSyqNL9tOMyFqHQt3NEie
0OU2aC311XGN2qYtAmztmvsTejOQyolymqtXeBixfdSCmYlyVXnsLaTQpZDHULDHkCivOy64GdYY
MoIDktlKElmJDHtgsIcFNBItMmJElRJfphWVe1Im2ro2ZLfUHRVVMDy0nzSDxxwbBKeY05P1yFUe
td9yI1/n+ABvCV4rtvyzYSiEbr22W5gpEDpIAjT6RG0Tga5AwRzXfUUgWDO68EII8tdtCwCxcIA3
fgYKXzY5WW7x+BzxNR9VeYcYqLHDbOX39wclhM7AtEyvouI5bGaFZB49yYyne3qAKUNm6LGAKl8x
hPMosEcyFpewlUcW+kftQtpeeHNRlxSNf4TlRRJq7iYmljCQ9jnsY0xrX1H8QgUngNah6nAwPapK
xlGflXb+BlIBRAF7a+6zhjkpXzOJsLrQ8wwzuxk0ogEq9Gno/Q22jG5VUUsmf63fp75R7yNCHtbh
zDsBUI7J5x+uhSIejYPtOF/JtLcj5+b9XRHsF4ukP9GVg9agAL7qLZMiB4eiP5G9hwAzSWV5DmhU
vjFBSdRPsedtUK4UYPbE04bd/IcYArbVmrz86PtjXv5dDUD22K/sVeDq0mEqoD/+P7wy/grXvGok
RAHwuUAeIQmoLR53PezxNjQzWJmmMuD0nv6TaRM0H+9p/fI4gi4ih1i6N1ZPPUmw2vmqZgj9rrIM
xrHvvlSdAJMsjnmAsDFM1rrvUfy0GPEFh08oHh/3/0IQ07PlnUrPb+O4qH/vp2GEl2IuzPEXVpNa
Xl8sQWQ/G1UIpdz7IkYGP+akoMPZcLnKxCn/eaFFM9QzOs2a3BMKvnYMQgZNtns8Sm1HQzoKVPeg
XQnZuFJdna7eym8oi5lm0jOhXHtd52FgiFidzntW3sgEy/kkH6lVr1nS9613tXV72DcGXTAcmjBn
Egat3n7JNbJ9mJOmsTJ1zXlC8TJSi8+Bd+w6Oeiq17dS5C6ABZWAaI9TsmGdAW6uGyPsnl6xNXKl
JWksJ6mH2a3Y2yPId8OucRqOLY/eLFARr8kxxX63o8/3PXY5kknXkT34qFjx++ZiZCwJY1WUzPQ7
XVzd2ugLdZQtEeip1IO8ErFTmkn9rhsgPNH4TdlU5kILZspcA5YHNx1+3j1ptR2tf0jbrSF2yHsR
35V0T4Sy4Z+viY0ZSIpJElywnNFBbm5rddeeIWoD/uDSb++dMk0UH0kBMF8cfXBiZEelBtJCJWNm
GKQvStIyeiYdvpCfueClCb/aEsA6C3+ka9M+9+wDwvQqZ83GTVaM0uaNv5rz0Nt/F5cTwN5XHcqC
5TadS70PUfS/GOPCH9iXZ3ztoJ4CQH4ywrUieBdNAfHpTI1Z/m1AKTGdGjWP0C3Xv08ArzOtkhPI
ItzH+Uu7hNhFCR0d/TIUSgJrc5jrRCwkA5ulKtMeaQUpLaw=
`protect end_protected
