--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
gmhNne2KDhR7d84xKtNvBrK4BOYWI/8OOSnZ85kQBRwxcAIeuwIQ0Rd2DwBAb3Z14xDwRv5pFm0C
TlI5aac4QOgr1miJWzzVa/NpzJoWrOVZm0ill2XOK3ZrrtY/CyWRrrP8kVEQMeFyawC/ZSQOHKwb
rnRyiSvO8pw2SR0WeUojCUTVCxAUPQDHX1dSMaTxuLG81TEwLKsKOOHwOdpFFOwENZCBwBcQzMNi
e8qmm83iwCCEf8JnazGQtVV5XWScqkOOZsx312g9BsFhy7hKzNNh6VwTyQ64uSdZDRZluj21FfMl
Q5GakWtU2RZBzoLcfvmQ6lbVHOrtO7mxNAlsDA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="XSktxA0tFJyUJnxropOZWsdXFNoTFvBmyYMb/CwiayA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
Kd6mOSvAYrKtN+UQZtLVz+BEp3d188wu0JC0PzX6Z/9n7eJBJm/qKsQ///k578phtkqsANGQIlVq
7IxD0TnOgpVfk6XeMAakDSslx5IaT3HPFBhypLHrzHViQ1yVCjD9O5g+hjoVaX++QQbbV+0N6CMG
lNnLiXmPRyQa/wa/LNNYDszHJ7owrVyCmWKY+PIURklmls3G/qSw49XRkJqCdxJBnzqUWfi29Uv0
XSYSxYcmCCHjBSbeO3QEIRx59rI7QLei8cKEMnjwAXuzh7fdur/0+FwlKewE3djbIkAXH98iXaAq
Up+gDQhv8UZxyjkiPflu7Rb22xCUwkcEl4vDjA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="cZ4Drc3NDdpCQrmQ5rR0m/IvZk4lJAZMmk5u03JqR74="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2608)
`protect data_block
X0ngnYKx8wpe4x3GiBWS9STPEaBwifDqiWkQndgUWuuGPvQF+Y+NQIK2uplBd2tMOdD8jQ5xhpRB
fQQWGyIZgZuAWuscdLBvBjbJratDHhnCnl9UUD3VJSSzD1U8fMYKb9UdNt2T8c1+QwfS2/T/8l95
l/Bs/3OcB5KIoz40xwAkRgJqBB01vKleq6lHubtIqBlZEmQe98gSFKz8f0WeGFJ4g1VeQZlUo+Y3
l+9ZTLvCMSujPKuj+Hi1oNCMTs8srKxKLDrDsXTeB5oPvfUWOrtd4AerCga9PJnUjAAKDMCYY1Kh
OxXXRLiWy5AlsrSZ2zGfaJ4BZbe2GxlCXP6SVZSDfnSc/aXeBFjfEggvIl98ofQ4ubjWiUoZZqgi
OIqEQRPiXF6VVTOYq8dmqiUaTOLIdo5Py0Veo9x8EsEYXEFrnLDy8joPF4wg/S3P4ZmT1d1TLdAP
1H9Jxb2LUgKnYJANP2yORF8fyDflIltbY/CBOV47w9MBHNvmonGP9Nw/RxHh4ECGCC7pcEH4oQ3G
JzrcYiYSB2wkoSBWSZErFL5y0cW3M5KFENIiNVPznat0EFAtd4+JF++Jiz6BIDXdNOK4S1IAGcxI
Md8P2qCZdgOus2fpLC/A/Ip8qb897rtT0iQ7uz7yDKm3Hpa3h2MC49kKhDfyF/g3jSlcdC6TpQfF
HclCghC0fjBncRS+ee1W1Hur3Nhi6qvtB+c9vNwItPwTUNrfa3S0SYh49sujAZi2UtmFBQ1cNnTi
BZ9rEO5zqEHoNOMghOlHPoVvriO1E2pN4W4t76ak8HcRvhyjnyRhW6soyYC146WvgeWjjhMvkVqy
0srQdnMXL5ThV3Sl3RpS9EHEyGlQ7hG+SS/5LTi/ruqSxBVqN9GC/Yxbgo1Xs+dFNA9E0Etk8Uw6
fSly3yoB2/2Sd37FBvI+SRxDeME7sNbBptYpQLdmgmsynWuUHK09GgMnoKW1SV5zJ0emBF7SLLFe
vC/ZpkWaLqlwHqsGcU8N0cUwW/Xb0uT8V5w4OtLVHzn5aijRJE5UEtqdrUimrkbTQPa+IDHjzSXT
nXCC32puujNuE+9p/Zu840RaqVT2/c5y3DyMgwegcaodabZseU2nbuiIa5VgY2nQNdsTM1NfihCx
dSNRKBoQHLKeIFnX0A81rAnRtrMie1iZ/fHYTf0EltLeT5wIgHLrYW24lNCcG7uJOpa4dVOD+scm
hnrx8un3CGsK10agD06bKG/8v0YPNTbSpSge+OWjVBof9mI4sEsg62629EKVpvhVJrVwSYXaUurd
cYJOnPmkChsbi8KQY+0KxCoJ8eXukltD3HslTB8qrOUMFZ7UDGPi9G3tCbujl25gR1sTicW46u4A
8DK48ipLG4SskmSjQzf3TDJynK4rFUVo01Plnh+kmXCwUvmUjUNaFP26pPBZmyx9maMGimTRldA3
YdffK5JsuW72rjmmsJJFwh5e+FHXveM8w8uGZN6qHovlsCsI6peXtzEOoCppp0rRGC1Id3AbOLHS
YGeMYlB6gs9OdGUiEp6kMArbUIANhw2gyM2kFLzssnA3PqkK1yWlVm26JKRsn6lLbCI/1T7yz+6M
UkZ3l4ltFz8WDS5SfUuju876nvH1UzsPkR9YF5pVskktXWFNvHStBk3aBU2tc69i1dYJIN8CRq/x
KmMxxlzpOFAOoOsHFkFkzwJsyaOkEuc5PgoN0DgwdmDsQOfpsVSWEJBiZf0PCBloINxTeZDuD7n4
SdXLWCZijAhNehiFDZ43yE6s35hoW85H2QWOMlpJ5WeMjDZQvLHHeF7t5e+p83955UKniUc/cmFn
GD78s0BS2BCSF75JP8O79LUOkpiO/tUTygwUyDElSfsPQqIFWpgCDwt2gwIHHsLSJ4hDZL0tTy08
4ln3wrGs3v8+WrNHzg4Pvl2/hNkZjRnsHEi9S2ncjlTXL0DOWz1/KY4o044bU+CBUzeKMLc278c2
n0nmPMHFhd5GDzX7UP1cur58AiJFOzK0AHyNP870QjwBxRO1QjEuEOs+ZIm+Ck3+JzHLkKG/TdTE
/io5K03zLNwzpgrIuQmdfxtK+PwqcUZf0HVic2c2YL5Ir8qyYbSXWyQqiHMF7MKAt0+a76JXlU2F
4JvQI8pZxnEBwGcEjQek2gr0Qo4xTT5XnXAxKRR8DR4ndCZ/ybRFb/fVPhZJtmRsa/OLBnhcY6Ak
p6hxsW+uep2LBO3lEyAyDapK7t0Uk8G0yG6CV6oaLW3eEcIpEJ8TTbZeL2hghJK2Hrwt9nc5aofl
KrRiXIKLqPYd1rynhAzXRpwz6vMi4xqFH2Gmt/TNDhy8FES9yZZt2yi2xigIhdzaauWW7QznpwLr
a9H8/9FdLXAG055EghYOTcOFgz/rkLySxezhX/92PSNB+gHqO417x4lSRE3gGf+Kol+95OEEa5e8
WecdzanobZC1fJW+IHGKgrClkpECAleOTFsubHvuVHpWcWoaaWRtmEluBYs5g3v20rb3tjF4iC39
vE3n8kZc89Itff8uo1LV3SAygUbSCB13uhnLJb5NVMfRdI5ZpfA147CNr7IVsNt5JqDCvNKjlMFu
p4hy2FQJOI36/ag2mg2rFvITvznR2qZKMwMbgAm97ZLbqmMwQh/zillZt1lYJd+08P5hka4zRD/x
UpJESy4WrCHSEWu1ROdq527Rx6scC4QK+vSWtFu5lEmaF7HAQZJBaxNrAhWrfkB13P59c3ShCgce
gMtTnVTKxqIqLP6TIn4gaFLXG9/Ydvupk1FPI1WUVBV7S0dl7JNLznfbuJg5kNdQkramAvTya+6p
cwXcbL1wc8QfPsulxvcMRNhE/RjkQOKB5d1zEABaWDVb7mn7n6yqfs+zVg0ZW3iAIEfRsWWPZn+v
JWW7+bQEKZOoc+Ro63fDkkXfNMWhCWAN+fPm0dsC6pkfcDhOSLIaP7r0hL7IaB0l6N507PQd2BOf
xg9CTvJncPchBPHZvrwwH7swVRPeGQRh7SSo+3IjIyrTxyze2udeqiNtxVvGK/LWvHEYQ/ZLdu77
ROsRzgEErShA+B/4MIoxY4kvc96MxCmw1llIcjjt0yZSnzNdbE6jnz7Gxlq4t4FyQZC8dZCDwsUj
8NIynOc+zfv92SzqMtyHhyK4u3KSWV0ciPGgRxE7rod8ChvtHCrpSW6dUnmklM9xCLpiYlyJ3Dha
1nd54E11PIH9V9KK/LAgOwE1H+HDQk14G7G7D30TkABofRl1FVcokJgZWVCm2lnmuXLUVmZBbH5I
DloSe9qaSFTZU52DS6pPZipbUCvOEdAMDk2LlrjAQRvMk+/JR1dT4loqyngR6EAcYG6QbLrtqG05
S30v0Vx1YaQOdusmroEevYpxh88l1tNmkzp6sPsQJdPBIWsGnNwkcVamZFfLYd75Sw7hpjQjJUGl
QPt5QzK9pvcoJ448skZqCjYgt8VrgzaBAZ1eR+Ds7IDIkeAzt3uyriPgwg==
`protect end_protected
