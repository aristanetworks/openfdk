--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
kH38OBX/XylEVXJP6Vhk7C50uW43TBZNTBCQGpUNuvRxRmMRHYX+ZR89FEwT4frsf+ylzBCs+3Vb
RsHVqJ3334EUuxJW3NBQ2Spr1qCbGempMqABx9ULlRUT7U6n9pPG3JT2ubH7p2Ho/snpNn8tVYcH
mawmIVOyXTbqitguIEThnefrBIKF+g2PxPjH/DHGoO8r2Gy1THxndAK7hfJWSL63OQgNjrtCP4Yh
mOH05tEL2Rwb4/4M692KL5534UY0KUWEwWKdxkT988iIXs9Xqblzi3pVRiKUC3Kl2seMP+Sc6nGG
d+VVUYaDl6QlwNO4/Bdz3TurXqcNYEAhBK7bVg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="qcJ3paajogY0zF+ZAs+Vxkc/MK36aEkwhMKhAnPF6zY="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
bGUiRgoB9AwxEevmOZCW+xRwODGYMGfMtALbgtuCvSZHIE3P479qIFsraod76Q037MXB9Z1tRXtI
5ZYfLAHR0PDR412rf92W2FiEhPm+11iFrHak27oNW82nGYKhrnVAv+FW4Q0gbCyBJWdUFoyiTuUS
cZv+kH+pxdUi9boUpL6u1hG+uCR0//LYnkGHk7aP6CChSdQjgvfRosmdU+4LWEfvvbDg8quwqm8R
rSHMoYyqTxXTEiryz3lC68yoeHlpyHUGCYqKsMtF5A3AXYufNmknZJK5tyNWkdWH/GOxpfABeGbC
Vsb8oKrx0fr2gk3/G1Er9hLpWC5WY26Rmni1bg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="G7PkQXZ5TYaBfzTH+HdTDvFukkum9Ig0UbfFUemRBcs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21216)
`protect data_block
43QSYeAYI7WdjNaGKqckTPJDlPExCANE2EkWThwYJawUH53ddbwLmMSkSFZb44C0Y4KiWIOcKqSi
utETPwB7qgYv7h28xBTWkT7BvCc1KSTK2eqoVHeXimZRPLIZu0MZT8MuZubJ/QSDq7OagHg5oDhX
jugteVLulW/2Blb9vbPL93Ik/URoa8kg22hVUDqOZO7UBU0HRAMMGcJ1uQ4nGdZ9VP8J8WW5NPzn
u9JuvyYGLh+2/FNNkXuk3zoeGqNWD/GIufQlFEq63qZJ2ahtu2ygqnQhyJmCZ8Oh4kXJtQSiEDvC
XJJFD5wm/jQ8IjDBbB7vTRX/XbYQ6ZrnjjcFpbAT6w2VQ6EzrR4efoj7YfPrZgkCIFO6sev9fldl
aOR/PDwXWNKo6ob5j2A21SwaAJO5cPQRQ20Iz9/96Q6yYY/nKloahHGXYXP5wgRbPkm+XRiTmgmN
olzW+J8Su9AOo991Z5UD0o7I7tmLoUbNvRSOE8AQU/Q6D+NByVEShvDyVLjVNpxLyq0Z8QTGtQwM
TwpFkl4NQJxjZ4oDB/CPPwnQCEt4Hwhbp4iGe4Uaw4lfnCUH4pdV9vZWhLmTyKTdzvu5ESS8GYtB
t3K9W+WdNnb8kQoY5oqX7yL03vtUkRJniDlJ/1agOKXwRmdPIZwoyV9LaDeXJ8eQyYUwOTaZNsKb
eshefiX76pxSbfDmuObSw/j/UV/CXJbEdUOdEVPxKPSgaAUxf6FyozZ+wnRzinzJMVC5SLJm4uoM
mu0oEB7CAF4Hqdql2yjINjAWpZfR+zdMuGPpdOnTZsqMNcQDWAswYkxlctXwju5QCcAaKFPeK7UR
YYoEnW+ojK/IOVGxfwh+x58jnvO2uyIAJH5mm7jI47VeOBPkK2zthvi4ExY3KKbf/LhJSByXROXu
5ZREAAodoMOhSx60IcWY+587nlH3dReTcz14wBrI4rnXCCP2g9gyp8dl1vMOuLc/toD+RPQ4LA+2
Ykwu4g3lWcDBG8F3EI5cZoMgIPOOrNV6bY3GkZw80yQrExiq1KfqxmKuF5cAixEQrZpTGbzaNbjC
faNZ7xgV3M331EGr0FFKU9U4LJtyBPdZq9pvYw4H/sFq5J/6CbvX44OsZpTHJQjCTIcO3KNFUKYj
nmKjPaEHF3o8f3tG9pP1+CohzVifGr501Ui5No8bDPyC9ip9V8tLVD7UqVkqk1cmlPWeIQMGksVN
27IsHLe7XrBiUDdE82PjzwvH5CadjvJj1xzN7aljNpE+J5C1g3R0/XFTdpXv+7MkZXxfJeBzbKVh
lXUfeF69LYtyK1Jv5WUHKu6tT15O7UGRVJgUh1ktFVWuywWUHjnGF3sRopehFlxKi99sSwyGSfFm
QP/cq4k1bs+x8UzEBp3ye2D2Bo58G6Hf0Z/fz28YlZArsNAPPaJofiQ0DquwSuc2JIATasGm3EmQ
+Vn9Bi+yP3lfmUYbj/PL69EvdYsGg0TqdFAgfWROnxqmfpdug2V5cxltjA7/A+TL8L2itMY3eRbN
zBWqApYfgFhT5JJI5FWR3KKaRvNvLOhK8WqWCQd0xEffzc3n4cBKr1Ngn+INvr9ao7+Q1ukpDAC2
FvBOD0w2/D+7bzuJ00sOKdTmAj9KcBrH0iaIqgWUoJRmBByqca2NUA/l7+zv2Hq5jdnb1nOkTAJh
RdWwWGeI5Lfij7NYrNqFdsdDb59QNzb7zsaOpeiV+j056q/IV1SQued27KJR+W89dQINVOux+KpL
Yer0u6wUU4IlYCG2P3fywhSg83EeVvzhHr/JJB07gjDOGEEAjOVVD2LgeNItGJSIaXUbpexJhqd3
v4fbSW2ZKmXlcTGd8TxAe85BtwR4ODX/q/71vu6hykPtvKTEg+l6cNs53YS5h7gn3UKbk4GujNGx
/SS5GG0vJjqICP3f4SoUHiH8DWoW29EdcbYdI0asyvGsqcM+JQIvCHX/X5LOHR6NlP+D4jR7adMr
2DnnvTUdVn+VqkIkOpXgP5WXldj//iCce+1845oOpaDiYQqJpqH5yt+MPSNb/2XisYDu0K7e1tN5
bPNZ6/wLjtYTk8FoZZ6QVWBN45pKKHw90pphCV4eYNi0U7/bEfAG3EdGPzK5wsGgB+hRtQL9BHmi
zUmulhwSltUdnwLbw/7fMJlsGZD2Sny2qqQixlnZBz6ZnbNc3vvn4sWfoDyv8DLt+p9/lLlIT/bl
PZffyfxSdzvWop0GWULau69DyMdKhORCEdt+fTUOOyJ7Ju3C0/wd4bzt32I7hwHPPPBCgqgoIhPg
t3CeXO+mBNrCELUHngvytKbUWiZmnumfzF1/Px+EjDDxK1wR1/V+DbJgWOLtqWvrdprPeBMzgGLS
pJvvo1sZj9bZ7lRUQP1CmxsyfxqkhwPhWKS81rvhEPk2z2vIe8SaNeow6fxFv1qDrjjobCR8woFQ
gjjw5FTh1gnCQc3YzvKHbZKtDKiCj8eogrOzqf2AtxRM7GsvVq4vAjbvPnrhogqF6SW1xmiasf8l
J4iTx/ENP6+W1oEXNM5pKtl36kolyiOvodo10juNvrccZqHOIAMsRPFgsymPdIgyx4E/8hNGd1H7
uOPQf2URoisYRRyuJVvEKwox/4V1Nl/d9PPstKDNBl8Gvzq9Boz3qW+2xPmDywc1gCOQx0jEcYY4
cZHmbYOhHlCHPrJOjd4wIcYy/nNQFskx4la6bwrgD5jFrUG7d7siVxnbLOi5wEMd1bgMl8Tmszbo
Sbi+KehUgy+FACgVN0hQv/dDHa6YuTsNu4cjUmFpmjm9g0I9cf4vQCpBHFtvRKxDqoKbutsp6tBR
wopJ3QDyUtjS3NlI0Qj7V/D0HY6gCkcP4n+JWJWuAzRA0qYJFvY1Vb2N/jonJB8rkVDZEmk0ATX1
zAKjn6r9cL/zpqZY2mCgRz5zjQYq8xmCC+cMvSUbr+cui1DBbolwx+2jIqxPFRuQGoyp5DZusocI
MYd5aRIwD9Xt6ZKdgahBkQU+8EC0kWWAUwxTcxRepNFfchLBY2Mu40pKZCk/KhxDVwcm1EKaEtCu
xvJSZRGo/pXCxbi3mV/Xtlimdzk0tnhLkEY8S4c+v3Oq1rLZSE6wtr3+34PQz7ksRs3jEx/Pqg22
2weCzEvFZQb2/dezhqHgB84WS8rAlnE+bFbkoRG4O8Bx8UnvpQG10vTutz9LD9+5wdr1DiKgCMbS
g1lNMjc0rlv6zZgojIrnWmgsmdPMe+erOS9B7pkZilYO5tBfKBgri87NEuXrLXOwD09qIco6AAzr
k0vS0harE40draZ477r9V/hsLwUFfB8GHfRSYGmRI63cXwsH5+b3PPx5/QQG33osoRj2C626MAcp
xgSEPb4ZwhkvLOkl6nJpUVntP7VwA49JvD2xs3A8bZMVbYIUGxNbOOa4Fn7wm8+cl0FCnub1SAi7
B6V/mkHfDz/GKaeE0abOctbcLwGoz/V8Lo/OdgbVdC4pth9lZS2W/syvv0BPQ9Ua0eCXD63C+3q2
t/ogKsIbMYFnNkKgqXqG0BwyrQhr3OKlhHE6oTvxRi1T5gN7Amgv/Ky/vtk7hNk15TOcsJShkCLS
J+BaeC4+XbnW/lU1vbHosHcM2Qz5TnCY+1KtpfFBhPASMDcY3sor/S0qPqUff3tSocepFHKarfz/
Rj0iZ0l7nzU9Jm04LkJq0k349YmGJdw8QjXX6B0i1v1N8yCccM41V6ZnPGLvk9dUat9fCyw54zjk
D1ZrPw2MhUgq8LH15IkN7C+vQvSQgkD7R10QeUlOs7SdmRdXBFpZ7ZFge+SpaBzSmyz4jnL4QcVa
nHHRjNywnZjH+ZH3IxDA4pKYKRuJRiOF/vZO0mfYUVnjq2FAPX/TmLE/YEXwNQi+a/XMlJh3Qxgo
/+TR9IJtBijQmKgqmOPstG9npJp3Sl0kNu6c5pi72qQJ8qYfJLDTi+Ga41KlXIVoyx0nHedUQEu/
3iP23XNTEB3gcQAxTpu0PP405MW0SBaiGQw9QIjn9bAgyP/kENTpizg1MNXE0nDTv5C/L1bGOp32
Ng6nhVtLobNYtAxlxLjbejXch2ooBsZJVt74MN547FBQI1bqL1foWcKfX74qRomre0fwzXdl7Qd5
573Ik0ckvNS2uvWfsTVWhaiTHoFesi2MkWUu8vkjgjqUaVt33eqPyeHKZ9FOazvs7BPkxdEo9ft8
G7XmM7WF80c+BmtBlCdMUosSuuugbRyQCY4vD02qHkX/sUFCPvKsU2j7FkTyHP8wODKNw/3EjvLl
uMYe2W1Jk/HMDqBW3I9xskq7je1Fr9OaAzjG0qe4y038l0zRjVUprouxMHrpUwntNxfB63mySWOc
Ej1biOd5wO8r/glUAjXe6b5GtHstX5PMqFjTlVaJj4mMJprLq6L7SuQi3iB+zgvMGF0wnAsRlaHO
Dz+xFYTEeUlLbyy5WYIN5rgL5eyHRcBCM36qhonWGaL5j4eDuSZkrLceLYGdbj5yZGIv87sueU3A
9ep3XOujcMw0sfkV9S48qdVR6+xGHBsMur6QZfMC1ZvGnzSVdp8i+1G/3vnSiFeAjRNTk40zA7z9
+nf2KHhUgFKOqm4MtsGoA1uEIFahKypnLUh1N6or1s6AU0hxDBqNgKUps9TE1Zza7/lD7LWh0nP6
XtmffkwcwAM9F8weiQdUABzmotiPOXF2vtF3wa4Rim65mqRWOtk1WzUIma1h9i0/0AAC3nku6egc
V8W9GMns3qiQFqBt882wPBuuoHCgQ8bcQ6ts03KrmWzhcuNeQsbaMwnd/sU5d1a7l91eAiY8bxuf
J4VPXq21LFJQ/tfMrbnXgd9w7v57Pr30qaOp/Sj3MhnibATUztHU0YpDM7fK1OBkvDAWXj6NMQYI
4Ku7zT2fsuBwrKi5/okGMOxrC4/J+uDcT1F0vwk9FClZ33lBCtJY7w20Z4g0Kxr9aRx7htmsKKhI
mMEYRCOJ1TeQZNgeGibNVmJbwq+zhmGgyxw8j7QuXfh6irXj7vPGafMdHH41PJLsCRthf4t1RiTR
Gczh84MVqzvv4/xsd8RsxIU/aHmqX0Haq6weEEKP7KDnJSVmVtQsBA6pF4OIuc2Yv7HaAvMzIgYI
isNlnU/iCqU4cbbxJ6z5zovlYPAWJ4PozKwI4Jq/ZDocE0my/vImn81fQnZyVNrrOTYZGF5bRjMC
9mlABLxlIl/3UkcAxIiM8e1dCCY37cMELiCH/S5uACQwAoHfJIIp15cYLOdSbe99p028u6jMsWBc
6RZ955gsrxyEV+XBFSoZyKKDFZ2o7mCKPJDxf0BMKTcV9MrCMAdVbGYglw6Lv5lM8bn537jui+uF
LxvaR0XUQHr8txK9iv05se19bzOGGAHD63JeOWH32cqxT8klGfvyHD+Fpiji6ts6nMs1V7adlOFV
QjviM39sv84kmEul+tQuZqiFd2Cb/COfoRmWKqW9O1Ksf0S1tdehpap3s1v7KpWEYnukcA6f/Q+c
YwFeDHvfwnZpcpTbeegASckygg1pLFN9xa59tzcErvG58HchUUQQkMIZYma4YsF3YN2bAxvGqBCZ
NuxKy/utttY3Gb+0VhJYFz6NyTeSlbjVbJfdan/289551kptKaW37GPkrDPhlkPKpaLqZ7hA68R3
Xaylhd9PkVlbabHyyS4hinBDNWA3TPL0B7xBSAezS8UqKNDNf3vplCkX9WrYBDKJ2ZY4SyhM5FYI
81KJjyGzzWY1HrxmuoelNyVlAjSpQOwWblWiShlC1yJALKkgIpUaB3OclQs5qHIHinVzwFrPWUNS
zzlr4AC8GDsKPeO/oBB9X4+Ln1VHikXz+whxppP+WP6lfeSuqFRNbhkaELmtwFxDFbBD0I3X3u3M
MCGy4UFltjclDXcuYEQExfNa6cd7jWvKtXJxtgBbt+WhHa/dE0voJpFa2PC03IgOxfptnjTjAx6w
qSECsUCzpIg6IdbmYPDJkQVk97bADjgiRC5dceQJbdFRljkm70psX/BBJtwsIpU9rVTKzGJDUkOx
kc3O09m8fZmcoCFpoev0aw3MV79VBBA/RPW1+AYj5grDW4cm9zfsaNY+2Yk+J+AqXd70dVaz7JlI
kFZW/CBEQ5jjZ+Is3/T3B8W0+sjPN6ODTlqGq6RY3u2ooeU44qmP/R5Af9kLusZ+UsG59EOXwSAO
b3OM+oe90KCf21POc2ikBxuYgPIvULYBNM4in3BC/TfwMquzBLbN+WxK2bTnYG2KdwX4q61JbZ0E
qT30Hl+z00EYRbvCENpWA5AvTx7bmovflIrJPfBXD/UvCnNf1pz3dT0BJmrwelExRs9hqvK/ZAak
dRtOuN+SeEQQ92qlMP2qSuSr2GYDhPCQrOdXvPAV0ziJaiggZl0AMTsl9gM5iymnn9KFYipLP1ta
/pqQsKiSjHqBWVIOa5PgkN1oYcAuPIs4lj5ZWt5z51VxC7eOGRGUu+IOdlzZNWXzHcfXbkNQj7WB
3OdCnY1oCszZHrASkJAUZxp2e/ZMIjcd2okYEc1srHSRvIIpilEdIgqUGXQw//PyICcSsaIf2CW7
P2/AGfDdmO5AdIe79HPuIr57QkW2IwoMZmH4nvqjV6rGLw8zdHNgMAsKZDQlX5DNRgOtLTQ4B/DC
qseX+amjY3OQoQFWrBc8jQ9yNzOYUuR5kt1S689r0tpJngY35qTjB+9GdhNgwjl3E7BCdkMtHGTn
8ziudKhwozMImLbuxc7Xp1F+JpyVobB+p4mGJOBVGpDtvq93AHBcmjGDgAAFu1tKnn5cXsD/xihE
ZQGC/7Ru4zVus5VKLw4QznCWHkFs0+TKloayPO7e0dEXJCjeOwYbfWJmsHmrU7MXG3A7oykYdWZb
PaLNNnhpmvc4Rfcq1WQ7+CmZ4d8hv3M9GUyQPwtptY8mGbqMFwtvsjpQGri9gx99YdcHrTD5hFIX
ESmv2e2nuHiSHbvfOYC7VL1ixeGW2gEEkkUkVJjUnpYnLtL/I1v0Ieg9c5J1Al64DzOs6AlaqRxt
F5N6FMYG6sTLwZXutl/JQ+c3Uassw6wsM6BhltHzUTqZyUV01fqfoWrFCqLqrEsVbNFNAG1r1/1u
sCUdzncqxVbC+g5DUTLteDkQIfjpEs8Y5qGNGCvQJBis7ZErGiAS3RMQ9wM0jYrtsPIKFIalnF+r
MbxdW+dPDJDB5xlI5eQ3Vzz6qfHAvRWcfK8xid98SPXNaE/Bm2x9uE6UGMqPlzTNc5Y6ILbfK1vI
oDhx2z0prLRRq/Dh+FE7Sa8GF2+BL0r776VmDHQ7aFwctIZp1pLBtjGlvouPaod8ycrcBTm/S5Ya
oM3PzTxeb+1VUtRWOTTIKGEYFtHzkk1jWFWjBuq0lsFS97+zc2z7hU+2FWBT8/id+mvhBtW5XX39
7DTCkPK6yJpiTp7daHsKZCLQFdkmSQhnxrSnnRgBGQfu99Yp7S4aIDPBwpz+QLiScXcjCuDo52ft
nsguvxEnYRxChAUEhDCGl9AkuVujFOAWwRJjN2SrvLzhPMhYSD9Szh2XpoFAA74rN7rNoBiGMme4
04B4aR/+sh8daghQ9KCd5H/T0f88WmREOPYz9LwK2JvAF8Ui8nSPqtb+UGwe4Jrikueuq6B+jYgO
lkgjuZ7OlZjm0sC+FBWQpXdQgT+QSFHg7KPebCZttTvT+PPpXPaRI0/Nmqu5YEQzfmF/2NgOD1p8
ZZL8vI3bR/jK7bd5Y494D6H12ut6H5omnWz3WXutW24BEKmxmPY5eND7tntlcDd9IlM2c+9+pGEy
SzB2+xHW39N9O80xr4JfraF6ffliy1cXTdmomfg0btPtxHX1LUCJmNya4uAY6Rhent1htxpwJu98
6biPGsk6h19RhlLLl1UNTV9iG7kt1lGjh+6oQK6l7KmKs5aPFS9r5eYEfE2kh/4HB8dAduUpm7U6
iLRDVgiSycHIh9dkMZmtrgssr8FnGfvazk8wAdfdkxhW0oTMhMeVn3YtDHn79SFtW8b1YpqYoVRr
srvGDmXuDuuxw2R3ImWAQaX3Sf00R5GtQrFO2Xfv98Xfaq93Er7Bc084saJ6bDUNfhQLXwh1M4wy
QeVOO/1Kz0vbXMJ1b5SRfJfTcYJ4pOUQiR+R0n6fMd4uE1ymgLiVh9Gtt2kCGiCOph3X3Yfc9uvE
FenN8yr8TCU21sBbfDef3qsyjhlf/EPap3IREnaT/1T9jOwzhAF1eETZp7tDYZ4hxXcttk7Vdq2G
WcU9sR42EbV96HuteUMBoiy5s8QWWXH0EVrpzrQGHleVk6GrXtoU+EIIuF0KGfO+HPXqK3il1L1K
DFHYkdGbHDE/V5NB/3SGwFRuAWZeMxk6Bm/EG9k3TvlV+wFAQjWGFnzNfguT7qjcOkK8q8Jn4mAg
aU/Kd8bBXJBC0tsFtoJrQTK9RF/Nl0Hb//puhcBXKN7sSgbKwCb6fjRBpSQfYzbvuj+rYIF1bNZy
FIFRQImfbizCJ4Q/1r//oilLPHr46ZC8J5Z6ecxlTZrSDxCZw/ILAi3cubDyHVVfpTcBkAMwmAgZ
u+eRwx9sUObC4Ebg3fc+7ThFQ+WMThCSX9tn9luj71GEJ7ddFuxDQNnbKySRznIqwn1dU02L3H9Z
K39ZKHcxWLlOmSoCFtsszcmXU+syTSh9BiFUNeR6bW8mldeJcQC1EwlmfGA3o+fwWLBxZCyFI7nV
pgMAwbAaIhXw5tY7N1NmZyva0UOSlzW/W8lnbfVJN/EepxueT1q9QN/XR6zYQkK8Y+PQEbxSBR/1
+8qd/s32a43GjGrvT08DExSYqmwrQdpwC5cWH0JuljL045JDB3fxgqD7NIZOvfRQtSlLYyFJwGa3
/CNBpIMENnuiFGFQXGG5+DCV8ReZO73Q4Nutglzh1FFxwyTFpHLBk1oeyhOlYNGP/aqwHkWFv9LA
2ReBtNklPCVru4doqg83nWghLH8tM1V3XffSMvkiKqHWZaL4OmlsRwi6Da0OQdIxVTmgcGHsEPvM
9Sf2W4t3DlcyN1/QGRxshxSP24gHksgEx93EohQIy+gsHKFeFC+Ys84iScWj2n+iw7zYALQ73H9t
e7gHMQs37ashh/KvbBwWBXP6N9JwOHmuuGVJoDJFNjB7PNGp08iXdNXSMhC95bFVHJ4/2CRaBtfW
ACcv8VkSzrokvU+rFylzjN9SaBpfB4IiMlYxqUBGg56EdsgMjdxnoYke6MVYZ2P8rJtNKzAl+4CO
VQ0F8rDUhqCM+vAQI3jDhDpFFbZt9nRwQAsGXE4y3n53JoOCLfZxVe8LSAzv9jAAuP4UjMFO1dUI
MdsyWGAGTZVaUmZA6ejyCj0t9s720LIFKLsNqQSG6tbCTUx/pF1dadKK7PLwRMiFCMLe5W4n297J
TGL+5N2SmXAK0tngbfz4vdYYlxjnsvxzW3mYWXVKZup/DlK7BhwqG9vX5PiAn5vlpXIXhcGCtwZn
ot6B/wkVYfTlLLdrfcVo5Isz004MzWYAaDu0cYBBP0HQw5mEP1Ab4evhr0bBoIrrQp3FnlbeURC0
wrZYhaZM5sdvPhK+pOeM8aeHsbk3RYteV2Hb9V9EtVohs+fnel46sUNhGmTJlFa247MlUUaohgRf
nMCLbHEHvrrSMfXUgXu3Uy7HBqJB8PLvhQeXS8YswvYjpBPW6+3J9DO+pxnEIoW99B1xL5aQf7+h
cweUWxkrFzWugQCQ/6ftd4hG4rqRhmiE4uJBgphnnGDVzff1KgiialMV2HCHRGUsh/BFEkVq6SS4
aMP8GbIGBv50LC9Fll6M8zhTBHM5yNFIuWh8q/V7GEg+p7g6WgQKozZpHiHWCh83OFPh148Ralrq
9IRC0DKUfCAk9e5ObH6SqH5uUGtWPDMzuspfxzr2MHTO8D/fxBpnS+sadTPbllORVjjkJyuNVmBA
bJLIjOMbPW0TV8a8UrVPV2oxG2O6Eqzv2vmSNxeiUKyvDC0HyNmKz5673Nqpda0/a0ZtnnxvkQRU
FnjeHvuYvmYGQgpQBICSuPTiCEO17aS5MpCIYoY3aQS2RO569oRw9mE2N1u77Xw4IHDpfRX3zpKl
toi05yvG0sf0dPYY1wiWFqxlFUbh3igbtPZRFlPWR+WAEV1uNd9jmBhcL2ZSJQY2C4u/qQLT+ueb
xtInv+4GqEBxoBdIjDjIPGA3VNKTR/4gmtYp2mPkmgBaQ7RSH+Lbtxpw2MiQT1/TUos/Wc/niCCm
fEtLj/0UMmdBEU/PETjhgR3PGQ5Q3b8ULy3KMRcGlmyMIyNG91c0Rr50s2hQVw+jiczNIsK0vWS+
UGW2/Viq0snYzZOHI3S9eJIU+oeEbV7SPvpjbQaIenxPEEoOXb03TlMdVe+JUi2hoIKte68R1/sf
ouJop2+PJspkj2LWW+lrCe2NdugLDWt4+Bc8ovHXfJWwnZ4sMjUiuWW9xwkh6mRPsVjRskLi/5w3
JVMxj/OrokjmgupZkfLO3QGDT0QQGnUQ+SNRv+eVrBxo3+Mg+iKY/gq5RcsBuwC/fOsrTbG5NXMZ
OViNtLG4kIT93v+ZNFMwV+GhMXFMmMIKxJNS/wcXbj9YNtnjmlwMlgAfjksCXigBjFTEs57UzF+u
ZIIAHe0myz5xQBLukQAzfTcWZh59gLugocFT6i3Tre4T+O0GqPGJmIZwOEXPODQGi+QlulG2j1mV
8/xAUbbCfCEISBun4sxeXx2ju5mZQkARu6rV4nFBUGhcbzPIu2GoIq+SxdsQbkyIddLNXJAoGj/Z
MeVodTZVuxfTGq5JXcUSoi+1EJjyN2aEL6POnW6i8H8Rg9y3U+fTCDhTMDF6QFcEyheNnw67BTjj
hbyxMR12y6YR56g8hQRWKI2uAhAiiRvEMZfgLKotQgrAJJiqoqIRZ3xYsXrmuqNGJzUyc0F/RI5+
c9u/MvykwDnwDVke06f2RuYSz3t3zAdMyfSsjXJLVOlt+1gl4AKyiu+1I65Y8XhMGSo3p+e/WIeJ
YlF3JOkI87vmAJcHUFfYdpkAawBlWNP5hV/EzUCYn5HWWSQuiEJaXdMiQtg9pc8ySeSKVME854SD
8ESl4fefvTPAF4zkmadyeWcN4FKG3zeSxztSzvQbGaZC7iE1owLo9vyRk+4uSBJq/QAekw66tcRL
Vx7zVzsXSnk1SKuaOWWk3m7hToNkiGZ6TMCXuJty/M1nbnGqcelUTkfYpwKPtUGsT0/lpnlTVjrq
HSlx8FM+cflHmd47IsgOnY3KjIzEPZa3wFn4eAcM3HcY+KvJ0UvtcbV0gW2nMI9gXtxO+ShWQiIA
N37LbIIilFyQLdmMrBroDicur7VCubipLfuoOGTF8Q3mUboWCnChytTTQCpfRcKs0qSGPQtcW4a4
dEhTsXbX/L2vyrcDyZ6sZlvKzR3kH7hioQSnvGCCwcWj+G06s173w4cTfIXGM1LoyuSxK2zR0WW7
ju/2ntoHLBKr7d0oFyH8IBwe401J+TH7EjMikaUXd++L6VjAwaT4xpupBQCgucFNvb5lhoOnSkmN
NHT6Lm7RMUS1CLfXPX9zrZFOL23++cD/pVLAwifK6+qDC3+R9MdGnE/hznaOHpd/Ru2kZR4l0lYR
/hEKTivQEC5QfwPU/W83xaKRV6/kl5QyPWgBshHwThjKXW3/oeUpJcR1GDStYbjqdSDlRZJG4FxY
MBjEad+R+6RaibGZzeVB57R99hvfX1hGim0/pBCwL0lyWH6+DZs7FXHDXZxYWp3PDR6p9eKofvfc
vBm5tM8xZGhIlQEwoM0MSHyOj4UyeUOLm3W6DEU77i+JBhgNbmDqX2AjmEAl2ASgyo5GJdL4H4wk
4+WJpmrjYreQZBEAN4ZZg1yrWx7n40Gt/M4LgJKIkPwsh8qFZ8060oFOKZ0hINZq8E0MksJPRDzf
WCTytYvlZ97pd6Be0NVUvq0ly8t7bNU/Jc8PakwjkDTbY2Ktk+oKDmg9NVEpsyZrNR7P1I1Hq1tQ
L85Zb86cotuXoXudNuq0BWDgkps8VQkjA6+QIK6cuofnfCV5RxV7x0pMhpZjr0MhXAUPaSQueKS9
sXoK4yU2cXA3oAMj5KdF3PCwkXjD0pk4D4u78+DZtG/pApyneC8JiTKBSNFYdJT+ea2DtDq3e35R
NKvmdH5Owd5NsP98WsS1poV7DSR4elNihlEqxxDppr+mbjT4W9OIRjI9+SsZXyMVO5NDJRIKF5Tl
oJyX2Qd/9o2DcHRMWEcekj1QHbmeFEOgv0Oyk3lZqna/M4nVf7qhsSLF+W5Z6EXdYKxSSRu3JEqa
Q34PXsuqwgliNV5i6V789L6Y1lCx9thjt6Y7UOwpGBiHsNCngO1A+rKNalrOHftdj3qyh5BhIxGD
e0kPca9fn/rcFSdBTUuKIXgTOXM7SyMvCSUppKrDd75KrVYWWRCKvWJWvwEPQp8ySI7TmljD4MOQ
PdeGuGkJWfafjXZSwISxY3dIxcLZRu1oBLZC0X+WSVdP16Bd+xLvRvQIy1GczvZbFCMOx+0zmTBE
aiClVDGl1sWJukGDO6xchUPZi9sC4twFi97Pa1GLI3gKF+xkf/6KsHaxiH7493GfBHXC+PDiyHX8
5VCmGwAi8JK3jG5PjpMFKuu0OdxehICdAQsAqrCr1+exzMALqoiF3b5mqNCf3zBQZXM5qFwy6KhR
HYZN6KBYFUbUiypiTfgzbnqVgIAA32vgloFqY1wTWucNMm46TzVbyOK8mtJTyhFl4REJ/27lhtyW
hwO5zKrAA7me0ieIkL7lQf8sanqVq6rvLFwTfs8+U7VYVs5kc0hoy4xI+IS2TXQx6MgTL/N7a33B
OWJNmni4JscLfCUVla3ZPchiUoVk3hpiPHx9G6rsOI+gT3aLZFacS1mvQnxIYxbXKgYzfNyZ0Ko5
eFZ4o6AKQbiXLqxxoZ1butPS8+A4BibUq+3CbzyeH+E2sG0Jl4YG2o6saSBYZ2VHJTw1CawuHoMJ
SYWP3DKnWXrFeuO671vzDA0IA48nxq0kZRbi5b8qH6AezVOQWStnZVK0ZMaLtdOGtTCY2xudNtZa
kdq9l6aw39QVUzjHWM3GOpcV33xFC5PsNsDd9+ipAWX4JbQX/E8uXMxOaJxUPVZMsCjUsvvgsjHg
8o2OI5acNinFaY1Q/TfXumDrpkUI1HhHZwu3TSZCBYGpryQLMGajILWM+WVJUQzmkZQOpq5KLLTk
JbdX1M/56Ekweiw2wVg0MZwc4y++8B5MxHSPsG3cEJm3vuT0uF0F5vWDVGmlaQIBkEP2Gx23Ayuk
YtnHAaEoErk5QcWVXew0MV4iSuvCJyiAMk4hhScRdAW4AJyPmbOU6bgtiWiCf734JTu2y4SUeuvS
hNymZpFThN6T81laLKRvH8vNEwEwPsKHG2rwD4XuUCKgmyNK9HLsXTyutfItU7o4GxWCv4jlaqJv
hccwb2oJ8BHMsmyIQJvhh7JzXXPjDRcREVPxAybQSKP4eBoFJrmLyaL1Ckv9APgwk4kIfS9pP8ia
JyfL58xxQ/SA5JLh7f80OAlfJJM4tUX6ONWcvY7AZpOxkhDXANFFR7ZXwWijMHtHVdhE7Y60rTKu
GnyCUOhHPeU+twdLN/XjCm/huOMhqZ/s8Nyj15OY9DodKHM5KKHgwCa+kXzmLXp6QpYxrjAEMk3N
OtTlvvDeIsB1Wwmh7wGw82uCaRAVHyMoyjGP3Yxjgzat3BK3qQPdyk4ajrh59xV1cKvpP793z9MH
cx4DzYf5b04dMgguC3ANSmBcQN8fCwTM5+CFVMiPbcPApbkoJKyO5Yd2vhzmBmnUe0D9qNKQ/jS1
j2/G9H1O/Unm1prmFewXOt6WAFgNSKVFKnidF5qav5h+HlrMsnMx9MMk7gEnhNWawtm0hKvN+IgT
LtRyadqsCDTKTrNcrmYp033gsm82b+PKPU1HrG0+MB/MlY9DzDi2VE1PTLKTQSMfdJsHt2K154AV
cv0///1X13YWtUv9XXtFFftgtpaV6+CeUu/ybZS/SirMrkG60hpaOwF6mejgtaTEUAnRPM4AJRd2
M+QOm94Kx90qOlBSJFHgQj+FSNuh457O9UeJlvKXikFR13+fgzpUiMq3SCza/sC1xfi7vzhGdJAQ
kkHF+AeJ6x1qj2ew7apJwMkAbBoyjJXkq+0L7QHcq9r4ylGyx/+bwUAiF9FSfGHp0PE0mb8yCUuk
Cd2AtfSYktk9LVJZTEb/m1CHHLGeLejvOf2wp8nqb2O7HN5Z976Heu4zPyWtR8kWjl3A54We2mUT
yaR3BEYf8XUJDCNsBtB2G9VNrawyc+pu0vr3yKUwl8V7xkoKcS0yblg0KjActcDFwwQdCJaXin11
HDbj2xR7xgCux8JHjzePfAe/Y2APmSdtyQIRxy0oTkhhllw6KyWxBpcnZFXioUA7PKpwDZ8vwjR9
yTiwiY+ZvQvtvn73yeF4YrdareuK4z/EU2V/7r+CDnBVw26SGrcZ+maoEGDrD0SBZ88kVtj1AZWy
3Q7PLkxbfCXJsfrsDHxhr7oMNVLapqgN0FDnnusJp9e7clnPuOJu8YUENczbzwVAZHvZH6V2mNXD
eBs0j7/q5PDMArF/pt9fy9lO89A1731EBCORIC0DnrOHUdJ3PF+4X1aPaO46lEzybkrXBVPn3Vlt
F5Ydsx4xFOSytzdbztERe7KEqJs2DcTJ77pXK0HWWfKnnrJHCa1uUaJTEy3b7FtwVm0F7SaeP0rR
6lz/UJ6b1aSJEurG3UyebLq3vr/cki8S2CY7WGKIwIa48G9pSzRzkjhkLyIYcvJugUM1dX4PME/z
qam6639v+B9uf2QSK0MLTJNPcVz+wZWcibaYM0aPAzNVXrHMst0aeaej7+2EhjTq9rf8R/Z/sxl8
HbBrnBXwQVJg1Jb34hxZEKTbxJIH/HQFFX62DxgrFQLtFEmlOxcue3pLFpLB/P4OzkFZ1yb/gQO+
e1/TQrKPKOyGU11B0MNxDj3OlBLUujBiRi33vmOhGl9DceCKKOntiNASanwpaTld6bkk9BpdcBXD
dYdr2zRCJ2/TEFwEuvu7p3bDENu2FyeewRVMyEUY6Dr6wojxYGl2EYQjXXk2O56K76a3iAtE93NG
5nIMe+Ps+eDpmyAEe1R7dsrAheYL3/qKNht8C4XsG6nChQaUYMIUZmDmJtqM61ntAhD6Izou5ngb
QzmNrLhIioVyyAMvWKBUplWiBYfCG4NEPO82PgTcN4In7l0cYFPLTWOoEehS/UeS9KaIE0VTOyR3
RTK2VHg2PKo8y/NKbu5LzIUrwAIYIZtSt9s3S4DE83mFGcXIOSuiGJyohaUKsXzxpv3y5+oXxGiR
TgepTG1ctahKGmA3UeMctlW9Gh0GWMlyJWeFUfJXc8vK+KRFv72xJLX7m7fr4xraMhQyW5FDVXAt
U/lprIi1cXCveiDfQmHkYQyOEzkXAdLm9r5erceD7SidWCke8QQqkQG9KhDZvJQpqGF6iZEaSwbS
ntHicwpA0pGwnHQ9SOpgdyXWFmv0AuUajjeD20dDO9uogBqJkEQPe1CiXCOnW0/zUXTnIW4DRNXY
C3wY3ctPAW8KngNLNinx8MvJPbDbfdv1cDrQ6IK/NdpTHgBLofVljNMc00Wz6qjP2XFyWeDKBGJ5
tZy1yyPOu2UtwSJh+vbt2By3HkQnV9onwdz0Np/FlGJ4MfroGjTLId2wcbdKjiJEl8X9jF+P2ZTt
jOKLCASAPtJnDGKuSupKhdUaSnEOtD2d6MF7YFanrCIl9fSd3j2CEulTjRJO5TWyeo8Ou8Ru3lf+
4Gwzpj7GFg2DSvanrSPLxZ2nq08gWBJMcvlYQWc2Dr/9THE/PHUg8pdVDjNc0d1ov2jY0gKhZLIz
ootchNRzoIE/Md70Y/2CecGX7zxzwsBQ45Qpz82+AcU//x77n44wct8JmgPvBqN4iXgLCpq2+pxv
EcUhp7lUfwbSbK5BilGZ+i8JY57hYo6dbLnrG92St++8daQ+Ra15EHi8zYe+flQUwFyDosMYjlP+
j1KFHU441o1i5ZU3pVExZmkXPgJKr+e5/GfnoPc2H70n4PK4smFtDvCJzKD/Om1gy26hYiisHGiG
xv9Y9l63fTx6VVhgQRfGHbaLnBChwDWzdZXx2owXwJ1128J8yUyeV+/qEYkDDJFQCmwLQp4w3UBG
Z5fKIPZBy9gLfrNpMUE57fbXcIDS46+L6FmKVzL0qT78f/hZU/u9INC2gl4axbtb3jYQH1vI1nIg
Hpu8vUyy4UCtfZFs0ZU/UNHsK7oILeBNhHErosWOYkGGT1VcidkN19FMCgscmqRE4ypg8KVBi296
wAs6wVw2fDRnY5uHy7rDifTs1FTQ3XHsf7uZyh2Ib9shTMdbdxWHaH41bBMQE4v3z/JVwIK95dMK
6aBw8+lHgURl/3C4MTCOQoB0vYrXbfWdfSiIgJ9UVJDovzQPNjzyp4H2rRa8Lobr0Xs9S7YFbImk
FcH30o/bP+WmEOra1bdB8uNSWHHJmYbOLC7wgU+40A4cLxftI+9VJH4ATs6bLHZNmsHg+bmaUObO
5hLSqxTDiQsMzPqNUDN5tnQeHnPWB2OE0e3MT/FU0jQjdfADsQAS8WxqK8usADk4n48qtq9Q4xXK
I1M+KQz/s/JaK2bx2SAf1VK2WdVe96InziAY+SnDqz+2GxeoTGg9IQqi/8Ts5Tm0zG6UDf8hkN1A
5dMQHKzzUgsELY1gV3Zli/HQ8h1nelHiHOHfVkik4nXlS0aqE+qbyalaJ9KCYU1apB8k1zFPJkme
iz32uwazHLhlT+rx6cpIrJnj4pNrG77pje7IsvUwhh8PuuWQ/QI+EIvfELMWUXGoDuSL5GgOl0F3
s2LvyuD+2HfIl6V1pzI8ACQv5FhadwuC7Cpoj+st0u2g17Z17l5/agJFqvwsRplesatWGYGYzqx/
QR6lMxGL11FL0f3RFOcn4PgrZgnjb3NMP9gEa0Ezo9bueQs0P3oJljX12TeORERBF2rD/1kaXGCL
85qFNZzWExIz4jObAp/UUa8kppiSfgyNQB3SKVd+q3KGwpMC2S6nnzmErGhMgWD/5OCCzhCB60sL
MPh3KgCntdMtEKBvAvimiO2gBQw0gKDYdur2oYpeBMKfpQ4skS0UwlLxfP6o17xi1oPwsnVltiWw
VCFt1xtLmozG/A8s+4DYamGetMOSl/Ap04lTWFJHZjBM0jmHWTB/qakG87ff31IpbFST7ZpBTi12
HzWj8Ck4myOjIel8YvnOVLVl6647t++ysqLfqQT9NSaLTbMVKL451ADEqB5Gq6cagQKfG0+IM8yI
jDEFYiPburdx5wi30wZQtUOu2kqq/ssEI+0Zln6ZqwDw7HKxRRBG+NXrmCzB2y0pLkd6OEbcHlAq
4+ZCm6FAr8cJ8Ccas7VGBxzzWqWkFh1s33h9nxD18pkemCGZOzmdom0O8wF28qlV/v0sxIjc0ILN
a24lUwPzaN/+LLe31H5sUKuXK6WhdyaRoCraRIOobmPVASFeG3uZtfZvmD+qCmdhTRIEOwwyyOtK
7P2AtX/uytMUTWvIcIHovZmTi8gH9OBlPnKSCUYSi2XKN2ir4LHcl3cMcjUhTpevr461Eqk8vFoB
C8FX3xw1/pTRmnBH4jf/K1o1gouDEbJCwo9CVcXXGtlB7ZRny3q3iD9z9JPWILFZPoH13CGEf2hO
I2mtGvJKGWd3Q8h06YCnY9F6zdjVj7tOyU+1Mc7qld/OM9/vZpkagLY3dkk9tK5GFo2VvbG8d+S2
R+NUoi1b7Po4R6RVBq+jgK0LNpdFAtjtYSAziNZo7vaTQ9yqqxicP8Fz3tFQ00I9ou8Ud9UIduA0
tWTjeioKN/iYczIwwKhhOZ6h2vpiBhG39GSi5ciHlKCmkczldT0qcSRZpdo6zw5WG5uI+vM/lX9f
NKksTWkWAxurSQQrc0WnOM0NdKJ9rNI2wXkJTJ8iZP1GgDuuXYeFbgkmQtYZj9IOKq3uxHxDkgfM
9xqANLWh4uzXh8EBatrzg5UKRDzsh9RyDju2XibycYn7HgJQMT9VRHywG5x9UuPtDOvHHoJ5uEfg
vnO4TAp1c+neesMb7hMmZlW2ulTLn1y3zpbbTmZJ0fTUr5HVJgZROEiACVNC0PEuQ4gIa3dNyYLw
HeuL86DfiFRVxJnJowD95eI5NLVJF7kGlR+Py4Er5PBlrQPasoryy7u51VbOY8DCsbX5LXKzUs0c
9tnGE0yM5d7r/snnAd41oOi2Uxw0dVPtFtyLXrVG6sfUJZqxVMNZqISRFl467jjiDSHz4siWf8WS
e5mwDbyD9ziYe9VIPkUbtcOPb3gybzG2OgdJ3xswzCKXUEm6EGGqjKnlF1uh7PKqQn/1PYxT6zOZ
P95ZQ+PEnfvMUJgPw4bugJSrx24XrF8KXOU11PlPRvRO0ehkEOPzhDrbrI4iQd2eOMo4q7fUqOy0
874Ky7+O8m2CFJoBLSvyTq3631JyepSzaHtz39TBU4LKmT8TRy3z2BvCGrid9ZGO9aDOfghfn8Ns
dtGhc6nLHw4t3NB78UbaaNox5z6SbTRywG3lllnlJg1fJvYeRyQmMCLCd8vb634gK6yRK46V4MB4
9ywiI9fLxCfSAh7n799zifPSZ4CKbnHqWaolgz6V4iXnsCq7mwadJznF6FjKQSOtWn/h67UhaEax
JzZu92KRORmQ1N9YpIjKvCV+6AoNNsdQhffyhYYVw5QNoDemxgneYr5B4HbVEvNzT9as8funHGcJ
LeJrYYdFfzoE8QfN5aqUdFwlRscyznKTXvImrF2X4Inpe1jSeFJxLiTWobtwUU3StNb4Pm9k6l/g
SxlxyKwu+0YMbyWIDbHAxNm8v5trrbOx6WEtIlMruC20TAb1bnk4V66eYM8tv/2RYZ0iekWbJbpi
66IkE1s/XIN8e6wBXnKvHg6mlMdFUXCrnLkCyXAMSqiPc/fHHulLlzA082MnYchDMN3ERh3RzhT8
eQHFRUesJ5ma8KFJGlSMb/aOJtZPkwm2lHM+qqaTsIJrTihNEALtEj5NjxKdB6B7SRh7Uw32mqsh
1X9c+6JpGtJIXtQE97iAAzz0iCeD6sIW3d9Itu+uaCzyUzS+qWGyG+2PsgP05v2LtLDaPQyHOWxc
ASjOmmbEc6Fb/gBlQ4lEEZvoyN3DPWcHgAQDnRJm5vKQYObGi31UwHIuK7Hvz6eyNzmU3Yay5jJh
AYbWPTJiJgNM1caGSGlDKNnxoY7LKW5Y0RDfka/SO3CSGIQLaaQFWTVW5+XiEQXi0+qpggio3GEH
H+DeeE2sbq97BXvEuKI9V8AuFaJpVUS/yDjeKZS99pPXfjhUgg1AwDtCVjrMNizgNjpho6jsDZAM
zjVmQsSBf0fUym1shEiIM8EDtTJ5XH+DZknJ6oR/vjwZVgXvuMCT+fTD5aGvPbXUnik5f/mHg/yL
M4QtHpDU6GwkqZOnOCXybI8A2tMgFk/b37onzG2zzism8Nrrgt8+D926CuVmOnFjy6ohQbImJNPs
Qt3sRKS5eMUmQri5s3Orjh4iK1UeTVrI1UtLB5H3KT1lbbXuwSMYxVSHtrWhLRYzgyiX4bOnTEiZ
H4GrADbrtQKwVWZ10lytdGWNy/koFcmCXVp5ew726lgLgxJ9xHJB+0+FdgIRlT02ayBslS8EsD3I
kVgLEkISetgkuas5GxQ7tbFO54UoI5w9So1YPUHR5ozQpyIMkCVe/K/hc8RdERCALIsjpGpd6L6J
BUrry9FAc4LQJIEGCNJI04/+Fh7z2kAnLJWYbBUQ8ojeok9LHawgyeNS7W5PBNWTnAU24KbApikJ
fOZcfoeYudSba0HSdmbHLyKj25vpv1rZj5OKyjpC2H6v/j4gKo2dDpGbXOM826pS/DydnaIamIve
tQQ5nnoVVLAU9nxweLUtlsJvxsHNKAb/79Gd44HfEU9xu4VIjcxATpvjtLxInTNFeP327LRfIe0u
Sfd1WnWlwNJhJUahYKGQC4H7MyrYgYbcC6TBOcLwK6JY22r0U9wiaUMK4s8B0aKuOuAwjKzo25BF
GC4nDE4i2ltjOYtz0uVmeMgrsHuGUKjB4ZnMfvjcKscbG0oqSPtFhc3BQWlh8g8X65BAJ/dRokfY
lN0Iq9fq/50gdiGOcUYEHGQNaitNYK5yyudDHbzNiqKf48XVKxbZ3B2CNlhJXD1ocDuEam9Q76Tg
R7wsbCBPLLH2/NREMbWEu5cdpyxryGj80p1vmXRB2tSH7PKYq1O7gMGt8wKcHNtXEVYQSdnyDIR8
EdrzRnB06b/xPfmzwCRcxCeX1FpcAG/Nhd4Lici7lVR00X80nzjxLHxq6GfNEw04s/G+fMa9GK3r
U/DkBwTgNjLIs3FssTcvO4ymaECTrRpG5bks5cA8CWj89/9NzsQayviyv68LUuVB7pRbQBKFnQoR
nkMGB/rGMTERWnAJiNObbfihk54FctDWUscdeJe6qI8fJX6cCCehQAM6A5sjUvEyv/bTOnRhRVYC
uboy1P+rfDGlncuVaD/z5SEErwMvSXtJ6jGN7DsUGqMf3Qh+8pnqhiXpkNjI1dHKkelqWdzlQ5Wd
T7+1Rv681wJbR5nZAshQ/V0rkMMQqF4aOt2YYEJRzlloD9sAIAUo9+Hdjm3zeYVTr7e3yhxLfrmK
q4Fg7kf4tOyRSEeXX8ALwd7z1HaboeasRs10TAIKoSKVkaIb1ihiBs0pdTolguQdLo+UREGLdZgG
+zGeCE4W+ZU8T7CUJibNZm2raTck9+mb5IwQi1NQkN6C9hu/yXKeruHwBiyyc8exjYLe8ut6PbTn
qM/7kpid0CxhLhsxDj0wzr4ztsyOdC6ut56jWugHQcS3H/fcBYzCYawA4P6XxpajeofbTGnLQ2Gq
0/pA64iIj5zXBYYK0g5VP48ZvJIQq0jlOh2ibKCgau8QfIBUTJ48r7f3dDpS1e2QGL24NfpZW9+J
enCguIGiW7KacgKEtQk2d7JVYRXzPvKZnHtM1T6GT8UUbrDPYOCYOLp+/Ms5LQWI+e4wC78NiW6O
OUHShEVwysU6inxFPmIf+VbQlczZeNoRbC7JEsiXb8lUE5KNesPfu/AFuui0ZW3P8UmIavI6filT
KMdPSl5iQ6m3HkHgPkDol/l6rnSgcKKLtdMb63B8pw7diYEN6487/LyS4UJkpPTmzSKpFVfYi0it
DUxiBMEPbAeTke1E0XAtGrFBI85BEG6e/Ze0GiZMCB3jmGBNmAY1r/TGNYd1Ja06n22GNXjsuA/c
lIiNfrqSbSCr02cgQ3y724GA+PVWTDmOqX+UExapcT//023e+QZiKrHVDJWjWrQiUo5fFQsWqcZY
E6LpR9n6NMWjfySLpE/dJMsO4BVoUUzPt5iLpdYk1Z/7VekNHkerECGmLB833gmp8uCt3QgQDho1
PJsM7YfX+jMc0HPyn8VU7ZwlfNujLHmDjnCCdoNan+Ok7+PfnetQP0RCPrbhxw0tddxVY32/aLG1
Sfm3XqWL5KLEap1jbK+aq1GwSLYj6pu7FaAbHQDrItBbC83weTOD1XRmRaddpNCutoOJ0UGdQA4F
jwy2QjCYdZWGnqzZfC8FYHuaPU9DNmJqZJkRMEKKO84HP/yn4QGsb28PTTJ3/VbWNzXmVIQ29sI+
pl1zGn+LMPudtQ44M/BdrIOiqP3kN6sKA24S2iUajYqz0/FWbwhTZq4qyUpGGuSMHyBHjInYVHb4
UKL9HRTdXT7/sbUXWDxFeq4wIB25Mc3O2a6xd0X74Fp+XkTi7WRpXZCoGKMGkEHbAmQSgQXuM2an
YiUvQ4TTz/e0yd6aRKMxfM/x8dIzWbs3GTN7vzOi+Jzq8AmDijUIM/AYO05sNAEC6kWi04NGGeSo
WdHS8GQXhi5N0BtR3P4vnKcrr6/jTqzFbLBKfjunxvdkl+z8t+UvMpnuw0x8+Ld4G86AEXStcruw
aXWr0Pjsnp8iRjQjLXjPXhqqRBO2vcI3Xm4QG1bJJ6XuIhC32RXW8pTSpvGBBMxJ1MiphYldKYum
8Mw0kcuBiO1jSweO21J3ybYRonaQadd0/IxX+AVbvoT/+K6AAuYFVWtrBcSVZlnmrRn4r26WWlon
7yi0qaQDRaggh0+IHVjBiZoKXXBP8R8g7nfzoMPx6h1VyBRu9GmHuhZ3DvYFe/2mzg1xjweoK0Ia
ttR+dFgTW5ay++AiI2XrFQUV38wDTGVYE68okuj6Ce+cCfdAxBH/Q0mhEim+9h63S9brsb5c5Cif
zAHw4CdabQGqWYgOp0vuH5lLpqlicm8GFPe2U4+UFKOhAJQFUn1oGkC2CXRpCiW5eJX0AX3jc6uH
1bU2RMmhSZokb9bSmRrExlXeAjhcz7ou9854zm3PJaOSQDCteQz8/1yUsCJPTe9ot51F9GyK7KEG
I4D16isSwFuAp/4fpP+KYFUHCyQX3NVICp5lP3j9+NGXWV8p2G0CuQCvzCwZ3E7aaHVritr7gGiA
NzoJSEnucux167Lz42H24Vj9InFiYwDo5Zgt4vLZaC9btdBOY4dt5bsK0BFPr181eoi56fZGGMlR
iFBkhGOQZa3AbhAf7OUYveuSl1bCRVj675+XPtFcYRL1abQwDaPJf0DFas5WuLvm3fiOaF7G9WDR
HYZ2nzwRfVcrHGvgJHOlSX4g+eDpmbOUkQveiEGtP9+ogMg2CYRG1+WxhJDZRLeGiJv0/lONireJ
aA6o9DvgqEEor/iq7O/gH0HTHvmkqipWpJCAwMoX2oACwXFoR4jtXh4Q6wo2FQpa4hU44KiR67Kg
odd3LpSLg3g6ML3+TNeAfewRQtVCHAJBjnQoGK+ZdDtguLj4bb6AffjrZL/wL7Hk4KT8Gi7OPG+j
/ebPNAEdoToNUvFfzQry6sdBArQcXbwFQdv3zyOFvjp0nuD86BGtsFllZv/k/T81jT/IdmZgnTks
1+lUQoBMj4hAqPB8PrEDphjXCXRt3m7uyO+VeuyVIQH7H6cUi1eerJ+h7JWGh8bEeXjDvxWNHpMM
UCRe/hMeybgWQhhlUwuQUhzV94OBj+ZyOuEt+AUHSpu/55xVoaGnXD63yQfP4FV3W4Z3UCvYMhyG
WDsIaB6/KEdxxVjLJfu0HXqombAvBp+kHAibKSGb6tMkghVdyYzCbXmSsg0xnBbWnSe0QLF27AZd
wP9oMmc6DWkWnoDYt6STBdTTWLrQWFVn2CXbSeRpkYQiLrWhZxTrdOqOJizjThwMYSZD6TB4uoOd
j6RGsZLNI651n9HquC1sAnqGnkPSsA/Rl2GihqVHJLPaNUb/ADhK7NqgKGnBdkwP4nGQfjZvsF/2
4prDLj6/xt20Ov08W6Wt8PHqLV3x3qqmsFwSM2pEZZZUu1xtw3i64mVji1OGacfXqk5ePdnbAiD1
GxXlXlRMCxYMm7PJ3Xdouo/sn2mQ9S50liN8PgYz5tI51Hi8V46fhnLHWIT9mekVbVJ9dgw3b684
hLwUz3HFTQ25O13Ol0FdLOVfFx021roXM2fs2zRswBaqHU5Zh1FGRAQS+1GpFwSp94++YETgbIVF
XneFbMcNQAC00muma2AifzgcXxVaWvrXfo9ONWuHIv89RkCklXrlDY0MPHzazBKUZLLysqvh2Sjk
fObm4hFmxGGBeOqbYiBXIQoTxtn9n/LgbvfakuxNEkymAckGLY1OdXsp1b7F/I7qTIwJYwzw6RY4
j8z5nnZwnhkHaMS8fWuiKwFbtHj3kAjByGVsdsSmHS1AGGm5bDcHyUufbz1HgJFMLF+4FBK7RxQX
LfiuvAwuN5uijLP5U4AQKbLnq4cPotuNn8+bpVWtbx3p9yuMXpMNEuVuVy4vv4TgZAfDTpeqd8W0
b04vfUGBmGWnmXIKM0kMO0ESORzRgJf3ZjZ14CFmik2GL8s0T0E/Qo2H/6mvxXSF6dpcUijnzSpg
qpL/oo90YlS544VL0W0VVbR50ldORHglV1nFpJ3nlWWYedae3NPanwpG5TmKmxtJVwUFBptKa/ol
fpzbOcMyTzvCcZovjqZhLaCFtEPp42MuQg/ip6+0dMaiEP0Mj7ApgicNkQ+2P/RUlSjWZARcGB0X
FOQUuFeVI8PKWtt3tey9Aa8+FqkpWHLxtXO4yGIDOiJYzbRCmyyxJiPIsz5KVnP3ItmeyvOxNEOY
WVFIZCx+DgAmEOQQfCx2nWAeUn8Bi/Gyzk2wEVH+lqhbGWa6Zjg86IPEVDgfJgO5Zf4mei6tr+9F
UN9Sw9tQvIWBXP6qAIVysj8R7bYVGAStOkSvZqe0L9IANTa55zU/7XbGJidKQhnVSLk/LnMRcwkY
VaQFbzhL0VzvqP1YgeROEfbPuU3t3ml6J0uLZ5JgPzMeUTLLmeXuWRuHsbpB949fVru1Vuqi3k02
Savri/QI+dkgxMB4paWQgIl2q493G+agOLkvsqQk3VZjJmeiSkSlcPENUoptMfjivXhKLHjZqrTT
es9eZtAo5/txfES8hQmv56IcuuG+3igxv7yI/Xs9vUHkoHx5EAl0bML+hTeNqRWFLOhdUlZ0mkHs
vSWl2ye6IgOXclUr7WvCU/NBRkuKcx6XpQfLtODsS7Bqi+4xgqwJqecuVHKh+QINIvkRMREpjMgj
cX+rec6gQ6POCUBJD93996mQCZKvteidhtNbtS85KXfy8wB8YIdKheKzp0BKWYos6gRKn0qreOW7
NLgbnRTyWpJ0fvwYOXss/8QbMz8HA6ZJyICEjBAQhHlSJU0Q6wPsyPCc/ztwYm5WHyg8dO3wV5ks
8NVYMpD5tq6CNhAYuGVwG/Nnj4Sg2BrNf2ZlZZ9uJ6t2TwDo6H3+xsRzRHYhTEYXlz3AWPa6T37I
5cmRLAepmWq2AV8oGpE6nG8Ot0a834qOH8bee4HyFuqRumHHuPYw+M3G8mN6PThtOQYswcOiPs8z
ZhIm3dJkAfEySKFdl2S3shBG1+jUp1ddX3+IXUc2StSEUJH4x3q6Tcg+6drMhFrwzVjjZKK8jRNz
BwqpjPFAHmsL4P8jrFjZPQrEJua5gTXm51OH6arqV/HXICFfF8KMHwBLOq6ct1wk5bQ/qQ/i4ROZ
4jsfNcZ6QKNQjG5kZL7X4RvuE6GHizP38hAfqpxOMDvWi7lJt/mAwOY5xSyaVKlu4fhwsOEmnKCt
8YHPnTp/vtioHWam6dDSoXSeR/TCCsKXOxCdp7Crki/vqD2sh/BPm4xlHLhvxbZAWbnptetXcALn
ZNJ+bWr3NkeF3ogVSMLnZEXuybxGjLSqRin1aBEmUoaezpzoAR4xrhP9xQASMBCBFNTNjanO5kdb
QZd7X0nHqB+gvdsOmT+nbhzeeQvpLZqW5zi8vPvVUlUdQYyy3UT5h2K0V0kEU2l5p+TV2H57sU+D
DJLeLxAY/qMyWIBKQiZ2/vwSO9iOypNjdz8hTt2ZQspoXcjkA/U7c6CaItuMsrDuIO0lSbEUUcQ2
ywl0mr9/HF6iHZdb9aiBWQm0jXXbthFYko1p71SDAufnFktlLNsin4j39EI9ZwuqouNABB4hZHzv
IwXKtarm/AgrRfcfNN3+9xlA6QXkcQTk/QQ22CsUTZ7Gjb8mXdUDFJTGVefJ4LBpza5aarDIw0kK
QIhfLxOzQNDVkVu8eJegt9V4mlt71f4Fd1TVAKuiMzg1VOXNm0bDoGXFnF775yf2+wQd8V+nuIO7
/y0wOiHfEU+lqYoCoKtsJg7Zym/mLRDCmYK0Srcant2rrWjzry6ikpUsnWPUBqAsDi7i0MjK1K8m
Oa6XvSFBEF0toLb6/F4FctYHDnRkX4nTIJxqzXr40idlhDp6iXYTQlJ03YB/PIeUfNRKBhQPwlhS
8n3ABhpPDizBU8r5fxNOxde/jXgfjAiCHMQp3+5qC/nz7V2I8xjpJv11tVTQQzH2Oevbjl04GLzx
BVQ0bueUl07mAcAXOUKqi+ypFozcPj+sPugryEgsQ2HXnJ81VrBr/D6SngxdIw4z0Y1EvFP5jtst
8dHw5kHGqQX7kxgx/GpKoMlXOdwR5m6JVIr/tJgZ7Xk/1cJ0hFmBTBtgxJFeyO7c1erlxYWgYy/t
Gy76OGs+MUhh5Rq7rZkYYbYgXIqZgIe+Y/EElaFc+LxjdA0JLm2a24SojMt7ZkpeF0YuhVM3w1R3
IXUIqzY9vCwh+YcUMa37fFVPmN3IipXIN3a7hF9Gmq0QVD3rPaIjwcIlLXjh+4d8tOB/BPBePACl
tVO3n9sAus8/XG3ytvn3DuRlt3EfhLedv9bMvbmZ6qe5MtzzB6Xl7z8MzEg4wz0E/HkpOlJ6SccK
oSx/05Q4U99p57w/PLjDK8XXizkrcmshDjc9PAkmns8ciqCbUkE+KtosSeuq0VLhu2BsKE4timyn
CuKTviZtgMHWnhJ1/IUq+NgkMh2uc0KiA9vnSHKIcsNbICLsV+91QgoK4yk3auaw0fFPZS2gsAJo
ioNgSzZGsp+5FT2Gzf+8mhqwkiEVBhOAh6Dxy/fzKcHp17otG97e0dYMyQdDhNSUZnrQo+vFsUb3
6OR//CzcZ2cg/luGhpRSfJsllp+WzT/XG+WAuIV34cWFFxGy/bgi0Ra9oOVkl4yIEm8guz3w4T2z
zKxdj7srWz8yGfmY7x0V+T80BVMkCxFS1TkqzfZJbQBQU4NnjMzr8oAcOYhnWv+hHzbBBFjPxyMY
jwbkTKW7cCV9nUwRIQpDUjrfp5Q14txwS5odzCBVoZ9cRcGhvbDHiMWkbrki4rZvANmypdpJRPMs
tdWcycNxaTT5kPAZPrvBIfH6r+BgQhJK18/iw/+EqWu3jhbhnAAKyhp054FJL4aVZLKSmpuYai4B
zieFhyDAUE0rM7pdsYi3LsNPtbtYl6jMaFu1y6vaXeY9iXjPKtzMj18wfXkm06+9rY1FFNU+f9cD
1eSBJLtGKtOqjQwnJ7I4G4z3IjtIZ+G2XycCm2qpTQhzcC8CIZ1LD/rh3ZvTWU7XixwgHWb784cd
henxxBN422u2wXBZEcZb/wNnlG6gJJmVQz+v6MmBUJapFAa4IAWhKuwYA0tXKJWRQDXUxVcCZa5L
kmWhv+fkY1zbf6ndEUn5D7w5W5Hm7hCInuh2XiO9qoknALdEbKJ0+EtOVGT11DPV92VSfe3o8t38
QKjzBCiMqr6G4he+PAgoRUeGXOh33V4bwk3IwvSdCwvOpfhkdnQVqdkJWGJmSnrYjxl1DgarX6ya
UTskEzqsqltb9uRmNVmr+jG5rPHWD3Y5L7i9GNGfYPpGyI4UEBSeGsJq2VnLeIYHwd6VglWFRGAY
/sgv6flq2Snm4xxrr4jS+7+O/TBskfNJKXgbmjfz5fyvliy0nMpPFQG0WKseXUWZNv4sybFRt9FU
VEbVTEB774WVqUxe/BJpjvGXD4FVWFwQfnkKN4fN6p2hDk5VN25H5FL/FftrgJCJp9SfK0l6PxDW
rZHiZE6sfIcmZNDdQqW+NnnDkUk9zs6sTZmO5vNTLBZtrHJ45n22rOoyCzrocc0VmyXZiLt/1Ani
l0O2MpRELDw0/2dtBi3NWtk08xV3VnOLwZdslzwgcnUtXVOl0/f7waRmYxh/6tLIu/hRO9dIJIHh
UTDsBRm25yx/+3AUuWbxNjwNOrLnBKkExhf7wLlgVCeov7dKEyOuWbxSg861ptz/LgWehAMKgELu
Cne9tiKY+upcvZIbkrT2s7bnRHPNF5XNlkXL1cZ+LOMujHIWEKIiMGji1IoyhSNHYayYjCJYcolN
7RXamduqdbC/dWZ3GypvWx7is2yEEmLcydvyDKuoH0gf+upLIolb9DcF1IIAWPtnpKnO6G/zR80V
d5wNkkvkHxr1CwqM12tPGGAEs1m8c+4gptROXRCUqQKJ1U4HMttPdCW7qdYUW7qSrC/9GN61RkOL
Hbpe80sUg1v7nBSl5dbi9YQfm7nRc9LW6X9swUyGewZ5ZnMsuorLJ25NbkY2+peBzWHXzHgqhmdY
qmA8vBRB+WiREFeDMGO4wvvyhvWcF+sPsO8kyuFe/taVMpjSYxcwYQzSl+a9RnLdhfBKRnbSGxNT
67vCaFmf15GnvbCFJKrSiKpQnQf2Q0aHFrzf+jWEmjWymSbZxAZFCuO4wdVQBlnHa6QpYyXznDJ1
RkrVgzAwAK3UYEqRNITD5AtH41S5FEVIhFoopQaa9UySiJ8SpetOFP0xqH+H07LekGnjpqUjdNAB
kY0YkxsAejWyiNAFakCCz8/HK2ZhxsAYWOWCBxyD4N44/fkYdPqz/WkSr0AaB4j/iiQsvlSPNtfE
T1gKMa7CDS35yDOU29cLkYfX9qoXxsb67xqmgSHcB8ppQLBGWLcHfdPbHqBGgv8Fm8GqxKtfzLSh
gbvQHWtiTFR0NfAo
`protect end_protected
