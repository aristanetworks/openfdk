--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
PlztjPytuFlpEBo/l81P2XJSRLorQMF2yXo/uFWN+yfQXyN44ZvnvyWvtgDjqdVfnxyTpSfwh74j
N5UsMBtoQPrJoW3+4Xnh8DbFrx0PmoLr2W+Z8n43b9+/nAL4Y1lWfsCngklBlkpsfS5MIRWaMzSN
Em4mcoiQ5qqy+uNO7Sh+LMa6RhgWhv1BcjYmorXo1wRjv3Q94gA0yaGHYti6VTZTnt/9qxD4ty0j
E+GOdyjH+kpsSKwq+FicCnwvv0l3BecqrkEqAXylUJydczBKTz96X3Q6+uKrpIWf7G6dQOoDe2hO
BYK9hQOwU11qq2m82R0mwe4k6MVu9zmFEUvUkg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="13bAhMhU2uvbY+OB1floJynU4cxmgu55nRneodReUH8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
JC7hyikI9GuFxALHsMWzpoVxkQE7/rsDEmmsD5fazgiKoRrMMZSRe8j09vs1D91EtnIyHzq2kMhH
I4wuRB4p1qhDJUJ1cSjEZ7e3iuQtu+rGiDIcDZSsmBkiBQDKz6Y5sQD3zkQDEnHX06EMUetFDg3H
mlYJpNh8Ibi6moqxziNheJ0bKPCosiy0vpB9KsCtM6mCpaSPl9ByuVgPVStTcRmPoX+UBg0xZxsG
ZtlXXHV+l9aRi8jm4ORbAiNKY9JvmAiklKw5VcHcp16wjVLTnwB9n4zU6IeHYAcXNAXxgBkZ6qCI
hnQjfiKpL9l3pElJdQJGDlT4ZKvUK7UJjbcebg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="hXQkcP/gnHLN6ahCghKanc95K7l5hE5ORH53xv3qmd0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10304)
`protect data_block
Lu9cyvuM8wpwyNYPEONOSaMSROlf1R+Pcl0Km1LzlstMIhWSJXCjKSImzUZ8BpP57xTHmmT9j1wj
aSRfLkRxQhdsUEvn9Fx2mgRHqfX4ejRS/dPdiJW02qjRHj3lgcVblxiARy96TtbuZpL9cHUJWz6l
P3Dei1mMmIsxKoM3QbduENn7naSX6bFtPPmEoNDTFmhyeO0jHRjMwtGL7iftf2alKB2exE6WjGa4
KS13jFqH8VJivzBrZgsDyUV7DDQc53I4lVKUhPRq8MRySg8I0nMbm0UkY4kL53NcGrTPGULrkCSj
mChibUAgjwcSyvPzK2D3cocgXaeqNK0EDUH86gMh9oqrTzyer9AVQ77g5R0XIQyJZcuBQmOUJUlz
7IHzkOMy4hLKdF7d43Qwhji37ycpFm1ZMfzbuDhTg51rYTZ8cMjzWEjuf71TcvQFuOjePAdoTXN1
nY9KN9gy5YZQT/UD22j1gJHJaiYT05rIji+9Eh7x7R4jRHz8jmwlYBrGjCkiwOsl/pwJ3G4fqqso
Lf361qGB3QV3FbTXQzWdRHZGXBQ7xT+oH48kFaDbIs51Ha10tkQ7/uRESG7kNnQ+L2mAZAm9nLGf
YIkWHJbOQnSvEKNb2fIfZIkNnHAVBeH020HblPPuUdM9Yb6Srs72X3a6yHOpG1PRpDDsOxWBF6SI
tOSm3p18jlO5UOMusjN8V0U9+w8gbBO5c5xgeKbj7iSE+Pe71DeOvFfRtmFoaJiqqUXUCxE59fgu
ZdLFa0iD/GVW+k+DLO1jydijtkcl59ltgxsUhjRixBdpJzAPas1oIGXSSM6SNEBx/XFMnxqe3Jn5
gl0StK3+ffZ8GShRJOLfmSZMGQBG+et9h5ssCQ6afllD46bJdf5q8fjxn2QzDTSgkQAA4xrbSEfu
VPzIPe1laJZvkvCB87hrXWBdH4buO1o+p86yiFqRcPzbHQ9zXaHQnn/YqrcYsjjmfyjbypRd2SkC
2oZy7Cr6grOo9X/uHoWLZcR6NaMC2/He3R13klvKhv6H//JBWbcTsD2/FGjk8MF94bazbaDuGcMY
SUHtcpkrcgIsa5Cz8s5vARIWyXyHuNC/x69lDRe6yN5gAv+I+16sKEgZ/1I4xtux9qg3eTQBGheL
cGxwUTIOU6rmJNqslvxPl2zoAdi1YcRWQQDADE11KqHceWCeDXgibU0MP0MTYNraatrTt5M3DSCI
OAWVU+ryeK0PLSrrrahPZTUJEd21n2jbn5++k4ukgPat71REukU0AQWISZmAeIr9S9Ik/ANsSPuN
KGQg8geoCRqcvQanfXocSlwgJcSj1u+ytswsTcDs2Nycy0jA8LSI4WrpGH8Gtz32TDaUXUBSEZxX
c5txKzGD1xKrx4Cwjk2cZBMwOiqMvoHyEOJNygByrfiAexG5kL4MWZauYgQ1lu9jMmE04qVQuoQj
vkoBQEOtzflr05oiPmKQd9k1E/qs6zwh1d8m+nwBgm+qmMjYDTx9iFeua6Rqx4L/2N6oDUOZfDdz
SeoWk4xJmpTY+nm8gnAIckdxVHhx1+GXg5fxIb5qsFI88AN1V0iuzjT9M73/bXMMLG3JryfoQw63
oAU2b7QngveGvB53njZKFau6+Kjc0ufBS1w2W6F5ZcF1knKsjfYqg+wD1HDW2M1Y4PyPi1WwNQsF
bwGlAtrahMjJwfGOtwpKO7LOIRbHcqe7B6nPQOvjcn1kFyOapfrBY+iiTtDrPPR57vVn8NT7dzNh
iMgW3cbhQCYIPc0rUb/AF+J0LSxXFXcU6saYs7r6WTaKUHjEyWsQuinB4Ya5tevdUnFh2b9ZLqvA
lWJv7vNnmTCs890zFKXgq/rK9bVbNAPgz4yJfxvG76faDh/biOfZCUyBdHJbOHflEqEdcFvrOT7E
jsYUXlijDs65nqIblTSZmHGO4N8FRI15zcJk4BiP9usd0Dzkg7VC8mawZ+jW+GVDXufeUkLl6Ptf
pR0KxwM2FitJJE23ibWT4ui91SpPAG3G3hb1p5g+YpiR+6o3ZHNeTxRwatlqfyQfnOgFGIQCB9eU
ElvG6Zxch/m0qAPofj0lylEE0njH+uedZZJLbnIW68Pio6ySTV+GIMNI5uRAYx930ywOeseGTj43
YicgVyBAnld4YfxRNgFUcZAnRn9Vtm6p2Oeu1AMeECBEOLfI+aiLJWr5564+6Vrcy/iopb/pivX+
Ue6cNMMmYPPCosl5J6uq5fg2iy2YqGO1bzsKmLhrgDLSgVXA4UsQvq7JZY2nefWeqbxCJ/YedUha
cGgnt2WBXzy6bt50y2+RMBq891d+ehzJmufGz1CAwJOciTtAjzSpm40h5J4fAVk0C8u1L4ponett
LZeExObVO7+Bzb/ijkY5FaDWQqxYA6STCaz7GH81MiV/JIotiDIY8SM1QOrHVX5uHe/AC718Gxhf
is87vug1NQE5gA/fRYjuEB473AARthmm5HIDY//5Lyf+vcT3I8Z6R1EMbC7zi3uCI+fff8fkn/SI
TcPBim8ttNJ0/dtDT3dpNQLGPJkKMwf4bTUmWvDEdR51yxCSSuB7fZ4aZT4O5Gq4yrzRB7wcKnup
+u4SGGDwSQKEZpQQumVeZX5h7FWR3UAEbASoJCaWjbWaPCpNvyvjzVhgCnJBytP+O66DMdkZNrzd
KOiUjjeG0C9CAIU7MBZozdInMar/EBbtFGkQWmuXJej0mjBqHSgLFEXP0+iPAZzD8h3ULIE0Tx9N
/kMzFrdSS+Kcn4YJyzcUto28FZ7cKUrRrP4Ri+iVGRr5dm9Sm81itVQEhe+7QBKtCNkS5LBtGWks
Nijm8SrMCe9o1lbkwfIA0zFszpM8gDb8q6EAApGBTf7lOH2PmJ7EQ76pU+8LGMcG1bLk8qSzrhL/
hHRchyJkrnFXCGFjWy0KS2baIWBKXV3kCPLxfye1s2kOfBRG78trCM//ErJSKZCFTL+P+ESnTnyh
q2eyL8e8Axv52ukZ93TL2Pbsw+RxSRSvOX/4PD3bznc0x5CUCASqU4FZz7yO4jWwmc+HBuijtwO6
nopqj6oBScUHEu2U0GYpALriQYEJnRym/VWJqgHY+Y3BzAs13/LDu3cjsvGkG4lDRRowKMdc2jcu
Df60jWgfVQ8TfdEXqSzcp4biUOIjPKsl0GBdor2nfTDDTgBjlk3ag9NIO0r8a8JHGtL0BUUud1i7
CSyYy072nu0oP4DidLplSM+4RX+wn8jp00CPBQZTg/yLrMpNfftI08OJGOU5WYiuBIAu9spLQByP
DZcQugQlUQ6SuMsnXL5JlMqYQ7+R+amD+CPFauF+Y9S36yL3e8wJi2qeduFHjOhjueLxM/Cwc2sQ
+flmtVSf67EPHWxCdQSk2b9VcniTGqMYfPGkezW2+rXOC7ZlPswj/HaJgZ1g0OmPqT3NNGBoZzu+
5FZnIo5zXvdhPLQutLx0wSB+estTW4Zqwb+livjYBBUQn44YmFGh01KiPopJjGC2zUEj4apRi4GJ
Wiv/IUhDKaccecPz6itqO5lPe+VRJZb8QUhyngVlWWYSDhru+c16FRicrH5ZySYBOmXl9Lf94rgg
rojfY6B0nR50sJ6aLxxGpQ2U7xb7q/98aC8SlHbh9rukqc1C/VEVjxYlEYssHBrF/VeaL1g7CZWh
b2Qmyv7t7DtCrh6RrjPoo5Vnq1JA73aazu14FTOlxQILqIjvd15SgBiU/kcXuh+463CFk77UVOeG
w6V5t6Id7aIy7XfagtaE1G81zto7+GIy9YnMhGlFBT0Ek9/btUkbKwhxGK1akbEIRxK22Brnqzu+
y8dTzLjB3J5lquYdKi2G+rlKzqiH0nsQZ7ET6FtyhNV0t990IXZO3bNoaf6Eo+QHxCBOmCa/tRtR
M90FNRANbDatlfTs788PUjUDJGkpNlKS07jahludoBA9siQZLMWsMrNLdepM+weXcxVAaWloQ9bL
o7cLdlmJ1O8mzUNiUtEJoTJgqOg3HF2VjpQiwfCWDjUqtG1/enbvj+bToIu4Jz53aWIls8rarH7W
PjDuRokVMuQ2q6KBJhxZqVA3YNj4qyXOesjl+hHIBWQtasUD9hwDJ9uYcZzJLNkLIV0v+XWjfIaI
ZybNI374HRAWSmPskRTDvaJ88N6Aw5IJkP3DjJdzIB7di1Wi+Qj1/hd+pM708y8eFbr2w8Uhdw9N
/G/G4LcZGdaVQqowoRkq+KZ82WhpMhVYM1uMSOZko6B/rG1oSIxBLtpPIWZv/q5RCZoqX6aCagl6
gVVCtP32vFGvFa4XdtnsCLmX6Z7004ikXtC1nyUeXDcFzN2K0ZQn5FHdGxbfNhq9eCDAVO10g4bx
M+Hr1QAhE6xheSJVOZYximSBJAp2RjiJOi5MS9Uaf3Dc918BVaX8xK5Eo+tLxcEGeiAFXWgrjzbq
cKgu2IAWi0oYJq8VZuSkuD8/Y3ocSjCU6wSqjdn5pRMzQQpqtII5eEWeuIA8XyH7KciE1dvO/TiC
IDBCG5TIUGdHhUlLUMjFfAD7uPoFhVLlu7t281v06MCTLYvpkfP5eN5M2/6visNcv5DR4d4wNqMG
P40jxukuaGiPH/7KZW9LP/PDo+2YMH/IWBVkF1oido37iDkVEp0EkfE/WAwQ5dlEckgpFnapqYcz
0ESVZPZMfwMBoRICFcKOrcnOiQr7i4MGNtIgMYOIZArybsSECBoND8Y6CoNzLGi0VBpLktF/FgJP
iHfIUtpr9aEdI6bWRd5Axz5efqqiD1HZbectTlOzP/rlDOsa6NTgkn6h8TtwLLpdVf9dqAarqxjz
zPcINfIMHy/hh2SftsgyK554CN96qT7Z0KPglGsG92bOoLpEqKyi6Uruz3UKCY1hMzIoMZPqqH5M
mpqG65jEjqBOchb0nAo0G1I9n6EfcKySsXUHdvbVkPFnVVEzhZ+GYFNInd85c8BNdEHUNg/xtF4X
0PP0IoJbDMdSuGkqzDCNepqIu6AuKBnjop1dBc0xvgOdTIVy6NwdlDR7IFw1kZhDUKBchleGFk7R
bS3/jxO1vFdU4rRS17wmL0mnCIm5TyNYre/vKmi/JibOWwJomc59zi/mIMQxlZOP6phPkcz/cF7l
AwsENFeSMI60zGyQAYn9LuelES5FKbm4rOe7lD+vDD7L5PrceBo9WXv11S2Q5K5I/L7t61Mf2xTi
dwto7zSuYEFuhTgWh2cyk7AiyC6eR7ZhdXGr7ZWurWqzf5/Mt0XNehoIA18XJEym4H4Iej741AZV
H1+Z4zqaLPqwEHZJNxCNI5UViaRzvPuEDaxVCs22zpftSy5LrsmYqcUKg4iGu0FStnRLCRJM7+tQ
fVXAuUsFyGX6M86mA4zZ7xXhMjjxOwGhLWFJ5XUKUz17F00s72Xn1AOa+Ty4UIY0WQb4JIxhbjIZ
JppXiP5h+FA97IBTjI+Pk4ahG7wNHf3Ajrn6LTMCX52PnlzQ5pAUYsmjgqv6SVEwMuiWjhrohLJO
rk4Mqp09fbRYk1EfQInk0/2dxg9bu7xvm89c4AhUWGbEFiw/6zdrvvCprq59s/cakmYrxtEwPCbB
gDtOem+Re4ukxa0J8BFXePSDiTjilV3Si/F3nZMwnaNoupQiUlHX3gcwcIcAk8TeuHkYBpEnOSAe
ktBiwenqsjkfFCAg40wzj7kkRXVasCT/qahCy4SXj8zrbxGT00VEaEMng5Qp2J5ZONAX/onOzER+
oCYgpbf7R6onVohB0Kuxs53tQNdljX88issGmDzcsvdMZ9MdO5zQm4CqesloARDNzoUbGgE4doMP
OftjudEezYfAM0u7ZYNUpwL7fg8C7/zUgHhsmkpu0nWEGrreRKS4upETzPHbltw+CJ+i04xQsKV+
FOcQk5wHiTPcowlkAqEg9/RmZykC4TtbXgLwBHUNuuzPDQ+m7T74AwkCwiSvs4Rtka2q4xrRqssx
m70U46H4ekdkFAoJLiBP+GuQgFwQruyQabgcfnOpyDwEzqws1QdCWhs+3DqOuz0ZaTm2sc9tut18
mItpO4+88VzXHz6PRi9u5kIiLyEqel9b/OVFj1zNM0ncocza4FrY5F9hSuKqMsvBI5l4FyzMEtm6
fO14/guJCGieHqjHxdIMWdQlbk6RuOiSJg0aio+zsoOiNsQ1AJJfP+cM2SplvHScOcsulNjW70dH
9+BVLXGQJBVt6L18FeIQLdBImTEYaA2yTrteYGAW8FXWwgt2dPfmzvU/YDw83CS7irElcQXbwFgb
vtl/xCeZvESiQ2IYUYQcMFxAN72B6om1tiS1W/7Y9hX9bxpIaCU07YQFK3JC3+/F098kumkCpxVx
+QT2SmQiTEyzMTd28SLb+hiKV5PMpGpeUmSdB3RlS0ooyz3jAVTAkbonc7S01a9v+T4Ex103nArG
C+nodwR8ECrXvQU0/CTzBC+VB15F9AJBlhet0Fq6UTAG+Gh5aGgvfhCtxRGra/DQyMvs+xW33f44
0mAVas71blEzeQnar1+7124ZTTT2q77fTw4+25qlMpH/v3D3Pkpv9Jr/bP36a64f48jqavpbopj/
DQs6NMLQ4fQczVxVfK+J/PoqEWe8Wy5uCZckR94PzJ+yWddVn1xxM2ZJtWVyuQgrojPNynF00wJv
F79phQaxo/R32J1Tw/HHVspYME1cqnONoJwqgl2qOxKeT/pRKBWrBTiwAP8GHtcTG9DLRxn9PdBq
E2EcaFNf4OH7XRHSqnMHvt1Ii/iam8WFp0xq5ebP//tihOr4cA+PPbEIeLx/V2kADYzKDd8UvkQg
twF+QZjBMdFjpLbid4hKPcUNSfY6s8Bm0blnZYZNpg6Pz9gM9rSa+/n9o9YqSzZVZzlfd0T0Ci72
NxSfX/VPGsjS3DU9aWRRUdAUX8JQkppAw+itwvbEjqstNavmlpVjZvUTPBTCc15xvc1XqBjGYIbN
qT93FZAEcB7JrElyK6qx7mCY7rfHNXCUbI7f4UOvXkkFO8xpZFYv9GaLBPzmvVz08u2+vVbMd9Ow
FoENEHM6GCWeftfsFcCLhLACa9nqeOe8aoezsb/dPdiVs1aGA/gCanOgWu3ePngwDZh3xJbKpcsa
JSPLA/lWdHou61YWOOok/mZ8YFUhhiQvCq5M7KdVgzRxlvKzgRXnga5HMX5iswikL/8ZlvlhR70m
M9QjfW1A6QknMkjwNVIRtpaSrUp1U79OByB1JRNKbTCFUbR6mLiBdSFLnkrqteLTI29ha0u+On6A
fwXc30BstL3Rt2jp3DhJ1OL/zZReMc7bAcec6zfRmcpgQHGF6f+4Mh9/Ewzn5aJxGZ9UZcaUuH/N
YslZ8lZ9LUehmX1KDQR7rxezQgYOPKh845nQN0wjlVjAJ9pzGdMQvAihfjjasAbeo2kzC9y3xoDT
8PkOV4yx+9TVVPXDdDzse8jQirO1OUwNU8zJ/fe9NlnKeVWf3UQoWAcRwXo10uLZgbSgPwXaAU1+
Aw36JQLjKf6HidirskS4nB3hXACygKN5Y7fnOsutwv0EuvWyCUewiGOJdH9PfR7W7bhFJr0Q+L/u
7W78lxmbpZE0v2VFeSX1pJ6xRmMsAmscLa0nB9StKy41qwxiYBg+sALYsRj3joTOe0gmCcsm/b8n
SGMToXVuX6mErS07gX86hqHZ0iCMUmOzL0G9vEdAJrU17FGUeGeoJgw6WJW5lMumEYKswB/io0U5
qmlqOpNBNEH5tE5a1sJJbMnexYL5SUef03nIAlNMKbL5EkmeHA1o3saGoImTzmcws6quV3089W8E
N0Ulg0xE/p4K5fMB7bXkxqwzuPr6bPY1vNKgB6vcbOozALk/XulNwymOp5j4G2G3ioKBK7FS0bGG
CuMXXcP+QQDBVrWNy+ASAKDEWmclF74rfw5P9TDQjLttvrYh3PR22NcLxH0nkJ/1oVaByjaKzmMQ
N6OHPckGdANvJagU0eltR1HuwZ+7KcCapBWYmjg9s5QNw8kBbQA82VwNO9L4z+4EcbHOcVYfFLOZ
mEOKjDfU+iDA1q/Jq5SWt0nr4GlPClAyd+sApNipqDkSrOFKBJ+6HqEI73XABrxkT947WiSxWxwO
EuRsMF4OXJsVnAbcSmYERd75jAacVixO687HtvmRQVvUQnQBenMR4DMqsCIYWr2dJQtla7T3yWed
7YSy6KkSxpKtgqpr1aM7HEWgLl50tCEBm7lv+XGN+0l14jAJ4/fUhhfFMR+mTSH2IOg399ZIipq0
khxgYcOwyHj33DX0UO8pOlFpFuzLpmQ54BdilRCYMIxhnwsGYU1wEL9lDKbWMOV8lKBG81Imepoj
uACxAF1nF6xcFzupf5lQqbA+aO2qQGoHsaPqJHyzFDmaCH9iXMd5lZG20Fz0JpDuSP8Pa0jOcnJd
Upc5tV5jcTVIWLqox8jCbsZTD9pkqqGibL8cgQFNL9a9WCCmOR44fyaHAxtY07He4ax/cJEymFxl
//SDInUhreSZjiTEuzc/95YbTaDcxFnrPJf7ibdvoAVaTvFGBLMRx7Jo3i12atV6mHfuOr5kER83
g0zjI3pKwKY7S5/JOzcCaghbDpmMWBybqDTN8VYk/+tDosaIe+JYhfir4+VyZCR1AjZNUaLipuHK
dKe2qVeWrnn3yV372Fy+oL6GPWzO+cr0DNHLLYgsnWlSKqqdCUTtE2vc0EII/EsFpyRSTzvLsKP9
2t/lOThpkmf7jPDzzUOaq+1MOgMZIixAkmQZeNYmv0cxDuXPnEBxiFd6w9063Gx0WUO3W42Th2ef
qd/UBx4xoZhmFcslqrQ+33XNFJBg0JlDX6AtrIXbb5lU9ijFTaYHqe9rUXWPqY63ZKvlC1lG0iu6
0Scnt7U73tLsK9tYi3TrJexID5TMTRIOik/Yl4Xu96A/2FPh7cEOnLTOTXSU+4h2Y93QrWCnXwlw
XuyoD4ITVErNVlI4ecgn+/Ng40OxcywSgqHM8eNZ+KnGmDZAVQAYifBBWT2ZqqCF5HslhutoS5GW
4VUeIabVRvJ3KjG+DHnh6CUYq5kdjmk4RW/9SqS5w6snBftJk5Pzj2HC7SzrVgVREBgTC0jvDcaJ
7vPa0Pz4LAd09FcWITh4FYojF6OhPOypMecqIh/neU3A6niBtrMS4sgWs1cMIVczJbp4typgQg1w
kCcfXQffzTwS2hp4xBAMisz+XB+hH49U4B9U1ni5YMrM4bTxOQ6djgJBXn+ji6O5nPzBV1CzoYiu
8f9UAe95btLZi2jsrU1aFuoMTEAd+KIRyuKwDaCpRjCCVFLWtZXMGvm7bfqVMdRWZvQItydiqVvN
mu4ZPE5ZnPI622dkAkkKVngrLltvudn1s1mq1vt/5rqUexAGbjTYHEQyhmvATDPNoDzTeheso24w
zle1LY+0U5Wk9hPluTaYwfC2QL32SwKIzKXfwnmg7cFg3Z7IJrk3elNtPNkZ2erDTkfunPViA0rs
f4Vkps6YtOFumqkhD1oZxzs3rdtt3xG7KXLT10gEP8QphWW0lptwafP11n7iFQSWKNR2edx33RA3
xBWRc00NQpcbNlEJs/stxCdT+vEewb0mk7Foq4+WCYfhydh99vX76dxaNjjnhcj5iW9nAwh6z71f
gCAobsICnileNyZU8X8hUYupS+V98hI2jUnS/WJeJ4tkIUpXtrm0RZ4AFjaGC1XfPa5S6MAeogPD
4Ny4TT7DloH8gecWQ15MVR0+8lbG/qzN09vmYgVCppdBwFzI3p2yy/0rXa2STn1xTGijaGd33kiL
0+SMrJB9tMAPLanOga2HUU6WIRJHRMWKKmTEasHvaRPVlqhMnEWourn3cJ/G9PZCFFLF0/93czRo
LnLMbGd725RGAC7hFvuRmkylgwX3z/gUp3O5H+Da26cCjk23O7TxoMLvseb0FX55dEI5q021RTDM
s+JFLKb7tj/kqAaF4Yi4ddFaqNmC0xMD78UTnYVobKll+w2ts2Xruz6oDeKLRO9SSr61sT5WPmfv
2LFTq6v0SRYpLyxB2n55vXDsmf4KIZHBMMT440X2T8bD/Pk1CKmkYl0uoh2MEDrzPKmYhJLTyRRQ
FMYs+k9Hmg1ZpR9kUCq77nLDYMXokTzAfWkSzP1amp9vz7JxXkVtOp0CPbgmK8KcAT5mnzXDXuiy
kmDnM0PTbVZyQqX7c9BDrJ7Mh3t2OdnCaECbj/Yjrli5Woo+S6hcGw0ge3pNDmd8wLNcKVlB9pYd
LoLTtkvKuixlimYyBcNIraHPs0N68BXhSFJv+hmdFxCh55C9AE0aSMERhMn+uriKEpRhJIrDuI4A
Vre/BRa6qmHbEY4SGTXNKODudKwRzOMGEikDw5Ej4/0ACEGVtVyie/8SP21IQGxRKlZNiwEnXCtc
rtlSC5Mw0tq7EWYA3s8xqmTnEhqjZ1Dh18gmzMObNXkAsNhiw64j1AUZptbQT7JXeuVYj6gqDgzv
dn+tXUMnL+16AzFmiJkUXADwJUeTwjj1IbrpKs61hNwJpeI6SNrFUWMPrwumwA2/Ik5pZViKTIUU
365Bm5JwDqk/bo7DvYAMoPoGBzxqW7tVqE8f+R6TcRh8o1DyhqHh7uHY2X+tRKVvXzERBLnmsF7w
ty+6S4USH7ii8d27VmwIRjthNkNqtoi9294O87PJUK07ObVGPgK30by/CXgDsf0NcEebhG2SuKCg
nc2GenOhDHeiWxf6sK3PIpdRpTI75Qz5cuvS4pgRUtmTVFJuhyG2GRj2YuyNvWNt/injJFllximL
ayMPnHOCr36JU+Ior5yifm0nhYCbbbhvsna7Ywqv5w8EyGCNkqqYFhHLFtEUbMfQxIAq9Thlfa7t
TzseL8A/Ca3FAgW0SZXr3LZO0vSXEZ9HhC9VLFwQwbMc1GxObAx4Tt07d17HXq2yt5Vf6/Dil4Iw
+ElTeZ44Ilky/PlLtZ/EfbUejnLmuYV9n1TXzpsyde1uBnExIpdjL3LWUJPmevJa9jB4FhG69Y/9
JzwO5ZnQP/e+uQDTdLFUaT7CFhZ2v+U0jqbhnhNt2UKFvjA6PKYoO+wEDMU/Jyp7WXq5IT/ie/jp
j4U2XqFPNyHGfjEIyFuX43P/uzATCUG0rA6nPVU5j7aIfo+p8E5EFmID5+PaDH3p1yA7J5jOe9Oh
n+2B5QD9lsttE4FM6CpRjQFhvSMphetJpV6qZLKQdH5UqDkT8BGq7u5CroL1l/HhuctYL48trgiU
WejtoB8T8lsJywW/sJ1hxzXYkh7hUnZ3PpR4y5HxqYFt8bOzSZmdZEzZSXPsh3YG6e34zAnY7jrp
S+dihuTuXDrpRGHfph+wWNXTMMzR1ylo20BwVoznTzlo+5RPpqEOetx2bj7XVoxwRVWPGlkAnTfY
+PZzGzaBEyW7iolUEnCRtcsh51Aezh+HU3k6DMl2l7rssW6VuCuLbVnq1CyD4UyCYxosWHXbxreT
w8BY725CXR8vdJp1Y0Z+VDMeMl/vg/kxl20F1Oz2vzcvPgYxgp0Y+CzCmRFuFQacDkX3/hQv+ebV
9IO8OverQ4weVm3PymFEQmwSMMj46GyUXA8rjut4rav8KtEPgDKh3jg3pt68wQY3pHux8ISM008F
6am/v2o/cgfH9k4NgoO5aeYQ/7YagVDvuMjJ0pKwBFeDFKV4d/swcwZ3Pk9G0EZQbDrnzh4F4hAZ
p8JVyKuascenyugTHThqN9g0ci690e6qOYZBcK7xXPhlO2xM2G/o8eKmOx4obBuQCT17+18gTEqa
idDdPyMAd8VrEdVdYV6nWA3/1hsW5qqbKCqRZQ/TiaOGbdS47BN/drry89/q5wuMfohqyTH2jTut
W1uQLCyDModQJ/MLE9J6QPCEE5XaHMsXF4JhZoeukRyQx3yu0fwxQTZB4dkJJYs17USXGMdjFQAK
cAARDxQWkZ9vbHaL5IuaCjdo4YbXKmqKCgxVeR9YhrAL5jnakvpL3MhjvIGo1lCi1zSp2wBpgElc
iiSVyKWzHeE5pzAjy5I2a0F6v046sAphTT9MDb5C9EFdkzXZN0M7TtBu1V0nTtxbo2XzLZIfgTT5
MYAK8EeNl8E2oVP3p2yCnD8LEJuo+/0CcHz3med2VUU0fjr6UaOYllKI9uOhB/ImFg9cmSj0W7aS
8mN1yuq2CkjOwXWP/gq2iKVG7nY3HqXh+ee/QeWAZ4S0Wqyt965HBDwUKAkHWXcHM0lv6Nq5/pxB
/Ux4HfSLk121THnHoU0xLMfMsL49wNlOHlzXzXDJ0SO9cwEZS+eeTe2TkQThnqvZ0asRx9dKYgyP
/FzbyXtGk0oSEnrENlos5b58d9myezBHSd/BDmsP0iaceGV27xuESfzKIC3Drj3oy1WKiC2Gpa4M
w68AwfYByn50vnzMR4ILAGib1h9m52z2R37a6ijwvU+MkaDEyMFioA4bbShhJmU+6/D0LssicQpT
Xix2C/I3oXay4nYyz6Jja54QsA7QrLVlFuA3yPudoT4gyHhAiD6gpAmZJEX9waQpBwUKUbLvGWAS
5sPXcTsUdze9iopVd/wj8dsfIF9UQcTTLO+KMdLsi8vSDDpv8rv/h15BjgVejrFDfR69ukKFu8hN
uItrFN+yGsdBkztjEmosNrnEXBCd4mS0BVK2oYH34lPtCvt7O7Cv0Q9jHQehKi46SLu4BFy3hH8D
uh0ivpB54ilSaHMl5vv8QwrPBMWtHCCdZ9sPeCc3z0wI+YlmWBhdKTDeLJD6w6RaXMtoALfbYnnm
X7a29iZJ5HIxWkRg4WHKqVFif/gyQ7BoCQjLPYDcNW+pRAoo7SyIZYfx5NWrYDKSfZ1ZeSU9bDdt
ODQ3VT57TyWlNxX473vf+m8lu/UcLHLU09P/3NCLK7rjiPr0Ma9WwyCXqhQN2EjpykIvjOSZCwZP
4ms9COyTRrhWr+MomF6EfwRLEqLnKqjmaLnqJk7hB0GN2G9AGhw+Gvm6gNiEQhHoB8BY3O4gZsIM
Mw481GV2FhhgN0it+6Hj4GyD05F3ATJ/mI7tVUn4wdv0iUAwkAxizSlaV0/nK7h2KosqlgTQwdac
efBYOIFLXJslGyiVS6Ntb7jpPw/vj3nDgHBSabpWUH+k9nTugKtn+bO2kvyLeoom+bOABOhRr7TF
BmU6O7QeiKqOukTKQsBYEEbh9Jujf7S/u02iwFRhoX3Kxgi4szqWihRNlWj60mdaGDnb3sO0anXh
2iyo2AoRHJFdamzS4TDS/xzPcsOfxJ5ftzc1pSy9SlcCsR+2+NGf3rajA95igMr8sWG4G0a6MLZc
yb35esMeNAH35czXpOsJefrc7f7A0Jg1qXfVoNfXw6fRihq0UjjDdk/JsJQysONpW64mj/KrXcaG
yJWSrDiaE7hkl17CJZOEw3dLgfFM1kN9h1YufmMqafP8cB+0PNo+5YHeibiK+ocnmKQQfQVlQna4
gVhf8+dqXGryYoqbV2W9vq9KR5VZ9Zpyu8byD2YJwtojs9SYDhe3Eng2NKPnKyLJnoNPR8/CLM1h
paWS6VoBNTrpz6AVcMZrXYAzILSALJYzJ9zx8myhmvQH8P9IhHvAAqjGfawqa6ufIIFLOzgVHO5g
dn9t4q1JZ04uVnQ9rmYQ15zRFWsPvYFFze80v21SotNxwZ8B6QMPTJ+1FylRAxUnCr8vkXNktQ27
o3B6fZAR5s3t1sQGI4zDd1Ap8TZfaKZlm2suKc6dZTEm1z0qlKsJM3Uc9IyUOw58esuw5rx3tVr5
WLYHuA460FtCY4gRH0NjyqSWs8MhWex0e+gVEjgg1HpJ3Y57ceLakrHmPRM=
`protect end_protected
