--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
UQ5VtB09iJp6FOQulliZHbiH/jfKLtOXjLH6+ezRe97homvZW8ixPauF7zfv2CgHnwbUBoBkJA6n
YiUJVpHdSN38YkY0jQj+CVWAPgWbsimfhQQMLBpZymHGAVAyOcBYfl9XB/gxu5MFuT4Pd6JiWcKJ
7SVMAbOC5UKEXh8OjkYo3wkneesPeMv+5HVHbOJX43mhCH6vhAcuJIdJvILW9YriaqYbPyDzE1TD
gtN+6CgHGhqz2lB5IDXiNXBpy/O9Vxrp8Yj+seWJ/953EPOxI+aIjBQIrP4H4jdEnBb3S533DKEo
vGt57ZpEzCnPVcL6W0f6TJKo9PGdzYarJM6QYQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="jcjVRMswO+GpltkxAjKBZ+8wD3U0A9knpj5iVQ9+jnk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
WBGHVHMvH6czKJic6jseL7xW0kFGXyK1YypBxJzWjqWND0+eFFDyRseFO29/sfldbXfdCeKHWjKj
gZ6ZrvYFrcNEqt+KKD1u9kcLMiy9jyT/vs0Rak7LGvwAcAyPk0t1QYU5bbympi8YKikb9b73aTxO
AQx5Q+Q5dSL2L1sQa0Ma8qYtDh2KOOyhv7xe8pPgZNOeKChWO1BBa1+Al7UtTZu20ErQXkhYgI3P
nhWO0MCYpkuTNUgDygnnjII3MTiazBtrGAFoHElA/k55BQ8ONv7EQL8bF+DdG1IS7BLQ52YufF0e
QgX894iO8+QJgkVb2jR9K7DclevxsUCrb+ZE5g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="1ianvkmZym9s2FaM3r/uaeeJCDBacwpnOK+CH+/NOSI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10912)
`protect data_block
j3GQx0agBgInBCQqouNE8Jg+/5cEdvs+zQx44QcBGRVG3EyXKfJ3Gzr+uw38fonAGALcsVJJ6JtZ
Y+KeK4OT5xCKCsY0MPJI1VfRNDWowEPiV7qdRj0JWUgxL8tIB8YBvqsJZZszor68i1Pmi5wR+kQA
s4KbtsW+hTIEAZhyZFBTnGeIfFD1vpRxvg2/Prc5+EBScTKIX3gNLFbfkq5N7JQbVgW1JpKCIhka
ajaoahqTBebPD1+ZPVoQCf5Jc1n2NEpm7xli2sp4osoE6Uz1RFy9jUS2D7XqobuWx5hjGegflqzv
ENbIIPVbLxyttluggGkHkXwy5krWvRluqb62MPXbQopQv9Pc9Q+kylXl45Tr5ByeOLK8YoYvWAtd
kFKHVbK9WQtUjAcE6G0KYmnJoUZ0rKvdWPmiYmaVcjp0dSe2SzCbTymYe7WBfPqN3qcIOM0I9frZ
ZoXTwF4A41qS3kGEYBSUqjDuK8BuEpSLQzui3+g0kX3s1JVlQJQsKWZvo6n2M6HSf8Rq95QRJc4F
bopnBTC398hLx244by4RZE7Z4gBD45sfFNXf+fr9eBsFw5alranIa7e7dreLaN97UmDb6Pt/A3o6
A6vextzJtXLrR4g0WXx1StdMgARl0+dvRIuU+ivLTQr1HdrMFQsAqG2jdEWrUazbksYxGaJ3Orei
PCOK0lgsTSlsOwYB5hZbAQWSyQBngTrTDrCCWEx8cBB12E4hm9CW9ZRCleXqlIQPHCFMchfOczek
ybUPEdW0OOg4ZufYzjLVfBy7nkvg75TVSJ1Lixee5DVKbdtdF7t3PoPafnNuu822Yxjq1lP4eZ/A
qUb6yQD8k40kyB7RiWTHZPAORH2gGpWWAdHmrZ28dA59WVZxNQQH5Ny/aqcXWX5psQeeXUlyWBze
rqq12Sj9UPrhBlwtBquY6iJfUGcDQL4N4/FgnI0E4bhr+28zN1b2yccV7AWV0PIt45Lzxo16GWye
RaL3CKfr9x0hzpIEUwOXZvwqYu0s7S3/CHoT/wY0FpRJMYcGg1oaHjbjKLH5aD1BYIpEeqgYgukD
P1P8KHqJLMYeDODoCHhE1xPzKMVrvD0GyWwd8ZTCfcZ33DKZVG4TBeT6mgs7k+Fu/6oei2JkIJUZ
metWyxORFIXImrWlg50Q3iTW9aEVGtUzhqRB34S44TxYGLkscPFLTNGLVzkoqTCrjhgSDFunSjlD
Hw68JIt4FdqBiY1Euz/iyUD7bb5wXQD5H/xBlCEh8PqEZaWRlFC3lsN01QePXKMDTxWxULDFjbMT
Ecw1mma6m3zLUGb9Sy74vDuwoQGPmPkbPqAO48TeE8F7Dos697JPfRBpauLwfr9uf2340o0x+sWY
ZLl/mXnokRNThbEUOLDLmTnxNchvwzsUjNByGi66kifz2QMrxlxNq2Ki+wd7u4cuPvsupNLIJI39
2C/0pe18++Gew8PfErF4PqUsqWz0Mr8uezcSex0XTNwYEQ3aYi1g4yOZeZxyA2T7dBkNrh2QA3Ob
S4maPn+7VwhpelaC63nkUDoBZFa9cAnFLNLheEE5BkSuUfc5zL6sUchLIfepKcKatmrE/RfaJ4/z
SPVoKLpSCA84/eXTM4VEUsdCkAvNWEK9S9bHTR78uwH5X4yNcMcjZNVKKRXbnM5gkqojHoIsBMvL
UOwDb4zcs1f+BBd6c2ysZF0Ih5IhNmAjbpjpMBCPf/se43/UYlKn+MbWIaXOAEw2mQ/dBA35eR3O
leHwxN49v+sE6An6CKnuZJsjA6LnHQtDTuluoPjCUg1cm7CbxCvBD4oJ+CXgcIRw6WGMABFpDpCB
nijlBmD0UJ+bNOCKFJPw02Nvo0GdUcw9eTD/ZdQGwQDULs5GsUMwMLJLEhnTfKamgwq0AeUnZHDF
HQJY5q/nDHjQsqamECA0mambuhvU8oZK3F4l7xRtuVACybsPhbkhUY5YShZHQEGuBj3IsIZ79DEg
ZLQWb0SOIT6K64YrZMXNyza/501y352QHakg7mkbD2/USKJ09OI/1dLGrweIruRXlL07BY4izl9y
4+E8hQ9e3Tn/mqmyODalLuWs9crNZ9yGKLAYeSfVny9zkq7yoPHX+HT8Tt/DvYc2BFgQfKE4essu
6RjgFsvf89QexskJLJfXcI/UqMMHJjJ03gtoVtkEk3ry85MF30K5Wyhn7Q5BbAgF8EDttSMdfR2s
s9zoLu/6lQJj180yTcnEDeWWVqPOANrhNFWZN0AgWHes7MBhv/tArne7b/qhsfmWEU/rItC/LABN
YU+GGK2GNBpIY6lWDhptDih/wP0POviUJF7o5HloYDJWDdwbzJzB1Ov47KhfVVntZI+VBwnmaObo
1A2Ix5bVBoTkz9N5f7A4iNmcr5dHI0psITWoVuOUQFAwNmsYc8sQsyIzRTNJpii+eVbvt7YYewvo
mjBS0mE00llZcstCFNYeu0nOiPLlENb1DWqGCHqMoDKhd1OsvN3pklBk7LPopKsxOsZVwQwd5I+5
Hn0i2S3zQE9fEaxFd4sNGZa10UKaJjGUJF8LbobnUCfnEt61R2JZSzlLCPklJ22e9q4ZtNekSPxF
VHJucl8sz5J1SA00SOgnU1bEKcFcpB28C0VpIk49cyh2UJ3Ms/SM4CQXrMme29E0UPSnr3B9299e
VYI9+bTEKK321VvecJvezL6um0VSBmLqglmeJ3Dvge71fJalqfnwfo2ZFMtaiSoMCBBlNx97CegJ
08AqUnGNSoXJJR+iz2uExaYODUO+EHQU9hUMizIYqIJTMOD/Xg+auO6AEtpoByNw/pjCoNfnu6VQ
k8bVWwW070Q+lIF2XdTWl+7UWcLS2UBqv9IZSNk5QxkRSLCY+9BD0PkOFDsO4KLSXQU1zXZ99/CX
x+4r7Sj4hCUBDIvpykRnf1HbZHNpSai7phSbZlYXICdHtzwBY547GyQGIvm341RzM80rnZdQInJH
EZl+n9xk9RCB3/VzlmF2+w38jCAauNCMRfyfQXzjlsdcpibGtn2cdzgjdtG7hOEKl0fcVyDriEii
hAWOm9PDMrg39jsbxWI4Pfcc8AQGkcPh9q4+q6HLkQ5J4wCDbSm2EThgpU4SZE44b3oPsLRV63IT
wpLAl3mgGXWeFS54E9BEZvglGGtgyy7aV8OL7g+NMbqaxd/9mCr1s5uAnwHYvgGtR3n3zHc6zw2k
lSojyRFxLIOynufGjQnBjNZx9abs2UITBRuah08Oc4jyW0dJAWTNUQgXfzV5TsdeQxhuEMuqeC+b
wXAB1NyrzJ2DJ0Q0W+P5Fdiog20IhDzVu0oWjgmtdgxCd1KW96eTbVSKRE9nlO7ITtaOMlQAgcqU
x4gCmJK0DvOgwMc/vKVpBEv1HUmi2ZTCpgVq5zRUiZEqo589UK1UgceLV4uOWcvDKMVBtNPjB6GL
k1L+M/MReqW06TiKAkAbYT4oh/Ti1gXkMJjuAL/aG7LUVU34zkPkwzNWM1/I7LPTPNQhjDVuPLns
c1KjwEWlBHcSTT8G4kNpmxkBMhFTkmC3iIbPBrgHUoRFjvGOT1NbSvnZ6cnqi6o0JWVmiUvVe+OJ
oXh7gkqLGBj6Z4VJWgeQrm2/lDSrn4qKUTWASeoAo7T1Vpkr6wThRH+b9qRbxiDZUDQPzXpRQQ2j
cZUQY8LMiPKymYA8TSMJ5N+SmHSIoyIS2L3VkcKyQzxF/mM14MZKDqVcPCEhJmWHE/Z8I0GqxH41
7IlQ6arfridxWUmxvCfAAt4qMCqey2uO2QiucCHl0taHBUX2lol2iwxdMzDCmgAIS1ugvl/CiVrg
RIg8WS9/L55ou4PXFd5Jdbak3tUbbn1SeoqA7Q7J6tpcRXY5bYSlGoEX8176TCagWODo/7GpGRal
nhy3JP4bYTyyq4B2EtO8FcQ1I815Qo1NEAniiiJ1l35OD4oanGqlgIA08MyQuwmnjTpolPhsKBrh
OscBjJhHxhgWs6m5xZVgB3L7orjhx4c7YwG+HK7gGLrdPxndH6SwYUazGSYCK3YMXK1SBzpzqo1r
pyLDnFjFBHFZoPsFe4HgWOY1t9LmLR3jBPGg/rysTiEEZWIFdeV5UopV+1PcLHwRjgrGdpLkNnXn
56K845zoKRSOu7NYLvKJYvcRzCdxSJwQ14NhEwLQCM385e3GsleIx7z6QQvz/y+uzhDF3nVe4fn1
HzQUTvwqvdkglU6qf1IEnfGKiRzQRoiMo8z+hYpMjJVVgnGA0KzBHuIiFWOvPoxS/REZnGz2jec3
9qxyxdtoNziM7hvxXMcvgBDyQ5V5FcF+eRo32Abk6dsBeNlrbA4J1IrbWu0Q1DcuiuqPenREVc3S
SseJhBaOQrsAedzW1j+sSxTysJZ5Q27YNLqEHUNIWdXaECbMEgPiEXY8dsuqsQN3eKnMXltxuPau
EfiLnhcIAwkcK4yITHCHDT/FkUEd9MsBVyiQO17B4MnQieKAy0/zGkPXtwoxnGShHRW5K2HhHk5f
smw42lCRBuRpgL5+snPpwSRGeMRMPKtlKiUnXKVBQ270i6idWhWZg39JYYi6++PQCdknBFwgepjt
QlhlPLig1/BRwna5Fuz12gLmH2QhyO3d9HzyEBpZ2xiUDvWiyxelhnsvwIg5OzQzhKLISjp61z9o
FDqjPWhrJ+6lG/dkCsVbDC2D3EM6K+ONajx+x+TWuMopov9EtH02P2Xo1hFq8K51CirDVu5PAm8j
rkyCMT8N4ZMHQvcfwcyLbIQF2xkCY4J7KIHcQFwCedjd7eU7E0NDb5bGoVpb/Bp75I6l1ZNhROPN
yCAXppKPaa4qvYJgjg9pCLxuyn2GhNVHf5M0Nl3p5koMNhuBGjGNDTMwDTgJRW84zAzU45e4QieQ
ySGRjH0okxcUVVueWPkfaWxonQiUG0UZ96LFa1dPHHisuF1JcB5YJ+X2g31f/J6/IHes9fmb7Keo
t0aHOXMb0GqF5eYNlkX8+JOHQxIuTKr8Qa2eemlpRXMgeAMDGEUG17f6dcv4loE9BttzPfn6M1i2
OVYr66qOyngel0cMf5IfFeEUSbL+mcPPt8BR/F0LfalTKY2oS3sDO5cMEOQiQnO7/d60gxbvU00v
H9teyioRwcASzw55XJAL5xIOYqwgpz/VxvSYiDqxi21uxbfD4ueYF/iCULiBQWrUe+ScQHeIgmcJ
X1Cr6u+uIe0hyKrfIhuAvw6lixgyX5r9/9oEF/YHguVgJFrY9hiFwgE9YguyWse4fBMJHsP9JaDf
lpWgNAg4XpiOjQURUKkXXzK9kdKipNXuhB2j4I0cwtthzXvCkm6xyrQxHfdst12EiBPoabhUhYXy
JLPSo/ELRtKZhN4S1AbXH3pM+Im9FXDuSHch2xHY5rvc62G/DJhdViAtDF2F0m8tAtKlevB00oj3
OQfIqdscOUmtBZrll+8k6tp/IKk1mvIZY73LWbwDQJB85QQRS8YnXBHmCv4MHjsOgb1nqGzo8o+D
/Jlk4n/gqNy8XBNe/8MY0ZcghmbQ5mTxFPOl1OLCg0nzsxprwhdbYUmyH9i2wYOiT+jqPqdUM9YA
rXncqJXpAcz0hNkEgvk58kLtsgPBZVujrwXcu4hzemc67j5q97c5HmEpbCr/Ecb/A8yMSxa1gh6B
khk8S0PAGs4h0FNmjV8GowBT14w8il+AM5CS3zCQlHWPHA/yW9aP5DpqLTcZnuzKMLmg7RTI+ZCi
XDnoh6bOb9BUtbaRJ5J8lPkbaqa3msdB36qQUoNbNjZahheYGaiobYFm1xAjf7eK9LO4Md2smGRZ
UWN4ckZpPYebTdUej2QJpSOmQMWeFiSMn+RibA0FhY4kfLFnyhZ17ov+mS4vjUMbW9EHKzdQH592
eCHt85hY2Z+7VXOwtF48HOj094aItMPHAr2xfDIhH7Cn/2A2jzasOwF96SFRjRXa1UgIzIlwYgmi
WEEOOkxgndjyXOfbD7UOYqmUGuQcA5S8J/4zs3d47++25gX2V3JIPKILJCRmt3dZF3k3zWvOiMUH
cS9w1c3uIPDqE1AdGC7opKFVQsaKDFGHkmnWfM6+NDFYWTthZTqLUAYGBl4affes9oysJ8A9MsWh
9mS0XivIAsva62huug8jlIxf0xA+ksetUsrOYhj29AKuTEnV43ttx4YJQzMcVargQ+pG/nGm7aU+
V+Qq0pWcfLLOAmszjDgFonMVjxylA9279bmlS2Pju4V99OGki1+Q6CGyL34dO+z2N34zLzRKGGCd
5qBvkzfi0I/A3dbmdc6QbtpiUUy4J1XY3xDWN9LRaksZvEQ8VAWyHUyurh7KhoResbs1FGY2eODC
pxegAe71kA3vu2tg1jwHkqVZW1jMcAjhmj1gjQKRp5QESc0Uy/uFtav/pOT1haDrp+L9YiOfIe5J
pNoVrFuVEOQKV5cBZcP7aZFm06+NTegSZD+WQNX3HPdOiWhF6fKcXmNzAJ4zwhQfd6qaHOvE/Rvu
JkTaDChAW3BofQP4vmjR+sP/GroBVTtsCx3FZqPVjUpJeBuBqBntca2jZ7UpGnZ900EGVwSj2K09
vU50vT1Tbl+OM7CBwlcRMPAaSz+QcsDg53HANg/CFpLcwFJhI+i8J10pfnFLP6Ysa2j+g1HvL7ow
rCQbbcjE77SIC7Wf4z8owDzdH8p9bICGGc/Aakiq7LFqjN6iMsKoppqjmYcbOp/LWJKpZB4ecBJE
L6IHcUnZBBxNCZgX0B0ZF6sGvVu8mp04TXFi36+mryb/bYFreQ92ziQeeErfMk5U8HxryH/t5irW
vLAs23hPAY2hLBTrxYYjSfyP5S2SCgSElb5D9OB336MdCc7ZnkYuKqPj7/trz5sGo3s4vENFRbFY
ZmIN3MhCfoKwJBlGps6EsS58/fysd8j2ORCvuIyICFzA4HqgkUxic4lVrjroT7iibi/jwfbcPazt
nj1gQ2plYMANN0giNzfCw3OdJwBY0FY0raUUdYeeT/WIDORWOm4SmE3RD9CsvXyWKcrFYXrQc2ku
ikNloRq870LflCJqoxvbVsXRu6IZta9NpBmuphfxqzQZuTEzO2tvhQq2Io9Jqhff0IjMQqlOaOgf
sGekvWNIrMeJKMdk4oc7N55YIVcX78R6NukPYb9EX6haMIEpdyrclbuxHX5hG3bGmk5lQHywtFWN
TCfXFzFltpiB76KDCFrhnpYrmIK65kyNbAUdCtq5EjBcmGLtO+R8UvlGX5it25ugYQ48RrPHWvt9
FkAvnjbknH/mdPZwPo2vRInWfxiOvRGrQCVX3YYbf3sWKPmsdIZpnJwibsM7LtPg131oNExJisSo
xZxZZkiiJsgKNOk8zrV0bV5s9IHph6q23vj6gjakdZATnKRG6IJa7OGmGcLvM62fNeG6w0kVurbB
bHdP0P0qavj1lq7rxEIVyks10D/zht0TwaZDbnKHQYpLYnfyzjiyLgo1GsH8lqpIX7da8GqU47g4
qcx65FduQAXaOBua4GvjUHJVWXvZIJsYC5Z9phxseUTJnTMejvkrab7P4TbUmISetn9KLhF/3kmr
0O18vNUfeL3qkllGKzkHTDEd3LDP7wS9td3Ujg2Leu1KSFhmAjIbxNtGs+fFOb135XXG+nsgA2ae
9/GugxOkX27iT1RZcnGw/Wtb/dIKUi1RN31Uz0TVTTKtVetIIOJhygh+oxIpNWZTF+1coRTa8twy
4ekFb6XgHSGVehEqoWwIVRLkQrdrOjmuUZhZ3dfRcVGDIgdEaSQCH5YFI6/PniAj/KqJTtM1/PyE
wIUS+BbCcj1d9n5bIwulAJbN/5KnbSySDDM+nmcfAWyjmag3K6YK4I7KnTZ0DgWkuOKjS4NJZKKD
bzRNCu4v9by/COfwOWuhre1TEn3Pp/QueFdPuUbUiq5DzAF5REtC/7HRvrAkOUdNoW0Zn+5nuRHh
zY00/BmzW4V4rDDTk/OGyy967SaK4D8W4sxX5BF+toyPtvVV87e6U2zzNQSNdpY18+O0ahqx3if7
2+Y54E1/9oB22KfhyJWgJORQ3WPKWlmwbfz5O6oI1ZGIvUbHzmZ2MvRTw/xk2cQGK7trspwDEWl4
6m6g4cVJi2O8wfhCL5PEOreKytcUQvTXe1dyEXlweIo4aQcLwOe0AjW6SVqg2jOQz6WwTxnbTP1m
IZjX0TPxbRAnVDPwSDph1TD9PBsFquaxtpkkV7jzKV/vRRPzUJkkuj37VbYrOsDl6une8caUIlY5
ynVOSEbDo8wfXHpDS7tIciWgewN+kMf+VVdItGx7mQqJlGGHxjWc/Tf7CCSTTDT2QY+sTXFGYTIN
MrUwmFLHrSq+lsJ6F0WPKc20B2Km5h48FaL6yKIeg87R2KyLIicQUAbayRn+vq0Rl7FqAT3WVv4x
0jwCFB88TVwl3ZymKHqe/nyepP/sE7PILWrdVmVv47zYaONT2za8B0PJeoUaaa3AQY1koh8Fvlxe
dpnvVZVCp/2vV80c+xp75l00DjIzXj95kCjZWks8YxaALL4NClIBNU03HWBl2bYsSgKSrKjkv4GB
0BzwSWsWgkHOur7kMMj3RK0XSKseJZKmREBr1wCEXQxGDgpfJU1Aw1hxaLy3bLuAFbOlL3ilpctg
Dc0bJS//peIpqqlrtJUstwY/rvQpCtyO8My9S8G7T9OUfpEBQIAKt6QrYj0KL+z5rbbrRUBsOOar
nNpgQmVcY22RyyK7g23doqCfB8RE4n7wCaoiflI6Chpn75wQgwy8eRNPRKmiNAU3JCs342c5HTOM
pMMp3HLS0IWDa4CS9yZ+5Bb0xj8KarYgEnWXSM8qQ0M5OgS7LNnecJq7HiiszENJNWaAMch8GgJk
e0F915kOyga9PrpX4A3qt6AUc8reDGCMqJGaCl8w1HnU1B6zUVkCA92VwLfvE9Z7A1SPoAoQAEJE
4Z+caj0USaAu3z3MNqC+I3xOY9QHeBY4cnqYaJdKzc1hgeyPNsyuhQravf1DwtjSI4jLoYIg/vez
/czZmlLgcIKP+TW2rh+0Og2RYWF2eX68HNWadJ03UShK3TXsqoLLyGt5XH4NgzYMTilcgZW/+95O
R7EkfT+CrwONiul3Aq04V4qsyQHVGupD9OGuqpDCkcrkA10OFZ1N2xgHEuYoLDkf2iePR8J9hAGt
9dASGwsHEKE40DBJaeFzWMgx8pnkthZHZMSnaCTt7XhCEyA/+vF+JMO9oJHvekSLO6/AFd0ykZsk
MWswzhmrYvknQAmhXHPIqGZptGwUVHigw+T38FB8Pu/4Ias/C0DOTEdai6kZTFbT4/HDKm8fqh58
jC3XDh65iGLv2iQO4mHOc0KK+hBgJb+rYjS19z62QdOzSd0exYnbeEhM+0zvxMRhZ+B01H+lYV5p
ZgMF6Vt79aI+1f/Gm9TQkc1DKsAo2n2a/meuJ1mQ6XHiNtzcpNloeS9SC2OSd/66yWPI7B7bcZvb
zcBu4SxL0DVbeyruVtPzK8YL9XucEEe3vVoAZQQASdJP5022Iw0/ld1YFYUHHiRRWZUvhp/QKeYz
xiF6yxCOO9LVUbTWurvFuYN9SolBCDO1myv1oDfqkdcIWMOUNAqcSi9Xg2jQG3AHfazwxYVtNVkW
vu36GQ2MOg5Zh42510tpu8zmWJi++z0kDUKMFLdKQSHTGz2mLJ7JMJiuBvz/dJfAAsdpCbUkIsZk
bQX3QLfqIKEvweiA/M1iXHI4uzihMfnNlAeAhh5LslEFHFHNuKF+eR64uZIJSoI2Z0DFdfMVtjSd
1DBzNM1y9EAWFw/QJs/8G5CsDl/s8Xxi1ezY6Zp7Q2Uegizy46F9wObL0N3WKc4/mr5VklfwaW9v
CrK37TKaVc4/5KaVIdJDkGfTibYJnKARagr5hJDc6m3/QA7K2W8t2vMjjbXWdubuFMU5dURCFxeD
n69odbwjtpElvhhmTPOCiCmR5QcnErCAULWTJYktOkXFABFFVGVlGiQdr/SGAplFnXrjqFsWCclp
7+swZT3ZTze88d38Hc/GSgwD2ASQDm6hbF/HGzjRkCNJOElCjRSghFfijJUMc6CeffqabFeKd5EO
KAnJG49bdfJcmWkf8eKfVYREMZV2OnMgc83NmTQwLNs+Cde/DeZ9HvIEhCBkscpV/HRABuh/m24Z
cEPpZ4Nb/5eVqRtzOmDRRFWps/LgDKY1eTs0LtjQKjyuUbHhu8veM6NFpO6x/pBoqbezZlHU4cOO
Tgw4AHpgb9OtllDitvqdv3nszmRpjVNGKv8XkRVaIAFHe+7BlRmVDbWH+hNdrUCwrqrGXpvTrvUE
B3LU+pKMxDUJHKjjuU0V0dVjeSLvFF0rBVkj3MMV3ocyWtYPaOE022iYrvw4mtumop7V6PlMgnWk
oGUmS4i6t7LyzO2FmPvUqLF96Z/vPIIOZyo/D2oVroru0M7AFRhU0OsggqGlJpWXlRO5ixsNn0XY
rcq1kF123rSvD0GUddm5GQXS+EFXDz/pr/JmiIlsFoQATmqkRCCZMM6/C0tSo/Ol9YDeOPfoiRcN
ryX7qxmBygnGU1M0+VdMy8XB9vFKP2JwzbSxBtwg/2r9Bz2kDdrvhu7BRcSb4QuG7N6fCuhJ4g9m
N+lMYg4StzGydJGahrPrfR4ydMgB0VLMDE4KHVRPYaXQ60kihML01A2vpzFwp1RB8MPyidqtOMIA
V7YP41FGXnfu9IMgJ6xK6Yc8VVbpRiUmrfaxP63I+dymO5JH2j8dHVV1uIv95VoEJTXyHsvA/ai9
3Hyur99L20ZGYGkh4e14eZMGTzvCwop0SqSLH0phbGbtN3BkOJkScY18T5k5ZMHYLLbIUcBRvr6K
QyBK98FJOhSWlVZYJhMUa9pXHoAtcqGruSmSRWeiekRhuTM4qJNYU0dV/fW2TsphqiXCQFLKGaft
NdMaKI/X+fVMPQZadmTgnz1+H46IG1FJbtZMqGYvcNjC+LJS+Tclt+HrjtMqsj3R6bEe9JBLI5yY
wbSR/uRf5kD1CONY5DDHW843zH2PWRA7eY1drZrzZMTAIRlgscM9o+Zbpt3EQUpzSLP2RRsenD0/
AtqU4VvPD9c9pmxkkGMNu5CWwY0HAS8+eLgxBwe4Aw1DH0Klj0IsfAVEaRGRYT/BgZvWyKdP0a03
yGNnHCvDgzgioUPVgA/yeVhAPoNw6bz8JZU5FM/onJ6EzgKNsbkZQOu02B5+2pH5J1THYg7cy2ZE
51nWOGFxyuI4gr+B9/w8gh4eNgtTCWHzwvtzUc4D6F9xxIdVkeeCkpfIDgBIiBo9Tjktnwv9dzYQ
v3oeSWuExpPOz09Ob7uU8OE0EVjvgK8MDftxsZL+DuU8fSa2FCgzMZGTPLcKjou/62E5TC/s9a8q
7lkJh61P2Iv7+TYtGhHV8e32XZ9nBv3CIyILadq0tE89KYvNEqxtkPUkAv/TizLaTJB8uqVBVrXt
4ssfYHwkUZXBCxk+ihJ8JwG4x2iKJqHhf55bghmffssxLxFuqUJk3m6Xf+EPJ/LuIZdJwOsF8b5b
AflAKaQRzBNdZixQndSE2OSf1sNlMSeaw1aU/ds7cYF7WK847C9OGSFOKW7IbGw7BEKteG3PtzER
CK6itmjXP5B7rh63245ZOupuwi7QYrOel+SdVVMuzPpwgmcnqjtTLCoX8Kfyuidjsjq1x3RhG91R
OM1WQQD+LU0FBP43fxq4b/ZRCcXhGM+E89RCClJoZmQa8kKen7dvTWvDOTkqa9dmu3U/ve+bC7aH
tFVA76u6ZgrdHiL2Ni5JAzC2HNR4/yQl0jbrYfjU40w8at/yvoROC4RhR9UB44+nHegTnTWp+3Vs
BSfxm3G3kuu6fDjkFpBlaFe5jZ2ORsCq8SkkJ8lP4bRGKf4g+/G0OnhwXXCSe1B5Vq4D6gp7snjS
eh7DwuFBZipTlaY+e+wOBZ/wHtjzQdY4V3PWPFFmQY82bS8hfwOfa9dM+sFnPIWtw5gk1hweU0Et
YywhtYRFiBDog+qjhDrd9JBV+g0LzAOHlHyoAHfnDi2NsZp6Zho9R9StiLgD3mf8Q0stE3HUMix5
HwebNaVPY16XD70J0rBssab8eot7r0bUESCHFoHxzWKzA6sXFmyK/keJUcg0vRlqW9g2VbvdOGEg
CGpJvQMPEAX1p+c0BTzTCuYuG5aETB/aPnP3WKG64HWMqJWP+5ifP1AX6NblhHPKROv4refDoBeN
hDIDg96Tm+X3lCL20eTZPoTSrnVCu7uQiqJM8lhAULDmWsdGuOznQCi3W0T7fnJBX20UUrzaXES1
WR64yQa2dTphzGR2cibQP4JxBtgFLpqZSulyGk+5NxZhAd1qkf0NtDZz/y6ou5+mv3u488vaLOKv
qa6Bt58y/Su8VRtExOnMl3tTmDWHcI8f+/EdOgAWpe8pQtx1k3WmVlXikdiC/zr5ebedsTqHthyV
RYktZq1G/YaFTV5zCP92lECCSeQ9vI93oAh/5KIijWAvroxKDiJ5gdnFpVvOdcJ402HcNwGjL9BD
DAVO7pC88dYXM4ejuuBpCeeuRMRQ12OYKGMF9X8+52mJaPM0SWuV3V5op8qR0gBAV/PnUmPO3pWg
9vRphxS93kTTjuoZBQtHyyeJLIXcBRF4yBgv7E1t7cUia4Pe3683a9fBJY/GGxmeNXv9KlxzuN9c
5Iu3eHDlypvcwr3tZ7quV546KsAaIcQUt0Rutwmers5aVUF7e6ARS/sqa+oOXun7K29x+otiPA8A
gnj+D9AaYTc+iBb3Zu0cwTFGIv/NGdYRBiQzPxkvctt00/urD3tq13PSmoK6vyb63jrknaFaFmVU
eDqz2QaLonfW4IP0TV1UXmsjSK3bkGUya4L0xv9K28HKR4gZrgu/o/XpFPA9SPe+Xlqmd6t8c2v+
XyY71+POAbiXkqfMVl12/Wa3Q3xp6fGNVdcnp51f9yo/RoFH2ilf34BVDoQoGS3TrbmkusIgfUu5
Ss2WJB3IOkhWGhQ+QNIzcvizlCeSxaETJ5cKmQE2v36sJAlfqJEvIeNXSpX1UiMTzaM/DnB93Tkc
W55VNrlZo+u9JCQDnFTLTDuaasYfj9ftBMmILCYEg07R72WAHzqZX3Vsa7BJk9AuB8a21j87r8/f
33QV/P+4RuGiF40mLaLbARG/OXp1K3pQ24vGCcrsN9vNj//zbEb3rAp49Vg/rdR3lta8TgQqFE3b
GQCmkC9ffG7Ej/77mLRRcfEg4mmW4MSaWxHMGPJiBuJqTHLtWtzYnMpNxD8FukeBRtOsiL73krSA
pK+8XjC/0IIn2hLuehTtrS2YrShZrNvDu80Kn/UuKzEbp0x7nWKe7nBxT5pCkEJFKbcaNjyv74YT
58Hpd5n+6YciYwIfnBKKuITsha0znSarn4gE8e8wKCaO0eJkoTD/dQYZoPxG6dO40GX3b5fi+iS+
O+cZWkcbcOo2M1aVTEUcA82FF4VcaPKmA8ycCBW7jT5Udwgvho0vUenVmbuVVcrlJFCDsnpWi/uI
d31J1CFc8bZc81279eU5OwqNGdVWTEbHmGlOYZ7CNHXsgqSKCC6M25rKWzghH5JWDavoJ6XNIsam
p57Sc2Ic7L/i9PYPewVnxsP36Rt+kTNtbN/WAEBSbOQLwRPVEi7wiJPIFDly+CWj4tyn2zUKtaQP
ZUWp+Xb2lBJtg8fGGp2Ktgr7bvMqS3nqg3ovxRXKMDz8v09u4HcMWA+FxazNBOiWmGeLlVVJtsZg
wGgnc3ifXeK5H7zc5e/TtQOiNj7036KL8J/SzWNwYT0re97L7u3iaRnqSNzmkJ8lWs0BhovhSagM
guULN1bDgbCe5qvPIo763dcs+Xbb0/T30T1gxGDRBlyc3n5biXY+OkwG3Zvo6fCAzNcgsq6YrkNh
ewPI1pw7VL8B+U69q+DBXLIgayt1nxijgJ1u7dKUqrXY93MHLYkiPkH8r6rvNNV0VqZizilhfTNm
lYnDBlBxRINLmaZB8PIVYPYXob4kT4XDkAjnc3FKZxp1nijdZd8YUnR16qXSmODU1z8/gM0dKkds
tI4OewCqG4HAveHfmm+kpWxexDc9ZYmdloqHD9SN6IXpg4OBB6iuxaNUHBTbfC7U64mvnRkSbDTx
tKILUqpzBmJUjSOyWJtWGXQaDeZ5dGJlYtpFgdsuYFlJ7PWRXOMqx85b1eKXftnXYOcNarUXGcsr
6DdMRaTzpWYgFB3loMn/pX3oH0u2cE9XxxkiSCxR3ok7yfYBlwgdoicfNpUW5fd6h1opwilkVOSe
fRzaDwfabsFlQFyYcyHMIuGG29YGPAY7fOxKXtDAtpVEHPH079hr543t+zrTN7zTUmBTjDhzTYAi
QWqzZYo6gNCoVCV1yf0eFVtzOjkLUbplTszWPQxGyWyNCkGzMKqiuKkSOZTxnu7vcjOkAwIPTI8s
qGGoMZdgI1Is9V37sHL7ncFW+lircYG9eHF77S7Lo/Glz/vq9vGvgTmVnTDWUAfdPBP0g6NRhqvk
/scrGoBa0znNuGTJUWQS/B4uNrFdOwC+QTtSJ+KsXkwuS/o9uvnaqQ9erQthOahKu2fIoSNX7l9k
84oqu6GEE/AqTyhO2N9lCik+2xDSwC9MvQ==
`protect end_protected
