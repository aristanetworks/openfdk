--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
UNp4mfBYwJypGxSrCUuch2RvQ+PFA/qEd0RVAAkHgzpB5zPCAxZAuKtrrsIkyctVgnmULBQb80/r
l+P8Rk4aIWiaLb3h7YcNZBia8hodTMN3EucqLyJ4XwzxfSCng7DPSIVJ3WGJS03em99jAhvSfwhW
cBbi4WZy4Bu9jftUQ4OriMxxlIVrnKp/yPhi68XPa7q/tC6tugLgGNk5wwBbGeZ1q/NrtoLRO5WS
whKNwpj7Wn1L/cTrPFvqjhJKOOsTyeXkyc6G7i4atIUKvi8qlWGYTB+pYBEjZ7D/aWt+Yx4Rrrg8
ujbAq5ILaZuPnuqZLYbg8QDP8gWF2yb45KsWuQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="yiY2L2VwLKIUZCdmszXw1FNNG8F1UbEM6P1lkrvDO7c="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
kKa7UJlEFc7y/fTLwuOaouXofQwsd3ZrGB+dmO4I7wtCDkURH1YaAA/U90xKbZtM39wctNt+v2rf
jJb1MDN8/ZpmkXpcTWwIw1UbyJFknTj9KlvkizmpyJOxliIHrFYeSb1ZwWUFere1AlQ2sL1EXTlH
Gz/QvjX0JnH9GB+7O6NfWrHhpZf70cPbT3H9TSGiN9yAkZ/pWYfEUtRHne1wkl+DXbRZaA2DYLsv
NwC0aFsF/2cDPcGJFwVwDJCbjn1YKKF+OurIMH5BEWFIq/cowS/lPeUOYbGecCM2iyG1fzQSv4gv
xdcAXHl8+wDVCxM04iyqm+jyJGQ3smHdqUXLxw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="LhIMGWvUkGRO2xUuKbB2F6oortsZ08tvVDFLngSV1J8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2480)
`protect data_block
Ndnqwo+TcYQh6/G7ofrhmdq7nX6mADN1gPwHg4udBGI4YhBxsYBeaSnuMBHHri3E1r/wP2MSTz4n
lflCp8nY8tLAzqR8UZ/0cn6aRuXRfpXhw8Tt/S1/xyAq8Bsg/rolOqS0JGx1ObbgwjIDC9K0GYAb
bfEIOqWVC0TfHdP5hDDCtrdRFfFXbVMKboiYrM5ub3XH2QhF+q5A3tG5gtJzi6NhtPseYV8FBZfC
6tlxlz5gALg7QX7r+CGVSEitD6va2egrVGQED5+FA2DNnALxH9xzJSTWl16QlO+QBJPXndNkHb1V
lcA6QextHYsHzq1n3TAEizpw7X9j2I1+E7SIxXZMBPz/N9dDlO2sMZSh/VEv0hJOGKMSCB730GIL
5/LjqDQ4/pWlFmrnEjaDBt4obNoRUodxE24d3po3/QHQvYhK9L0aP+O/oW6OM2VFntneWQ1jTUZ5
BzkzTTjSV7zMA8JKhk+YyaL2cohy6wU8lP1VlzGUbo1p9VD4JluREmbwAx1lhlucccXa4asHob7m
Z2aL+qwH1YzBqlp/oqkW3fBgoOIG/XFKrst6+QHzLHJnF4OAV4kc8V5SpEIn2WM/xPTOHCh/hYdS
H+MJHaTZt/wa9xIpMtWh6T2KX3D/IKoc3gjKV4iqDF637+U70QTrQUeKqQ/aOkLWKSxAOCXDusMG
vKEgWWXYI6avAnaR7zbBI0gsQ7gtwiJq9nRKXpVmeEEhugjdJMH3wEFWcokT+x9nbBBGqNwGtl+K
aWFKVzHkxN9jm2SBK0kLaenCt2P+kQXLbJGzZocsZT+Dee0BQjfWDOkBtS0nX/E89YWEcKc9qtJq
ndyv2SU90cgv3qGEf+8/qfyUPke6cv48T2mmuvxNjq8RU+yrUtgJ1mvW1N195jmSxX26mf1HLGoM
c2kuffYH89ANGKvfxXkBgYlNsAx3IvDgkdyv3pztwmfC8uoks2Ode1no6UyOmskwCuPgfsMwFNlP
f5s6no2oileL3YDgicoA5KmVyo40oP0WFsNF+3owJHOFXdVnWn0lJB511uxMN71gzeJWQdda+Vjl
sJMjXIuV5dso2cKVr7ne5w8vH7E2xHqEce/OXgFis3TAA+naZjwOpXdwHO4tT6Td70uzg9eumUdu
K2USP0rkVADRENLO87X+jMtMJ1IOPuNtfI9L4DtQLA62e0AfPnX71wMagX0S+Lb6r/7PaxYW/e0Q
HRcEpuJ5ewHC5L0V+jBuh7/YgWdES+qcZvm1o568IfjWsmI3CVPKa6OX+Vs6K5pSQiKtVYntAs+e
gSxOs69atxrtMmMidqHgWOLSHJjBLAM4ppRfYBss4dU+Qe8BniQdNMmDpwnPbuiOPrOm78fUjiqK
EWPr0zYbwFtJoDhI4OveUbwtj10SyvWKlbtUenJlp5KNjp7Bip0A9nczw3uyPMXjDVT/8DmF9KB6
U3BVak43w+DrzJ99LqjefIxGs4MyJH332L3DuWlvG72YV/FLKiUzhh/uoYa+I6tBXVLGFkQAvei1
LBEX0ix+y/XXZtIas/FtS4mhyayrRLcCNiLFstSw9dIw9npOGdI8K3/EdjRbCv9D//HB5ptCgi5Q
0Relnr7a2FiR56ruzU04ojTw+7x4JNeB5YpK5sM7b6Jl+7Fjsl1SHDRsYJkGZpQzWXixJGncq1fb
lfTFGsDEBQKfKrxXDEUIrecUNp1xaRvBQx+wWa5UutUFkugZZQ3qiW/c6ZKE6O1T6MULHd+/0I/O
2NEpc2dKtx3sGUSVMY+Wybfu64M/V/Eb75tk17Y5uPsnCc7wSMvrpnRUaFv3YHmarPILhEfcknXQ
b8i/sRJnD0maVcLe/nUqfV+O0k2LnhI90P8hMCWjHCiKQ+jNJKI1PFSENFAZsuIIJGcsNrD46oc4
+rAyTuNkLv5pX2/Ky/PhbAVwVu6JMmzYl9C+LeOa/EysbOF3deN778QPN498TGFOq/iisx/hkdG5
JistbpCQ0PLozIX9g7hv/YmOH1aPNU1eSk7VxmEh+HhHfQ0XMq5jSUUE1uYi+H5JifokBiv7t6C6
VurrY7Id9oRGBuBxXLnfGF7Ukl99llfSdpYGfvpyM+4FNdqpNVPvrZywquxqnR6at/DgutuCUeO4
7YeXWFPJnFUUu1ag5iybR6Wmrm0qoKjtdOKMTeMGjntGktMJmYgCf/os1fvrnw8UVIed5/hyB8E2
NTp0qPBsyGgjtbucxGZotx5ZaXNv9vMwSqdomO6Hp17l7E9g7dTMKF9b30twpf45P10X5jLfzEdq
09h3M/GO86h1zYnDcLBfl5RG19mtUkz+ntVQ0/wH2+WaYLaRMo5JWA8IBUwZNNNa2EBEet+SVO2V
BDZPmuhFi2IzerGlnwvjlRdZpiCXSBZQi1ccpbqT+u7+7lkSSMGC9/yQUyViXkFXEV/PBucw7TYi
TFtLuCImMjY8lkpkDeoKowlVHUFodiAFmCjs6KVqrhjM0KzwAMXNAEjpAt0tWkgOFHbilNw05J63
dA8C9zPCitXRTUty0Ptr8tpCKqmI6D1DqW3ws5eAwcW+ENNUmT6Qepmy1B3Dnhwb+yZi0H9bkGmk
wswljqaVfXlimG+du9uZGA3RbVNccvJo53noD844waj+v9DSx28CLorkgRSH3oxdBizidx88SXFo
95+VNF/uF14MOAwpmiGBgwGez1s1HE9TGsEhOPud3z+osdcRDtU5huB/hGcyorBaYmSz4HuHAHn0
wlv94rmxhbY4YOE2NzajtzrJ6sH0JKH+ivhXjDMtuAl3ZK3q0Oq6K+q1eIuCyj5StpSOx4DhpNZ3
Z3+ErWdbQFmhMJJA72Xa/KvHd9tMio3VA4tci8YrK0fl9pZ9w7ksJzZ4daOzjHgHAklXsjhk0sPQ
tCpQNCvp6WvKEcVS5dx6nydSzxCDAOo2xEObAJzigO9BSduqPZeVkqkb5v9qFzENBDvyGHgbx7RI
wtwnXRH7pGxXQvH2ptWbzl5fcYov0Cvi0fOB3UyfmlqILCq3uhZSPhSJyQeU7xukYkg9OkFEWhGT
D402PrgMc3SYpgSNqCEUfOunC/No1Wfh0+639ls6Ke9vzQHiTcG8qEh/CdolF0KRSgYa2pYQ7HPj
jQGwkGdvoYRs7Tjztp8fMbKn+2LuQnVp8jX8NHd+i1AAKlQzbv9f8LBMQFH1HJVla5yG9DMBIHpb
1/JGNUcX/OMP0u4x7yUE64qAnLHBUCoxQz9ANWoNuxqlYINgitlQnE6At0u8RLPdnJIxQ7CgrZ4w
JQspxmqOd4uA5UT4Y3yloYBNB/BHeZnmmt3JM6I=
`protect end_protected
