--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
H6fddWPUGsfO8rYPt4Vle0Tm5g7nWw+BReLCbPGYVNMJcY0GkJRRVIAkj02ykKgWTVgShByWEHwz
ovkR1RUt8FgexrMe2iiEGPmnCEjRULxa88Pj7dI3WkOROdVbh5ktTzS9BgUiGFLPr0X+45PoBGf0
PtgBnvo737PVo3eGj9KjCQBjIScIPwKRqA3YRyhICF3k+9mO1wIx5JzT39o3sor2N+0hJIdh656l
IRnmaRZYpNO68W1Lkr1uBs+LUXfVoM0caMvad0qOa6AU0KTIPg0FctpSQTsUutTGuW5CAYR3uUwV
yp5nMuMbPTMPiLrAR/bITxP21LxliGdJbi8VIQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="iO3270o+exrcKTurKUcaIXmNlwA8HGZoffZc+gEVbcA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
SXP0kBpw5itKbVqyMtseCiyFYVfVJP575nd8Nh+WWxmoJUSLlT6OSF7Kq0lRxMlPSXBkCp9PAUUT
4foPqr5q8mEzUrav7HddJEGAFwoTYXhsyZveXlga5ffqcdjqgQb+Z11eP11z+nm9kABhcv79SHHf
FsIuNkvDV/Pj8283NUU1dxMVRPQ1NUU8/v81+JMz+DLB4XUBKphmuI98nEKgU/UsVWr3NbL9Yfgs
bthokXAysnV0Z/j1N+CN4pnY2ndCK+EeZZN9OijEEZ8hTlcmPvaDPyPzyBILbPrUXefLXejUeiqV
PMVT31ATQLr/j5gXdmxZ47DyfAWG4o+pXtD3qA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="XO854qqilSEfjRkGjq3zOf0U04mxxcnbJdxHBmTrUMM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3888)
`protect data_block
JbuMVFFEy0PLKEJgVHAxw4qKkdWsgbj1/dNzrSJel0SPEP5c5+YsSP+aGfm2BQsU09+H/YAypBDD
3Rm26RC9QJYWUcE6MsSboLRyEI0mlLuObeJD0tlxu+cobIc6AucGcx3tu+CLmaSiNo4NHm1wo869
H+tE/+n/xRoLLYZ8v5jKpdsWi+iqZYliDamLa0hOqaoXmjIqIqOiqIIFlo4EskIGH6l6tAMe5eTb
RjEfDBuaSSqW+5r/+EMVY2E7ZgBF02DDXDHutDfvAZzlY1ksg9YefkY9qc0COhl97npfbL+lxg6+
jz+HbmCYKP9aJWfAwY8jN0vpBBSQ0SgwXqbVHT5qWvwkILwXrw8q7yicUB7GUryRifr4MiPhIr8y
yGgqHpYZ8sMrCkIErElr8pTzzVp7Us2lPXkNXc63aPOL5BlkuoXed+/JRQoi5UGbOepYKpVfwyER
8PaWyx5TbfTCcbSk7eEZ6C56UGYHVTQnrN/Yr8HKrC4d6rFZlwCRzLNVKME9k2LU+CnGmqWkYYw+
1Asz7G/CZSR3k69F6x8CwZeTPLrcivDtrwur0DwgXADjlKyMbMf31r6+f5tjBbF6VB/9KIJ3O3ji
JN5vNGTkMlm043tzzXITwFGs9A6qdtRW4DnM0/FRO4v+MwVfIxjYEHRvxtMzSHj4WFt7j77Rm4jj
Nvjxywuw5IFUpEUg2gOVqlwxIsmowR6l3Kwbj/GGKseT5LD9Xu7hxCXLD+zqcgtMiQzTgy6IJU2w
v8YHC1YmuEFhp1+vtzQBN4ifDNEIWO3S0pDbC05dyhLwMrGxjYYzi5YAh7P+cTtVuHkBDss0haIc
29xQ4fWu6KmlbILZr9t8ZxOIVxAs6Rq0AikbvMiweF0QUSawNIFJ2UFvaGjOmq/EC4RwZUlVCjWu
8h3ZbWWKW9shjxW28QsC7s4koQVGgDxbKwlgVgtj29r8hdZj2Oiot0chAKxlYllHjTbgmUNBhMV4
fKsPl5FJaaVh3+eCGG2LnX2M3vugd492Mw5USM2LZf6pSEeoJP0AfPWM+fgB5ouUWs+xf2N7i8kk
6bzEIHCRhFWORZZkz7Vi/ryFt7tURVxkZodiy0VmG5GZMeNs3zBRm4OCCIk+el6W5112LPkLGnKR
LrXtV6MTsoqhYUmx2mlVqRAE4/lzUia247Qo+Jw7XahUwBj22kGabew1GW3tAvPaEKLgV5CTHWIW
gOHYh9tvZo8uK5c4AkUNxkk/g8pwExBj11rCCa4X6A7wxmS+hCzDhAcrPiB7sfJoYvk2Is+E2oCz
UdwNoLJMSxzL85u01Z8PVqdrqJ6XuOIf1jZl66l+um1HjzcinKMxMrafZvVikPxaRDohM7ae/2Rm
4awsUoBQQXt7gMU+8x8MJpA5muCGnyxGNpYdfgq4Eg+u7wic9TVV3mIDj/khuhiQsz534pMeZ5NV
X4g5JVb5JIXXhs2+vNjyT47fK9zQ78HECC/Lu3mehzyswG0CXEDvxmFR7lbmKOZEGkCoZcoXm9ab
/1anvIIbCIeKNB0WTJoiUxNcqn+ByTUYE/fn02hJICKa4WN2pWlyF7eXEUNbJfuTn7UxZ8/JkReA
xwjSJz6zZGjnhtINsSmOu+G/gGp4/EeNvHcGvkpMRW6d39ZyX0ipF5fVLzgWMJfIbR0JQ1TC5Jxo
jgDoJJRLZ7Yy1/sG+He8CwxgZI1EJ3580Xi/oUXqI7XgxuBMIttWy2EzJc/DMCyw0wibtVQv9XpS
EAUbZJiuCtO+UaVXI0FPXcXv3C8EF6AcxsUqMGIYM8t6myndALqXA584ELkbmWyaiP/KrBnQD4hj
PmiYKxgyC/b2AEwSSZXzA3dpv3zNKgBG11in0uN6JXJDXes0HJbXX4oCTPZ2YMOmkwxra0rYnZ/l
72u+HXa6HLYdakWQuJPuRvUQ0M6RElE6Yq7P3fquK4I+kIjeiDXesJZpIA/YsfcfZKVX6sdojNZK
Y0lG75ie2yf9hjrUVwR/Gio1Yq3BwwLaGLEpTxKDlJ/bY5Uzd9q85qjloAVoNNDkgn65BAuxOyUB
hbJY/O0eHg7vgpwLsw6RGZTNQ3eGMk1A2SR9GFLcp1Lew4YnSSaFlNZk/hhNMEmr4Lb+Skjr74k0
TvlsX6K5o98z9j1qfb/e7cW672TGJ48H12Im8Y/hq7ISOavy0W41jQeCUy5vfEsg1DaWQ2u/FTtf
3S4WLXOtL653IuRumTWo00Kaz1/eLQxscahXk52AxMUH+yNt7FR355Z3Z4MPE64dDhgNGHAzjm/E
QEws7Sf9oSFu9Fgm9XAWjzBgoVfccDkLfQU2vb7jkRYUZOzbmIbA7XKgLBqJwK69MbYXEX0ORlMq
D9hATgcX4DCjW8KoVbw19zeyEDQNoKaoBQwb5pPv07vTW0n+QgxGiIVNP03R9LMhvRW06YyCllYR
zSrhwuvWG6A0vjqzyYEeWKrTLkHybxZk8qL9cOQmo+VR7SPiu1Djolt/MEXUDNNA7BUs3m5zF1tC
ql+0iSSZj1usu9ERZSjtSsUFeXGromVdeTqav3kuEYtTvaZvhlZbkX2uLAt5Dsj7S+WFLW/im9Mi
rPBmEp0OviKFHIPf2deOWaQEipPxIcQ8bOs6kN0QCBYwTt+8NwuQg37kfERjW7wNiPX6ttqBaMMh
Fglqgq8D3mvmyJntKsl1aRjnzMkKZpaS5aB1HrBplJSBU2scL2bx+JT1ZEPFUmw5tfcI0HHHuY3O
qDMEjo32aImsFuPK8sWixfEr7K6QSg9zznBrtcrf4hYkWax/Vv1IfppBhTto5j3i+1AbRwLpX/j1
KmNDmrv4Fhph1i1VPjCEo9WEzrmrj3JCjPE69IuMwVtfSR3CO0haz3oxdzjwl/YnPKWqXKgjntpA
j1HyRgtBcW79IRMp5znK/1piLZxn6aizwx01R3Ay+FrMKnQkcARiKy6yU61zIc8uq2S/rA97Tc5H
YX44iFM23Vho0EPxMBM2MegbkvSFJqH5SdoooTQMVVsbmyeqS1d1oki08ZLu+vl6UuTstuTwazZ9
c2rbhgDkOODwA+YZyTihB42aLrZKyxqp6mxRB476SrW6IpdCXhbsx55vEboYHVvv2UH37BDHRmDa
HZcWHWfQy2xhdsrEcWzRZ20nEST7JKmq/2MKW9dy/B5ozlTmVkRaYD7iNEuSLiMuyktYINhGt4sA
pFUK1nWu47UZCkxZd4D1x1H8wQE1CLCi8ortBJaofxtwA196YFr++HQyzqfPlsyBThDk2L3Ir7aV
Dqkih+ijW+bvUi7XaR0T+Uqn3NbQRSzYkdXB7SvE3B2bh6lE0Yl/TUoYFbk6sfJW0yceR8e5kdsx
nA/q/HD/gxcb3XQJWHwon6nrYgW758XDAv9YVkO2s2adttY9imD54zA9dR8FpUGQrVdX0stcWANp
1B4oSSGdrSdfxV8KItpzJkuL6abbJfZtecG3e0rHIk2J6NujfnSb3ueLTiyEBpkBnOg0kIKn9Uqq
lbCRr0MJPhwSd5zjRfZOdIWg5ImKTwr+SnJHE+Hqu1skgq9S2zqFdRLK2go1Ib7PSsFib+DjGsPp
HjRDRaBD5bnSWUVrRn6K/0QbqRCrvdM0BtdyX2bJHzjIkCriRtO20IbM5DbbKkQCoG0VkepRI+Mr
I9tFB4xToc4SUt/vqLHpYjQRGCvH/PIbYdIPrIlYBKpHU2dE18l1Rs10AjjpOZ6VT/CNb9ZLHtJQ
poByanKz7tQ7ccR2l1mcX4I64dhzRGrYRe7ejWv2uoTTOetSmF3JT4g1YHYr3biDbmZkRPZXIObj
XLv1FNjturDCnuCJ694PtOev87t+6RaVI9ZNjdnlwzoY2r7jiwfmIRrxQgUrpN1tqiuTo70Al5QF
LRFyDFLWYzCSWTfchXmaVgqidbcJweulaXP/MUvE/QpncX9nBF9itnP7uQaxXkZdbVVfuwV6CrdO
DmZ2E/5HU3QrZDhTukBdqAdDxGkgo9492C2q/GaAIZDzfXR+/gaU3JLlDnirT1yeZP5IByhkpspE
u/KkW7BT4+kOlcPIjvvb8A63/pVWVaYpOBhCJQZVpwzlCY11Yd7sznYI3axUMs7Kp5ECxGIIshz6
Cvsj46a1GARJHPm8CbSmdiKXxEML2zUbEaX00hgnhX1RCLIuk8yKasiyIdI7PcCoYv02rMC6DfnP
X0lAiswbh4FxXWmIR0Bn7ORLVjCBX5x5HN0h+eEpVqsfGvECm4ubo6JBlsoiLGe2hg2+eFca/wux
Xm/mHn/W4VlFxb+K56TAXNW78iA4R9391FhLoUUNv1dmf1zzUYOOJDywnuXVlN9s+Qn7O28BquBg
VoEamUqKwkMpS12Jv2XiPOhEOOhUotLHgsJlPW7YLAri3ioGYe+ZMEDROyDGI9+kHkS8dokkXlok
h9yuOPxVa0WCrG2ESontwazzjE2c21Ywxk0+t+EA6BBo0QhjLfDvc2XcrO27CzOk42DOrnLp58+H
zdnOrsjXgF1euImzCU5QdKISvcD+ukrf7rGKPn4VjWTpH/1XBKryKzdrK5bhKdDrvG5RfIGS3j6a
3nxFMdcECTzHAgDizAzAB4g8mHtuIDfm0LIz/fv3iICHeFnQ0BHnhjvGEn+XE21xVDQr//P/vWaM
spalk3XC5K52OSlSON/kqUtXMldy7uANe0BcRFJHYPOITTVIpUT7vJFruP6mXL7g0dTCU0v499vf
eKxObRx3KuolMYuTlgGR9J9VND/8sntvFh0wGBU0w83WMTm6QmiupN6vpFm/FI+ah7WPpdX60HCn
M8HP3gjPQGdFzV6UeKcohQ7II9OYktgRQdDBebaqlyF0MZbExf2MZuvaoQr2j/k0owxBKJnfXtny
VXaAnUUBETQtTM9jOn8/BeoSaP4nMaoPz8hpZzkDWLgqrCnYgdpgrMxMjbpbv0RVhyuv6G8noadn
Ukeo6NirAob0b1saFkaDt8hvJUtiDUnDOAaBOGi0u4SEucy9T/b1ZT70uiddrjGPw8hBItFIanfZ
Bv3Jx4imW3oG+hsWeH1GTTq8fddKFw66i3do84qLbCAbVgl8F9a/yJyjF+kSUKC5Ct4AQZKYybtP
fXeeiSR8lcjl0M8hJOpZigV+PTg3dz5d7/ANUKbySQj4W0/EpCCPkrWOfDtk1OWAkeXc8eip58zc
jaewbtxiiae1aqMg
`protect end_protected
