--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
USX6b7k0AbY1v9dQ+gc1bxUupfeGTWVIS4aflSGVqkeNtzWpWvV1uy+n/20/LUh8dChSDaybyBI3
hwcQJqQ0wKeCr+hE8avOR3/ouNG/bTfCuiDT8ZPsl/hguDwqQszsEcBsN0vwJ7VjMs0L7qvolIkD
sOomNkv/gEN6rWLqC+w5cVQ6o/UsmL7Ve+gSLtiRXHdYhy0v6M64+DnSDVm7uu9M6YtkB17kGwVo
cENfInQbeECG+Q00kKbBF8xOgm87kN9yP2LZuDzt68Nxjis9v5jXmh+tFUD/RLm6lIR3DEyjHU8M
plzeCnMvXfhO6YiJgf/LwGKZjtbxor9w/pogdg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="0l6q7haBJDseehTXP7QmmUm29me7Y2jd8RFXcs4LVfY="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
UvPdFG7QZEaOcdxqPH7PpNFxv6PMC2lktDuyjNTM6+CSauYMqgEmzMeuTmqrIPtGppu3tV6bDYfF
PsOVrmMEdVJYVCFUhb4TInqDpKgyLiKkNeG07XrKZ93EAYTqwoqR8tIIyno/CnZVearFhMVOjS3r
3vrYFD84JOl3SDsxglgU5Gd8f7jqKJSK6vCxoM8UKKf8UuU5kTH5FrQo8JLqBPdg+WjMisgzdoZp
aKpeWOoQNu7oVrlacYezaYC6s4QWDwx0L8lBkKe1KeuKfm/EmFbQnnA9txCXb0tBIZT1TyRb2APE
xF7dCZbv55Xqwh5ILOvTrdwT79AEqN9zjUVXbQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="84GFuA9UhsdlKy5qOwxtqTjzpRU5Yc790/0v2ocf8JY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3888)
`protect data_block
CSHXR5Pisxh8dCreI4mVobEApsOn1CIJKIfOp8MglcPqsJ3d9zxTEci6cskb+AI9ZwV06amOR208
XKBIPQxHR0OpqR4LI5YYBrxHyi8/UZP+k8OnOAC2BFgcudKLeqQUY9UuRb1RX3znSd0Cw8BMdhXo
hoXnJLfu/1OtttEoZuOyKaNwyVWI9hMPN3cL3b2RaZN91vAcu2d7uw7SQ8j+dLDJ3CwtagEYM35d
ypzx4LKaeTX3Qi+jMHcYHr5ZmLt6HlV3/J4WIu888QfmPX9vS1vY18Mp3b6oCHvKyhwA3mEe3TVI
GuHSu9LFF0uepWfYFL1MF4g4MtAa5IXNriV8HMD6o8oSkKb+q2JUk5124DIVcxGlaEAJ3lICNNJQ
gkZxlswBn3uWNj44vZAR3x8up/OWrryRkgKLhPpXtaVa72LdFk8PvYYSq1LnEJgmeZFu4RWPdQJV
i4lONNLNEJFpd5kFjSXxPzPOwxta5UZlazBZbpemCasj2YHUx00uyiUNTyTFAEpPdy6vs1yhtxx5
qKD4HStiQbjG2p3Nr7iykP6gyiBn5tbv77uPwPREPAOLSO8rwIDeKd/82BwE7ecB1XsRPTFRHn6G
fhFs0NlUCB4ltnYFGxd0/toEpkyWyFFlkFXDcSSX2/I6FDmk4m5Fq/QwB8aUHkZ8YbJmXeYzIvT7
CZk077/cZZyBa0snTa4SpPGKwDv9jTVpvVoMRNo46xnwLhCFZ3LywF78Z0fXwW6LNFA9fExu8h08
lnThJTY+xnozsyqoT3uYcvDLndD27hmkbO+8a8HDMuZjqoQr7N512kl59UkDzv+M0Robe/G5QJA8
G0FYYhwx30omyyEj9AHRr7iMmPo6YwR3XjFZG3EoUnqIYfhMD7jdpp6lfui5VPDpTHFcZPHJ+Wy6
AhEmZ8vMpj8HSadO0AQHVwc39RWzd0aNGFNB75yIB5IMQ7puKiWk237qiQ72kgtynRKGFPLcA5ON
MS7AsL2GGmLqfbyIbA3UhJ0swpHZ/zae8AHwjMHRKikYVolSFAH5dNZfbF7/zJFdWMg7H/G/2SEX
p5ZMmI5EY4juw7XTWR0smb8qdlwy/rvobHnHdX6IZCkt4+z7B1tLzo+qXVPFJz3FnIE4dEX2Gvo3
RocK+/jkieYl7QMfDhRsgoDH2UmcuLMAHD/3Y7zcrhsdgzdtiNcjtQTq4z2ZzBmvfTA22CjwcsnS
S/F1lL1IIOm7TeFNX0qnK9CU2LFQELlVuhcupR4H1mvHbujPy/jgTPZ0tVlRQsEQScdTCNM1DPGS
UXfqsaZScD6L/ZiyT30+Td1zztk7CHs3yjjFR0BMT5qkhFarKVXqe/eP4GIj+rw3nCKofLVCCwRo
/vCPyLuG6Jiwmryd2DOlA4oziuccYZxSotjNwkNni6zl6wG6zdBokOyFggggbPo0g+WVXqsQrHA8
MY+oi+WoA6xk5AsiXeum4Y3L4X5XXQ/A/qcoC1TSqNQBbh8voK1k2PVlDpbdSJoRcrJ90v3TrDns
jxf3GhVGkLMnteyAkqCZVyN1pDN6+Opnaer1HBEqCfHqyeJhD1mFlkXOuZKzX8kzKi8Fjr4lrGDz
+80f4hwGx64n+rYW94PmbNp8AOorBTug68GTQxffW3mMFydt93mHs+axME4OrreuFHN8YmEIuUQ6
aKj7RP8g49ylxeLgK97RLo6koRMqoXcfcD+0EN3csfanHLF672Hfub0qITCvoCwVUJJafLgTFmrc
/OTahT5H8TD/DOGXdbnlUQS1jLXDmgKkB4LUa3u1Xf4//rWkfsB+hw5DEi5+jMD6NeupSk0s9uch
w1Wble7lYifecxidKgxKoDTc7r2cZAjhIpt3aqBuOBeqwGaVE9BFfuU/LOp2k8SUMUmbXiyOBXH0
erXfC94JTXoBbMLRxSeefIcSX+DdF2/kWXMKjCgLKESQoyyZj99RF+OHxC+D5/h+/4Oi6noXtllh
uFPg8uX1LxJg32742GVDLeP2IEPQn5HDkjNgH1LKot21S1NH3KBltPjKrCAV1k0jDtaw8ZtPyTYM
nNnF3tqAuaMOpFlfTNbIwdTeds8LS0an+/ukzq+PBZmxDiHHL57UqOLMpJ6GkCubSNefKjKdiaLJ
b1h0Fe3czfPuL7t6y3gf+PVNSeLVjlfU3m9ONUNfZXhL9J7PPaqHQNNyAovqnbI9g2kjz6QdHcS9
Yv3//HYWsNB328EnlYjO0KEbYl/3mRsa1niACZ/v4z8N2bIqBG9VhAAOyN9adXpHScCCo6udKeLY
/bP6tPv1ZPyf5h8cohVEWI07BrDG6nM4kKQL/O6cPDmtUJBqNax6tMmOPtk1gPrQPWPPmyfs11Hy
3nJWY9jnJt1omNVroPlBnp/Hi+SOdBnWHR/6Xs/3JYh5NVeahRbOUr48DJuTJlhz5hct0djNGGx3
1LHLXvo/ho0cl4Tnyvn4rsnrs1ArIyD3RAHiQa0dKn1vc3/gdCCc5fHoyUd/W0W4eWXxFVeb1VWe
NRN69S606NpfI9TSQ1yFnDaICW1QH1X5CXlEb0L5Pk7yUQ2tzxo4jJjSPDZFPIbYtmpPiaWgO0jA
YdTnOQbGu9Xvj2nSiE/AGws8px7NqlPNqoI4xK/vyI5Fa2Df4s2ZhAfl1aI8NxXFL5L9NhjJ0XqW
G2kwWbO32xEhOveMNhheb+FzS3hYmG5YkzeHmCOjYKN8EcB2gkGRFVzRZ7hTR/5ELEAULzCD4Sb5
FZJ8JMr2CGcBWthNbgFMxhx7LhmmVHGzY73Uv7A2/9PLgxg8XKrY8JPIEb+CvrUIhlyknXbgkhlf
pKIBjyfa9AAC+kWLFjWNHR2MY0+DeBKUEYrGzMRdlAmRM0JJHQXjYD+ee5pLPH6TYXyzdcuRb1jO
ozZvzRLDTw9NVimfkUr3m6PK6DufrQeUWSPU595+F1/LXLUlwSkthf138kW446zKjjf+W1MJNaIB
skI7nkx5mzBYJqL6NTcbs/zrkirPTrAzmQH39GBqgdZU69TJEFawpWZ7WOlNNN3ShziRVtao8TVp
K7etLFenpRc0fPR3I9eRgPtXKkRUqx6JmOzJwPgZSw7QFBKGNXHtdyYvobnAPb+OHATWR2BdVpF7
Aobl3qqibfJsCzS4d18FCIaTXxpa0DzrihW05GeH6bLZSlVAzOVjcfT9sp2SDqMR+CWDT4Si/tQT
NRWhzVyYK6XY8SvNnjOelRtZdk0HH8Vixtwtzt/VsvkCS7nV1vEqjHaicqxLinF2W2rpCnsq8vCf
40Iu2ib8KflZi1KhbQw+VQR+aRZozc0I+jqW0Kelv0zvRHU7qYCP3JbgxsLICUROxhTzjLoHkWMO
QuqNesBBXXIZxkgliXztsyBfsUdZGmqzzvkVe2GlNKO46KGWo2qt7usLHZkRm1S97QzDL9QNigV9
vqU5FSXNb2eApxX9u+QvL4CQ8nvSUv28yiIU2HOCSNO4sYn94++PpUE7Pap/MjvX76gX8tej1p+z
xFKrjzOdTzptA3g4KQMDm4hHaARAVDJH4vGFZAkDn5aP+i9IGhA9fAo2usS+O5TXFdMHCwHaK4NE
315a92ZrxXBrstkyYHBr7Uy7LiudrKXTuVUzJn3L55XqNp+fp1ff0yAqJYgnKdbRPVQHTZZoU0OQ
Dgg2tAp8mDi2ij0T4UsRxb2r+fRDbr/vP3yGYRXXSAlAKLyBKT2inH8A/fc5YrLsFsflqoh+YuCn
/MJmQNhBGJuspG5YFP6q7aOsFvMlyy85rmylRVgOO0WDDBzDHqCY10xEQD2+AqAbcm2ICr7i6wHL
XhK0f8MxUOCpp09GsyK3b5ktdpngsupRG0QDbD0dfcxRCwafdbb0aLc5M10iSVgHvW07eT5rGZSF
XkHufDOgClNvJrq4jzmMY66HWK3cbE6np/n+nLQ2cbq4GGB+foupEFs3YJqyMMgUf+6qIEFag4bD
5UjNMStP6i3HafhhdWLpmPso59dKLBU2qmlKA4gpQTCYN/eG+//2dH6MJ6gkwKTwDY1aLBqHy686
QHDiN+S2Cpj8EdagfXDsy73PAmcWELrTTfAIufgDl91DKc7H2ErXNDFePXBFePzdkBm7RnieSZiK
UOHbuyrKfASP6SWajn1qsC1g507x/O22xBwmJWGsso4RohM5dRoL0Mhu5TOBnRPMoa6fivpmsRxg
fzBCLxXQ2caBw9+aoxZTmsHDQbKw2TC4FiAxs2D26efCh3ePeYuXMiVk33jwfHICKyTFdG/26goL
mj76FsBadxh+oBjCcnpB7SuPqx8Yr5AAqzC9XUwZ3sdGixTmnLXYFn6k2qQ+miuAWF8mBA/mrsgG
UdVvbUOOakzTU2JRo5tuub4ufQ0s54r2aVzYDe0x36veglHjnO4Tw5Dgpm/rgHqrnTVBsrY3Y+uR
CtS+D6gdlPBsTGXSP7vCZsxdsqRBmV3p8nTyUNliJJ4jmyhdqfg6YCPw30QTu3LU3xLyiWlxoD/W
gSAsIICmQyCVXMZzb9/8KEzWcdmkv/TQW8VkbF+8wM1RM3vUGPLI5It9L3rrfLadhciQ/6OMooi/
YX9Wjqy4KCpJkFNXjnLZT1QmDEkKHTwG/1ZAozCpPpVVidSWmLojDjYJJlL1hMx/y20PYd1rCauq
Cr250UOV58irtY9F3pHW90mSvJGM6ukN/WzstSULUS8sxDqFFLskLH70uM23agceAiMesYOJVLDn
wDlJv9ycbvPsL0U5MxPxR+QH+HwqG+9ZHxjuPsViURdgZjaIrzrCNotPoHZpmwy49Bb1M/Z5Bbpk
rGEJ+dcrtgEjoLwhTrq9y3F/c1TIDriInIoFhfBHLQQ6LFxTaAINBRxTqlYI1dn4dHgImK/8UEEq
wMGvPmQwaYuimmFjgH5gaAk5WI5QYQ3BFkIqOOtOEI319LvUfYpU0JGkt3RduXN19aOn58H9ZGUK
qMzpo1ZtWWb1zyu+mKbsLVxVkytdqB+2uy0pcDbY7K+3s9BEOEX5RW3LGfKeXuCgfkpydgVi4kvh
vylbABO3JsnR/+5EgI0rWjn6uOtirxNXZOYltsPLxo920fh8gaWSNxJsuXLWH3Y4YUn4FVlmLbz8
H/hjjwuj55WzAbvN9daFx7shqrzIQtmEahzqpUjYNJPnkXtbZtW+y9dFvHIlsczrwoj4sCTKDE05
9tdQdIsxYF2I0W/G
`protect end_protected
