--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
bS6Cn5GEHHirFiMtT0IgrmiyqNne6UDB/UepC+DzwBYtRTctK9YsqJ5qRwInsni1TNyif+0c7CaA
O/rXxvt11gUg2xN3ZbzVPA7mOWp+Q+XPkLBpt0O6p18IKlcrwCYgLTxNN4zhl6x9J8phoicHPevL
HlHC52vqPkCbcwuWGfNey4e8wD5RTG/AnWjthjZMx++pqSetpWOBCP61Nk9Dlf2RVXiuok3IUZOM
eo6j4NqMiPD0ZH2Pyts5dqmM/bsUOW1mUlpXwyFWUcSUZo4raJ0dbOAyEXxtm6MLgcjbv7436Ubc
VaIdI+3i/E3aFEbZFaklVvs3GPRl6uqBF6iTPg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="h9fqTjZ8pMxhEb+rm2XqoAl1daewPsWyfEuHCtmEUcE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
c/o+A+nlAg+KvPhsbTgX1YburmF420s0eUecM9CBtUA/ltuxpGNru5SmRLdmFKSuHfhaDtL52Snq
S86BKggJMrTTe7E3laj0erCZzoDo6iIrkWM9fKg7Ngi7zJoufc/ya5fG2zrHQD/XcztjEiGdqZgr
Rx5B2F3zWgNfEHD+VSDqe+q8uGlLMyo4HGIJ3itZqfoU6X6hQu9Q8ifpGk+qUW3pIX06DMlLulCP
GMGeDaNn2YugQr/herFfjF14CjNGxyWQdlu4Fe3kWzZ/WvE41CxqJ/fiJah1VrJ2aQQKK0icnYfZ
cS/OxzgT7PexRnhi6lrFBWbwROs/GbEv15N06w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="2wFC/LIqmQyqFXPJmceJiNTrr+E+exwR52oUkRIbqtw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
zpgBUmy5cSOBcoIm3TX/SVHP73lwdUQJCz4Ttytpk0gN8GLw1SLAMB/JoOSIpGA/wtQY5SA+lMXC
vTb7kmDE6CvKc7+fogv6kGcJWejZfxqT/jIAVYkwIbSG9A4WjaNzFvXMIQe6A5tPLI2OdvGTomci
N0/UWIa7htX1Up4GYQpHL9o6grrwGC1w/QbvNzzbVMzizy5SsycOdYVHcalZvmr82mA4sJP+5/lA
CiMLfxMwuBGFggbTU5pAepxWXu5kZSE2BqiBeqzrTy+rjvYr2fNuZi8Q05SdpbEPFaDpjAkEuFy8
28ut+NFqAgbuIOZ/HQHZX9UZlMX2SY7gP5cXc7YdVXb33L+Kk0khJvkv+YcUqcSJl0Ods4qYtGXg
nFQ/ZxExLf+xSK+r+pxAjmz8ppcRs8NcyTQv313wia0RmyD+6yD+xTRALBFCzGUmuJnpQFd4q4UR
27TiZGzCK3scYA067y6k3KorDeumhAqVDhI5yy7cQHoMDIxB9w787CyEUAPkKLpVDKImu86f/LBI
JfCDauySvGRSeOvuhlBcAY/HLBoq8ZsLxH2zklPNk77cmVoK6KzU3tD5NeqTCFP422zamNybf+it
SoKATl/b/yN5Tje7DA89E6P8pMBgtlSRzc1899DBMonfJkP16Bln1NI4f0XPZM2SzK249QSy9+dT
mDkgdAW8cb4d4mXR3hInZYkZdlz232z8W75PQDwKj98Ng4xYe4iBIxgpvqfX/yh6TaAM4jG4f8G1
8Kzc3JLh6juy4WzC+4ykvRlfpO/y/oS9iCvX9WBg89YqSKm887q45KPgBGiAfdUnWDuKqNPScuIR
s5ZYZknMivpgoptkXjGOiyxZQ3f3bHkLib9az6n9f+AloBEZTol4zxrR2jClxvv+ErgAXbjoS6Df
bdc01J3xJp4/a8XWix2kyoceTDqSZtare84YdNIW3vX4yxvRqDqrKl04lsjmXN45OupiBvEoXrib
iU/nAH2esdL4oSzpGFQBWXm/ALgAJmbQJbrH3m+KGfFsQ7++jUf1IBfMyfKZjLn05pTt42JG6Qxh
PMZPXfkyNXIW0CRHsFyiY1o2FD2ku0752lrC3oLJEsLxxLsdyGjU0snDPgi9htV9eHyStK0R+E/d
pwD/JewHU0WTyQ3Smqb72YqB0A/vAg6ClNR8apt9i3/won/A+LEC17wyDiK/K1eiJSviZ71RydCh
4o1OjTRTiRAup0AaLHvw/jRxlm+/Wg8vfngkUo35h/m5/0qTXfsOyXOz2KhDjO8dIbq7i5vP/61I
B4oDtEb5vF7ML80TuKpCX7+NiPVlBHUaBrNoh9MKeHoB1ZB5wXeeAqP+Z1jJM6qCJF8Grf37lwl9
eMtb+1eklXBRDeneQSS7YVlHswwmZtQBd9hR3NN1sfLcNiYDU7BcoRtaL5mGf6TEPHkgFOjJI3DC
CAGpf2gacv6S2bti028vJ+RrsVWbgP44PU8q9xDDFZhGiLHReAzsVL8ZG83FGR+ZweQfln96vvGL
R9FGAUNq+F3TXdjHR2vmYOjAeHJlbmqyxs13Y5TVGKcse5LwSXnqSqmlOXFNQPcZJfxUbEZl9qKR
fgHsb+i66DFvqYnPm+krD5ZOYt1vXdsOKke2j9PahohFlv2mZdWXTHvNaWoft3eFvlKjvzvKl4YG
vTsDwdHaDlsOKhKZtjJo2OFufI+ogHUiV2aKr10H0ap74MwXCp8HQNiwkJBQ4ekbdysIcEKaZv53
nHUTJOtmyAs4z+IAoFaeSi2knajQI63deDd2nUzQQbBqq/k83GsNnM+/pk6Ny+RpFmMNTI9HxaGa
2lRvGh0QxCYl6dYG8kDCdKo3fF77F4NbVFbLkC8ylhwCYmAoKwFqJRKU2swdeH6y7kAiKTqUBldH
CaW03zE89xNDnAuh41NSwS0CTz3AszO8fu44D5FONZkZC2vy0nuiKzowgsQGdQ5tTYiMOP6KQwGZ
wbScY+1YgoU0OhUhgddFsWxur4LaG72OsY+OsekYevPd8sG2GJsDLSOkUylcXk+CI5jkz4HIK9qc
ZjOwzSOq2lTfyINUiusLKMqG95Ftk8J7LhESIW0FftD0F6aWPaa4tPtiI/x3JsLZXOBr3PAd6m7A
xAPKCPBE0AZ00Q1mFSOtcO9Ab2nRWDUSojuuXUrRKySlbZaLjj2ajlH11utqZkzQsZLIhaOmv+oZ
mOvoQJvMHFkzQrkB6HyrHMYYjCV7jTdavhJelTYFwCiuwXB/ypGk7I/HcduUnL+CzZd03tQYqe4A
oQyskk04jN3WPCMteHxYrSFsZQt4RPUcRd6Csrn4Fmdn62diyZ+moobbGzIvBAwgx35uZX973NEQ
8lsNsOAvzc+NEeEw04kM7mTDNL8o0QAcGSOIqPl6mN5x/+NGjXHFplJWWyt2t+nerG7u1FEOatGM
WAMJCQDLBRmkWC5HQxTu4CqdXl1sIgV+PwrP8fn3En00zAkz2GlG2ia/6NC8i2SayuMWK/AzxIuz
FdVnLTtNqA9ksFuzU7Z1kqJPTxER7P9Z9O9DK64IOTJp4CjH+9LFLBOSLn+0dVRIbjETcWtd7iA0
JDwwgEbfPYNvmy+Cf5u5FaS+8Y+4Dd0Ug0tVUlnQTVRcjT3GwmxW7akrcvDgX+mXlUNMNEUuhwy1
Su1cPGzhpyiddP/p435VcbBDjJdejNo5pXHXHVq3jymSOH/ynsQ4g48MEfGno87ThOWiA6JoiPcc
kRh0PHNMaOra6vmBBiudtGDbA8JANpcN6dxj7JJWQwrISd3az3FLhS+oNTYJawsPlLgyNSS4/YIs
f+AWJe5fe4xl4J+8JTNr5tBfWpHxzBe42iGWJ2+rIbdOPpuls4DtCp7SOPeN5tFf8NDyifKV6KNF
V+/X+uTqrdjE4a+74biAPuHWtc2B953zaJLqdECWMC2ltVX6T5t1HlqRpWpxF7yUZ0a8ZseyOYqy
t7zD6uiivwdcszOaQitMspADiM+cCGbwr1Ls0H/AnIBEY+Vekz0YJd9dr1opgCwrJ6OVoianJl9b
K9sZn/jpEB4iILsWl21b/j3AmH4/sh5hNCfkhATiPjXaDhvmUZSKnYDga+RFh9izsm/unHLGTvbu
LP47ZOiu++EOCflNzUZNAbnPqJ/8aBsV82SlOD1RHCL2JE3CaVyqR2DX1+D8e9RRUgwE64cBmBqU
YTUkNS7HRe8PAnoplxZcK5V/o51nD0k1FZVJ95tV9P9iAQtY9tyCqimhZkj96ZoDtHJiIb58B8gp
xZ7YbTDTrxDE5iDV5W3lYOvNXh6SPvzeNXLfvwlDsntebCQbhwlXO3A7gxrGDcY111zd3rYI1eOs
QpRCuAPEst7mLDpLerPwrG0NQviYTFtjBpAAeCbSbmbxzL9QQ2yb1St1jWFti8R5lsGNAmIlGgJ2
5s6uFmmAJ6vWBqQY4521Ksvvv8qRGbO/CIUDgeXP4UZOaWzYpVHIF/H0gi/8Nnfs1leAQIl+KvCl
/1rLxAoCixb50vF1uRMHNes52yd/yEDkquQ7doRtzvZLdNgWXavXxF15lT/WfCf4uxxaIxBlx4SR
mdwv83sekLkrqFVR9Qlr8Pq4jiJSN1zy1W8Mv3Uc3owbsNIRx2NboqGPWL4qg87lBDV3/eVcQ7QM
ALdRplzWBZBvMB49wOl7x2HfQ5W4fJZe6EEMig6oIcr4YwheYyWxYM0DcPf1wSYdfbvukPCUC3eH
giPBVM9jZdn8NODE1uRiCu86I3tBUSU3rq1V60Z0SLcn835S7fb7dF3HxfICgqmeWqSNNrbD1EKa
yk9/SpI9lfux+q3V2fBkt4Wyk3EIX5ih+92MEuMVS2CXoC/N1cmClAdGmjRDXDdgblYrbdMKbN26
vf5zpqyvExnqzUHNEY0ZBDkUvDtEs6FIwDnybjnqFnu8lmo9gLqsKwtGZfZQO1JUH8o5NFcArH2T
WJ++uRFVuqBVf9Bg3AY8fNRs4s8xF1W9HoT9tO2dvPsCwVYC8rV48ImCoUXKJZgI2heH4u7oaJwK
CAgeuS1rF16OumddsQIhKtWOiJi04vsjH6LmDXjYfORvZkqBDIHdQe3nL8vsVxgXY+NFvW++MUiP
ylrYSzjZGeUE11Pll/3K2xmSjwqAiEsz07u88014cWHe7jY+5UQSadEEi4erS0Ktrq/id45UVEWL
xzngNi6P9l2l+Ja/eRC0gEK8zInKA1+fmFj//Mm+yPbiICArY2vVpROaIVHbbirDLVQYyyJ6E9+E
z2FzcPnmxj6Ag2R6tmtr3dAC4KR78tIbp41+Iha+F2YYrpetPHwzdAtmKierX5NJ4L2Q0JKf31oL
MuuD0ETdWUpthoJ3dwVVWlnx42aa6D66WiF4E8zwaewGpQgrHBNyeglRhQ8FBJAOVO4JEtxQ7VHw
uwqpx0HY+l0vXac6djJ8eUMNrJUqJq2ld3OJMLBog9cRU0QAwm7oenLySPMrPnXUJvyv2aTASSat
gpGeqcdLk55KTtcvthLRTzfcYeaImcDJJx+f7j7nviraChZfDyXklFXBZsUNzrp5Xo0Ew3uh2Txl
t0Q/JOvkJkn82MUW8ep6ySbcXWkAllEJnIfNd/hoA5KVXWfhdtd0f52GWsjiT0aq30Z5ttigUr/v
GPJFnRQrSQxu0jTGYXbQkV0e1T9SSgmaBBw+hR1ihptddwiNBe9n9qoxTcPyoqmGHVM5XXtMVmrk
Nzew+03SnXob6IO5fWHHYTzmMhTaxcTG2z06ZvGVLv3/lhZhgYYd/JC4MLDJtyvQVx6i1DOUqNfr
ep5P4MmLTUAqpY+Hfg1ppduxvAwyJYpGs05Dci8NILS4PqaAPsfJxKF0FolTzDZu43QZFxlqz0i0
TkfVGyxjaG8BBBAEtKTsloadH+ePGoWu/536sepoCtiRSN/J1lyOmLsMrhPUdl064QzQEYevjwAr
cQmesY6rx7gzSTwlVPxRiSvaA6NLImiF54Rqwz16tuQJLVTwlc+a6I7ewCPBCX0Z9kOFpKBO7uGg
cnfSFpaDDzwu6/0JT3XUK2C5iIjaLW7gUbiCYScShi6BCgY9bOdiUrKUZBH2dubbKgPDsM0wE08l
Y5Klt2BijJeYagHUmRI20FGgyWztYf216Wda0fTJxVjAmZXV+vQZF35OIMqY/9un2bVsj4NQqZFj
URYc8ok2B+HkTOheyu2VBu8LmWYehVyYEg+ITDJYIvJxqq7M1XqZfPt81zW5Lp6KQ/6BUwY2e0BS
8a1sb9DrAoJeZqpQmXmgV27LnvYh0z4ne9XBTKHclciVDKgCd6O2s/7u6Tjd0x4kIj1lhPdbxsAP
llAOirh91kBmy3S0OKvprap19pxEz98rMCFZ80yJGwKDL2dax5bDq+4Dlm8CIisAK47h8KkULdDU
MrzeGpi9w0W3MeMHnhrKIpP1lKM1gComm6TbzJSx34Un0pwhlqeEgxTgk1Q27f+9fllM69x8izMr
WCnCm0yXyDHYtlsXVUXRQ2me93POv45IHDjmuMOFNSsXWDo5Mj3+TMHmMtDGLIv+bPTPJmdK0a20
vOxQgZwNXNrPgoUtfolhbp1ZflA8ycZw9ebDxfTPKtW88pnKzc08iTynyWfPVEg7WfOSEAhs8ioU
HZx9hoYEF9twpwnegBwkPhs2tCSnvu6Udd0zFYF8h75pPswtS+BHpdsFlO25BfRVtSnFxlFO2Km+
LWLlm3iRT8ekUoywTI5y8gz+FL7bWFDJP/PfPKynESyVwlcWuRiHd1lujV85dXd0OpPo4g658stZ
kFSa6Kzn6KP0CVgoUNwiDnNuSbZPZ8MXgoMeErT3VhHiPy3l79HEe53xaFjEqAi1TfHlkdU5hHsj
2d3DzNjLhbjRVlof3afVNyhNYZ9V9ms4Lv0MIleH9tKHeLX6QWiQeSHIHCbe6PwPg3VceT13wRwr
TpKqtpZyUsCaSx1ZqyzEUb5tTlBm/+gkofY7BuOE2ra7x2yWnTMWQ302dXZI7Jk9y0N+mo1OXwbf
bQup3qB3q8yBTMenOnjWvS9Fy9pyW0A2qX6i9rITq+ET0myVDXs7yl4PgjcRWN9vk9W/RydhaVPI
CGX4ao8riVYX0KVjL1qfY1Fb/4V6dCtrRkIOsLhzlQYpm980oz6Jn9EjTW6jHO1+fZbljhNHCsCT
gzT/HYD449oOlpaiagP8Xs5FvxpT9siZHkkoW0Haj6V9swWlaELDy3YmCX+bPgsyrcJXvBSeD1T8
zI9unWsO4VyN2gT5wSmcKqCIV6bW3BBNMR6Hvc9pUKuA3iXemtNoEfxOyqMsUHwUt3XBwVURjUuw
im96GwGTSHTW1cqt7+ycDr6gR0Z+Uxg4Hh6zLHzBXiNvCOf8TBppqLGG6sF1HBMbDKwq0NmEnTvm
G1kqszmZMxLyNkK4eogmjmV5b+N95YOimGsIwaMopU+sYBXMxBjsvkOD1nhpDZP0KkicjkAcEC3E
LnD4ADyr3KbLFXEJPRtopzlizbm5VfMXejMnjJsIiI2I2DJkLVOoozP+QTcZmOfg2tYgvThdfnid
WvWd5tPrtXxS18xyJ56LHlopdwq0UxUiIfRZA8fjVIjeV/PvUAbY/6EB63zjsn+RZ9HTmO1UjAJJ
vNcoKtcCgxVtPRGOSrP7EetiHzXj3Ex3E3o72d7gb1Mjuk5XZLj3dGhM6lV0UxvqGGpGi9/CbxLn
s/t4/7y/d4zEyB7p1pH3aTFE99xTNi8CS2/0etAH41syGeghTgORsojD5eeTSnxhMb+MZnOgNmyG
WXIWPiaMDvlbUZep+UUfqIs7Ex1r/N6Nh3ynZP4v3mBye0M0fkBWOfxbWd4F9eWMucdXaHkfufQ5
Wk4sumHKWEYlo38S8MpuLHKeq2+t4fiVF8DShLsscg9dyT536tLzNm4gozO8LUPbQlhpPYpEQJ9D
/bh/BXT3iSyAHpRGg6kOkfUrnEjTDkS3I20RWDZn5+yrz9Ei5LaerXPjgpb6+KNARfP0ac4lBQEk
k9QDCofoV/VxvOg1ufKSVxZqO9y8uvWOoczV/9ZaEUfMFbXIk3UpqT+GqIx9ZqgAJmySGglsPnmi
lPGcTQUe+n1PnsY=
`protect end_protected
