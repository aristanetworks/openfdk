--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
dMGPDJVdCeMvNX78m2ONQhS9vgIdhKpIlrKQZTUmhtQvarr47OPwH3UnDOXQJnDym11yfdlev1HD
sGqY8YlAcO3RRbkwD2JpVMCiajYgbsYSz38k+MVOddkFhpoVHyymr8jFBEC6uZ4RI01ZiGLdckbk
mTgl1/yAxwqMpp886+BNqMffWriWNKxotRO3vzCTvzauN7JVmzPhnIiSTFfNhJqnuzFb4w7lA7iu
xoJA5lYk4D8Ba+qRKR6loDAEU+cUh7LPr9vJ/qHAMOj+tnUZO3HyDn+3fhjrD4k7U3X6ZausnBgr
NSMq1hZv2WwPiRy7r9ns3QmDOVzxKVqIkTdusg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="tarpIS/8bbSdGRnSwgAK3AjLaH+mnwTSO9ZFLsaFrIE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
X4ILKUkWNAfUi5KCvM5eRRjdrjuEOO04exkerPOjxjT4uh+WoWWJGol4TnK8+Iy8jIv1O3T635gx
QaE6VWoyjZea8K1wNBMNYXmifeDMIXnL6/o/dgd5Z+vNZQwfiYzd+jprRR/fioRWfDH+iFSV6itB
MAEMhpsQ5w4PZyO/kaLM3VYGi9xhItgK6szAhlLCeADrJsWNuISd76kWXSTnowRBye66YlMmmlnP
wauciBEGKy60HPSqzmQeRQXWHN17dIG3CfcgihmZ8DFv9R2/pcQH0uV/vP4nAj8mmy7Atm/r2Kjx
Mnyc/ClqBO5WafHN7hfw6hbqx7N+Opl4KJbO7A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="A1wQs2vCn7WruBnjhFK9GpiNTXsyo8qOdxFrmIjFlcg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 61728)
`protect data_block
+gcI3e3C38X2RhN/hKwasNWLp83da8+0goiI24fNSvtTudP1yli0YoVDL7wNZmgVKqrzfWZPUVIi
q7gBUbRHTnBYT4p9ly0IOwxR8L5naQLztm5knT4cBAZstyouL2Dix7bX1g1eGgHZ+3FIzmY/wgb3
BHJFOk2fdhyC1/4ltDw3ewLrude2qD/tIBZYsHivZgMR8cv74fuMU0Iysvwi9vThnawbytKVxJeh
RDos4BdARINmlMyre+HwEVL/wQkZQpK/I0B6ASfyiYgIfKL3afZaLQYqGZ6LvAuV2jQMW2pfIx36
F9BKSw4KjZgRxbcBCehL8NvC1hGFenfinFMvIZYTIp4k9tbELGs9OjmfxkIk5OqR2btKRSbvDOin
OyPZjPeH11k7bSZEpki8GxJKFaSnQDV9FYhYmq5KPVU8oZL90A14f9webeVUs+qyFUUd4XtQTSqz
rVdSfoSphLiX56PYuKHyqhRhz5K+vfJOFuB6x5Ef7Tl7BXRqoqrkG5AxPqDYQ2BMGIvxjadaR1qF
oDiFFhCs1J0kMQVfgcnbeUfVkh4GD5d+q7UGGuf2JmE/QSsm3Ro9g63XxJJhO+00hzWyJVASv82A
MsE8y8V5LkS+4MZwaGjFPAUe4EQnuCynR0dXP60ELRB2C59MUpXn7LpEIKVhVgeBpY/s4aPMDLxS
Ht7JqMLtxbFYWXimNJf1twVJG78kUEKXkxc8NhqDXVEnKA285eInhR6XOLz5rthuvL+majYVIHNr
AQ6Pu7ThSmow2t60i2ifR+OukTUK5OWhuJbwJi5zT+8aEo1nAzj1ytMIx0CPpa98mmkT3nFEuaTN
DJX0ci4v/Ayn1hEMmTwGT3RzSN39pd2FnCwO10FZocEOzO86VMODiKTIe5gQSikemcQwx4Jpe6p5
wvD493+2rxzNqPOn2LEA2nDdQTsjUtwmkvRPCdaj/aPVGld6W3Rttf2fKjbUKoU0XTfs3CsePHma
GGh8QJDIH3g6BGG++hn2sB/iaGIw4Z/Omyg0sd3wux2atTJETuQzPG9kbZN+GWeGeV4jPjskjvil
ZCtb6sv2S+VnnAdGJ4ZohFNDuslr56GskokFpPHfhJvsETGAvFG7FCcUTFMT5Tc59CvwK8X66LGM
hs805zpP1+GXm3lI4/j6mDAMmUsLuQANjEXFcNe5pyiEwu5JpMMM9oSXUaUUM2YD4CKUt4Zjdgei
Nd8PARad8ODzCTNrY4YaioYPP45cJP3jFYQdgCcerOnsPhadwX5u2/HITprLh0W1rFKZvupbsbfa
ur+4N1yUZYujgzbyrcioGZJ3SB86ZbJZf9JBY7mEBSYgxvvby7hVUGhTPtdxV44MJYxDoWqmWETi
sFUTV5u1vKfYCvO3CGyPK7ruke0a5/QG3XyI+sv+k9frNFsEB+VuY5qM2ZgYCdoA90sfJbc8WbOq
KiYRrt6O6PdKFwouXNekUrG4TFjg0KvF5sEkLABf5pU/rMRNNg/xhOhG934RHaotd1oOvNA/1blN
3hsHDStN2aMHSkuMzedEISorgheAyfwDouZhQI2RA1rFCW0KNFl0iwr1g54ttS/S9ENEeKyM+uQO
RKkyRnMvyjwEtrpiu2PWS8GihzE9OOYXtXbftYVIYSsO6DkgvVyLrcK+lClTNcO8E+eBeT2gckAT
VYv4iXZTYXvBCZRlS9mo0ieofIBasRM/agrjoknlrUiN9Wy8ggr8goprDaet+NYlBIJpJN7KCpy3
IEp/oCZwalBoaCam3fNfw3f04RLWO6Rm3vD3x9F7WaeOhH3SLZ7Te+/YstIoxFixo4wZ/W7eX+ok
ayTvhsIaLrxZN0XLFxHYUmeAtzHY4QCfh/ryh0Zuhnzcj8BMGlKKeTtFH0D4Dp533IfR7OXqJvlB
1PtmsAx8H+2wQGB5vuogl/fy6jbfppzoAfcVFPIFEjkjiMeq9P712qhv+FS2MjPQhPfm1ari2lr9
7lUp9W5lvBHfl1ibnKGiz+psNyz+ILpb45CBm6Pk4r5p7xbyVbIM5H/1RdbnlQ6oPzlvfWrl++mn
U2ApQrwfHEwBUzxo/JUb0B6Jdt4sbWrUt2ggp8mnBDRceaGbu6I9G5Le7M5IQja1wR/+f7aGcSR5
vEEwK4X1GT0efegMkziY2AU/8THZwBNa82gKi6aNcP4NrucX+R+AuSxHjrOok7xaov98IE/wWa1R
x/2U0ztVaD5DT2sKMTiKHtAVG3//dP9Vv8Ar5EXXBTgMzcslqRMNHa5ad/vMsxaQ/cwfdPzsksqY
9K4m7G9EtXCHsyY7z0Xz1UpkN+KEPg6NQePgaAoiUAz9bWjuf/UjyiJhP60LdRWikp+vKQZgpEU7
ZWA+R2jGNq8J91Ym/OgL+ZRI8PwMo8M5yBIiBNOHkfk5MkqpZ5yicCcmTX5akHOJEmrfFYXnNMrk
3kVtndwy9d8VH7Ii68QBknFPiwDYREGYGpfnsEGltjP4qNYUgS3WhTrvT/nSmJfNmLhCjy6ZinXN
bzJ2suY+7LlDanw1DtmfsVGQ06YfbBmkrV/xwoJnAScdg7XrbYX0vGLZB34+2IzKHpZfFpnyvhW+
6450GSRsELCPQRg09Jvss2Z1pUHAj9H2ZjFQMwsPfpfe+NoWMoFPBASjfs0irSgGPsOmDqkfP/tl
7RDnaJLmYAhyUmN7APfkRvEF3Qp+73Mh9HkSCjStsMT1heQ4TVyUwIb36TSoS1WHRqTZrG6dVa5J
itKofR945V1DJhqcUFIkKIaRpDJSWvI4iE+2GdLhx0GFATkMuQrmJoS/3mMfpUplXOavm+HX7tDZ
HZnYiw/9wHPEbV4GVtBSvuhS+PF67tvAtk3j5fu7P90ie/4ozoEFF+LIfLv9ciuyOkb2OmHE9aNW
oYKPcW4xzt2Y3mgKSGXMV5yfX2shcD+lEHH+0ljUHTJqIhjNc3KOK2K7NaDOtjve9yyea4eyv6Hd
DR2FYm0IiWfw3O8PUB1HbeIKR+42bNZuF5L22jotHVASsgTIo06L4TkkXdqRf03qYDwFIK7WSzjW
f/qe4u2Kti2LJghwDGcWfhKuZP6BrfuG0Lf/sUKaEBlAjdOQo+46dKRSrluwle6RGqANBCa3d8Yr
GlLIIGPmovLHTIGlfrt5bAjdYQe6ienEQLk33+6mkdG5pkjG9fLPLeJ+44P5ZAejXMmAwSNB+U5m
mZE6E/v1xfsx6wn7/+3KCkPMIemJuX3S7ub88jZmL6LvuLd9KHERwhiF6s+jd0w6PkCf95YEpYW1
pAAngVydb1SdRDpircmpGP0LEQoV1eLsEM8R/ZPVbf/iQsFWCgda5MhgP5xXtkVTd51bWw9SoiYM
fMUFuCUo1sBx7d4PWXWXM8I8gEsIfQ4u0AZzshfQIobAR1W3eMwh39G5rNURuIU4KHUYgepIvSeE
RlO3THNcGwh6fg4CMIwQHrH5ud7XxJKYT7S+VrDw5RNaWouAciKEH1TsIlcsxdEWHuklTup/dlpv
R2voKpYHFFaBMYfFyAixMuVwkLs4QvtcyJsC+ily5sfOl6uak8jxjvyq3mzq56MmiUTCWMzBlKZJ
4G1mYfC2Br07YjV17Nzyw65jGkU6hOyCyWlxzdRbwa+WOSjg8ekJ0PoP+0kgH/jrHLGMLbEuMW3y
pdhQLEUUH8axVztPAVgnNbsUt9FWz7H/BJYCY+5cHa0M/jkxkON+wZmF1W5aCFZ8Nym3cUHAsyuB
QoVgJ6MISAGnsmnlaLUZEuySgliZoyae7Uh/KHbr22qvR9+Qt8dlVKrpqptkFG8Vm3im5ujhMQFS
9EK0XtlWtq4OxzSMtHvhzHGBM830Q7ySp4kt7e++lqLJCFKcE9QhyvHinAXpnk0+qsZN1gxruxKu
xm4qkKb5pd0vQh3yeV2z/Lh+PXBueec0JYG14O/5fxPNTn7MDfgtNiAgWs0UKoKf+eh3dPmax+2w
q/F+DwqDk0BP7KRUl2HioSv2iBtaU6nr+grhADWJwh1fsotQO1fnW5WE46MB2fUU4mgNxZ65KDz7
LM2HHYdxfeX3hmVi+E+SOnRNsStfsjlNeWhqo3uAjtJrEcg1coQVGhWkQwydSYOYouPNT0zGsT7t
x6V3PJKvsL5oH1tV3495G49ArhRekNyDVf5IGLxysiGHuCjPSua+AJtx4Nl3mLtxcVctFqrLVWe9
KA143TctMiJF8sJXefQBlCn1W3sZNyzANCi9dBYDhGuw1fHlT5djKIgdJ2Vy4K0/MstUuHRCCzfS
Xdh2Qe0WgI+fjd2fSGu07MT1g+N9bNE/yquuAxG91Za81wz66Ia64QsVtf2cQcqicIsP9AgKz3vz
BXUwW55PX1pRw7b588Y/g72P3UlMtOYLBko85E8MbgwGoqCS0qfbDoofOxHXcayZLrSZkz8ezjCI
QlnLvK2HjwoVQQzncgUOXgeHNCG0uce/z2Lc0kBZtD+wN9RL3noYXpnRmBdvCi3fCQB0FwbK0zJS
iYdBIf1aWolgAbna5X5+HtG3YDyRuzWQS5u5A560bR0DkspI9vx8TxgwdGsHkLEqjV9XEx8xWJsW
yv2GU5GX2Yc1vKr1vr4lZTicS/9Y79KIq5DJXysqh0kbzCwtLuk6/8ODW/bbZDfdE11NHI1vy3xr
7Lb4VKsSCPsRdJTnLBD2FiK0U6LXazyCZtVMgI+RM5ffQ+hBprGuuYrnjpxwBDbRC1wTU04X6bi0
KOzYUNbu7UH9apz6BhRHvZuqDY7wBd2dMidRx0cFKY4TvXx+rTaG2oHbIZ0Tgoo1WKIGKjpQguAI
6B6GofBcjuAuPCCQIwlJOpoXy7zAkIRq65EcHtyBqv0nHweecP99xHgr7RKdeHV3ggJp4Fn8TLC+
lSW+8pfwNe0++pInSyC0hNHvkM3NTrVyDdcPbhczQi8H/s6sTP9luXgFUO3jJdQA3Pw1LKJ7NuM0
nZ/rkDgqMU0Nxarcp9AGjxo9eW/I+LSPZUUxDxI/dlo9OhG7POHbV/cuqlivvt5tocwpIO4AlFg3
EOCx8VCaMWaHLbkxNC6B4+ciOp4xt3NTUrSPks0hR7UrZfgfRUYhgkWUOLu4FwmsPpUiZ/RBlD/X
fr5aA0Zl4Y+zWbp6PbZ+SMjCiK3JOTnb0KavRl9s5k3H007DZGypdfdWXU4hffPAYzL9YdbDC8Ld
q45UonFwck1SXUpwJnxETqGIMAzqzVm+Q8gIRPLjY6cP8k/P2S9qUqmL/fnfrYDuZiCJukfQkJeu
qyboIR6dS+7SkkiTzHUBpt7LFhP2J4kTdA+EvpipqLvOo4vswOMkEBzo0HCzDEdIKceuP6/dBSDf
FNRmeJZK/JQuS/KUeJ9+pWYx/h2aJMfIt6rNvnk7nY2Gp8ouqbA3xkr/1uanAMn8nk79jc2Zeu3P
DfTHcqFoMcbMHujFCSHRZf3rQyLsJ5I8opwitkRhJ9l+g15XSpvyv4lpZ8W4ip3EIkWOO5zwwtL1
ZGUGoccteCH729l9U5wgATontECo1cAlCLYx2JJJMVxvqTADRTRUc9rEhv9/0dxGLrlWCQWIdwvp
UyL9ki4l25cgzSN3SIW/vymwAMpIP9xkCdZqhTcfXASZvVDB56Ia1Z5Tu/Lwvt9bT9EYsU6oK5L7
VdpYzcu3+L4ovntm4b5H43bjYQEH54t3j/bgJRJmLRt8O/shcdbLrryuITSKk62OUU/eiQ3+HN5T
trgPbPdZqq0FT7GXnentLKCBqjLIszBdX9ASI4pLCCPIDPr5zlWI03DDxPXUPM5HUB0aijgjsb/1
s8oRmKghSG4rR6Ktfyokb5WXiVLmaOT/dfxg5lAmk4IE1d4ix8lU9RmaKlWXfH8yvBxcSoPr/3yR
3zicam2uJt3+hIFgx+4Wb2AlPoTor7kUgi/RCrkZOqm+nUfjC8XQw4tgSuW+nh3R0K8M73df2Z/v
yPyFFy71lBEt6+YY7xHVHHiUi1B3f/xxaVrJwRio/q3k46sNOJ9eBzbI05BfBJgs4zCGxO0wZ/mg
+jzJ38IoJSPhDUXndycp7YxpRfO7ubUzL3FfuO7iJeIWDSB71mBdDJ4vopQvI11bTsHAY369iZRB
QffT14cmXRJB/knIQaYtCevYArLo+83AvGxtOFkrD2suxLf7HNwSghE//8WKDY5hWDcmeCkoGXFK
hUYedK/IZaSlQbVdydGDIuT3bc1mMSr/Y7icSs3wtnRDZdMbctiKU3EVYA1ng+apNG10jJMBe1o1
oYbfu0Q+2ny4pUixjCzOPAFayYwCuPTbxKiX9fU7DrbskBmSNdT89WXJ9Vwau6m2gtCcfvkGKKoG
3yV07xTeVqv1CYNlbvmMaRyfGduzyhJvbTL1zdsemFw/T4fO4m60uJz0Bx9hPi1WQXV0I673ICRQ
exmm2SYDOiMV8ozz8PSRKseb/ipqpSbqw0CvVzxuXlsoyGucJ+fw+UbppsUbGy+AA7RcvjrksqmI
qgu3Ag/OipdpemXVRt4J6pnN0PAXqu5DZn91zEwlYEmvK8KsDf+fv/kCT+/+WA/FjPOvt88rpmkX
aOj/bcavNj4QvcsMHy5T56Lj7HrDgZoT2Muj3kWPFdLiRtCL+sZLHVLYM06orQu9cNdQVct6HAQq
nK0rC6/M0AIzb9iyPXGM9c6ErnP3LmThY50saq9JAGtvcgnOlJAWYvyf+Pm5UPqctjStaVPI+xH7
lLxAxxh5AnBendFKClFuGij/em0RfeLZla5KtCUZWteLjdt7x1iRT7T8MclvixDpDCZ3OKUVCYWy
VEpeYKK7KZUIygzDBhSnCW1z9/fEll/piIoy0UK0r9prsf4omhFkUO3oHO6kz7jMYEaN6zZ56xZw
VZ4Oy/gG6QBql4/skTmANWaRMmg9nfbu09j0AYlcd45YCK6m0IXSb+ALeoyJqiujQ9RAGXa9pe3L
uRTSMbYBFTM7pFBi+mYFRxHkKkkDZ1obdQO/Xj7rxLN4YSx6pmVejPiwtmVRVz5csbHuG9y2u5b7
PsuTjQVGWXGLzqwG2G/qaTWCEB4sC6EYzfI7rU4208ut0fwyPcCtagi0JKikqnqfCudX2W4mlDKy
kgxxhTRG5kytWoKhk45IjZuymqujbKdADmQCr2d0KSMw5r+eLSKv9a8HwbH2C0VQ285dPu/XahoG
a2NKvZ2fPY8opq2c5qa0F+8riJs1aTMj1FKRIO4p0ajfp0P27NvSs2LGilLt5Xy4bhvU5ATxiS0X
tuZg5JMenJuSAParr+LUTWk/o+m2wMeISJ7Oik28RI4Y0vdF+ZMfiCaqF2sH/w5Cww7GAKT2HXHN
c6My2Yk7FMl3RvBGBmASMvTbJKYmJpj9HC7A64yhxzKD4uys5axZ2GVN+rFiHG2omotkcXwWTERL
RLzGKUb5WeN9KLJM789f+OSPPuAeG+u1zubf3LfGURA588EmTnEQTl4hAJaa8y7Vrly3TSJx9xTI
hlz99GmBE2uuMtLQGg57DKeDGE9VBbZBHC4syy+LbB754WDRTXO5xokOEI+WNLDMh7tS6OV69k0R
c/TnkKLRoy44Pymzblou93PutwdacZgnkArnHjEvg51S4mMgzFlRNVfH5i57ueyNOQucm/a/gTit
VA7FwBH5MinWKq8F8MR072jmAdJcPBlI+rH8dlaIt6qajroqHisJDVjwKr4//k6hwGsRTl0pzfC8
Q8fPbmcXX7tIP86dvWpBB1LA+FmSA2KjYahpSGqlyKtlbzh3qODTgf9Byla04Hs+5ybA02/+7wOJ
/syXU9PDZWj9PdexNA0+gdtabUE060aH11RnyN87+6o8P3KNR6EfR1t+HMV7mxVZT4RDaZopfLDg
pkGH05+4EPFVJM0I+O28iwgiRxILSizKNO87hqsdQJHyn32xI6J0XU0v20QXly4V3yEXpr+D84ia
Giv1TyLp8l6PfFDlvfI5Cel69y8/vCP0JNt/pQoa1eO906gHgLU+DxVELz54QkMM848V9DDbjU0t
ReeI7HAvY6MFTwGhnxkI/m+WD50d9BmyG8/frnc0wqOTez2yfaHtdGz7gRAD33XpFrwT5gwwonpQ
TfUnjB3TdKvzIALFuP7nphDQIGXBawUUO5eN0KSCLomplaFS3UjxVgdbKIxyejc+UUBElJ++x2YH
ZV7444s9FVzKNnbDKjT2nqea6VKujBvZCypkxpYddksHaWpxZvKIT05xIf5AUoem8zU4inCpNm3+
CfEko8a4gXOoJ8Wu0ZhFRmq4rx63oIeWufb4iY066MtICTLRhWc5zPU7q+kgtG5QxN4QBaWaghDz
cmGiMCoE0lu8fLvMG1UhzJC/8FNRwUf2T5KDUelX/XFt/14ifDLpw7U3YKHxfnbdiv040lSV+iQx
rvMqxM9jBT+Z6KG8+S6Zs1egNHFqJN9LNcAQpRqjUzLk/f64YtOdE3PjLBli19kqbue3MfUPJbh5
OjrmCD6a9CZXrTtb0HyKQw1k8UUGIkRUvHW7DC7KWq/3XbCVhtPqq3d9LRiFFuCBzkL637W5tIIw
dVuO1bmNYsN9DOu9GZOy2pgl6wZY8PjR+IQ1rm6QQ1aOgYDsPTRch5dEpzQZmTC5NX4m84OIn0BL
WpkPZYa31vpsyMyy+f1RVToncACwQxiURzN1a6GS6sI7zhniEBHUEkXed3XK0bPQnTXH4vFZwBuj
d28Oj75YyrBQC1zUhv0VHhnJ4lrws6VVzzsdNxSMTE4VoRltXrj70OIc7kInNlgTCm5HHvPHJ2IT
v2v+iqvgtTFMRHGBmR5f+rN29nb45qpm0Vv3OOnTgLqie3DfzSJ73PgjvrISekVxme9byRhkOjZa
2Ye1wezYgtLvPkRKagwFDD/6f0JiXzFMwit68qZ9To9UbFy9MRY3SXbhMHBg9aT5rMR7jKmmC6hM
FXiQtAFPVy85/vsWGmnYyiYrdsGZVRdhrSNZeh6sSoBlLXnnr4Ta4720jemiFmtlIUV9VqN5nj8w
XKHtnDRJiiaS7Cy1fCIR9OJe/EY6KJUy7DRjfqUWkri4VfyLok/rg5BXSvThAEkOmPYACPTifoY3
XSUIrBhMMbJwddf4bYZxOiY2cc/zzctiM8w4qaO8h9ouE6H1CoHekVeiYGQRWwio5NVL0VgZ93d0
0iLuiyhABbhDWvkKD25IFyJ390fMrdtiPkk1kQc09QfWNakQppRHSSrV8d6SBtB3NUaSAq/f087S
7c7NC00pnsSvg3osKQpVwNfrJOoetOvxNJBPrg5ZsSMoihWkfeNw5GRfoAyp/fDDH8u+nsK71LoY
r8Z3jVBNTCSvMcaJcPc3/Qk/qhw5TDCDnzTJWGooeJC+4/V/8HOhM09Bs6qTUI/jZwxTRpJE0E+F
78eXnwii83vGOg7BSuXRWFZScetG8vHm9/W31SEEHrez3YJiSOm6YZddJ08TWjkktxzX1jDSLSeo
Mk/mH577IQl014bLvDcwUZ+zURsPA65TKr2ck2SqZFmhdNuA0vIWtyaPIwUgwUXgI8UBiz+HTSpy
WvdxjagCuwB2QL5ZDFLUZtyewYBBETNcr/qbSmhvi80h9+YahPinKJ0ynpY9Bk+V0EGbtO7rCbca
Z392kx/o/m5ce52ZejBN9PgLKHHMfYoKhQDxfe6yDODEqeryo4d7Zv010UHxYyk1Rbuf01/rA872
5TPal5NcuQckLW/nyjrojTsEjUqoo9pH8DsmD6raLSshicsMYw1EJVlq9GxL8NKHFyYgS2//j9le
SSO4w4hEZeCdYfdnLsQB4Dx589oHXBpv6BhUaMMIuLmF6tBaXG/KkLEhgJawZqJnurYnY6bTYC4U
AIRR/O43O91hB7qZyevqwFzvW55wHD8iGSxgU4N+7vKzlQifWUl56Qw/L+c6fXN/EC4tkLNDHuud
chNxfi3cWcFs+nte+sy9WDJ5vumSK/3DmmeSPrmJrWZ8IiGh+alfL6XHF1qONrnphM1uwigeOnIi
oSCNSbNDi2VExDJgL/wZg6xGEqqFke4RLm68Ib2dhbA/p/KNKhNp7XeaXw2sv1ZvZfcrOjpyQgIq
JAOJYD2yJTf8f4wcf8eU/jKIqCxynUsqM4/Csa3R7bd1mb+YDoaJRmfOQxwgau+/SiqsBbzcu9HG
oa/+jFaj/jMJheOW1+6kGjOMs/PZTqxkDk8JlEH9NwHNNX1p0YZGXVOsfSlpPBITX8fnI+OQLgcY
qjrw3V0NOGQd9V0ZIe/cHn6x8zxl317LW1SU9aC0VylLIPNcY/aiehBbW8WyJ/MHHfyjtY4xn7kI
ZG0QMkZaCCJ9vcK5b0+2Sp/ORdxCNUycsuZROq7oqaOKVxWpE0gakF9kvugZ6mzgWR1IXlSMLLmj
1p4zL0pSZZBesOJgU0pH6MnopDBKeuK6l78YJrBIpw9X/+K1quG+eGPordvoRXD8i9/1/TXrAwNO
ubJ2dU0GHIeB3hB2voFnCcxvyoGgutcuBLl4qzDm+SGdTD6nb6+VDRcp0EOHINvkl1kghhArUE6p
5CO2wDr0rUvQbxLmbY7JMdd8+xWl+26TaysxdT1vabZ8Sj7QTwwTIUPvARXihlX29biaFWAUMAoA
16mMmbA/8FVM4UNWkzHS5KPcAqFIviaxTpMXE8Q7iOYyozA0Ge327+teqE6NPt3s8hP7vVp3XTE+
23m4t/7gBJG/hWKO6W0hWCpPMhM12jg2OfpQ7YrUjOnMUGogwAWrSaVE+gfJsTt2XkhzYdVL6Jir
s6WVnKu6cQ+GRjmpeKfGTp0tB0bzai1eC+ueFdw4bNODvd0wgYuSgqMGs8ycYk88A5l/kJNMdE0j
7wvR2rwS5o+1tUisUSx8SK9x64TYv/m/sO/o9CCJYA09zXIsuFI9ZZ7kYI75EKEWZTOsbysveyyV
+8TLcTGzcu8qnRWnC/FQrLh749N5PVcQ2HpP7WtLSwbhI8+yWJIHX6OIR4d5paf5nkpKxiwDSSSg
A2fnqgsd0uLoPb9ws4S7Gyxj1e77xrp3L5TD3FFljhCFPBd+URP72vR1UOnxGHmB6TffLTp78WoY
ctsx9/30raG/fMEc9WS98Hbu/QPaEEifBATTzXJOPUvoj0+iV6OUuDn3JyVVx/mzh/uebcvaZkn6
ZA4mMO/o0keEYZzNEaeEZe0ssrsymk9Bn3E7cNSPqDhly87pjxSF3O3BwWhVEQq8zkHh9ngRZwpX
G1WnU9FEZ8Jqz/59Knus9WP+2EOEYJvPFgSRY1E/mmvZO6GspjCvr01eOLeTovd/KMiYB/M/PA4/
tiRK25khHImRHEaUyw8TBjQ7aV3SBQpfp3W0Z/k95E03plvzqyGb51yjycbaiGm/Bw2KaIrIf3mk
U3owM3V/sr3Lzltlh8ToSdmYJnryXg3LExtmVpWYhX6C97sXywK8WnU8YdXu3H/561EmW+hpfUVz
Gob4oXKlweHJy6OMqxO/l2nRsabnqbijQeQE3wWagt6hpzkwUj1YGxUm826+dbFxDMd9P1ykrPfK
rhFf4uHnuMifbE3cSw+qB1UveDRLaXY1Cus2GV3OxCqF518aSOUzFyDib5XCfOUDCiOUxp1rQPgG
OA1Qxr7rPlHNlN8qgmum6HKz84aBqnuUpBM5sGdCrOP9PpZfKdMewNewnyN3iBJQT4ttKTG+nSiV
5tlfN1nJijYg+OrLGUk3zb4roBL3YMxRgxfTkm5MbrrHtxhBYxx3GfqPrstInI5wq81YRjkOu3kJ
MHvpuCkU45yOKkEl6zTQksAOSi/V35Pi8+LZtl1CFOI3QDKpOvHwKvdDLL0U6eVas3NiSlbHa5xq
uSggWlzthoE8I16WAEVICSDQtfpMm+n9i2fIlLPj1i1x71BcRH60salO9ZFcJid1yAjs3gXJsuzp
gxWZbunZFSOYAwSnptappFiuNMi6AukW3BO8RxjqXuFGxDVfo5EkIoZ9Y1HINyLOT25IPTeP3KGp
LXW/pWw/E1LBv8OxPa6/zj+VyfFE353pwThuOOLi0OHIm86yT8xOLF6B4rpdykCUiS5rzkFHCF4Q
JjWLPLINYnf0htJfjcoutXwttUox1FGZCciMt2QeTChSpPf04yVA19x5aWu2w7PP5CaBrEME2YwY
bptgzXvc56syFtXPjjw/2zMUd1yjarNQVcV4PQux53+KVJQRVxad0jk3tWM2xKIlXe1W0ldfzN6u
6UMVX9d2JpcehW1QZoAFkj4Pe5q6+Lzg4uBEOV3Tf1IjAe4O9GYmFvvjwzo9wcxm/fll6hfeNAvV
H7Ul4jwz2+Jnaq48HCKQML3Ut+q/2mSCgGq33Kq0jC8z5+ftf5Pz4Isvb7zoy71EruEaGtp3VPSr
fxaBuHtQcGQtdIWCyDKMYAP0HtZKhmku6WvmBA2v3IB3QlUc+yoDJ+U1y+mKQtfC6RnHijVPIgZd
4RhdBi++Yo5+r57wJJUWL4z4N3J++n/9LhrhxBvhb7nT5zNfJT/Uy2wGJ5++sQvYQnNsdrQk8fTm
BbSnGXnElxwICMcqg4a7R+PnvsJj+7400PlUU5KNpOdxfTi8L1O6kX0e3eYVbxkktTwxG5F+Lv6G
O3Z8+oqTr4tSU8G+ekjfqEG32REmrfNp72yLLWilRDcZL2REPWJtwq9qjsXI9GKv3XTTb2rDKtUB
tfZhaXIZe49OW5qC7SRSY4HhLb7EYaqqGHbIhoYt/OfSlfOcWvHvWIVQ9+YfDp2Z7evnIlbz/mo4
HAs3B1iXJcXZHXIKz8niMbxwbrQDqCZhySKJLqiEYUQGszO+o31JJ6crKno0bTZ8AtLj6AsYZfsR
1pJwUvFbMWQjSgtAUHJ5jl6Uf6FZkudSoDbGLWyQiVsVFLCPij2LaiYsQQx6ucdzzEpuQW5dh/xO
wDRlxuTmv5jdN/x6KwSOZi/RBvsIhBUO1R1RdWfiYYuKn8w73pY+qEThVfr0A3CnbHfhOUuwlZ4T
aoVeCqtsZZg98ZyNMT/f8I5dIEyu2QQ5xsd14la9d0cxnUZGpsS+nHahOzUh924x4igROa6vXeu+
Gl9O2RBwMh1BAw0RNRLp9QNRtSbVFzJVqfPk7T0DqrShB8TkpxM23Bq2nxW0/e2vNMW943d9PrI9
zyj0b9hZD24OsUrJqRd7Q2TdUha1krbW2xpdYKbPhbCYtOP2G/2tsewxEAu+7kuTf1m6KHeHLh4E
JxgIYR4AyTdnVYXCOR2bmu+0OGtyxTK9b1prtMavn4mCM5FO5E6OWZk9Nta16u+dXfQ+i+kl3oMU
CIlskoNkopA8V7EkRcbs7gpdq3+3FzSfySD3JAauYbmRuk2Q3Ro8Sji25DSTxGCbOv4KT5dZFZ55
WU75RFolLXHZKafzmHXIvvsQy9oLF7lwkkRDbesggeg1KIwds2vcoA/PxrlJVa3j56vHEQzWQ7Wf
qX0qoas3ZdPdGqEP0nW5fXCiKKP6YHslrdLchIKrvy2Qx+npRVzwD9fzdmwLmOkFEnIsRp5inZDw
HR9fTkXnEIlQezOmQjR2pToganTyMlNCzUf0hOzvv+Je11Jsw415qcg030xV26p4fkL1ibuPjEn6
BENp3ThrB8EDH4+TkF+c9QAmjg2epL1irh0qdnWLWq/yfVnNayeFNSgUf2/zkknW+oC/DaJlXSg0
XFl4v8LFi8ZNCE5LSdkigZyTC1fRxzG5sXDfQa93q/ivhSTIi30ZHpDbsYzic4PQoJaujSyweaT7
ynWaRGwrDmW9Ttl9gsyBFkT5l+4B7jmf7qeytsPGylaOkftL1IHG3gZiZqEWBadD+4nMTYfuCMyu
XofCy9hUKoud8q+I7OlU5bocF04WPjF7SOD7dHiL0Ez8Y2h7bwy67c93WHg68GWIXz806YK3y+KN
MrtXkY6wx/MmPR8s+k60tsv4cgMPpeoxGJQzw6da8po7zBQa07cho9oV1vWVaei9MtFZqSEYd3T4
M2TMfXziS/mFi3c/KiwS4RSC6KVXLu7m3s/Cv7YbYcJZYOfUrJMaF3XPeP2trsoReropKbjPuw4B
uH9K+FEntqsWJsUIrV0pf6uBhDZ5aHz97DSmNf2OpTa2x3bWYUDOpBpOnObIzgV/+4KVEkROQDpC
ySfLRFC6LgBdqGYBaQaIbcH0tqWBKVr7w/Vd47KUXC++Bx1drif1xhUM25yjrQmE4fA4proyv3Vb
/g9lvZTke/RbM7NrtY0Ywev67v8p24WXQJtOWwykQHXxl1o6cWdxQWZ0utds9x/1VRwhlObqXLCB
Nm++UyLKH2jSKRZ0cu+sW5AfAyVfbDFzCm8kUrZS4uA52q5lWbystbmGeYax4YcepiIAlinFL36O
8a52WgTCbVcJ5bQiAvM9/QBtkjTR77v/uxBcFww4lVmex8Nisglh0PN0Fkh9nG5eLXvjIjGqmJbx
XfwjQafUQG41HOoUD3qrDGQBpDQtZm9ZcNBUV97787BksFqUUII3P+zoa2pVjsm6vRm8qAa6m5MB
XHuKWz5bAjUhFosHpoexJQKozRYZ8B7pj1fwPqrJlF25UjxSBZFuyuyB16Uosuw5NIIUjVxi8Es/
Q0xcH+iCJqv5SOwZi3fbrbrwAiXv7EZHkxPMz82lQ0ZYeYiNT9WUQeRg87il/hUn2MUJlrKMGesi
0cjMI/chvqiO7srvTvBcYD67rHUfj9kTTbsy3bTNG9RkoTnhN8Yg/FSDrKfk2U+sFe5WB6t0M6W3
Na8nsKENxT8fukY3l7mYP654OD5ncdIE2eCMUJNf6vRq6/degiJ51lDD/pB+cApQgRK+w+RDe9T1
g0JG4zUmA+ZTnxUO6KpmOxiiq1l+t5lVKKo6Wclht3I+9c1Bo4GnJo8sXRpCdC4dwaYI27hocdDH
N2Mamck1v0jByeWhGpavGaiNbcAeoi+Ko+YKeRqv8azeCgxVM0EcVlBUeNSyNh3RweA5yV1apMYM
kTo/FO2ArltDh5h4vhZMZ+YIeD86L8Iq09e/bU7nLj7tgO3nN/v01NvBTGRKWpWyKxopogKOX0Pu
OZ0nowO0iKtpTxrghU54eLbRYgXumHuZBqkhhxdxi0I5y11CZzlT6oZuofMt0odhnBhzczTc2j1l
eXPbxTiNBI4uLDQZeDw//w0WuhIIqnufLw2lUsW53HvTKhoFC41O1hDhXrq3VwgPMKr4ZGDQ2Cdq
6QKcCtXrbX7hLoZQkulpwgCZNeur0sICLjilFW4g4Igf+0p/0T1jMXeTWnHuexFr6HDcqdE0QHRj
aRWhV2BwLIbn/MTcv478TP65a8gpGI+dR8f5wvXL+L2NmtuQY+1wopJLVO7uqRplKCSv08Yap10U
NIqCiqj86vAtXiPMuHWRTuOW2MOUxJyjQ3vSQP9uNSS7YCXY/A7SkGXgvnJ5sabsm0AWOgdM7pvO
j9dnvXUfwy/rNR51wM8Z9RogXE90etyM6NLt7yyXiRwgK+NktMPuSZngoeJnBBEjf7Zh0thPMs2F
3THqNwQyn9f3BltqQflVjeT5GEOWKq7l25NIjfidtGBFiBDWMRRI7MilQLry7GGIugzCP3cQE6FY
XR+DXP11JnS+tDsV0MdjjHVM4HDEFDx3NfgD9BVnm9r5hRIMn7qS890f+t1fORx3M6toxseIXxi2
HrisnFn0WzGUeBn1hCRQFK+eq/Yw7JDsxmBz6E7VEyex4a4pACD7L9HRS+nN4MIziCbghOynYQyO
lQn+J2CBJXsD/M8PVAPFZND4RY2iPMIUtGkN9i93RJEu3qGdNmYg09JlBlX7QxlySanUyaUpamRW
XLCiGrMhMgH8JITc6jJjCbV9V5yAbZ3JOI+bxnel+qY4iMb8oVYDV6nQHXm8tMeYdGiY35KJcPgU
i2gAadqCZCTqUyZDsVRxvYgJny75nOQ/SGfcFQ+DiSaiDs/jgQ5oAIyfYk04xPh42GeyEiIxWS/r
52NgaENQGpYXo9C1CBL2YDlDo2hvCj2MCM5GZcFaQFnesIcPVnrD9tOch44maYPaP0rUhmex6n0O
PImQKmbecInkazBTyxPOyWMlR5P/nafFzN1YwyTRd6XMNQO4bEQX1j2hzTyxZfQC9clXXEUvuLuH
6UJy2nLbKOFaQVzexVRH21ujLaW0YFFVGuTLxOmNkdCBMymo0VrZo+zOv4+S1KeP/cKP+8ZkRek/
sGEibK5HvihTinsuACAz20pbnYm5ECw+MnjLASkQSndlUlfXA6uyS+9z0CNfnTItzXVMtc9iF97C
7+yZkoDL0aJc+HNqPnhDa9fWn1Aj1ZQdU/H4g5KGzJn8Qki9d777EQpTKOnPH41EsDuc9tGPHtjT
sPwVKepYE7i0XxoGE4KkqCyZTJ0VKC+TT9XW6IMJhJUxYaLzSu4pclZXFjqVk6hqyY8k49Sev4cP
V/NW9Z8Bqybaa6jbYall61013zwvryceFQ+YAoeoqFBAo4HLiYBlaGqj3cIsfukO7fjPRcw6yLvs
M6/OUfFtWNTz0kugCpLYOECSMmh/BamNlvpqZZ4tn+KZaiqJJn7GxXFaiM1wYH5Yau+uDe+j5rQr
wiOueIAy03fC7MgvDIHNzLByWGuU+N4B+SsERddsXEBMGTxeT+iSkkTQTIPEunHsUfhAOXGh1e6a
s230y/qPrUNiwHzL0OXST1Lgh4f5jInKdmei959YvQ4WOxsvpPr3k4XMxDM8xMr4icCpSRcheeCu
gYh6QLI+Dnf/nLMm2zRmbCnO8DvyXheWY9d25+HCCpSGkUcXPu1g5F0FAfUzYkwy1nYhelAK+sWt
8DMVMWomC/WvGOPsXJFKASgNdnBbD4aX/WmSbKtoUOql/lzfQvQF13KBmB76NmtpNTTi3HIFCGSc
7OkI/ff/mITbGErigxGC+37covIUuhV3s65q9MGLClQIHyuzko0CZgSck7MYgWcSDG9T06zWO1U2
JeAIARK4fYe4M0CFKPUc53EC/0uGjhPM6N25OVhGFZd0e93v130PdTOidpf5CbzzUSJw1tWfSfBZ
OKjVcYT9LmfkShQg+CoOaxDWePzyPA5EoEY6J9/1/YRp7wTDB+XZFyzXDYQvqUXh7iPggvnIzLDG
MOmmURJ9UdI3YG5PHAf4c95HWMFt44hXzCtLfS75XrH+CnwjtIBR8e2e6yKpuUNBOyhaK0VM1ZG3
WGgEKH9u9poNolRoOH5+rQfwwW04P9fL4uS/EMKtW1RP/BvClUXKk8vVkuSRGw7MfH+ViT3FrKeQ
l18ToYjujVHPhPaDisXgt7WO0e0MTX/X/Twk483DH3NjhD9d8pmOvkFXRk9Qsd2Jcu8AyXbX6kwi
TjICTPagpAawOt2cOeVmz3c566vBKaPrVkpQiwBqUqzV4jP/eBkpSnq/V99aqn9MS9fQSYYcz2HV
5waR4yh+ZnbifJpJkd3+ehOj26/rEe0dTFUd14LqqNwYMJNfU5I92lhxU13ybxar71hPrA3x68m3
TGLnOfow2oVNlG3seJmsYCJxla5x1SQP/BLD4xD3eIheuG3v57ftiUSrRVfmcvlR6J4DdH7xcJlf
InD3nRUYRlzWozHZx248GOSiHvq5SVMQqrQ0N6bahL3dgu1ctL/k8XeVDiOuEOqeyKRxrSQNtK1C
1kOCRTEXVFLdkq7IZPGlSp8Gm6rHCGRSrlhBYyCBY2Fp5mbJ7NvvDAIgPc7lxhH/holaiTTY+Puc
tRa/2ND25KrPg0urbmkpzDDUJKrOK0Wf1q/iYQGh8uv+85x2ZsQ6NWAh2O6msrNQ8klm7v9az3T2
+a9qg3rjilEdKhkDoBsIbUqyH336QtD0VBzXUStmVpwspv5OCkW1b9BOz8Q5+acXNIgV1dVPud6M
CoHVVOdMIej0wQJwrJnp7H5PDQThuaLMYGiiSoCp/E1t4ATF5AEPBPlxOl/6LL9Ln0RVBOXwilU+
knEhvxA7ebdFbXND3dNTX+i7vMZVpQr7klxXH6UP5nSaPpbqhPh6CyxtUtdt09SYa6Q2+P41/OGH
JqBSjvSS69qRWpygLTT7TEJQ283nPZm0f8XgO9lN6gSjrSdjfqZKWB2LTnSdGXEfGhMMcipNqhf1
iitV4D3KDB3FVATJzyvUqRsVX0MJbwGgEpxOOAgnABnOhgEA0KGBUvaNx33zwDry9sP3B3gDEYxO
v9O6YR2xUGyyUZipp1yjXVy2BVyMOA3FG9UMVPKF0Y1GDMH0s6hfnS250c4ahSGvSYyMyeJbAoAi
ZYEotOe8cNUEw0ipE+AXPcNWp4f0uC7/mXW1z13LdqSoilgCQWqbV3S/e2IHOuPafpbAX1X/BYjP
gdkcwypr+jAy7SfXBapVdxe517kJ1J4TWvltD7a9DX8WXvnGTK7JwtQe2SEMdrbYLzMZON+Jjfrk
8N97aqptoLttoORU6bBe4QO2Q2C6ecAuSHc1JQPXDLsoCOX0VGG2sRlKQ+Lux0vKB7L7NGiTXOuu
1n7wRMPu9oUggYfanJExOZu+Ul7pnN7R0Ks7hFKO0WdxSmDRhD7pW7MKjE806zxtR2d6BW9r7y2D
7CREL6da33NgKCQ74HNJF/tR4UZoxkdyh2KO6RUjuh8J52xTqg/vp4JTHm6vYgMe/9h1EldRsyBm
3nTc3of/GRTnbXmuNPNEEgBVZ2DxKXYq7GiSRd93tvG4RZEIgCRitkgcpRiG7NHUcLNY7nBh7baX
XDjaFpPgPfqvdp46MTvOz4NTKCLRu4uedQHGkNBSg0ZQnYW7nOzTyBz417k/d53JKYlO4EJS+1VC
IkByxR3cZS3tTn09y5FWWWisBs0hMsgQOyqjlR33pxjUcm5gT9gphaI7c2XWbYMXvW0zbF5xlehA
7NG7PC0h1r9sXv2SvmYy/57rru8M5+Se/4AXwuWQZxqwDxMG1jCq1KXjx/IPO7O/XVgJ5Vx1U3nX
hntwWIsoy2FmKIg4LuLq2h7T4DsaS4nyUc3mksTxMNp434RmNeIZliSCnJnscm3Dj0axkdJqnG2p
0WczQ/G4di8Be5zB5tG/VZQWc8sBypsrJn4acdgI2qS78zogHdCrcu4bLENk9OhYIHeQSJZXn45N
GUz7CCEEpUDIGgVOFa7x1DdxCaL1rU3b0980GK3Qt3Jw9d4c1bRxyyvQhwNQuHHcuJk/lCKyZTDN
/tgmQ3TsgxayAJ400RMup78uDIkiu0uLBt3+ZtciE/O0yrN+qAFCD/Od1sqT0MpY8srEKGhTPYH8
RUKDvc/yWOoPmOkXJ9ivDr0chjnMKCJbY/d6PhdWrqgW8A3rTcAf4rBwEUEaJHF5NOkrtptz1bhI
CqxWP4MviBIgsbgcbXOi1ki/93O4wGvB1H5BK2wqad9stFo4AJr4oC13p+jOp4puWqxwJKy47W7z
LeTPdkDi82pqzLOTSf8ZV2LaTijeKtFYvqLHssCAj4nWKu2+6JR6Km0CtuuaWq8w1WKdCDS9xbUU
jgmpCtkGvpc1QujcfKzPz2j7NPDLeTlsgx1sxN9abJCjBXOuWXklLb7dtozrkXJeNBJqN54jSyUI
JJbG4KmODifGoSGCSi7GWzXvdCGrI5jv4U07abporE/cPpVQAShQQnjCz1QWUsxaKFvidJJ80ALn
6pVX/rX/+vCLrrNp1WIP9dTTeJef7sP6GAgsPdXtGy/x/rDjzVH2tRtVcQ9zUcC6B5ncokSx/HpO
/y+c5dHFDmfAYcohASmMjiTlvlF2UmqSEvKDUpNBsBkTcTfuFE7u17kOiamWc3LllhLjBIL8yw7v
U47LWxQfPHXHtjodPqweYzEHV9ntDyQSxqnTNhTpcxUKNN4A6wfmIoNxZdIdHJDRO/tfoVeHVtyk
Wk1SmNIViPcXNRY9OkFuL5IJsxEvGQO6WujJIPPCfVY4C28F+nJhE0GAsYIowhFNyRZeyIVp7ynr
9+Xg2sVWq6UtxKC6AFHjllFf36ZQM9pF+7yL87mpibLMpt0RjtD3Duak9wirv/iCqzsPKUPsSL/j
a5DL6NUwqtqDSEVSrdMHBykzOoA0YQCa8SyKaa9ryE0rp97fJVI0AyUo8piVsuNWILKWKoklQBQC
RKk88Pu7o+592lCbN4hA3gsXnhYD0vPZ0TU50SUBnwO5C67MS9HVbEZSSObsdLrn9/GyqLqOLyIm
a33/yEfsiy56Zgkz/pZhjIUyu8S5QkaoTX9QXDzJnx9oqio42dvh8MhXzp8YrnwjhIP+wUgCzZAk
tDGe4PGXsnFOu0p5U4hTU8+zvK7Sfk2xAHUbC7buTs+HmxlHL+85vCGz+ecv1z0Qi3FGzeFlPSiN
Vle0tDjUrBZ0rul+yh9EtqVTCgWDWVyLDVqq7cQaplTLDiaS90QD6KRQF+O2DHni4h1Txfd5dpCy
d0gCl8fqerRlcRO8R+ziXSEBxe7hDpL9gBpQCUO3wLYYJWTiCNQ+gVyiVTDRnTV9JbXxyydpq/kO
QlGrjs4NUOOQd+LNrHmJ37Bim1Ksv4CmGaOweHCM2ANZ8Djex/scTRr6FR/SgaOtYPRE+tgXOj9B
NhK0cT3710CT8uHNigBoZZvpmFF4LIA1Ro8Q4f5jsoJXB67zlaanpL1cQBylzUoHul8okJEjurS3
NWNewcuZE1kd/2tMa06ZBStHJ5pI/yoBbahecKSwEoXHqKNtUqEcDnUX6ehRy0iMW4/NUyKhmwod
BqcaoIuUvx/ceXcfJEH7uT5VRa/8aIHI65P81qL4liZscF9ChDUBAbgGPFr1ZeWWRGfQsMLlaPb5
K7SBHbgaIRoq0TrM5m3Y225hHnUgTV9mOaKeNAVY1LVNpeaKzOun2mPozhUVZodcqKkIdLrNb94L
vvVyQ9bBira7O48ZeFcaDK8xXkzrP3FA/5wZWi2WIFyrsFavN31zRP5vz+fFNWfp8BtaC9mw+o4m
DlfyY+iejB6IGOVTY5oxtGutiwmznznBcgCQpgCMVnIyP5CGBtaqM1ad7t9oL3Sm6DQd8f08KlqU
v3IqpG6cmcZIXz2H+CycqqMmpUJxTsdo017sqW3AnJAg9wZOTkMu16EzG+EIIzBAVMj/1+uc384O
Iu9XKnX/4xvOCQOPfZtmclEDoNm3r0WV8i657TLX5zXAcroJtzJWL+1mshHj5F7Drtq2de8AU+fx
bHHlcpJavAx+tR0kID8+8aixYFNzyqUp1DGcnmIAstWYviYb6XyUiOZYbqNmyxVGwP+Cr5c4dfLm
37ne5ZZfAlwyV7OqNp/HUvI1wyjfH0xvKAjgM+WMcmr26A3YBtVUx4boQ70LDVUwdDJ2BziJTLRW
XRMRX67XYC6VbnBo4+jNwVJ01WquGi+Z9bveuCiZXyUNs3CHQXIqY+xWe/31ynSTNLqkTYY3M5rG
BkD1Q1O/XUUWUVAOcQOxKPXapRGfyqFKFRLJs88A427O7lcmA87tv40yt2kpqZI4iq+26oL/ziRt
7wGXJmaHKeJBR8JaKc6oR4by0jXmSRHMT99G4CXjytWTJTOEzP/XSVNEqZpvhRb9KsDw7PBr0jeg
aWdNchN5R5y6LxydbxIpqc+zVHCxsfnEBPDVQHdKTtVrH27TRJJNhi3FL2p60t76hfASqYEtUTfe
qwg9accrV8srUgVUg2TbtPTwc2rbK3mopnkFtHWTYAXG1QExcV41ndgVl+WwZtfJkhEAUkpvLLq6
rUmMKQ9svZjohA9CAa4+Hl3Z+asIYH0dnsWLAFm7j/YdLfxLTtjyHHK6D9bpJuJUHeMe9+8UIvSW
0jCc10c146nbXGbZpTUhTwLsDa+F3U8+H3uIUOtTUTpXknaSMv8WxAbmNYeyTQT+hUhqCKLdatlC
zK8ODYEN9v1M2gyAc/dP8yVUIz2kfjAonbv4fTYqCR6pA95ZW4zlSAdBN6+v07OCJHOKqq4BCy8T
yedJnHJli3DctTLB8pwelFVEO/EFuhld1IIpQPXCgjNcZew1XlsrZOlk5Bib1yswtQHjUnaP/w00
zcYAQspW2mt0SWDYpAmRBpNxc6GfKsedxc3hzOvI1jgkz8JC6+BRYQlKWVrETD8KwQLgwVIwkPOL
LrkZ167vETwpIZF1OkBD7c2QUGfo+ayoqRfFGgGMTKx+y71eGTloiCvityA/SgetiIwgANJccOHH
Vwx33DHFVv5JTp4OZ+hheGzvupbQJq5XEStVFfcfe/s/uyXXTYHyqcZKitoUeYNd+iuOpdVMS/5M
4IuPvFsxPYNAk0TEJEBQ0AR8c7soOx+F8zDJeGNG2wafCo+qIA5FgS75bhGY/8rwZcpFPiKSYiuR
D842jjwivEHlxJvICY5lxMiEITozdsN9WgTFJsmDXE3L91LhXMhzqpHou/htZzIC1Wrqha2n1vYx
X4GMp+R7P+vnsEGzeTZjQBFl82OjT8UbogTR621DlotHPCym/NRfZ26HCyo1peY50tUOOGOdaRNH
uDnQ1tOrZHkGjZEEWTJH4LQHRGkrVO1iz3dpEenmQ8X8VClkZmnf3zVZ6dKv8qyBaV4xcgZ07PPd
rgEskE8fFcRK5FA1u09weCv8ooLF4QC+/PNQYzPfn2UpfD/ZL9VJ+B5RjsfutX29Q7iMj4j2ea/S
upRXIpaRuM0yFxn7a6OMtHYeaMC+1Cx6jGJYe9lkA9FqO9fSOHF3hROjfR/JEMD7YDAv5ruPBv0y
zUV22ZEdXcSuLhigMabf7qMacCVcR4tABcy6KvfDNDqQLwWaOaBm30RskZ5+kl8qUeMMO0RpuFuv
5+w2+a+LaR6VAhaWmM7zPFZtp15UHzv0nao9xvE2zjmo0r1EX0QxAqzQmdJ4rNh55c+DO6T3431s
3VWoW7xLz5AOAuAC/s8OhYWnlfuq7cebcl17g1yWXcHDXkChgB/+q/+EfzYH2kYGA4OmjnXBYQTr
2UKrWAWFHRJIzycsFMpLsrSaNmPubXkdWZGEDo170GqLLuse8kmU17vP2azsSht+ZDsa2bSnyrFw
alg/5lYV7Q9V4a8++Eh85tpteEdKjO+wBh2389Cmn2R3qBJuoknuw4EAHCBkZjavKbv6+WD6f22O
fMUEWLfZ0NEiAdenFaXs0hciTz6FqxBNbiL205RPad+BTA2jomx7FBecJjWAE1YVUs74+oYBfnqf
wc2dZcUEEF25YHIpMwst716JajkP3L7wgvrm1jvhT0gPqZ+Jj4RCsnbS2noJp1mcybIQadW8tRzX
QxFzaUevytv6vTGyme0GBS0kB/Umg7hkiX+842RoUsIh1WL8mBmlp9l3VEKBJaBKfy5KT1DXquOl
wg+5rLsA8ATQfCRC8RulVJvmxKPIBrOy9SBpjcZ2BA8Tgzstu4He1oIXUr+B4FOpMwaCCZQP39pf
AAeYF/YP08GVsJElER9+DlRWOa5HbWIgiGvfyDtKqbTMseg+oN/+vRznePE5R7YnnIuvp3o0zKeW
syfJh6IHcHVctWvcj1kTj+O4Gjr4pMY/Kxe+GdluqEvN6Ojhy8UUkCczJQ9owyXlUMDfRINzD+Db
qt2fIKOTeI5o+5dTbz/Rf600Ls9rGNPygXtIc3jFw6duulTPdfH5vcvP+8K4fzNlUq8S908WYb9R
Tmxxlumqs0NBv/frbuZKXBlEr3EUrWV9roJf9nETST+pu9M2pzOBnSAw7hdC9O9fk2XUNTfAd2Wr
qRyhXaGQBIs1qG0VB45A/ndOoo/jO5G5q9uuEcRn/Q2yoR6IQcsUROWYNLS0VdIXR/52IsG/dTCQ
zNZYmpPhC/aoaGHRxNNTYXq/Zzhu7XoHO+6aSuhOgD90+bvk8Q0yyjYod1gsCtCJS1h2mBKrBZ5X
VfNCIP3JhS8B5s1+zgl5OItkQ0UNJP8BlF5UQqhAXhXIKTyFn4gNHv8fyF2CVqOFbvPvukfC/R4k
dDUuxDZrEyVY+uRu+EitSgqQimzlhgXJ2EIzRPLT7Yb8HI8kWVmBIUT5A7C+6xlSgeRPVwUbxeqd
6xPrAxLcqcPcLFsH0RNAoo64gY0EH197Gh3YQ4epeNXG50duwFz7eZpF3vsUe2OxO4/BbSRzFEWE
q/oLmcUjxG09u55tefZX155wYR2Zj+N8UAGkuUGd7oXYx1OxRdkWDorxwl9iBB6TaeLsHnxad508
dKW0CCXe4rBhAIoMxxUXaZmDegS73AXybToEf0yEYxeld/R7uVlSKL1bCVotbcFqKsEeOFA3u8Xv
1fFC1zUS3qaAREj2rWIuRcR9jrBqsyqNhEKFVHA8vrLD6c48xVoUUymvGF6Mv9rnuvFTUaD0RHwx
jMo7toyVJDBkKmHZ+zTfUS+VvY/7Daz3Js0tGAJMAKHmIn6hPuNbHlb8s3/6hZ+P5aLney9AXy4O
ktnjNevbYa6qB6BvS8aXZ9ksQuWnJ1DXbZvRL2Wtbh9ADtcPi1UpNx73mn+ALZbncTzJNZjbNqg/
Rl6EqwID5Hg+TTzsFKmVFdZUqJoRSNkahn44CaIdJJlpwSF1pF3TQd/D8xxj1LttK5mzSaBS3I5C
PZNU4PRkBHltvjiuTPdR4IKmZFHEeNDwr3Xi+eR/nZb7eizq/JngZX154ACu7GYxDCm/VFSX0ExO
Ctq55iHJCFamUhDW7FXq18dbkmw36B3ChWCDd07yuLBnzAKh53YYVCdXylWHzeIN0oslg+J0FT53
kx1kzciinCfC0983A24TU9+OGs4pw3HYln1Ig6m1NxLBSHEYND+DZ+nDOgJO2BH5SxWAz1G+O3Dg
RvwVlKRAjKccb7kBFYBRUDaPgnN0P1EBmVgLLSM99UUKi0oq3pY4uNs/ABoHuavkU2/BTaKPrt9H
fOnXhySsECGZBlBlvhrwoSpQoEmZt47FLmwaO0M3ZmqxSEiJ8iqRug7PFdyfai8KcqNTc+dqXabH
ERV0wyj0ClL/w4k1R90jcB3JgXOQiNGr7A/YBIsoRPIwefIP7f0zVluUvCucPt2lP5yhAnPjKo5U
zTMKq7e1PiQkKvpodUN63Wd+OLiD1lTsoj3Uk7D7RyVyDClq+grzDQBvdjkjkvCpJYPcuJlaGury
zwQon8sVC5liN2dkI5wbobyQA0NXdh6CHad0g0jEBZCGG8tqqDmUZz2Nm/Z29OKF9dZzTE9VlCdB
hgCiRReGmdQsGYILbeSKvoIFxjE4BA1yv3FDmW7nD0VkHVjHPxUXfgW347Z1/u0Z9xvmBqdX4YAS
R8YxoJHmVRu4w4vVjTkNmDpmmaL6RvObde+0eG3xVl3qz7vfZJ/dbcR6eoztbSaN/ta8vGythUT0
8JO0ZWP/cog7AiCPOoCQuQffbDuKXNgUf/eUipsIxqQCuMrtYqDjK8zJxp+Phma9fVcAV5WuxI1d
tKK+M52NmsVn58psS66Cr/YRok8pZ1ur5VQPoCDyzzZA4bz+Njz2r0wOkSYoBDK2zIECFOs65xyw
vj/vBQdu+Z226BJeZn1VZUebW+BAjhsNiJ25EmmdckBDHu3+lG1VxUUVCRukZ9BVhIZpAKeeaXkS
wP68Z/9lEnvX7xYk+1jDqA+7xLlg08lgVts6ntRd5VXCASDiNotrA8mY3w2PlfNZXispYvh3g6hZ
iQbJBw0KcAiuLa9wdGBb6alw811hM4a9L+ymvfp623QIkhGl4BoXJM2rnnAi+fEKSFuV0NcN1lCf
oUnm+EsFlG9HoqtTOmBBEMnUYpeM+KG6/MR0vSzkkMJd4bGH17fZOUX96mk05Jt3gk9fPcG3C+7i
ZmRweCPzZSbPUKQwAE6IN8PKsogP2dcteOlTb4cOpYgFQ+NVPCW46yFIsP3JMK4gVWtzrWVJfKT6
D0T/QrTTHJP5/TNnmejED4uDJCjZbXPEwy3VvU/Z3CPDpwrpbl6xVA5ruKQn3xXfyzLm9UI3aYzs
qz/gPXWT54qWRZtmf4v7vBNSRwLAtSUbHtDZ4nMN8f0WDQdQ+aoeU8nzSuIIK+VTgoiz7gTyskYE
2Jh7DU0cJm8kEHdxsGBD2NZX9SZLcTBdxxIyE4tz5wxaoAktpcxQj51PIUmlEJtwu2CDKbuGq7iC
9dvYe3RcBy99rh6SZFTIvPqp1TXROYNPXDEnMObuuRerrP0HdUnFgHa6vfHh9ZZJaNf8AOqwOK0p
gVn6QuLuEUCDQx9qrPnUS7Os1VTPKuohMxA+IVZtjC8249NspTNeo5n2QiRRfh/Q2fDpe/O+cabH
BDGtanQkWZ/qPnASxuPAHU9nq+Ke047HFCgAbbygGlEtp28VMFf+TksWhpTjjdLec9xcj/kM8Wki
zW58iuuopPpGm7g9FkiTJh4s9NFD+bGaLhNbi15cAahg+aipbfBktE7+KgJCJMnxj18OkjDdRylE
gun2OOWZ6jBkDGLxIu1LuXkDAVZXu6dvLIy16Q/c4rmwsNwWaxKJpk334E3CYkzFdTvsPXMEH2oq
KTCXjlf2shZ7R7XAj0RadcD8WhpY8NaZ+G17sCnI6DxDUgnwQdr6fgsyfB/nHDG7v/i0VPn6uGMo
eWzdCeuAag/AQHUfb8mE+2u/L85iiagvu4cYy8CYlYxHBMh7EUF1e8U2WPN03MoDdouLqutuvWuq
KRqK73K326wPKMrmAjDR4q6rC8lFikvmryTf0HgT7B+IzU0bO5pKlY7NIsDtugCczWLrL9xwCn4L
VrmIeQhkM+ihmv4pU5hleHkRLWOOa1+kmnMxyPTySsXKEHfZMbmacsTAeEvcobcbCUzQ3cR124k9
YShkpIqQggq7DJaBmV2k68ftpgtvmJ3JS0vc07Hk9Lv+EkSJCBAYfGP8b6XDhM+bzhK43erpa8O/
rSzjr/YxBLB5K/mxdWAgol2xlwqyLQNWmTzRNOZmksCP8PfQDvkEbNKgzHyzyhz/sx0JSFP0aTYG
rFvPHLV1cB04c2l4m6MeuSTv/5I80jkviK1YcFotFsdnWrNTehdWRJTsFLAwJlD9EgQ32yTscsoL
D3tbEYlAKYskEQcPbpagEBGEGYCKADQMpGLY40TnpFCu6nmebfFSwWaeDZTPBzK11WUVAAfuWJaP
Zo1TZVYrgvajb6m7qKGLVw7ERgTaDeCoEu0aJNatpbF4g2TxXbGEquOoUSxIP98mw24IsBdPrWe9
4X/fq8HlTn7vqrk4caHCXkl8B5hDctWgLBKqXCUEeTXSRQtOYpZgwfYmc6t08YC3qq2PckmzJcXq
bMYARbAyKIjMGRupOplP+DFXW2/Oeg10J2LvRfyFgr8XK0IeAQmbdm6nTMD5Cf0+WZRmpI8nZak/
LRllpK7O5JV7gjlFKlK5qhTr/sm9z3kF5AMqPCpb0L9qD2bIDEHzd2+oGaOsoChtrKs7xYEgkL0H
u0U8fE0b2QnDO3vLngBiZcR/o9PLHiJeY59EfylyQ1xp348ng0ODKXReoXhxm4ALD+0V0ibwBKaj
NV+I4Kktqku1rOCIBUvYT5WeCK1ThDGxh8rUNf0ZcljHYpjoPlKe6zQvxkZ2IkwIZmnFlLeYYUwt
n5JjZ6q8CoqM2sflkdOK3PRHvhcH3u0239eI9+VY5Mb5eOVkcTlikHEtX+Jry2+4ofScK1tv/G6K
aW6F9kmARkIIc5qvD2yNVc+L46IlKiPm9/b2HLha0S6EDCcATjEvWpCQpYVsKvYR1/TrnqaEf8s3
t5i3Vjr/pACxCLK7z0r3gTwrMM8CYHpMf1CiVZjlTb+camWx+F9N8mEqqqWby0fXJdk5tAueIlvk
k8JnrSfd5QqE58JM9NN7OkLB73roNMmRQDNFt4h24y2gT5gLj569dNf5yExJ+dzhaLrumTe5ajbP
2ZHBNN6jRFeNnnlNYj8bdbOmoL1XRt1pHrdL1Ts42Jsdxp/k9BjKjQixMmuS4FuYaQuKJfPLjx0G
3muI33Tki7y2olCfDbqWEXweu4hGzIbvplC7mVF49ueYsdtESlEzIa8uKvDIqm0l/8MJgsnw78mL
DdhES9nf+Kh8QYX46GxrwAvT/EtlHLZtLtT1ip7iMHUqd/ihZV6VXEkfS7Fk3NN09BsqPRmz7U9F
ngT/pWz09evwn8tduleDhYs+YbacoiaQSEwcMANI6jlyDxfPYmKYMrkOuvLi0lLIykVL9m+ztxII
P+4m2dhgng3/FK7M5jUl1NlWoUCWpI/MF2wclhBqFjqEY9t0hEvhUzoI5F4/7f12fgEkiAjoXyp+
nDNVLiLZgdSEhH6luQg2JfdIlwsIKkLyXhgtTvAyumQu2TLGL0CKn/i1rKTDBZ7WqkM+YM9wiTIp
eznuksfuToJDC+6Ki40HhuSwlBqCuT8x62qXuoILJGYZsAIyj/02H03QgelhPgD91kxd7iY+4abV
iJ3IgFi/Q9lgbEsRJPbnMUr/217ExSHMQLWiPN7y3ZYsOrpv0ADQ+3Z1qPnxdB5d2Igh/yqz0XIJ
7+bXzmWLARnMBwa/SU5vDDHtvfRDl/AFfRw492cIyEgUa2g+cqYRHPnnvdRl2CfoXANNr1tNg8aj
h26q2+QRdXuFnrypAXzgEwy0HloA8/8dEnUC/lCulyrmOHUxFBstq3rGZZ4XHh7QYdOmsoLOoi0c
Fb8G6GZ/dFvBLYNRV6cmg5mtMjqHgUM2MnZdWU+dYG/cSF/WpnBnAHxkHBl6M9eYIbWC4A9kOBQv
cSLFGZuPr2E66HnQzRp56CSGCvnOhD+JX4a45BXHFsbZjU6/f/dmh0ywyHBG6744bvUG0LqTNMCC
cMSRpdxdMVcz+Fupz7xDbUb/ggESoz38QbztZ2UkEjTyo3n5EvwVOhHMDifTnQ2Xc4kumI4xgQqZ
XF9RXXtl+T5npjnaJ3Y04MtOZUy1I9O1VsS2/lUa1giEZnaEGFancc5VrNj8lIxcRLxoctVCU1cQ
ZWIt/XrkWfc/Os8LUlE0EABtxVeZufxYcskswrZy3EQF0E1nc/QB5iPu5kNxRVeXrVOv8Js2zeOv
mStjqlyVPZWlm8YHBaqolVjN3ZUQDkXm94E/i0hTDXEBFMwufb6HTsEmn+fF6Hkdar8UgmP8zrt7
9GgNJa3VIqk5NMwAMX5B9LwZDGqTz86qjJI89w+EdRilEu2IMs5RpnzuucVuTgR6VsELS8wCGMDO
iw9ijk2oVZDqZzft2rSCmJNeoD/kDzPSZ5OYMoL43swYRwjRtSleOcN9tme6usiKUiJPh1ioXKxD
hSTdShsIdJd5oqIDtrQnnkODVjlb/7lgQGWTtqzNAB0fPH2eF7+HDMdQlrd+Oyue8IQeC1qhSQsn
Zpl2p1d/P8P1QoschJVd+Wulk5GqV9BtVNtISuhWGh644UNia15MeOvQM7AAH8pArB8Ko/2NPlhk
MhMSiNo9DYK7P8uovop5Y4J1sfbGfC7AojnYdGZ07GfST1iKfTqynRLTcMh4qXZmhdo+WERpFxAf
ZSEWXztJiDHCKO7sSpn+UvhMMb1RX+LedXa7PzSyLOHJompNiFM8XAX3MyUIViHzkDC3yX3y2Z6W
bYkEBGTjUr2MIbVH/iylBZmANlv4m/P6apBvGlHpSgZ+G7h5Qf0BV2pv1dw9wcYkGezxAj1R5OcL
KnDQep1CwHrJSuPApBVhB+ir7ujrOJfcXFQSE6z7mrqs1aUzcqOxymDKjWIM+mh57C0T7M890WJG
m7FnxWVWWNOMVoxD20JOF9C8N3I9wTo4T6ZTd7xN+1XrIbs6sHFZd5iBmt/JfaO7KwJwRMixr53W
Xu3xYDwB6hVpYtK5Jf08DMppcyQHggW8hCa4/SKz2AlTRH4KztOKNQy7869ntMYTER6Nh3Aa74bX
OO8cd0QUh57EpZHYOeTn4cqIZtKeYRXsxQZP6T+wd1Zca7ik8zZazWk48jG1l7n5ahAMRClNqyXX
bv1jDkEAe3Gj/kCRMMNBWJk5SbkKxHJpZderTVxUsjfZS3nSJMf/taLiQmGDQdfdYIq32a1bubNY
5XrrqgbhGsbinPfDsjfQej9A2HpvY4MB/laFNaRAPkLYWeY8kyezyFEP33ivvYVE7kDXtzD1m4qS
VXV5gZ1UCXQ/7Nd50nYVKqbWQafNt3zh0759TYi0q3WIcIPwhA3Zzange2WCvKuKC/Hp6csHWEeA
0EUhu7AoQ4nwUEhwAu9SNtc6PQjUWJqZZd1c/aUHN9m7bIOqcLgaPW/SEOIjB9gs0sy+aaC5Msxc
8CTrW6dLYtWjJXP6F23BPQOwvOBbYHytmtqXoWjWPkdfevTqBrFBlK1E7TZV4JBVd0qKoivJYJpA
C+kr0A/omd7wi/me+2dpDAb2Q3eOULshbue8pQqzG8OXVOvzF0OawbQHW+93Ec8IFEmElfiGamSB
j1kJGch3aF8EZgAnWMLPMW2LtHjOTXwVTg+9rT1OgEDDeX0/NXMmBPafJwA5JSpAl+MKWdY7k01w
jcWXfgltRC2VrQK2WRUw1NHgwoNODICD+v2aOrqJEDkRbEx2VWBVENEuz4schlXTbhUENXtT5COt
jzsTL6ySlsMCig3LJG7PCOza/MswyIxOU2IsbVIubVKbVEtnetx/BCte9954Xnj06emL7eOEdM48
f0eNDtvC3uWoG3uhDqJpuzb16TKNeIMuJyQyvrALZMrM4+BPtH5dREldhYgey1aHyXeIo36+64Bi
ZwRPmdHyHeNDhI27C6tx49xNtUnURJAMfVi2H08xg2yENR6PpDN3m8KS8T6Gsf56/fkA2zjiVZDG
c3ShgqUZAWK4q5V4VKaVQYDIpfbWqB1V4PPokhvzMEMSOdgsu5XF/2x7yExBl4e8zC2E0tmycuIA
UOrg+GV8IoGvKcDcN6sFVYOruk97cN3A5Mt6pTNkNb8nliedR2MYhCGF+mvxyKNDu7VKgnKJUQlo
fPNUZF5q/PDCjX3kUBmvE2DWv5k2ZJ1TGh98FsyjgGeYWMNQoIVSKaBSM9hqZSIOTQenBtqZW7h/
MuZuLlVLXNU+2wX574dksRnUpUjRzXVSUBNTw0TJLeAVKmInVh3dBsKp6ojiy0IeIT95ZMsIjS2Z
orNIgjarsmEbAoZoy6AvqTbK++gTonNh1RVN/NjOLJv4KzVX/EoKopPgJnYvHcxqbCCKDS02Am6v
aVUJb8pnJ6YvipSmcLwPnUOAauFc711GfdJPxaV7MefaqnSHyt30qNHgzhg7nGPBhW1uYELKpPtu
BakVeb7DvpM+6yC8A2X/wqSPYZSaYHzQ8pR7/ZdBlZ/hFwuSB31ZBBTsoG87n7vSzuCQDJ8i7nHr
hRHpoLCpPYXzpy67NQvaaLH+lbVTtnNrvW06O4dhRL7Sbbd8B8aOk5/2yMIgAdzW9y1iqZiKmLBN
SiIijDBTRNTxj1N09LnwHyKIBzy6kewOEizqWPWS9Ghe9k5XsDsn98krzac4ZdqnQaRwuKlozRFC
u6QEDwTrImhubTXOcKt2F3JQg1pcXPNL2rQoXFo/qCsoapnDJ8tXeepDf8LPmxS0BMmp7Wfb8m+U
0g9ywsglzQWTjH1Tx+B9A215sOHxR2us8bKeRN/RzXITqEicQtnFfAhxkj/6qR1TzK3K1OlWKlvI
7010F2hxWticTtfj8kTsxW+9U0F0ulPk8qtAUroQYj2KekKGbzQuwlCI4dLWm1rrni3jWGR6d4/a
jt6415WWkz8E/FT97BQzR23Q/kKaoWCw5CmRHQ/ba65y2yZiaUXioqGd2olyUYlkHeKuDUF/kXB4
jtIh4ZCtDu4+AKua5UAPnwATRN5lW+gzdlkXmmR1hPs/eXIMd5gx7seh/2TsalCEqN3aWmec/ohu
k3itGOgAKWmBmyoeyu7R9rBUZzAPaj4mGZzgtm/sDi3JFJFVS4uSeOA4hT9WhCq5xnHjmf1cvMnO
G2CGN1PMbwzPybDFeFWYQJcdvLyaYHtSnt3Mktg5smwgotd3MklRvL4Nv5DljOs16Sf4U/LVm503
gzfnhf6hBsS62QKF85A4qBJ8xl1F4b2Q/hxMNr+/otw+gFUdEDqi4dyDjyGUR5h0R/huJ1DQLC4F
ktsZcOvsU5pgmCvkrdO1pbynUrkxDJysk+TiBChqYkEtPclmf1Xgd1ocDGTJNrJ/X8UjLKOky5y0
G5H4uHzQ9qmgCt1LZcfhoDgNmp42LltBSB7fB2vQmWyz8JdA5Eg8m2N+RrJSVD8NYQDtff/OKIxm
OlXxiyWx/LFXPNRRnTxC5RpFgn6MAicsOn6mhdtwPM4d1BzsF5xCKyAzr+ZvLm3w/5Er+1WxDHiD
ELM72aatGfe+AVkOgapMltlFcNC4f87VKcA0RBRvwuA7Vk8Uj31sO2SHCwquCv0dNuV849IfB17o
Gw0jdzogE+oPzSWnp+iFL9+5Ht3QU1ZVFWoE2PDlC/DrHxcw2ka2qwKmEwCYvQji8v1pJ5MInNU+
fyuYuK9yIhAGKDgXzwueZlgAAxdJr94c++R0pw0UBljCsN3+99lVFAiFT/lk/DYBVu4VD/dVNCcY
lPpYrkZIOxWpBZyqSZku4hd1ylu1QbrEPbj9ASexyObfCxM5YCG+UsAvNjHVr8wzU6jpfZLwTA8S
18Iv0sDz9JFzSLmcSxnp10OWCfxxdf7Vp1y4iioPFM9mKac+7q2Nv5wYxOVvNtnIQMfs3BNTa81b
w5S7JS188LhVO/qQ2aInO2NxGIRi0L+By1EKnspJlquoruQVtE+nvI1gWAIoQzv37SnG+Q/bvOq5
JXKEcH3AhJFjXaKctpk8iepVjeAEMrweYThNdgbzdTf7w5bJYEhBmujqE1wZgvq37lUSKQSybqfU
vVcVTHUidqlEfMPFaEM+ePnps61kYAhDK8ftpsKe/0LwGtGvoTU63ws9G9q5d32KxSIYwE5C7Ig9
5/BNrON7wfYpiyYE6s6AF3wOwwn4qd3eVbj3CbRfl1CWuXQmaw5QveijRxURq+Cml2pfBQ1fZaNf
tjRVVgq15ZR7UWYo049kmIfwLfcm1BpOQtadXJZDhRnPsmTR05HQLqQu+Cgn4Tf+ZbzFUMMNZqwp
STgyVtBwpMXQ5G0P7YqGsrGkwNTx4HLDU4lA1nXl4HnpJpg7+fu58S1eqcTEX+Jtu96fcltAioxW
tbEgeeUBtRIwro4lUmXQlQd3uvjtLChmLfIU1KefWaKEB8k7Ujk5HHtRugMQeybvxBYbBr3zsGR7
ysrZnBX8QlLemvV3O7a9LhdaZ5DQTCUTLIlon4e+F3y7JSKDHL4csaaFdnXi/shdaCWBaqBaTBdu
g2DAMip+6EgLOfyA/tw1CaaoDyzuT1JGesNkuUXNmGEHTxCFIgqsDB3mgqMXfmfYz/vxMBwZCcZj
Ltw2vRu2URNtarULH3GqodvQ6G0F/btI6DFe4flMD4alcZ+/kKQ7iEN+3asGsBPUf4ukTzbWm8gm
7PyR7mCPHQQOeL7Xk+gn1OZoOAqU+eYpdK95eC6pKJIQHOgovYsuSTUeLBdDvcdncELQtNa5M/3x
jqgO+p8i5pNnYnHSttdTmWcrhxdQThci3nOsrv8N2BD32CglL9OCDRQXJ+njYV+8ngITfuKE9//C
XGG0kGNSjS1e8YwobZPg7XcMUo4jmnSL7oFDW8fPw2fUVv6w0HuNoaxSzky0DB5G/JZgPmA3Py+j
cNh6+rTNKBWwuz9pt/ey/BjIHEIcjE+ItRX3ZqHubX3GdUaqIgheyYXQmeUvzSdYzkv48TUmaUhv
J9AqON8G6e2Gtp8v1LvGQAsHW/YiOoMQ9MsKfulGoKCp4FHjHtTq6m90XtDznZUpyD5X4t9lE1H9
29M4d6HO8d+x6FHZIcjSJP2wWGa+1Gs/8Al/vuN22Cb/zek3k0T6lx9nhvSP01FG3vyxqm6v9LmB
sZm/s91FNstPkohAFskVV50wcUkGwc54mUo6UbvuuhPZdtexBD/01DSSne8gS3P/VnxQ9GHDevsQ
Zv/g+7FM2IkCTRIdUyWw29G1pMAHVyGfwu+OEyQD5jvWoIKCTUXxIGswShuxyfk8cZafKF1drhUv
pukfzuMABxX9zgDIjzk5N71jv3kooRP/fBpeIg16NLhYy8AgZAWw/MSN7ThlS+0pfDn6M1diNULI
Uc7J4dRSqPslJsZ4QUbdWeC6L0irntVrzlnbnsJuq0C03f4eff7eiobKqYWGK0NNywcuBzrnSRUl
/6xRRCqHyHxXPKdUqQiBbguJoq8rEdtDF6I+YFoPNq+0u9YeLxCDv9lUAFt8OC47BSyAtl7CRIlp
9pxL/5l8hvqqcUET/MDwJ+2g3tpZogGGmKtbROBvuV3vz3JdlsiJDJDqw5wJTkQZnTqM797bSjoi
B8oYPyIIZZJZpnX+0FxIa7nO8Qt7kRecZ1rzdYRzoeuie2UPgKsO53r2kUFzusWpcRooZ7ANxtoH
2OkVAlUh1+yL9MkaY7i7a45t9lxpPc8KqE4f0pLh7l/kfM/jPAEbeyqaluVYbJNLtB0+LSsstA1+
ML5aNcF6Yztsqs+EehzWygYYy2H5FlzbVw+J8i0/nuGf4RxhzbkLYi+MTn9Ri301zCgY+R2UUYZt
waAgnUWui0+kprJ4Pa/M9vndsxpUbKSEnVPEN0zftxyCiGKmu7qqDnhSP8jYQyawjDhzSn/iBA7R
YcEkfQos8pYSqBV6Ei1PiuAhdoUS9jjuyDqAySrH93v5hEjUx04QXu4u8fKhxEC7bvyqt7yy5s0N
Kq/5lh0wNMwaYickJXrlHYuzevMpGBjLNFuOGbcTDNXtphxyQJsjhodO0ABJ43HHKg2BcMi/gL/8
m+5eNVg6Krbl7mSUqTb15bwznu090bPRYvrKujmdy8sExXRq1xWOjgZzJFztGSMQMifqq2t1/GSz
h1y3zeols6ubsXv5xwC8MT7sVhJpfr5ha93IpUXbFs5u6YqMTrwefQAfdjVDE3JpeRjiL/55t3d3
YuzDRnXRiluMp2DQlBFQ2qVjZMxkE8HcK3PZwfbqP9OKZ09tBFYDXeh6TxJOWlC/p4rBbk1H1Cpv
/QneELBY+LkJS1XAjv0+lpIoN4fxzHD9Gl1mDVGKrC5oK7ckl9HOxW6p01ZC7OnfXyC9z/cSg9D5
QmlCzdOp/t4gWQLC9R+B5srfhhBBZRVq3JHEOfRJVLDQWvl0+hJWTOyovaQo3F6EoBaMe93oMHiu
+ZiC9yqknAAfjP7KXtaR3d5oXLc7cOUwf1zkMAZUfcPDF2otRxUjMNS4Ax0NmEw2/tsnC95pGMCD
PKcji9lAeC5Iv6uuhtdTS0yvsEZ8FjxsMjyTFvs/agorWqWwBEREuj6A9bGZJe8N3nbGJN2UbNTi
sVHLN18d6Z+AbySdJh3z4A2E8NENNa46eidzhrS9RtuH9iGS8rYsflZYbueBkmRpP8vNHTHiVob4
Hfak6fbQDDhR3HDN5KRYjGqxb7CN8tgVxGknRIXNdOORrZlSrgPSE8drMKeF4AMymFvqfZO5ZWwT
ssVTrJUZ/r/cGAQWynzeN8+JEFBCg75oGlrP01AdBB4LYzzHZ/fNiX9wKifXuTTEJ+29JXnVmws5
T8ubAjuCfNy/2xqUN0+Y4NFVicOe2rcbbVDnnnxm9C4TBdUrUZNqF83KUFeGmaU42sQOgD43B/Pg
ovhErhO3wpgOT07pvJgD2UH4rK1ubTRB/MHEV1epF/KOZpeaNEYFrRpzjIM115Wg0uVTUS4Fp9Mb
EIv0B1xlUPWHgUXw/oBr7Lte+uGKgeoZRYz1fLAZ1uxHj8Rx50jGPoZJ/S9JMm9QpFnBpTynkwBQ
bn1O9v2d6kJ6LWOxL67tAjf/xp1Cnoq3YafSw9VKQjizhob2CkvghZBU2A/vG82FO1z4BIKejI/H
TOYtsgsTlTCLf74V7TKUA/ANkYzvvjWI18aIVlFlP58/hr/HIS3sBz3S00IQguMVEHf25Ivkjuca
DeCQ1cfSvAwEPTJoyOHGy7U1akMrmvLmrVBSQ6Ltv/Kosd/I9Hx/U6Mdf7CrVYW847gavE60/pKI
CikFfF8KYdTk4qRk1oiH/9JcvAA6JldQLhqrolGBgh37o6s3ugqaJzvZpVSHZN29+IgbZTGMqZuD
xWHtKt7R5Cp/CZNdoRXh0padEbCoy8MH0yvbgONdbjrgcw/hx42ITWEI/U0JqsmLwvFf5hSdB3Uu
s9fFeMNldBC6by3kLRhtu0+6sSHw4Z03Wln2JR5TvNfoJkaW1iykJ/LQk9a8Z+ryTVACglIykXJn
HEO8MbyxABXCoAE9CiYWcdmJhol5MnODfbkfjlZwF2ZCp5GGotSmx/ZpdxCXN8FBRQZ4dljddWOd
2Jl3BZkS70zYxdt3Nh/MzHqz+AR+UiY7SiSH1ya85YUQQE7LYLo6sSPILRN7pBlITN4QYFCzoVAC
h9jFJw3s50A/eKiZu3S3vlMsvLYkTMXk06YrICsEbOcdIZ7DloRWhS2y/dcAat/aL1MsUhNjyH3a
cyy7BGE8ekf0Kteyn5pRVtAB5myayw/EdzAA4370lB9Rq4yeDLxNYnBKLbyh7Jko0foa5QktXw1n
sICYHz99hPBwL2EOFMXmB4Iz8yS8lVMYiJIv68lrYRm5czG1f0ZPZHT7zweJIT1wiFcf8TLSWe8F
/iFInXYQ8+dG3hgAskrMA+miQcEXp+S/f8qD2pikPhfk1RJ+unhIR2g00oykcnc410citKR9cwTu
dDe//hZlA2oB4xUyZc7okGAW0IMIxe4ovxyckEmrcb6l+4whBhMsxjN7KcbnbX+RxmibBcP3SlL5
zimikC1U8Z/R6gUVFVufKAF35h24xF+1bdjzG0ZTDfOBz6FrYg5F6kdqU0qNGRm0bZuBo5nlVWWz
ML6dU0X2VusyYmzOnJhuwN41yMmjkemzM9NgpAjrHuLZCISpVmtbGNO/v1l1p4j+JGWX08ryRSb9
tkHU57sRhpniCUtJ4VYhX5+ZG6YMATqpn/NXA2I/sltyn8JAwHN2f+nfHGmSdzMXYJaEZ5ZVUzUm
CVecrszHM3lQ+N8TPLaQkVkp8OIABnbFOKI56oASsEKJ7UsAjyfvx8jzE/0HdiMEkTXO1+F7+mx8
7Mmxi8PKSue5ycn0OVEFtIMgHEe8NJJHVE3fqkpKzNQwcRtoK+KOVOxKsIZJx1SFAuyiC+4+4aLN
qoX+oR5iUQYklzAixqNQx2wcJzWuxdUFdflZycma1FzQw1HlDHwWbxaMbsoqTUp5RhCqiogJ9J4a
c2SxKuuCXY5PvS1jjxScdr4LksrFXRpObw6JhKbAR6unO2PakCEIRCyCpiScWzVpSMRizNIFoPHL
TdOPlMSZjtCo96JvnNy+xu+rmNGT/YHZqRw2cnFZphEEzkHHbDusm7clltBcfFOKmxEQl35teTvL
ovxl5WDkyCBuZdf9qgkxBIsBXpoU7tlWqlRnUPtiqpzzJ/UnmKYd23+poeOceVJunGo3prOuXpGX
I4rzOx17Dwo6YsBbsIW2np29yDeS/klI510IMdedE+M/WubWzEpIwWwmmjEfEAzHtDLEF8wbY/QI
cfiniNcyqy6TW0QcKvNlhkKa/aZCRpjfyBm5LH/muQ5UJy+E/bFA45yZXG9huzQfCRNAjcgMkUVU
ECNYHB8NDXrQKtEC16CkidRlYKKu+o0lF53IwI9BjR21CW29rpIc8JTq/Oa9S40Yg8kL3qm9F1q9
0gCXGGKYQJMYDuCJA1NHD+84nbxxfiyAo8iACVtGJ0mSDXsGfHw5XL7o1DRWlGQsxNf1DNyZYC80
bvjGYkRJ7b0zF/9Gz83WCwcUrJFF3hpYWl5hWr4TiM0d8b4ONgASZULAZyfjvM1Ljm3/rhzyJyR0
Ph8X13e40dhTFu/6akQ/UomJ/WljZxJQsL3/e6aHzERsOJ4jakF9P7gf2sw/66kzLhjE5v5VKlDJ
y+yY7mCk6w/mC5X0A/U4AGumY6ya6X04QLMj+2WNQr40d4u6ga4aPZeQs8R9wbJwqOczBjoQvxcs
qhsN4+snStTRPrDfhmAdojolQW2EPvl2Y4b4eEblLyoEOq6CQaP3CX2hE4hJEonzOsDvq+a4ZHcG
Q7ffy02egZCu+ddbvmANDNyZTvSZFAzCZRyBsLP50ax4dG9MnxHoB2HwrF6HP6ZVRXz5C+kNinqR
60cTV/1oTcqdwGuSxjoCzrI0dQ6GVI39Xw5zMDK9u8YzjVsaNFMUKs9JUguyBworIq4ZhTEmDKyR
Sm2Sj3FZPiDfN9WRKbJJz54uvVDPhzqFy7s2p3Wke1sRtccduAcJUiUDR6gZlKpfUvUiFiW3PZaS
VePHi8GlcnxQP78vmEKIp19dlaY1eUibmT7eFyt2kk9170ToO7zwIXw5jU83+TTR74DTBRscAcwz
qVNWSPjgi0suxQIA3ffqc93KDO77FudmP9EgkVpBB8MdBLpO+pHECtcmM3BC6RMfju0hx4ULFBy2
gi8mmEyheAPLeXrowZdnL7obgwc2KOwLB4Srq1O8EwriIV1GfeqHQrQB8nyt+8gArvasTm7SmQ2S
LSwJ009kKMC2TcLxxxxyRwFHqD+XZUjlZGcx7boyKXjI7Hvgm6t7JF62ZdsSRAk7FrUAU6wQOSSG
zlXjbxhNURIlLRe3Vdee2cvJo/0q0T2ytyUFZZAs+baMmP3ERjOVyiwTo6F6XIqNE80nkOPqhJXJ
/Kn6kHPqkn9rWEV4kz90Mk+FaQYGmV87w5tMOoXqzaF1YQ9QM/dXQ4KBNIYrZ5kDQQFv1MNn2ME/
lBwEWzW7TL9FjV6J3qiqgDRv1KqASyKJ2PBWH26iHcq9+Xucua405kcyxKMFUXxaZbevo+W2FbYA
A97ySOQytem6G1rXDI+8B5SBlHpwheDdyyeG1DDi0VLnTZZeH2RfiyK9vb+h7NRx8isoKPh8v+1z
nY4sBsBgPpU1vUAn3JQcYuQrH2t1C6xjzQztzfK6HzhUEhHsEpfplLLLToZBTkRkPdJY9/6CrZxg
Ky6qeLq/hJICSN7pm6s9Xyqtxa2mrj4oKkLoph2tu/SZDtzo04m5HEk/0My66l1AA4wl34mKI7Zl
kPK1eMQBj56yHAhb19YO5E4K0/yRzsZFuwC1YBIDth6P8vyrBBe+0ugxwX+TEZ1YGxsOxkq0/R+q
zusC2zGJl2TalZQuHno5rvuAqmV2A/GCBO/VFpoFLEmO2Lr9tYelz8eombhEKCCVmiDEoyBfKThe
MJYEtBc8Yda/SY1JpCpxU90OfvOeBh7L5q7BccWoK8DUDf29gNnfCQ3C1JQIn8FLIZoCRh2STLVf
pWL+Xe+bKwFr+bBubo/5ftRDcOSPTuBANIei5VVMXPPH+lAlBrvbmmOloldwQzYKqAWwksZJuWAc
5nfgSkxCmzu5AYriQpomlGZN1P0+KNxf4gPfZf5S/1lUNiakPYcBsX+CovF3ASCjNY5mkdNXY6Ub
cUIKLSPFCVAZa7DQNBoZOKS39bf4HDXkl3Taj9E+QTtnu4tozlYTw/tnRrg1rQZSpi54YbkMR5rD
sBdEwNdtleHD45HgqbwW/uEA5PXwjEIPL53AT5ralMcsgc8kc6BkVbhEEwnIcrAwWpaMWmzHRBDq
t08ItajKF18JEMNN2nPPqNt9Gadn+NyUXhmaUbsOv7JIpWEiK2miTdkabBdKci86C62PAmnoXXd3
adsZHW1eB/n7goIkLKbxTCyUcO7fJifqun3OdPtl28PYMB+82Zx1wbiTbqD/4tax1hQOcydRUdec
4OMJ6bz/zzEDKL7r4urPgDeQXKvFWbS7cAD3z0bSiQqdY5JxCtYX1Yh6nHTCougaFZb9nwe3EnI5
/EUuatG+Usrzka/9OfEWeaJ9ngW+Y7rVUKpwvJP0YFbHfXvzWTGI8k8OK1qgodpK05UR4SP9xro/
/XBnEuuFhpqfUabE3pi4BVLSYzpVoXKfdm2/cF/XVG7R7mdBGgA3wBInDbDD0y+/s67CDNr2N0LR
EHjgtpRKRhycHHPO/bQ0Y9iGfYGNlG6gT4uVEfnWc/XPt5DWnrd0rIJ2FRD69RysEeD5++OKq7Lf
XvHIKkcQWOTilsiFDDgm7M22GYxYp+XRneOCRGNxjJLkJSZMH6gtdYwxgWoflofWW4v5Oeebs7s9
KBgazeoj+KIQMGNC+tPAYSfwIcDQp0GMKPZZvcPT6PwtA0UhYpQdwAEGVDi7Lt383rWw3pMc/1nR
J1lppl0gsm1IjC4ZxhdLqt+Y+02bDIo2MPCM1KY+OZS9+1Xy1LlsntYQz3rKtdrdjYa3OBj4UntG
e9Nfe9CC9xFpp277nWaM+KpCrNpRYfqcOOe5rIa8DFy89HxNg71D57FhfVLJYHqzLoCrvZ11EHgl
nou1C4I5+Loo1O49J9HtzGrQk+VcdZAntRkCzAgibdWdcakt8TEUAePzp4OZtnI5wNU3cC+1jVfa
EZdx7CXS3j8HTQhams5chJTdfp5jtw+qSpJ6l3xWH15lf6/nfCHKR7+BaScwS4/DYrfXowGb+lxY
q1DTWXyNAgJw6DfrXaySpjM0oaU6y74s7lBwouqc1pHnkhQWx0dgfihlTxZsOEUaj9fx0ddFr3n3
Nb6/SCVkMcef39kRrIDtwTSULZTF/DNUvjvGNFffsPhjNfCpXahAKl/9t4SpU09jSiz2tILBtimG
00HvSB7L8r3UzrES9CW2aYFpGupPCuT73agUemTK9cWsLVil4p2xDNA8DNgfU8oaTORBkkqCRLtZ
PuO3ZQwDgHYs0nVnhf27BtDBB8XAxtdLiYuw3pgSrgX5zvzABb/7gpY6LizOgFNMjsCPXNlFPyiV
nhmY8KwxnCOQEhLk6x6jqdJnuYed6G2Xfk0sqN7DMpt6Hm6R3cRM4vZtrPH/3rhZ1sLxZ38UYWKc
5UFwbLPhnu4bHQcID3wUUdDthwrPy4DleBpWBY8N5yPK+D/Bm6sdTb6VtCO90tqtesFNDjHtWzVk
EmyQ77DmMJ+ccJYGQEvx+GV2+UVrfsm2jMyXOAMvMlcwgPHUsCc1+4qjpzS5mUQ9DZfhGwlcsLut
XTmmLFhq8wbpWl3Ias0qcu1LEBh5mpMqw6W1R55RNBoZu9VS6yGtIqlegjBfzXnMChEO15TITkQl
lZc6OtvMAFejBsJ0XUD/B50JAx4AE9HW7lLfitapci6NtwUoPDDkI09GEkISBshtVRCpdRReJsbF
JIB2cCrfuT3TMdC4VEG+zjkwfac2EnXRpgVXIR409RPuUk8dFZEvVBBJzbLvaIX43Ew+MdvbwLwB
KrpF9f5oP8INkvYV95OMHTwI2t8V6X2rPw5QXyvsjh1duZRy59GMFS+3w1bHBkBs5IK4TfzM/wua
zkY5USU+AVGkb8uMjqdtq+RY32W2ZVs+R0T3z64jwVMJRNVaBHHKlx1CcbiIrOFVZJo2IfLg5nxr
BtOZG8+/k+dDFhf6RglFZtAXjNv3tzz6xKbtpl+dlXT9sCLxcIUK+LDeKmWP9bVMiyBOZdPfk8JS
nndGLlm95BaRwhQzUbikHTv/TMAviU/IWnGJYOMl9Sk0AuVEIh9cPxv2YFwlUl9EmUez6wfUeNta
AS+0eMsZfnJJ8OUpR73ikoXVPYAY6Z+H/fUD9Px59SipVRoJEemKMcyQvWkWLywYN9eicvOGaUYB
gioCPtkXtuQsY/GIt08e5DvPcELz8bek6Ir1U/ZAFTHHzP9tvNakdkbat7AGIoUgYba1L8S7xg9E
0kAin+/4kcNJ3JXro8ubQpO6SqPhDruntBg7TN9jJAxjkhfZ0CmW9uZkk47LlKzJTI/iCwQ6mJle
abKdtoqUyWom4LhJ7LZnvc+fBbwsznUWm7cPfpuAnXWUJMFkTVI31ie4uamAosGa0t3Fj5WwPKSk
aO4okjT13O7Fs1uwSlx5t+RyGI8Eu96F8oEdCPSErP26ZH9r2FlJB8WFAaTMySN3tVi0TMfbnPIH
cJKgIHOHyy0APHHZ+acYGW7k55VA9Sryd5A6NWOzsjNbHuuHnn8O7kwVRSg+xxd9Omfzbm1pJ/DU
8uXI9aNLo+jKbHWynd0jcUHD+lhNg2m4/3khgKbJjTt+RvShbk67wt7BI+RW9W0IrFVMVts/Gg4T
RxgsY9PpJEApw5a6FTNgWjyvgLw1cPIWkrwe2qOp7Z7VHFP3G/cMscgyt7KLxbHNO3YeXWwOj15t
y7dB7s2NADtefiu5m5xlvYciv9imdXMMDBiMxkyrwPws72nnTrEytwLv+GDgNttP6C35R8NA+eIb
75P62CNZbB9zfkGFSrKUH+xIsg+kqu3gyfXqJTZCDgWELtsf2O3YwrQlig9orV74TIJiC1ZPtC4H
lofwEKp2o5xERHuoWeOKfaM05OcRrdx7Cf5eVUPE/KDI/0XLbubDEXy4TrfP7Avik/1y4J14qX+u
fEvLC33MWTlKgko4us6yf/jLnIxn0OVtK7q4YlEltG8VnzOO/fBlsyXN3TURrk2YbXTbthi1KTiM
2HZjIH+hLO1JmxDzrnm1en6Vd7zaNLI6J5sCOVjbcT96FVeYFTkRk1tGN0sj/QP5UIXcegP9ZmCO
evh8lsh3EWJSlTdLxcZbj7AZxKBuuT1W9TAj4NcDDWIZxoElnUJ5KZKJTDjN4XcaDOsoy9mgr8Fd
PoaxaTDdXytNDj/EiWpDgZWpSc2VbjtT1G1yaiOdxbosNQLGTDpqHC4pS3/khameB3KQ57NbM7PV
0ld6V3xOpnbWbxDBd4+DKyaiNukT/KpXffFSJPqg371UNCI+2kkE1qzrIPtcMyqPgAWTJnmp1wJJ
fnySF4xfCfcHVAL0iIEo81dU531twjW+2QgPmYCaeOwFGfbwEmUbyixJh92pmfdxB6MV+f6yKQQK
qxrKMEfcQgsajtP/bnf+t4J0+EpOJE0dOox9qmK6qIQnMqgfgGWu199nDpqyQTDEsSxCuHUoWoQW
rBcTkIi/N/CH6OsRWChDkPm7665iNoHOaB4r+3PFRXHCuYCOD61Amc9RPar5TLh73xhiQW3woFSB
ZZ/MTG/0DKZ/J/vjJ5TyVEvclUh119h2A8Wro6Mb8mVpz5L+WjUDXgllNaGnuozEGA2Srb1nwyD0
+vxE337yXmBdD9A1kkxJoayN8LoKdLZROr4gsppnTRU3FXDaY0suoIJbWY+NFCxo3rH8G9ZpqF5S
5+dRjfEgQKLouozy4yQNlUGnkVHgPg3Ztqvd2EXIk5A/S26K1uWKWijmfTdj2rIJjE+S1s2QP4WB
xMJnTV6vPYIpJvLCw7LEOApHbRT2Qgx2nMuU9b65Ipl7J4noZ9gl5DEhjKywctjdLAasgQOiYfCl
czI31ynf+TNpOwzzDD2mqsDr5r/7G+BOXtdN9FJx4ZTggZUg8DiFd0qpGdBy5RaTqheuBgEKgg1Z
H1gsju49pfYt3owBtXPaLdkPyOVwq4G8eYq7QffIlHImEytWFSZriLoe0j+lPEf9K4+iHHzqzkGy
nHWu/I7hVUi5kIbfKsMpIBWjRa9WgadmypHxm6lhUR8vVYWf85zYSt/77z0YXhhBOpI8sypcNTON
ifTE37hhHtUw1CTQuOf9tTDrqogpmTGwaN/Uf6dxtx7JM3BM7g3tGIAtV2QXSBErCWpOavYWadTg
gPwg4zQxwq6RoRx8GnFHWu6Xhb+/g+inuqS3ZLGqNUjO5yTbn+VTvP41qEhWieN9Wvo6VJ0KK2cg
Fs9u2+eNiau8ZOk9ULjeZpQ//J2Qs4oBgkf/563nu2yzGf5nMHNk/NL4dE03OuHXP8zyRxSvCe0J
Wd19qAgXnlfJ3LJS/BZDDvShA5Fsjyb07iIzwIt2fFvUIPJeyQIEo+NSrUAOqmAYcOV+xqVy96Wg
wNTHWQc6YVmrcS0VqlJhD6PUViqVuNnSPSn33QYiFo5CU72+QTkFMZfVInceyj0qhtDwP0ORBENU
auBeFqxQshL20sJWTwHpMq6ojTu5F/+e7q4S5fkonvR/JjzGyEg0xgPFVBgRW7jWQ9zR22wbNcH8
mbFjYQuEtP7rhiV3FNeZp+7tcwiOf8Zgjfj5roHDlzZBsKf7bW8PbbTibgzVNMLxAP8IfzfVjCEz
HGjOpC/P34DC8M1U0OmaVGGSXxwXFo9jf5d/wIK/nBdCwcVpnY++PZzlMeSfUawIsH9nPswZYgmA
kEkhMSVyGjjZW036CQrTkRj20xeNNkTvh5NhYceha5lMpTGlsX6TdOXNc08yEvkD/maSE50rmOpY
FTDor2wK4G0y+9oYMEjao3JywcjXeWoVg8p/mEZSAhD6gUUc+isGBz/CTVjYHDNeEjMo6Hp+WycQ
yie8aEcC85UB5Bj28B0t5zN4l5RKgrwNdi9I7jJXBPTANdez3k4zLsvnW1dCK3KBZhlX/4kY9ocL
6wETLJyrF2lwb8z97XoDlWsTTxuUvkM9RrayocVBA5Glse5yyAAXCIv8f4SHj9svclyAI87Xy7Tr
0Z8E2t59l0hBaCQ8dLAPoTfMjLgrHQVxC4mATAIxwEO1FGy85Y30Mgv6zfCI0NJoXyPgrsvv1HWM
SMBBz3gtK+VFLEaYVeuYlwL/0VOROBDqEXbTvG8IZ+yZfle0WP5vg/i7qdAnFxTs1ucgSSx8hH8r
sD8Y78qnhVEy8VZC33WLm6EkK0Fzx9ns5RTChcaL8jW0perAYLzJnozgGaOvERJuuLV8ewV49E7z
l9/Uj0maWEw0blA/7KoW+gd/w2Kk20QOSc+4weKjJ4rfu5gY7OmHwmGSLBrA/3yKrtIeVHLM5Lee
H2nUds8cxcSLXknDWAJrW+pD+mrGPa6fCSG8vnB1SyqU1FxIXW5Q0ZJlDC3ynhdaPU8HceE0l5Mp
D9IFcGuxv/fD0FBbMUkbDnVx0utUIcXkdmw7WxML3LpVatc+OwZiXsKKf9RqFF5J/GTYX9V2Opwv
2xEUfIjaYXEz2Jv+73bjK9CAh4ZDZxEf4YhoVOwxtI+P+6M5v59Sftaq/Jp1RY6iehF7BL9n2Ehu
TVoStmcXA0CZwiGJUzTCU0QmU5PBtp90hyOieiChvVNXiaKSyagjqdBeXs6a479e4kE0Wy3sxgx7
4y/tF78YJofaF6hLxY45nox1bsJvsOJuWgehHZEhUCJZepoGQamI9FG492MJbDBNWhXYJo3cU9tr
D1N3unSaHgxa9h8wCscF97P0yblctHPXS1LBlGmQjkmy3CQyU1o6Ad/bxN/LbDmQoINZ7d79yntx
ycnZZwXv0RnYuV+1s5hcaTlOgNo5vccg/8SxLX+rIKlXQ+aK43ArxB1NhzExkT3sycroVdNHKjz5
dZ48BX1iNnRPuJO5Gan/F6paJabYJainwYOfFXPmMC6I9tz737+/tlxmZ71KcrbjM1NLFnsnHC2L
uChk81Xz8Qe4YyoEcTu87E7tTbrm94vpdiXVrsGFgANu2aQdik3Oq7xYa2ISTMeKMZtw3wlLjZJz
b2Zfk+3jOnWv9XdqSsYCXJ0byoJwjBZVKWZihR6V+3ktQLqrwEJwEXZGMRLW2dmNUC0T6YWqcNHv
o6gc5RUijKTfyA0JOWOvsp7KQon9m9QAT0ldmOLdIxc0L5Th54SrVmMLgkfOEO1PymUBc8OZ8NbP
wUPhDLl79OEHe/al/5GTyPMPT9o2pbA5Al1jSkCZhkK99pJsGSLTQ4PDEB24FzK1pozywxoEptk6
TQBaZ0BKFq2MXSXGQrp8pkI6DX3YrLdzap/0Pzkp4loJtweQA2aoMLTfL1oWjijYOTFLNOmnz1vK
PrEeb06nno/zF4XdmfoVx52ANTHySxNyzH89fZ7AZYQpEiin5IXscrz6oRYIp2LxjZsJ56ovoQjF
Wd4M7TqVl5nHjIkCi89zIelhNnR/5pboU3/vivBHfU1Y9ISrRInhw758BJ0sMq4oW4ry0Va1kSqB
Nt+P9vqXGOYnD8Z8tUSvk0ueqNHPJDjUogW/igiLM0Rg8+6MqQIEDwEqc6i/GIzpfyIDwtw9aAYE
AyHRxoKI888gnapzq2C8iFsW8sITOToyf/3L+LX/xanvzeZOlQHCVpIM0dJ++ZblRbdHl4Yvis9u
fxnuru+F4l6FOzi2CXYtEHi3UL2Qxhw0Mn41uthoYZZCtPnRIAHUW38UsKMBGP1pQpbgE0opGmTD
YQPsjrhsFVsDZLAYX5GC00gDe7ILpk4EK3dsyjKwWrQUDObDtBPxMjTfsJIHkghPy9ZBWH5gK7AJ
aO4S2ncteL3iUjm9TwsBYU+oSc7XDfrajl3kWVKBwYbC4FPd4L63J0UyqtF2p/Z7GfRPgLBgfrNG
JfLrub7XYQlT1e49KuKPFxViYP9d4eap2BxONLj6CZAk5NbOsCuKw6fJogLuoZ+pb4z9A/alIRqW
w8dI1qATb9l1Kwp+sjYgVQuCIMRMawbJka7jg+1fMiW/IGzFs5wJl/JBB4tjl3kEnEuYakste5Fq
MAqbMgxcjHAYNkGZm2RYI9ITAIARIQKO/VjDY0+PrlPPQDX528ZCqBjn/I4CSOj6qPbZjkpqof+X
gnHmyR9XLkIsXuNDAcN6HuaAK68LCVlzCvYCVmQuq2oYaP2XUqipxcs9R+XYrgMF9185xZEBFu1m
6WgHUWRRZepQetPcbDhdlQyqVkQKNmsxkVVWmee1ACJRHgmSAtmcrLB36yHwicIIqooHkN7MaqV2
7bo5GzAJq9RY7/Xre2fU6jGC3R/4PrBbb2RGQ5HWNAKIEwOJAX67JLElzpUq/8yjQCYQEiGbw+Mb
Z7lvFtshWhdES267wyxm5FCaOT5IhzjXeFS+lecKBjLnLUKMkF4NUME6pV4Ez4nSc2WQw2jY2UkW
KYsm25qV+OkjQGymalmxBwm4HlwFwkgi55C5F/ku9EYyNRSdFmev3wtc9uLTDQAylEXDABcfk0A4
mhq0Ll+ABBCxIAGgw5vjwZ5KCgQ7xT4gJTvCn+4KclPfk2sQmVmdM7PkbskcupyRssrdACufsVJo
NTlEB0wL6WW2gJM3UcAzUpVeShd6TLyuE35BzaF0zZM1A64Q0k9zZNLqiXMr5eqxqFiZzgh3hJtz
9TIIfBeTTLFGT6EmxeV5aLEC0fXBKxvhzfzvM+pknVVdEfok3WPfljzaxJbstG/vNZPHVtYc+IMZ
ixvUSIu5LPyFhvX2SK6yl+mZKcmHpz/JhQdwwUoVa4cV0YA+GlNKB9zSAyNs6xHgxNH65ObXZIRC
SuYrc2qAHF5F+2vGIU96KF64ItK4Km6Bc7G4+5/KiAuisMn0pp/TroqDH2LQzH3jrOBS7R4Y1fHF
0u7IYU0zga2uujyDUBwZBjvgRTUhsY694/FRSDOxgekBss+z+7daEb5BFFNVS4zS6G20v0M2STT1
DAwTYQOcy3Sd34hE+y7p9bh6fxIn5f/SnqZcUxmhTyKx2HzN5Dp8aMFsj58vTbRzCllBkKhU6BOE
QN1uDKChM9M5HwCRG9sU9ZycS75cxwfDw83nW1wAvkovEQyTjv2i0bPC3y+fRMVfpRJEobBXnbBs
C5NMRfSxME3a3J1Ytbfj378CdwaexnqbvMqODSQl3/ZUx9k2igPtJtpBV0tOlLeK4ay+j9vELyQA
Gy9VrzpISEv5m+Kfrhdaz6N8cy2PeQmXVCMHL5tAfnX4p+BFDz9r2OqyVrwP7w4eOVPFquTfAXP0
pKvSnkUp0bo4r3BB7rMSB9ksxBL6XPbvDVjLX+3FQW1TK+lz66gDpsnm+PbsxRwOGjwkDCU4ORWd
06NtlcRmtMFXz2hYK7jFub2Oj5fRy3CRiJBcMUBcEFnJjlnRpLNI7QUHXGaF/0Zi1BltgERr5l+8
0LnoK1LVNIMhQ6n1r7T19DOm4DUQWKYzg/GUJ44JusC2kwd4bxa5bXlxB3BSq3s7cfumKIF+gjtw
yAZlxWVCY/s7jG9jLeGJU8zseSN4ovWUwIwKexX5o1BFyyRl1Z9pXXRAZQ27kp+h7U8PItuDM2ef
33NVYja2YYiD9HYfRwsSk3hkfDbhhdWWQhYRj7wXCa4pkXGcThygfl0f0hnrM2vgvF+k/SYSD2VP
58FWpEWDY/rjiB92LFiAEljKzt1b74HFu/h40MF1kKTfag7gxtrL/K35L9tJ/xcY+aXK5d3JqXRe
tcwrxfWQuRDlAy+1MAZbEeYqfV+UH0xQv+vIz7Qr7f/BOvLJB2eIDqBu+VMBfIDVFAjkq7jYxDzk
0kaw8+SPb2F1RJYhZ3+RW0Tc6oq0e+JKpDAT2GHxdqy7OUn2TpRGKB0a32cW90pk/Nq+zK5AWhNC
k8H1q6tm+gC/l8r9I9JoA4+6ija6ghdW0JzSHIXLRBxJS+roqgqFBHErCy4yc1FWJ6qDp2AiQ4HK
Fr4c6s5Q1C44/52xhy6hdZLcKHonDvDNHq6bRceaFJ6iLriI074gcMJ8qciuhYxFir/R3YPC/RGs
nEPDljPH20vWpFt6uL2NHITjK0gpU6S8ZNmXh8udAXN+x8gprxA+fjX65/Pk4nTMHxa4mbWRmxJc
BBKDB/7K4/kETF4Tmv8G9nCJv8BYv6VpEIwmBxzgF1pAKddpIric9BMPsEgKI2dKF7R/hrM7uqGG
+iFbN+muctGXb59E9EVBwGX64ff8clO3yN7xpdQ3JZci9mZf6rjziAwh7jIg5q1HFfaO0yUoHuE6
ukiuN4OWp6xLcQqRR/P2640ZETzafoC8MSBdzf3Z/lQ9J1TDkj/pKrPus0QN9KxvUTzCC0Zwi9kg
q8RN5r7b52CD/5feh8rW1SKLQqSW8zdb2n0Dhbm15ASqHaoRA6WXi4Eey7g9ibGQD0uui0SSXXHc
QRTpvxgW0/btlLJdz09WF/XsAkAlj5oUnnpZ2Or8wvGBKuv/oZ8NzU4s3nOkBDXLsAWwfBbSKIzU
BX3PN/wgY1LqIOwY3NbLoy+GNaqImOvd5NNxoHmCwzSyDCCjENK+GT2fCbNKwGm1TylDNwMK92CA
cL5TUCss+Xbva+eXdpSFKjWyYQTfJtL8uap638yuhwDnmbBdr/nYJdbpG9gHBE0LvW5mGreytynk
92jh/CRS/x2Rg2MdxFpAnVqQqarUErZRgzAlE69A9N/Kyfy2kXLqMHikHtChLvJWHA6CvxpHVvMw
U6qASZShbfdIygYDuvS9ydHyVDVQsg5tlXex9tJGLfg3BsHrlweJSWBL8BnbwIH5d2J79hcuK97V
tZP1+gIL3Il833OvyW8WI3QbppMuNjeyfzAmxc2ohJUPst/Dq1dQLh7Q25BTd7kBKG/U6jYzCR57
i1WNOGVgLvGlKuWVI454C+yxc2G9bgq8GreZJNi/Ps8JkGZTOf8kyU7OHkSfJMCdS/cznX3EDWiE
oDicG9DimiXOthLRQbM+rP48tHmd0vvSK0YZAO/UImQzp6Q33b55qa15Y7xXdcin+vMI53qAYoyh
ezC7Ac10zqVv/dtKZU0IqU/INyw8avaiTNHTGuA6z5tW9sOn1X8pWFa8eMfd+l2cY9QNFqG7q1X4
elUTBSYa+wI/r4mgk8P/mv2gHttBI8XMv2uHos31jlpg3fd+OI1O4WvXmnpq3pKNV7swpvS6IVWb
mLW7AZZ5ImBVOt0Lj8wLKRYsKw4fFkTE2dAZscblUhEq+wg0y2/O3BEQJghmT01iQ7MX0lSlesa3
N7B7DcWoTeaDToHIJFlSRc3CL8o9u408Osahar6Tu0CLvXIiXLHhJ4pxrEpgNtYcBKW/UpACCTrb
cLNS1zkPDHQGSlquf11Q3P2M5t1ZptX6QwYytnuBJ2vE2gJiT/MM2YaL1Md0+WQ/RwRG1x+DtTE9
gVNVyBSurhAyYPXY3cMjsUEWdQkTf/ozXzUKWDQGmWCZuGKaDQ/2H8ESSSFePL0huSIuUt3ZHf8f
RcODRboV8D0XjxK1tJ3gPN1Nspi7vP4Hl0QVUW+u7k+AuXgRP8TYlvErG1WxoL/Y3Oj2fiwhPscx
WXsE6ALdvqRkpdUbqYWmK6qWh3QJmATPohmPJIUbM9rxa7/t5CUGmfHFkK6dVRZd//Jn0srqrSeY
oPcpNFIRN3JI0SNp66bectCrVQXSXqfrNMl2MEjOZP+xrVQ3Z4YHqmSBoR7t2icJBPSWZ5y6GGCD
CXy03ufItpLG6DNEq9ltTaVd7USYoTGoQJrNIG/8e/Q6htlN7odR3OSL1xeXY6+cqrXkj6nPCpWH
R/hgnZrD7w+MT4JJHcL6Q+FsqH7vYbZDlk1MxGyzIrWrjUzluMTlIr8PKGpoD24JfpKZ251lWLNt
rqZMzmCnOMGNbp1W1Y5veWjgSaEy0nM+q+jLDXQumxioQ6fcD2HANUrXY4O80ZrpHfdz/8BXoyzi
EPThmI3tFr8mM0Z89dD5X3Ccq5T7WikAKvHma2F7ci8h35jCb+mFf/OAAfzLB9hXa9WKrr6Ppxvb
OaN0JOX4beqh/OIYJg4G9MBhueKJUmlX2xQmEthXNr8e8MNWYU0StIxLDb1NQk0fnF8s+HS4cH4k
qEHx2KznRsT8EbS8VZoBhdQ+uBjRHytWwEkfi4Mzgsr58QgF02IYJJT+DZkHbE7EnQ8bZCj20Jyv
/ORly5GI+IACPhiqyPjLSRER31ruU1yGfGKy1lfUN1Jnt0U4BJFgybHgE+chQZY9X2AVGS8cgzdP
t5RWWKyQY/QPpnE/jHoC7LWenQx3693dfxufOxiKGeLFaU0nWeUzwW9KIB/Nud1NFxoIXcvqK/vq
I5eZlWumMPBnZd4lt0b8/xcnLfjNmwlfsiejVvo1p7fpJkkfGFA/S7BTpJpe/FfPwQ8BHZjsSgTh
f3ByF4NDfJtViZ56ln7gdV+U5WsQTgUK5TdaIy55+O5C6EqxGe7Uhl/kZlnEQ9iO0iYk2EDvQ2rq
LBJmwayj+WM94QstSHbx77kc7nzLQfJV57xVuwfbwJx0JXLgxVuHARXM/kVutuTNYsW9QNPqRE2h
s2Bw+fF9a7qXGdrEXt8n1ddTMQYFX4soabay7NXC6UUqlZ3HY+qV3OseO+QpZRB6bVab/jF3XyU8
BMbFR6J+wabk8B09QXSM/8OzSiHjurC45CzM7mR/dRX7LeDhrIttzRy0Rit9cuZtmSU/XxXHuWl0
HWOH4zBUr705+znLugJcelHL6/vE5CL+Rqpjz5HdksJyd32PEKOfxCAY4TdVrzeFOTGhXDFPW9qS
ieHJVVBLHSwyFxFi15dVhit3NgrFubUjdGxaib9mS3X3e4lSSrUtA+URSKM1Z83sAo4W6hR0VqR0
h7ohAQCl4pwO8UjqYI77XcDSnhTiCRJQ7Ls9gIJ0IYNuTWjQ5yENoN2xZSCkvvkRIAoxrPf9Eovq
xGvWq/94FEyGvGXTGqfEts2lBzJcEmJ51RNs8kdBoWH7pP244iW2Okvlbuqm7mD07l1Vu5KuOWsG
Djvg6V2846a6A5cb75OPo+jnd6q23+ku5oeaEe7fZMFl197+Vpmsq1Uy33uYjZxatbdFj4N5cOJA
wR16WBjiXvLhREUsPGr6cg1XglcrvkOkpNKNNQzCF5PtWCh8myYFHZTlPm83p9Tcnn4v1FDn/VLk
W331Zjeo2I0xnAl3FdbMhVlvIyiNd2qKRl/m2w4e/W/dH+uXmrDFWlFaXbFz031dzYF8KhxBjg54
2I2ZbVsvG4e7YW6r0vW3pAcvBFq0h8UB93VPiWQcNRI4ygwJmfIH87yDKBx+zSJABDtDrA7trdit
frQS6JldXnAzyrGku/bWHz92QbRIo8fp1NOyqLOgmJb1DGDvOFN1Ldbgz2pBz4LqVzKpDQmuH6S0
idE/n1k9ntRoJLEuNfxBjaQq+q1AQTGqwoNZzi4JmNkc1lS1htKCXdOYSKtuYH0rbhQnQTuKoPsb
laARnWxY84MAovvFvVkD4NppAEOHQyVylSlRoCxgmBWT7GvSWEuzr1DP5vG+gwACsseBNDGwVatY
ABXtaj6vdbAmlNdk4lbWqapQPqYuTc52wkV1H8SS9QgTOqL3idCgNXD4USHyP8FWAphEBBgVjM6i
DdeExxeeiwm2+OSvhXHL7w+eA15aPWXLvrlZ8Yw0jONqTrmRLGblFPNUQh8OzEZbm07gcGsx/apl
AF/zpzosQwnNv9xNW5UiaonjBH904FQ4/XdJ9J8kUjAts360Q2gpGIppv4EwcnWJ3I8+C60lIGp/
Vrf5YGx0XDqIMxvgbqEGKdrJ5IFAjHdJm4WU9I4rgElHcmvc1FhYCZWADvJPl+lyOyJcmqvK8+Au
cAsrnpik2mYql/ZLMiwVsq/j70s0cy+HTg13Z607gBMxRqFFs28CBaTeAA396QwtwbOYmryCD27Q
JGOeBXH3ApvTZedWyrg9bKMiXmGYVo7tENarudhSLglRMLLzURZ36mf5Vwcbw10kYjvXHJ+z5ATq
N/dTyMb2Je14r2GE+S5l1LL1DIkMMsSIFui36Nc9nyNYY2+WH2DKMVK+WC/v3ipYxhU2xaL/gDo1
LuJsrVyCgnVsXGo6sN7YMnodsm/WrjdcuG7go3kkCVp/XMdJqQNv6w+6VeUkEqwWUeb3GhR497KJ
bLJHT9SPsyLiyuf3Re/QTnPxPdmce12iF1ZdVV1cpYWklv1ZpOKntIgE7jLP70lYdOJ2w4kBWDvs
/DwrbjEcP88WDYPxN58QTLEerXZOxJuyizLCxpiiDrJ4cJtzwqQwetVIaYCpL4JdN4q2/oTImt3c
BzjsxM2QAHOQo9rsZ5x7j0sG1LefSsgG+M4jRL2ACSMgAtpsfLTnsLgkKw9sZPOAsPzKkrOHrKP7
S1tcPgHgPNX3mxrLw2WvQuNE05WfFkPWvQnuVRZy/rmOzNnlXdS2qKCyk8moJ+/8hs/EPnI4esub
6sNjrrOK2I+q9auFmueG1OyKukaOf5r8e34NbXIirLbK7FLoOFJhrhyfynN+67JhHysLrG2H0vBU
zqlB+0Put8Yr7s2vLIMCrtEmNgwymxb9urgkUroedm4ZHZzRXcxyCCaTtwPlQt19BwqgjfY1cawl
tG7nd6uRD4rZMmO0QK4FcP07gFsE8dQpZjOc/o/ogtEag2LKnLLX5lXjKukmONJXf/xbCXQF3Hvm
d7fCTJP8EmhvYe+N5b+7H6eehPZMIMgPxw14QlTCHwY9G2WkUus1Dwg3fWfBCq58IqpWmtNyS+HD
iCd/mNWcBqTXBkJ5iMrmiIdeE5EzjcZ3rKsg1tK9x6UrtSDD8rkrInS85UB7Jd949dFmMd8WjXpm
xdoxEVy4gTdwQAoDBQwjarCU0cfDvkIJdtsaB0lPYbLQvMjJk8eUhGNuUrwgS0xHMIjLsq8BwMyv
Q4h8/EunKc5SKuH5NfAnrxvyh9dIrYKPG//NpQ907kYJPgZxJgzYely98MnRDFEcThBGqTqxVHYz
V77MUZU3NnR1dxyRsQK0BYIxZBoxthlSzt9kcemxQKrypvloIh6022VUdPXdybOy0ooW3qI4j8R8
HjbmBJJVDAKa/ofJvTtsny9hu+LP+LglgTxB3MWwsv3c/H6SWvR+Dk0jNMkb8VNHXtPOeT60zxVN
9GHZfvYLuJEfFuWlK+r83+BmbXECGuOTKkUaJNyJ8utZXjNX7VFrNbtr7EwQ08vnZS+HW0Xkr90m
UM5dByBOy/QskRPjlI8VTn7Kyhele4+MSKTVPPxP+TI4N2DZfOgN5hb2rLM6f+GxAFYMln+xzVbf
Htsl6SqoZpYOnimjMcr1aV42Hy9AyuxqlERKvGc2fOzxkuiDBZf0sPGFIqGt890TQnsW1/wKpTis
DJ5GByo3DHQmzVGdS7nP9gEE1dXABFYyrS7JSBmXik3YoISYNMalGK+BZJaepZ8l1R4wRBF4eTi8
yFG1bdfABj8m3kNmBAh7wiOBwf6VFsJlTrU1UjAtCtMjE6lcBl7SyqaesS87x/Sj2AocxKOP1Tt3
+GwjyI269zda2B2E8yvQTlKIEZXZZIvbPGKL0mM1idnFRL2p7JFaVZyVur+0hFG3YTdAYy+9vWty
Yn9X0iFV511boQFnkX/7NWBu7ib7rPXJuqm5BHO3Ns+YvKk5Mk0eippiChYjZSgOhemCkvVgd+6T
VPCjJN3e+eu6t1u60AlR7Hm4oTDqTPJCIKLia/zROYMVU0FI3mmcDkFgkDbosj9gLhLxYn5bNNm0
aNl7ct3UpcZxUNYjuYHmyU+cBesfW1+4VwOIcydLGVwxqVA+/ideo4gucwmoScplHp/XX+0+7WHg
c096mBkxdq0Xx7Q3SZmY/odCJTbu94/VnL2tRkchNKUnZi6VbP+FVgDfTpRpL4j4XKniDL0zsafD
Tf3T7w4043jQuBc7sQhfY21U421yCpS54S+A56UiERmHbt7JOS1cZyBDfQY/tTGVududcMyawFaQ
JLq0Y5OFBnHhNM4S2OkJk11t/HUj7VWiKFcJwex7NjlXyqreI0oln2zCk/BOAITa+KumCIAcL80z
Jh08oS7e91HvfKf1hwtbtF/AwuU6LnJOPIQxjT562lH7RJlva+GFeHfXEXd3odJ4jQJWs47tP2Yr
jXa2nOTIMOFBYimApZoDrJjxDXAtkystueI3OkNgQwq2GbFArkKv+/fFm0fwKbNL1Dkl1g11SD7I
U26j8QXaz6OG0C7XhrzwydK9kDe1jau9qQ37uj2Ny6ZzuEs8JvLwVyBirs78VaLQb7fxsHAvczfH
SHUGRCC3U0T83izWCkit2XmCvW/4DAvd4K+HnMN0N2bChth9cof1QDRgKM8zt3Fmju4adIBibocn
ppN5+x+41JxArvUkwSUlnDQg5aWMRYg0a0vS8CnyKN0vIPkrHz5cOm9XKWUDG1j02pVIffEHi48o
3x5GGbK6567KnssLulV5s+qDqsjAWyp1geeEyQG040kytroQ6Lqw/cfx7sWh9R/c1GZCYGP1BgPF
jnakW2KNxFNplCAl3vI/gSQIRahLDYpgx2KtkBb1va0IJ6NqeBNhnIArH84SWDqYo9SiRbBB+oE0
5KtRvuQ7PFSQ12blVLlffL2wfCPUD2yRQOjDTqROQlEjHVxE5Mz1kvalzKgxvsIHq9tn0gnNI5rF
LreUawwipX3AlQFN4ZK6qkbd95ZIhkdhGhL8gId291GLMd/rGRjlUXwZyGrFci1xXvW7GiWDt4TB
okzw77FjzviFriPVumrqcpzobacGstmvI+NFOWo1QdDKLFiTJax2qptZ2fXYaYr2/6Io0B8wz1oH
P7/5ObhMkeEzJGRAhYHnyy3AhavGLTyPdeK03l+zufiuBgSjcZDPR6ctsdZBwJCpqrtAD5GK/iMU
a2VQEUQxIT2knRGz54s/dhike66VXhTc8dYFgmd30EcbuQY/VlFN2qOrkvVfOO3eqZiWDouLUzY8
Di6DP9BICkiybF07hBykmMF/6ra0qfm9nqS7C24KzKvcP5WgSmEez/R8fJdnkxO0KAqp5PuQxh6T
ZYGGUlFom3970r00v5+w0chszSgf8kW3RdMwapJ0HcLi3brWuoFu4WBXTvdn3o53bvxD/fkaHK1D
IBem3SUwvtz/0oenoj5tgsRgMJbIpcF2XOYQ6b+00mg8GRMw6wGif/gXH+O27bVjZcddjN8KJsUa
3TsJCu7mqlKWhX+HrpXKAtQpamGvUsMp2LfXIiGVUyNkz8ChEfCwV9Udf7b04H13iAg+iV8jmk0f
q1dHtcwZ/c6f1jPX3VT5kXQGIYLaUb9qaZWHO3xlb6A6r7zFk+bqWNmN6ViCQOaZd23kRTzR6a4Z
IynAQJ2QroviQj/ftz3BEhqTlKKspMxwVl+x5H7vKPL1/i7r7WC5gZExMwGAhD0Dgcrfo9zx5wF8
ixxKf6QEftm1pNYIyJR+9VRpxA6ltYr95nCScxq5bpwDAgCQL9zHja4uuSQazGv+vUEjwTzNGjIZ
/dVJcEl2s0SyQrZc7xCyxyQmrM4WzkZBE5+nx0biI+i84j1dQFecRr9cGZdN7PIYKApupb2V47+R
1NExRIxtZ2jslI3ZatWYTgx6wD4K6wdamLu3cOzpnE3n1Bx9+eQcpBlLgBDdY+tBHStQl2drwjX4
7yJBrGJvBrL5qzAVNStK9Zb1KrpMmT1S/i1rqQFl/ozqk1hlQqWC3v2KbVWHLhaCydpQc7lp2Z6h
kniMyIsh72ZKFeWLWO42MNz+eNPcrBYZq/QS5vSooWsQv2Yx+A1mj98ULq2/bA3ym0z3hrG4ye9x
NWE3q7PbvUOumSLuaJ6o9FoQQf6XyMHBqGAANezruv+w0yhNW4a4GMA+zWW1IKqKQSW3YT+VVMrE
tq7j9EBbmaSjgIx4Wa/XE9tfrfnqh6MDoxNibxdKeM+xWx7xjY2OoG8cfsOgxKb415f60vzWCTfA
+xxnKdu4vCnYKJmt1pSmZD/6M04mlHuATRc9ZsfvIfjyoFmQohqPR+UcT8qLFvfGnyY7QBxhHi28
BGyfIU+4MBQwj8Ipy8ZUEgKty7R0K6IbU2wybCP6DKZ3dH05hkNwJ0INnv0v8aSpxwTSFnAm5c/C
4ohHJteJjixzswYvMWmdKWBWTOQYdzSDAqW9eeNe0NY5Q6iR5lL3yMWj9OUjSkplUKvVIU9Oj/+/
XIcRym9RFjBH84LQhElQoWGASMNLYa/JZbKx3V7Rp+LNLznXiEk1Uq83FJE/lvWwDW0k29txJ90d
xdqsocfZfSh0shK4qfm4di6it7MNE/NFwFpeaLIfWG/sOoED0SzNOxPdewv6u+3xZ8K33hjj9F3m
mw0vCVGR1FAVbneSDAYjRQMZyjhc5lL0aL2pYu4jAq9Cl9wfYzV++Nx8YM86NdD1QiNQDnqzSAjQ
gIF9nP/AJd6pPDzTn1db2r+mJ54jDdoFJ1NoJKYy7skxiaAwlVVwny0n0p76jBl6JKjeyOZkYvyX
u8PMHzD7wGyUNPo73GH0kNMu5cnjpDJ+TTol130PTCmoE4NHGbLnt8m8MbD6Hyw6hVy9sf+I4sXx
nnfMgSuNQwZILo6Cub84Mf9orwAnG/RAGm97Ab6jgDovJe8xYapaifWaIpMLorKaSxsk04qukcMB
/JwYOGAZ5xgsMf0s9SoiV8yimeng80P6NezOrUV08xKLK2BrBmlTzqKNddc+ST64D/ZiujWfNxzV
pM6Lg1x85Fnq6mUadrpvZiU2gPr9C5GAUdhK+H3vHJNxkmC7n4+gEcEctMjtOSIvl8sLD6ady48n
IZ2wYv2tnk4dWqmYCn/jQwjegOCNIXJN15JoEkpMCn17hh7Hmjpcu5CTX2tAtT61qclstMCUvhWs
pl066aj57wAv4tcrnY2+p5ejHFx3JHtXyGF3Tgup1U9TCMF6KnNYpEH8XFnlrrJR9yzqE4br5I96
FZEtwFL7Ulzyu5A3bZn9yWn+Wwwq5nwYojCxczT1BwZP7Ceh2ud6ImKu6fAhkf/urW9wTf2ELLWr
cy+lOjt9FbMSm2kmFHDbqt4ft3X+Ov8xNeBousPtK/kUWGu8jvTAQmEisl1w5wwA+yky1dPHuZ66
C1TogXeSspsP8rooBNVcmYBjg/Y2zsT9IU+4YCjyCS1BBWEjYo9hFfapMObtK7/1oErwTW3y4ojg
qKksPWbLbhEKrFZPbLzqXFNSsG+fhidra1vSF/LtlKygdd6xTOlkt8uIuyc99VPJSoX5pfZDNJqz
MIOokQ86CJMgZ3Q4Lpq4/HZBN/Wt2U5ODI7E0vkZTJiRrW3td+XMb5njPnc8DmBDB4Bwl9KyioMA
NPGEWAYxjEwDX4ACAKi/T6cpLZ9wdnF6z+uU9XmgaE1Tks210b9df2pxC8WdSOMGHIKanQ6fcYpz
nx0K9rE/vqumFqyZsGQGs6YlemVDf2Fogi1dpCBuiZvmlnDd/cCs8VpI2FNZED5fye1Hufc5+kQb
s4j31YJrWSjV7j2IJbWwGGJNNiQwZgJxfUPvxjRnr9S4wqlZzWPhxyrFhjIAe8bv1Vmcz8LtmRCP
gzMO/kLzHEZmCXqtci7N0dK8WW3wHei/IkOX7pD+lnc6ofZT/FnrTmOzJsSgXAQZFQ3++Ju/u2FV
HXpGRmQiPNC0fqw5h71znepiSUYu4pob+DgpLreB5H4JOMTyOwV7AeL1FroGXtH2W1ls12Rwpm6v
eN8rzSVAcrqgwGS5NwyW0quENMYhdviIZw2quqKx9mGP9TJEQMSHvw72oCn3/UDDxUFFXxBeP39J
YNPx/2VXPZu0eW2HWH3js5Y7HNcp0HAvh8XtMRw93WdnNqRwSc7db7hpy8/hw5UpAWN6qkIAGrDc
9wZjvYLtqxx/dIxTWgHKCSKvw2sez1/Bs1fhqkXeWiIjT2TV69IfSIcfqzIjtwU6oVZ6A79ZIdZR
tSrBS5QvyHw1c9KQQtyQoUaJauR8sVD8RBN8Tv+Dz0xWAAqMBLm5nuELJ8UyfzYbBphfYkpjC7Nv
wyDdFq3+7rn2lfil7hbL671Dwqg84bngVp5WBVhBNK+9Mfyx8Oq/R0Q+CujT9AxqmuY5VArG1Okq
pg9RosWb+0Zn55QhD58q6n+l51QnGBV72UUusXQ+1cONo9jgqo153JE1I1nF63uWHSLGefiNBRq4
kJvXyKpvYufMWZS/IuqipPWATgsBtCllrFr9Tbu7OBOC53yFKmLPlhApWKrV1Vx3nv48ywVmc8N8
UC+yZAOWfA29foZ/3V+EZDlgApyClSj6EmEwfY7dV/ovSgu8My+cZHlT0Oo4nFRjkXBcOJqXq14B
erwOjapdm3fi9SihnGduHr4VsutX+BZRHLoYH/FndWtyFl+O43YOrVX2AWHJz+fVXHffVHFKoaRu
oHsiHK1XRuVgM3CoTThS/DnRDca9bgZ6qLHQ3KnWV0jLyuzc+K2KnGB/Eb3ABiT4mPXm3l/TuOhv
NXKhSvKurV5UBv0T2J3jBhoA3xkyS04gi8MJ447C8c2L400rJcJrM00T5RemupgOSGDIvgHICVx8
cMHZ1LngHrAYWOScIBbDdfvqo/jgPaLp9dF8ItuEXUV9Rom4o0iD2wMIc5cEjfRccDQhZGQBK3tt
rHme9kGz9T2z2xQPXthceX4eW/FlMAHHLzKRx/V4JO0lxBwWDR2GkzzIl65PTPSlzB64hVyOU+pJ
Favm4Vg36upGoWZja64/rtEhQWbkBXlSs7GKI+FD2D0xNZ30cGHEUzrIW37PUM0Qil5jBfXWc2cS
mMhWeObC9122t15V9seFcvEThPSMai41COgJuuHlvWg11tPSbh1rKHlyaiVoIfee+nlOvUZiZVPl
uEOYZtakTOzU2KS62vPU1oQB2Mc7EYc6R+r55awPNafSe5lR6dVme8YMKkBoKY+Ml3N+sY0HfgFU
cBgRflMuxr61kssNnrzwxTg4iUlgGkpp0mhFhp5j2d/VtnpbGTQbCFDIj9cmpoe3PdKWt62hr1Mw
QunCHDyK3vj2avP7wo7oi44oU+AF1ny/H+4Ae26NL4vf4RvJ5YHNKREZw7UZev/f9YDp2qEKlA0I
p2W9x6EASYUKF++i5+XCj+cugNpB3wLplTqxFoFg3ruNdPHOZ22HIzMB1oHsKViqFv69W1pEvdMd
fqUcfun30V0Q7LPLeUIrj4zHv4gM+5HwMm8kQKDOE4XpAGohOXFJAO2NNEdykJccz+0SpybDh8/Z
831NDPGlBhVWZKvAVGp1VuolRgSkosrahYMBkpibx+3ODkb8AKpte4BBzbwuACeF+j3kOF5HI0RV
4/bGF9+CUhZGQ+Enr0r66mesuy7U8lxDCXhCYV58Lj7YCC1OX6MILzgOZ4110przdrouRoFXI4qu
ZJpVaBp0XJnnLTywUSROcxvpA/4V/AFdudpM2XrrPTNoZbDbc0Y0fW3RYL6U4HZ0GV3fRkLFqHug
qiyueus0JVY8yhxDOKVgYMK4GR5pikSAis+uFjHIEzJwkGUMsfYUndiC7i0xWQ2tWGhL7pYGryKP
JLtjJlmhwKxL31mmLlqfx3LrNU6ylLXRneCz4I3VUGTVtHbyaHViyoFYeBT/NRWmwCmgb+9G/n8Y
8VzMm7QYpfbhcza5J35kMnz8YJwKdgi+bNFCD07q38U1WQZ34hJ/rGJ1Z0YHHyrSgPiB+HeXptkZ
VCmsa9SzSx+cen/3Ta/v5nhuJ4eJ9viCczCIa/o4RcLN0VhBoE7Hi9Q1Gbout1CjlH5yti40d952
KX67frjU4cwmbqFOoS1McL+cJPTxuu9GNdBX7YbfNdWO22FTbfeTQikGfAxrgZ4ceLw/tBw4LKQ0
wPL6Ge4+iTfKf2lkcDqS+QJLBt52Qee5pDzb/RHxCtsTBlj6P1egiLThsmYLQ3y4F73fdbhDx1k6
6Mj1Xx0QPNYLtCdhuccrGqpdT7QwH+rtrBXmK3iBzSrTIorJfiPxYL3s+p4fvfDiWFklFKnsMgWO
Vzv4Y8HkmGBWfgDsSsqzPO/W8PG+hLRDgOCZn+9nj5peDpJE53oHyr9ZRy7NMvnyYPMuiWJ2cdLh
k1SyZxBomkOuW2KDONVxr9AFJ0hex8CABkJUwcSKZ265HDWHaEM+luFGm45doiv/EJhC2IQNv5eV
uNh0OpB3SvW9oquslyyYAygtOi9JYJo0JtAtQA166AwMRctVWEIbAv0/EMQGB6oeysGMaanpV+9b
hn2bI9cGQ6dje+zscfuuR2xmZwFgSMkp4lZNR4VuVMDQ09TZCpkeO/krcbOWIi0tjAF6xITnqzce
lDG8rdPlpS+DoUEz30fqs9Y5LsKVI5/70vWsCUt3hwMzTtTKEzvvDiynBNU4cEbA8fkI0vIuiar0
jdwOiq0gVVCVcWJ7JjDfLWqu15lx7MQzb5z0hbpFueJJRoBMw7K3kBCd4QFPoI8x0g1Q6sPNCVQK
ywyW9EvERbtWwPjWUP8kcR/NoSYrcC9mzGYQzrV8Rh+BYt+uJx0vo8e8nRDPIs65Pz6EviZhSP8I
+FS6XbOU3DVBSwJW8LMT+NQg8qry+W+/7VhEg5StPQgOFaFG1uu+5PF1Av9VuucYsLjl4aFQMkzn
aYXKXPnl9f4nLHIg9iOEer2JWMLkf1C8NRdH3lzSil1ExmNpkg+VsGu0VEqiEtwxX522pUJz3FVx
stgVuxtTVQzNF7ge/jtgjETWtJ6fa0uFa/infONvShpmYsTdKYAXLJ1STt3MC5C1arnh61wcGIpD
uTjYEAxGtyqRazGlbBPOIi7XeSviJhmU1LBz4qbBUGaptqUwCd9hfgBo3Ihi5tv28fsDMd8eOZQw
e7KkGiJTaSVlhnj/WEhNudEQrowk+p3JOd4HTlmRnpiY89dSMQQVpCIiHxaFYTtYbQoqQiF7FzYg
k/tGu+H/XIzxsG7GsFMOHyFssCqV8Ciy8hZyZ3AOpXM4XFt0WMongdc0uhCJo1E71TJYxJpYB3Ko
C7qwgKjNuLx+qHOIdFVyoxFxUDfU4eF6oVxZrFw62w9715s1v2G7jwoHg93p+3sBz/CsBOeJkAeq
gWDz08fp8dMBAYVmNV8l3gpOxTUghDDua34PG0H92zCjUl2mTC+GlSgRBM1/UHeQsNDNODvjGBRh
IrUyuyanSjMP0XhAV02JG7i2OVb6jNx8lBag86jWTF6HgS8tEbOH76nS8hRAwMBEr/i/yB4KZAof
pQzUzzDlgG2lr7rJjdakaLu9LC8oZIi9zoljImSB2UxfBaWMCiiw/5NNyc70F56HuNccW4C4yZES
8v4RQC+Zs5keuas/YgYkYPcrdJkx+3Sjsrwi+hMFktGPF8JoRNHVeIMB7z36M+qjlUmZljecaqZd
1NVEN3QFXVQ7qCGUSOmivxJoJgCt/1JspWnnvCMP2ZK+DBYP6/+/s3Nd+mnVaOtsnSDCt6J19Gpu
pz4dwZZnzvshy2+6q4xGAOIbGo2ElVDi92mmLAMEbtXfwP2rF4SPZjOTvkRbttdD0vKMrJiAP0Sx
QWFCqoaiGXQ2YM1KoKoQVMUkvcirtHnLFFTM1BXxwT5ppmcj6s5gaO9VlDz5G+FTAP5o3UFLGEIf
TOeZB8bObOrwYzzG5DetmWQ7zTwujyHdRSZK7iq552eR+8gkZA/1Ve9OZhWQgKjMxH3BYy7LY4Y6
ObNSdPe5IAtTWYB5o9jhtyFXvbW87lOuZGLtKxGOKNvUA5JIMNPGstE93Mm/XuOxp06tXYFRTNUQ
JD+oSD1Jeqx10WDfWfS1QWVAwZbCiwnxQ0hoWuL20BQD81DQumYz1B8WxocPA1R6ciWEXnUY0aT+
KPD/pNHr+J4OmpsIKFX3hDH3HW2BnazCkjtx2vzUPeM7av85EyCq2JS4ufvtmAPJG968zRpXapCV
y2k8JBzSl9Pge6zSdBdzL+Bp1ZGU7eHyJpw6K4JLFojdDQ8aoAUAfng0foQrkA9ezfjdwtEpKDIT
v5edAqOvROl+Zs0P2M5B/SRibBQ0Ax8M74oJF3xNBwM+x8l+yGi8mXbBSUnNb8l+gSHTMCWQCvMs
gWnC8xFCFUFSpuvWc8+K6bSVMli5kAuE4MWOGAhstRyEBdLwTyPpQlQ32mdjq2bVD5aXvr6Y8/AL
dwcRJ1Ne71Vpwsbj1RRmSkIh0gF2MSni6Cis7ErscNMSrRsAgO/Avar/Wv184LuqRgX6OhZ7Zc07
eNthdyZjIeSfme3tp8HAP/TGDv9XnGCRGUjUXcKmUlxm68MIfgzfUNqrBdFagmGNozXdldl3qdrY
GML6l9nw8F+1zTtwIxGBSTmM0v53YZ+/+3WIIWdg5mX+pwfHqbLnqtM6GZTFkbi9xF/I/4fvhrdA
P+oDrXz+O5wrRZ0peF4qYQSoh0uB2U3s8MHDVvmMXS7Y/iXq1qG07GNdri4OJRxIIpVKYllsuOj1
Ug6s5rEAQJ9KyvPqGa8FGNqkcJWlJRxS1URHzZTzfQMIe7Zv2zx7aa92fdUvZc1RXvKjRSfQBppU
H1E05fXj8W74Y9O93E9wReUW3azsV8BOBy9SG+blDpGTCGUd8LDqyNlQUta0u9At5BG3UQYw27Ov
wVad+LcvwYVjaHhMLykR7f2h268/xb1gVZxyXxB7cZW7JF3uaBNldPfAUSe/hkOVaK5OEsjHWfCj
ySKC5JHSvjD4ddoS/KJcck+ZwYz6zBHvIYfbXMcQgK9ZOg6Umhv9Z6QQzdFbbwwdkp4aFGTRUur8
JX7wAQFXOj0hN6Ybj4FsFWNipiSoU/onWqeCZ87o6tGY4nv7mhHeGsHN3hOTvQJi7nE0PvEACu17
CusXxA4bRx6jM5HrzcAbc8gOE5RthRmZexnXYaYihKJo8vamBDVNAd1Rg2H83z9licJTi9aO/YgS
Ug61s8ASJZaKmjptq3if1/mJGDxn6mQBcVHieK6pWZc6c2CKV6hE0YxSWsnqSDZr6k5Xf1GCMIwf
4iM1++L6MjqSDL+XgwK1BGxYYi0Yxte4MZq9XMt1Y65S+DhPduHQ/fC41hfHHYhABI+4kccn1vUn
B/Q0GCt7Z4CVtZJ8OsZUeFmri2OVnmxjLHc3pZ0lknFcKSfxruaDF8iRI40xPn6nQA7iV5LN1thc
aBJLoPafpEkcCDJYnJ8UMVUjhPMMcqwc5hr/u0C/d5B6X4P27K1TBX/ylPvHy8NGYZ9GbN4p3qEe
uBp74vLePjTxgHlEmFMs7xpEiAQONueRVcOSChKibqIgSoFnF5H9Fifa/PAUK/5epOXh8ZRTY0CK
7JBDZ/6nj/+z/9RuoSM3xRZ1syCHGAq9KhI2Bfah9F/ZLb+N05aGslNgIgU5qFlEnBc6dnXERoDx
oLGxgWMUfnvmePNFRT3JcPowO9MmVa0fIGgvU7UbnGApmwSe/MFFMam534SqFHhef2kIOC8/XKmW
LlRgrtiFlapHUZ1KjOsDnMpSKepICtM4BCsPFwn8s4eOV4onAR6X2Aa5JBKhUez1TfplrUWQHWdK
WlKZuge2zwxoWtBfsBeiNVhY7pBHKOIxGwg/t97f85+A7HB/Rnq3C4zDl6Tni7GDmuvczALqnlU9
iVDeAzuYJ1X1y3rejwslJpTEDNdD6xxJEC+PLIJ7lRB/wRjgkqfB3Y4zIqottutfJFr9nw2f3VOU
mfT9m2tUrnde8NKejcIEaxFFPnMnylB8Lsi3/mTn9jnErCBMixnEMNEplxpXYIVm3e42Z9cu+iVS
BJrjUKSf4XDEhES0k7eKCogNsdagFBoPK5xWj+LyF5+HepXG4TSes3Tw6PTsLB1ScGGidy8/GV1n
E0M5pn6r7tbMaqjSbhj4slTxStd0UVeACVh5c8cGdAF079grj0+G1w5SHDuq++g81+optu0RzF2j
w4ACdm43BclxB4X+v8qauHx5bm78fnoQaomGeFJs+9hhjYOSfbPmZ1m+H/NlvrwyNGoOQcuPUqdN
mfnqANLUXeQwnLErKxmDkQakZgJ/LKikUcQGE3PJ2qzZJDB5sQiazUR3pxGUuqAKhUgPqC+bDD3f
eRZNGGSSexE70gSN9mQCrjXkWBP/ViEl+RenCIN0nsCpNeQ+pZcS+A3h9pTdBwVElvvUTQWxn0i/
GCSKw2lItMt9Fz0PgL3yMZlw0cvwf4vPiGeZD25XkjJiuqnRBZj27twY7s4N5XoFv/cqmMvkQ+x+
QEmHmmxS5fK6f3O8oJXYY1G0V4/6QVVMBspt3ITw9RzgEHHl82pRosTX9vamAR/WHRHGWb27DVgq
9QROX8pGT8lmSpifcZr3l0M/FCx9Mp88/1KKuoFsZWMjdWhCcDct6punTEir1ttOfwYbr9IN4M2G
/IR9IvU/+hLAiJiFOrZhm79bkdUK+FEkiy9BysTPCN265r6Cua4nvQ3rc5gk9ZGI3m+k6XJj5wyj
XmHKUpiNUf78upHX39YX0bq6n6LoVRWbaYoW2FKBNfQiUUN7g8Q/YZNZi1TfOmwnAG/2s+hM1v4X
jO0tA2wQJyfKRHrIVmsLpuDk+4JHk7TXsARGRKT+87y9DjkfaKMbFwMUOZ/P30s1+2tKUC3/v6bx
3YFnCaJBVVfWJnlCTXifdFzzcOAlAyY/28z2OtThBUbkr+JB1GiwNnZlBHgMQwDyNJoaaXNSJWxn
R+EyKZRdenfDQOpjeyqbGtGthaPRi/w7/XZRtMhtu0tbAfxawhQ9oJcpiuB49OWtg4RL857RydaI
zJuPSbzMRSyrG/LQ3pFBYbLWqfZ2mJAS/JRcUuv4bVktM1liYsanP/HrJH8/FVCaqkOYHqGkgEf2
noO6Gc1weugOeLAorsaHQnYOR/t3O/cjNM22toJ7r771fkpXzNH6TcwwtplknAy/s2L6k3J0I9Yf
sVLk9D5YAv/PKa/+W2F9z4Q4ztkXtwu6A7H7ZQZeB4ESXK9tiv7VwlCBCGWvTIEqyYx1CIAMR/wS
PgAqPjGY3ap23jmjL+2Sm+jUHrt2J94CUa3X8hQ8Q/gfH1A7tuaeyeoHQ3efHKllyoBF/bcEZa4G
aQnjternWtKG1c8rzfA/DgcvYpbAHE3+w3vQhd+InYXUpYvsbSYOi/3Ufk96sFZ2wlUvtdptdL02
u+zDTpMBQSL1ZnYVzaDgpAfMF5CYqxXnHiZKKhE3Mja7as3us/3L6OjPWX3/ZNMBT1gdD+eudK+d
p4vlnV0mDtjn2Wc2QmGltBbJ3D7eFl6bYXIyG2ceMQlXhGgyQ1gPVchNvUNQd4ltQbmTaUc6RP/P
WZwGsDK8mjm0T7JWyoexdLZnf6lAk1HZnxgmlA8OaV601vrGeonm3URxdKXYfWQykH79c6l/6eqw
YZKxz30Q8WwGF/L0ObQEGvAyCzfODU3t5mxJJTDByYbb7OdpoD4ies/1LJ2e5ft6st0CSgD27GDP
u+Jz9MB4J01xWOHlK174oAdOhlRFKzZTB/bPgs+ADyrNHW8kWIB+Igplxr2wno3A93WdXswk0GIg
KdxTTR1JrMq9yiuOOV4v0MmqVhKEgiworQn7CREcs9rHjUxnAzeqUPgNRaNIaHirLnrwSU55/tfu
xTdRbvJxNv7sgt5KMcd/2tbb7otVXe+n0ckNsuM1cXPRWRJ82p8768BUNnVl9edq7/MnEh4SVaad
J8pg/X0dao+qnT/8Gn8j/RbrTX4tNrcm/zZk/fuGkhPGZiDeftci/RhiykcbbHiCh1Eogx51tHmX
o7L61O/SkQ4Nl6A3E9EB4x6mtp70oDP9to/FBPwCA1uIPpoKruoilBXxPBrWtlKUobNnTNPX/DHw
4vVvqyZaAWE9ItT8WOFfrMYCrgUR9NfO/x0ofDM+9/kXcaJIHBSSWn+MiO00nOBbHIgxZaWLzREu
2dvsSzrUWs1TeK1tt8zvNqVIeFcPjOowmk42UEQ+O7iKYhR66Tgk97SAgF9jjTlJ429F4y8OyLut
y3we9UlJpHw3Co5wA+k0O7MY42KpREGyU3y+0jdZ72kv9BG/ODneVr56XbA/jbYf/HJsNCZA08N3
5wjhXh3dRd++3bKc6kda0+KQcUSI8STK5TpJVbY3c26X49hZMJLYn6RiOClyANeMZvaEcpSneC2/
SvhEpbr8Zxy1MUaqwQB70SNFvcnhL7JZZBHvB0AOWJnpIoszELffNAQoEbnl79a0A9BZbaPyxsc6
DC0vGs2lPiaF+oScfcff3yPdz5krFoGM3s6hhdecLjj9aImZnpde45G/c6cW/QIAy8Zl5SlsXrGs
G+W+xVlZ/yXryhHlKS7TcW8Hh1sJt19D1HGQtUb4t7mgwBvGrekAAveeqOYi4dKVXWpRoBKbV1CL
evl7rv/13f9wSufCYKLcZGlCHkhP/hKm5EAoCdzMw7QGPdAHkFBEwPt1MPC8OG40G2Pmo4HbQBsi
0N0NdenZMHnPltQ10XPp/pyf4nLYushiCK/DhzMzBaYoMFm+ZRbdolTBbuHxhSqS7dqegL9R/ACu
pMo5ylIkr2e4FUwz8P2USb1IRfyP+5rNg3hsiDiykvMGaysXNI/ZKA8IaobvC06WquUhzdgvqSw2
ma5eItGaByfB9bN7frwCldi8npTkGg589vv03Oips2zZq3MXKe9++JRUVsjskIqB9+hPyUEsgPRc
H1r2dFZoYyC7OgV3I3ylaUAMRXg3a3ya1nQDV1J/mhBCzYcTyHQCM/cq6Zjo0bYD+XHs3cZN0g3a
cVxK/KW7SRkSB3E+0+c4a4TJZeGuNGXEEprSW5ZKaevgE3eR3T75pKkA3YhBNlPQIhTV2fnjFKtK
+PYkzPwgpmz56zyotTW5DOJFPiG+e0ScwW34tSnSpdpU/hoXb01tiouOyNYjY9UA23D4o3SPC3SU
lJEDV52JcUCMOYbj71mPNjdETweQP3lmjKaPDTXXPQlqJHSJzSXGvjnXu1g/m9NU1Chg59Giv5dr
8Cwtjt1B8wRaXPKfK5WK8yl6RthJ6VEuJxyMUFNZ6Y8Qy41h9Ayr+CXzxPIFWHeaOMtz6UuH8YzS
uYJPLH4j8UcJ9tWDg/Mjrs7ikaDCtRjBFT4TgaCy/BZlpBt5peTX/5rZE7o3qGAZqQ+jKn/XPZmR
DM4a5xFbDd3GV6zi4aHfgnrRvamWx6MC8nG9d0JvohgQzmd23yCktKgexUNOnqR2tswenBQtT39d
jP0J4Ixl24qnSxdwyGZbkj4aMY3PbcMJZRUOBv34Why8Nq0BI5jBNOW5uRFxN2YzpT/9D3m8bKmj
Lqkxnf3jp13m5sPr+/tbJKpoG4gwEU2aoR5ZPBr8J1U2swTWVpRDSL+MuGvqCIq9aUaMwAxverql
1cTYDGql1cij9paSNUI+xzxoGLF86a/jMhZxBVlkYVuzi0i1CWPSZqFx3qKdGSVq4hdTNcv0/bJh
AtDwxoYCkrJBug2sP/lGx9NmY1qm/8ZEE9BqqPGU/kuWkwrrb8rLS09J42Jye5nbFGoUzrMlScAd
lc99VcvMqmyEZeAFBJ1VVIrzWdO+d2DKE2OG+ZYTlXrA5Ae4NQBn3sIK2EVHIBShk8gzIoEyaF+q
dHfunOeGoKvJKwJZiJmyafY5fQzSYb5m1WHfBrA6ZeWb4yAw5eT45rFKB8ARICG43MExJGR/Zjg+
Aj2RWrttKMjCkQSj1b7dvCxq/gAfwbFmadHig4N8vImeuQM9YhfgDil9pn+mtFKyFU4pzCQ0xFDu
awUW1fTQ64cCx35s7f+F9zCyhmBAuUazfis/FdZ6EIULsdjI151mjigjsFsjpu+jIB+ZAXlhfbGG
kNjZztmjBj8wArYp4QWf+NBQQK6BDmKJoljiIBxmKZmkulQFugQMsTCuhJGY1frHdxNinoNvI0Ye
uN+fKeM1laPX+7yYrQbVavsaO/gxCEDIw4oyjTGNFLZhfDBcMEqjLgW5sk1XiYW74K5TQ6eF1baO
zfV2tE14m2FsOvonwxTzLT4vJjwlXCjQF6DIUhx5JVMsG4nYZykf3Zom8L5/6icdpKOwtK1CqDui
CsAOvT9rr9UaZu6WsZpDEy42yoJzRGKwxog/Yz9r4VCR8ULzAp5G83Q015VpJx2DP4ILvfHJjoyr
WeTv6HwpA7sQt7kZSSe16mnTuDoU/MgxegGK22q4ZybpJhANg7OpWPU7QdV+K4eCWVD4JtTajyoE
b0fqNy0Jf15Fda3v/8QNfcWL5QIFfdcNWR89aAPjpJaL91cwOfxC7pT+bQvHZlTSISbIMeFfCBuk
cWQ0qdrHXSPkC/NClUmDnS+ugBirBXMpF5l5A7NcQWcf783NiHw67WZo7XEp1OZURgLzPuPyHEuO
gGwBbx2j3/fPCbKQddTRCmQkTT+MwkRlw4STPuHYgyKDQ78SRW4qRSjH+Hw4soGhuuAaEx06ZKIg
DFWqMWvVrK9QQxI0MtUBvvdkVcnuBeHDXGY7oJS3Z923fnGtLCXp+aGWJPRQpQxtLckIrBioCCtd
5SvJJ7hoVrC3ln6skgNqGJ+TPbHmG3F7Hg58sWIOR3aft2oZvGD6ObAbenq5fTdQkypq9zoWyK8A
xfwugvW9VWaHkQUp23hI8q9DqUBQiDqycYWDETNg809sEzonWOFjKncqMDxkr6vUbLqydgD6AXx+
faF3z8MiewV0gYoIDwRsc4XGUuHbSBhVb2wDWVIjdbyUyv9Gu14L0sNgf6LMuPs/9U5RYspyW3JX
zxh0ioHsIM9c7XY+J7yVjYxNufcS71WDB3zEIAk0bDHobBQIri9Q1v/ysf2unKvZlhD/zMy4STf7
gk3aNdJZ7S7diSxj37gEbzl4RXKngGwsZLq19EEGg5x1Nx4OiP0QAEtscZ+NIA7l9ljAxGjE/MsI
yxDkypTGx7cKFMdDpUoXTw0+Bi/pm2PhY6cwwDssMF3xI5PJq05yv+OQLVvdJ+7rqObvo2eETpeg
G/Go4R9AgOKAEG52FlPb5H6uDUCWN4yhRjbrWTxCgj6y48SHnSyHm2Qi2o8kxi3U2Dc9Uqy6ivPY
tO29x30T08bcdDMnQEe69LVwGziI26htcziG2rQjoDqrRAgoI//zPsb4b4UiuOEBdZ8+FfgG0Lx1
yhus5oSXN9ozO6rZbwsuTTaBYw7yV6jf/0NG73Rh6VJjLiZ/kcFRuxCQgm8ffxa2Ag8do0Zxohax
qpdwpDW4tpcLYGIdkN863C/aC9KRdiUhj2XhU+0O1TNFC5Ke8Wns2cM9it5lNMrXJCbuIVXPbfjY
O7eiZF783VoZ+8x5//qHrRuX5krO4wN9Jo9mCOPv8G4uh24Bc9KfmVwOR4mfpwrejWDabO5ORFVj
69aZDnwilhNXF6VGvII6eFW7CQkJNPB95dZ1vvdL7JRRcIqhF87L9kXcckVcq8VueE+drl8Si9/o
qz5D4W1amVmZCpXts3pdHKKN69rmlrC3oMzVWyYkzzT68vhttGeIErg8yVk0k1vdcat6k+PMOuzB
IF+j6LSNZprFGHCFzl0+3SNvdgNySJAOIlZTydrubgrh+l9/j0TUfLMO9tuInIoqVsg1YQQ2hwa1
V1Q5EZF836dPGKk3a8NDEo4hFcaqZugcdCHm1XovDQdvOU35I3h75alUJVyaBv896Fa47dqzG6yT
t9Rz6Es4iWjmsheuYzdIEJhNnj7+m8w2nxVjEf9Bb8kI/uSDZU0CmSKSemrw/wOMpFmbE4HcuNjG
+KVri0jI1DJ7UZnOQcM+x+k/xNpEz1WPZ2IRZxNcTTX41xQkmNZJd2EAqdHsGJ3ctAe7H3j3AX6F
LmA0d5++kOh6Lx3sQXq2CLKxkRqI9eLGPtp/yZqCgdH64nwMt2ktFUpK5tMR9cyMeRvXM/1Ry3nC
91fyaTv7qjF1dYSl4lwNKnaQz+xZJv6vu/hI4WGxiez0POtfdldSiYBDy1tR1WBOE9953s7ObWWp
WkE7JnhxNWb1xpGSxfsKeo8spnCtrEymwx1hz01o1cHqo9pYKlq9gvF9a2+LTuZHE1Q1oPf2eeZE
W8D0mx9uEvO/tI55FcSKYcMvMAPJnjLJNtT/VBXNXOq1w3a8mmpSI5gYhp6d84JbT7AvZ4dasyQ2
F4SXEHV3M2qGCcYvIKHXLzTryIwSl9DPSWwckG0IafBJj1fQPSaJZDIgxHo3MIwPeWsGHoVxmH5G
c5bgBwQLSiJI3ehzkCQ8WaF3UORZebdsNYu8knRji7x0WQvRGBUYaoXa1IgP9ofDQUOgqRKFcHj/
YK+hFMdODBdUZdHKDrneREBzMQ1oiHh38yYHiqFJjZ2ZPBxp3D93Kn/G7i3LNbr/PzTLQ9gv0dOQ
BpKaTzzuSzg4+gPO/yhmq1/R+76P3K6+qfuojr2ycOxAUnTTs9uB2h/LEKc+xl2uxSRd6m/1lGDf
Q3DZfKYixas6zv6SJFJcVTkBLBxSWIwXd1C/4Lbk8LAQZ3UV//LO/WML/7OYENw1dk21fL6UCuvP
dyr290FczMe5/Zuk6kGRWpzNvWL7SuWklHlcC/lwVX7Ws8GmE+pcw68maHgFsk/MQz3PT1bvvW97
uYtC1oeEKoDejwGRaJzod8tM0jb58o01yvEgHW0BqpnXQ3OVIxXY7XaAr+6KPvF2gRvhmQPvLc8i
mqiVTKTqXbGJeK0ARn4rUiettxjlSkx5vkUYt0uMcrOfETOJEzG6mU00v9DcAvk0jMtruXNXbsky
4Gu1cjDxzcU3czL9FEUIV7qv/OxsvqeLbPl70C/dUyCeuQSDlO2FeHLZAKuGvo8USmXF77uqtNhQ
FOvMOHfkoEY+VwcoeWYBXTvkaWM+BGZyz4VBEFCQdyhLkN99JrcrZas1ceFDRKil8NjOj7aMHbq9
26yPhK8fnk4YbS0HQ+8yOqItM6LZYLA6Z/8SJPsr7HerSKXYgSrb4xx4ARUMZ6wiGNNgDa+uUTcI
7osHEweRVbm0xPVSmXQrftuN2Jb/h8pOEKbZ/jc4fwoMN/eGnPKqxEExWmqSpg56KdIds0fCSRoK
vv5LGBPdWysjapkbarJ2PrFOkMOjFgKrgn86W5mbYEybuI+1PxTKIxWyUotHMiQ5zFZVdxbEqdkZ
JnfBEU1ZqEdCBsnlzqQVm7GIzH6QhgXToAmnxvb7GiIC4f7iipstgPU8w5Ckm/cBVdGO9yxn4sPY
DikmA1n7dwh9GPMJKvQhBL0G4HTT2ToJfa9U1wK9BQIXDzpYLZj/bNmKT0EnO4io0iEkxNkrRoti
teTwugzn7BSHGeb4QNLKldgdEagQccteHkx2o9X3LM30f9Jvf1tG/VsrUVpsripiSddzfQ+nni7X
PGWlqvNF1ey/NUjnlLgRtfmjZ5ggJRvGjKhloAnv1Re/HEKwNQo3fU51B3ZsMpv0Zzv70UPPrkmC
xQp1SYqPLMD/XPAo63C7QOiaH7RhyfTNIlNoiQRA4UikxEUoxZJIek8/6wGVD4TmeFaevU09dHFH
CjrFxiPPvc3UaQsMOmvoB4Aheh26YCSJH9rxn+OoNuF03iVcHI9hVDOAFXDW+vMaN57xcFdkEs72
8Fl4pqdjwlbyxaJ3BlnrTVDtcIhiuGKCL7+CoANj3GEKXZXY0diYj1kbeM+eQwUgZJreC8oo+JSc
UZmcBNPtCjYrBvyMfiT/MzjdnZoRyD5TWsylmc8bqibSP+JoZPmFs66bhCeuxSdpyZHpQdJjQRkB
N3ahA6QOCMt4QCkpr00aNgCdVliQHTAsOS35NT5NcE+WTSkpG+s1mmk8hNx/35EZf+X0Kh/5QmCe
vFK8yHASQjc1RmC+pZSSemF+6aWuP3QBNaHXQUY1EZswtpKKy/dNSdslILsiZR0KT81G4DQvwvFj
H38RemMF1FAX2JTdmYAz1jdFff6Ygu8BF3IX1n0ShJe9LaxOMqQ6OFrT2tfdr9APKRpmp5uUgy+l
MYucIcKRS4YVn0oMOqrVLiVHX9SSHsRllOongZv6VuRxe1LStuinfD/CwXbIAkPd5C1B5rmlRua6
HoXA8y2TtqCEljJX9Mks84EXp/jDEquROdBKX0uGrYZIpvJ09cUctuHmysj9wMloiEy54GgD9eVA
+6yvs9MFzFVxn84GUSPoNg/4QFbDzTD/RM1AXwV4ZyEnMMUiPJibmrooJMUQrnciSZLlnvUMXILi
IGHg+3sPPmzfosUmA+3AJzohAxcmrxneZcgpH6C9xwCxaO+cWwxAOUGWH44IN2Jodc5ZYLCDwZi/
qnEgtOrYAlKWr3b4m7NND0XrIVyBKwXs43MA9NEfHG6WlYRfO32HBv4U97Hx2gzjngwCudatJqH+
Za94yA96D8oCT25P8c38qX+li9Z6Y6jXvyR6mjtTUnlvK8ebP0+mn+BuQ1owcZyZzKRMP4RuW4aV
tCs36HpKPH0kXoc+TqWxGGVn2Vt0DcBdzkxLEzLZIRkPrlKhabT56/H1VK5gfyn6TLZXU9shu+fs
Bk645uoLqyxN1VSeerdxbWC4NsFt7Adhw2NDtybm/cJk6VXYlqZdezcc4xmFLHc+VyqJLlbxEilV
lBIdT7yNSypvgSr0bN8UJ9JfjKfY1KV8Pf/Zh9qIWm1DdAa8xeFEfDFRFi61kcV/+2IdG/wIdE77
QXtYo9psPQQSshPMUnJVppgLUy+NB/vLAq9A/KATt50D3T/xkJDCMkaeyihjmPu62KZtdATLK9RK
h0B7fOdOfXNy5C9HrMHGXr2RK2lMJ+9jIbVEtC1irzcuVPXSkZwpjeqsfVDBSIFEKXYAHiE73kRN
qc3+2bVr8GrKkdo9HEBTOzuCyS16rU4n4CT8fxRh7QxrbfCslv8HAyED+3V90AM9HFs5QraisBjZ
HZZaQY1Q1LnfQzQ2bfxhjD+2qFLkrl26sz2KzIHBeu661DfcEIonJPgz+ugxGkkNHpV2OCM/zMCU
+5LzyM5HQOg3nIOeSPzKj4TjwNeXk5CK+fDIVVwO4zh6RT0YRpP2Ooo1JkCttx4euTmWQeOjWjhi
m0ANrv8vjGfJe6FXw9V5sC2IZ8wIpM3Upa/kbZ6zY/V1cCdtj0OjfqJqiAI+hMZoR2GQrEM5i1v3
etrln9uNXmP3ANw0zFSWjknn9aOY3yjkxer1Yy2eghYIXfne1Mw2GDIaxZOI/uLxUE1iaz8F0hBp
N1AVXc4JvZ9zRiw7N0pIDJB9VQ5GwiTIhvm2jtArTRZG3YxCPsOS0Wb/d/uKzxmL4bu3+9cFF2Ge
Yq15LP5YnTwYjEtNBKJe7SjbeMtF7k++SJE2wALCkAY5uDfBuCIQoXaFss6U+FL04Sp2GADOHxr1
guepwJFgYSh0DYyxjDOHab+e7p4yNwtOvie8qKg1wzWW0ZrugrQt1yRhHU4qvQVCQAleup89tMQK
ZP7Ida5JNtQK7PfS9cBaAQm0yPHeXapbFxJOxaeTdw+Qv0DGPbOJvCqyWwE2j7WZ1R8n8gQKK1vB
KaSm92MBmncAssrCDmajaZmsWqHrexRrH/w72N31PHJnlLrAzdz+GfULPhPSHRItjHiL5F8KzLah
lPWLZTswl7tkFJUuMf2ZA4DZATm3EH/zu2CFLGWGtEfyq49NPKPJ6iKWBcFBXs6u0LtqV/XjOgl/
F0w69BA0Z6AN6SvhRnZdg0Fpjxx+pGqVxW7a1XpEacLr8+bhmA4K/RztXRNkWZ7CitU8aDCmD1O2
D7cKsB7gVcqucAOVhF2inotN9ou2Cnk2mNTuseotdUuP8q/+eSYzd9gKlgcEFjK7i/bt1NAjyXSe
WYH5YMZUI8sxZSgsToO1Ppo7PcScGElobwtyGgJ3y2+Tjf75Y1eRn3pNAPJkxU7+vOSdNai1x1+m
+WKjdBQhJU9UV3n8vR6NlSy/yPX9eyoC3PyCasUvZK+804hIxIqzlTaWyQfwU2Bgt23xEVYx7tam
wHjgP/gp/fb215RpVRJAqTUWB7aSxPQgbkl5S1K8JjzX8oXtrUxFUfGPTAd/zNPmIFnMuPStrcFP
QSSfTpGV6q8y/Omlq905/KK3XwYwSYwjbJ1jsfYZcTPYPU4nzbcMFTIXR2+zNKrYF1lFQE7KEsMz
+M/iTK/WEO27/S74sjG0FyzaQxNauZvpk9OaSKZ2qz2hWPhFTx9zg6Pz1dpHPWcQTqADXz0Snirp
LcO/uTNjjzMD4c0rG8H63xiK1sOrPgIdKTr7Ce7gLfEy/GKxbzOdQ2uUS0jRLfOc+Qely94t4FWO
xkkKzlqIpL/QC3y0MDeqq0LCMPn7Bb1qPB/zd7NnavSTDWMPgIRDBtK1+349/yUU0oNwVjo/y+/y
+JRM+8hahf8bZ1MFbz4whB1Oud6pcQwkVUO99arFZTC3BhaLeRRzpBZOSUuW5bRY+PM5mLvGBOMO
pwMGDqnDUFWnZrnEW7GcRSsiZEMbQnSPoD5w+sqMQj1LOmUxOv3Inz0BBoaHAI1xXO55c/Md76u3
nz79dKIMSrMfE0Hkpm743MIk+6xH6ronjNsbhsI3TM5iGv090ZxzWo8dsVzT5v0k7jehmoiS8Mup
9BeWhygkSB1K5arNFTTA5AbguAsPUCgcKH2wCrmP0U4CmsD/eTAt+tVc0vl8E99DZxAtiMzl9E3v
qYg4RBx6dufmAwE7k0SmRMW14tprB0YCXK3hycuzAP1pupn/WqAfe8oFRJcp7gRgPnXtYiHQOlN3
rjJNmxBDxftLD21J+CqRtN2IMQ21s/o1Sw65E2NDx+z/yikzn0aumWTaIaFeU+qFemWcYkE9+/I6
E/l1YuedffQHNgV86sLDmyfTLPnBT8l4m7s9HSt4db7ILNUfjEbup1Y0U7gOObwQJwTzkyUbKcyI
2uMb6A/0zXc98xxVf2iwOrQdKVqlhGrcG+JqLzxM0YMeAernftfqqBRxV74JfKUCfbIq/1+D4MxQ
Lk2NFzOq/iKNGE40pNur1v21kV6fXAJvCRLSIbxzpnIQmCidlp99TdA1ZGnYTf5ObULj91TOZ8MN
kW6xP8huXnCCaMDJiwpvG6DC45+X1pd3ZXgzg3+VeTwUoiGJKmcHa8cHlh5vcrqOxYHr459OFJGP
9IOOyv4HjFNHXjs8ra46k339cdvMlJz8LHy2PdvZacyq2l+Q13FZitXODNAnNz+WfMPzk7oRwUOz
9/RyWZ93fkOf4ovjiz0LWGq93DtrSLvZtoU3w0xgWuU2bFByq7CRf4Bmvv6DcNF3L5tICLtyt11g
7+wnW29W88kR4Xfp0rxkyssQADQiMlRo+KdJb9gmjXr5wjVHQF+KyTTToM9KQrs8Rw28VySRlGe0
2VHY5YVjJ/pBbjDxuJF5v1xKGqXNs66/QT5G64LPOIqFn5jphIAv/pAsxfrup5Thg+VLhsoxK+lC
cOF+XqhQkJ+D0REyHjNcHHuMG2ibJJkNgOmCLdlaxa/yv8nGURoSYjyFDQbzK7/iZcWpDtOnOSyU
GbzGOws+ikyfm0rTQ3y28NJZuN/C9oADxxYV4cqyp1qUty2GTsZGTiuMnekZ25PqEgvpE+tvq2/1
n0YWPXpSGjAk/Fkik/4+PiQpYtLUlZwlV0vnD6QMVIbe8N8/7Cn/4EtUtSwgOxuHaa70sF2162B6
mMPM/NhygwwwFobPKteHk3tglIKOdRS/FvCkEr0xKYHldSHoUhs4RbO+BfCj6J3KeLGTUYFg1pS3
l5SWEoMhlLWhAU5ne7GEQXv5Y7lN4fFwQSI6wSBVMoPIvi5jaUz2RFNJ4UMEY0d+X0N8AJcm8spw
WiFMPiF0AcVROsWX5p2ryglFlgU1h8mJQzTeO+rs0LJdFzzZwFRE0+k+ZcmFCrGGghdqR8Y+fcol
AY8+YLUFJuTAfjvgWGAvZmm4QhpD3LoLL8s05UBLd/xWdek7YPFRLR2vs6jTLvK+tZSbTIn1mStq
0A3iFlBYEPllcL54nXOvqiRfkUfOIwtLTale24JQ9OW0qGlH+aKcdXxZt9NNO7xLW7orTJBoL8pn
PGbP7e6A5Oo1ttjHgeU6V6I6Hw25rU5iY49p9hKWc3ysz6uD6Al7y9c9XWo6mXkbO0Ilpty8mbU+
2IovsrOmStdeMGoob8T4NgbpdjEasurfJMznB/Ol7ELiGcjvNjUyPnSmnB8AJk9gvp1QKSojakWt
a5vzNQ2X+suvgJlMyQMDE3CFS7JnEOkyWAUsBz1uFKbHi29bAvCJ2dounX/+gfRLJkN1DAw3HiXp
TvfCx1z6zzdBjKSwKufeK+C5Wwue/aiQDadhK3MEOLHtrZ8dpFvhawp6cAZvE2xwn2SAfi+SDknZ
G2du7pBotHieKy78lEgW8K5i16VBths1MVYrzmKP+sSt3FWWK0TIPxosykr1T/77Vdvx8YEP5N7r
UebdhSY7LWoydcDaaYZYzp1LYhPYlWEKGBl/5mLj868Ydw6YQUjwheyG5SexRiOhWfyuC5aYOZTo
E3yONqwWlBnzZ8sJ+5X0Iz0CF1Mu1WQYI83QvQ0SVZ5NdJZd/VXJoDOpyH8fjIwSBFVKVUdzpfye
NkKMnf6b3qFRH8hdBZsK8nsK1mP2OCuiZkqSiIRogyAjk4/rJHT/BTnHln1O2dejuhwqauzSt5EP
hXJJTjDi/Xmk2FBy+1V2917mZmSotthV/D1OYJbn7nhgtWfjV3MffGXsnW6kCnO1rKn6TUn+sJvv
s7LNsi+YOUvUeZRSkAl/QDnMihV/zgXL5snX6IRE6N/obJpo/lGzyLSkhDMQIjGE2iVKvlXCXfzu
WGNY6p+chxuBrByoyeEE8vJ2BY8E0F02cmRflxTAA8jR7MH2lifG7RbqN/HtHsfL2Poe6ySDrOoB
g4QwjLP+nHtsJ+oX4B4D0m5GJtYDZotSpzKIuIoJeXW3z/sMkxAWEoZWcnLd0Jd7uuHVbDIqonZF
VZc7SnWAombb/kbMeRVf0l2JTPylCafQpsqQSjXcVNyfKPUb7sLBfqd75BwYGVb+/voj3QNbOVdn
tHxK0fObtKApwepmT6MTRn/eUzytl3CxOT74CFbu1N57jdZf2GuAtes1mrM8EVsb0PGwsG3k+znR
WP0XGQQgo3Cb+wM5uom63Pztjo3OePc/1aPCGO6Zxah3N3n7v/9XKdCsXSztOQxa7kbCyVJ65rwF
VMx2sV7sYDLMZUQgtcXmZErW0ojuWWvHLGxXDYytJ/M9f1KiRNcuxr37Mj1V8h5kSgRz52NtMiN4
GXMgFjXbeIeYS8HZ3UUPP5zup17GzXud/v8EF306ZdZqr9LJYWL0AU9uFpUeDzo9dcT69GtkMjpZ
lmSK1EvtsFRk24/84TVAlPn4RlSnaYvkOenpTtbun1oSYiPFGe2473O5ZxqzcKvTlDJ7yLEc1F6B
6jMKLoST1yTBZcMn6a2IZz4kzq1mRqXsv96AgiiBFaSfulmGbhn8HomUByK3UoOnoJqbiSdugiZf
Jc2M5f70YQ8kh3Pil2/f4pzWCOPM9CbqKvVnpbLq6oS69/GZKxHKJZ5LQAEGt0vT3hwpAXhPepS/
zLLMYOFe6oTuMJ6X3Q5FTie7bPC3hkKjG9ualJZZSZvc1tn5YU6Wxxl/EhFIdkzlvHjBnUxJdhmI
dJrG72qbyEt24XeVPRuMHx3qpc9Uvk1Ur6T4Dg5C5T65gEzo5iu8C35kv7eao5ah2FU8b0D6x3jT
0FDP0V4YHljMM4QosPawzw0Zsn9rclwGlPUcJnuFd+dPNfvJymbp4pC5Z4PB3xlAc8+AT4bO6iqm
wfmbYBh1k1ofM1ikqghjCKi/t9x/yjejyTQddTb31kdlzS5GEWkGF0I0T9mIN9mQg5YKrPxMwQ79
kqx6Jz+E8SKYB9PCsOC5CN6hPzFemoA14S9kkLZOQGbzeJo5vG95N1xArdielPLnTVpzDJWTKSSb
m1BY/cg/u/1ezclFoiwFoEk2XL3uF0xE/dN5CHzfmYq8O0kQ5n8fTXhBPsbcHH0qrLExlMdk5xBW
9HuaLtFTVNFzTcom5mqzUo6Q/kxx3MOugPwuk8TLYulN72vmMpeYLk9r1FR/aB6AVQbLm4maVstB
BW5AZJOlGNJs9FmljnXyCnT18SjPwozqAPZONbhhchvIiN5TVfH/x67+/LXGVV0VD3VJ9+pJCZMl
2eIajryf7NwbAI0Dh0r5WEk6ZH/W+qTRUMEDZViM0UmSv0VnP7CGQ8d1Kdh1+9edo5FN70nfGtXN
g1TjdCk5T2OMuQ2XBZXoCI7X08mWY3qpb5OaR6SW75J1w0iEwswouURJaYWfiIu220kI92ZNcdUg
OqXz9yZlUIfkdW6EpgwEv4DwRdH661oOwt4Qj+klr4+FJPjI+Vqh50nT0F9gpa1x4sRjCeWjGnOT
/W7aXS0lob1PrpFm3+0gwpfmD4bBAw6Ap7u5gYh8USK2sH9bGLRo51zfkPW+xLHzm/Eiw/iS7/Vv
QHLOMuHT8bi8bSG93q1MOt0oRK3kqM4HCDe544s/HIzxJ8ogmx7HL2Nkz4cELZf7dQHPfcgf1pST
huqIvp1HdNs+zViVmO2KJkrfTGGy+lUygUjd1XswCTTl38tv/4DjfBYEgm9DL4QmBSAHDtRUOBmr
snGvzJc4LJZU7j+/wsamRK0kbRAwM+G087UGSdlCR5/JJaXuu+NUASV0ngpdSNUrQRGNz88NdC9P
hdE/RGHCRz/weqAWD234GbpZKGn0Z71SXfaJKOOUNOvkls5dPzCtP+Dg9Mq9joIKRrRfHXxnqfOF
jSnLzcjw+fWEyTRX8cnnkOS7Y7/EYcBthlI0kgktf5Xw8+1f/V3ELUUCC+UXbWA/5ekeHVkQCq/0
QwLpQyE/CYnLMb5JIwa7KJ9zkJxcHqTo7Xj3sjRQl/FGj1IttmRfCepv+toGeSArrpCF4glOMXpR
kTFfGK1cXTCjIzSz0/vbLNsjSSeYzG5dFsHT5Ih4t0dxTUFGyurGdJqarm3dEg/X17K8Ms1Uhv9q
kGfmRPlT9/F6sBoBTflvJSS64uetOBZF++kWnsa0ub11hOtQ09FOyObCml48Tkw9yEFqFqgbhQCw
ccod2W2XH8Ih5AE9EqOdpYZ6S9JbqjO2pqnELtJ7QyQ1N5o2aLD9VGweLveCPvFbh0Cdm3cP7znh
OUwJnSptjhjB+cJeDhcXRQnRrOiJWQ36O8Hm/Rtfci2XPwFypma/H1Q3cKOStbq5AErj2FDxDyo+
JlJx+jJIZwZDdgE/HajX4LbFGSRzotiL8ZShmBdjAYuEP7dtyEHy95M5oOiQuvZFZcNOaypEPJdM
QUhXkWTDJbt02y/vlJ/ssMJBEvatAbeszdTg0eS7a75yTDALZfs7hXXSTrgzZCE2LAuCQOa94DfC
oUMinb1CIPG8ubH336+0rfX0t4xh1t51abU2GklaWLNsvdghVc5D230lKTnXG618os5AjxO1GWE+
7L5g18zIGLE1VPtMeozuHmLAvOUOcipEOi0+NI+83cvlAejNhv3gW0X8Ycs/sc9ia6H8uBp0XxBv
fgisfQGBQVvytDxWx8X28bX/R9B52Z5izuZzOdp94v95YnY5FRqd11RushJIUXAyU+Sm43v8bM5U
Hr7YsTTMP+bqZJz540yLCBr3Gvp+xBMgw/4o0GsTHoQR48MH8GdlL28xokPigjl6iggBxEs4eJAY
fuPHR1TnAhLh7BovLxBqS+eLxwr0hcY5hxCmz3x8anV23D0ET1glNB9hL4sEGs/opj7sktxg/Eur
FFwNHxxGaFtyYj0WziDLALm+3qy9V3nIJO+7DMhojXtAa+gaXzahW2k/6NO83FOE79Fs+fvJDoKn
/5JEbXvRhwgQ/PklODgL6HajkTmMXSGeMkjpLVS8udpH7jm+3DDyROAgqYLaluvAj6QdQprsiJtI
E3Jkk9RonQUKO5mMfkvy2yVnuyZ9GvEOjF7P293GyChGWPiyOm4f/rwZqQpt+rrcBUevXhRQDitf
hA9aDciLcEGM7mu4KFBqfC5qiqqQhrKbIispBC6+I/mQrE/Tc1q3V96csCtpo8+iegMfSVFWUvhV
kdfrr3hJ6wObJDkcJbhHkVa57vuDqvS3VmQsO6xAgFMn2HxEv/ZeC8nmF8h0t2n4isvJ3KEiiFxU
XRtJwbRySZAlcWN2vtGmqzQIY8oXJV47E2I0mLIqtfg1oTuRUwGuLcOHwXT+5Iuypty8+mg2jjqw
oFnWtBMjYR52r7Mef0eWM5i5CFzNgOckUpx3hypy5YYlwUXe6XHttklJ5zXCXkLBRq+08DuBGaXG
UvPJm6HnoE5bZNeIQbJ9HZUpYc6rUm/YJ/ApCXrjEHZt0yrdL703Kak9YwHXx0VJoeRmWoZJkjgL
3DRS8pHbqwVFuNHKecY1a6JFKc+k7wlq+IyeKWpG5M7iijx/j8GEAIvqPX67s5nnhYnr2VtRdl1g
VuRbE0Tg2cOvs+sU/QjGPAC3e09UBcPeiM079ZT4YZiOmXhu06laInsS6iaP+5XdEN2xHa5NMnSt
d0OrdfqGLo18piMCoyDm9EX2j5D5kUeh1LCvKmnsSMz3P9AWQAowirG6Yayo89dFqrDPn8FvWJfr
kP/GcyntDxr7nQrHygDjM8dGPCCTaq8NhhLn1L+xbqqJO/A4oFa6l3ZE+75/NakhXAsJPmflaY/D
ejPSiH7/MChKr8Xs9zELEE5a76vghvLTkPcKiMtagRiMjoDTGFkh7tgXj4Cttt9qK1pXpsu0b7t4
5hGk5OzH2Kr5kpd87AMJc6zeUtTReXp5sY/+euWaGDWh3cxRu5vxFyhRAWhEDz6Zuv5lNBFOeJdr
ma9nwJ+sP7echkX4BZfx2rRRNFWvgE8nxdosyd8wNAdNT+dz4tLofkvf/ClCqG+3gQiGUieCy7rA
6zqgI2z1QXxR/+9O05cIwfeZkC3whdhcI6HlQ3Pv/33cBbxTtldKcyueeK4AjxiJCqihUa3soycF
k1gdjlQdTzrWz9TfPfhZmC4Sp8O3UURQfStOi+iQ2ji1pfADQT3xJMw2AWbJ8C6R5ebOsNsgHsz3
A0Hh6V/HqXZ/0OrC39Q3n3hwilD2ge191Ubnpr9E9dUYM5QPMPz5lLhCnIjY7d3TpW/Eg1ShjbpU
A6OeATYM3N6oA1KqfElWVBy7yodySv0Gki/dhRnqbdlEq8/AA/hxYVQEMv/fEgg9+lCCjtbClkQr
QATXd7rQNfJbBo+FhsxpnN+ecd7ERu2+PGsjokltTP5HTlXiBHGZeS/Ybch5kVREFDFGPobI4NWB
wh+KQmcLFOVHQR8kIqvWULHprRg0pkXWzNdpUjT3GnXvf+C7Ux3Fdg/CgtAvSRaKdpyM7f2S+CRt
48yrAozIYzw5lmLCJCPINT+rLPONgDCU08EjUOHmzVy6VoDvnZxxivHf17bCm+IYYyo89R9Cpvzj
ij1OPB/RStNFmk73Ybstb/fWdmeSCSWWGf7uzixK3Uch7a8PzeZXSSbFO1hWcO+azDGXAHPvWgKB
yvstImG8WIzKyTz11R0Co4l8FNigncQjSInp+CLBZvhrBhwhynitp8C+1tnj9mn8fCmS8kUB3jhi
f2TeNwZIQh/xhd3r0li0QDk75h1PC1FlAsICdJLQRHVMe+lOYsh3MOn53/PAtdgCzJjpCFT6f6zR
n6hw9fHG6yH+3BIZ87Bc+Vva0s2PBldk05NF8vxpw6x6kRpG5F4HMPciksnnpyspq+fyhJv3jiNV
Tb888rTDCOec6+Dt3d/F2RHL2KSnVr2KqgZ0qEDF7HhupfQUi3j4tUTHG1RnFo8oUaE5vNQoWcTt
W1T0bAHzblImzwf6xVQOzOVnxkNVl49xvF8tMJOfyb+CTkNUzbTiN/Av8B0U69J6zZ4/AOtPmR1v
1fkDBukA/RyYW0EHWwVXSEtYdf9Rp4ThE/Qx3A284t7F0FsFTliJD9GDxF1aVtB25Ap/U6lcHKh/
JmznKFuZTw9CqxyD/5MoCWAcuSlMM2+HuOtPD7I8fRAzOTd443ytSwavfwxHYjTXd4ng6Q1S3aIH
6nf0y7CqUytSBr5mNLWvlVMB3Z41l/rz6ciJpxVmXnvjxr9XDJBFHYSc1WbjbsZMBqcL5rNkPzF3
N2bEGhIoteIdZW1z/A90GcVub1RNzfaqUsn6v5Y3ZH0Ka3W8HK4g33ddz7qCF5+Fdpcnbhi6O9Go
ut70MumuP1Qi8FjK4ELTrY7FloemSVt//0Asa5yW8TOp6S0jPGCL6YRi1bsRVnmIeW1+4S7XO2zK
Nwpfui9rbBHEzRcSShLgZzUv4bTg/Hx+eZl3yzqFJp8rUZff9fDFI7veusRFbBPPH2WOtmcH
`protect end_protected
