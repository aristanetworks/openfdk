--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
SQsO7iyp71OQvdoA6VCPjvVG0/Qr3d48EGSbANKIck9dbCzxJGAqK/CrRrZQEkpDCa5j3g2qrXFm
6bXkbY+UwIw+h2wuAxXoHvKDbWy22ZVNeWavuxR+avQGMCnTp9YpuR7v9XkNOcGSGN1JrRxGEsaB
bXy4Nm+T6RUlx4xnTtXtSH8uaoyg0DkLTYmlvGEjWPx4B3mumC6gx8vGI7Hin21bZi7uWv2UxGZE
pLWqrUPpIFN+nfKTIaTvhwn2AE+zj+0kYBy3YgO3TwHqU7hu2vVTAniEAqe3bq+2VdYePxZUJALy
0iyp8AuwX49q0BWl7I22I6EBji2hJ4rQomILYA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="P+Fy6c6HxkpTRy5OabcfhLgDTWKc0w7b+aIBALzCeBI="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
Q/U8mukMZjQksTxXORqXM/N/LjfPry1NB5K0DVAj3b6KzxPgniE4N/YEyYzjWA5rBuG6iNXCr9NO
UkaFSVP7Y2vEcW97CGSfRddXOG4Y+BguFPaK91QyB0H5xO74sBQJx7TZJW8SspndV5Mc13d01bEb
J3zbddy7rHWEbt5IukhGRc7m1QiKyG6PaKgLoVmPKOpwffSQwTl1+81pPGVEGn5OaRZEKjjh+0q3
EVdjtkbtcepIHwx0HcDkpacBVTPPokdYUECO/8ZTUu7VXxMHqjdLyIBo/NInIGAuGpHARUMNYWKn
kiNA1EHRTDOQi3xAtokNu048HE3OUBF+geRRAg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="vtI/gn0H+oigcRIvu8R/XQa94pfKP78zw1sOPdpWN88="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8688)
`protect data_block
8zeV19TkzankjwfGfzGPnBDUIrEu3lXnvliHzAeWASfBcVEiJWaa6cUNu26LffzPlv95xK7k0or3
urOJfIPF35ZUs6EpfK6lEji8a6pPXdXC4lmk9DBoiTEYEA8N+AzJ+PZAAR9Jm64EAzVQuPmpUbTv
WwMwcz5geULOlszK5DAm91Em90de8Ber1BQLhdtybf6uIGya/E6F+bCDP69uniVQ248wKih65myR
bJWoMSNGwlj55br25ffVwIESJ77EeK+M/nGq0P/utC4DaSmfELbEVfov9BzHOaDEFqPZWDmZpEFf
mYnc63WuwF0YV9NVif76TKZGhWShbBLaGZzK33geTPpxtQUp54k67yhix7+pRYV1TSShoHFQgyGB
K78akE5I7wC2ZhregVlooH4/N0Dw2ZEctD2/8iJOhecTHPDUPAb0PEAn0nM5wFKGPgGvErA5D443
mVh4msP8rqcIPaapqCZ1D134vs4IKHGDeJrHx7BMMnApHRHJZntoW78O+RQLbxT2/iC1Vaiu/Xc1
PDiblq1SxPiGvekKPj0mBCrw6CaiuZ1zaqH29qPdgdSlxGzN9uJZaDakfyViwQg7Ksg2e5bb3TvU
nSwhcDWaFUtHL+JLXzgsFdQf+FqvLoFHu43ILP338xqlipdFKbCaIxPsYp28E9xNqeJ6ODfWkGqB
j0vTC0p762NP3S2wQE8FMByWYCKr/qn59IKP8DFzODDKQizECOobg+DE2FtfsMIhH2329yQgsCfN
pdxtAw0gTDUK/71npRVNT6Nzaj/S2ApdOEs0xFhoNhXA4XJRtzWKxTQNLjlgpSloLKr7sE2ZDldt
EEz9PNlR94ZV0G3uav5Eak9IYZ0V/SbzjFuZds41tKaVxvktwFE7whSom6O1uZsMSKmVszah4Gs+
vHE5cw9WykjQXjwJQh9D3PHvSdJ08mawXcQPdnKV+Om65fDK3Nt41GZlEDfxq/nghSFAcdFXtgGs
4dgPLkRpFJX7wo3y1zF54EIGwiwmaa4hQcFBtgqNsSrSMz52zOXAv+Cx8MIY/FHdLghSP0M3QIo9
dBfdFtNK3jsrRX0ztKW0+jTZibOBIAh9OtyS5PwWT0lXhfer9LU2WN9BY6+/r5OpNr45kNqAHzRB
c+ljSxqZqBswTwmf1neN7tZThCgO7pfo2OjUf5q4kks14BaINYDrj4uFs1tK296VQYK5m2y6CDw2
n8d6PFkpjZT/wQvcQYlwkum1w1tSEsKOQRmm05EO4XWyiUsopAhhv+yM8isrXrJMpCfcR1v1VrsK
18eaNLMh00iRpaTOuM3Zs5y1hMppsJMOeE8WZt2nLdngx//6RGo6HtP1Dhhw789g67qCzyOHeRXW
W+rOH6dth7i/oEGm6xVcUjkOZi21lkR9pRnYGj7rgTqJViYqUEjG8MSjZtWrYJA4uJBNi46z7o5w
dirPVz67pXotoSZyIFo+EUPHPm/mGoTBuozhdykM70D6uUsOID29EkMqHywGyAn0tgOwChVM3m36
4dACdGvN1ZomrFX99xIFg0SICNiE2vGmNPbEkQ/Br+rzB10AViG6lZnp1yyntf+z1j1HCBawtbic
BJ3Ko2a7ULNFwRdzhEujMySxFnqOPuivZ++tBcC0uioHHcoQ90fQ4GPzu45Pd4TUQ7LB65f8PAVK
7obv1ykxwWTxWL4DMjCNLXkd/STSAMy1a5g0hqrK2FD0yYjFmMIP4X/sQsNaocWBrSRkvVFQwwjq
d7ms/6QhbrY9QzpGca0n03Nk9AHMq8B7iAty0vF5AKGDlAlzwfiMeslhY0+qxcQKSpCRThAEuwmP
YTJ2M+T5DSwaa98VjxyWf+ymRVe+Xv0Hu59UHBqAg7Z/rcC0gPL3ImJ8fb4doO6nqVpRF4rbcXCd
wYO+vk4z8X7Oyl2vB9qNZq1fSu/C1uRdM4mzPfkC6E1mnlKELT2Wbm+EyadfCvTUufekdbSg80sB
JQpofgNlfAatRpPOBCuLFB+xQTgncxbGb+fUQtaLK2bF+P+q6Bq0sDtaoKbDS/+CUJJWLKQ5ONF3
RMJ1/vG66RRpImD5NpyPhiCgYHaD6i4WIa957kR+mF1HAn7Rg2wurPZxL6ON1bApLD71geAjo6BI
l5xQMyEXJF2tOigvAuf3xu8GR9FFV4jWNsrG6x9PRJPfSTDb5GYwCRzVXRsRKSWVroP8SsKmtnE1
Cfalx9Rrqplh3XP8l1b4Ps0Yf7KOJ/n5LLXMh/38QSqfFZRT/LPF+3EqvpMoOX7bMydepsnEO9XC
XBGxW+Vp7V1c+L9YPOV0HYa6r9ZgX6CCvS8WeEpYD8BIFz86c9D8d8ZosniRd2J6pjHISa7x0I+r
wphLY7FURzLk9J2FLlO+VVEicRL+pDTidpq43qRL3sU5RZe2ZUGs2qTO4JZnodCq5SrtCEOdrmFh
S9bA9SohjTLl8l2hsYlLjp0KZGWB6loLPtPnpafMa6ne/pYfxh6hGkvN4Bi1Yesdq49h0TmSmG5j
hkXtfQm9suoZKmzQdzvLpFgUHLss3RLG/oFKddOJie5dMLkRuyI5LczphV7kqpvK7/+rbNZ4htsU
UBwYf2s40W9DxmJ/ER3HJeQpgVcARY/UiKX88Z/ip5TnpO22L2YhnwzIQFxQy+zwvH1xyYNnJjT9
NwDkt24E0ePSy82izthS2ivwBqT93+0FhL2H4A/ZHcg3FyN6jJXVLXlEMAuWxX5CRy8YYUtlAzgm
Eo4pB6bDRLWHYUONQIDEIQzbZ67K9vUlNoA1RkUT/Q5s7Fmancu9gTt89ZvW+WyVzXZaw2JX+Hvi
Iw/EHl0Mq2oYWYteP2njJ9hyu3DbNOOL42WUR3kWCkoZOMch1THSWayZuuaDyg0EqiNhNxC3YXAn
B4tDA8d15iCYtiQb+Qn+9ZwS+XhcTXT5CmGNaIySKafxxbKXWeQwLa9eFakDkSco8tZIaGlUTFhY
tGC/LVQ/a91aGkPU9fz+6CH7VYIZj0Eg1TVUbBSOwhg6Bimo0dEz+iHCv85A7aB5js792GwOx2lV
U7W7cXLxxAb904PjcQhzPEMtRPTQDPUFg0USjnMw5try3bEJeAv6y6fHYmZrTyGWuDkxnQFLkuVP
13tCaAyh3vWSCCaxvSYYvaA1qhwh57axMjUMqQhUS4MQiRyoDVCE5Ma13WFNB+JUjdlWNDSOzKzN
9OwjTUGcOP+yADnBgbJtF+IJRGBnXkZIOdhSh7F9UqksTfhzPZhBCU1vLUBqg3g8P9XW3EIwF8Je
6oExrnssOjh0QKXhZrqkpoiIA/HNRnFfwXhOMxzADX+UYRw54ZQ/rHpf2l/GttgFRUgDKuo5Shcb
0NVu1zaa3ed/mHgSwaZmn9UbdNWe0ZHqj1sX6K3CXawx+aTyO3yASB2Hdo/pbCtRtTpWYedlNaWx
CBNHULXLJRAYXu28lqmgXR/an8yD2PcANM072EIpJKt2J8CJkNOFpDUcfSoo3QdO1U3JE+ECk71a
dwX8s/Q+75AuyLwJ0D2loARDR71cwWV9sz2OHMaU3M20btktTOlM28yqugl0gLg89HtGAHoFk2v+
D/C3ov9QkG0WiCrHL9obPAgRO9OYfvHy+DO1J9ZxBM9mX320YaS3S4+lgR1PfaLHoPCwqbyMYKjM
XKjoBucKlX3M75937WbHfXM417fch0wXDvtWqso4XwFI4XUO41Ry1A0OsQVmOXjqjHvXOtn1bdpe
8x8q7de003OyI/DizdGxt/TibJbtPsp+/51Imroxt5tyBnsiQWd+RWNN1/ttOHsH0Sspzu744B2g
1kcUUbLKUnOgTGob7fvGipcFk4N1aiKVB48JRl6f1T28uwEMQXFEY65VVqPdV5FLqF7Ero4CYGHh
rHBJ+m8Oy9ZpXJAT9NZerSp1l4JZnIADmbnxjYpTMik+PY9Xks/3JrsFE5hltlX6edMwuAa2hChs
qEyQMIhEItItomh2jIb6gBW0OhL0E6S/PtdDTUE+qHqhLK4i7D0tne7+xOS/+n76rtiiourgCIoc
AE/e5KLEWWNir7QSF0dwPkfcaFs+ch/y+1oVnuyMzilCTK/qNYGiPcKJNltd6Nj3lm6uiL1MSeZL
YZi7l3uAXcMidxkxcFi9jEQdgQZdoHtQyPgfy9siGBQHluMf2R37pnNh4FPaNRkkBw+Wb6SoZ4d1
ipOVm2TWG4133LuPhYxdXaGuN7qsxjVBQsiLLigfmjQ7Gc06IbLd8Wi6NtDtHoMqQgYS1x6obIOb
nQsJG5QIwjr7FK69xFXtlVMHxKTBJ9cQPzKgJy3qGbbzP3W/Lo0KKZ9ah70O18nucym80JFOqu4Z
GgzbWzJWsekmsndsApuLX9b1hPcYJQQ7UI5oRUqKgdzzhOYP1t0QeYXIuWSTZhtIEOJM7lf1sbp2
NDCYxEtvnQMo5L6AJ6jzrJTBh9FZ3fgA9xjE8ZUAsyB+PyFLXfkdU6ZzkgZO6TLPon60dwaokRrQ
fqkfU1fUQJIpdKdKR15k/kyN0aaP9E2S32sQfac7r/pGgfZzrL054HC94xBtmjUYHxifRpYTSxDj
1Qa9xqn+/3y9jUo5QkdoD6t9l2WvKDJud/MpulG6u54U56YEoknwK88Vc5tz5f06e4jLkkTynOP7
2ULF8BYlML5fZp1WV4ERvv8b8LRfFTZowrFdg8Ja8D/Y3ldegrnv4QebzvcOhPvzS0Rb1dioDeuJ
b7A+RgGQ5uqq1Y0pC3lZmfPOMrx8tlHOSJ3TmdMkQqLtn4KL9crySW6SFU8rThxE9RaJ5aWKwo9b
90WlfJpYv5cfLRd1qKSlpYWp4r3JQii74IJY2dtO0zmR2jQeHVDWLItKN1wAV7sMFgiLv4jS+Wh5
GWvNuVSP0Dio8iHrDsw5CcNVOmZMMSYC8NWf1mkQG+lkOTtqC348mPMjAHqTfMGNMKHcrlJRpo4i
gXSvLiymSRDhn+mzrn1w6BycnGw5W3asbxw7GFcFbXTjTTSYgp3wesTp8kp1eqGS67crEPjb8b4R
atIbZJnDnTCm5rfS1GJFwZYULQEDRTEiFzj243afZfc+IIsAvsUwG0aySPW9h+mRWaBWGaQ/n1mp
Pu5oNEv/W5p/i34yaoHzWGLv0bA9MdV7n0DTa8Nh4RDBDjsbSuEmRuYJ+bj9XqkpfpESjLR2SF+1
Hlz2p1gnk1yU34KnqOmYXaWj2bpjNesTNmKisd32/uAAiA+BRLaK2ApdIRvGYhUggjoyzhLIoX4X
QkioKPu4Ynr22M69/EBJOQTFEpBgy2ondq2PepXHlkMR/+75c3EYBjZIbKoXHOTAgRnP23mcUs4Z
34CdIa7nNIeXfPglpQW7ZQigZR9yVLQRiIKR55fWHz/5trVMQ2iQ2/iXSEb3WtrduxselP9QK1I4
spOtrwGe/UyWbBzpTTKb3WyGaKPGeZTK4/Hb382nMpsE9cERwVYCYCENZ94/DuzsjDqt7RpEh9dK
2MIViM8SKdjCt1/SCtJ4xwrmlY99MLru+NpOnOr34uIiWzdvvFJ5dcyhue8aZN0bY7nQTRPpeo+S
zDATTrp+/ywSEGNodGi/LRoNeUMJyPzWK8l7JXBHudntRZqoJYZ8//KxdtswB9+q//BJpb4KRGIP
GSlmSWpbEad7jUt2lsloP0ERhTqy9dtgqudwzFAf6G34JcmT3bXXRx32d7BBuF0h03rq9BdmppoL
qQAeb0IsZYhKEmv691ov2QI+/HfsFAThoqdUikAL8Q7EhxZcRu4wOgt75WL+owJoyitqQM6Hi1Fr
k2H9yRRHaAHteJYMfWgozZqJUIqaPIB2E2+Ux2tu/8oyfWAvoZRDwXeh66FEvNnvJ9G1DrOEPnXF
8va8Uxi5hKodEeByzYHuaTGrLQG4p2UeCWzsEq9IhGAgKYnt1C3Y6lK9SjlfVq6NuTUE+4r/TACD
UFWf3hLRa1V3F7BPm5Z+c6EiLAG6mK7ieVceImqEtiK8NkjD2pckqb+5A8gc6jegPaDrWukWQsbA
jCUEmXcyJMGvvD3Lg5lmiMMSq9Zxj7WVEs6rQoHxXVygnmnkwPFoVnJgc2N8l+FO4Dh2vp7SSW8b
e8RbOOh/7T8z8PFyFzJwV9zTzXUiK1nTGi9GkAjtjGk9OUOgAWGGko4ZceSsmhppkWpFcsEXYQPe
GfTvSAW7QFbMeazJtQxDJQtY5L3OM3eay5Jk9585eFs7c5PypY910PGPHRq4IuWMpgR936D5l4ug
lwCgw7SPhKrgQx1Zmu4DTmvgMgliMFFOLPRo7edpLGFIKnMpf5/jKjfmD3xK1sJJHx7N8DebLNuf
oS8OIDPAPLKuGCi9Wym6BN6MsnNnxQ1+2+f8qbDEos2WGGMrQUC7HlfDqiCF6dMCf9eN0q10TT0b
iqDWiqatywEoGzoFZ626ROPJTvokprwYMJVBx6pabbcg8k2lMKa3V37HS9matZfpTHh7rjzz4Sm6
MaKPTHzPtsIxwPnkNBdgahCkB3j/P6QHNPP7SJZLDJQ76Dlcitwb+k+xUoqyeUhkymIlA0ThhC5l
ghdQi4zbUP2FjTEptz0Gdhcnd4/aF8owhtSh8JTtSTaqpKejEGv0fwaPXWTM2ESaPmdehpk/VECC
/YFPXQ+6JvwfRJs6kpoE384YGqvxKVuuMLjFxQg8KOqMLI4cxx2NeKTDDH90RHVfcXFaBPy/bdqU
z62alGokkzjWZnZiN5W8RQLbOE+csM14XRFn+5qy5qOpLK/0gd7646OjA2GPXNbVCWuyDgZvhI5K
d7eFVUQkwCTLEdgwbgp7SWRMHyEOToysP2TW30r7c3TTgSNlTXs8a99Y0pJfPBxJytUP6ikEu4qZ
LdmIlOsIXPLKo/TPYNkF9nwMJ+UM8CuOIOi6OLbmf1LeB9LKXa1yldNfU4pT/ljklYLl8oRt0+BZ
W/qJheoJfG9JwdmAVTC3UADiWrmC74Jgmr2IrdP07KmM+uNoibyXhpCJ1gPkt/x0YoqH0VyEvwgc
j/1c79lsKmg623bjojGpJYSvj5uQGHn7xf7cmtQz+eQSTDrpJajTIImHCWP4/jo7SJ7z42n/aMIR
yGvhvbeFSByLiv9wkrvWCoyx2/1DxRrRZGbKOHo1OMc2JrEBU4JFl+7CsoiC+xewSAzbsUGefuXQ
PzlpDGw0uX7Qj2jgaIMgedkGpAvcDm0LnVctdqYgC/6mDdkoPzSE2SArREzszl8mItxqrmg9jD04
c7t1L2M+DZZXy8A8OGBibJIV49UvAbX7ZQ5DcdKvUIc1sSqudndNsoQlm/wHt2z9fm0i5bprNYf+
iL4dXj/YrScLLXzTHa2ih5tDCOAwQ+bdRhOQpav2Rd/zcTAaCNTAvJ57YFEvkFTIX7fNJAwmTKhi
i2cQuJJnV7iR9DFVu9FLnvCM0CsQ5wuDS7Qv5h25jauEEjvgeEuis1umLcewD+ia6QbRXxnjhUv2
jiBfGbTkzoBF9eMChxcGLvUoyxCwNJxnf+pCRJvzx9fVJb8EQaiNJ1ZtJtfYwBn6wL5GIM+B8nVE
izJBOZMGeUKt4087CCUxat/xBKFCSe7VcU6r7MVDn0UgyiE1lLLTkmtahTyxQSqnu8xs3Uob9FRM
7TDaXFZ2IDe3o4qMa35mA6wNTB92p8aBNUDaWRT2lMrbLWc0fIEy5D+lcHR69pgapbjRUTrXO/w1
QmfYzUqHcWaFdpQ9UKHqYa8EoKDvKAmx90Jqmi25Q/hR0VSXxccWT7lzZ8XJV0qaWFT6IbKjDVY3
PGHvxrLwesdgbjD5S/gx6oLE73cYwY+UOiEN5T8c8V8UNlIm2SPa4CP0uC6guGDKorYs2ZF3EgvN
dnE/AIV8yOG1wPgLIwzORMYWpjGBBjeyHK8wpWm//zSCGjEvpy2ygsu3f3ZFEvl9j0RWWdKZYT1A
vvBNIc47Oi0o5XqB5751lH4XasvU8xrhUJlkdiOsHxyR8m//AoQS3+S0UeAEi9DC3aX8is1ycvV0
G254Vhiwv/JchDlDLuWb+f2D7/1GT+stK0Z8vsfMiqXL8f822YIuCdRce+wFjvJZ6vOe44j8Lw4K
rf2ZNBrNt7gYrf/wXXNrHgIev4hJctXPJxG8pxQvv8mm+M/2J13/7EV9aXUjeqIEPLym0oh72PX8
wKcmv0UDOFFF3c6wEwc2mBKeyoQr8yUCwSlaMked3iY2vsuSKmqDKOH1UFwG/UOHcOwUY1xiSHIi
C7uVaNVW7PLy7moxq3WtO4uKKeNLFD9zG8/dqzE5qvCLiUC69sJd+k1mOwqbhpBXjsqI8haqNbKf
I70J47eWLtaqHas2+jJQP8sYeF9f3dPSjg2k0n4+fhx60Gfef7R8qAAGot58KR477tXD7KdUBSYO
HBazYlwqtRu0ZKCJ4oGIEUsgG/0Fvwymn9yQZUfyLByQ96Dwqo3O02Lz+YKbIkI4NFhjiYqFcu5M
vd1bS4t4nxgw0AxIXUEscfUXnmQkQrj4wnoAS7rWggpa2UoJzfoE8inswPP7GS391TaqqRsAYLF8
GWVSNeCn3jUeFWIXrMQplEZHYZc94Xd7sKSrTLVYel0YEf3vZ8aftMj/sKV5FyVVsB6RObOe9Tt6
NCyprnNIBnTnFL2+xxYf0AORYf8CZUCb7gB+Z32fHorIYupEiDQUTDkEQrtUPtMme/2gL8ed7Urt
x7VXAav9AHOeegMp4DCtiXdORMo3kplR5TKKO3tphNWhoXNvm6hsJrH4v9x+mqrNjNAC4lMKymXA
s40DYcNArOSyHC2BMcEbdlWzhpJI3W4zmC4TLhLKPEW9ro1pSAHx0l/lI8mROxwaZ/IiEWAuo2fC
pc9mF4SIWnt5NTod7jvOzfpblVZRUtSU/I2aeFRmmbHtTnGu2nGgfmQX5ehuIrJOi3lLMPhXrGB6
hAqFMJd56/aWeA14Ovi37ijb3l0Qx3xzfS2gaFeuww5GeDSKafU41cOJssCW/Xz+nM+MItdSZdSl
7X7jGdVbA/X8AzJrPlMay28e/nGt5V18OVHdPU3qJ1Y1feaOT9EouQHUKmiukTpGKbUkjtQYdIzs
npa+C/2R7KGq6aF2r6LM3R5BReGx3GujslNWR5cW8t7CIklf7u5k+mKc7cT4fXRsDVh9vjyEbntD
DVn22upm0e4+p2Lo1Rb75M82i00tRz8BYGo2gbI6huntrqi9tFPOhKq9N9pxALleuBOX9Pi+gnzI
Waunp9fIgZ4ucS6u695vpVWiF61CUpOlbu39Q/MIPz+e3KNbjmJwNEHcmpVtsZtnpgcY+DU4EIEV
qntLSzGwPRovAxsYKasLW6zF/0AXQxWrRIlYWOw9ZZs1CsrDprlSxRt9n5ehf6q5JyDWdfJF7g2K
hp3mCOiPD9ayOoC5RYULgx6xTSGJlcG1w3B1YE/qHl+55Bf2Cf3QqG33S6k1Vp/ji9rzma5QHT4a
gUIq0JHLh8l09l246VTyVQP9SCBAX7Jd4R3xFd4n+CSXrsN1knNuQzs7wsZsvcmlDMQ27GnIpKSP
stsMT5BNBhqI0QK/422TOCRVLlNcdlz1tjPf1u1ZLM8S8D7EjCEWN8q/AdmOpj4RujFuX0KZZJyP
oLTadpOXM2sVIO5b3LqC8hIpboTtFcwXGTzFbq5zxMO1wfl0Ptfin93JaRneFEfbP8aSkSEilFrK
mQ0EoHHVZ322h62OMV06Yyf4lWXegntBNXYa2ahydCQKsePHUyLZMJfyKbhyKqaxCGEhRzn7Uoaf
tJrnaPOzhGyYz739zXr33DgCmWy8vIq9ziQC3uFnEw8fsggZVGU/KsWIldK0cZpIjKBqG3Ug+08K
4nYps4ZG0d3ogEBgqVV/f02YEPdmfOAYbdkBcOnoJQJUhYakIuXCGRPQcx7Gjk2tTX5aWAcM4tIn
X/5POwQF3S9JujNmIDBxL6I/VWh+SnUpuAuovoR+XJy04Rr7BnnQdBxy5DZne1dYRUNcEjpKFW0A
REahe25G83NE4a6pK6BLdCSUO74ELdw1QarkEuxUUZRSCKHOvea0+Q/mKDuPBMzE41Xun2YHdu2k
l/OxFLkfu/csxksjEJR6ydinzQ5huBxDGUMWLO2rPG0vgKnty3vQF7C5jHYkZZHjErWJ/L7227tT
dhrLgz17hRq4wBf3nurDnvcbylbtmFAl9uwPumF008cRvu3mxdGyRnw1n2OHDMNQQyz/wGhPvleL
9R2X5VNjT9/45H8Yq8Px+NnV8YMNu1guS2fxZ9LXspCWYa6ZvDQwO3R05ua+4Enn56htRw+d5PkD
TnpnlT5dNXkNbO3tSDvvt434APHsvZQ0U7f1/1zeSaevMkWJckBxl1/+J2hIzDckUVYIEwdJ0zKK
J4Qz235erdtRD9iZPhuOE2UkiuALf1b3aa2ejUMQNJ4CQtjYklagPKFd+cQWfRTgvRQG/Cc7cQMp
CMcUGXvZh+pO/VLoejMOsZVWky7H3Mtpsfsa9Vne4NzcALE8z6MytJxpB3wFYEZzQK5+eWtGaPfI
5808xYELMErMEYsVU234tOFmNZT+H5JCXWqsWzaYCLh9wJbpL5d1z/YfGHSV8vuIXO6XbAmoZ4G3
MFlaNoAmoCgMdu/Ed6+nVJZC4pQRN6PZmRpmhednJjTAT4y9OzR7ujGZopQit5uGS6A0CNe/YdwF
vj5vEcN+a/hdAcTH7W6wygp+f2R8Kn34LxEJiJpD03wzzCsZLC+8hPUqCyWNRiIwUqABd+tm5lx/
wWR05UhBdQEX2t+6blnTdzCAk/LCpZjJgiFqSpzJQYC8jdMOOdcEAlhp+u0pKucj6GStieV4GEwQ
8jX5FPTfGnDAWRq/MCAtbEFugiDFlfHAjmq7wdU7tS+hhhn9GJ04o5kIggurRoUl9xNaVf5aCEXg
cI00u2CJAPOs/6Y2/vft065mjz2lP3rH9ivyo4Ke5zoZqZJSS75/qi5KyOiaI+2AwcLxjr4X/GTu
DeFtNnTsjbb8X1xpc9PH/38w5GffLyXN6rzQQhmnaGR6lRvGMrBm/cyRK0+caXIPDmR1sCnPbu58
XSHabs0oTEf14HzNVMfWTAM6vEGE6/9r+dfewENMtMG4gBxM0y/5Ap0/qHfGqyN04ZoOzRJqP0ws
vCeUe7mOL3J/vmUSX1+9zn0Jopi+TxwghLxcJ0yg6fcjku63BxFK0Qs3r0Og49KDNxCnNSlJmT33
dqDaDOgLfuO+Yn3Nt7gXrRBcDL/dh94yKIEeQqxhghXmlcatUyZOUhfARoielqIRVHdFz61lneSD
b+vVI5JUtHzEtvvkhVCBBEcajJUC8gzc+S+CbWhDwyoGYO1s9Hux6zDPgG69UvtFEMh0rvzAN3md
0HtZCrePmLqH+NdDEEVxCdZEAT6Mb636ZU7lzSHMg8au8uQYdiwgolobwW5mM8M0SCfUZI5u+j+c
2k/RNLpSe/nFMWaHTsQiCgOb2octPloHsmMHK36OgI9hOA0Cr9CvIuEonEg6bwmnjfyNuRLmD9S3
HaUkWmSp0oIKuq1Tr8wACm9J/Trao7AV0yDfgaPe4FTopoykF/rfJREDTiwZG+vugKXXyD0kbF4J
xItfKf5fIRBV8IXRIN6QeoW28hoVvacT
`protect end_protected
