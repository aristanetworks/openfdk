--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
CL0J2uHmeylQjZpWtWkR13wiFUIWvAAy0mDIZIua3MD7oaEDhtGHkt0PaThXDdqdXrHI9hfJNgem
c1bq4lel1aHeqtG196sZ36L1M2oo4cps0fv3h8zgRUbq9yqkQctjoZ8LPygujwELa8CxZa+8sJ6W
4YnunltQoWAuXXK3Fs/6bJcQkOPTKgeYH0Wp34o4fZ9C7zvQRV3C79LP1+zDvRWMESF3z8X1Fjtv
i6h7J+pq60QXKldsI1pTJDlnO+/xg/psS7aMsNk1x5PHCswjafbU8LCmvRwt0kxSQ/gCyx1i8SO6
KVd0zxM63qRnEsm2NkpLRDWzonysQ4dOXLc5Og==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="BquzYUWHJI9bvhYoPYZjOsM2E5zVnpf3MtJyTAfukDs="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
n0885VpedqF0rcZ/Vt6uM9HqCNbqYfxcnFQfOC4a7Zqodj+SydWSy/7ssFTAbzQyAw8YoTpezyRm
X01NgP/+Q/4yTxPu/TY0pgC8iIUaXMa1XY22Qrlvw9kdkmEpmwGPiOksbBrviLcAZpYkkphP5Hg0
8Q/ILt6K90DzDMf0/GJbZQDN1cVkvWMshAjeWAmnwuynyxxvS2XvOUXvA2Q02Do0n2N5rgOYROZw
I4LGDG2uu9VV5CGVVA2h6dTH30HOxM5R7LFUK+tYvc3AVlEFGtp0mX0e9KrjrzjX28hGymUaqdar
utKoYTI6YbFWd6lv1dkgSiqeAABqAdzHF0nWiw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="REijTQ5wDWCEeHP1Y9kLOqzdB0HTcMKFek3yGE2OHxs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10912)
`protect data_block
BAvfHtDgaQAbiTL8G1RUU7kUhTIyO958toHseGxTQvOThV8oN75UZYtQe5e21V21g4Mur3qTBO4b
qZuaF068NHa3Ef448cM9gjN82Q49EjAXBlKXbUOVXi913bHCEM0OSe+MpnyDriclp0cKJqnSFPV/
ETu6W8r8D93f/fnrqtuByyDVjRbHFCKEJzJupEc3FM4iMzeXVUrnnv5m/zQMlAqS07kKDcmcMOee
5ZEZgHZbqJpfmkubrppOsbAhIglUp3bCnVhbuvwzGvfHocTuIvdWTy/rU29q6X5xV/vP+1insBs/
VPIKbdsYCMD2ntB01soacgAALA5lYOO+tgNQdnL4o+QaQaaH58g6fNMEGv7O3ak14RXaMCCd7pV9
GxydOUIM10DWCy71xLEhfpIQzMk9LoS5gSAJD7N6lCV5/b7xLarljnhTec2mDjNXhzZwkNM2boei
gr4NyU1J+zK6XzHfIiGXpJk8maYN5vhgyXQ2JudKifkVplYU1tphaH6pCvqo67Amolr8btpbTSsp
Lol03I/MjI+OVsK6cuLw55yq3aX/CF1bDBGfhiz88hyC3B58ZxfnyR/kpZCA/uCcjgApYgAoUWsl
CgOaigyZRZ4fru7mQbf7Yz6L/R27cbgWOKPN9+Z/oIwxiNUJvS7rxqmdlBAtpaJ/Qxgf+1fVulkr
JIXVi7PBGlruBKeCzbQ9as7sSHGIHlYieARihEYbzx4duTftOc/Dn9hbju5vesl3T3SIszXibeUI
JLCMKdi34eB3YbugjTi/Q6/6B4x8ocf9tWXnYjCpt7cbE/4Nsd4MCi1F/wxp//SAgCjSLjCauL5q
wAdUt3+dsaXnjxiqa3P9FuK/nQRFmCxl72JpztofcibHmGllRzDHUHfdbiJR9zEarTSIlRW5lGnh
zfY73AjkVBo0DCkDGxxY6f14VXy5D99MspHU4Mf5VJD4Ui1b6VzOM5K4WNwL7uF3v2hNsma1sD4F
wTCl/2Xc3vI0Zn9R8TOE+A/DQBcfojyqeCFHuyVOobZ+c1zUZoBisZ9J8gV9XUY2rThihap3b8ys
mXQeXLw3zizgD2JnUY4D/Z/r5U7WjkuQJZRjTZBRtj7NEjVHTBdZFkke3pkGc2tGD+F1cBATNM9h
CNPE4RQEnZ0nhM8PTvunx0h/vY80q1JAgxfZ5chGcdlmKdu7VMdli6zDLnrqiL3zbZmkqQexCMta
IT8PBJ6oIQ8vs+9HLZ313NSF3IUximzBZRWmfnBilb4aPp1T7EzRTJp4cGpn/67hgJ6ycH+I37F2
JVLJPlqZdOkXW/95CayUJ/XkkqedqDnmiO1D8DLpwCWR6Krn/qF2K9xb7zjP0Bv/V8+NU+1n53vB
UaGKgPAV8vpY1I8APEzoIrYzYoHnJTFc7S1tfldHCbVujHX8SgkUhYW7HvbeAaqQo3PycMpUli0B
EQRFRpCD6PIEJ+k0YMXH3Gmub/ULcgrAoA+s7xLPU9/ebow/p+A+wjPgdC76kqri9WzJi/+0VpjT
mLHWmCCrwU9sIle/PIIW/6BNhXd0pY6fK4fD9wGbR1046mwCc484CeM+K7DqESQ9cPpWzH+KK1xe
4hQ2BDq0VpMhZwK74V6JMHJ71epVszBoNzYd8ivdBYZ5G8PP0+rfnk5bY1yOkBq+IE4OHfWv3Bqd
7eQkCY3ZMcprNAP3g2uKv41+FmmAQbkE0+P2FUNU3NEy/xbYrNLunYKOlS0zIC0O3YVwGOXcL13m
XjDNVc4kB2kB2B2AC4t8ieNhyMuPrH8YxeoNzHWCVofpfr1HVEaI1oVgxvr/DGFg8J6G805BQ9yj
dPdIHJLRd3PDsnRxlhnSM2SA5KvV4pkIy0Bl3XY0mlNsK4AghN/hP3wTXWzQMIyyjaQy20Lb+gW9
Nw3jpS6HRiHZE7dYBlYDnFEdtUUY4ZXezKb+tTKJxovJTg1YvNr3UC1DJeoZzM4GdGqdjjZ2sUVe
zs+1Purk7mk49vuqtjRQTT5J5z4hlu+S5DQF3PsxywGM+9Bvn4kxZ8S8OqTA9BQ5updIhtWYHjQ6
wT5bFKlNdqqPo7ipYlTusPlumfdbufTWKOmukl2NQBT2CjiL7Qhjsc6cmTOSG7TYX1nGYhFM2ZbS
Vh8y1UnvfPuKXYbxvu8Y1o3APuOCwOmjrKNyPw2nreTf7ok0TxwYqag7hu6XRACZB3oISgjKEaPm
bxpvb2LQdWR3n4HO0/PqawtBBJlv5CG5rcdDmu1VNuMweUI+vpQKb8mqaDJPo0lLTQuq95cqAcqq
NcyhB28xTqgVPWI3aYtqzK3MBFs8cd1I36l1IhWpGnDheK0qJsqMLlMr0hpRjQjo1vrL0Htsichn
GOtvuIDeKBc/d0dFqsGR0aBLHYOpM+cTUSmdOyoXEgmohp93i6YAYT5w9CUVRsAcQuEMiyzuf7nN
HSNpa29F05xLzs5/LHwYlqmABi2FZeGW2mTT7ahjyMlJySQJatkzg0At4Rlxt70emAmLC+UnTTtm
FgXxBsML5pGMvxwhjBApxUczParLnJNXCXD9Ri07PZtLEOWVqbfRHZD/WfrdyDeEOjh/8O8NIQS4
wrwRnZRgz/Cp34B19IEE8ha3PcW7xqVs3BdHtr9vx1yhCE+IRMHzsHey9Qs4dI00FmhD1ZZQZcF0
u35/HuYtqhEdb8MgdA7OBWMZO7yhEFhjhV36AUMGULvh24oe5SqVNxkUDRp7AKTg2nSoPIiz33D/
Dix9Inol0I5hR/9q+RauhCPsUxTuan+Jt/Wtw3i4n974HO/pso+/jiioV8OH4hg6QbNGY8sbZwIr
VZgLWlIEYVwtBneeuYD+SM4bOhWoEnFMNK6+0q8Mew9F/UQkdOiGLeZOmQXY7LGbpHXvXC2m8xi7
dCyyIWkCKmSuH9FZDQHfWcHojfFIKNzLmmI7+Yq3afMwWyqlHfPQzoO75jieN/FwxdHQiIzPZb/V
kmCHARb1+wekRwSUGTPOUL0L0pDSS4j3hsIFQAFw5Lq7sFVcBWEpdOeq0a3AZe5dNg/dtSMW5AFW
EY3Sh1nEkPuqiQ6U2mbr+ChsxywRcRabGTu5Q40KtWt5vef2rsmDG5wXR7URConnWKPLjzBj4dJ7
+PTR2PxIMIRVE7lP/lDhnp+edvtTKru3BSnIM1JnR5flw2wJFjYVk90V1Phkapwj/Dab91dzoLBY
roRsnTDnfEid4+r+QPqv7KmKawCIBx/PUiYqqNQiq+Ue4OmLRziPutfuqw5TabppdeX3e2jbe/2F
pOtesppNvxB8G4qnkoDi0+az6IATkgCEm19hTVIc+To7VKI7L1Yf7SBUqN7TCbRXbR5/yIFVguu7
y+RcgtBeLjgNvtgK5dERUrmnoueQAXdck1b5/BbCS9++brTLftzNXnMt6cko9yBdL3EnZL9o627x
CJu+enBpBVyWr9p7q+BmohnJBvf15nxKqYvzC3eU3ujAscJoVs52bLYhYTMwoSUzOwlW35ikb7FX
1NY5ejIQGIB122EJ3TT7pxgQLoBEA/2Ev932G/mvzZKPUsrsF/F9BxNMRlLYnQ5huTM+5f5oYN+t
CuMzyOY527v1roqGlrXwFuOfox3A684ZelfGwC081f0o0hbk8alIp0QQMr3x9A2iYahkGdnjY8l0
LmwAiJ4/b2HEP4SC8oCBRCu61Bd4qhOHL4ZuYTBwwHHWmy/87KOslGIfb2dZxhebyEDEd8qbwzD/
CEaHcZ+ewwEOkw+vnlc9NsQ6DZpaqvJ3bbldGLJPBdET9z1iDT9risKBh9wHbaefh5jdo8OGJSJ1
isuEnFY6w8ImQnjlIBrFlSDBvDkA1vsA8WpIBOHDxGDEk/dtoDUEIPO6sr56gTtVzWy6/KZ5HRz2
VlM5g/Qa97Tz7n/oOgTqwPCOctdD1nBWli8z6DKy33REolk4KBuIUxSbzlF1NSzsXMFalCfcXrCl
Cfh3sllDL/wboNdqZYqvd906pw3br91Ktkg9QJl5578/QV4DgMVgMMJDpFjg9ub0biqSlCTeuLQ8
rN6jT27aUarmP+sIfzd2pmjXZ7tS+DPJ4uLLywCo+Ql+fj1aU0sP7QQ61kZvxVzuqbsQQS84Qn4s
ZxNWtoHbtjQ5pdf/JHYFXgNBphQzjkhp99SDuSPvFybTELV85V+GEk3k1oVoasRszbIMgkCfdf1z
7fbKkewRwhwNjrcbMiqJ2veRxVHI/lqrIDG+XPxW4AoT1555vbX/Q3HHCYT2qOwKGmTZjmp0A1cq
GZL0Cy/GNFynGe8vHHNrC0emG3qMhjcl4OKRWmFcZU0SI0ofGQWK+zkJbkrU/TKhHfHrRzSMlHlV
GrIUZFovXJt9JEzvOelRCLyKEGv8dnKJyujMNqrqzH6KFh4YniRFl1tGWVQ14wLDhLF/nhhlxaRl
HaAa+u0PhwVhNB0Pdx9kJDzGiUx8fAOYO9R/MLWj/Ng7qE4Z0qdJOfzCx0BFwUem809O01C3RUAI
OJRAYocIJNaZV2GFsKutj0IpiB60v2v1Xa+2jFpC8It1FX/vZXdnL5/IbMfh2LujZLGGoQ4IHjTe
9BNlMMJCr5Tsqg6iIKeh5E5KY+Da0zzq8H6voJxK0/NZJsaqhgLaUOA1KMwMKkgdeM3977veiWJd
XCzzFuWkISVGtO2F2f7KBXfjH785JBnsIDe+XGCxMLVja4LVljrp7nGgmSS5R/1/GQHlkN4Q79In
fgMd6pMpi2LEkjbthkzu89hR4oSi6xVQypPxSXwVosFoMk7sTjyqwhegba5VWnFnZs0yxZxNNtfP
reDTWBHvOT3d0/fjU3FDx6JWTOxcLLBAYhwv8bT94sk1IOP6MPRH9cR2xaJ3CH9HbyW4MxcGMSmb
8ZAeZJ3+XRQ805yfUBbKibAK4G4vwt7weNQLbqn3PLNgn9dGLuIBoykftY+An7L5319mPTt06pEO
GhH8ErXM0Qp+pvjCwRECdjV4hNVdb8OFz7ikuWqRfTRbDHdkllSxSQA7seCtJ7Z9rxQctYAvlPhU
RUPWqXdUlxvfdQZqGfm8b8D6AAoHkgVxjE+lrbFg5EKhAM1etBGg1EtaBsg4H66GSE0nxKgKvMIz
8JdPJXSNqj1AjZcJNKB7+kFHjqCROHKQh1TtpVtbGoPbtYR5cjORgWO7Gzdrd4ECGJmyKlrMhbPc
F5i/0xbSsbi6PG4CHU7eNO87CngYSmPhGxRlz0bvbWlWY4zmAi/dIepU4TLf6cTzXd1BknWhmPs9
CTPl+ozU5M0+rBXb5pCAvvbEqT0BAdBEzU7aPU7x7w3sOrnJq+a39bDhfMNp6S+0IElAvivATTxg
43WN2pDKanBZYNv7cBxfE8wKcY6Ott+uPvuiCrxUee3x2xOHNK9hVgqFaasqqyDTOZuUjOb6cVAi
THoepI/LEKDhS5/TosrTH9IXokhnrDjGkhWxVz+qD2zIRP5DZgyl/duijODhj/jWldNJ53SdEWGX
mjy/UYeJ6j1w3xVBY5x7fsyALfL0kOvI4/Lim/CXdb2s9z+faG31+lgHs8eD4dMMTMyYEO1S9dWT
ZzRTSrLT8zHEjYCVe6eZcRC/lWqCXukHHeZ3+Jgso9KVlzpoq40PRTtjCuc8GiAy75CO8056HjNP
W6ur5Qa3uKkW1ivkZOdoMTRMrOSPyj9l8gBU7J0VehXzga6aAhShvYA65xzgfxxxhk4Xuy+ff/te
aPHF3o9NXQWenEg+nQqMERIcHTvkEOaelP1kyUqYN2vYyxEPG7BPq0G7CA2xbdpDPEx+m2TEcdQi
4+9KjotFziw6bnOPIkGsw4mbjUjM9LIjb/mHO7k0Y6osfvbcZfUOqKJ59Fogp7jch9VjrFz1rKrl
azruoawVAtwm0TP5qqFVUjtoRbdJ8KJsPx9cjPzgkKVQ+t17fvWyh9llKx67cjNoPYLcqC0MdJHE
0IbI2auDZ2mxO+M3o4p7IcvXG0gankJSi3go1Fi0x/PLdg/7U2ZfpAZQh702j8aqrDnrMH0ucju7
3Qd5HRgy5en8hlIf+EG/v2PXUXi0rcXrzlBhjU1h/zgI2a/ioJhX2Y/9BpDZAcFQ2Nr21cF7Zhx5
R7QKF9hB4rKvYCBoXtmVJIPzAHW/RZlSEQ3saFa2GrayqL/5X4tnWptAQTzTHIzO4tT8y09qgTIx
e7hYJQepucJ1e/WTL5Lw8GdAf6UlJG6XrQWQ3JqiWxbkW9LeVSp04fNwfKqkxH6QIVwKBCEEARei
iL+9+wfoJNH6BhgpcddoZ2A0V9zsIVvfMyN8jBRbAfX4bqyNpKmt74O4eOPhWfLsgQg2qSRRITpl
Zo/xyR3qxhApt8UetBSiQDy5pX8de9Cl81TFIi8IkFJFfzC6HV7vQxYH3w+RQXRzsOQ+GVetJP4j
9xe/BbP44k+egNqF3NeewDQOXwb2hecb67eHPJi9g+dk48uqfwoFSaS/v4+Ip7krU/QXJ7DXxtsb
TLUji4lEH2WCQK19T/rKuAHxgvBSUNgi5acFWhDV5DeD9xVFnMTExz5TjKpy0O4dm05rz6q0SaCS
MqJzmU7g3UTRNWj9GuDJthOZiX0KrFqhk1rO1mmyEcsWe3rtbXr6hjqJ7XgMo0KR5ioBaTDmgv2s
Tx6cDor5ks1LwmqxKWIp7n72JxMjJq4xs85wVZuEITZotvQJ5nDyPKCe69lNfcPlqIQrbsNjFYON
qX9inHoObnWtXHfp8zNxRkw7KE1nB5K9oZb9VxVRNX5sm/Kj8Nd/8U34O/NQHFQQKmQovX43Jecm
wL0HwYtwqPVxaSCJJVWi59bU1oXN8FsHSuc/Jsyd4DA/7gN42L64Q4m5z6T4IndoZJCcvu5tl/76
woC7vlalZepZPKq/l7r88VctT53EE3zo7PNOO40TVqYrMUy6eudTm2v3AOElzy2va0aqqkGwWoec
FPxcCqw94WKv9ffC6RSoPHR/+gIObfF/p/Pj3Lt25/QqFNMd5VRygPxxj9X+ROpQ2hyNiGh/nBV8
mg/Pnm+T0uHzNTe1oNFAD7j922VWP4UGJPnxiqpilwueUqV5qXoTR91i+ZGGjFo+pXkvm0Vh/C3U
LBM2aHVxF7NjUMPqT5z+/wmsxQVLGrQ/x23l71RkDuJX4XQ+ACAv94WAbHWQ1YhlNdZOxhmC0dm8
yb9I6yVV2wqgMN/4EnEFPz/1wKrfnuC3r37zfaQmSlE6c7Hrqf41sGr2JaF6YBDOjSmiEr/vVINm
aFNzSIa+oWQ/PvDonKQDkOXr10NilewA40fZUWN0OBL0erpnPDgKCqU7OsMpsfCD0ezlnMvFsJKV
6f1OyvKzYJ2YyhljAyBGmEUFDAL5vviOv3Qrq6slIH4Q6C1Ap6OcCvF4uQovLLKmp/4lJIQEDB/5
SqI2+Lbv0Ty6wdtKhMas2vvd6QU+RLTSTEcoEcghiE4PJYcEMIoWkUPidCDhOiZZBrr9ZwEt67GH
5xdgtXQijp8moNNRLOzb8u3Ch/tGGeOx6xdsJdhjlDI+fAs2/avUpiwvollH4lU2BkRY4qf/7swg
NA77BW7rFZgegqhQBRXsX2myrQjUFih0QpBxkaV+birlKjfdaNwOwVQY2osv2AeIllkOT8iHFdya
fJbgg7mbx9jGbmEU5EU55uUvyAmhVwxX1874PBcygs7vG8/3sd+eezp9dxdq0S8zSd1JL1ySP7lf
pdP0ijFJ+S2PS2/rurOWkxC+CQ6SlwJzRKtoQ4LzO53j9WEDzP+dfNgyw/1J4U8ctSiFKN2f1Hyz
dDKqMEMUhjfqJ8oJLFsztrENFI5l7SsO4DIh4De3wdTR+M53Q95WCTgfmi/vKDg1wo/pOVXR2ac4
MX0bTEYDnEvc562n1Fccrf3lB26p5p18QgAD4NDZcKyXz5+xvF4GlhHNK1kVVQgckzoMcNxIaKLm
UQFEqNA0yQaVJKxT4M2ADA2d0LZWc3p6TWf9UkpAXjBrcBcHCyUuvx500VtQMIAfiuN5wnfbJgjr
7baPx5AfwE1TBHGmywEAWjdfNDNTqifTU8Y9ghd4dFOlTqMpbDK68A6ZPv0rQgYw33RiuTq3wi2D
vm5FKBfadqtMshM2cbOae3Tv2Qcla12wbFPGMS3+rP+lXPDE3wH/qA7BgMGDDa0AHlNfDXpw9VZs
TTsgG7mtTDCLLAiZR82ZYMHGwzzG/S/j8YMugSKTuLKJaWYkHcRxXmfe6vhgKMWroWaJkrjO7ZFt
ZeP2jO3vKFsM7RnV6pjVn085olqdilGnyfxHlKO48FXClLbP1l8U8HWeDooP8xRH79Sk9xp/vEhZ
vqKKCO+af/dasllW8x8kz8qcgVM6dpeP80rK530bGgfyHUkomtwcrQMCG6I6UMb1zqjjoT2jCoEx
0pGTDSMHZRbSn2uhMbcbv8EDQ0IZ6UEACSxtmdK44ue1fNKVOLsQA8o1kE99CbYmC1yxEV7r78f2
nX6YTiiLWWvI2cnEqMR5v5fV7EFAGsFGk7k5phTWe6Ue9++DnSIZ3qL67qioX8Phy0BaVuvQxbkF
+tWd+pYki5By3ir2OQenrurZB9aAKG+ihNtpJ8U3ZLdoemc0x8sKgWmlSdOmQi21VYuXKtTsZdWy
dqQhOZ748Mb6S+qUkbC/J0pPLZYYBXf1ZTnQ1HReVAr4vlmA+caea4If/F53SSSFuHFLw6bkwLOM
FNF+M86V98iwkpMS8yh0Bm1LQ6SlbV1vXFNNf1pOUawS/lwAJu0f6jeLTADJVlTQCEA1xF2x9qPo
VYzUU4E/XvvLI5dGNcnEV2ODNPM03UQyhVQP+SLTHHIiv0D+8FKLpsgWtg4ZNcoasSjKR5N/zDQO
UFh1iFJm/f75BtcWbdpQCMR/RdRT2YQDEd+Fy7Zxljku8ZH68BTqBRNFZnXUXa7aL7LML/RRHBUE
2O/hon/SnXlLD1ktgzFIAGCjck5LbOs1SGDMv4Kfv8NE7QkWV7rJEn+un5JQSqKBzqqqCUk4mVer
+np24ZsBPH1blXdZ3uMKM8qqcak5R1mTo++wc7ItcN4b+nD0rN4BEAA6Uui/PgAv19Lf+W1kuoUM
+1vsoA+R5GJSVkHODO+okNac1daOXp21ocISZ3g5JygItrXDVhz2lcEO81Tu1N8+d1986hF9Eg/W
13rArBBHL+iPZsmlS6H0uv8wc7gN6jOlcq3W8TLuGyCZjEtLzRmE/OS9uJ3EChceCcmGbHeDwWLk
denIMkx5BXES2O8MiXzPStvTgM+p+P5hQMjcuY1ubXmfphWW3lnQlovLqAfmgx7UdgTT8ncf6e36
awwZ/e1TLqv7joR4JWT0ZgxMKxShz27E9j3ei2RvHxPeLZkinOm9fAVoMl2zs/Mj0+vdX9od5noK
ahXjxL9csoOTfO2Wtq3485FAlIztqMS44PJ6vTaMyLj8GkuuWW7anJRuw4HQkY0lXWJZk1xarPaD
82pemuCVdbQu4VdPkV27T6tkQHQQGNucq3VsuiMQSJwhCQ2Ad0AELimUzow1qtvUCYOksCGVNIa3
02Zd5D+4K8jnoPmdKLmGnAOkkFo5NNJM0bBozAdXEq0JEbPT3mspfP4MBOwMW5OBrLv8x472lCMg
72gcdsx9HsTp7dxA2o4gPrPgZnAPW52NOetGtVjWaYZfdy6QaHtycsdNuzh+Ov8iy3VT8qA0GhOj
Cw2qIEG6UM3eCyMV3TDYlSZ28ciQF5Ds/24YnFMm2M14KmlDDgdJ72jh4dfjk1K5tdcNsbgqmKsy
9vR/4gAnW88JfvMmWhmTbXHlGxb8frobX9tTuqo7H2qPjPg3kcUn9qlW8KTZ2yTmYyP+Is6SbRiw
jM97uZv8CG6vZ2YNYswfaHkzae4SiX7OgH3z6NrX1FmUemoqdt9qzughjEXa+2Of3BQOCP+qSyoM
QfJcxKDXU17aCBMLqw9ArPjr87IxArHmHuQzCurAhmMOqLrXLT9UQcA+dyEKGeKMmpMGQfoa4gTC
02VX1C/6w/dUJMc6WuE9vNqqcARDumTIglFosN/EgRDnrUoHwZuOH/l43Q+885caKmpK2W+Fp35K
/QhmHMSDx3+UvVG3r/cbrEYbniJn45X2e2lrNUcj/h7/IYC9yfN6cDZFPK1K9YZ6fL26dYM7yScr
etG7ZM9d6/z7vN6LIyPCyELUL8eK4u41mkiq4PaXREgpp3n27/TdTfsT4w7a2Ovt1AOCdu+f+WKI
kzcJNRS6GRgTJSkwrALFgz+Jyz8TIIzuCv3zPDou6jc2Shac8ZC++gpgT0AdYVSBxl6rLUQXng4f
1I8CsNeeEc2Q7YrEk9zIrx5WOJncPrzGpSin9nPJHF7u6s1DGAFlSID+n9nuRG+Rf6VK+lygYCnx
8Of4M/k2ERJD4wiAMzN6wbVR3QxgLFItSIaQPzIgKbAvO8JBAOXpgfPV81cWhYwbC38czlmBj9oz
/B7U48WoQc/5elmw0KtHWpC5r6s8ykpwujv9yXr1LufRdVxp2AXyTYiee8Ybd0MNtG5F5UTHCaQ4
HcmA5uoZba2Ksmjr7fZOW90ZhkXY/UC00eicKaUViHRnTrAsp9M06CNtp75I6C3yl4HIsBbl4Nfm
tu6H+5mYvfWxheKKZ/Oug+39OKNQJCl1jeCWUBcqGLrn7QfOZQTFcLq3xugZsB1byLKpVOoX2Br6
yxVmWVdZOtdwX4490kX1tayUYSQkZqsBA7gVQSruP5qhwvv9PQfalaisHSUJaQxcqXJZ8nKlhoq9
4ltqA33qOhepUFq+J9nKmvZQbEGYGsmTdlbBQrDlYEuPmU4v+1FYx2mLQSMr/3qnrW1fgj89dkfg
JHA+7lmj+W68egeU3+1gZhpVd+p5sMkcHegfbxBXp7SHQLVV/PWgidYxPHnAqrjIWU6zI2cxvgB/
0yaJ0/lSre7apdiEieqT7xQ8HyAXUi6qD6n5LzLKsWz5IgvT0v4xTId89EO4ckIFI1BB3zO4HwRx
nL7vtnTpHGGEKuaTuatKq7PEER+QyGObxL0OAGpquFeWXscVGKaaVvh4e4TKdEIfkbQ5+p7jchys
KhfDYwmpl1FZZP1h1wcmrromIC/6ZUJhoLm2uaFSLW/Bkvk0lkc8wjhPls9hej4JnStfLuMXEf09
HAan26tgk3Diu4q7pIWaXOQZrVo8DynHn3zFCGLTSlMdnmuoD58iHuuLfBsVu5nqjbAYDlURYxQs
1CSml+X9NBmO07nGKd1ZhTEFCOEDIOt6KEwI2E0M72ulk05+0vtvpIgoqt5O4uCbjzm15gv1ZHzV
u3h/vxGk6Azh0h/Xt7mOmjo/o8pEtKL94JrqV06f1/bvW9KFfsZogUXJE8c6GXpdvwSK/8BtHUhd
9VaEPyA1H+t6ZH4r2yuA2hJKUcDAC5GSnTgEr7K0LyIDSmYDSaFTeDqSxGLg8Q3iCzHp8rtlx115
F8AUph5OzsD1Uwi8IdI8hkM0xXjU1/XzTNF+N9MuTImb5UErF47Px5gTXcwMJcS7ccI9wU57D5zh
m9IwGkQkeZd3jHjfA0FjstSK/ixv25KdCMmNRm+fG3CqC9TjWy5u4RktrSZlm8dAb6DNUp8FoVgv
oLdOJa8wXxj89iIsad3rHC7QUiNxbxmnqAnLnNjXJOptCraSZ2HYeOZ2Djb6sXTw2l2ptHuNaGqo
Boi9F2sbXVcU7oa84P4plieLxC3436ctdnGPmBskrJMaedJrZv8lShtTX6Z/GaDuzRrYChiLskbd
dHEDUGDeWXkl6YdvoNgOYH5M0dNyGhv3iZidps7z9W6fPzEuiFSTZty+Gygfij1XM7/ZaASSOe3C
e3OwTatWpud5pidv2lbFMLABSyhI7As52zSokhAbUSc6Ff95XwV9sZnmYE644mS0KIjt1Ez/Wg5M
d9vFfRTWoKBRTXD70nIElcedXAS+f2SlPq3J9gZnJZ3ZxRrvi85TqdBC3Oz2xA4SYiROgrNGkAE2
S/sUHJIE0y3GmAo4PiKXBMNVQskDGwVVrJI7ThhKDbKhIhiWdjDyIUnFwjngeFWN8NKsN0fA5k1S
MZ0B6qyFRlvRu3QMmowlmWcgR+T4Y0e+HxvcSw08xTjkJaYp5RyOZSoS1pb4eparmjtXJiKrGng2
D/gppyDDBtzV04fbndAQkUa6FOntAHluLd+djvKUT2dHPFcmNQ6RYbEmgXYqiErHsPa0vOmr4utr
fMHvxNoenUeUph1zG/AVPLw8W4hzzIZB1MVXQteHduLG3TUBO8K/H1cKzqEYg0cX/1v4MVpJ8Imv
LQEAjqNbaMv2Gk14XnWoJv0yzw9r/OcdBwzFEY9xVH+zrb1s8El49/wwszgKMNblbBK0fKRzO9nN
ftZGacm67+Ta3/OOOT8qaGSSfnpJT7+tmrcstwng0ZufD+vuMveKmxYeoIisdTwk+Z9/2smZMeE5
l0aNhpZ0w2PEChPhfhq7cXBPC7Z/xHhFsSEYE/+pa8zrOpZgY5WW9ZmVsyJEtt2q28i39cWx3tAC
8rLSR62uytTLT5Cu584N7MUJ2Na+Nzqn3owRABr4COmJCJvbgT/o7R3ZzmtP9xhdK57trZdcqs56
8gso8n8YDap0TWjmfOG6DRTPG51fgY/ISiRF5posvp9ho57LNIte5Q0v0nO5dow2GfWPIpn0BX8O
LWT6OmTRkAm73giLdBMQbu6JHMI8eUGV/F9hTS+lL1OZNGZF+0IT/EMTu7qpsCmlfgaykqAqoxi2
iBRuiA2ndPUaobL1PhC9PiGMhqd/UXnUbsybyPii1fXyC6HY8Odt0YZVp5Kon/C8Oh5KDRMsf7iN
fph6JTEycH+O5gGbwF0ZkeBGbc92kS0pTshZjCyd5wTkh8wSQItf7dkJu2DVbnGYAfB+j0N64OA5
jhh7JHkPGaBORGRJngtcRDuKl6v/wLAG+D6ZQxSnwsxHGw9fOM7IpLPdrjMgQ6HDJWtmXjcQfmgc
Ac8hWR4xzal5b64f8rUmfdJ7BqGSE+Boe9GeEmApWIGdPfC+ygAGhNHCnGuGity6hVqrU27YUwru
ApCHUFD5HzhWxuvs8H+s0QvOXEs0JQX2vI3ghv4BDPdT5XjzQuZjz8ovdwfqHkdjLiS4163JThGR
P9DmaJSLa1ewTEm6O2dce80w3iGLTEIybl+hUKRCsXp6+U08WRgTpe0eEElEsoBxT4+L0c5w/qfh
KZkZdmYJz34+lRvQk7quBfippggrkdnHDT++VKsUA3PwyGl3iA89SQVZpIydnG5DXSW8ITqaRJUj
GXkFquKoBjfNoZsSmu0URVZY70hhILq7nqnPJEO748G7vsK6qqMwiTgnjtHVnLneidmBP0jmmMTX
FWFtlwr2CThmoFVsgNOOZKxAioKnO2jyuluL+Vd9EU0kpE3H8S867+AwWcpNEsA6dpZ1gvr1JHZo
BuFcxExKlFdt3NwzgGgI5kfT99EV1SVwyu4T9eNZa3i0FTwEqTfBiSdhprXg0HN6wnAfnu0Zcbur
NsoAadpMHtKOvam9n+yHT9j4zd2XjEKczS4env/rPskz6AFdgHVQ7i+UdKP8KuqWYw489OResWEc
dc/6Qprlx/aU3q5UIbNs3chWv1ApgdtgsP7mxTxvbrE/+WkMufkqppXfacLAwnnZFZHh9VijlcmY
UMq4p7kYnulouP12/acL0iFJqv3LuCj7JcAbdNxCD7mhEhsD4uu9lxQEOAg7985CODyrmY+rVEja
DF9338YXajbF/evCjr5xjEyL0uFz+CGDBtSaQmanO6/lQXkhQ2JBmkrDC9djpX+o3cGxG2vdpQg6
Ml1YX2+dd/yyFaj+t7i22f8T9Am/wrqGcq2zolAzNWpK9J0CLA50wNqfWB44g9YHsIHBr1AtOGxr
mSfsnzKBP+X/fZvHeEhTPx0JiTIBWMj3IGpypB8c9yBoNrj/p5cazpJSFJFEwD6U/nKVCnY9gZeF
Y4g0d+cBa//aZGNgLK3RZ/5NDmpq9q2yQo5XpVRzUM9S461HhE2x9ulYWJo5ZmWemV/nveDXiN9m
RKXbr1Z+K9gwuGd6ljusRkB4/OiW3UGe8e9Vjqg5PO9rDKnq1s8qpkSGQ73xG9zX36DtCd1BFePz
F17tLjjVR6AvMVXWKbPpSKH0SCplsqXKfkoL3dP6oniiiWRpNILsrP86OgXyYiSO/F3Wdmz73Iw7
QQrgLza4/bYd+ljby3k0BQAz/Blse1/QDe7sQkXYYFnNmnM0BKiTrf+r7jzkhK+V7iTh86VuwKH3
vexkLCx7FG4fO7Fvi86e2CCyXW5YlY4XaISMUiAgqvvmK09BgTu8QyYodWct++tEArFU9aZ+E4zE
IuwVOQie5cMQ31sfBTLOmFeMGIYON40voYfmTaZsuxrQPQGYycLoiP60heaBAO/juPk4dVYVJyV7
/qoA/QgmWBDW068VLdZtBRDrWrTnDAqRmheiSH3VSvdIvhGsWlGz1n2ELBXdnQkaj2D59R3RojtM
YrwQVLlJAoVf/nH3yCbxPQcK9lFahjJPsU86dbCErEgsY0tLLIOAjox4PDnNDFo+pItrZNyU3voD
qxdf0dSS1PLv88eyhFQWxD31C14rh/PtVg==
`protect end_protected
