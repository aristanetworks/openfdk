--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
BfdPHLnW8CW6hrg1es/M9VyqXbAgdbn7R4Xci726Tx2q8v23VAN+BAdIV/4EIfQG4O+d+EHK7YjM
3uEbk/cqnR7f81f/vRZJlIK4SF3p+lrlPgGP9lDxJcwoWWunSLs3MqJyoMN/VVDEEeag48KQOuuj
Hzo+09OjjP7Zc835RQBnk6Dq3Awpg4aMr1U7InVLhp6qow4biQyLtpgacbZevlUJMO5E6lEkqEfg
SlJpt0rlmwnLnZsiYyeQQUaZZ6tlETReAH0jCQ6+Gcq/PwK2taqHK4xFj8vFyrMP9u2fx4L98wjZ
rj4WXfjbyStoYxBJKlQRPBiBhq2XaJ2vK455rA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="v5nmE9Bn3PaAabo0BfzpFblQ2MmiQ/BnpcqfdEc3trU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
m7xgl1PYjoowXGT9E6UyKE7EstiIZy4lthR/plm43XYolSX57Y2mZlbqlwr8vTHuI9C9R/2o6yZM
ziqJxgEqPYIEJY1614HXgQX5Tcmp/PPMAuKmG0Cl6zoCeE3KCD9KwVckC2y57mwd17UtctguiBwg
dzGiF56hhIgp6wcekoWdgPRG4bad+bhn+WqQvoVcCU4bEXlqa33AxBUlKVHMOrkjX/057FQJ2L2s
N+nuxW8AaIvs9Smw8PMYGIp0uGSb71eD0ch6iKffQtZI7qHOgtyrLhTpwOu5HhoGedtDYwKCto7Z
WZOpjj0xanbMm9Uwqzijr+WZ1dUi0CmFxLdlvQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="zsvbjd2Pwr0qTKG6FKvisYbd1hJdakRlhN4dmBudYyc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
uPvYEvGuFKBHtS4BCV9uI10cBCJL7oIHkVMI7Mx8d2Yx4hIHhNAwyk4YUoZx5LY9vlhl7nKedEEK
7MUZhoXWKDqHExVUqZSAH6YOPakpUMQMvvPo7PDJUK9tIEju/XV71Ke9A1rL2MYryrs6zT9Bc+D7
bb+ZgHxRylC6YsrbRtcN1IuLJW7U8zin4YPbhAiMfT0+PXWda8cGjDnnEuaIeV8IJzHNIIKT1HMx
WLv6y31Vif0UxnYGRIGM4TpvDtby+5j5ZSRFfJWm144KmFhxIOXxxEjBTqyIeQEDwNHBabAn0SEh
EdWZUdlOm0ldSuseUHZfQDN+38rSBAstNNK5EzStpkJ1epgocOkBOCipFjyX+KHSSMfbOkvQhssW
B8CcFpwPIYCuuDIJt9Av5dyAIZcTzVTWdBWjvMAI81R9Fb4UWoPXxkIDlPDz0iwdzr9XHu+zCHsq
pKT2gwnc/v3gPYSCOGTsGQrJICVOxZvp1VEp3exSUHpeWeAF626NLBhEB49vPjfV5bbFHDASBJn6
R2Q5kADDccC4yIBMEpmvFLaebPpZjoEefX9F/MCTSpAyop2RzOIKZZ1pqicmaOSTzsHgTa1ha2C4
pjnIIeRzHxtXKj8EhIohJkefmQKJyk+XpP/EtsrjL1KLSEd0ZEiHc5WzcbSES3FckUKhEksV9b18
cDPBqGqRxd0mRWs+MAxZs+EGJ6hqFgwZoE57fqSXUh8c0ncuPBCUb1rVjSq99d+q+eaON5M7PYhG
SPbHMpsSd20vDhKECIgXUGtMsCfLDFNqEvtm2jLXlHgDozwKbA7D/zP1II8+qTWqAa6O1VEwQ86z
fPDt+TH6j1QwSMLyzhJ1you9yHlSBchHFLkwMkoJfFaiK6skqhTb7d811zpsyDMoRDpXzyF8f304
MgZ805bmQoB84PRKDsm2DcaTE0AnfjjNarhPyiobKfhjOg77tDtl7zT5AT8rPO3yl0M4l0v/oucn
pLCSntwxK7U01rMOASl7z2Zztpcl8SNhG0Hcm2VyiYn3Ahe3DlxlCfr1Ffug6SZ+FeUfPZmO3ZPO
CJsEjbynBdItkSyzEgNzbrkcPDz5Pi3E4OH6kgMU0W+nGEES9Aoa0ffwtAIkV+seqByRglpMAQ7Q
fbtVrtyC6JirA77jJo+z/71ZYFkB0BD90IoHun3NJ2wTxDua9fG1SoNyhe1csIpwzWHTdh7r+I0Q
+6diad1vyiYCW25G7sgaNODiC40DFjjnmt0aI+M90snIslFYkus/gz99qZk2FIT1O7sWR8nQat5y
/2rDLBVCaIsaZYRBjQSdDdag57sXIRNVbpzmWnvKuv9viaB/FMQ9/Kd1mBv7Rjk4qc8wwhXpM7PL
WwNBS+o2mQZMuTWGWKoeE8iGt0CHbA0fTwSRBDi0TQVt2KNulICtZU+JpfpMj/9y354PyLBysv1P
+YPyMOE4IXPD8i2Aw9J7ZLKjracZ5wIjxCiI+bwAzupSxlUxMS3I51EDn4uhvLjaheMOGOvALIde
smNrq6xWIxGge3PJZyar2NT6waJQp6LseWIDhhsP3KFM3uQTIuIPesBdZWjq+pKczib0SezI/qqE
iLJMFcG2Ek0mIvQi+0tr9rrESmJinhSgXs2/SJfZKlr6kdbo6rithsmbUmP8ZRxxps45jow46vyB
dYp+dKscby0y6cF0XZxFH+SKediQUsCiDBVYrT12MMaUzkQNwHQ3A9Q/GuDzDqAkmSgSnWqIfrWz
ab3/Tybt2rV1ytWs7wl+QyAkW2+Ah14B/5dl7L2QqfDj/Jssir6LULGh94RsTyInwSMR4jgYoUcS
CSkCMLxffrA8XvfGY5NdTXh57aF1NMH1ltLKfWd0OUIfJhU/YdNa+iGDqGRc8uv5XKQNkXx6WhoI
8lTo7641atukhF5STUC6Mm146FWMHNbr+YojZnI4VUKrSujKst80jdez2cTVEpxLZVWF56J/ASLF
flMRqs2jWVriH/VSE+pVr1Kzv5jtxQ8yR91LI19YbWXQ8Xf/d4id4MISwO5sPgFOTJ3UDdiOq3GN
u+a5GgEPf2zkzlKOXUP9seyFLZUe+S5N4t+T6MODyh+Johcsa5GY94JL9vW9g4o/5c5MIVNp72SQ
/5Dnar4ZMU78djLcacm3wZPeA2BWSyQdFB1tQZXczZ81MV3MsONaBImUozl0NA+fcElqsOimTvir
R06EwOpUqn+YZPSLJIMqhEWZe6aogmjDXZgevGaUVtGURntnsPJggI7IoLNGNweuAhgqF3bqM2E/
qm0olT7EPPbH1NH2Cu+v6kBDVmxlfTsV6fKKlgYOTnXiET3kQLXHgEWE5GtmoulT2wnsVIf64z9V
9P1yFHF2/FPE8lOrR4V6SZQQGSDaeWE9wXizSo3NO9+TajtAlAu47TcfT97Hft6RTWVFPO0OCPTt
Ba7N9Ja3iMvOF6AqeTynxRpKOQY9b4JiCqt/Trwuoiptx+X0vGiS2g1J9zociQ5hIH4IUkTBN9vn
7lKF/Y1T0kAKm//l30Hi38Ghia81n5RoVEcvAhvZSWBBC942pHR+js+sZbsrff71JX1KXgdltqEL
ZinZSsP9yGmYhUayEp9or1u4eYPV3xXflYVrxcjIA/OM3f9W0G40gB3wKSyY94q7AL9ynVWtS28O
jb0vpDR6milMYFaucSxbiZvS93cZgWC2V1/DBbBLzEIgi7K62vPXjrKUR0+pBDJgNIxIJgXv7u4n
t0ust7FjhpYkoFa2iKG3/OQi0Jznmkm/s4k+m44FM8uMfRWawvDcN0yxOlZQ8glBusbSqDOBdho9
xvWt7mi0GT2eLW7dwCKulJeo04O0OyfToqOk1HJ+P3XBn9XzEeUZYLGCNjOZvMZaQwCndLpcTze7
2k8666w+F0vw/53PXNls4VNgDcmEDw8F8ffmReRt9B4li1RXo877ZM9CRUf/KD7LQcnmotkN3NlA
yQSFDG1Myzd/6RSOEVFEHKwiaN8MH3L9KvqNQFLrc+3hL4RodRolWTVb3SPwUcn6ZyrPJ62ioQGr
hYDXoCp2mTiDZARWLMWrGbH99epclI6AbyhDq4P7NYxmgYgW5y14R5SBrvDAk6ipWWGa6h1YJjCQ
Yf2Pn6O1X2ryK9cyu/FXFHsrMdbNje4wjWPxDS31gcgJC9MLRi+ZjpMUR8kaoJEjGDoHPfgpRPDq
erXLU0h11t14na4Atx5hYkkf13TZNnHoCgJGdu1ddrWG16Cvo75xAvVeWtA/ykuqPhP2vQsD+Kjd
ddMTo2SlG5Ru2C6ZlUYCwayc8BrgD/wZ8nez+0qs/Sl5MQtd35JXCwMQbWdXqDPIh6pMJt2yTY9d
Lo8QPbHaxvdyarDLDo+kQ6d2M1nITeTXD/osvvo+FUJtk2qhyN7NmsfIA9z+zq/0E30uqPQZOtGe
ypre2D9WwRAnHG59JTn+uPXRYIQyQyc+ifeWolLmAtw45mJbWb3OHDQNlNn/Z3xUQ9SW52K2RKGP
a/b/p7DAfAQ7PFtnLJSXMafbRw/vLmXCP6Rx1kweM9wTgnR0bUoQnq9RQf07XAUyadfFkaEZUMpR
9w+zuIochCbidU+qXl5q145pfQr6QJQcBouGjBEgLi06TQuFlkfV7Go6pt7cYg5qB0PNZnZR2yTK
CHicL3nU802gym6L8MBKcXWvUTSNaitLpA0+Ozyv7VXQ/jm8pCe3CP3Zz5XmxCYZfj5CCNBV2sz8
53QVMYSCYSKoBCkaRXYKZ3pSo1knotUp4nBW4rntURxNeOUk3bDn2BTG/i+WgUFwVThJF54VN3+I
5F0vAs1Yqz6NgMRm+n0QGKfX9daCvX4DQrzPsRO2B05C7VWtPgsfYEbp9JsYOyMjh+Bi2jZZiFvA
ZRtXQ6TBXEd3DL2n0e4p2x6abo8Ms9G8ocyo6ldy5RChsvmchhQKslm4SInn6+tF9J9hfkXE8AQ4
be/WsQEitRoW5SagAaz2a4FtWrW1Be0hGg3EpS+9zGmoP2dKmZh/AdKam/FLEx0NvASHoyxRA3vh
m7NCf7iIBl3TLKGNG0YjXHHP66rf0UhfLRU5acxGSzRFVKsK5+K8HT4lmDmFBp4b5c5iTv/MXsX6
Sm4ex6jHrswNphZC1hbwsMnezrnbJ8NcQ/ZRzzsu2BBt27cnoyFS9N+0cQfuCLIQCO3gXD6EzBKQ
KtbMaUy9y/rOr3ZEIlWe3GVpCYkZyAY37iLXcPuoUVOt69X0j/GjSTThK6M3HL5CulW75IoGWKNJ
qmnVEOHSSeQ7m4g00PvP5cFseFcZZETdo1OX+6hoJR2V1S/AE9wGpN8Ci/axO2759GtykDK1BPZA
o4rhWiwU7g9hbhRQjNPVouXT0heCLcA6bbHST0MGtsni+fflQ9li/qhvMQUatUT4iEje2olBYSeu
4BIPqS+FpyaEzMusIo9wFqaMZ14pXt+MQeQW4FKGk2zaCTeKG5jHYIAAGyBolBxmMtm6a+ti6d2i
vWiJzsdhtAjGBSj8Nl1sbffvlwtq0BjdiYrMU8DLP0lDXVnwUM1eD+aGvyeLEgLhiCgXnyf8PVBt
p9zOa/jqQfZP6c5iYxikb7pSq3J003HF3w+gZ8KsBG4hn5O6h8CUTLiKJBaxlhrCIe1CdOjSZFnF
PDO3tey+N0d+T7H4TyBv4hanQ7s1HvBdNiMw+1DEjFXQPCrgJ7cymNOwlZWy5TKyGekyNRrmmtGu
ec3Qr821nTeqz9yAlbTglFCGE4TgAL8OQUPM+wt5h662U3FZ/WBR+acradVzwbhWPiTGZWo2RnGK
swUeO3W///uAK/jlaCsfXY9WRWP4YlwevBzFf2UPqeJCOo3xc1GnzqSRt5PapGIM2lQvB75KlLlk
zls54gHziRpE6A4sFEbNU6+L+zXQsbuGAwzudZdlKhL/L1Ue1pFBS6pq5yetDGWfHOpr3c5FF5Mr
oko5rK1Nq84JE7YYeB0lDlWt25DU7hdVztzYE9TT5x8xQ0LfVGzRTSrRDA3K5GjDDZzHmbfw1ARD
HT2EcKqpjlxiqAzztNTxmEPNZhcxhyPGV4eFv4wjKLPI7yZ5EX4pQ/mfdll8nTlWJ4CdrevlSvgH
VEz9bOts7uBo2mAjs4oWmUVVZFTNVj/OvvpM+A4pAJFGydDKSRDXIIKv2INkOVGfDhWfzEkUjuGa
GLK4z6dUfLxAwsP4PCCkjFDL8J24GOzmvdTyRb3jQI4oFzic4n5Kv1i22iT+zb7EHxRlYsS6yxVv
0z3MOOZ2CeaOTEuTm/2K/jupww3uG1snbsuCwXxgKoHfECZ5Kr8eP6xdCHSfQiwwjlE55Jxxf8FF
xZL0J0SIlqYk2qfRJPCPcNzOxrJhl/hquls4jE82iznzNrVNYKmBFCIrqJU9/M4ADmnubg94Q1j8
Vl1EtTYpBXuVxFpMb8DuuLbe7VKwVtWR4uNywbf2uNyn9oC0UhKwcoLrje2B1m2RjDP7G75ZAvhK
bpxSL8z8U37PwTCdZ6O9xSwJWzhWwwMq/pzdli/FkYoDPu7bBOimjh7TxWOpE+XQID88Q2u87/oR
teIdbHJVMYNC7oIn0ghg8sydj3vHoyuuw/BQm8MK7zecCsKPkGLucWmfdjHJmu3OXDX1rUvHSDVT
MN8dw5dmJleY5aGsvfdOzAZ9iXudPMk+pgo+H8psKG6gsajqhU4T8gG4MKXDO5MHRXyMVFD/ebIw
6SeCk+hB7VDUqJq0TOGbWOmiqcaZddQqkrQ+Z23wOA3CsBVDi82uhyAdulz9f/yJBAxyCSTG/KEQ
ZOCZ2GsZyx9HeLFWgQX4ONJI90N5lIqJseaijjekhr/FxkUkSUDOq53BhkkyCd6ICR0nF9EPeMc/
uo3yD/3fer7/6M6k0eiL4DHSHW7fWQZ8pUnNiIUMzoSUNknATBHcaODs+0JS6k3eB4E1ISs0uPh0
U6P3VXeBboSsoyqwU8R7XvoMbNyeSX0VyttKEuM1wdwn1miaxX8PMUHVMx2DVXh/sje1XNX5iqwF
B3HpQ1tWyVpSINNLtIsC4gVJM/aeTlARJy6F1hCrftmqkCvRwtx3wW0KV1Vi3IXZR7aEhjmvf/Zk
Cnttj59CJGKqOKVe+KScn3tGIMSmHvBVk93s0to6AN1ljbTxKktzSA/D5GnBeLF9+D82/BSM0sQA
a+0Rknu6JdTCEElSzRZYV/4RZM3VRS5nayKzx1N6VrvPUBxjDnyR1TDPY/s0MErh9Zmw/2+27Hpq
8+EFJEvxKPgHt+LNtUKg9ckjxHlZ+OW0cTEx0XCpoDqelMzJJ/Sh6YDHXDMNnL/43wrRNzSXy/7E
R6MYc5xJSKTel4O03d+RsWBmhllUgMmFBgvCZInuFXTzr35xTkx3562gplqme57NpkP+sgROmUMn
gqDy9Odn0Q6wYSheqgoRKjfLNS5AqmIHyuynWpekRyNGcYFDcCvloZSyDJ0y4qPwOSuvqgKpIhw2
83kb4qxLJ4suZjwcm1lWRtxR5z2CnDlYMbhewCFdSMQYQ3d9T85s9BuaNZoDsf2VZVkvZc9hlgxB
103itXXSPDsw/be/OxtZgRck0LOXAnQ3mkhDoMQ7Kl6c6jkXdf/yu6fDVqCRWgc8y9lQhltbZj+L
Yu1lvMYvUNFYyATsnAtNRMcj4kNsqsVu0gOqtHtoNpP62PQUppdjlA4mVbSTRYgj39Ceb9ldnrwk
4AepHwr/GlYrlGzJyvCRiERuML+DluAI9+RvqrP9TB9Vu448uZjr3tIHqwu/ZewabHThZztja/d/
hmlUDexQWOFpdgM0T22rFTlSqmcIHC2X+6gi+mXUhQsM8Y4y8kbGGPuJ2y09aVCNP2QWBOODm1Sn
8u5j4eR2ZKwy1kLnjKYBVWMMbFnZKfCbZGE26W2sF4Zv3cGCDpJLfdEo1oSOt8EPGy3R0wJ6fCCj
x9e1hH7kUo9gSmgmSedklHRdlKWGklerzeeoI3UuHn+RuWvHmQzuJKxPa4GfJ2Mq6qv8hwv3t5Lf
rDLSTTSG7IHzgcu6kycVcYHb4LUK00nJ51Gja7HrDriBfOhqBqwKg/T9ifNTBQLgxM66V+fnslx3
ZYBTHp6eHnKFop4=
`protect end_protected
