--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
KwLLE02LlfiJaOj1tiXlK1A6kFOZ00nZWZbM9+v9ErL9YXOagvKdiPzo50PPy8roTJ0ptUozhPr0
rRiv+tnnDEqbzkCHQ8SP03ExX6AdZukzhpgPhSfDE8wZkBVRHYvAhLMdJVbDVn0dPDaKt5MdmJgZ
8ywZ/Bv9dKD6yfPl47hHXkZk6Sj47M6irGMG7L6Sy6uUCB89k0aN5tqQei9GC6TBL+qC12jLFkp4
DSMna6ew2jzZZMT2+limyw6GPez1tYj+4dtnaovFv7JgIIiNaS6xcod2Ao7bAopNpzBNO6C8Lnpi
V8jAHyM0WqD2999tOjsWXThZRXlSZ0bWBprWDw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="6WGH5o+yhy92Fce60AZdn+RywdxStaOsPQN64nXeFuA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
lMp90cc/zD9/nShekX4txf+6tyhKzhLpyeYLzgRbaG4TESkaAy1t7vQVAjUwg2OkNhsS0KbJEvkk
4qpY/JZ8ozYaGUqZLA3bTDYXO1OKHhFCcupFNnZfUWlSjXayBjUmk4LIN3oqOccgoNXsjsEotf4D
goY1ZpHy6CKG6fagY0PHn4mc4Fm3Y9SwKTkYCxWeApgocIPH86itUNf1yOKIBLJf5ZYra010ZE7K
TGg3zXVTHHp2nccFVzJS3Ao+F2we+wx8dGqcITzpT8PIK/FuWtBMUp9ztnNv6pOqBVt9Ih8/qt9z
hjYzj835/qV/wO8BG7434DdbDUPTAdyWu9Z1fg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="KIrmHueRe19qI1ImGa5+epJmX7hD0rFunVbos1JV5t0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4496)
`protect data_block
NOdp17wp3FnKoLJaty/XG7hQ+Kpm3jbKMGCboFyPWKmwIWZpIrX6PZb5CJsVAeFYf9Uv3ZqRz1rH
+7uf4GlWUXUUD2/nBnN5AA4NfOkuMdOfqu8126J6Ck7vG6QXA529YaqmzpDDmQlMV+MK6xLOZgpv
9KvgOGeFwdhnILAJ6ZCcSZeHnFskPM0BS3qYRxSSlIusHyXpeKK1+QBgbHyEB0r49sgerM9/II9p
dsWlyDIovIr8a4JBoMGtIeqxQ2kU5fX9ckpVEPxrpVFTV7RBJt9YtcQVmpKTYodAMqBzWaPQm9/A
L2ZGBDj0/bJHppvYzKhlo9eniuojrMnVazNAR5Mvj0RgC89SsgTd7XNSQ3nNViCGmC1XkkwKcS94
2+fwNWv8fDgeueDGzpiFVpsoLHlp8Ak2eiThOjyBbXYCE6yinyR5HEZrWtDENwulAe8DtP2HRgWA
D9XHkBtPa6xUcjMqDJVkaGkhlzat220BCUsKOQZTkOSQSPPR5Xl90sBQNb09tWVzBt3FwU+tfUuH
/IBUAOYXdbvBcmz6SrlTonOumifsx5lfq3UL+vKAnbYXyxJWQwB2mweOiM6m5KKp/XZ3ByKlm8gU
wdd4w4dKoYAOOEtgG0jO3KYTUHCJj5G6W+Xhp/6uyUEY7/S9KYb4bw0sur2Yw1DAOFa+ASPHs4Tm
KSvqRhHBcngoK8HxDl/sv2W4lInXlWHhnA5baEW/oNURgB62eeiVKYPgLhmeSxPceussRNpkjEUD
YDfttRITLBRExjNdzmqlEY50QHW6osgwAVM65Vz1Zt94OOLGx8JUrAzGeXNMf5fSsfnNfp2uWQKt
iiMHUQJstOzDukmPuGecyypdS0p3UwObK0HYU+7cRhVbagjDqIw9WN9lJBJo7iak2AF8Uy5/+x71
EERQXgqiO2ogZqVfMhOLc3Wb1evT4rJ1hrz3POiGQjavEGq0RZ/30mWrpkkCVlpNlYkPA8Bu9JgS
SWQjAT5eAhly9UKT4y79Y6bJJM3AzHKhyVuA1ri1dH8FoV0mUXHxVlut8pjkF8e08OVySsqcOjr+
nl39z4F2OO6JJYwy9TfncLWJ9LqqasvTBJLja6t9moV3z4Z65ZvgS3CPAtVbdRrYs3TFYch/WzI/
8J/leBqJFWsRlpVvMHnTdBlpnYT7L+j+wccZFYBmuToL+JTNKpvqXx9oPcQeHNgV2msf0SXV/qMw
oHmTCyQOp5mpibQ9Ce8cPUGfUtMbR9+XVXoHOs1SwQ3xBIYqGf0Yac3uPDZDvTR00Mj4k9S934mH
m6b4Ak7JrJGy7wkCENWw+H9QevttcqF0cS9UJKH5S5fnPtTP9vmKmCUjkkbglKqMVH3xnbxy/W7j
cjuxxQs43Xid89OrsyZGKj3kQchhmnbQESyqHTu7nCrazohvPUZEP9oNtmMIx3/iWKmSJwBvLT0I
aGxfuvQkI7HmRl6h2lHcC148yradV6yyxMexSie7bNN27kLMQsANdAE48R1CsT36AaXX0V7Gq2im
l2lzl32oBxwv/PuK8BHNuJUfdY+XuwAZnmT/2a6x0lnM9vwL1CraU68wj1odiLzzFH0n+eGhMJaf
5X+EJMP3SjqznKgUcpv73HQ2JdPDOIDBWFV+/ErEsNg3zkLGQ0ivobN02Pbv1oOYoif1jhzVXyk7
UqeHZkeZTAttbySfWqjpQxnXq2GZaYULKegjGMhqRoS1ldh37kp2wQwRVVhCxhoyGdxLSFqp703+
vZoxWQzTpSPlqUopwbzCcLYOIKWnskU5u4YLvm75Jw/0CIAQHo4ujQh8MLRgufq001KzRaRukdTh
DD9qdxpi1ekkISs4GUZzw39u8DbJcnBwR8Ajl7E5h4/GAT0ttaxX07qgaEMjQkFZbuaKcFLSqE57
vzHU2FGnHzTYKpkOVzBsMqNIYGkMOm/NxrR31I1YTX6yE6rXe7eSlwLEcethn/ydS7tPaoh9hqeU
C54+kV01l0zHoZWor4IRhZFKM0d8zmHfBr78FE5FBU9Lw25SWs/aoQBNEXMWK9uaxRD3UCLnVyAh
RTAtTNBP4h3Sj4UvKfB9e6KyBDvncXN7r//fslNYd4T/lDPoqREjlI8YMuk9Rwf4ONMaZRxo6X3L
X0Ge7RjYo9eRBFtS1Gr+Gh0Mb98tqD+8Jyj8HqqrfADR2DjOE3JguHYkBNtFHtYfAPxqgwBzKqB0
sRSkWpesoMqqNJCjKXCDdYt2gvrXnOaSjighAa5VvLn7PORdWWlVLHlqCs9IY3XrsdH+UGoMB/eQ
ih5WN87lIf1EE8sfnbbtg2E4/nyHSYGlbBOahNiW0lI3vwMS7zCaaimmIvPZd2DDE79KTYk3ZVE/
Vc7EiLvajirOhDEw5gX+Ru1h4w5aVm5gy7SLZFPQTZ49nlrKD8qqYyXYCUPe4rvQq4Kb5ogHhCct
uAkCkObC8yWdHDcKT+DT3ngrn7BYFFAowEdQt77sriMSQ5o8PPFtDnQAa0DP+kKhdyM7Zd5OWczQ
FcoX/crYXrU1yvlKX1Vcxy2IiCp7xtpKEwv8Yefv5tG4qraPCGkK0tZ06TAb8wWo7BzRIxc8SBUn
2qPd9NkOSH7It96+A4hvO/i/GMFUAwtI9NzZyr2Drpszu/l6bheEi2N4/Ued0zlb35WY73mTqLxW
+eIWY3esW7cMnI2D/3v1x/fmHtWtgeim4QUKH+0MQ+agrnIPvebPAt2RO1vx/QFVNXf5F/wAobNx
y62vuqSjgDzeE6/cid8q3A/WAmBgzIA3LC/KI3FhcBp+dTnk3EwtdH97FZp9IPElNwjul0PVRH2e
okve1Y6pNxpcNAHxBEp9DFjaF7KJIaTweTUHcpD75WVreANtH56ps/NeSj+mBuIhBcs5ExfDF5w0
Op6Ak0VmhTX7Jj9NyOyR+uQfOxHb6FKNPRNQhsWRNy5n2gdhgEwfp83ryGqdDHEfYJmidYkq8ano
VlW+Kmk1l64qJD6kQYTgvnEcuhX0w046+1DmGHkLil50pda/fp9ht2nq4LLcrdy0wvZGCswggase
XIGopRo01MKdFA9vb8tFDNJODSuhnKHf42vkMeUUbFz+C1QxFGe2ZRLz5tuMJrdsKQsd9rQEtUj4
uk4NTJacYGN0qrGP2QGkcCFFD+CbZNPCW4PzGJfFfechXkGbcZ9afVJBByTbpQgyAW6Jb5NlIu7X
IMyt8MWZW9RU3xTvFo8bnzptS+efvW60Hq6G4k9t5FQTEGfdo0SqnZokhhEiNJTilIfWPI/OCYTL
iE5K2iy/8ejNqoNh/hmueyg5lhNeZOqJ5STJ+PxxrBuKesOS6Zne1T/MjZw58Mew2kIOF0Zm/7XW
3cFWpu2lX4tntjYyJXMRCQ2t8lLkUMi9/4dQjOsIeUVGHYdZxRWO4IlhUuEu6qZ7MWXS+tsvZBJj
R25hvjLsd8Lxlpi6298VmE3W9JEYVwkXrkHrsJ9NbGlMD/HA2rrFJg1BbsSO+iIo1YgyBlDk59Dd
Gg5On5RrJHaUhnXnhY6+zlR6aRegIsHaFwf9sJaIMP0SaHtI18sz8ZBxvRNg6gVh+ZxdftKL7jW2
qCDdMAkw4QFGx1/BtsGX+MKkdp8lyeuf3ONkTkvJqG+cCJXhQhXvqGK9tHv12KHOsGHjbQtNCc1y
qYxXqXpS8UZXqjpipEWRyc+bq99mwp+sTFLpsllRCSSaeAJH1Oe5K7dLEKkwitD7B6Dz7YqvU4c4
99jpZJpWgA7xbXUHQbgw4nRQHljMjqcuXe24jNH1plzyR7Jen699Ywtc80deOnOF8Vux/BKZm0lr
CRBiN6qIaEm/o0WlEGlRMJnszjuA6bq42Ofr38EXt2+9uH1UmGyZMXFGKjHADWgbHZF8rTWlLitI
Y50LufQ2U8J+Jnu8ak8dRVrsQSKWlLNjsO3XzL+ZXHxL+/YsS6VrFEE0RL7u/ENxH8ep8qcWmIhL
wq2xN/q2uKTc5xoVBS+gDhZz2/Su4sCiJ855ODD8vxo9qdSEN8VTWLhvQ+u45OeSe0ulJoYaLahc
z6cSYq8v5C7yxqHKKrZBRyGx/zLlA+XJqsySMnm0jy9smcOXOGdL7XQkZXEeLfl/PKIiaIN41cUf
p24cAQJFlJB0pW8zIkiMEcWlSdx7QOcWEwZktVVNxT5i5WdaXcxkSlEO0onKI0+0WZsORbMfQxJ9
0k7Xpd9UlAhUk+NQSZjrreMnNT0oGlHWvrzZg1UdoL/FBC8mWxxUKtyqEDE+jhacnWpo/HYGiOn4
KXLEpBAStTw9NjVrV1m+M4PL1MsXdR+seY0wcnuiZ6hGO1P/RsBOavQZH68KYkS1yquNof8UtBw5
fuwroncFgU2jjKfobMzZ0urxDd1LmpZwXOybPEhUQA3is9gVLWuXBGLyAcgczluuTVUcq48HL2gP
s4YJ50gdJ6puGc2XPnWAvUf14tEIn+gzFKWHRYgMoggXnyJw2L7ASe6pFvtWXMxk8z7HndYyOFnL
/0xLz/zrpj4B0CZV2Ty/7QFdKbHSRgje4iGejMNJugtxxQ3MRzRHrmYNCvNpLuC578kku7bYxUMs
pzpTyNAorA32kJdmLva7NR8k6uxZ+cHNdialNOzUbfqnRMIL82omDrTO4CDxForEefs4gJ/+ehsq
ca1FUZ2tDIOhIFkEV4hZClE4XvXRePcjs5lqPoaeEnpjHkJF/T6y7MWipX3NxhayOCeYs9EPv7qX
0VNEycJ/3xCQ6jgt36yN4N6ECE0OlBVSOTQqhmdKSjhJ+ROfnAVJAdi83oFmfe2IsWikGPYB1BYt
xV9XN58kXN0lfrNv7Jrd3Mxq2qqoW9DJ3kVR22JsM/2AwkAvE+ccR8rpiI6VL+4x0BhCUajkTNwS
z1o5DKEJ6fBbCSjaETiDTq2fycEqCRFinZPkej6vmVQF9klbhAm+C2+4loY50I6MFayIzJYMYc/w
urEVhtL8KCbdLHLjIFVU3/Qp92wxt92VVbKOjMd6vtZEk1ssYL+0MO+khBnj+m5vDGvaUPd2Ga7I
D/U2GopqpmtlW1V3pk/0hWLvTzAw5YyyoPwd9K9mLSyhxE+/t6yefVHD4REnoFKS1PxsgzNTk3ky
eLt1MsITlwwIusuezA9wmybYds+YZZWQPnml/K7i/RrYwg4NZlJkq2UMpNWAz4OK1W6ZJZnK7dOE
+BBMI/lvXSofvAT0Vp3UwbaOyb4AIiQ3sIoz9G73t5+Us/u4lT52leYriANJiPQXSVEzBvvLrgD6
/GzfjQDRBEs3lG4u7wCeOi7D4LakUe17hx6mMk0ogEiGBbIh/srxZlKkOMXFkrt3j2ZPh5HsZKIh
9WLWw4xsI0iJsh2jN6RuIFMEMU6lmpR5DN4lmjAtYPI8WY8OHPJJp508r8ISBq5sQQ6dqH7zExuX
OmO9VEq62IKiApgYHyRSmPLNkxEw8rl7IeNkNbywbLYSKKcrmlc3Na2PlSM72+wqcCuSihdHX2UI
e9ge+2TDofz40GJMcr2ay8EaeKCr+ac4dQgzTF1EDW+nfC3OJ0L+f75F+2uRJhjLp+X43N6WkNV1
gEFotxpWv/uJ1nYWG2HF0T1cgPnpGW+cMgOzgU0TTZuQ/V+lzF2orjirHR2qDl4zW8+3O4SHtAyw
TqTyEY3+hxDlesSsgTcM9hC/F0KqxoJlQNs2Zvn0v452m/6z0ZEgtXC92n0VAg2j5iUriAotbXjJ
OtWka5q0ee3ID8KaS8JKv5FXWvhWC/2tnLXNOlMaYbORsxg9f/RUbtlUAbPsP9SCZZPh7tnnDjyt
+8edKAy7U2IskZQEbxTU6LiNibxcpkNsy78cTS7ddAx6oCbb2AZVw8Uu5VxFf0w1n9iu8bFClT2d
nb10TnPuTxXWOIrUqMZOXyrjMO5ZMAjBnTD0hZjKtD/lMwUBRLomd1DY3d5mADMgh8yJ6ejZMdCh
j26tswzENTdIwkSjM+u70RfbNNEuC2HiT1Cq5nG9JYQ3WQ7ZRbYZi+vP/GqCmqQuGqU=
`protect end_protected
