--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
dl2i/qZUqQ4SEQd6YPgeNUvQXQZCv+dT5uqjA734aW6YcPFwmYnLikvMIYhKU2YJIoFGHoqy9CrJ
sfVZifKdkY1TFV2pzFh87OEYX0PlZGv5PaHKaJ0z8mtNnEd5j86JnlJe5RSjSlhhUtO8nDHVhqVm
NPkryhx+D7x0pRHjD549JexIUxhGJpxGYCHl5nCQg01O3q+UuyCqil439qu5aauIqLjYdy5CMNc+
6uvk42kMLLADB3F6hXAeo6v/ABnW1xFJgD6bm//qfw+wiS/2XsCurSBxy5vg1psB6j4WBJos5COF
hW+3v9b4AqNQL3RdbwwEASO21MW6fO0JBGDHRA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Dw2/Iw1G/VtmBoaOm22lgkTaEH3RjRbgy/NvEbkBiSM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
loIAv0H7H5SC96qitkTsg+xXhH94oqmEJbZBbqgWHHsVi7TkY3URQ2zZZGSGtDRh2vroNRhAs8pH
69cgRhuAZibn1Quw+67Aw3iuGR6X1a3uwGjtpSFKg8bNu6Mvg4HH0jYnU6/T3j9BjhpcW7RVj2w9
1H7kTFY/y9PEBp+WKwb3dzC6JA/+32bYNiCU8Kc3vTaZ0tbkMBr9qs9Xs/pgB4NI//zadRHD8Rya
abV7gmc6mb3FCRr8n3uqdQtC3r1goUhaUTwNJDL6C94JGNZT7I3kb3gCOtywFXxLlGbDDnFV9t1t
PNvENedVcaQ8bMDRgUx9QDhTxLEyual0JbKlXQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="uX42T2cK+wO5RTI/vj6CeJUmR0pbjm3+E7guZJSHfQM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9440)
`protect data_block
EU3pKkgTbawLRt4XPkOXsTtZhn7wyp4iwbcAzQXcFZZQ5DeK9Im73paj4umr66SaCQHmLXpvDwIN
bOxf1la1iK3VxJUGxVSdATenLV6gBdGsH5rsKQAL6BtIZG3LHpQxITHIIYtp0A3MbqoHFRoDTDJw
0Pv6tq1PiNTH1Ggzc9fVEJLuXAPvXX7WLMzlUNIv0eevqoNwt+t1qd9Y5XAade8u9sVOe39w+W72
eSS8ImbhIrvIlVC70vT/enmEoKy01kw14gD4pc95mODvIySDh6QH82HUR7CpyJBTmTHc/ocR95rX
fEs8tyvvjPNWPVKWdP6KiJ69hyUcaJE7nSATlhkGT0XmhZtf+grA7vBjMIrJpi3F7nP524+MEWZQ
Txyiq/OR4u4TGyjkni6ad/3tvbEVo+4qfchQwzIgo7JkZuBLqLN2p8B+CStk8Sh26D3qCjZ1GlEI
YjHUF3/3RFpjaxkDi1/5Yq6xlYRJ+rUobPM50JGtOfcXm3SGvX+ew5GFXufCCAkLxfmMGbXQxCau
TWs0CXgxh3lLVJ0EBd1zKCDYAqcQ1tvnlc1r0oejrxcyo8a3998dzDhn1baLMkLXCprmI0ONwwT2
U+MMA4jq0UVv4+lPbMbGcIx709S4XE9XdA7dR7PSZOducBiqebMsUkt2zfhau+U6h+Q3jf88ElxY
QHYOHpy2nKZ+Rw8fx8/4+v+DBhRmdVaPbfIpI4CRykj/YkLr7ylw5wZsqDc1oq6Crk9fSrLrIUPY
c/Gl6ORfw2RiNceIAZ84HANl/Oy0nAqLZGXbUhQQZf7Ov5ZPtx5S2iWVYJndcI1gTM6dWZJ17Atm
PtPCm+nP6WW808weQ8ZvN3EuqyjrRM+g9eU8KTelbTge25Kvhf5EO/Ui+OxVJvxTaV20EeYyiSs3
poR9iIkvCMztGPje4Pbbb7w3S6Ud1d2bULbnZNBEV9i0BNvUExGqAS1t+5J6eZ4YFC16OoPf711B
Hl1nR5mnlwJPezQ9a8giKVoVcby014LzVF5uVXtINNJKe8gxd5rsCAbo4Sm3b12x3dFRpaW41VIr
mSV9Sysdvn6+KNcl4SdLIwziHgjByLP5Mou46H5s93MJzwcRHvlTikeEdXBC4Jg/CuNkN8MrdY3F
kmz+j3aepI33sWMBqRPHDOEbZxkz+xLujTlwtrEksBCwLhr3m2fX54bSvR4eSq3jyScGn/mBnefa
+b7wlYVfiOC/tZ5uQceLd+AVGjgSG+I+bxnsKR9fZWpWpxSofpkTGQKnYyrCjxfBDBB76u8+rZ/B
W78Mqy8yzdp9aRT1lR4TbsfeEFz4NsREetk1K4ZIwRY2yJzX1kJsnfHhZ0fXk3XiRkFN01idapf2
zcg6UWCKhGWvyZnR14aDIpT1oCuKWtmnYhnewNIsDj/S9VtRDWCsArVfCwoH4Q8FpNXOhX3bFly0
O8Eboeh8SwRspXq1GyED1BjVkYBb+LTG2F6Q1rN/WSJvwqNlr5pXZ6B6aCwmsWfbI9vSDc54CIBS
aBVpQV4mTPv9HYA9JX1OGM8RNeS0PlHVrhvD4S45PuQLk8nJ7BFkvEVlk9KTTGc7NrKSUOmpQ0qQ
Wc5BZ1ka9+NLvfUyaQoOEeY7qs6gVIBLFnc5IiPvvWe02T+Z6fcayEB10X/AlW2M07Uk3Qx3yLVn
9Spd8dtobvIwfVf/e3S5PSTgyqtH0N0XFmbRSIGA0wWaYVsHzyXZuZxert5XLgFpwo9FL/E9x1ff
J3hGAi1fj5ilpZo4NDW6+N1tUzH5jT6zCvatucSXbxIhRMfETVzEsXFEZkgQWGFXa38TzD12Q2nw
SQKGOBOWYq36kbd+VTNtaQNjrsPCgtBB7XGlLRU6HdZGejEXOMGYkAFJQnc7LUllDw2JedmXtMAd
WG7lFrbwllUNQNOP+z5GC2Ykg1wqpDWt2ysc/B1aIYXftBxb5FyzdhPFnZK7zP6CIeH/9tcOqDwm
5rf7JF5uj0Mte7bN6lT8U5rRftHvtHJwb5E9KwIx5m33MbDgKDtwaHYWFWgvOTmTS+g1hHur37ml
sF5xKW5CaYRk73tCnlIOHwg/0soy31DngE4dObEU3T+ycV7JzoInrZQu/Bj6vGTZ20yGwPq95w7S
pK6A1YcufM41/F8U19xdq5/N6upPltlP9pdrzAhAPWwq6y81Bw5fcLbPbzxKLPOAK+0FAF6iZJzk
M5Ybn26lTJUwGSSRcNegWDvJh+qOcPhGdKXLk5KyjeAND/Jir+aZh5Q5XfRk0Sx20XFh6NQb6+Vx
JcyJ6jHZU6JT456yrF/9kyqs5jTJoW5ofnNUIQW+cuDQc9jPJ38ten1gIaR4FhqVAOlGK1L5nhoX
Ri8JaDiEXtlcyuy/yD8UET4xDXP8WLOxlsL4ViCaQC7i8plQ7QlkeI6dK0f8j5/7UxX3pnC5eqaX
3nqe191y7tHPoYvG+mnJUaZUtxE8/ifeCWLdG2eObeeGn6PHif4vkzdDJazjb/4Cf56xUAK9JmZI
p9wbiQVhmlO/8EJjWQnxxnR0ntCkRqCglvg7Ijdxajq4f+oS3JN+olDc0WR/Av89vWRYW34+cHzd
vDBXvJLOQHMe+S2lTYyIXjn8F9959YB08ZcNZPGwO0e0U5UunXBuU+OLUEG27zfT9T5k8W6JCMSw
YyB6s3K02iws6Bb1TQHjOj+mO2s8IHIxTbgbuLu+D1j+iSKaTvrr+WwTq+xknNNNzTNIIg/17eOE
mMoYLlHAzxMiaPnAy0t2g8sH1oeORgAVPWnS7Y2UIlsbgbvLYMfldrx9zw8uK92otLiOojslM0S7
CGq+rHGkUn6GyiIs4nmH8113SenSc2Eabyzy82NOGNlbBkrlTKAzaVNAGVEl/YaPTsPl1nAWJUtG
vZ/r4cC32rfybg78xlOC23yAdnx4qUrPn3JEqvs04Tt+/Rd/SGw8KJt6SexpX/4mBxPd11VtF0QO
fU7v8vyFbXNoxSkE2Bzo0HhB7Ec4GaQNRkG18Pt0HSXdWCZgyVttsIuxFglG4lYY5XrDnd4zjqV8
Wmt8SKkKYyFTMg3dCbUo30Swc6JykPesbgfYrl1eEB4Y4IsfJpUVSA9iPKs2uy61dJb4AYDs7Cmi
xit4UrZiLjYGj6XW8q64bmhjhYvzKvrKN1H4sIIDBJgdrtwQsifG4R6KLABjEFf2Czw6R5InofQm
GOQgpeS4fKfx/sA1OzvHbARnFd+41zVHy7j+rZNVM0Giy60JOPkRT2Fca+sbgTeedniOFMmxmFRK
myhPixOOtTQlIbygeaQRdyjWT3YK4qKPFm1ZBhsypUiRqmzkehNROIhKPf5sQtRwCy1SWZwMkRyw
P9yWRW5OC2VnYjHNbWKwJ6tUIrndpddIfFupd7ttFYQBdIwRby8uYkLds7AZ9xn2L+J1LWLeMNFF
yp07PtR5FWKErngYr6hWXkFFZkEA2AykrwhmM4dxU5RSjWx4MbYx5U27Z6lDwtguZ7+tc8S5kra+
wzcSm8T1xa+NQZHLXXsf4eiiCT0cOZ3GW1KPYZibfkSMe+Pips/TtRpu0P/bHQoQfc3IHV5f1A2T
FIVsgd8XRUMV9iaZrfxK0cibbvy2R0f+qXKr8cOa2vxxbaM8LBVopftkn7U6UuSSl9Q0BSScfE/I
eSg+jOUWmpBVPYT92r7Q9DExXF5lBnDtmIKTJYgdM1fmTSeoRO3Rdo6495ohXJGn8wT2IxkmqxGf
yFRWPgRVbQuumDmFMgFu5JQWd+8ct8D85MGmEAL6IFvFRV/9LiZmxMhiEOUnR/6QipK+IQvOPU51
H3uYB9WxeznIRaOImbODHfamMvS3YmaZp43csm6M7bVdMOJH9TfV7zSj9xP0YlUMKSy67IPYwRhM
+oG6iqf0NatQZ9gN/sj9rusmcjXKqsqF2fppnf8VHr4ptJr8ASNhD2p9nOQC16E8E1IP7VBNmRDb
8S2NG5pvdSd6PhIVRcECGEPXIk9wgOF8NWSreft31mGuuDzhSB8K+XZ/WWns9D1nsgRWZL4sMsIf
K9DchoKJWOjN94hW6Pv34nSP/Dx+eQRlYfbN9iK4LGF/lkUxfxJSf7WVEdp6iqPLkQKZgf5Pb6U1
ChxxxxnVknLT1sKIU9XYBwTohC6B84aR4jl8E2SZQMIjxDdlLB62/yM9LVK8IdxdrvnQ8nUi08Iw
jAni8l74TZOA0+bm3NJJPHrqkeRpEuCEJcbdizu2AQxoh0E9skJPrlGCMgdv75jVG0DSLyCL32rO
JbdebPQGqff9ipFS38iglnyVDI7xAwtla3RJ79ObF0MT3gWq/RnVZGDY3xtHj15h7aExbJGka7eo
23YM950VcnWeKgCA5IJ9ipQoof4CM4+CTtLPuMXyULXeH4a4Z2CMa92/u7phL79TMJ5VcSahOBbl
C0zLxnfymqfg5m5qvauB03h1VcfHAI61UuAnmJHzbuvs/iLkoRBvwy84Rh9oqX+5h9HpzTGmqGFR
n6NWuJSpPu9eg4f/i+8ekPhRtcCQGsZsT6KrfZTdgIvRr+zE5Latl+6zBOM/m8b5VCI89uGdOO/e
roduENmuEbivR0LUG842NOtThcDbqgcs1IBhfQVIAC/OSUmbw3E9M8hZFbKKNtomDEXqBLCDs7dL
uU8olRvgp8MylSOfTjAJtzjcr2N6X7U7V+sAbutpz2dewaaFBHlSR+0t5Dtj7CJ0JIb9ra8xMGar
ay+yJwcVgmG3vessh5D5fMnFBFnKTP5iuBT3FnX7krhKQmbj1A0HnE6j4shR09SieYlXEiJKG0py
WBgdg3Qs5QiHOlfzt4aTgzWkxSpkalS4gzb/Mq/zXAbDoRrfItt7s+xXUi+a/mORsftmi4VadwEE
g+nKPajOqEA2GWJ0XwVFq+R6Hs7jlWa120NQ+fhsRQIkr9K0ji+dUYj4fl5mGB2NOIxET0UCG0Wy
mlJzXb2kkqLdn9vnbItwCCUNkX+HciCH5CPvo7qyDiQpD4C76aDrUf/hJtim3vXoSfavqjwiNO9r
ER3x8vvhbK2jetQEWukknspGh1G24eeg1iNBXwtOEXEwsVd+Ag38L7IFy9pj6Y9Y2NXt1Me8cWAi
4esULDr8f2DzsPpLL0R6hX6FsahLEpLBNyRum/qxMHnXTnQYyVW+FlBgDunmXqduKoFMczDC2Yi7
vD1N+9HCiyd11XOjhc4u3B58B7F0hkHLMHRnRI/Jdb38FyMVI0LmEDHn+wwgg4rTzSOwWU3tzwtK
F3+yhA1C8kLXKohcQ7Ccxt1UvjfbPdJyghUFMir6rkXM4+LdK4lTuk0zpm1seJRgQ0bdjp6Mv/38
aoAFn58siqHWVzEdWgBgqmoHcuSaFDLN1qfDoVXIak8l533GDEPIInMk78S3TmNaed7nCOBDJFHV
9x5F+bnNu7tZ79330rW2FAtlyiZBO+QdT7Q8chuosvEqhssmrtHu/jV0iRGZ2ijsh8GcudTaVC5r
PbfnclTonSLDW7stm4O5okPylkKHdO5yGAv6s226KCS3ARWBAsCRNhqN9C/VT4yUoOJCPycuvIP4
VHlWMPqVxP8f+8HslXyYOv49zpvk8LhZnhXqSwfCKC1lJ6ngzzNocMDTqCAV2Akf6AytfKT6XNja
A2IBBAf2XOlQnLHdH4y/qcKljZGb6NzGjtfuwaoAttBaFw7XCbuJ0EIZWF2FnD3Ye47NXMshERRE
TV0ohYaOcJbHPkAXlynUCvWdPQKiBllf9Oo7nruNzV+v7GEgkwDaQOkvfEJ7vIybzTXzbQ45QdRt
CfO+vl1co3D3c+KQUclPKsG9WZP2T5gq/Txcm0hTXJ0GJhd2+tR/u7A3sFqyM6u1+v/Ipm05mGsC
wv3X+123LzqgQ7LEVuFs1h0y+yivH8d9Dq76NV7ZrlSBbaKWAW0DVJyP84MaLvTsF8OXpvE2r+TV
ixFLLBbR0sE54kCca2i9MCA8ZgW9mimafI24V+mXWVI6ZhZT0VVQnt71HivBmLH7buJcu92rElJQ
vjuXDxDT+Hthc7CFDpF7k9ONbXOdyrCfgDNZt+hh6WNusCfr4BuRAjkDNo+4I1uzFNpF+mIqCmN2
PYwbHnGYVxhmtAB4ZD3PAliNCYjWx5POuykthopvPDOsIDlLhu3b9Dg2PVaZUBw0llVtgyLg1U8l
YTmADwUPnxMdxHycoX8hkzubt7fHBzzVgg1+FPpI9CU0yUWl1JHRV3EAA4cpAyKw7Y2bwq9fKWqL
uBsCgU0oYKnr2z+yS4LmOLjhvpUDksFx/ZWxAZmZnYZJKlQ8+uNI4fCBmKRraYk7fQgTPTjDmgX+
63A2HOWcg9RIHdujVmxji3jpDPEKQediLddOq1T8I4hgy7rO7LaOURXwx+pFPwU+BSCPygD8/ivl
9oIxn5FELD0bNmwxn+jArVWMjXTL5xny96gMjTc8UAhHKBVu/qwY5phhd/C/rA2WP1DD1/sk8NxZ
Hn+/PEPmhtXnpXWJU+ar7oAbJsP83zqcY3IQ1jOKxECdGil/iocgIqV62xv+wtJ/Uz+Gt/o1XTpN
QQa5Gff5+yw93cZwNxH9/4w95eEDxNgy+3wr1uhfCThvjUQIj40WvA9NesIf3mPaU3zwXuPPNs64
GykjOJnnwKZX01LdzZTJRiEc1pyKdrzIPYHUmXbzaw8kt7f3VMMRdRbXjqT8LQOSynraxz65ErYQ
Xm+4hcgsMQc+vDwoqclzR4L163oyRw2LhHOnGgtwbrzFNIe/6EazVBTe30DQeV3CWmIr73BkKsVg
Q1jnR5l+wZRNIbYXHXuni8/4g0lvbhql3LnllhwreP58ajNk7BnY9u4sJ7A4ocREs7nQE43MW5f7
GhRcgOL2FpLg08nuPNVNxyMb7i4esDBgOJKS6IbS+3rwpPGaNlDbc2gHQd4shvNsJJJYHIMBChMq
quI1P3337BsGHo5LR13TCRo4+x4d+nZsvNH/GrI3j1i9lauw54r9GUmQ6wlyomn/izxCYr2z+pu6
SxJY9kqXU0VeY9K841m3ySMhfStoPFiEqVZg4rI+7+D61he+eE1brqlZOsdO+UKZLYoI6I+6SC83
UOnWvy72xjC2VWElr+dhFGvFAg6II/2KR4SMSFPhhln61KzzS9sV37FF40n7tDZzeuc68h4sxM7Z
OjDo/IBQ8YBWecdGGaM40MMGAs6l2nxcKTjhaEKYqUr4endzDBZJP2Hf8vZM43PwBWU6/tVCbg9C
MRfUrtRNajf4/T/UcIck2bd4Hw1VP4GSBc4vdaAeT9jLnMhbET/dWbQt0fHv2to6oBUp8zeC2qPy
P9aRW4jK+kCX1hgGk7Ros5PQlY/GxuHJ4r3sntjyaWmXclI/dMIOtGx0drCqwNTtcEsyJKW3ZzsT
jZC4ykL+Yvl6Yg/+tkCyEchHp2xLS4nyl2HkGVZpjmMg2zPCQ2mlvjmdl8Hf5qb2Hhsw74T51I77
oWJTe6v606TqCbP+Kta5Z13ntssPosxgxD5pHj1PFhlKyUe65JwWezoKOATwf2RKkj9GCjkx4980
6J7V32i+uRIRnJ+YHsm08wbobLgG5iNvFncku0AZjumbbHHOiUQBOx3dzW0ZXTfBMql6GCtuCmiU
srOXwB+wh06XP4acs8Iez+OwBsq/wBbrHggyCjM1RcuYxcZBDcLufRQjZou5rK77vOIZ35cDpNDU
l5At9TS8r7lzND5Lgm2cene1Z8tbFcJan1jHMvy+cg1Nd7lxYXOALspN+Iai6YxT4+lwLrQW5Grs
fEugfI0M4FerEUDHE5yKFECywNLwEiaXJBkKA0t5kCPfUvrhXYXs2Zl8sdAsB7Ok7A5jYXkGKWRT
YYcVbuCP1xM8hdOgy5HJhVTCHhbtQHA3gZ8sKfnPtk6/k82HuWHILS2lynao66iQFmlznrKchZhm
qlyO2Hd0aH783Xi/bJbQMxNWUnNelbYsloKCYtV5gdNLNsTZgl2JRkxw+kpa8biRLcKszgIS/r49
oqK2Cf126NylQCqpRoNkIfctBH+NJdCOMg6rTDIqY6UXJZ64TA1mhUlS/Lkz6HVCWOQUhrocvczs
5sv0Sc8Bmj8wgVKP6oXfmTCqivhzeJ9AuOohAN/U4nL/bRosMcLaUJOUe1nKfotGpse2PHHYKgVf
UoeyFT3p6O4TmFi2fDblmse460pcEno3yaLL4yqxzCemf3wbZi4J/4hQJWWr4d82TnUyTq38OC0n
tjZ+OisquaSoQZdD6pP8P1nFKOgJJxFWXNiW/p1hFI/6Kt7QqSfOeoJzWxI5VuWxq+d/6kaol/rv
dbiK9ySG1/kSEyw/sd7XKl+tYpuOY7EwOWDz/kXTVEK92cwe8DtPas5z4EmHzfizuVdka2MNEsL8
5sFeFNANN+v4JvKh1SwmqLzuCZGd2qY5U4aAQ38inRMCoUGlBc+9uP4a9WFycUntJB1tT38JUx3O
xxO6vcO4Os/lGRDGYcfCE9WJLhg5Q7WwihPK7LUNuwM5EESCQ7k94THdAKRpY8cRvgdxpu0uagdF
tA1KlJGrU3sMNwsVqWng4Fbz2HAwvdubcNH1sMeclzK4BjG8up0LDHWvMCh/Ur49er9woHcb9NpE
C8EazwNQiacJ8rdbnEtHCZh8Xpb7iKwmc/2Hm/NrmmvO/bmYckr9e+gI4OgbQR9NyDpH8HWOs8R1
0jsS8YPRMWqc+wFXbX1AGHPjvYNfDyi0p5RQGJ7im0vrKqTo81OnS74QnY4Uy43SHPRgj+wZlK6x
HnB4enBi2H72wZE8qx0td6mTQjVs59uNmy46oj26/ojTJwKOLyyDMvgv5TDCarD4JbMKVQjZZaRv
drMUTkZuedxdMldY8yATxyPwUoqWp3rmiwq+fpB8WNQHrS606QkKMaTMmcPGJIXaeDVSXnyj6v6Q
YvtZ5fOPLPzPuAY+hCet7ag9Ub6BAGtT7yqR5wvb7jo0Wa8o/STPk3IJcIlPqc/QJNPXDBKTsRsv
0XrPVUt0Avo4DexlpNGoaFvF8es6wn/y+IU+75e6l0b6A1JbQumbGurUuDLl6WxABXHu27r2o3MG
IcCF0KcJbUykemFREgTOEnuOa4Jg0q4VNMUQw97lFiNqaKKOmh1ud0zJMkE3R5LYyrUgaKh/TIe5
c9OfyGneTt1lpOfl+ijTeVjYiINt86RDGPy2WlxHRk6f/kE1sRk4rJptXS5opvz6v1zS6Xpcf/a5
mTq1aLYqvq3eS85Z1D8YDu39Vg1Qk2otSannb6ShSYWymWV/aH7+oLNUk74Ac0MBMUZS/ZW0MSH8
Okz+YVKPlhlPjJ5Vv0fJd+S1H33eRGW2fa4NdwfOX44VHheK8E8NirIkfG/VgaG9HmmDIusyo08S
fbZwgc4HRC8kQbp5oJ7TMA+7ya8jD3Nh2OVTb6RAZhBQuJEiuJ5sg6iBMoYZ48JITHt/zhe1JDF3
rpVIUVyrc8GDFJhx880Tf3/ohghEo6jfMeJyLMBtIMEMiZvkciCBXwyhxl55PHwa0IiakbAQapMu
ZwH2Mlkt/jSI/4rNd/BgnNAR9LDEqu7THTYTFz0yXMPwsQo75awCRCgR0a8XcjxYpEt07xALzTlo
ErtLY4t7ojoGU+FmP+cyj+dKgoKunLKijiq/jkKzu0BC1QZ1GAfVV0fANfP9MIKqG159ukQGMZKu
Uqfe9VLV1Hjl0rXFuNLT+RbZ2RECWaGCPytyOV6YfgYub5m2M5hWaghZwhS/fRPbyH/07cSbfHka
7LQJhHRntPQ842ZgFJ7OuPS6nJksUwuuXLzNAS4izK1J7DNW2j9sNREFTRlBJXput3fV/HbVJkt9
U2L0PrUdGj7Zi2xIt2SLjtmQlqgnhdUpVX6ryVSM/BH1PsEiEaHg7YWWhxoJLPeMLyDgNjqnHFi+
qQkvMKi3WppzHJQ4SzBwBBQQpZ3xlLUY321XfuOobV/w78KSzpkCYvsagNUC7KiDLsF5wNf0Q4vB
VkJ5mlKUByfJWXAAvkKnbQZ9YuU1Dk6/v/po95K7bBybASRdPsNgMjTBqBCpTqJpC2zgzwJ5Q75z
M4Xz1m2FbYpNHI95n9BFr0PWIAit3mDfLgyk8bL7nNXvXMa58bEMKFSRxrFa0vQBDE31kbyZM8II
ktZDDc6uny7NgCM4xq77IMHU2t/KcZ8KbcBUVDCAocz9r1IrP6yW5J+28iVSXSh38mTXd3+oiTqC
LxfZ/hE8dzHVjp7pYUQPUlzQ3mZqXAQ926MrkyuXb5aa8ULXykXpvPpDSfWudaJQkiCi3KNqATys
v1FxHrH0/dMb5gY+I8BBCqVm6/ixI380sc1gxWh//9w0BVcialqhpVGTXTQX3z6kNX+TApPRlX6l
tPgGnwGjjhGz4wXiZ4NUBnCbXyZHRK3TjkEZMyobHUE9yPVKsOMHlGpDIr0X3wD0ZdDO/zGQKy5j
0ou8ivCaiIgv8MWvsipBUVg3I8nNsuL2oolD0oI4uFJd3P0G99QY5wAAsfZbK12QVrkgyOh1KRp3
PHMv5S3+L2N+7g17TVVZzFdGcxGmZybaYVkxaXEAJlPLdDTyf/vGq6kZbw4NXL99xK7LVpEuk4Dy
sENQpX9QWrogHQvUCTsZQl2MaJZehsuujETG5IJzSeNMgGDR6Zgtk6sn712OpH7MiM3ovx6wLscY
n9bMV0/vp9vyWBK4YJ9gwCMl/AnFPYdwTYQ+zLaMdirFQCcPxKQOlG/vIeuamAu5IJ/LMoeygM+S
4cTulX6/CiQ4F4LOn73ic7bVHvuPQxLsXZqWb8SJde8bhGwO5mwGFMCaJaEnjR+IGi07vLIkn/2j
sS2oZBoijy9Rvaqm16XAjGupHl498kffgGlz+RqqbM/XZhQDrFEQlSNeMZSMiJwppByG3eY35soA
GotHc/sMwjGrLFv2AGaOSyQ9Jg9zFNy0xF4WqtRs5xGsXehdLpN9gVZIdmnflmLohBDFNdQn2xhH
Di7QjLkOT0Ca06A8wGk6VH98NxwLUZpDxPjfpQpmhRkBgPVq8JOLR3av2gfeo2EpDtTSaO69+eO0
FbZDrHsBrNl6C+Y1xUYdnfgDDHaF0PVQsY2PhvkxhAmA9TvTqCFefvkudQFPdaLsBLddz2sNwkAO
SJPtgFe4MO05N5ZZYq6a5qK3tN/V/Ep39cGQiHlE9hu2TJmHORkrDG/qiVSnbN7zCbGssuXo9L57
BH8YmB9s5k7EIC1HHRwmSRbgrW8fhjY36OQH+zDbgvUUFlVERgitrt6M7nMUpZns+HdpaApPORBE
KxiIT573DLBNb06zXY1++ixTUj3utzq65/cxwq4dBQKqsRjvDJP5mVPfnsrDfZTddKZrKOJMl1I5
X7nQM6zJovNjvjn0CNFpeCkbAInt1TP/WcXuz1jmBOux4QnXSeurT4MrH5hbmh4Po4QWiZW8k6Rm
/mr8L0IrCS1lripUcBRr/B2ZhxP8HCfTwr9/RaZZQSnyxrv03hFqX23s7WuJLzoLdfjObHXn8RiN
ahYTeg/u0vXfSvui0xNCpHwKCWAzf0l5rnvEX8Z5RT+vV8wpYGG6OQq79XhmXJxf96+fGaHkQU/0
0I1gL0FAh6uagz6Cg1uOi43gK4KrcolXVI5YWVgqp+WuzfuMcOc64AyfCd7bmS04OIVOUu3l+pZb
byk0zkh2gx6zE5ETFRJemay3z58yk6pQe0O9PMSB4T+wICZRStXReDqEgvOlnEtjrua6lHj7lJ8A
11htu9cDrclhqlY7vkroHMbN7RIQB/7YZ8uC0C4PfNmdVfNOh5h4Y1XdqHlkMzXKGsFVir7XjZUj
usDVcE6fhfMc/o3Zj4p4Kbbi2AWS763BBHRmDg3opJsKs9MYoLkDO08tpV9R9kL237AqA3Fwmq4a
EPs4qDU7bz/IUbazX4veZMasAf5b364yc32lQvDsJ5ASAq6BoQIN8YXvDCBGQjiqjBhlHdZfOd0P
w1hCGN2hQkctXWUBA62Q05rOMNoiJYCLKgd+j1DY3hNB9Uw7OoNdAXnPWlSiqznRZ68ojWssD76a
KYuFAM0p67P9ubX5skGwuUF/KX84VxlqcM2eDb153Ki/Un+32bV8H3PiMOGTB1AEROBiMqAIZ3Hm
KEVM6PWuQD3+2j3hNirHU+QcymHQgQbf1EekNWUqAPIud39PyF0P82ZRcc1zSAGSiKPbNwngaQsd
0YWVrgqCnj1ZY91xiEziB/6Q5wI84ybx5NT8pw0U3uBQ5RBEXlM7Nf3OXBETpSC1cABGl7CNxAQ9
q+7qvP4l3s7mZ58qBYrvqhOoFHu6pxFxeYzAl8bzdh/UeHuLnkXod2ebStG4BgAoFXEGrsIrkV+F
0EBPx+LWmId0B7Dd1FGtshWhsqyruyI69ZWowxEswlQjEsRYgUNwNpQ7c46w22K80/cSeaQe8Kya
74gnx73RXUWK1c12MMFmIMcIGwPhFyWS0BJRY5YvzDeIGeST2Yscev5i060yvHU3JbawPpTqpefO
Km6QUVbrmXz+oXV8HmxF4ANRAZaS1jDmKPiIun3Vejpjfcx7fRwC83XFuyPovpx2YH6USW+iKo7P
ORzy8G3YWbOXz7ubKcnyc28AoGJDzI+dBiHYwLuwez6NRWs=
`protect end_protected
