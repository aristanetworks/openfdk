--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
l34Nb+2zFgsx9/2tjBP4LOoGskdFfsy0ASyJSMEuaxDFOzFmO1QOPkhu8iYLmjUZVVAPPj7IFJac
JGd7qcoTcWmnAL6kXXv5U9axGSVI0zsguueJmriy/f9OSKgY4OsRQpmkUhLSLL7677+AiSpg2XHE
Y+YW9r276YHA0b9EQVzgsmmg/BzAikMbb8M0B7Z1z/T51DG+RaNjDExfCzuZSNgtHiJSCciz0VlK
CehY2Zw4PCdWUxstsMPP9R5zTgZhNJQf8rTiCXRSMOEM9vOITi9YPE0lfuvfqApM+3+pa3irwrbY
CZ42ruEMEpI+IKooTuwtwym74isKlht9yp2yUw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="THXnjK4qPmPgNvh+A9VsadJkG/I9Wx1XNYaMET5lLj4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
DbmSKlcmO9fuB5E6LyFWG8sJJBMWQxfuzmeQKhyPHWhKlTAUXrlKbKSiQ/xXAiSeR+bdGJpWatpC
fcN3xbHi6//x2a3wEyyLkYpyMloes0GUcl38IMxKq57VoXn1DwlfvaBMGgeVjD8h9lY1zYe8MVPp
q4rLrwBL1LA2ZJ0UaEroe3+qbKCW28boZLuB3lZa7Eb6TRFVp/3GpBuWcpcjX9FeoMyxtQ852u5l
IzDCr7Aujm/0bK2W8dT3j0TU8XMjdHbeCRyjJ8yz7VlPFEqFYX2JtkXJEITHWMsdM3VB1exWQZC1
EXOjqgDriEmgPjTltDdpbsoEuAGVV13wpQ1QKg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="RQLe4LmigZ7DTZB/pckaDiAp4aICstLXjXL1OfAOfO4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10048)
`protect data_block
MQLWZcAqvIAs1O9DCQIRX06LDTOmAcuelnP5g8UQNv2he8RkndHSybobLP+R3oMxQAtSO4WlssBk
PLkyZ77y6JG3y//OlDqh3S/qzU0fudYeEf9R0wDTucimazz2BaSA/k2ihOnHSoXi/qcw1qS7ZaZo
VP/t5boz/dq++hWBb50E7mMAMm4u3XaSUOsc4+byF8tVmL1ojrAOPOuwOrjtcP13Hd2QIfe7ZL0G
uLgJ5MTekuDs0/j9oclF/nPebKjItX23e2q5BlbpJa6tfDZrZKAFZsYkYb0PCpvy1ajKp8b+Gkh2
bPyRLkGcrpnDiev2JDFJg5McVPbdnfCAcpZWMp9TK885cO6eYK0a5uJjCGg8Dx2u8uXFS1U1ne7d
rU8mQ+lCneZENNej3gTtyQdSSr7dysMETd8F1IsQErDYYM64b80OXLyv41wSMVSo4RV9JxlG+0Uc
td96l8/g49vq3Yuy1ohHyeYC5LhuXvLw/cJGdzAzidJtg11Y0AQm38slW3tRzpbr2B3fRxcCZpuj
8eFoTI/pVHTG7mypl8pSisyP+Na4RdySxRFgHmcJ3XC6qbfhrNyt+Z5e1NxfCoSlJq+5fuR9GFMI
8MkFBBTFmhsAzbYSQD36IizzCPwQ1vLZufhDZtUvBRxatzSwxLEtYx2yfTmYjo0+yAo88ibtM4/g
6g0+mjwCWXGtsBZB4Q9whDRXcA1DF5xA5MkyRHmeIBagL28ZsGgHYNzRPvxE+R/IBtyWlB3lv+h3
vxYDodIhlSDTtMpdVhqdb7gi/w4RuLtyImO53/IiG+espKQZ24GbbOcKLPYTo8RTTFCGo+NUt4Rl
wp08oWkfPP5iEI401LGulM7YKqYGW2SGsDYFOHfaAQvVAEIuHcU78Y17GU2jResv//3O95fual3+
p4TZezg6VUVQPFybP37/F8YaFtNMu1g7KQ+d7ijTF+UMPmjGfS+WzuKaeESnT18Imba7P+Dfrg1v
R0XQ8npI6mSZDtToaq9hVLA7FdVzAUVQlNRsB/Lq19iuQdoQJSntubp/PC77LGOIJdBgZK1h1Exm
4c44Ru2zYU4wbSrHkapyOuzVK4Ge51nWL9Zn5GXFk2HqXu+wfeKlH2jRF9VoE+vf0xEGuNSqeWsm
NoWciiizgHPN5Hl83szq2tl97uV8v59OWfeu3PZ1ryFKWfHBdH2+8bZMW/yzK0+xwD8fcFsjsglc
egDYNe8IxGpr3i9i4pCCWincQqZgziAFmZWVKIXIf4TqC1pohLIX3cLmzV4o9rp1GOfvTWiMAVbR
q6LrGUni6ljDsgKtpIUgSxEgQeL1FKnZXByeMNI6D3/Lh4Cf4trwnhbZxiXiXfRnhBqL1fBd+E6h
O5LnY/Gh7xb6aAhhYjWT5TKYJb9UnGK1Ra7YeFhEQ4MgVo/iTJNOPHzVOUQTFizHloosMsLFbH5o
cKgJrnExYv20cvDM17W0F09Cna99xsghwm3DwZXXthorArE5KLG9klfq9nfoTdClg5xrbMqrBFNq
HXwwI1veI13fRhg9efTKgM02BId7atgYFXn6+o5n9fS3xkodUfUVvxg0hP8Z6dp9ft/bR/iaIysZ
CQlPDCctcOiBhqrR5xY5FX6H4VdmziyN7eBwA/KBwEvmsCxtkUe+1eyg5Smn+K+aU9RupQWWTB9X
JkE8vtFypa9CrD+CqafL1iBA3C04meRWSshRvZ8aXb8Uiz6K7kSSF1fUPoV5Ngs/hz9AzxnB3vHh
ptlo/YJBb9kGxlESffm6r/eO1Tv76xuxTR7RCbNFNcq84MHYhERD5UUTx+vrPWh3TBnVUiuNjlIH
DR0zzKBGXCC97xlqvkiDByDuOoR86Pt+A0aMZaymMScxsmQGf/2VuzihL6V5yPcYSrJnRJHypj6m
d2Ea3DQCadbe0Idg1OlKAWer+YkvYEWXa+xFX7qHZjRqQ3HaKNQ4k0dWyjLDdol8CboX+TFVvrUO
qHqGsjKsepz9yJX9IMlKbUCi5PIkDUjY6enggsdUJBl4CxveqS6nHVTANVdT0R58MO+gB6DbW7iw
5InUOa/4/7PAqzE7NnZ5KvEJQGK+GMVFrpos8pBUHfGnwrNLjDOQRmZXM+GoAiOVre3HEmAsG5k6
ELNaSQN4w0ypWY7bMiiVonUzk8aIbOmGm4hOSpGB74r5RIkYbbxwYae6Ym36i0S+j7JZ4f8Am/vw
0nq/KynLaKoA5BnsXmGWMWpnw+ge4pNjrfu0VqMh43UoZUCtVtB5x/RLZ4H6P/Xwd1XOoOAql2M+
Jy/no9iaEzcmLF7j32YV91MbCAbDI2bRiiw73t5U19MwvT7wmpXj1tz7aP131uP4sp7tuDRQfAJK
fP2+pM6OW/YW0+fBuZzZNEV/e7hish6bbFhlPILb4V/t7LuZmGSImc6FtlHVqPCHKSO5cGEcUGzM
+lHsf1UZ4zyGemVsA4O2YIR55KmJozvHvlp57T4OefPweaOiP1d9DFrmlJBQBqbgW9VSjOa/qs6z
1N4pe0WYSl1I61KbfD/iiO1BcxbaiOnHhJzY6aX5UVjw30nnNFGo4CxfIoLKOGPhKfLTJ+NGE3fm
wNwfc1cBsri4oKP1OHHdhyoX7smIZfK0mMfyRzTquWmF38qHhc/Es5i00mDXCfjSWRzJDh1gOtiL
k2iyFyo55i/0eMGQ2ijjnbU3sQDw5XeAnImjFtocoeYmV+dmKsqLCB+9Iku2VoBuuasGFqy0F7oY
hSIRlRyX2uIZlftoiFIFIBZ6KlnyYakvPM4j1iDIbmkPMTNJMFTYH7iRSUGffukzHk7kfScHoQGy
HJrOaymth+/fElJhGllF6zA1SzYlz76IDuCdRzvJLAhbKCUwk9wr9EORqry0KFlsDfs9DODW0kZX
c/zIMfLcef8pH2r5sDjv8TrvI6levkTXVBKFGcvYD3Fptcdcw+XPeih57A37yu8U7cj7ZLqupdnD
8b8UPXPvQ9YixKIq6c17fgj3QHtfPDuJ6zZo6rPPxeL45MAPiTXQpfFxtl9gpQ9jCBaaVtFT87J7
bnl7uLok+I3fdhtubib/qetq9lzHP+7U+PrVS2BSpVL6TkMLaGUzuXBVRNGm6avzYYGaet+hJxfQ
v2hPvtqK9gS08TuyptgJTetIksnYgJfEwArelovji2mMrNTAg+1H1zw8SbNzF9hXQfPggRuBibcY
zoBJJSlLNi68S9qf2/l1WHmT3klAndSsLm4LPafoEog9Gm0r3NsQUPueGcsJOMmXjYYW+bi3dYtw
Y4E4GtAFOVOxfQCHSgBz2y0huGvjwEdmINtSGBobaroHyU7CLhfaX/RegnWBqei/dl1GLdJMwr0y
Vw6htGBRMnPp8bbcbn3aS3rKCYmFz1N15qzBM9aXPipaXus0ROdYk3mN1i06+rvUi3rrxb37T7EA
cMFvPA/75b8RCOWMKJsTMvo2Ju1X0TRyFo95Bdz457i2tibfWPThz1SMHbSs08/80WtCmJGD44MJ
wpIpdnU3ECLI8HmHFo9KMpJxiZ1R6LEQw/cdiq0nKXLs/GBqXvhaWSyo8FMOWW4kZlZx5RxRqmEN
mvXRd77cUlvhnI6pEd0XYP4nHdOxE6MkJvaDmvv8heegg1n4PQcgpSN9c0cHMeRdiBvg3sMUefCk
7PozE6M5HXSfgUu2CQvhREgVoIGU3VaQKdjq5s/rhqoNDZrims43CqoIVpfYLet4ON7aZeaPOWZ6
4KPzJfjT5T2jO22YaZZ6K20z/C6LKCiD+ZEOhBwdu5Q4cKrpRyux1zVhkINaJvdVndK4MsIkmSjD
7hUWmzYdwH69ncH2C4LHTNtvVZY9u/92R0tQ2os0h1100dZuOdu1bDCEfmUEWhdnQlbIFHS+sOGS
wmI3FIEAjZTTHZQqwa2NXk9usQLAaQUx3+XzXO4kbSrI1amo+wdkse+KH70I0JYN/mDBOw5471xD
h0gVo6Mu2cUY82VnkJ8k8DOHSylHPW6z45jgB/0AApX2zxBiF/EIXrWC0wDQXcJZ9l9pbe+zAZb3
jrptTzLuJjCBRZoVWpl2+P6iA4RIW6X3D3D9F03ln7oi+qWWckwsHVbi2oc6ne1UfdEqT6QsS37H
ZdkHpLq8fhCZQ61s797Wq8QweH0fsi2IaogDdMcm8sL5CTYQvJuNOA7oXZfjt05z8BwIbqp4y578
beavcU8FR7/t1XZA209k9uumAbNUwG3hyUMDRnbd7pDn/kWhE3MTjnxBmI/YNG9Y7ibSebg42bXV
dt+QNS5liIh5ZSehm2ADg6evn1ULAVxtbZlvpQqRXBXg/fYB3riUCmQcWKDxZah7pAhMJkF7WqbI
Uj4CCmsdz9iSCEdgGB+Z7buMU9/FekVwDoL5LsDqVk0IhlcFtN7VrKzj8JS5rHM8fR4Bi8XrHwg4
8lAoWJO588efMQRNBowXQpM7oYmBQF4p9trznJbdJTgQmiizbIRiySU65oVSjTn7JN0D0OLBpSb2
TPfMhX7B9+HXYv9kQK81qkZN7KMU0VTzVfhlL6SdHq4KWO3UKqhOzov+0GP7YRavtrEZW0vqLiaI
L2TEfhAl4MbGXxVV9nQ3qcFsMfRsdHCEYwFDPzQIN2NxtvhO13qhVadALnqZKi6CrLlNacx2Nfnr
iJ2ePTgLbdHralh/PYjPUTZzK1mlTf0SRSoXJd1+BiY/h9uIHFVDXLtzkRME7esTAkBzI4QQxEz9
fau1VKdTx6JGlJrmPOpnC9YJjVG3PNWTcIwFcZDmVhTFTRvTnwWmxCUb19jwPiQQnG4WyufoMzmv
HkYF/pGG5ZDvsBVIJLxfu7DayMxztKRf2QG4y1Zx9VuCvL+S/16/E2clYh+oRl7Kr0yTwtfubWWb
fxdUF+VlPxWTDpcHH30tHTPjvtN5GWaxhRwaDJvxxbUeZAQpBe9vWfnK3a7OMVyFFmAjBtwpeyPN
vq1rZrvhpEwdyWtcW8q6uS1otbtbgqRKv38s6g/ZmqCLjXieKg4GtFhyUmt7Y60e8OW8/6rthy/R
+VYrQ0X0r2cEQqp3X/fBEF9289aUCK+PQlDJZN4aEWItccF/Wwr2GIVDgUwNsJZ9mCR5kmi3ubyT
7VjXdU6i611PJ3hrcgvaF4sdlyargvMDoItaKWNo+88Po3yaVwEpEt5Ynv9snzyavzHS/xU1aU3O
JdAaOl2VyELVHnPL5VCXu5aHC9xGeLx3+AkhRHBegBq0O6lnfYm0pR+iPY/FUs5wImBRTyU90dRb
7HiihUn4PHtISYxVUgFV4996Hsq7yGU2lr4harpfqiUZixBHew2KANd/nEl/+twhNivx4uUmvqjG
U8bZ4BkEZBL1nrTRPB2IyW3dfk3cXkWzamjzafwXPTNrYkVJba4h8HXWiORvi22TVOA8q5/Piiy8
00Bc7UE6b6l34KVuQQ62NH3bHE49BU11sKFaPeEuEToNzb4E+eGxDlreKiZhi+oPIsmFDH8HOOsj
xndOK12HQyA8ZkYc4dj8mW9ivm27qt6F31ITgTgZkmv/3I6yMPqvhoHQo2VvolD0yIMSDsprf8zt
s4wPbsEeaE6R9YKQ3HYFGvVpTSahZbOhx7Q+KUt6aSfA8+a3CiQmS1kPU4NpZ48KLVOEw6FmS4Hi
ADHAJojxHfEMUrQ1vedDIDOY31HQWfE/3nCAZk0WKHU/5R2WvObj3fGAWJFbdtEJH6QPiz3CYpw7
NhdHbdUYAGmJlAWob24lN1DHM6OMz8hY7GxMK9jAE7/bV9vMU6J4KPPuo3cyggGMAypmjY2U7GDR
6JTMzgf7lBZWNKOttrUtKwKM0gcdpnkyXDnhBzpJorgNUn6grqmqrqpgElL0o7ljnJBeXDUT6ikC
mrQNo6whEXJk3dM50ASzp4MkOuA8GKY7vVLd9M4x7YYxxaghBmvhdcb/9txAAWNUlITg8LpzjNFg
CervjnPIDeuHwkNzJgptGsGtsoMk+xjX2XekYLgqYVitASwa73NA8F3fd+QykHSjb7uhoIYFSoss
bG+QQpYMiO+JfUVmmYdiZeSMLJlJ6GSEDbRCoHOnHmAs7VI1HUCs7zsua/fhJzfT80zL0OeuboUn
FIrc/Z5V/AI7QB0TRq4ELvXWjK9e9yJ2OzoarAGJ4PtEBPDocv4uOziIuU27TwZ4jRjT58FrqPBw
DuAMKZ01uizQRLI8PDAxLeYhg2V/pBwKXCrlyGNmKG9vBhXB+4xjaDOng5TQS0nBZHQXydqK1Yxx
aThRxdcN1gb/E8zY04JALvTjs8h9s5I8V8R0f0qjxfeLC67w2hlNxFL3Fu2OJUI81G+fNAePUIUo
+YUfCAk1FJj92wvdmagHTw/nlrNFF/eQhbDdJVY6M4r8iS98g+t9hRywfTVcsw5z1oyisidFTdKg
Z9fkITFrtUrO6UPpR6EA2SlzK7shtWldzYFJCNpOVR69zLRozqQx90z+tttFxNqSqVSXqIj4lgKq
AX+L3I6q0jvLqKK56CVXFVVmYYe8SbQHsIFPDYRyBOcbUV7deiNJ3X4/xREqzqSdyI5cpT0LZtur
E5lDqnuxuoS5zPSnAnVKaxwm6CcAX9ihIUV746p8Lf3GHKkg+8UkO9JGbWnsTDktYdlhDvhJJu+T
byxWKdiJep88Mcv/Xgk/s7lmtllk9ofi8MXoUGS1nXuFktYlUg1caI+3QR8Dg1xDUcoBT+bQYyU2
3Oa9zDBf364EFvk0jWH6uTAIWPzLbhOV1JjlcpRUB1R7tjCNK8SCU1WUGttNd5KfqKVBCG3F8H7A
RYXfABaHu5oPAEUuLj6vUBzCZVC99uI2MIs3TPkYgI4Ws9J671VuDcqnyqXWJf2rnlZ0cL+BuCpI
tDTkCdFpRBS3hvRFLHVLOAlB59sOuB0u9vFGBgMYiD+FDdvJIvfJJAZbx6GTNnDUTTkVhNIkxfxG
JsnJUXOdRnEEvdUDcM61TmfFEwWwJUMdKA6trXWO4Ur3YW/eLpnGpqc7IZPAObd7nQWodvLPCnap
BzLNr8teMr7strE6ScPiEs0WoPWSF8fgIkMVPysPy4crfacwSCCxWMNiXGuHVm9Oj2gEx1bf5SVu
V29SGOHjZ0+Qo2leJh39EhLUsDQkKFPADCo0XoSP7ZoQAomOQrNwb7m9lFSKEza/lDACEK34qSUM
3pZjLJW91CXWCZJjjO9riAWSSvJa8yvJk5Ns0iLAecPz7nmor2cEZRfat1kigSiZxLOKvMN6f1tT
fRTR70JXGVmDUKLOnJs/U6TnO6UwleewGrLCVpxIB8SyWzENhi0MwhotwrKcIYqlmtsQAXyBiLIp
/RzNtPQnhij9DU06sjh/sErjrAXReNlfNvCVd8Ayv4hJyMCU7keDwekcyCxlq3YyMKa/wBeFxEFd
JxCgwVxSSfjz6HHVAdukyE61UgBG4fGbAn2rBt2wuqyKn3/H8KahNCeBviqukOpxShBfyv6z7oRj
zLPLoO9Q7GGOBKhZl2gGczILBok2FlJycIqo5CN2e5gEVapM2E3A/oFa9aycLMxBalvrKVZp44Pj
5aTsD0PqQNfniH+A+jX0E9EREl8lvLFqRvNypWZ8EBPjzPF6UGabaWL5f7fuMf4Haq1c7UkXv6ST
VavHZRxgfVJW190tOgEgM929mbgbJh7FPvTjxWDa2LEas68aQqgmfKe9ejXqbJB7wVQ39OejSrFE
g4LENY9oQokvsTEYGtqAU3sID2rBuclIXBPRD6WUYmUydXDDHROHGw5whXWgV3CeaveaxUMezpxe
4YQ29I+JQOrRh3bNVrNbD48QF3Xh1wq9H2I3B2eJkJUMgKh5feIODV5EPyPcFhGW6cL/+UwOetFr
8NqwZzykpwggGQpH0qlfrJwHbydnoPz3vmI36/cXAPaIAQ2Ox5lkmZcwiqNtd3L+BGJg6HZ0Mo6J
2DHuf199vmMlkfZo37ACMa7xMoAVvtGSpE8L5pzHj8OYLZrLi/Ojgb5qJxpgC+hXXHxWd5i4J9IE
MyECldg86NHNI27BQSEe5gtuhJgB/j/s1/uuELV2y5KvVEwFFhgrciIcKhOtON5BWU8czQxiXNuz
3MUzYYrKld6pRtoYSP9sVVbntg28ypmwuEkt+2Xehah+g1fPDkNbb9KqYy0QD3cGuHqp9SlDLOgB
aVO0ueaSw//QkjOwrpXvZVESwzS0Py5pEaXa1IfcNu3IvI6dmp+HhQFtVjCO6bG+MxC0DEfltf2n
GUTArl51W58Anmh2QeBWq11kE3PQEYeuevDIbzdXqTVWlhGIu5BoAlQU7BRVhrLxFDbN1nMpFzXj
0kzK/COiViA3fnSI9sg9muckZShzOifpRgdAm5tGLVSFR+Q21De2f6T6Kpw2rgYHVEhm0qM0rxpz
S19i167AGpEFCHpPpFu/qTaxOP1UB13n9fRb0cBIh3il/Hw4BxaE5iXQqsxXKG+X/B+3WJ0cSiYL
gZ+z4a6HsPNXN2K6iKJPgWHAJSLyR1lpvwW5DJ+GeEehhrnqc10CyjIU1uz/nEWeBw2kmIcQGEK6
FADFtT+HkAH9lhIha/74Yf/ocGuWrBoOX5rGAluHti15SesaoDzdvYV71x7KGTCWXT8RusbmymPY
/yIR2TUWjD83ttMBW5UIdR0PbGtVMgbqzYek/JKV4b/B2lv+oowZ2n/kpiPCsM4hk+1jIuJI3p5D
oDGEPpcAEd7vTL+IfkYVE0E+DnhVYH3MhkEkre0lulEi1ycE19cdkIdj7QgQ+T9Uuoeo6Bn3vfHX
lnAWpvGGgX7BFdMHb6+tVrSlQUKwiVMyZ7PKxhLVv7SUzZAL0zKRjfXjsulwZMEXJzkvm63MUr3x
NaqTNREfUOqlP5BwjZCaeSOejXWhQGuUsnsknpDJwMTTSGC5Hz/16LFxkr8cIrlJKUidGyjuH1QC
YznPIOnbi0AQR9MhO7KuCBPxtwv4uJCAnxcKUnOWQkVYWW7mysm4ERM5AfgQEJWN4GJuRleseFCD
lpK9NDCHBYT/da2kkv8BZMXAN/jnARVKVMODJFp0vosnZj7B+6xYb8gapu8BpEA6Zik/TbFdIos+
F/YxnM5H7DV8F5PCdHMHknZ53iCb07IKTC/fLYUytwla40gDighjo7N507js3EExFQ0ZgRBnt4fl
Q7xZd5dmK4TSCV6wW5YAZhyK3fxhfEwwCWGonNkf+U+ul16ndDPSmPnqL+Vebd6Adnq7tAa7NSJe
33acK+23ajgHcmNI8eBxb9PnPijndMXAZeOy9LAiaLdJHMdF9BLu+L7Isp0ywxe6VjvOhZ0anoyi
inRueXoNaRQu9h6HBkU+SDNE/xuH44q4R342eat/rn3sbe0c5Oaa6k/Y1zOL693W/frODCfS4bR2
aTgV07ergdQT3yagsSWtpeKOVfGjL2nPrfZXVm/f0aD13BdGNC3EnaaQ6Jm3AFMqkWFCRDPk09Pf
MEtKljdPpDsvyUYjP1kyvJQ3DzsHpjeeWkGmA9M7wE/CoqTEvuNnrzLQeqwwtmkXoyxkMv4QMOF/
4LLI5t6LUJfJWYdIqZABkBi7bfajCTYCIOh7L5SLhXQeKqp3Zg+ewcsp6SVBIDYeTkHYjlCeFWSx
EiDbZMjdw8bgwof/cbcFu9so6H75lnL5nkY2OL5kdHuqILFpn63EAHa1oIAhXAriEUDsXZkC2DFm
nqqJfG6wIyptT8qzxLtW27NHcixYW8v5eORJsDmlOgMImoRy7x9uGja2rxqsRFiBB1DZ1qVdfx7t
86iZzToKARLjoE8xERWSMicXuaFY7K2a4UZQy4NeUFtHTJJJ0rtbiape4ynnhAiKt32gk/xpdKNu
W/JBDSs6CL26sv6lPPQwUZ70zXPYR2RMaJQAW8BI7sLQcmphOG/uDgBEq9mqqQrDg78MPkYMYe5i
j+t7yDJ54kiarv+p2JisxSDcuFGakDc1TUj78BgcswgossF6RRGPS1nFQ42XZAkr+f0wGLOdj5QB
5piJpFnSK5kLYiuB5V2Jy1c9qAhvyxCd2Sp60kZvqiPve5UM6UiboAy8jzliD7CZM2zpT9KxmZyy
1EtehsQLLB6xFGMy6bBip1hj917NXNJrz0gZjOSAg6QK7uyc3jTMa/om+YuwJODw111hG1gAiMh4
kx9XRjFUiu0wjPoFWO4bXCxouuzS+stFTMzMfwHdUnf7BJGw1DZG4aTF8qoXOreT3HQnt4/FD4ME
PlVg1surLJ+0ldaethFj3Flx4plot9V2/zSva4sy5tcZti6rcomSdZvwhvbrIqHCsZOLdxCZ3efW
5ISl6oWszXqhqciDaBUTcs96Q0pRzIcy5Q4mjRjVzRDq+bLZdUTmBtNY5g3OVaYAPJb0OtKscOYe
awdepR0nCfCbJle6911yB/o/NCgI74UBQaBvVz4fTcstsO11vBlPBmFIbuQzUHrq/6gt24axQF/8
FZuwXsRjjVO2RD5AYQ1a275XhRcKDQ6vOyFXi+1hfatatrz7EZSD30s5dvlf9m0z/piCNiMi5Lwd
g4nRA7lMQCBpPSyTLTtSpDtRZxsOn43rf9Li4L7OUzN+UtTeiUyisbdBO8gYNrcxVzOPcPBhUooy
wIoAF0/ozrbwH292C8HEAY6GbwXuODinLlFw9thim/KI7UeL4/xHettTYgqrKRJqEm5T2c0Zy+Uu
vSC2J5zi7mgSUGvR/C+ExrcgQtIfawQRXRh7srv3IlLjAsa9tAeagLgfmG2/o3UGYAWbNC1ZbGR9
daFVgE+OKct1Jy4puXtC3/m1GBpjKCHhOCEXTYZl4kpWJoFoQK03WaKE5HLJmYXUDpbC169VxZTG
Uw24crUh7J7ab7tVG9aIF83wdnHIEa0dpZ27kcbGgxPkLx5UhpAJp1YrbrbRpTTvBP6PtY4MDUPr
vr3fgCaJ2KjsOY1aH0GuKq1TtiqEqR8H64RtKM1gq7kEIdJkKpztCGn7Njyqfv+MuZYoYQtYe+Wr
W0CEqLpMoecoyRTEgHJL5MUeFEQM/zQPQAKoMbCNsKiZb+r+LgcK8x8j3T9//fyjweMEw7HXqU7b
iNe3GXUbo7zrt7tYHAzhyhrYEN1VbX707Dro2FSn1zDUUIxNudqjGH8BDynmsMCrnrFGWoAKzvhQ
uKMRx9cHLCODf6K5y+vIoh2yfC577pjBc6jT6BMdcD1RTp/gGPTJpWuZq6haaXwFugi5Ru0gZ5KM
WjrehQ3rEZKibhr3Og2+CtacT6s/KiPd+kqX7G3Y6/AirB1VaA3rDdmz+fU+AJrTkP/9K4MIUQSo
qkFK/Obp1A1pwrv9rZCMts67OaVhnbuuiuzNxTbb8iVfaZqxQmeDuRNVFa2eLDd/4UhxfY3588gg
eQsN1XoLp1QLEvIodpJcvaJvaNvW+9LYTNrRqUgA+RBhzdMMPjGlrvecoHNp+tYRQ8AKTbVboj35
XkCAgC851+5IPfOaiIFy/W3JsovhVSnmYFT6CLUY0SOreOEHf+W9JKKbXqXkOovn2i4Mby7dX3mg
A3b05WbQcDNGeYRDjUdJUJ7WPV7ISAVAtvTSrPYCbgXp4FpSemBev57ZPNwbX01pvoCTZQgc1FT8
AXDLLCZzx8AUGNVKYclSTOFnO078OAc9eN9A/zikh9kIr0bzlTG2fEMgujk4tHTl3/+Qf6fs8EJ5
GCDheciscOBgKaIixoiMoGmN+tvnVJSdTVYKlKw4049mRntP/GyO5PF33JzZoByW4xfbjfXmRiwX
fdQPTTZiXU2T77E9mnqBYXxJCtAY2S8GjywfwMAjmjjDKBKLIKyRi83d+A7JniRW19CLhsRxVW9F
XA9MhHx6U7kdrCMWg9M3GLlQGoqHTCX+JhqJHQB6vEZAdkPwovyc/LtMzW86+9MvKJHdUEK9Ynm7
XbXm0Q4zCHgLxN+gJw5bdSeg3VWA5oAk+kjchP7SG3mSZF/MAVpt5T++t0vbWTi1r1zdI+1V6Fof
WKMkDCOb0Hgu06M90G3bPuupTRuOe7T7QujEdHH8IAA08HmoVZAUVOGfA3u8GOPCw2VQIWeqGcHb
SQ/Fe84OW/bw/aPo/+Cu+weO7ECW+OJE3kSudx1qX5Cfb9uIcDOiOdD9bWdokTrzoedryYfK1Cvl
tz67FfcgTNsF+BPiWykslylDsfMX/s0VzSoXZKoLB48VzvK1OFDMo2DIQqVXjcDx9Y+7lsvjVpkU
2fGChUWUuj2Achk8qux36jcFXP8RJESBKvER148RqQyvkwEY9M/ebaEEtiS0scWfWm/sr87imA5w
QA8NpgX4fyF9BlzKwdiUGi9IGw9IRNwYXFvLzcGF1urefhARUXeMTWuM9yRy0F2QzvpcPZss6Y+c
oJOgSy+fMDaHk0udDtlbT29KNqxFvaXvX6Ws6CFfmAVDDQJhDfYrKTB74c4JQZ/RTKyOohTaGkb3
A/Qht4RS4n0FL/znqrIF3qmUlJJEyet7jcIYzYtb2T/Pzo70Mvxdmvqw9glt5AuJjjDAAuVXT6rF
QEZsPIjs2wm+S2rJjiG7MNNpAIYpo9IvSJIeZCztEqlqrHVgRikHQ/JyyJUNOTb3PYrqmgYCZ0U3
4vnOiOqvDGJtYHiw/3Uwi0Ywli3pjIED2DX91ejn1sJy8Q8C6RU4/2JmFleNJG01FWSMdjGQ1O8n
kiushHkootbqYntPyP7bkbhAGa9f45GvR1LpPOpr8MLsi7WdmTKo2KbhqKPEhXBRR9LUjpBDkKuK
cXMiVN7+CWtxBJ0YXvlcCHc0zhhPYuhq5mw2vL/6lI8d8kY/IvXu9zHhCjHbyY9qLKR0qublzX8Y
eSCL7dPwT7tL2D2sCr+Ig5z3KqwDTy6+yr2onCI/3BEFp824wp/L2JtnNXRhDxEKjdEew1+FqFGp
U1Ktj3QFHuyNUc3MfYvvgEMrV0O39+SIZobzgG3Y9VvCQLNmF4NjWoF7qHDx6YPb915KDsSopBTj
ub9bVeaaWFywU1wwpK5QtZxBmRpk7fwW8tc9nTFGJcFXenAA17Nhe72k5OGat7UQx2H0/FpaHNKb
53M1xGANDSJBGNdisyJFqTLYyVk6O4qUi9KHELAkA0y9BGpF829TsGrStNICdFTrX6K8q235K6rv
3EdH0Typ2eGQc+I1OatEAjysWOQPp7ok6LLpxd/yBQRs3q/0/YfjR4i7qZZzi4UDi1O3lYCt3yEd
puZoJSfS8vzfEn7de7wc7YEP7SlQQDzQB83CECsDjph9Oz5114FzRam0C4IytQKLbw1neHmE5hUB
MTpb9arIFxJJj3MZXkEnrbkRbJoEoTtoatrtGZgVe12DfPvJnXRI144B8jGkYAYmg/YP2No5W724
/Was6hrmQ1EAXbkLZOJIZDC1PucKvNx5Zql56IKsEunXPxCn2B5jX031kBtsXQ+EDsQKS4a1PNH+
9+HBGmCecC0jTrPlfAyZyg==
`protect end_protected
