--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
X67NoaTX+OQ9Qp7ziH+L0kxpIRpUyfI+KdWBnl4oVqaNg2+/4tQV15jOa9ra/+yS+MzFc7mEmHNS
2nwgGJmRFIKQUP40ejdgPW7QZEqzzuV+52yyJgOZ6EHmzbg84PJh97ftIjS3piWgVtY3+MTGcit7
lQvizPv40U6sDhXGFQ1x9K7aPSTupflkLgcMrKiTXPEsFiMo9cIMvacrw/fDl2bnermxM5q4dWpK
PyBlG+n30juwLHzJ6FOAxKzaQpRlbiNpbisW0v55L7T0jpvvOR/NE/cYS99ITmCUJ0t6ucp0QfTn
+xlz4QLJ0QAvJMDnkQQdAjDcm6oqJXV3xScQYg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="2mkrbTWKpm8tOME3+o5L9d5yv6Sg8DnYs/mC+yzb+XM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
JzxHCClw2m3RJIFtYqLduUZo1XxKaOXU92cj34lHZLm3Pt5+jTKhZIOZbf1+LEFpCZ88Opzotznc
THw1EZkhUSYLH+aDsEW8S1WJjbR1DuulbXeld3frf8BSweWgjniR07nmBKu1p/TeOurcS2hhQbU7
82XMVHA22f1dSTprioi56AikuW9CBG73XT0aYUq7sh4Qx7JCkQEFLzjwR6kNyOvyGEYfj9s7UtI4
P0CuqnbNUn37+gKEgafXr0p8SzuN2O964PoxUNLLAhT+9uXyJZlMl62lHZgMTVO1iDO3k07afLNq
mBl2VEC2YSEYe3/k5tGGBzzoFnvsBOG/Y7mp8w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="SNfoBiZDG3FBGXhrSDHKEctm2BB590uanftKjDoAg88="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6624)
`protect data_block
bL8XikJa7GjwbZI39w1vOcGfjRI13z7YVIrVRBoJ7f/taBn0+bgWDjXBkdTqWoi1Fncwc43HcjOX
6yB6MfNMhvvm+ZEexFGyGiv+NrRZAT4KAd+yxP1qjkA+mMvYUk220SIxoO3rENezutY9D20bCA1a
yxkQxL9bIMRXAqsAikGks4CsLV0ta4NPEEBLsOsFb+NVKlyn0ApBh1oAVqGM0m22g/li6q6RH8xy
XVn28q+Y9ERBQo0Xwnwpxf+j0XD8QFvYp5je4PLJyRcozHuHEag4RKSFOHGPvHfOmNMWk80TRUg2
YeaYCAjaA3DPrHVy7G86y8/IjHTwVJkrkwkKxvNJpSMnn1ehnvXA6OrLlxY8rPQKG/ziRqezTJSM
XJ3Xksl+Hsl72LhYm0RdPKLxpKUpzfktjLv4XTlv61Z+sEdYvWbEqAULYYHQxZo17xA5EsZXGoqt
Ww77jbxk08a+VvVPpDuJxN5E5wHUsw7U6/AwycQ+G7HqZamZbT+rlPyd3prwyes19l1+NPgDptJf
j5ECtooyenMhkdzCELm84rKARrek6m2RGIEkQXC2DrsjJTrXkNdYY0TUHmjcycNDtxAuX+wUyG21
1+ZUJsfJzt5g45m1Nv/oW3usFdp0toi5+nUuidFMKAIuNSlTE6+X1igRizNU7N88tANR3LG6DrHZ
lS11pY9CUrD1Y6m5UbbxnAL8KGL/fgamq19ZQh+IiaBCbm9QleOMP88/WFQv/mcRdNzVaH+IdqWu
NtXQXIPFvZoiZ9OmFZZqTOhXwQ7zxi134OhKIkCnReOsRkEkB8ZSRw9r3b0RuzV6ddY7RC2YTozH
z9CfnU6JOXiwIfJzMqxBjh+p0DD3+TreYDBSSDJqUCdbCilcE2kVglvPS3U3jRMXUyYY82w9EmKn
eet7xU2lGaf+JGi9X6LReStrZtNXU1PbHUXP9IZarSWAuSvdhmxdrd/HIzKsgmWxBJjIj9aTaSQ1
BrGlA/rpCFpplYRJJ9AE5747KMOkvNsHDS8nL5vkQD9pZyKRZP/BjiXv90W+p3KqHVQ85vEUHze2
cjkMh+I8C6Ka02DPglZ++UIZ7X7vQm6WxQbxpmAzNbMahAsRyigJaA3RO9jP3LpYLfphg8ggUfrt
dabYkpAAnAn4Nbwm0gRkns8sD9dnfWQDLfyUVv6ldJ/4ldS9K79LmONKuN4YUK/4/iqd0ZZWl3i3
wfQR7A/uRtBJJCg9rwjYMp95D9scy/jrHHjnNBbXXyyzwAmS8PT7ucYLLBxygRA4eEcqayTeYP6w
Hw1tjKxeAoXWe4shXCIOFaXLgTzZ1NoIKwyl4PDkSMubbCQi481MWXKURbj9v9ZxI/nA6Av99ZiB
N+O0H4o4P8jdP/hG6pwW4lQh4fEW6wk4txmdpYxHAYj17kDC4pPqLHdWSNUQIS425fNVY+6nwyR5
QwvYAitVxeI2FRWEaqxGgFhxB60K+GRjgag0Rqlu3H/10Y4/MdhXNfUQtjXCIT6Va8EP98Jtkcq0
5lyvbIj3IaZ0+PHbk/p+RaHx0RaNsl9kkWooGrq0fBDZbiFvXacRrSvZOQE/CzUwbWfxixv0L9nV
9fAITaRFEB6oSfKYVxpbb6psfEEyGBMlSSoSTaWHax1U5fQAjrUo4s8IvkYQu4fwPZOKuUc9gI3J
Gf4034DISj6T0w4TcR7mgOwwzwnFAuTFOcutU3BQ3QLix5PJI3YDmsTKrZ/zlnpjp+xi0ah8bjHS
kp1FahvU8RJbYzamfjtWDyQYgny5HBhJJwWFbOxxYpk7CWp+iaxlK95iWbXUP3oieWE64ROI7REN
85gtwhIJ2mo1SWaT4npz4VQrNBp2xgnQOTWd35ijaa6peLiHHq8Z7hYXIUKxQW+Qyf07vYuEg0/+
METyyUHIAIdVDemj2Rn9Wrudx+gCb3QKzmUN+av/k7LGQAO8FiNZgr65HZk+j4vr1SOSGWv8p9qr
EBqC4i6WmeKTIOcmiHIOI4FZRtiMrLLrNo80qzWgaCSmdRaqCNEIJIIr7A9RW3HhdhS6lSTDwMpg
WuRDE8grsBhTxsWWR8DZ6GAr74O8iAnw3yE9rBWkgVKGnenFO2Jh+ka+0TNUT5mG3bMr2uIZC8qZ
kMLT8Lck4+/igswa/1BSKyBhtONhmppuAXpoC97MuI0pjld4YyWRl79tahMkC0BrnbJDt9OIdWyN
L4Nq7YlaAISRuF7A62y6ilQOMQkcvjrQmQvA3/dDCKIZndLqJn7rExs/rYnazFSwABv/32FIHh8F
mAjgCKxrOBeunJk91QWGhMPfASRzpZMmNdJMi4cbW3BDBJtqxW9RfCxepO6BDbDsS2CFbcsmn0pK
WqXRfzP2d3AaPsmp0LI5CVW5DVpgICwfQw74NPFVL6mAZxdy8LTJXEY7dPeYE1aomLSLpxVtkN2c
Br9GIu6f90t+8szoH2zQtkA/eieVzxu8XrE/NU0KqeeOhz55DM6w4IatDC9WCDvT73iD0FNM//7M
3Q3SAAwivQ4qexI6zwmrxpYViUT8I5XAcz40aGbzKhIUYgVFHm+/VaOYS8qo6KfUZA9W/V2NXQB8
ZSGfOPLeRXeXorRTyvlFha2JNKvk6sXXAxshnuaq+FXhI21wYpB8CqSYJt+anFkciGjIRqdg3x5R
7TTL24yDb3Sy3iHGqxE4+fFmUyP9Hv45OchAcFz1LMqvLdyQAEBNwrIaZC4D3t6NZF7yqi7/EQJv
WcCGwwFnvPJ9qdg7OdsQbeOjlwrddWjEzJcaPfwaM+GEjLHhqOyMUDqh9jsnvFAklRDIFUUft4eO
MqfpFWkTGcLmXqESVVTzMzSaZ54PUJbl8zV52EEPGS15NzBVHqUFeZUAXRT7oOP+eBLnWvA1lKcC
gX5aiL99HAT+aIPbAprUlInAwXvapOgJ1+l7hk5hqp8qSqs+r9FuLZ2yQ0VKEqZzwYvh7Ng6b2DC
CtxTtDQM0toKI1Vym/wvIDxvBEkNEjDZadYYy+0xxIPtnLIzkvKEzf0nv21mff/F2Cop2JkxDAuD
CbLApPOZHdJLBf3BS6gsAD+U2AMZDXHJBrH7PzrxSDXDlPAyBWhKlz12162mma8A9k7oIHz2ZuS/
bSZTo/PhX8SiV6J1+w+Q0hyGcec3gTiipB0t70iGq1Ub51rbWZKwWuFg9wQWlzSxTJZeTR1ArZnb
JhAJG1/wwoQ9oFZCqbtbtHW+0q+yVLbVSBVbKzhUIvdy9xvHudzJJUgnCn+DxKTCg6rHTJk7WR44
fB0tmfspXdjkJaXTX6JCZYpEXW1atLHnNiPbmyjBxoEO/u03tR2ok6ap1G4pHAVFYWmPuXNXiO5D
Aogrx9T3eFR4YtCBA18GrsCZi49vJ8+sU3n7tlzVNpZY0E3L24oEZlakUuAUEdffcjvbn2/x5mpp
qgsw5CPLhm70Psp9x3GK0ey3jWOE8b9YEhQoGyNCcqXbRH1YKOSn+2tbjLYxn+ay93TOeHtYOPUa
sqTX3olp/qCIYoyECEPNCOB8MdFvq+U3fN8np7mejt6NkawdyzLexHd8w719FGHzcSzZjnSKfQQp
1LD8kIqUDgktgKqNMvyO3O9ouqBN4RVpuTaxmgvnr/JwCtlHAG8NXtfkkJ62b/3SZA/5v1x+YfPu
mNTx/BxBxYV3GzUhno3gI7KwQAd7F4/3oG00wTXPVY+nZeTQ01DzUMfmureQUFKdXEuCIXkIyjJD
6PwwYnCh4oDafKoQAScVu9n4tjRhfycX540w8mG0ELkiQlJXI+93zY8DRMis/c4ZRwMVbbqgDHV/
k2y/RP1gAEaITnh9uym8P0EC8cFpuIVMASLrgObQjA26OULpo58R+7O33EOcg356SAdfF9Glqo/d
XO+TxHWA2BfagI4jKCroCmLUvsyOeAtS6Vt5dWKUG2aW7iKHasq8xUZLILLo3pJWwjXsMg2RBhOJ
XmTN3rtyW5R8peMWMEeqG90lVtd8hec3CPtwa5kSqbJ0bpGeBBPSWS1R+or4ek9xNEtw/W+VRgpR
PGWLxvhhtkW4rqnY2H6WbkWxvbG8B97DPil9EEDmKNoe8CsjrUebx/KKIlIasuwOgcTOKxCIGlbv
YJWXBOuCfS0zlIuOGBIGV7KgFqcxTEVbxergSCxbbKkJ7mgPPNKANozW0mEGhh3EhFqDjueN7rUZ
pL9KBMJFhou/7C/6T/Qxq460E/BOkxUWjKmEiQHHMc2hyNU7ETY7ga/nT/3tyZf21qlNTe4GzHlX
SWwtxmqBmmRiL4fmZwQ2EeW54etHvaoWBYLa2OTlLdJuxu2HdnSckFhvwvj/H4PYeHKEUoqspABA
P1kUBmpmfkN6c50LvxYpNUMPLeztRBbUMQuK0gNRH9YOIgGwuKUzF8oQ7gRcFqNNqm672c/O5Qdu
naciN9cLCKzL7UUNxET2mEyvPt9x6Op8wNmjK1l/RTGcSGp2DF04ryFNY75lJah+dyL95ZCngEhH
r9lXoQPaQZmr7Sy38JJr4HiQ9+iTSEJ7MmAnoshNVwrFI44aquD+cK3qTX+4LT0ct6fhjjwcNWkk
OXtaIo1lb9VRrTVmy14LfH3GMUcPPz9AWEXElxkARrmJUw1Q/CACkonZIQ4CAJYMTtGgC2eNz/U/
ZuVe0SU/HVXE/cUT/cxdaWmrJmkXfk5cYuSWi7b56Nf2n/9mkwD391lr4fMdPUwT3/HZvNi/DtqN
dj9mQ+7tz5zVwLeZQotmkbvU0gCQPEnlh2D2mLjMKdLfZbPNeNv4Wsqz7A0nvqdwQRBjCpvBe+Pj
2aNm8tWVtYaH9YVQQZQSnG+CyBWiQ/0XkLW5OHxQI7UbrNLW6CEupotoCUhg3qcSNAzw6ZDUn5RV
uVInI9eXWFK+2cUh2Z8nh8H6GmKaSaTKrkO7OJpPROx/w7q2btHS5AMfr8YPXpnZjJ/2Mehbmpkj
pi5OjmLAsBc4kK8sCgYZMZBFOBM4c658NQNiaz6tNBkgpjpxFP30SRBvPmzEahvQhQjafCJqDexh
08FUdqgPZmtnYHQbazpTGuxe4g4tEn3ies5/3eEQlUr83B1Z76WHjGvgFxMfQO1unT9PpWBSbupU
OMU9rxIJmETxb4phOKQMPshtrl9nN9Rsl0xpkv0EBffUPprTj4SVpiJNYIg27GvDg19212mfSb7q
mwnWeL2UClsO/KdtURyOv5eXSdQ3RZoxIfI9918Pz8bUb4us6MuYNIRSEmKClANvsh7wB9v7otDo
RWfmPtKOC0xNo3ptfIXMAXOrurgC45GXewB92mMi2l5MtB8a+XjSCZ0NgRi3CMe7TTMVg8MJFuhh
lW4lRElYyVFo/PshYrsMiUhutq/m14sxwQCmTGwBc/huHqFQE/501rQrSvST2CbY9P7yEFHb/4KY
R7oowDvJq2MMLkgLfOL7HDLh2+cTaUUuC60pqvYzRI9gy7d2KKV7WTHBDFvjV5hEPBmbeWiOSWaW
3BAC3n+bprHp5MrX5hqrZe410Hxa4dymKCsPCVRxLN9dRv3QFEt5iazMeAt2UcQEBvYZ6dO18CDL
qvKo9mZL3mU/lJS4buqrSX82R+pkWU+JXqaL9lJuO8GgBgAPr7m3IrdMHaBT5eW4krwpwi3NpUrR
cT7515SybXLhPP2XtrQVrLHT8qcKKe5YaIC2zwA80Xzhp0tFfsrhZVDkeulo2JJoVOOrBISavHM5
3NQDG9mIkc/Fnc1zS8oGQEqQPvWAdkQD2f3zA8TevpQkpBMZUrzqn1aPk7Y4Mrbf0BjABoCOIQfl
m1oL7MGGzsrxtN4v+3CaMef3J99IYSOsiy53ELBjH6cloS6tadJpyXaJXjuTYwMMLJq0HfCAzewz
yJjblbA+g7xxo2wd/DrHtyLb0DIzcKuvvpi6UTIra3PK5puftxR9P3yDAOa0QyFTnvd2cZWSt6nP
Gc7VRFFSQc3sAb5lo0+MgjgcOI6kht5/8tJL5HgVUa6CmBeu+kFpq45yZiazi5oIvw37kflMGGwp
Hmd70tiiOIrv9vTAPwQ85OoDNvjXQa6ESosgKYuP7bwGylM6XfTc/8sB2iueCkAbFLTjFaT3Zovz
3ReNF8movUpBVKi3NDeeN65K2nKO9EnL6qyYbWO97YAqbNHLm0z4k1YZazEVSPylR7g2f7r0Bk9k
bjjv9LdAI7WZBuvfBkCvOOjJWRJ3BguKxkpmQ8CtRUkQfY81LSqiX3xAA51rv9pHC6aoix/0kwDy
2zCeqZgonf4K9Bt1fKwuUr5P3TYUbwmHT+1WKzVpogmCJrXN8JNNDKI+4B0v5CMy1R8fudXx24sH
L/7iUhKR28X7fE+6skZXQtARbOyfdRvEj7b/UclkvARDzmQuY2yKuKAgULsV40R1D0niOMxiGjxD
53RMqLCXiORoiHPoG3+OzmfpKz4j7dnVRkNehFUggRT3CRUv/4N1WY0OvduwZICkyOJfdm8uJeeC
mtw9u0Ca5bpJmroBWZqwEMIQXigI8TDTN+8g1hDknhAojgzFVqycM9ml5CR+gOzx9Z6FfvrKnaXQ
YLCusHRF6YRIunnv3Ctk7mQnsLHF4i3muPb+d5bmDRUtQ1fQ5ZHeID4dKMztrCnU0ox6JCns+DRY
tz5qp7BYcCXKR956sWjRnnFhmzwRBTV3DDH1D0uQZvKBXDUWn0XzJALtCR4jNH0z4JRzWW+nU3eX
dh7HCPxGIjnH6q5M3IUm50RBxh5Psm+XslV6SIZRsNh2rW68NG/Qi2D6xQRJ4qycxSMLF017zrz5
V7A9s5CridnK88wbqcEgEQ3xMkyFeBwc2W2dxmfY4uKACcJnTTvMptIn6GLdqkNaQnwfskXO01Vt
14YyDrvYsw0GEdf5iJphxJJb0EAQIpIVXhoWG2X1TWEZgWqeToPFA8dxfXvVdvqlCKatFbIsKCSk
FX25n4LJ8Cz3NQBzcMFTftTtq0CZ/DgvO1hKAmA2s0y9XXQDuHzG+LMAMie6jwqdpInqpE9fVEXF
BgA251Yag01P7fXhLLM3uqwDmElkdNOViLXc0oyTWf4TQZZ9Re9nODHo6A2nctkPSV2hMTciEE9G
u4+LOAHOTAFLGn4vbFqCUSEcEhHcPC6hiMQ5Aqrq9VdU6C65amHcZKLuwy2krCHI3KNd/j82wIXo
nvHqS/xaFrvLPjDcLdo9EQfno9Kx0SmnjGBNLWISYm5o/qEctSbrE843QWJGjotxRLcbeShmfmAV
oHnOyTxbR4gHl/dRQ19T6dYHL9W+1nOPL4RaMhuAg7e+dbodaK6U/YxObhRLefiU20K5xV93rjKk
rvmhkiVKSZdZHelImk19V0wPUApNhCDsyv+v1qx0dDbcKopHFvkE/mH2oBKqrzs+8HXij0BcyOQ+
i0tG2ECFGpgaTOWuJ3lux32bXTFiP0aWhWDiz0s8722jmPAiXv656W3ROrcoXDZCIfHBDF65idEZ
0UO0ufORIYNalJMXO1bsYX8QdLKx7knRbf4kMNZ4tdymMi3i4mX/ARw2Yh0DQt+zAnfJSYWNKGlN
kA1yo7jHzJFTwm74m36vIpnpEJDdbpCvXlWY8wT6W+UNC+jCAPcVAHXnee5JRQsq+TrkYQiAd6f5
mG38o5s5cKl+AP85AUciXVxcvsTcXIykChQIXKzb+Q2da/lGSFHLjT6vUFWSX8QPKkbKbvq/pavm
0F1MU2H8psz0BeS2v6i1KDqzpzxL84S6vX3icFhF6v2H0iA0alHwEtcqC6cg/F/U5lEn/wblp34Z
fis90r5dv8xsJHBLyz+YrKZJPyYfeFHHXDREaIdGZnA4fxsMvsmih4FiXraSmCx2r++2Y2ErWqWg
lG/mWaAdod2DIDIbxIgpqc7r/0516YeqqelRAxlqkY5lDt6HgyzRNwNc0E/zPkxPFRKUG+NhIYne
GKLpikXRpragb2PqgJbXB0+mEs9aggVbRE1JKJdZmrAK1VmIxkjQIeh+qpuvSfOyuz6YgE1fSbzm
FON/6xEog9U2GKZkKyeVM9/q+UvZ07+WgAN2R6VY5aZRCF/rhlL/Z0qJw15BdF8ISUNAsYoCfCfC
LhOLBv3o61auB1UAFNhx3NLSsbosqkCGOxAoQENVf8+CWsojOJ/Kh2U9rK8tjOAfFTWSeuagxyRl
84ZTkutHO25Er+dPPe4UNy6B40HjAp7h2GXjCHIFgjCCvH/Lws9vO968oKnXyr/sHJn2MP7mih+i
Sz10+O3JfAjJFqnB1PNhSxRGDUNu4kG3CP7AJ/ZjGgqI5l7A0nYaxlJxBOQU6FvaZT9nXSGJAzVm
UdflHLJyq0WnJ1PShiTjw6fTIZ5BzPTtPW7MkAeg/GFOokZinkZXaWm8glnKaTCQaCf8LTG7IXPV
b8b8JQuHdyZyZIoBY25TTnyBIuyodhKU1wIH+zR780a/FZ8SvXcLYGpqBEW6hPmY1mkrrCqPHX7v
fUgJcR1r583NOQ2LIJtuNNHD8BgayO27ohqCxPfNZqiKyaumuCz2RzFMACEkRiHf2RP735groyFa
1MlndtqqQIAN6sJZY1kerKtKLaAcNxy0mZ+gz5DGL47aNwGVrRns79LhBirVyF3/R9kOiyMOjL/t
1ri2pO3Tq3k1SDxaN3tTiNAW5hrrpUea/mHUb/YZ2XkRgFMIvdxpBhBAmvdiIJzf2yG0o/+cwmWQ
sxcDlA5GnnhfxOBNJP4/D52S1yMPME3LCxMaoL5bG6nDMpKvs1hTuRUzkpQ8wlyKsGooTl5Rikmd
INIQtlcpgT0Tvn0c26w+vzvEA76sDUPCgtnVAyx+ogg/J7Qn/jAYFqwSSuCFNEnPgU890S+/7u8E
Y27OhuAjLilf/YQQ
`protect end_protected
