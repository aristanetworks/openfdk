--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
IeaT/6jMnLdCl3p/A36jJssqdOxvyLf+SzhQ05fU5UC/nTn7f2dismWQLk+czQdBN1ySA/xXW0Om
jMKBRDsYDtcfP2Yz+XKilhYM6Y4WQxbMdxausIoQlMnkykIi/nq1zktd0pyUoIfmTIQON7NlATYm
a13ZI16wzZw8YFYarkqpkZNqhU6t43UNpxlGWChvAffP7g5gLnBvrAtsmIjBpiIFTj+zOvk3xOGv
5MGACP8tzBgoE9J9e9LeJF6D3WxVyFxyGFNLjlUT35zQ+XL+DGz/Gz0THubz2LnIE1fbGKNcO6tj
LUi0vtDGT9wb3JVbenkB24va2H0LRtCHvokJMQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="1LQFOKUN1bvCZc7vFP75Ol2SIHh3kx9MTss8NMLOB9A="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
Zdy3SPisKV6pkHTpO7F4ptlqJyGQ255J0AyBhQUpKokd9GZUD5j6vZg5VueKROXkKG6sa1ccknC2
Kqhe2AoFKLwLgLaDfgXqJQXFEw1gH92M5ALk2trCAGsAU6Y3qkCZP2B0mp8Y2gQLFZ3X8EUXMNEP
KfiLk3NF+IFdXbLyR9wsMt8K2/ziqCVz68jKhRbaFrSqSGq4uNALtL1FEs7X7HJoFY+8NJddpZIt
0zFHkHyv097qpFzs5zNTLMaODfzIDB53+QEQAHk0ibIWDGFph3Vfa/O2I37ccyV7JxpYbwgoX0Lj
mTTaqsM3Ez14NP/ucL+M3DGVQEnmVTKkvrzIeA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="0luwYW6N84iCGroKwva2eEZUAMyj2Hv3KcFivYvkFyA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5184)
`protect data_block
NQovf6Jp+RlkRiTs7X8VmE1w18qClb8ra7/2dxuerAGFatFSeXFXBBdz8M1mRhCd+g8E2onDpado
Ty813/VDk1bp/3n5GrA8+W9eVSRALr+/THJM8Y/mo2pSsfgj0+QFUO0iU2SXrv51qINlSzt4hkwN
NdPMkWbNSxZ3bHK0PC4ktbSZxx6RrZzvN+NMdLRLSOwaVoq7cLCBfj0JI35rEX+hPnjYRHzPrRQZ
rL8ZJEshIR2R0Tc096j9CrAboJT13UpvSLY1NnwuB6AUMrQb3VqptjYFbP+//USSE2zBd3XYDFya
N4zgEfy8S8Y+a1PE3aqHgQgg9BT2MH3CIlBke78eUqp3W40f4Q+o7UVESZKnCNWLILSzGVebbE1q
U4TYwu4Rv1TkprWk6f3BTww7n6jrk2fiR1JREpwXNbhUvA5BnoGLHeydz1pW8CCm/4ehIls7qLZL
8KSDD/DtWsQKZ4NrUD8+Dr5h7L5GrK5tKgcFMNTLilk5//lCikuJaUy5sFzpHLXmU+YnGZPB9vTx
fXc0d8v0KWs2qRFc7wfUqCrRwGwn0YVm3S+2pZ8obAn/GfGORCnlU3UYK0MkuCF5yIs5RTFEVAlw
gKPLr2KJQFlXgBmdxrjbsEO4A9YlnGfQeGjQM/Ywum4DOPyGjL+b7cCr1zoRHr3IZMjMWqboScQt
MH5qjeWWTGVRq/UTDC2J2vZuZDF4t0icoVlb5NQYMAMLDsWFj3U+GiUP/o5DZZHFu5eKuzf6QhdO
+k1jhu5Ye1oFuGr64t5ZYSR0rCc49WybhpHj+shTQhAkUzzMXupjvgx5s2lZ5nYVwpMKcU9Hv45z
MjlE5FOZa9cL8KCFZLcFAx+oLTmXPMvcoK8yk5uwjqNDn7/0uirS4UVIDfgbnducD59rS3D85W33
ME7YtIyWH8gmkjwK5zQhUiVsH+90v+RtSmFcTdVk0/NWdq/SvjPDdjuNRZsPHWBABi92pfqH7nt3
viy3AnvSXyAG5554VS2XFwb/TpG6kinUdBL0itXBS1zvfyRCt66G4jMOrGYLDn4NeFTI15W3Ri8c
iWenT6W4foAVhRpHRSk49mens6t0eCwJ69JV+SSTYww1A1mRtdImV3dMEHdrph4Pum33SQLr4nE3
L0rqD+c2zgD590uxR5wqxjIFmozUBtVjEvWydvoX65enoLibnG5rgSfa7hA9qBus/+1WsoH/O8Hu
wKUqGoKdvFYLwUjGNd5bNBR1wWGe2KmEsxAcbrnmlZ5kIFDI5jVxXNURo8Jg8CqGsSyhODUZBy85
ccPQejcdJiXc53HeT3dqCBKAO2Uyo9pX+ve5QabXNaEhNXZMyFv1B8APwWjbLQFEwdxtG4dXoa4a
bN7A7UboPeWo9K2m7TR/1ruMzR4yQxkl8DBvuro1GSzJL3fg6Os3HJd1sKZvf1lAiqXLmVG7vat1
UacXbLcQvVay/ouSzkYRxa+T9Das/lyyLC76tuJpJvDmu7fFvuWbbKt7AzmBAOoALQsJnhksHEYH
cz9VOwLmrgVgCxfO5p7dtq+32GJ8pZ8p40p+AvsutgTbzfik/WZVMcM3G7ttS3OJTu60Rw5GSBL0
1THYOnxnI6WbB2RI1dhiiQUjRGkBgkKhrP7PuTgESqogiUYc+tEl/YDMFebudDddnJkCFBCmeMza
TXE+y8A/caoUDiaTy+6T+Hni/lQfA5x0p6dc62Y5RzGvnulz1r4URK5vAi+oCWjdFR3rMIFIsRSR
pK5g4n3laG2Oi2qTBK1SbhjVxvFjP9LUBttgNhZ9LnmW/hL2tJdYDe5VLm1MRhCuoLQnLG6xHlAQ
ee41R8DG+MGLIotgXfYBf9d3jjG19rAL9ri3HHj9BqXs/PqclvcDq2kHGXaJuxfBcUyNBZn04wM/
4HI7HfcnpaqRvvqod/MKA6BcM6vSHIP2nsKD3IaKC/94jH/fvOGBrM1VGElrhHduBiZZerHZ9VKU
+NDRKMuGatDtyeANi9mzd0AqFIrxqhsf1MYx5f+dJ2v1EQ7IwVx0fk66JMCGhYXRkjKVFoTQkjY1
ZJxcX91IWUy2g1yPKu14t3O2HaxQqYLa6vEY/BaFrDp0o+x/0VNUYMtVqWOiah93OPwOkB5qPtmX
TUXrQLJLRyc141t6QzDDX7C1K8QR2oI6kmWSF/hQRc1sy/eoPdJOTTL1LWU3rD+ZkyzI/kmDslvX
01DsrPEEQgQAJdwdcKb2Zm1rfw2WcQvCehHJ4INhPSMD8wu2dlmOnwCllu9hjeLqPpYGpaAKc88b
3zUXk3jxg1SAzspfA1mGzK9pddjWyeuWiPbNZB3vRE3iGH5kp1lqLk2aS9XYdCLuuUCsVXY1GWXR
Lm6I6VY9M15MXpxNm7TZNooxKya58TQHBObpcHVQmcylU2mAZ5GlPNKOfw2h0gDbZj+L1fZSDl5y
tWhwwj+T3dJ9gkepErwieiIkJplLoaupIOTZNXaqZtuVWUGo3W4JLDPHr/jKRbQBND7su+WuaFIm
zSxuol15tyjvAe2hjn2bB21JgNle0jJ7gpXNZZALEJY/Rz3D3RwSXulmdvXFjc3xt6d88KH9Y2f2
BVzRos+nuCfe2HajiroIrf23uMHEa7+XLGY1aS3ydwe49uLnH6CmMyxPLGQ7K+YXXSL2Pdnr7c09
wV0zdSLV8t625ZOrGz0Qx0j/BuJNtRLY1RjZ/V/LX5tD1b6NPQWDFArozqDct5c3VHXjnrb3ozk8
AKjs4htQJDiTB3vyNyibP5sPT0wXc24/n8TyKg8N406pdAOhcgoJR+bpLZSrDeAAujieJwWG5c7m
QtNgqXvwoT0MyFdzYAYbVMA8ESqXQdDM/PZrN6hiO3kDkPd3aZFgEoc6hONt+bbWb9akQe56cDwO
dxCpkcRR4U4nQDOYkgwhC0W7T0jBnxJIKd4Cohquy1XKfl8C69isHXDP2dEMmW9bDLq8LtN9MDn/
tNBRORKI47rUxTVVysD0q9miXaxwOMDn+Cx6XM25W/XU42icTjM4UDK2F9OzME047KjH+qOLAeLZ
KPbExiDGYXG8OGhL9mVpQ5fGaPF9HXm9SLg05wc7wdtcRdcVKPbph6GloXr0jz534R79HKT+/bYg
O57riMngAr+hk+Gwp+lgAme3+yYW9e5Sodw4NZyKWz933E6IHQ3z02RIEejoYlwVXWR53ucQ79Uc
0bDNg+6Noa5wduo9Sk6tdccv+UhlGzwhk4x3dECOTg3Sc72+SqqtO1EPLijTodo/D3ljwuVFfDH3
WJz+IftYtVOwjRa6aEojB2Um7+xqyo9eBxfwD+WlzZrqruBcBk37vP1FoZ4LrWyH4594+TLr1IAu
d+wi4tLUXLrGzwn4h1GDpqOnylbU8SEfJW3nxQIGekAw3wV16v63rGGBDaNjg3YGznTRS9Rhr5nE
qU3scIgDXXVBYDn1MeF9X1+WAX+Sj3uZoMJIgilOZieCoPpRMhQgjU8kdT61ctw6wyGnG3g4xMwh
QlZecZpljpLl79YLSbWKULYb1vu/HHXliJWU9vFoFNSEEZPzdChjRRDGBqLeSdpQKG/qTpMwymWM
jMiRTKJM1+UtI7pd+yiEtNgWA9xn6l/V2smbsSyEFKmo8xafsXS2oVhswdJUTtZqxFuFwy0LWggE
W+IMB0qeDA6L5MQiRV+0uTVeTF+GWsxtvpjvOi81OFP9laoFtaVtzZge2Ei0MBueJfeJQX5Teqjo
IW4qTLbdg3Y5Mh2gNMEbyy2Ts0roqtJhbcDvoufcB1LlL2lZ+Q7ahMbcb3hSVE1c1S1VKKAB6xGP
u9W7e0EhEJsQXCzibpxxfgMQdPXbPMMT9/PPFfv+hLfYwyenu+paN6NKJp1vAh0ClKJJB0xA4VQ0
59q3JiXoJNavcmewRjZIAP1NmFVeTycau2HkDEI6x9+131sQDk6ncyi+XXjH4aAlxLvr94+hF/Zk
cUUDfe1V7QppX+WykFgL+ALonp1t0Q+QK7k508F+oeburtNIgGD6YuMxZ4imiJpPkbCTHvSu+Kb8
RpVhpe9RSJoqg7s2Zp1CNqaY2zMbV1mGqpUqcb/261ixUhNtphcQ/1zlmW/pYHIkkzHvXAilVmV8
ClHi/+ooFSOhhZY/wdOaXsQYWqrwGQLKZpP1FXw9pRRYzhC+e8BB5XKHf1UoSLboYi2qgxUzNauJ
Xax6b7JEMOigSbKcXSERFlYaMGBOUaF0U2zumAlNnbzC8/x1LCdBhb/43WNmpgZnHvcwnRG3/ioV
rsaazT1T7aPafM2o0w7L4z3X07YehBAls1ESe9ABxYxbTEVf/bQGGgJGQPYQHUSX1ZwJ6sndAoYf
Oa0WTylehRqqrEe3R/FR7DgY3IgLwztLZ2beZ3JESKHVDV/ashmEsgv4Xu4X6Te34iT3/VQBGlRo
pCmFVj/vykuPIllGbjFzPCDnSv6sNEJtOzjEAnCxFDLk6zdnBoUxgIKfB/0bwkbYFr8PdiVLsWLU
+CwwFMIXjA07Fr+ADl8Ele50cpdOuwYZgbNCEkKRBWZuMBp/WiiPE2gMaEuyMKrkxTn/gPg0BtfE
dwNxNG3lo0+YmSo7aXwkoVAEdjPx2X7lz92ZlG7I2g+XVpwQvHsstdkl2Rzq3CflqxZ9vgn+TFmv
1ALx7XfXlyVvXQFCFGiZpAILJKxCW6gOERd4p0dh9rCjQTrepD+O5+EaORSt00TQSjkQpEgGxeI5
HtY/ofGIVaTuuaXKVoo7oxxaEJIVJmD2HwYB3LsNLTTkWiJupDSHL6cN0KGLGqrBsWqFomlpqO2s
KOseu2RqgrdtLZulUm5RJl++jBZMoD5Okvq8XMQicI7VTxh7rFY/1kweJM1eeIIp3FrIY5PsYusq
l0MjR1CNkRKXkIm0mBmCGgDWz3qrph9KDFUfttWNTz+4oHlJQBbttXv2Ep6h9TPxK1lvlhwLMn4A
mKuio11fL7u0PTU5cSvHI3UbyuA0kwyBuMTmNO1AEW/Tv8guhT84KiUA/GfMAE8UWw3XT1eRlaN7
a32rjPN5bqR/epPfH1wMNOn/FsxyJbtAC6p0uUs0ON0260JKxQ6Vs51t273rvCBeS6mhui7L/oVf
Z1T4Bwg6zu2RINwTgKdkOcy1k959gQ3N7hJtvuFVaY+QrPwbRywbHhjzWUQ891gxQOXN4qybLba7
Q11wKa62dHJLD8QKiwCojm0cSaZruy1Df6VoHQgkJLMjZP6+nP20njv08FLtF3kBkeNi2CPAUMKQ
S8SNAyIc+vOmla0UPwJ4UPZ5fZ3/tAs8URmyjjcMlrq8s/KUrIZ8MHBjYzkJ9eiReKWslYzBdHk2
hKwYGwUHkqUt15VQzx7RbtUHU3ZjQJyt/8fuPUcANRvZyDsGB1ZdhKKNYmIHy1pv22/mOoDHmyJ4
hr6GUuAmMPk2iy2IRrW4aluiLCHr55AYdoFKuNuia/K/oXcAdUtQds2/g/kSFwGnssUX+Qrui53i
n+Dw5tXe6/tTZI52Z0qa2BG/Upyl3tR8j5l2ZV1a/0OvEBLcqZVs8hgG1xkJz80v89jRrZyAnVub
KkCWXknlgDHpM2+WF0TCTfQdkN+wTTnAiYQifwkVVyk8XmxfA759NFIJnCLxRtcE0OLlCfqTfdFg
y7r6gJT7kY3bam35DsYVyt6H9duPZvnEHFarkKnlL+QoGQdcxZPtxwLskSfQqhSeCzdV8dKEXW14
NHW3h+HlY5gPhWAS2JxYtm26SbDOv6f+3jqjQ8YZ80qcJ6aZK1v+2R9CG84fxbofBJMww5E98dI4
MBuiabfEqFOpzKq+0KzwG6/1JHoddHx7Ag4RSh72bcHNOMi4zG8VxRuT24ktzdUW9KM3jxWYj4Zq
F+x73sapCoACLNtU3//z4QufSA5yGeSAU0x1FXaTY7O3ZXDqhVszA3EYoypnYZ25TPMt1mGcy/cS
YpeXYa7oortMA6vBcIIH4bFV2FD5hTp+wpwY4x5sCiTg3nsHsw7hy4L39muvW41xe1yrQYnlOBRZ
JBge+SLXJqRdGQb44Jw55wlQbGLvf9Xj1grzw0CvUwZwYidjZWWCexpLhY4bo5bE6VQ1WS+4pXle
uj70wpOnDDszg1PO7IwWdh6dlmxI8PX3YdGP0VM+Uei7CX+HUDa/xh9uMSS2L30zsiqh5Tsh9+fO
jw3WJ4q57D9Gs/5ZXF0RQpa+R5Ze0WVkEASPjO1hZ3NorY41Yk3htZ/V9QOxFZY2olbjtWui9qfg
5Re+AzbfZhIzxflJmnlE0OHi4vNggSh/WWzejIRX4v0NPoGVb+uGYAqttQG1Q1gSjkXQARQu6VeX
Cji+Q8bSODBKJh59nwbtMLFU/NZa8rXi+CFNZm/eljmGqjzRBIdosdHJfwjI/vyMRnb+IsTjnX5+
GYepRYvHtfvpoH/XRranDkF8w98RaasIbOLSHIV7CFcsqAo73TziFmIJwMrn2HXX8S8Mochh5e8F
hD4uaW6mBUp1zgIGBewgoQcqOSw4vIdpKYnlPTE77+PmqxZ4edzUpmF3qitUQW+poYIaA4uwuXae
REMp5JZ8IryURDwkHKuwvYJe5T+E4q5sB7HdSJY732Nni3tFKPdBSrPlkayocbfUUwF+eRA65M9f
t1iOlW8ZegAadIOFoCa56Mc5DHKucXtJb1GSKVkLkSsL9xqVJzbUoXv7GvtRqwf9l4CJy7jH95YS
zi+yeE4O7jXRQA2J8O8JJlvaajMFXjD/+1D5Tl/asZRExRz7kDn5hxeOqER0/qUdAmRcYdnu2tUX
axzfwbRRpxOuSULfpDW6oX4yM4vOKWfFa1DBWZeoS2me3d7ZdE7aLp9OUOmT3zRbGP1wCdyix3zN
3otBamQ+1qAbOTvQxaiMcKIEwH52j/Uzoi09oJ81BDnRO0WopLK+/iMjpLFIv+N8GBoVxh1c
`protect end_protected
