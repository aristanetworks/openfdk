--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   duplicate
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
CixZdNSaWpNMf+3ERcOaYM/qACicoLfP/SZoWcswxw3bC6eKIVMOGEIPwoLSm2J61KakNArtaF1O
XtvnBDrhcVQuzav2HZRBAB8EqYAyN6JgF0Vo+69vUeRANG1lj7JfShYwzyA5d8qwVRWCqxD2/FbW
HtinALIhGreWzlrBOJI8ZLiuHNk6m6uQ+ljAjMhYFJcnySLCO8uUQxpw2bPiapn1M0LuXT1kMZtI
kJruXAFh085vB+HMbMM2lbX+JOzusv17q1dchr5O0BE+SMvE4la6Se63DQTUoFcI5B9PNG68x0kE
yWB8Vu4yI/0/G5OV0TqkdOh0Mmyd9W6LRoUB4g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="NPxnXPAuSwdR2z/4TR98szEAzd+F80Xi78fdKafa1dY="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
F68ya4zu4hEcWEd6VWziirV/tLQ7iivCZAnnWbVcGY6sR+dicLZ0Md45PphlFKtNTyZJmXJm+yXI
FpBJRt4Q/dlj2vpc8tHqC8glaHlH5U1LeCShgdDCmKSxdD0h7l4BXYqo8cs4QeRshjOHnnRHnkbf
5fs2VNIm0aCPl2Fq6Hl9FaOxRh2kOptZycNN23RkcOEkTJ8ws9d+sQ+k0j2RnvuOuKPxTQ399o8c
3nySuer60eyyRx3ilJ9N+ZDGVYcjThtAstFrpXicf2huQo/2xV3OerSwyDtTqS5WDMC0SryL6PRF
YhOQahtPHKMteMVkFOtGOPNeI5J+lRgHsw3PyQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="NoxNW24jsBUJlBbV2RXtADwGF1Xs9J88dgacF87dkT8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22704)
`protect data_block
vLHKs1k7DohKbhawoXzGF0QZQvDCHjhOioA3YFEOZB/Ixvi/GBeRV5kPYTHjgGpTY7vr1xqES0Qa
QPuK+cqT/Dakbr5JUyewb8+ltFOrDPW9oXyKSIDRG5m3xHhuvblfdZMkQAU7Rzhz3WU5QZvMIAKI
sB62pQjZ7QiXtFQE7jcWMP+kuUETzq97bHEN3iHwRXFzCEGg2BA3pxsYuitll3xq2vM8/y/UDAEl
uYkiavV8EYmYiWDdFEK91p1qDd0VFSR7Fxg5DhPG8KU7uTQOa2GmY1xjoD8K0dx6Drf091ZWmFLL
qkNzWVxCa57QxnkWPfSweMJAAgsbqoIYyUJCGSEb9ZMN2EnEuTtUwt4HFT1lCpewi2/aIofhKp06
6m521awjEOb5YozOTdMYoK3CjaVE1QFPwZXyEe6WUYhD6qgvrZMHNfuthVBnh6D/c+40DNjB6uBI
LZt0aJHaNVIRbBr+YymbDB4K5PXm83cs8uc+du2sO4pCW7PVOAfG9rQmTzruC7lUyKZJWKQu8HnP
YT4JVMYD+rX2qorlEaji7kuVAkTzZB+LgosIHhjZXXtCcI/7e8LP38DoeetPc+om3KkBlBiwk+Ar
DX3arkiZvD5+3ErJAtsvhVQXwUsbUvGKl+VDi8f898aFk2lyrN+zPXISl7psT+iw/pf6uBZ3HF5I
ugks6/haDCiBSCbqrlwpoUYyzMnwiEJ08AndxbTZ1Yn1+MHZJZoLzV3gT+nVDV7hEuSTJU+qLFG7
DJrXog+rFEWDCEkvkfMPztV8uav3h3mcu5D1LJJfCOJISAvRkmlsWyIwBGSrJbtYtaELOHQh6id4
yHnugWxO/Bs0qD+AJuQntKlczVt8rrIJ9twohxnKo39L6gQPc9/K0tQN4DqiflznMOWAK0FvRYkB
tcmc2Wm7HYhy+ONgsMOy0+tQ+R7D5mn8qwUrnq1mBpOoVN2+cKVsSPI9FJYzGN3BW+z5yRiaOvpN
X7vLYDxPIcUNxCIa+w4meADxKLGf1d4QK9NAkI9CKLzT8+v88c6foHvEDIVfJvwbXc76ztwioN3t
x8ufW+nEpFVYGaRoV8C90Qw+AhkpoiBtN5NqNsOu9GSYG4+G+Q8ZELHZqOb+I/eumpZbANqsSMqD
mVprJoJJnmncv4SC573lbS/6vOf/W715a60PdW04KiJKSv3sgjeAuNkupPz+VIwPmAhaPxANxMUB
hRYpzn4mUZZfQxv3XbnESMgzpjrmBbCHO4Kpfxh6J19r95R8DFzReUORfaQSmTNImMSzEceDjlqS
eNk/DLhlhyV7vLgTWEM3M4SOBPocmhio+rPMdske8o0LtGycZJj2Z4becD0sCMjr884sA4Roe2uq
y/RqFHnGPpqAW59xYtui6wyOtEfYThC+I4b5/hf1uXPCBrsfytpNTaUqMezasJoeTb7ih1vUlzrh
m4NF69j0Ok49PPNsmaqjpcGQ7G4w4z6IHH4R//fy8POyQB3apnzSbhizEcxA/T+BaimVy1QYVD2n
jJd1lJ1bMzjYWZYEyVOZ4DLu9XRUY22ow/6Uzll1XU79JXSwKVWHKzBjNikIS0hHYKlZZyJgpOyR
MZbm8TUtpYqI7DAtBbyEyaP/B6QvrBMe2AsfCESFRn2IaVFEnDQjyVETvQo7qH7J2Pz6kbDFezZf
PfOXiP7Qb3qE6GAfI5mWQwiv6lA9S+bsEcAGwUyw1oReMH8/LnRgJSjPImlDVG110W+UmTQ+X3T4
TWCgc6PtGdW+xgzaqhGb1/KY+BxoxMc5geFu7Wvsaax72GanQRh0AeU5Z3OYAEMNbDKZ0LXOZhpY
4wPao68vSxKf+I98Z4Jrwhh1Kg6swy4Ofocf+m4qi73ma7XDt3Lmn+6aMDACZfsqWNZ5Eftk3t0S
Wk68piYgf9337VeKCWFYC0fWCTGsWPeP46mA9dVlWzMMXnUFd6Vhyx1GWy9k576AFoFl3alvO1Mv
cezR9SVuU5Zd0PYoB6vji66kP6l2XuE6c13mGjjFOQBc+q8ZJMgUaCP5zA8bPoe3oFzNRw6t7anv
MQQw5WeKteFgWePw61qrv8iievxN8eYClnDzzBDwcLh5ubUC1MM8+oDcF1ox1MuSJ4VIwN7pDpIQ
4iANq0k8G7ocN520/LV4qE5zVlbdXrkV/cHpysK7VKiBDQnV8Su7pbnBu0yC+R469vTDHvwwGFW2
4kevoAQWjoXF9k8ShcBQdrtWTelEJlJwM0mqNxi14gm2LjthPC+yDK8w3H6Dpo5r7hwn4HTZzcBW
jN2dr6MFcUAGNCaVWtjdrYXqjwcqtT+JpyO7IX4KwcC1cbVHlKRpG26nH99sxTtl7k06Gznil2wv
9bPJbkiYBSg0vIBuA+6Ctvex9iBq9ELR80KA/75ry3w9phezJSKeT1b8yY23DLmW6oPVNLzNXHne
2+534fgD3QHdgmxocQi5Srhp/z07jgpxe8f0lBukR0m0Axy/NySPxye0UAM1y/+mMIKg2Ll0WXsJ
RDpvHjX1Z2fJIp3T7xV94ptACL5sNqTA1Lev5N2Aq709amsC+btKrU0FToh7LWqpbLLKTBw+y0kb
tHSM88JEa+j+wkWEcfUVHgXtez8L2QjmW1ykgYCTL59xDMIqdSmB5xqbqpx2tFqy/AUwg5cvNB9C
SlFKx+crZcPdKQqXUvYhh8y49Z6+gB61bX5EFKb92I4VqciEZUjbaOFEdX1KYP9cjiSnDG4p3dL3
kIP7lOVesFB87Rkq8jhvn8qL0Lootkt5+yNbSA9hA0yROSneSeHoVZD7PKj1cJePMqTWZFv4nIV2
FGBVSgkgVdYxxIg/R+ouswvUdzQbVquvnpUBtbRJRnV+dJ8gLqh9lLhSQCXt789xeBKRSa95stSx
510Qu4ftQUdWXxeF0wj0/aQ19/ph40ApnvaYe6S+s4w8xzFd0iWCpG5LDkAMRq8MWBmA1OywbgND
N+PVb3EdcYzuWhZ24XV0Q6k7n43KlC97u29eE5zFb8gp2uDIIVk/kRprCpD9s0MyFO+bgZ5BXfHV
qvr87nkX9mxLz5GafnAHI0i6TUfX0qx1DnI3twSdgoFcBigeD+fGHCtDuHu3pfjxRgN//AzY12lR
aeLwZwvTyd0d3zggnAkKAHg6x5rY6rP/KSTALLU94UBI8TVJgGRaI5BkpsJnMAtNpZ04FtOQLg1E
lx9cBZK5VHq4+4YzAn13Ne2mAKhz4UKwk9o+sGsLF9k1y4hNNsl+lsds5oW/ovsZ6+X0YDOLBZj7
5hyDNf9ArxR77oT4Znlz39PRWuxx7yqG4nmASwJvens+OmJAIllUIPfaoP3/Ps4LeUQadVJDiyAX
1QOUw9oT/wNWecOu0yOzH4whjlOdUnQQVyzKhgDGmwds6/cM+o1meMWlOcDptQmZGf6L7hQo9nGZ
5RaxpbSSW4SCIrBmBWILaOJtHy6DskaG5oTeyYA4hOh7fp95NCcinyvFfW+VYL7A2fy5G4T47hPA
DFYNsQo7BkCL9oYyGVLqxr+S5ws+BW18DaMiUElTtTFSradvx7Lf5v/iHpN1+I2cNqRmwZZ6xP/w
YSOxA0UTUL+sXlojNyp8/CQqn8pbzyWWCQwHLPzydQYprO2C2Rfec/xazq/TJ2jQEXS0Kge8QGe+
ZkBb6FpFqLeMpKM58CBZ913MpweTp0GyEDYJgC+gNSmPvKev5Ql3wLcD0LWI/3K6P/pfD8LDQXss
CJd5CwJ0ofZF3AYVt8hvdXBpbpQKJGbJxilO+kaQVnMElu3DuyP6n37mZNkv1MdTSJ/6H5r+Uj+f
KaJ/Qj2wi9LBVHDc77tweC0CvN3K6cooURbO+Uo6v4Kdo/Of0u+GOCR3ach/8vFovUsbErUmmra6
Af3M6cqgnT/Or2IK6/uWhOu7HsMjbDPe5UUHCgpPE9NRI6cSU1IDLpQV2TN4WIqtP2MvEOTmscs3
7tQJ2SjVpJup4bARTvDXbVSKnbDYBefxCSIMl1vskfl/5CyaarqFgZHBWAsS+69aYry+U2fSVs1S
5jTy6eOunIu+IVNNXKeRodyndXD+W282Uss4TqDTAup9pdvGNjClm5Lls4u0W6uxb4WDb76CBLF9
3EGDEZXQ0aEjFoGVCTq8v89oi/gb38cbsTsjV9r23RVnzTqdiO4jplbNrNbnV0ZtuoMiQwCXDGQo
mJtifECOcpX5yfCsY6XLBy1qtFaHWVEDY5LA6koS8XLSj3VpCnXDnVEndVaan+ebO6Odi4coAKQ5
TU28hrw2GQcEgTR6FVWhgZtWKsv16zBu6uX9DxpMWjx0jUoFxrpotApwl1pVWLeUHXAH/FDrCHsJ
IMZ13COlFACeDWO7EQbEoQlY6LVGIM+VJ+gJtRrfUDZvCVca4gC+fpFdcw9l1NtQaCAm2ihEcLjH
MBCgzCnU1rM2ZOGVxoLRFD1HNuuZ52lmF8/bIZ7jQ4pmBvfCA+MIxxyy7jP7fUIOSDhpGVWgRb3l
HAgGsFfzwM4P8VznR21Fxkfji0U5fudly3eSjCoKacv6voAi+tRkDi0Pxs9NSORD0rHDDU1TEtYK
h6aGpEB+N46KtAVnpbh3nmDRbOMakW/Re5u/7XQlcfebHlXDK+YFWqxs4fyduI+i+kDfsycawDJ4
cV3QlLa7FrkCfArl2iw3lsTIMeiFzI6fnxzvROHpJT1ERKgRA0L4dRgyp/jW453tyMcHiyqPB+dH
SaTyfSbbOGSlfG53IcSOaezyYRUuK2VrutTIq6OTX18oeIBoZUddF3ha6yJvf6kLh+wdX4CeLiPF
WPfTzyk/Q7/JykmOvK32k1pVcffwWDXv1zwWEkht6ZCv6K79IsPSb753pOSZ/gUVQmDxZzrk1u9g
0fh8ds4ilszsB6CvstzosWq2szlElwrtE/9C625rJv3ZaUiUpM7jBN43MnqWJiyy43esjCi3wHH0
YqkY5VZMsC5lAtAvCp6Mx1VAPP+m0Oll0FegrPxt73Qx0xeUYttKylCZTonDKOTKDCWnSiWIwaL5
WHPt1trYustQHgJPefw/bXXhMPMME2/dpmQiFfl9dFpR0yBHb0y1gdb3QaLvwpXrg9ZzilHyTi7i
rC9qLxVFc1WCQg0lK0ewGv8pIt3JprLMBlP1E6pD7YTc/nvXunppahVNCFMwJ5DhpHgOk7M12LBC
J7qyq2F0LG8RCB8Zf3cjPQymAJZ6huxgOgpHxNVOMCj8zLvFceM76cQkGiaR2zlmXlV+msfGyD2a
kNU7O6GGEr08HImET0i+RwsYind/C2mk8xSB4TFmglZy0xxex+WuVHpm8CJJCgx241wRDEEf2Wlg
B1mWvwCDV5EFJzDy2Q8DGAH9eW395xNAIYWY+2B4RyVP/USx6LyFlVwk9x7kVFAo3ExTliFzGr47
Gta7ytxSes2zU/wbzSJcYGsxzbfgfRKiuMG3QnqCtFRiqGmdJI7TnA9S4cEm7XZfVbiex8JG57ey
p+kH6FDnGkaODuYIf8d2IUHB8f4tD2WvXpipIy8om4PVZaPORzB6YuVTt7CD1HyqUMENFdjErH3l
aSVcos3AgGHTndLJge+tmS+wZfyQkJwbSu0pIUbB+qPKb0q5XSrQi803lQyMff9TYGbqk3ug7nE0
t30TRJxCZI+je0mEEz8InEas+rkzNt4Zejv7pyKBB7L1teVKwip8LZRgrqFLopTtxLs0AeHIYygI
NrS8zSMR7VRXWt2xF8HE8JPsQ9zfB5pKVXrRdSFQvzFJGF+FzQxeyVm8muCJaZDkoe0HmOErUDpX
iWLLNck4z0gMHLY2Fdo3SRaimmBjkHQCcg2eysormsduqpEJlZd2hghJhhNhIUf7pW8P2Z8N8Dab
+F9UCBRFhg08FLz4ZNqG4YMe7Vqfzh/Xi0zUMl9yiDrJje5ho06CS+5WYj9RSXaGGb1oAnQB2ygn
tG2+e1mD5kKuQM5xTZDNylG9k6sQ6gflQna6cyw4GkG9/MIj+qH1kHyO6wiFnrfl4NXMka/F8npk
7sg2dVK8K665EixkqJfaD3vlr1a/zHGXabAUcdt5fXermliOqOWaUz+lgt6EWVGRaCKsRbok5YSt
584blywqOKf+IvxgOoH2WqD3iqpSi9Fjlh2OSBUzDT5KlawaR9tJd33stfyryUD7WW8jiAunVp3V
j+Pov2GhHaM8Yapnvm8LVABPC0O6b22p/L9yrfRBMVUmMb/fenmYZ0wWQsOVJkJ6WF5AFKPRybCl
HYn3ipjsbECVb5VBWpUx1XzMc0MKBEnTWXuTfC6GqYcBufu9eY2HY5gUEToIELr4tG7V0KfVjC+R
sMNwXsH5N9TDW5IG5Spq8FvzEaIbi8ZGQ5d8Sf7JZgEeARArJ7tIzqoRM6qufDNU3zPYIXIHzexg
hGaG9RBovfflSLiaTZNUK8E1s08Jha6ymzFo9NvBXxq/UTW1M+Cjdgo8IOhZVIw7k7J/yUsr/fv8
inqxBzQ/d9nNY+8s6MY1eIT2LKk4vYPrsG2t5i1Q+7UpRhkbkQT+/rHsREDLNJ8EtC5W+2l7bMU2
iFv7Me/xda0jxf4WTm4QCwHJ73LEzdfd75uFjlPtqHXjs9CEoRt1lEiWguOnxOmdm/B8AQuukNwZ
HO2FQgkvz+FtMSwTJbzH665m0bmCSaeFpiqq1OqjLkwzv8w/negvH8/qig1GFl5/KhoIx2RTgin1
G2iGaAiql2in09KsBdMdnd9kN2EevbkovTIXQ87wzZC9+SlLGOLOQqRtpLEvhMbOtd4oJAa/fTop
mNR7EGALsbMJ1NAcpP/11SBPmu1qpsQ/p9L/fhadEHB1a6a2xeKfgS6sxwpz1TVeiiTsY2AneKSR
EcgCnCGTvusTwIAQSsIwncBOU5Syz+q5SsiIpxKwLtLm3m1Z/0pWp9wh2D5yl2byWuVtGYR5UyQk
qVEuc7WqNwRWLw5PqtMkLvNmz94Vp+qMIoL27NuTo7WmUBmRExGTSbGGbGPJPonZriipuxuM+4gR
j3VfOBB8sH3V1Ii1CK0sYOHehah5lUg3LasoIdhtC3sD54GpNMLaNDA60vLQrC+SyTIPQlPgYfOJ
Ebbhkx+gmwW1DOye3zjcuQEoDo9c7eUna+uRTraNbFNLEtfslPFfKnzN2D7iHS7VROlr8u3QhO2s
2wA6v3oiGz+/Ltd5oxORnRpopJ2UoOu1fP1rCyDoEFHjz0momhdbusrKSJzONzK8kNLWoawS2kkd
AnnaDj8Y/Gajh3XGUZ83T3tcC2ONp+SEPGedp7yHKGbmL36T0n/+BZA0qbR4TuR78RWR0Ohvu4B+
v06rN8PjhADDuaLKBKaRwhKoAGUAeA/rfsC5AlV3S0BDFYmxi84UAbubE1Uw5q+GrrMjobU6pC1W
fGcxSS3l47kuPeCsuk+6G0J1bWtFw3cFKfFZIrlcbegsRTIimjYSFz5cj6vMuB3ZiDgQ5tHDw6YW
q7TZphL+r/33/+H51W4WfYQZYyFALsDoQr+IorK5Ay1jc6FofVWLThAw4yZQoR5k81PZLaMN8/lG
LCb6tdKqP7MsBVjZz2QTdnvoafcPUtp+faQQgrS1PXgLua/hzqkwWbb1GVVLjYK0f6jcWfuf7S9d
D4xzxTWeoKySVyImu/BkK/zu7XnOoSwNze5tpSsu5eUFVmQ+Ln/iA5BbevlY0jVZHaE2wXG2HvqY
iIjvAmx+o3Qax6uXLvUfvWXUnq2bzBcAlGpqAGXC0Yo3PopoyAmr+5D088DoVGbEK9cQdfOdAC+g
fOCQOGI4mvZBe0G9AXJNbTwC/nKf99y1Ra9ic9CAxOzzwroHV02V69gEsxtY0hoTY4sgW/HPhgv9
yT3p/e/dVQHrKdZmMlI2+6Mt+NjJMXflj8b11Np+kU/Jg1GsC46KDzIFbIffQ+xJJQO2QS33Hn6G
lB4T7Tavbn9CYI7+fs8UkUgNtFKTIoerfVhOqhmN0tPlKQBOak1ccff0whEob2cPOOkDGHttk7DI
jPRtTeIGgGvVt6tIyK69qxrbg/Fw9go1g8L0qp6LfUuWdlrt2CyFriGdzhenCiBb6C4Ya5uaqZ37
6tI83zDly6DgWrr4t430jufHxkCqPSnUvH+v61KfCpNgALDNH7PKb857H3BVsH/3ST86Z/CmCQ1Y
XzkmfOwj5QHxZ4qdXUe/aPqcE5G25U9o0CAWb12N3xT8fq7o5krd1FJf6wP0KxNE5kSUm1AdVgYp
Hsaf5phzWlppsAfRw9N/1nkeDOEqajtTBree7d84X06daTM3AmB5AvmizsPTleoeN9PuOfCg3RVb
YdLTunsutYBerpZuoHtwciEvxWXco7310nj3m58jYr0Z/j7d6mRRQZm/NicuRa0N4ut1AzpXKTtJ
cNEzyw8Fz1HLzUg4IKvKEMHvOa6trYv2YfzOUYa0vEbQ4/W+8cmZudA6RffL4auep5a1jP63/x6c
xEFNfddVMyNi00Gv1gaIq1PB4Fu5o2HK1gdLH7e6WwynbjZc1BcLs18w/Y0sw2lVmHlsza+eQVFa
QfyOP6pA03q+FD4mL1o00KGjApfX//m6YFU2ABsh7fXAf18y2uN25I2BxveSm8PEeJfcrfqj/qeX
gqjOPOn2PCeYQEKUxRclyrqSHfvgxxJP1B1q+lkkAKcwoXxuePu2WSDfEd20D/6yKWup+JbUF0MH
RdcNQOlEVm4SrK3Avf32GdezLK2iFESyLuPZThGYlzt0tYQgsDdwmA/tRQ6PPNsiUDlhn9msRax2
ulzm9GIi6G8hox8bvRRW9GaVFI24Erl5nGCQQB4MKwFoU3A4u1rSdHfgbbBUZKlNk7lC3aZ5fxQN
snAtwYuawOH0CC8md0lV8L28ADM/KoiJ4dFW26M1XIXJ5vWHshyv0xj0TW5VDPoPQT2YWjG9MuXQ
cEXdqDdaA1h9Ob/5M6tT9SLfkhdgT7WN8W8YMs8Mstg352lkGaZA5QuO2/SFn4yVaG5gtbDE4PG2
AWu3fXg6aoweqfFiAek1uliHZpL8/pJkk9fpOgV5HVB1/EXj4QTRAEsZ0QY90nnaENlk4XGnZR7Y
ZU8/6OpgLEZI8ptJcXU4aGjNNhbSMoIS1rhEqGHGsOpdHGUHY/XTpi68QTOxN4wK56JM1+KLniJL
uE7qBVRl3PJMz0+UxF1c4NaApUOzTV+2YWoxaipDuK7b9hHcrrOozojv1XChijg8TaqJDqNgKvci
NQrZpMcYeFIUWWXcp/nLliwTFSsvip3SFYOGW7+hbCXF9husGawmwDVqnZBvsbx7FDuHhuDPGOnO
lmi3XnUHV5Vt+Dnw6ywISIcvX72ff8O7WdLL9cRi56H/CNlxVi/SQC6d/sr+Hufo7NLtqB+9EYos
FSix93JoE0QKgaxAGyx3WwsGLpB/eYcL0uWO5izKPvSLD+Mo+Ubuy9ylsubKwWKjYSh8Z+HIIXvF
sH2GR1Ss+WmVVMSjAE6NFHWWWJrvSR30XIQdgz9qUtEMxcbLYvLShqNAF5GoD8YUoVa3Q+e13jZv
jfAhMlyM9gM03fAlVDdciccmtW6kl1zwz5WPa3ZA6xWTYwICeRzBNzMxyo/yKeJaIXd/+PXf1tOo
u8hmek3/8d3CM+YnWi9frUfL9U+Ijon1VkuWKINMaupe+MmF3l4IYd/8TY7A5heI4Ugrpe1vTUAU
bJbcJvhyCYKcmthM7HQzAA8Tw2znmXvm1GOnUC9YEcru9FWKlZKXqoTEOVNuSjtAk11NOs0AWw+j
c4O/Y4MFTjYMd/Q39H5qlpwiaUAWsb4QXVbkw6TJ+1NW54jk+jGoX2tlw3YZSgCl3KQUxW106/HH
L8xw9Fldaj5HeXcs7aEMx2PjmEWqUxXVhjqlrLhTQLW0TE2mCQBy0sB40VDhIcLfkueHTBSzSFAh
ADzh5MmucM0o5witb/QgoczbvRH3gMXw2A8NR/H6axULB/1Ue4+EXqzo0DIE22CVE07bICqUQzn6
yHu1Ta3sGr5i6563pgsxS7fdr9jU+xS2XdeZNnr4eq10ivVKtmdmuGZfkAzLDEULlEVlKMtDBPHm
+eX3vCbxI1KWVJbRGRT1UNpn4l1ab/CcnY74CnH+WPR0Fbyx9m+HucaSKj139+ICv3+Kv0nhiZ5a
B/wp/O3YbupxerBDJ5FlfF69sAJACOA26Qb8iF5xx+KtZSiLWhUZXSJkoxXj7NwJtiirAfTLWjMf
PQ5TdQs6pvGRxdHqFSkWcjpKG1sZkHLOrl/N5WaMBHbbHmogMHeLeyQ5N9SEMrB1u1bJz1ChRqdF
NBl/1oII9JLlelD8orsHV594k3gmNIoimwo/DUmBvRL1czmKxID/vwEttaW4g+ZZTzf2rQeDtEUQ
WjvR1oydwUtVrFC9bpxgIGflAGkWz3vEM1zHsNcY2Ou/gCV9elVWLx81n9IgWeC8gFnyVP2hkB9R
kjfF6OpU5KmnPzxZxMHP1a/7cbJw2t/FCJNyKE2TbQ0BxW2U2I5nE1yco3LmOAPD6ET/Eq7xzpOI
O9pGxPzCYyKcAlYqi/tOKsBcWKz0h4FlRwIeH2PfZwO09BOzx9YJHi79gR49RM0Rf6O0HCVy7rpQ
cgrTQ/0MSkp6S6sv39aBxk23gzlt8OP6fz2G/c70wmwoTv3vs2YGbqoVBURlfF7RZNo3+g1XVELb
HXC6ersP5A9hcuQWrZLnYU+xVb1mtniTRGRVTe7Z/tKZUQ8/iZGwBP8howAtgfRE2019ls41w7tC
a9kWGoxT8AvgRI05oSWafAH4r7mxg/zFYgiKwL/a160c5mZqS+/fIlhTLEpcZqyKA1WvQ/hFndJv
sDDIYDMw403ZF4vQtDDTEm6C/Uxx0w3MSPXXMQNURjnWet8JrwOWtmIr1vVicNdARNZcHk2YHcrp
K+pCx/NydzMrwDMDxYvSw0CWOR5uQkcHSllTxhhDi7RCno+q6E6Phh/OfXL2nyp2x92jgN1CWGoq
wbxQs511U/AZ5KOoTtC4eGih3ttN+w/Rzl07Tq79PucztZveEmXWSCeB5yqcvmw4mhwvYtXSeEMC
lKakXa2QPMdx32AojDHmLMv6+3MDQZPi7oGPkqBx8+HrJDTVzkyjdQ3h3aIt3EDPaWj4+hQMNiBp
LFw2RYDcmudZc09SQeFHLSsJ/KdY2LJysSaRQmVzThsYMGwR+QYvW/VtqBeN3WZu+LtW5larelkU
IwSCgYJvAlksKZTwl9azMSAKMBG7OqZbGVhHto9nKSwj69yUYbu6qh9NVKoi+GkYenZRhTsQ39MS
MbYgNPwlZFtZRfkVMzPIKVzT1YSSLO6PZ27/Aig807Vz9X/XmyKCJ/OL5246Lzd7SAQQg9g/JSHa
S9Ifq4TvZQiQ1jDQJbJSNMCcB6tqv8rp/bn2Ew8W6HXwrbxsClzIUUe7MeqzVHDq2zlzeUdbXASM
v3b41JnSAzIFoASJmyaPrd03ALXfGjonlrc2w47k3SzYI+QG6qGCd1UY6/PVwkXydOp+GKMmo+JR
pSqqeQ8oOZGFlPZVmCV2lN0EQM9gUC0MGRK/OwYu7/55vavRhyoNamGA2rtSEiXx+xs4RE6kchtv
2Sb44ZojAgXvxrUKJZnHr10FT1NBGFNRTNkegTH4tZ26QEsjsBJsOJWDPhzTBWDZq3aFEcUpdcbx
ecICAjDJS/HS0pMG9tKsljxMmS9h4nlmSYutJQbldX9Vpoza64dPsaxZrgsa0Pvrpssy1J37YDuu
/5uI3hmM2Kd4WqlanNz54aCAwYkApO3MMKvUDpspQvU/vVRpYm9Lc+Z6JyDD4l/mt1+SLjKGdMPy
ALlpdih2VNkoG5yS8aapKY1FgHl3tPWsMWoAzJtnQClsEGbRB0BE2IZ7YJLRUPwORFYeXJmB72GF
yYg8CPOdAITyrH0VqhsJw5HJH8hWVY6KiaIYNasbHzoInfB1x2Sapw9Mqi10eJXaLKQ2NCsWXzMC
B8MKW3gEvKqm9sHqldQfMXoTbi3NRh9i1p3xzPYvIwSltNAPtMqq1qowNND7qbXHy5lk4dUeeCAZ
+wnJqavYAuiVclIqtkWNl+DarIvZHVcCJP5+D+xYC0tz2NNVeE6pI5Ugk3Z3Wh3V4YYGfFQyTSJr
chEvmIu+sVXgFCJxb1nDqpwSHiUVGpWgWd9YUK2nMCKyr9zMMrSb+zWX0ex5Ey5LPFApqTrZUuF6
FnjDHSXZyPMDF/+eKSokEB3NKr5ss/DnpNtuB3dMCzjs3ZtXd9JrWrC2DEzZy/obtgNu2hYEjQoW
67Uf3EUDTsZzBjkiIpzqLIW5tZGvBB/LvN+0/QdfJt1NsrZqINLxIyZoleRq6nTiHErw3dJpkgg4
OtDgE5t8sAFEkiHwEJbeLfhP7qzCmswus2WeXDcGq8YgonJGiH21+CL7SYs3+uRCLPzXG95qvkL0
6GbHEaCVae7wuMBYHPdrq5KXPvkLfRqv/E8sps5+LTHPwyHCxO6j2oE9CoXxy2bTAC/7X+1B5ndk
9L733kl1FqSXQUF//Mz+v4beRnIBC6JmfO/V5ZGLqQ4kYv97yMLsrvfVfc+BuGk7dXZqCgsR55Bi
3qDOivwsAl8kQdUVgN9HRbldIBfGNqoDOpfOTiLPoL7Uo5zwYPW4y5R4eu+JLbL4JulQjMmUTF5k
/eesxkdmQbNN6FC8+v0nNBuF4OcH3QqwVxjsgBTKHS8NtxjCZ3uPlRP6SByV6ZlfwVg0rbz9yW4/
12wKCYIvyHr1IMqT0/H3YigbFeOAww8/qYRmD/WkILA9KV+Ay/hHGYryM2kgq6WPzIjj5JpCbcMV
zdkLq1N71e+PvbY1I4FUHy0VVvVSAZqh7j7kx0K9QPlYqkYDAJD2CWbMhC/J0mkIgjk6spuW5uDv
GaDnZhwQ5+H8xeEVAeFtSjjGrxqGwDkKYQIXsHIEJn1gumAos2IGIrwRTnO+QZlZoqUbUITmg+eC
Z+EM3R5j8oqmLQqj4Ow0UoIkUxtPA9lW5YJe2Zv0uL1L+NKcWQPRl8yQerhbTfCDChCGAWWBj4pQ
XNjRKhATOCdPURYLlfgjMnqlKd+KACGyH0cr6y74/EuPnHamXmT+8qUVIEjbEGyusv9O5JAVVNyp
/6Bhl8hRVVtHd8B1eMpXz4WS0OBbZheDU3Xw7R4WFDOVBKDo7guWd9d+knRTLvdfpIROC7EfPZ6p
3OoSRLVfdcFrMwtkLZRELj3isAu1ZA9+oR2qO2u0M9v/uV4UnzBkWCa5h9M3XYG+CZuFuZqlR4KY
qkrfGKYoOfH9+OvcY2lr0QfO/wcnmCAiThlUUQ8J6gOIXt03KLeoC61d2XaqqxKhChuvicVSLbkI
+NsR+M7Mr1BCGvtExJSmRTGkEG+1kklB+bK6A/F7qdqcOaAhAzr+DxiyqQJKAhVJCLAZsBR5zVso
tDJoWJGQFzjkr8euV3p45DPznRCALm2HRRxFJeUCLIWpAv98/1HDN4YAPKFLAUlVB9fQInzAu6xC
v+YmsfUeUH7yOYH9suAKcE11mIqaXF5CN8bCF8XWJjMSbKmVuZA8rOnInoF0CMi2mNQ7PJy1ZS7o
h4FDcBvBxvBhl1/MrbM4iigR3vzpaaBnOApkE9V42qcRwffjruB/s1iRIDiD0PEvyz34wZ6soKbo
qb7lh5KX/TwKO3ovg9DgN4pdGxGk/OGZycfv0iaeXibnqAxURlOlou6NoPUT39qPKJWwzfsnrkLy
s2smPDtc5QVXWDMlbcMWnJ3UfluUeUYHiWCQzJTMYYN9TYU8yvWedS5EkmLA+juTTZ/Wh+2yPLW/
4C3VIltYrbl3/YwKzQdTMMPiG28Ooy0HxeqdOGfIXNd1RoOoljBJerw8brA9aiz3Kirm5/jvlh1y
jbyAnx2QMvDsHK7dhgBXKZ2gL2ZoAgP/YhntNgBtukWlYP2fTYr3oYFhAgD+vDrEyVLYH13x3Aqy
tNdrdEAvaJreOsUrP5dqULn0xk6g+GmjQzWUPIPuhPwoCKRus0Gthi219mfKFP8TEd8dhvF6RCwG
IuHkdkY8P6ezcTGcbXQsjP3tEFG8rO+kbSuzPDlK0vFH4oOsSveJf/q+dhEfIKYxjjJFhXcvRjQd
p7EbKYLFZQsPKRmSqdOV3NFAw84UNMoPof8CfElXMWqFZxVM8Ss9Q+ES3xyU1y4tJ2GKlgaYI6vK
kd4OGKdhwv6mHVQ0pn+nbbHPJ3JjkwksOJP6a0KixXvoaVaR0DuLDeeE8GXZs5tNer5fLmj26gyZ
5YxP/GHdnKl6ebftg5hGVf02TDg1rXMPLT46hOf8AUpPpL2P9KrEy4xaL+QWrexykAr2B59WD3KJ
pAezbSgAoXpazl2+P92D3m/sBSgko2LB+sCRE4ZdJVCEKOQfdDV3ed7nnvbSBdbvAtzjqfJHTxOM
owd+GK6RFDk08IO3hpkmbzRsJQEUCAHdn00wGtXr1mQdajUqsaPpJHQFS+lcU+6+MbahFGDrBgrs
4soJZKohLo3cwRugLxX7O+5pvRCBL+/GukeZQHOK9UhietMbsmxBuDy6kxNWpK090sBvi8Z+CUwI
5urbHn4CkEbg0GMX9zm6QBkaxH8XjBMQUNKnyCPkCQLhkBHoPWOZ9ZvshDPAABWgOtUjpWuDhsp6
+OOA9xDuxNCF2P6slXZprCn69pNf40hacSB2heGJrOywfbO4I6s1fqKe2Y05SEH39QCzERtwbEHa
XMAfI9vkNa/PKK7I36apMGuCoDpu37W3dsQgi8IJHKFajcmSNd61F1PNxsaWnqMPpsiRlZrA0sjT
vGWtMfTa2RSzsY8dn4Y0s0rBbEHFx2rGn0I4eTfbZGW16efBatw7iXjYEcrBuVHA/hgb7tjDKsqw
ksoH80RsQ+w5yUkEz3IMpMi1HqGSHW47376MOx8MiqomJ3IpAh/CPpwn+FFr8FE5auCVsDNeZ8wS
jcesxZKH9kv09sTEK8L+IF1qvTh4LbLAWDLtsRq+5q0R+tXnbQnxK7GKEE8jqDN/RnYAtaXcZzbJ
9GmCM4nP/MC53dTIZSckiRSO+cf8xpuRXQPwCbJDNnTPTDtCxmcoen5bXy1p8igwXk7KIKJ55UYf
yTMZI06ATGkzwrtPJII/57S5J5B7WzlWxOOCqforPWlBMOp6EBjrfu6me683SAGdVHbGuBL2tu34
JI4+6vZmCtib9tXzbZ/NStoBNhdnOp+QMljrrr8rhQ9xi94ghr/WBBuZC0W0JxnwJ45QDsEY0Ql6
mCs8GvFE2wi3MfXanFFCyzhsyIIKKk7Z3NTWD7PIsQfQkqBHL/xdDPMpqC/vM03kFTColWgWAvr/
Oyei3FhCm/9q1YwRdyk8+Cpga2b+apZ81W9KOUprjyhA1NYPRGt4FLVKLN5O+gaEjNn+Aynrd2R0
IAkGRLW2yQU4W1wIgtPn3C+Bo2h3HmxWJDGGI4O9kIkHVGLRkbuiVxRE0ih915QpiK/RIWq3o25h
HyECx0Ux4rrCXY9aQyCPNnThDQcymPnj7Ro63sWH8h0P9I1HOUA9K8hqnIesyMQ9KqzmQ5kiRJu0
x8K6uIMNrQ6WYEfxin2l5wfTomeVkIb9MSWcXEcJxo/VZ/7VT1hKoSHEy1r8iwuyb923+GvjFeVR
PToltpmcEBzGJXuERppdHXBWaQUkicdenjTfRqD3eCVF4qN9zAbDSQ1M+dGXpnOofYKH12KO7CHE
J8UbMV3BAVtZvOlCxtH6XdR4QB4wsso8t8pHRrfiozST+x6/U+Xr/rMPaAjNE2BxDXkulpsoEYPX
pE/k0yY3sTNyNBWrSZulBrfJuStekMxBv85li5Vgrk4DmIP8vvB3oi6524xQM9RkNyiMf4DvjZiG
KYh1Cpzoi7Fk9Da99mLvd/9xgPV0fe32za9LD9RIij1Cpia+LTcIKcEjmG+fDRjXTd7H1EdB0yks
WqIouDURfGec/Bag/Zu9PZmkYJlTfQnQsNNNCDAomIHdeh/F/Ditkd2YAeECCkt7qViY3tTp5UCJ
D9IVXd2+FFLakkwXWQFnotqri30PnbU86FZ2OmPJyYCDJHQe+vdX3UeIAAWlEgetxc9XtdJJ8aDR
/56R2O+f6g7ql7AR5q/Sb2DYCYC++URw2HGyvE+DATtOy7m55E+yZcJXT8dUgD38R/M0+lKzSYXw
2Cwc0VxxhcWuJYtmjP2Jd5algw1qsGK8fxq/uyGlwKJ081N64AcwHrFXwRN/tv5A2ic/4YeNjRo1
3bR5V0KzpiD5vpFoILfNa/61cXiSYnWGGsqO3YS08DvtyC+hvQfDHtT5zpxXcoU5ffpV1gOhe0yp
Kc8s6R5BSXDa2/LPX/VDI446qmo00V7du5diyNU3lufVEiuZRp9OoauuMy9ps7WochuRwfE/dgFM
9htuf1ONnRC4mYDGLzA/wUaYUhSwwpR4bIanLoK5M3cWdLY1RRfGYYj7m+hXdOAz3gcD4t8kd4mB
AfsSWmRSaxCyHdx5YY0ks8aAJrFaGryW5KemDJKShmH/iNz3ARRLDLa3rgJunZEneY2x4JOCeFkR
/SCnYbaiDqUMjy5aIiqFGDx8EvDDICXYaNexyy0WT0UMYM5OcaDeqEwsHgKRPC5YVC8LZbyYGsLY
C57vicT1YkeOQEOxWHs11vPsuxWKVK7qYIVeTVdpeS31rm+rajNWUOY/8x7eyGeDO1+bPCRJMFkJ
nb4fJ4qeoki0Ri7oUmrWAQJH/vObHP7vb5NqnWZjjpqlW4jHBno7gRQZrULLX2ZuosZ6gbsUKqRR
0MonwVP0caqNkzj/zsK405ubGwear/E5CPhqdeWzUNj7VWfptDzmGKvcKg0GJ7NOGwa545Q9FSrH
p2YS26UYzjmA+CX1mo4k2IPX4GgMuzUwI4DvcDqFcOVT/yKR/7a/Qa2K3QzpL3JHpBr1uXWjLHkJ
yJ5+0atFmOLXeRQ4cWwM7BiUibUbXrCka7fJTy/FVr4+gacrdcObtnhTw4lUNId2nj8patgvWiU4
M9SLbcsFY+nT0F+a8HhuQFfsiGW7FSQJ53Hh++73JKWM/52Ey2sSkMT+nxs0+YDdQLVoAy+eKR6A
D8cRZtEtGa2tQPcBwxLm4kAH35OpeMD9RISUEXrq3qPVB/OhQ+hHe2IRuh1b3aPCxu6lCb7uNEnB
10XqeubzXmEoK9W7SRJaRamf2SyKsYdkivU0TzHkAJyqwkHjIGUiyCkihn1vT/NLsD/jgBFkph6t
1Vo7B5hJLLWBOBOFaIzeIMu55Q3HdmXEt1AQbwY7aduLsSdtfF0SV+dA62dSn5+mxfl1eKjaA8z0
1gPM1W6/hZF+G83/4IdlPDWofVzLs2fHOte83V/6jPcLIiBLhzuEZgZC7HUrWaXQXZtYzAgrCov0
Fow6H8soiJp/CVLHe0/ajW4koMIBplFL3COlxQEQJgvKeYJ2wzAxskTN5RwI4UbuOf3CSAOC1LTa
TJrAWtGND/fYIJco46UFUtpB2pWQXZMm3hJe6BOkrSqZGDxqPymmo9oz3xV5wW8PyzpzhHJCLv8I
gc7EzAoDO/kFNTuDp0Zq0KOLbUfcwMBazE0JlG3K8T9dHkKmVq6yGOZV2SUpRGg9UKxJaK4goVi3
Sv07xnZggXyS6uqllTI2DYPLlt33zdppYIkEzpZTD+odpJCXWOBECgxAKZNSdy3TdSLfz+rkexpU
hAWYxGhvMJnvBwRJE2YBKdVqOE4O/B8ZSlKvHYq5jN6ynstxcRI5vaLfUkTOZqjvj3kdYYHeI/92
o5Ddi4h1yVN+L1FI/BnNgs4pGNplEQWl5k7pH3i/DsaeY+7UbxRTk3Ln/9BKolJfw2KoN2j8EZOM
XuS13KOTbKTURACoBH7qrilGlFusHwMVSmbE+cfAPeeuyejoeQo+VSiBQP+7AzVLQj5FEU204qYc
03791lmq+S32bh/BRQL7Wj6WSfHyChXJZ1Z2H8Icwab4CX2sAW1heLRuR+k1QjJ/HZWz3ehX9S7n
OH7Oy7Ah/wyGgVWldIbuEyz6OzfKF6qVTL6cl159HZG0p8SLHchm8LJ8N9n+0cRAGSB/bZoNzAwe
zM+eLkURD2eGehKH+jNPqACmnNBR87R/vysWCe00uU798s7GNa3mHw1DUHMYVEKVwrL6LOVUab8U
JMHkukX0NhNa+0cJZUVPGbl9v8Dl95uzzDddgESITictF+MXBdnHnYJJN+iveKVfbNLrkdN4bpgd
v5zV+PnUBH4jprJX8N3KJWgv7Ngq9GFYVp2dLjdsLZzyb2J/3ggWDRTyYF+LbrISy6Y3GtPprbg7
OUedrj9eh1uCXBr0CjTO6IRC2uuhEw41u63Mq5en2+MOKPQhhX2AbR9d2FK763BCj4iQdRxK3e6a
iE2gW/zCwwO6FYTsZ+DTDmjp1tonpbK7CWP/6tSWHVpbFc/nr/eOW3pD1geA+R9o26J9jkdX2eS5
Z4pPvnWbdbbV47421Sy9gYxs3vphhF0oUExzUE1Us29sFJUKTNoK3eQN0nlkOk2Ei+/jXgQpLmzh
SL47c4PyVPa61xhCKLjbgLxTHeP9E8cowlYSSIlaIg5xsy8Ku8jMpm6+oSCEIwoSefk5b4VXOvP8
tzTjidfq+IZViSuwfPaaRwCsYD4lVM0fQoKs+EpIHbWAsw+MrFWpwWEh9ao6p2tXZx1BGCxZOTB+
EAGMFIt6qlqpBmTFi5oE2MBL/WaYpQPc0jb+hlE72Sou7vwOk0cxe7+sQvmuZP0iwG649KKLf8ul
XqMIHAlNXtV+OMpQ8AwJvrv8GyTt9AtBuZGS8nsNmU/XFfL7RiqpB9oAQhMIS1pLjn+2DFX9BiS3
hTwTqzqerjLOs+HWvVsRGZ8vRU7A8amxI7E+Jhxw0JhgD3RxPmWVBBJtE4Dhb6Dz8LttC0JDlmKs
Cjb1vnVo/8+BIhBARz8vx/EGkxwa3f4TFaBo6VA9rpfYa3buhW2M497z4MQWNt93CQlCK2v+6Rzq
Vt/qQB4b4s7OOKRL59de8y/55rDdwxlva+K7u87NVwOXo7d9QUR2ToUdhPxXyskBp5P2dTfmJijd
Z+qEJJQXm2fe3yZZ1sxx30dLUBT/jRVdEqcdKNQ/yxNa6rBKtRHOGgTA1LBrrTdXQWP0Ulc6L53P
LNceyL/yS6KAPCciiwwv6vHWLqLQvol3kvjTh+8kSyMIhLjxdfIB2LoErfa6RWyZpSmlr71KZzu+
ud6oy2TxPsYQKNt0zDeKzvp5Yv+MHEkT7k0OnIud6jiidJCcuqHyE+Ek4daSxZtTcBsDjZQ+9K5E
ugYP/O6ZRIEKzz41wk+IY/JM81eSZYuD+rKcGOUmTIoLIQ5SZlR+3DrjSO1kSX4b5GSjATrgfN8D
+K115cllc9/AyqFw+0kpJUdTkDAMYkLy1sRhW4uRqu32AWdzOxi09HISVZWZ7z9/KwlPfuX1FkmW
HdqmDGBgc3DthWHwWejLTENM6xLX1aWjM5Pc/C0pDnNwGeNhWOjZc3FZsu6lYx/xecgQKLR+oms3
1GyEA6ijf6czgT/s8H3cym2P0WrS9Iot7QXYYHlQkEKpRW5iBPpNSCW3tgJ2MO4af1h8L7zaPX41
+QR7sJFygH6KORvkXMlEsK03dWf851nfkxVHVnp7jLW8LAUX1kZ6j9lT65j+xoVfY8vNIbys20Tq
zMp0PiJFZROIoDpZ4MlCYJmXHyPjTaabFEwCV3PXP54eXDylKgEQjpxjeVnSMMGdWMhFbE7xE0fx
S2jW02BKQQwTu4Xg2V0Ve2Wp94ivC26GiaJuuNEzsHIXDbXl3zEZCusZTX+A0fs8E/0xg6/xoQa/
wE8FW4Cb2hTx8sd0BZvQN+86D2QEO7uy1gCur3U5EOvm6Q0mqbcKAXcM29bhROpPFZDmem7IECuF
sc4xlLWwdNKjbQ0HvFQv0JFff7CsXzGwawUzfFxfZtXqdMAsQBdfXrEDgUokt8p/kWInJKRr2y7D
Xcdaa3L2aBZci95tMSm257IKTNPdbwG/Q0od87WmzJ2Bpl5NLrUuWKOf6McCpciOTJgath8dQXhJ
zsyd9gIhZrKr5R9HuZyPbO3Yr4hH3qbOhJMu3/o9NnnTFwznCCHMBxiPyyMbm6b40xm5TvVDzJ7I
ECiplA/aTRY32L9oa/phpAm6fjX4dUloEFiGJzIsDJk9nZqt2VZhAhkQXEpK419o3vZtz9O+s3fE
2ADN6A3dVgHGKRBJ7lFCzYiySdbG9lSeuYQiSlPoAkArceP2VJSqER2qcHxVWCsQDXIDfGLSmdHg
xofzzu3+qDrbIPXlr5tXms/AEBzKCuxRNKv9CBrk7lotBKpRbQBeX/VRHD2hl1yYWe5GllCP1xsu
2geI3pwloCTK6N+OC9S1HSAckLPgVU+UIw0GbARDiUMbsgXarrdiM1eHKkQUqQzlHLmPmUqEyKop
jHFlvOnTY1I+KCD/83fcYwup4kQ1zKp5b3A7n9/LoRGo5Rtz2lIVOkDtg1mjlq+vc6WFSpoM56JN
uPeVSpShN28KmLZUvijp6VppkT+7E2yJHtAdq2QUN70frydr0aXQ4GjRVX4E8ZNSiIZEkhsyA71I
lk3Y7xvxZX9ew77u4U8qWeamLtJkAG1f/3MdMbiijj1cwM9aGddP6wlBHIWa0szNC/eZbqTDffg4
5PJWNaRG7Q4Jvh1jGoLtcn8XKL4vwEljZ82BW/FNo8kkGprrUvOZ3FUmIxjzTEKLkquPYq4o+rsc
lzNj+tUOzGbF9G+7D5rFNN+0Sm6wqSbi13KcclwNrlj5aZh0CgUiZabFcbV1x/JIlLPwZgEGam7f
P4tqZlTpcTj+z7TUeUM54D5Ocmek8mWro9ooAfuy7WHTzEkGGqS1o4doYwFNX7y7vbHugqz4LYIo
7wgRw6EticyYHO8UFqcN899Ocf9cbmgAK3CK+WxjhbQM8hF7MSlRLha2xEw3WIyLGgnHzEOhuLsg
sgxgMZv19jo+dSWjggzP2oxvAvTVfyvAA6hAEWx+7soUTF8cpBDu2zA/P5lAXrtZV/T/yX1I0tf/
te08tsd0603a0zPdbiWVTsNpsF5gjNcXDh8KwEiNIwGEnP8xUKdmO+x9Ndsyn9aglUb1vYJqf4CK
R1m4R8uMOjFYaGE9PSW9BPv9TM6Vt4TLmlCMBL8lsmZ/6zb0QY/G1H9Kbo0tqfzoT/MWKB7suADc
rIXf64hHyXXILmpPBHOwx/wdxo1Pyj27LvH80rMSzbsLmfqjpI2dzDCzfGvMJloGyFfECMC9MKQ0
MVqwjvev6oFJZ5z3GEEsRIfPb93sDpFiz1qjV6Qma4bxlPQv+t6tb/65pqCMqV41C8pkuBVLeoiN
KfQvLCrWBIfJXYziXlYmZ8y6Bqaj975pAxS1U7D3iBXMZmyVHPK1A0TBdv3W7k7O0T6F+oYRR0W0
P1ovT5eko7CdNFtgWt7ohTvlEDG2fymskggGZRpmL/POoIG1Incjxv2LpB5QngvgRgJiSVGOOOjd
JOBlcCGlON4/zOUUX72uVHo3lNGJMKBB4CMroN4sdo2L8LU7fKr+CPjNuuwI1piElmUQMLwdn/6X
YmnmtDLCAN4U/EdVTZTKsARQUAlWUfRZNQNqQUgNr6tnqOc9L9Jj9y8KAuFR3QXIPQPiTuUyQOLl
oQGqWze+ry73cT2f8xf/9BplhXh68BkKyLmm1ncF3/lEhjuRrh9xvG+jMe5KQ+0LZ5XRvf+QLIBk
MD+agr53Js3lPXwsEVlPeqppYB5aMBwu9xBCx8gXpXmYC/dEdC+88HYXoOL/1nUEr7O4Ws8HisLQ
EJY6tMKaqUJ5myUZm/RTk4dBaRZKRaT+OEwjwkB3+H8nlC1CbNNH8ZPbNeNdrTPuyFaaDro1iGi3
cH6OpxVxJURuoni0f/A6wrUxgL8+tzgdrToOefNA2tUMCTFccviwZAoKtHyFHjn55dSExgR6VZK+
K8zTS8nOK0WhzCRE5WO2uK7w1BPksNhMsDsp8TOyl/BXdzKWLuBdU73aTCftEUsNwlCxeNZT+hUg
x8FdiWIlYdTV7uMsblhWjIMpPPYwTAG+rIYfIM2eAUGhIAjAtHutxoNCgGo/SoimY4XGkagok1ur
t4XIxnirtL0aQZXvwUrbn/eCtRD08AVTOAUqDzQMY8RCPpMpU0+PBXi0S0RI2j+6XTSEBgSRXoR6
TI/qYVVFm3kreDfBilGafOyKnmeeUjczJGfdEDqS9CYMXmXYAqe1fYJwytur8CxgXx+P6nUd6CB4
T+OW4qFh8U0FVv+Q4NjMJtqt7SCtGGrIQP0kainE0xxaC6rcHC4o27fdugU2kinZAH8mWZg18QJA
5j1hJW3p+X+gkAXozRjzzfNnjPm+2ICN4588O9m87xP45Ak8pfvQhk0Q2CwmWxQJ+fjx8voRcoo7
H8X4lTBpWqHKamSxvv9lBd12/k3C8/lQAXztXlDQpz0Ks9YFRcE7NJBMTnWW1Q3gwQO/TwGneYwp
7RLJ0EP8gXzUyVdyJxBnJoGgJjxsZdRUs9SsKJ9VRvcEdCPxaFFTNch6w2VfUOLJMLoFrIGJNAsQ
9/+Vm2TPIesFq1Mb9AF/P+3rkT1axkxMJ2z2pYnVzvdot7EtGmHBJ14GfF+uqS5pHVNPWG1sEtMs
yd/4HOgE10UkGux+zCaDYHfXfc2hhHaMomuMlLFzxTBG9JrHgx7tQfE++XN4b82Vlr5HpQkkgiFs
hauL3YvXVuliQyZagqMNHiJozAWfwI5EUU1EIodSj7hB/qSqhYo149TV8x4PtQ8USWCksnpwN2L4
OTrFy6L9RyMiE1CYmfFha+QA2ZA+5l7CNpmiOsF//N9NqS8PFCGRJ6kLz3dXaebcruP3SRvOVyVo
Y8Zs3XXB/EKjHbkqtaSHG464UfOtetKRgmz7Aazhw6PSFn68KbJThYuCFTLrc516FPNo/GBMxPnV
fmdBZlrRhKwpgBaYiWiBk3lPUi2cpeqd6JK5GvLgoiS+VRvM7ch3Cm+lNUZtrYMbzA9g4qoIfN6N
/4e3wOX6t0bjfsy3zU0Y+EfN56p3xYs5oHif7yWKF9+ci7jvdPW2Vo1rS8XM/oeF6e+/ZrFO3WXU
fn70m6E5CDfeRd0RW/rSyXVQZmw7ifwJdTeLJvHZeYpcfvu5MtIfJArCLR4t6rbu7KWiYOe8Mccr
Y5ajmOneUvyO5rkFK3M0goA51scqz8Uamg/xGgmhvz+NL5mEIUIvuSN4dJkeQHQ3MucnvXrg3iad
mBnUZuzRI1pW+BKjpjIkDIAp9ahExjuk+0ja1fP3YbysI5F763272PR3sIBcmO02rVkF/iE8xpYC
icWfog+p7hnUDefBSygMjcpuaxI2rGtED8NncfQy+RAFod9h+2UQkakzgvle1AxkHrAvWNzxB/oA
cCz7QMt8Wh3b6Etpw6cRzG0hDNTeAOKYt5rY5TwUhhKFPJQvVjtjfoLan478hiBMnvWxTvtSZbMY
PHCp1BgcV8FRLn2rTOUjZiQH2YB1ID952Y7xprGcfoud/Xo24QOpDwwedd6AGL9VGphzfqnfkyBY
waY2rMUL2UKObDs2GBX0VgoSXGyPlyIQKM1zzvODvtkVl7MQJXNmh3EV14J36/z0AwcnPCcxlrQz
ifbIm0iLEpnXltSDGb0O90invmAFab1K7xJSM0JSr9V3P7RDa9IwN1NJBLHF3kIDF68SXe+aixX0
U16arSfrBnSm0LtnIr7YFYkUvRlnu7boSTUl5Qlcyyi1RIsZbxZDkEAJ3VXwSMHTMBMlpOucpzLf
sFScZamnh2yo1ICEqHUeXXLlUoNJtBMUszLSe/Uogu0ArKmWtDFO5t3uSui3DHx3STBM2QByJ6uO
MNF4kOX3hyIju8ETzApSoR7GbI0rfil9o5qLqJNyX9ryDw7V1rS0lCL8n1SylHnkA3c78hM0r8CW
IpMMRL/Jjl7bgbuWbpe3iRHX3Gd1zDbicn+2Ap2QQpBpoRhXc3WAj3IuhiCv1sVowdbTWvo5RGZK
S0+S7chJ954mYAuaWrY1Kw9EP49AypPH8zT0zFNiULRDBOi5AAobtBVQsACiRUgsUCUsY+ulQ/YV
E7HkGkZKqjpfiz/X2fGGR91CZBFxmIC6capxRcYwpwOPaAi+2TtTqOpNTm4AlpA2qSz09SdqcafY
FXt/i2PcXZthd/WFFaQqgDAgk9Emrgr2uhrBuMh/3cNQ6xScHQM4yZF14KeQc62SwququyJvMsQ+
Xnc9oBIYmtMyxA2Frvyp5COVvHOJWHwq6m5dhzCBX8Mv0DwBQVtrMObkjXaShS8tGas50pUtG9Ps
NeVh8f+mVSJOHsFFaOMpLbeYwe0wTZosFkOzKnD3b9zyL76E264gdxPWmTHPgguhbqFDjopp/KQq
6hKwZpPFZ6uDIDqy7ilwHHjl5df2s0k0Sa8uWIZonhGPXE/O8698PVDHPTOyR2+LQ0pcJ3xMWIrV
0WsLoYyWxcjRTPb5/sMu3zPHMrFLROw4Rg0abub2OwidUSVHUEwSOoJ5A8bMMR8yp3G+kSJrOxf/
dwS11kqn52+J/EiUqlBvwPqrbLy8CULGgTSVfOundb1Tq+fyoJ7ULxiaSGWrq/YgBt6M3l3atWRH
fREExsCgL7xYy3Z0k6Lvy+GLA0NAXaCHC0CkVdb/BpWHGaBYyVhInuY1Ba9on+jWpEN09JgmrV74
RHs5MzjxXeBvY2xj7ciVg8g/EBgapoKVIh7R91EZQ4ChEmJJyrT/NF9pZfqiD59FHkZiThjIlSJD
C3dOIG5ITHx0r7zcLFFHMYw0MDuvVhG3ziq01ctaWpQJDSNAb0gxfqvAGnxXkgpBo4yAiLHwUb6A
7TZlbfoFNHhuwQyeSAccNZICE7WgtQYq11/U6If3GZ5nBD1ZZ1renQJHxQmMsZgqWcoRv7eAmbgI
irmPOBSHI9MVQZY7eRV2ytd6zU60RFeutrSmWcP0V3eXmPVm2N4nYWOhoYar8e0tbVXAXd9JlahS
it+5z9vRxeG3+jPg8plSruzxqnFlzOpmAJWjN9ZtlmykwVPGrKzIVXwmeaqQBEWNVnH+dU+csB2E
bt1YZJ1+BzKGlnDYjnSDQo4V79v9c0CSsJS4ZvbfVjIFHqpBbhVG1448xZM8fFvVtPUvt75q8ZFu
Xwakge6nrsiiqe1riErh7LHbQnAJjxRaqnBwRWG9Jv9mh0oY6979PlLciu7iRqRgWomoa0cRz2vQ
kUPz/gGD12fi6AxZ0i9RQThI+ICKUW/5hBGwtYEf0aqAwzch1gn7HDopy909TPcscpfQgAqnaoEf
qKdRvSD7Q5q36iowZsOwVHvgIiyCD73W4ls9OnJ/jrSFQNeVsRCnFrvsAyj3QNrl1vmR8UnrJ3hy
rfriTXPljSaPjw1KG3gZpmjP6SAnCBJS9dRIoeIfiZLMFgq//cdozP7WQ/CGcBrGQ7LApmtYP0Eg
3otVr9VSo4grq95j49i4w2O6WXbA0Q3aSL/gM6nsNL5MhIGe6rcSMnJYGY/6WOmlkBv7Tba8JMC2
qTX7dVEeQ8l0juOLRY7QZ3EeEgQK7+20t6DNn9Crgp6QyZsWSJFREGPv47YZm1uefjC53aJtXTuU
zIYjKO1RPZE1Lc06OJGvjkfQTdOe3l5TwK6W2thUsPoXMzPale5c7wBvs94pRX/IXwWi6LolMmJO
h89WpC1fPS3ZsXqDeKk8ms1IA7YUJuVI2PyUmDljKyBn6sRr/WqX69k4bZpXihdwUmAcSgfVaf8w
z53zsLUdhdxaSGlWkUGRZ4bmpEiUSG8ks5ynHmFIolBDYxx24Z05Ke+QRqEVfC6CDnNRLj9MVcOk
f2vYH15dP09iXvJqisxlSx1xQCaGh1kwNsvW+Ib8IwN82nwURnTP1bNTSYnWOzvEXYVNwLERUMl2
RIuW43x7hnmdTrqRkjnYJcXkmlvdkYJMwAzHNI1M52kP6qZATKdaoSRnwFZtBrI8MdrVwHO/QHrV
kFQINoNQUPdXGXmHtwCx84V/fU2AFnHb2ueCCTY9crVQmVhbSdw4GVVVmLgb5Hj68/aGg8Jly34o
o5O3LWDn7tfL6ktCnmMBuc8F/ND4w6nH/NVRGFXav9tJpgxEy24C9ITLogshDHgjNhtrHnjwOPgq
1c8Olmkmt1yocLkoZFa/pMW8R4/CsBmc1EqBKnF5DhJdIcJXJqBO/nNnPKqTpknGNBX/AWqodWeH
lETidH1EEZNYR8cb8gJ8MXoP0E9ags1YDaXGgPz3/FnAE4PkC9aBkLovh8q5Z4aopekKcIrmyNXz
aE457+4TM6xrPpQgm4YIF30WtAVzNMXv2h9452QHTApPJfRXXycZnszN58Tt4Ul1WLkp0DAxvAR+
gGhJRzeAGRTXIMeQP6DbxLES07vsg9ZZeTPcm9zzPd7zZ/8REnOUGfD4+KKI6ag/5bgumy5lRiPw
DOvfNzsirT+w1ilF8sCkLhP52kX8YCl44M72rnxLOCz0/6OwsN5GN2YAKTQNQn6neW76l0eogzdK
glaX71TaaPMVeN1M2BrZRo7Zf76PEJg/1U8uEs3+p+Fl9VAjPJik8H6Vw9IunEJX38C2kXz3uB53
CmyqoXyAVgncLkmtk+WANFhrBz57H4mR+7ezSo3BbHgyy7c3kKhyVuEu/ojS3ccsDbk1tH8qJNXr
6qwBliKFj3lPKPqdZreaFrRAzFhaZI0X5XLGYanX/UWBn0upGF0bBaMGMCFXP5h85WvG76OiPy8B
mepzUOutDo0/x+tkHJYqbhjLmvtvrGBblNH1rbetxa5yaCxTsIoBniQtMK30fvGCXMdjHQx67pgr
Itqy9Ro+ta5SQyVv87RfMGpsgQi9P5FR1fIGwvPWJhwJLfDaC3LYx1LQb6lqvk/QmKmW9KkHqY9s
Da+jmWF+VoB4Ln1NhXLd2bsurN2WbTDNP4MdHyLpEz/zqPNR3870k9Y6ZR2HRiiM749I/ns6lKxk
DVS1CNUv7F3F0M/gWh2Olni9496qZOmUePfuMOWLVkl5DSddMjOeUfRCeEtIJI2wyNPiW+zgHovX
ijqozrLpFHcuZ8uj+Klek0L+ZpLZqOWndFVb2VQv1fpQLRXKERN1z4XW1Cs+4cc5Gtx6/Q+AgeTb
OdudV+Uc5Uk4qTg0XFcI91NTBbs/5y2Xo4cD5PsELBnQ1fN8enpuBgLnzm6tCVaT/0CoY8Lr/UEP
HMGho7Cx2NQl7hqBXrFqdadVFq+h2wdYX0iJhqfTfC9vI0+egkaXmg7ZYslmeXkBvKZwlNKUayTT
NYXO3ISxM3Kw4b+C0LkuV6vLI7SA9juynn6s6qI0ga9U5WSyHSU1Rqdgo0N6Wx+NeA//038sBNKh
g5Yz7h+toKDetc8T0bSSkavGIX7MLEXFiVMM8n8fHy25SN6eAtg+GfRhXpqbag44UQYZcjQQLdlo
P6bhxxS0akWIQDZpntIQ9EOuGS+eAXsT1mQwFqK4NPAl97BpX4jRn9oOeS8rRzXLhqJnCcGOevwW
AiuMms9dhbFFkbEbZu2I09NaOEMOix3BiZrGsuzRzhyFjkUx7zJWR/pBeVM8mq6RrfKQmH4K6R0r
Ian6U52k8Z9WbdvIqsHVB7vTD1G1ZdUPrUJtJlpxCzKyZdQA6zcqDJtZbaXi4ZQfrgg8jSmB+1Q7
krxOJCEFnjc6jZRl4rIgB3yG30cMxksppjZfO7EkX1jQgNt6q5eTp61mebNjCaYCA7+d9CGPFEfx
O2NuX61UQL4mwh8S8nwC8D1t2LUxzhMEqc1CqO2yOJlGaj1qctbKxYFkPHa6qUaidjhHWOiDGQqJ
MgTz6akJbIKUR5UUYN79/L3WLI6NrmEYk+hzOwmAj1eHdLw+rOxUhxR+el8wOJl8SigotPXowCJq
qvUfo4O3Z9i3snKQXUl1rjvEfGbJvgxGkd2nBGcZpCVjCsTBk6QAvMEZA5VobK8lvQGjcV8X6CCV
ruZSsENkxihsNuLiuC4U0lLc8euFpODD7J33RGXSWvE8SCkWcTwt423SSC3To15gcAHeOSXVhSXT
SunE/Owy6t3pjfp+76jrbZjQ+fNjrSfhh2rFm+pVDYZEXIoCIqgVELbu6gkrHY7Nv7+y0z2n5ul/
suPh5I9bRRvLPemSCrNIl73Ce/LT1pJrAkA+rxMFjfoOe7CxmXUmiKHkrjZR98xf3eH4PMzSO1iQ
n50wbIoGf26fG/SaXQazWk7923tUevsNfFUgciyLoEAcLTdH1FyUESzNVkU0wNwJ1ihgs6PxQXgk
aVVSliKFzPRt59tWq1t2fuKVUqcALu3MrOFtDwNmlWD+L0Ql1gAu0Uox0kgQC1mFzn8Q1cEfXbOV
gS06sI8hodeNMMossIg3t7wmH18kaMFs6WLSe4GSeLjgpfKALs0rHnCMyz0fu7nN1H3pJc3qVwF6
sdddnQGPQ0pO3WlkK6ttSq6Kp3tOPqaifN8EKT6XkYa2Pl3O2T/9qrD1fghVDF5dyVwSTb6aHmRx
hYxRdc6bdH03nJajZocPKRxAh51KJT/1I6Pl8ROXbvXx+z6sUlgi1YLDDAqC72Crcd2teax0hBET
t4e16iC/VuBX05yFrgoAEI5Jmei+LsxlgvIAic5/qJzU82LGTyilrcPwmYhrDn5FKQLivdUA50c9
mHM5m5AKYI2pulVi1aM62tqcvwwnsFrG8gokmav0d1gmieOUnUfIDka/w25TsAn+zesfdPQmOqDM
JoUKAbYDM+4c4e/OKn+cAXmXrMp+xEiPzm+mCeZrrSP4KeMHRglDHwsswRMBxdxJAjRx1YFCUsya
QMskq5D0LhMTCpZJqgNtAIrrLScuvIAJWbi/5ihS5tYaCn/BF4EoVWX+cY3AzeAdFDYW9aut4BD7
36DJpalh9IZQUg/N9/WVZaX7zoGnjAr8rqQL5hQRHiucYaK3nMTVdPzLEcegUODN/HzzpRkIjiNv
rTsWqnRCJeVWdXwtrh6lOOBSvUbyemFPtrQ7vWWYY6Oh1Qh0CZ8kOnxtK03AOhU58cmWppey4iOG
tFb/17tN4LitmV7pk9I3BXYxZ05S+6aEu9hAYnNcaG9Pm0tndO6xnrjMD91iaoid2zKuBDYfuqQZ
xAioAvMf/+JIm7QrXerqRMr3vtD+abAgu98dkPdsApnqvu3Jip/h/Db+KVJyFB1gpQbnF6r8cNya
S7k1gp8uEKz7zIDkTyjoJ23ukiskX6fOyZIRUgfgtX6wEaPnA4a12lLOZlDXNjbnRumOw9jzYJHy
5jOeBI+4NJnKAT3ZczPXiHMlMZuQ0DJZq+1qvr23kgxCL0XVoK8EHS1v+BR0yhnORH8+yNi5mV35
GE7Jois4AMVuCaPJBhZwTwpX9KoftwLE/c1miNvi4cqGgBSzAClj+y3L5BJcLEnHib5JwXi9QwsZ
UnJXgOQVfzcza0ouoRDo5VoOymEuOXL0QCg7LGVoBik4Bj6lPjv9qpgTWhUpz7m+8nIW1xwpKkaF
wG4lbg1wbNy6ydgxfVA648hBlv0jXu+rwpE4HZuFp7U1PUD3Lpd2B4Z2qIgpGwZ+5S5q4P69nImH
ZTAVeULWi5JgiAY3kkPOZ8ZErn24YPN6aPcbGPTh4jrRDFbqStae99mhFVxXDTJt6y12qwXMUY0a
hlMhPZ596KUwTVO6wlhTiP2vjmEYKtkSYsoU6b6pjIiLNNV/C8oBjJuwdDY5/yLOSBbH6tzdJGKw
MC41TVaCKSJ7OxfX/8kzw7igbAP9K+QQuqUy5wXpJJ9cGhEApjPW8AyEfLeOl73rg3O5+GEmlOZj
rt0E01OVh346U+e4T6LoJzesdtDs8XxuJqgGAHF4m8pNPM83UBXxxpzNCVyRvQFSvBvH7H1U79Ut
vAObOOF09yXHOFKeKL23KzrwFzhz0nfbdPoyMTs+9YgDwumKrh6ProodEpH1MHfwy1UR5GK+RunE
UKhH5EunRVhzmAYfWB+u7ROUJIFIMukknWQHb9YwzLBusjqUMHWqpEJDcVX5U/RzxRaetOrlm6fS
ze54G45SIUyeod2ZsBhzjlxZ6+uW60bF+PWJpQMIjlVlJ5Q+n9WUlEjhyRIA1kJQwsnsrPR3N32i
ly/E55tFOsgbXhdIhh7CWBbMoUphRSQPLwSl7gNBDL1D9ME+Popy9pbx9VV/52+GMh+j1AB0ERCf
Atyv2TbjGaEOtH5DjB2cnDuoOg4Er4h9OSxau5Ry8a4KzE1RiCo3aXVLzEDTqTN30T931p4295os
Bz9fE5IAkee5icD2quh6PEp+5iPv4kCKPxYO2D8fqptqdPtlRlkBXTfq7poUJl3bB9zf9Ee4YAp1
Lb2kT4uld4xryYdwoABBV+Dz
`protect end_protected
