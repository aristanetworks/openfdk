--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
UeyBFZhRcMUHU3sQcaTWeZoNs2vdw7SoMByTrv5KNe/yv0qqiyLsgZNQHsyhLcq1Hv+rLhmKali9
OTKzM364Ajn0vU2sxoKJns3oDbA4ly/SGsYdBo4xs5+U0+0739EjVdGrcA6Dfwf28464nbiTRTnE
GKpCRvtwwKzzTfi5xzI57CFSyuFlTICwWcJTgAaS9XkDL2RR+HlWddp8JX0+6+xh1ew0lVhWnITZ
OWaFh05baqugH8C8v6PfQ/qXfDPDuFG85oIPI0Tk7jMcNqiLwlVAuHL1Z9yuLz2XhdkB7sAfMgkD
GMcsJGjh7tHbcU8ZCyL2hlqzxJzlXINawiBPDQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="d1yuhnF7mj3/1eJvYSlTW5rcVGndS2+tRCVglftEkUU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
SSP0Y/BKLfm4omTc+dReo9OFvs9CT4zUCrUSGDAkZpzWA6YvHCwhK+ss8I8VXaPS55JZWlJpon/c
II8q8Qgdo+yhemL3aFT/yAo456JwfxRPhtA8iGhaWfuWzs8aDnSpukaFD3Gat+diigT8e4eBJKF5
IYhU9tx24UwzrHkBkZX38JEJOas6CfCUh4ca+CIS6OKIaUK8g3YkAmbFl5wU3d8cMtRCeQSpvCWG
rimfgV3GByMCkOLUJDSEMVq/MVl0mZhIeRpUFU6xUbxPAY7KxwYj3ZKP6E7t6yP0YJVzHYb86sfQ
fpAoksWY7YigNTIE668QaPx+qLjK9Lf80pZ+PQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="LoXuaIqG3MVRoPESlIGtJSY/TmBelkt5tZq5mHYD14k="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2192)
`protect data_block
cF7xdgPUmADCFQKU4I+f/m4Wa8n5VaFnGpq4TIuykzQ8xq8rFO838fa0E1QP3Dtg955EWF/7pAkq
vRmPKoxvCbSgF29Av/CXiIKO0Psfx/AcRZTBiRYqy+98jw3maGpcVWZULF9z9UJQVa14B8DCkNOl
RhmAXB/oBDzSnlsjX2P2s3mUnYxlM4XWpHFaPxlsVCcS6qwBcK8s+JtgePUIOet6XGwRL9He3Vlp
tpcKz5i7Qs7Ypd1Tj7C5NIxdSgG8B/bJTpLAYame2Mj+LT9G+dLKfwlrVy16mN0xaQu58rW91AX0
XSAj+f1AzjeBPVHY1sk6ONZNqP81jz1eTW/KSNm6eHPI7EDpbsAeixuq8AnFZEv2CIWo0rWqo4YW
oRcD/4GnFS59Jra/feKV5/izqjYWMe7r4jQUQ87QtKgWSZx34VB/onOMJMJWNoATrqT+MrJIGBBq
JFyi5Ovivm1bcEBVLJuqUz1+p4M8VZL114zoSbDb5J9pqjUpskbZXB+dhtbpkTCnukwXikZ5yepk
D4gzLBYOsjU+E2Ls3U6/q0m1UIT0vgCP1ti81wKllQXXzNHY4HGo0J8Dhc4vpKq5RmA9UKJwv72O
00NORhptr8pfjS4iKLF03dioCfR2i6Iy6W4Qput8fU4JKTLXWwRLOfFRt9SqIitl/tmIE5kp7dmI
r/gkX+Fuj6+1JZYEyce22nP/D3Ug8GvhzmUd3gN8DY7IhJa10e8WDA4OT8ZhTgpH/ZS9TnlOnZxw
pqaZ0A+IZRvi+DtIkNrXjyJHVoQ4at1psPRKbW7arLR6JLvzmSLFlcLDct0D5Eh+PTGFVrSwqQWm
XF1vxvdI4jPJhhXcw/2O2AKOgXkMEwGZJkQKqGrz6mDimN7NDD9AGbgAf0d3Beyci9ezpqAkyk5/
ecz7XETf+iV4FsedqmYoztgrjlmo/YQwZ56vh1u+kCwTbllZPTgc7jcBOSxnzJ3C8eHJ2YocGDsw
V+XXYcfw1F10eLGE1wMrPln84RTtUWkghVNxJa7eSCyM0fBdtf82OzjCLuBuO09Ohi4bVFd5CHAF
mknc2dOG96tqW//a29axOk5bDjnbuEe5jrhrwg/wHfyvTbTxXscOn2DGL4hgON7f+nmO5lviK5Mq
5iCIOwMB0+xQJ68wwNvFecORL/cFPY8NTtC1Yjt3A+11IR8WiPrBsHwoTXAoJZ27kQnkI17qeMNf
s2VjjpaAeEFq7fiSEPdmouEhI0bxWwtkU/XFO/WH37efJA94FCrMRlsNz8H2ZHVhWia2ILnxynP9
JXBM5j6mpsy4Dkx0ktuOsqWFqTVzKqJtIdI2VYTWireg71//cYW+HisbxfWNYYQ3PwNNQHuqB95P
rrFFihM3+tInIoFYFxBj1rXv4tzzQxjfvSUU1QgIp64OZSjE5mEA6T4zgTwv0HdRosWv2r3UEndJ
QwvevhuyDTdu77IrqO/wSBo/9Eb5aJjR2DuKRGhAJU4rxU80rZaRsVgvFU4FUKzJaqswKg8XO35T
dbk+1+IYGzd0EPYGXa7DnhzI8LeUexZQ9PoH7yjur/uVUpuq3NwoGVbAyHbLx78Xugf+p7xKaznY
iBGyF6OHQjbGjpboj/Nw6V7tBr+t4GwZwhVTPk6zEwSjH6Ed732Izeb2KWGVY/Q57Jy4M7O7q2Mj
d+4IR66npyIu/y7x2dnIlYE6K/WtC3J85eJ0x4xoEl9gmna3kF0HwMsiacocQN5AG8BSaEB6WSkb
TB6Nitv0ANhsSCcSKx7FMHUw2BengW+SAbCYiuvQpzU+AipGjjwrtsmpVK0hhD5p6gNLBuAExyE7
JWK+5mV8EBi5ayu1TEoii4MVVTXhrs5WiNAPg/P0LHbjuUYr77iClN7HRuyikhOykM0v3Zuv/aBi
K2F+pcA0n8FWsn1yJ45yksvN5gt48BQVpHXBtuD5kyPOHpW1J0Mbjxk8DuK6Ajc2jot8VKXrO5wD
s7KN71wM4i/MKSRaQkiAbGY72A62Fl4IJZ++wQp1Ij30F56Wbspz0KIZ3GdHi0GcRL5XaS9a/YV0
ObFvO0jPB4vyl5l1Q8gZCfP+PqNWPy0dTLQfOni3Fy4suNW7ltH1JmO8t8lXuqfjeCdFRNLuv0jU
oBOC+RqW3YEc6zajNN5HhI+w855d96vQTsPQIKgPxhTEHx+jAIEBzcph8lz/1vWprbmVJYdVNdG0
PiPrmhu/UZRJaa6Vlnebnf8dybrEfa2khA6afYmPAnb+226PI+/YrcXe3/4adQD9nHNi/aXuEPaE
G9cXArIT3VTCaOtg7yjwmUkFcayPms77aQOwlXjEDAJoDrCLR6Nwle0LJPgja8TOi6GNAKewcgvJ
jymZ9CA6JbeGzDEGnZQhIGhj9LxOlZM1C6V5muPBQlSIW64+T+FEtUQjkeNSRrAV3FKwvPqMERd7
ENdZ5CgHW6QZfMcInU4ImfsteNwqKzgdKFgu7007ar6wfD4SQ7RZY/XIlNVFCD5ocyM4u2gfGAHZ
KottxhkimxvCeHCdqDYs3omMGme/okf4SgAixR+0N/rfz7pwniK9MLQtLcwauTWwlUMAFxlEK7z5
w7O/8PhaWzcMxWom+Br30ue17lWgM6W2UtuVXmG5/rndSXc+1+5e4TL+Doh37qRJhzQUhJnYyGnY
eqzsfO615ILtJLjVkNYAWBYKRXf2GOG9S/mN7MsLxeTtcM4yxRN+KMDMclkQZRMD4DLEGhfrLzls
+2b4B1IODHkYu5wJ3F/j6QU//80FGNifN82KHLS3cKBRSlOt6eG9f7syH2LJIc5PqJ0NNLxG/m4k
XJLn/EyeastEf9avS7B/LPZRH2hLwBuPf6OxTLbvphFLjhZp+0G0E6NMEd3IcRH+G7BMUxZPYo4c
gK8DSP/tNhkADj5xsjsW5m78VxaJBOatLGQ=
`protect end_protected
