--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
WPzPMSm89iyljDe2K5K9lGosqJVqnwCX6EChW4fjySBue9P3UuAROUB5luYd9mACVyacX+J1cTSG
h+Ir+jd6AxcK/OyQ8MNxVE3qWYiqcYIH3nas7fk3c82oWEA7jFJWt5Yw81Wezc2oDkMSkpjT6fB6
lX/ZReJfTrWneuHkMgUxEZ1a4252/e3EiffULfyw702tW1/shc58w92/bgloGnf2Tp9sb/cg5L42
bnEvimclkZCbIDKXED8SVQVhZGCOl6saohNFVWlYXAyLYAm/ARQlkCrLMhnO+ZEzCuzS/kZDsH1K
PgeYxmpicBsScoXozCcXcsG4QQv0XCiA685V+g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="h5WwKxQzeELKLRVqV7nUPprRC1y084b7Fx2BeD1OVHg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
s8EoQ98ZBHQ2lwnWeBQJzXlh/IIDRfX7JVcrGQsvZ/YyeXVU5PKtxaaAB6w2j5Od3WH+hUMS5YR+
H2HEcRa3H5ITVLLu8DXGcpvZhX2sK0gk3eQqxc4sL1wQwGNg2n8Z9ap0TP9AWwYoVVlH4Wc+0pW1
a65X67VFNxwaoTqJryKqa059tIQeRw9Ho5GBOx3QPGpbxVsbUHPB9BHOuWhvjUDExXDrM97eWwzi
b9A9cjmCoGStnGx10Pn7kbuHbw65tomCMAgHRyYJT03PJ6M8ZA6SyN1Slm9l0caFIv5R4cP9W6v3
861j2j84FtlGfVsnPcDqnS5UN/H5m/Y3RF4FzA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="/dWTx5toOiOZ8qLUWtSvC3D+TNPjx0s0uy22qDUydOk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7632)
`protect data_block
L0SI5ylYY3SrOob+pwxAgEX97jVSlY2Y7H9nChjK0TDE6qzhvI5HWoaMWtUUCB0UZ4WSa2dj6KoN
wjRa0lPcXVXohyABdv09FudWgAn6NcjIycvwuz8FcpNr3+9g2fFoltz4xXS+PZHIQtqgrW9+qvGT
+skNBzaWGJzqVNSpaE9EFkh78E9VWCMGYGzdiN0Q1KqzKh8ekvxPVX+XXl6tLLjhYmFOnIvc+qtV
K85vQuLWrFQQuQXpdF5yKU8WTzRSC3giiT/jj24o3sBh+s27+EaD90gnnykF/KO7GrngOFgOSnMe
vUQ1YqatGky/1A3gu6RCJrO2+D6HChvFWJV4ImuOXrgtz6oWY197ONaE+BPUgEelisCheplv9Bvc
rR1MQz4bQfCXU8iIoXV+dnK6DSVVxBEA9YdjB+DZjk7rncwGYqIwl15nAffVW8378DJ4SKa9phHy
TQz8dIBr7QtRZMSAtP8nyT8BI/ptwalhoakqWs+KHXwluu35A7j94slGbjYA8L9NGeZYcUKep2rR
ZfGCawEaNfpVWWZ8s/7w9VjKnFzEk9TF4V9pup8Vi4AEEXkMqAQfMUvVgp0dngTj+m5aEonvKrHh
CaghdzcU+x+SwwSkLO3rIKTLKymxiUU5MxMxYTlSGdb+NJwzvSIXyGuUbZhy7T8wp+lndlEV8n4e
H5jIz8t0eaUKoRIDbZsbrgfwFFGlqZzFJa5FVW7yGDTWVWhqY00n10Q3UEYP2Kbb1UBO2on8eIHN
V2w0stQqHBeXXQsgQE0ovGTY02ZPgGdhmcCJDRIzVjlbsvkwrTt6SAHmFJZFgGmPnKX1KA9wPUyl
7+RDrBeeamR6+Up3l+YHE3UGAOxbNgOToZ00Q6azZaMI5cYspmmyftKaxUwvNZVppQEptVZUjPcx
S2lx9dhVlso98auHSkkHiITw8dyj7J2j8D2Fkm8BftSPXVfW5IPmF7nGPeErzaSn8fk/F4K6+q99
0xDYMfNC0mxnLb22C4ekCBOPzCgXpu08NfqSVc9MFS+6vx7cFes0PVD68DpEgvXVelDHmq7/2bqV
OOqc30lSjlOrxdMiwyMlF5SDn5K80p4dWlkXrvoJp0lPj9e+f+S/wzr8dLv99GrQRCmXmunDUP2E
m97qBKWhDEAqzSYvXHXeQV/QV6jJIY3dA1Z4ghEbLukj95pznaP/z/oGaYIbBP7R2p9PAnDyUQxB
KbPi26WHZB2EChwj4gmKPQL8hZd2+c51RT1lGMtrAmWMRI0cqQJblQZyVQty0NaD5tRm+6xhnO3o
kEKFMmB4Z/kNF7/i3J8lfquiDBB39/5543dB0w4MaLUgKpFMVdeDWgYMyu5eH3wCzSSlPRgC9l5N
GNEwBJBUO8VsBsy68h18XEOnzSVZd+J8FsEDeY+GFWgg3J+mk0igD/YPBkUQC0pK3C1zNqYiZdiB
/zCjCxIs9vOttnXQIfQzOxBcJgmf7rHzpEw5HF1VON7Xh1hq+3j/3BCmHoz1ry9EC6Ba6KBE38Pd
xHOrFf7FL8wDBsVntxCkBZaYSEtktxozDqPxwFIFNDmj/pIpdozkcvC/AawJ4aNlFQzeZM39YU6l
ylpXACYgzNWzCQiAv7HQG6+dC3Pnsp3mV9lX847Hzo7Ds8RUnWQ9VNWz2Tq+20xhmxWdxhogBlxH
Xenslpau5gnDICvyLeF6OnomSG1RyWeR+6B+5z02QPk69wvI0JwQwMbMPq1ALrn84z6keBQoj4uY
Zg8aQaBKuioGmtYjXEEdL1Loau0LTJzydtbd0EFR+HDldhxjyCgkfkipYHg5HFyAW8VaWAcR8Zwc
M9FvZ6WiFMieukSC8g4AXMgwawYn8dWwIPXa9XAbk3wdChv9cl+gDMk2fu405WAKP3pp1AxGLJE1
Yl1TuMFAPd/fgkCw5oO8rDkOwByMUj2OdLJAV2ij/HvaBLLtvCTHxOV5C/hLcTEgd/t18S1eD1/c
p/NWTPzakt8b/cjjzE4Rzi1pLLrnmhvaihzo/gPRx2uM5YFOFvNYETE//aAM2NA5+ZM9ZIutsUl2
GOJi3Q6DK/chNdaJj53/Y6Bs9KKCxW+Idpu1IWI9IvcacJQuKD7OBbiyR374n5Y9fuImSBSGFEMS
K3IxCMcFx+SocNkkw0LDD1H3QEIrfzZdeKMASjdgl1vMpjxiScR9K//BbHC7P+Tm6gRr3ZJb1X2D
s/4UflzRWV32uxN4yPGEeor8vQV7G2zm73ct743pwPXZx8ZkFWnutlbz2AusuMaYYHMqUrRWSdT+
rujGHPpU+s+PJuup5GkBZpJ+NjINMCRYuyfikNL9ZWWquVa7FBRUnVK5+wVwQ1Zrr7N5MXBdBvdU
u9l8CpdG24KBUi4ggnxeSJXJJLvn/GcnKDOfLYAVgXFmHp4XaU4zAAEAZ6L9oPOJs4/ZOaHx34e+
GOHFsAQNgdqfzXRu8S4jmwN6tLSTG5+wcOY8GajP8X99JudM/4wa8BvYWVEFOfJdI9Y/6BorXh11
DxJxzV0KGpPQPXyBH7oolko4GQ4VFA6lqP9waS72m49rFpFtxzrqYUBeOINmmSU1FPfyH1HGNEPN
KLWC1GvekwWRX93KtOZNtaTt36kDQ5LjRNzGOSjclz0uIc2INPffE7BjdhhwTwM7Al1uoRk0XY+w
FzziqYU3SV0o14kRNbByv55pW7gwFf9xZZtEh8cD7IlwbVSljcoJ+ibn94TXOtNiS275NT25Kvld
3VqZM+VF4d+eYYtIUTeUGUi/sclCe+XHg0FtUvWJ1X2RmFFipks738rp1WUWTwkJsKQCY2a2v5md
VXI/vz+hhkLKKYVezKp8JghcfjKgpVj7JHOYJ1wcyVqIBRC3bmLC/OYjuqdjUPPDiTUVGkwxIuus
kO/2R/l4DdZXt/IgtijLp+gK4gZkAMCNAy4NWvkg9RtoxQuGBTILOiU7s/5hHo1Gn0sWlhIVFbG0
XyaRwM25K1BiQW0N92bViX1p7cgcBstvczEniDpZ+SnBrACjS9qjWRMnU2oslE5cSpXRtQ/+oOl9
mcUdh6bBZe9tr3Ge5pF3B+2X92czYIqNtgxRbH6NVeF8I0Yvwjtc5JW8eKb9yiItMWZE99Eyw7DE
q54UB/HaF/ZpYtvS7+rlThQgEL5qdgXsPlYPKnAvA7BHCDVWaOIfcj8ImHzPkIbQFZCDnkMYTu/+
OcmUeLy62KprH9AAbPX25My7aFlhLYeA6+ds2aK0CDEfNgQpNP6mVw98NWnbazZsErzh33363/9d
Lg1a4FJL+S2AYSiiCAUlzgt1Cc8vfre+9aVXRyzKVVkDtWwKRiouOcSWyMVgnAps96pSXXU73p/N
zg2iR08TWNvnhrn82ZqGdgyiXx8H2rC4PvIjGBQY5UcOG9XpWGLlGYboZ2Nc1W/upOsTUh8yu+ps
K7/JecN4+QLO8T4FidNQhvS3b1ApktbxZ2d3WnyD1vvHM4TG0GyBrI4o1YvJ7IbICp62ifA89CUn
yOg2fJ+lHbcltxMW8wLr8fwjOfelLNXpNfwrUTmxGDmIA+XSueQT2gjtj0A2cpzDOZCxcer8CCI0
CgWgoMP3XxdchDq57yK5P+phamEXz4ayWnxnbV/MLz/kMPzxVo5l2oensBv+gAX4u2aOpbnHIxZZ
u+AX50GAsGuAB/1rsHSQkr60z5DyiEXozK+aDrksIsbDCj0fqWkiXyj6VAsvrhgdv+7k6V6X3M/A
4cefnDy1dcczGMMMqpRrun+PwFsqRz1rSWx8sMJm4pSlew36nmdBbQsKpVJ2q/AvHzLfk9mueWxp
xXkeTI135rCoEDcgMpE5yk1b4V9WGc1QukPwBrXNa8LC+42hsFf3qkX2rGxSeujkuZMlB1OC8GkQ
fBv4/cW5DGBayUI+7jwikafcphnasj0QCbWUd0z09Os6CGzUUZSp2TYV5rzmY0rWoMOtlJm/JKM/
3yeLQS6GjRYFjKiO9jg2ff9y2JoEfXbpBXHfntxElOYr/sLJNzihQnhz8i4VrY56vrV3rt2piVto
lm0uJVT8TPyw19I+r745SwEWq+VVY36lc/P2OCQgTPwrVRsiieNHBxYcN1UgsuB2jlEV0H4eqvEI
BNJ5/Qi+8HYYxJFnRtzZ5kJa0ecqraMjNAL0uZLzUosd9d0vb/o8Xr4q6V8FpCYfqBOau0y61nvc
BRk1ucz6VG30YyY4eD/+aIN6SmR0tDL6Bjw0mZX8F6gjmFwunv9GcxPJJTTPRkdHFjE6a0qC1pWy
THBs30zYz7iiqJq8rC2nhQjFyQ38Ny/tUJJqmv/me0kOVrPCqcckssqMJcOWczKh9k8nKMCkmbjB
q00bftek47XQKHJS6x3mLN0m1zWyMtr+MgfW+khTrkrIOT/9494OzigoetjKggv0xeFmL+Vtvctp
OqaK7m2HKLlfTBIY9ODiJC9+AWfDAdgovvYnvC2l4FhfjwVsRIhSpDavXtSJa+wbAJ7RFqJmfGQ3
H8VQROaM0GUg0VPvNHQzYrOwrprlueEDLc6wpY3nNEGHfFWC8DM2cg2Psf3Y1luFw5qOryGBp0Ai
5d1AMNpzaKC1oaJLh1lZRHd5zqRfgZnPxPvbEdSEzKy/9+0RUcFXalcWkh1oKE4FJeZMjVeC4ClF
6awHS6U9nOQ8knd2kApN2aLayEd9icioz0W6vvWgmfb0g2Ca+FEloev3fgmIzyk5k3oyeGtHRe+P
hZFc/CrhQjeSBmHs3RotBD/I5qEa2UTMTwmk6l4xn/FWi3hfYTK59aWKwaLLCrJg5AZ14BEx+hH3
3lL3GJ7bd7xnRtBsyWIOfIRty2z6QmzlNX5dKU/3GMTi3WvJzMN20PSyuQ/gAq7FMLnJtm+CeJcN
B76LmFfDJB8/Nhhv/2ZjTrhzCpzH4xCg4+c8HEZy7TDm7Lc/tzJAbqgmOBSqNp2Czkj/soNo//kI
5gCU+kTrmCAzPch9VvaCZz3NhqVBh7Cuai9yWiC0nm5MJJcqKUWrWHz2BVpK38s9ni8lru2oz/vT
6rq5F4BxoPyFVxuK8Qciq5dAqnChFg1AQtKiwaD3wreJ+zmPE8uEpwuebVKKstMOu8Cl6Bs3DsPh
z7ASf3Vo2dszdGZ8Fd5JVXdjcOvKc+OODISQW4IbtzwrQxchmUOyGoyCbPn0n+CwylSEPTkqJIOn
PQ2PuUwAijL8eaBXfs0HzTOFz7QmyYjlSrl9AkBJ3PNF0Bos5PhGeh/sJoQfNZ+5qwDN7RanhcHt
YPuKzdwMA24LGPcLVfDpu5Zg34RIzwgGTkVf0bEg870i2A6CN4YfcG0NaGlp3IAB7uTYEIfj+Hxz
saEQfSASFGe+qRRMfqbzkQ4SQa1mv0w5JIbm14TZeguH8LZjIS5PgKx6I5RCTnshk5cl9DDTO7uG
XOjXB4sbDn2OsBOKp9PuMBekEmeGdHM2ozR+iu1IULc73exzEpyhqIYYNRNHvzvIy3AGOQF4uBgy
JsI7ROTe2oyf/hj6PmXG3HQJjtj7cLLhzgnUfVuJGJMVP9s2hc8J6/7f5BVhCGV0t0q6890bKY6k
HqOsNoc6xOs+paiMDZxG31kIsAaA83RYpwBvw/54mhbeD28RHj94HVgSwbpbP3pAIVqJZW2nBuks
7Pw9k9ESmZb2BQkVU5DcpNo2hehZxitpRhvuEUM8YkbY72baHHjDqZ3BEZJkYFzFZUR0IrnouRfN
FnI9PEyybzdWLTYI5z24paXUvX0jLdOxIybEaIbqR+JJpOuszS8TLBuFOImd78iKTxpcVS3SgIIE
0zvVCjB2Xl7bNI/xLGtJpVQAH/F+mFZ72gFNAkOR/CINd8mDeuSLjndlFomA5HjfjgBJg+Ve7ccq
/vNq5mVgkV6OH/Q5bCjMgil0sFmqXmUQ3EmUD4Sk1L5A1agXF1bTBup1iYscUhbUMccz/SIcx4Xm
W32iwnVLp42umGV4iDanOEm/I0GQ5odEqzWo96TawhJzdCZsTlAlGmw12YkCLpqMbeMorPsjeQ3s
hutds3hdex3M//fLo/YBMFsnD7+BIKd7xpsZt3uIKZ9OsqvH0nijRqKak72OyOUqCv+9hgz6Wuus
mpVgv1cA6IaMAe/xK9ATC6Kdslo2HMMK3tYehcmOpap2vcSrt6HONuj6KJB7kb8l3oU6NLutuK0N
JnVo7tVQ/hAQ3dL1mx5oOXusnU88dxWwXKOh0qIIRc14YAv6lm/SBtO6Lhs1vJgFN2fHRaw1jCiz
2LOLdp22UL+n+64vbb6/Q3t43y1N1oRniTQG2nsKsjyRB3pSe0kud4nwffCWeO91qXYaMfnxvXkq
+BqAtYL4TUvAGmUBSEzkgzGy6xfJ4Y0vEZPJR6Pl+VlnAg9E/3LZEAiZ9vWEQ+pcdgQgzOd4pGk6
iZM95vsHaD9g45aeg0Bsf6xCQghsoVnyaL0JmIWsEAvR8onwW80qpj8qNpPWNMJkrKMXOJIzpNHe
gFA/idsP1am4pmSGYEVnEbmBVlfYIJH/rkyDpcMQBvxiaREY3AKYlF7oQJJz8xIfFsgBYscUajFO
8+dq6dxFIB0Q9q0Qe9ppxLQCO/xE3GAIEof/4lxSJTbVTZYNClr7VgpKkm20EgBNkH9mhPoMgNVE
vM5q0R3EtjbCHMHJcBIkQhqzU1LCAjBDcJuZfSPaWoIa77trMieHbMeDzgetbe9nwb2yRDeEn4uL
+TRPmCPcMQ4sbRWJdachBtAzfa/N1S0qoHnJGZeMEoYrtDODMJcXcWObktjat77ndlEvBSfgeqSQ
gLtgv0lgMCJQPZbqK4ylDxGuZhgeAe5TzKTvtw7XLzrjyHfFQfTC6ZJRr7PBvqL7PKHk2//90Vpu
MwRWpQ9BH4+f7WUnAXWKUxpLk6tcje2/wfWFXEK/IJjsOAEctNCcHsXslXHhl62x9fm4lRA/ep1i
XQqds7xf2sLwLBOK8vzcKFfjC0QzVZa/KFaairXQ2IPmqtTrsrCelRMLmGejo3rhJ1V/epyUrix9
bv3+HOcqnwqDzGZlQDhb2Pe80lfhUoPsA4eAKfc53rVP5q45FLT+FpL9xFcpmnRL0J3xtiKqEQZm
HRcZPWUrLhUvXCbjvegQTlKbtB8Q5wcY5CQHxWL+ffx+YR71kw4GWzNuCxgIPwk4yJJVwZVDZdS7
uykjihM7JxQvyopz1GWd16lA1E4WAA2mUQA5zRf2vFobLpaZgLnpI9VDjVgiZzgG2pD4Qjq1GKLx
ou+eTcyuO3PBrPJsk973/RSN10LflS5/q/F4y5Oz2TjK+o7yNIq40V39+D915tNKwrkzWfDpPx/S
fFXNcPHofvvGDShpN8HSLWghqyC4okp3Z5eWQHkv63I3INnnzemEK3Fx553bk9cynd1a/C5NsA2F
wi/Z2n3ofHXt1Gq3amNcY3YvH+KxF8AlqcnGc6JFEMM5hFM4SYjcyImH8ip37eWZPQM7yOl80Hf7
ZfLtKm1ZbNRrotksgxTn8lF89QW/aUOYH99BUGyGh8E6AqB7p8BJI1r+vS6riJsKOqWpnoieFPmE
Lr5MC9kjv/mUD0LtNhSQHPSqDDlbj6562CSzTdKuQLrZNYY8Ux3iR17MAZP2tyRJ/f6v1TvXvu3m
x6FkqTlro5lcO1NEfqCwKddfVhNA/3j2uhPo26OMITsfo6H2TKAvLavJmgaVazkd7o9lvIVQxsUd
EdeyTvE1qktSVRxypnfkmcaDJ58ZBzlPPfxtqYkzzvl++fFXsX0claLaXIf3aw1g6HjBFSAYMEJG
zO7Jg86AwpxZ08VXDspI08fUh3t4+TOhDeq6C/JjevH/wxnkMj0okj8WuSwpG6o1EwrsU9bWENGg
URicttmauPcTC4Afyif7n4gkbE6lc6Czz4A+sUiVdwwgvfjqMmoqArMmQWz6Z1Tg7hQFgh0oNDmR
XLa4PUPZkiqu5AMVRwmYS4XGVK1Ja3nfKWgWcKluz+S7ces3CuW8nsJhrj/wUdGXMjPATFuOjG+o
Ccp9oKwiaPlb53FkTcvXL7DeiNTs76ZasVRQZBfFIbZqFuTW4qQobuudKtAOHi00j7MlxYvcEnO6
RjDR5lQ3BJxb7huRfhZNGPpYYG8upTnNDvn9T+XyDfJU+sVmN4r4rNmX4oLInzj3lFFUdcezm8hm
pMpwyS+N2Gp4lwidtXTYgLaLoYKwJbZTuqjC83BmYkT58hLpkccWEwAQv7J4D3x/GkXuG1kuvbHD
DJ6I5jjWmFAIs6719WHk+cLNUFv8GA/T0aWPa/JBj/NUN/lJw7QnF/i38WoHpEafO4EkIKoIhqkB
Y806yu1+GRdkt4CQyawtzZF5WbQc4q5FCmI0LZfx3pc00u9blcVuUXDibkzZg4Y4HLFNxBVq8Lxy
/Qlif3KMWoKqogRBH/BsYcd8nfDF3wtsuA/jCM3Xuy59/qRM6uTo4SGqlOa6rapvyddzDMt3JcfO
ian5DUTYDPCd6bWGGoyT8Hgiv3GDfbMhG/WVmeMIWrl+KDZcEZLu9tDi7Jq+A3VnFElIu9B8Jtvk
EkIvvDMI6ehscTbYYNceb3ItFrx/m1ddc25lK5/2jdw2rfihPUgND9lVIu93RKwgej9ifigN1RCt
ukUnKqQdbESNcedUmGJn7EYsRChVP0qdaquj/nCXPcNNHVBJiJku8wXUExKuY0qiD7hYB9yJw8mS
rUU7jpPcNYiNJGsYdCjZXiHDgn+g99mOzoYEJJXZSjb7W2g8OBN50smY3454EL3e7Zu+QAABe0ZE
pkkBiMU4y1nsRS7VArPan3KscCtmcv9upnpFQYCMHmQ6MwDBeD4lxZzXwv5NwtZj0DAc8k3YqmPs
iSWNYds4x51cBAeY7cB6dII4ryA5t6pZYweCSyhLzFkDh4eQ5pQ6UqorSd3FbVpLupDeIXxxn/KV
Oo6kCW37fFOMiRSN77SVsjAVcSDMUTfTzQGZFz2CS7v07J1B5QSeFFUFrYDLQv1oc0aVDdTfD9bC
Bz1UzUZnU8JAouP7MmgIaozZqhG1Pxc4wTevbwcTCmGuHD7tZIOMm1kqTU8Vsxz/mFIhAsw5WLEj
v3s+/7/qSt1kkab39iGikQaX4+lijXaOn0sFmKtbwoYwTovRIcE4rlovP8WRxTR56C3+CIGKiX7y
ZSIWaG80857F2xqkV5KNSlOpBUfz0r4VVW4NNLm00Leuy/kiZFK0fJO0ReGu0v893kFO1t5fCZQx
rQe581yr42NYqqV/6l2RULHvEhIxlieWXCwT52Gw5tBjzeqj9FSMPv0EZVhdF8BQcJSraZm0gQUk
xHdrhnlLzmB3jQg86XhIC0BxCQ7+eSDKw+mPaDyaNu3YeJKGSHDjXqMtVpISyIaPiSNNwNEfjGaN
g1eRhGfh8jER3z5NqhPM6b0Kqi5NwpSE299bBlFWnEAbA8abvuir6UJ75XoBoEp1GAlP8mrgtNGI
K56bGEN+pveoPkLYcSdR8xeQHjMrfZa0MMkmb6Gqy1Hcs+/bGffE0bwNz2iZIM/30cKYWq/y9pll
wPe/PqPqd9K+DIiiEIFYd0TvQ29cKrvstdZcMfOu99+7tVWQ72Bq7GGToh0DSC2poDhIjf92sbt5
vVqR6V5FP3UX51sWrsyqlWDiCnvaOb0m4qwMGhribGZfpjxBJA61HbkMsvY2q/CmGau/85PsIQwQ
NS7teGJ9Tv8jRxTGC+A73K0nA8UmiM2dmu4ANyKjiZnaAaNKPtpMvBrHcDL4vZDcMduPWoq/Hk/t
6ijxSsHqpxCFu6Rp/mW8rDJ3jwTxL4BxR2bfy0e6Dgai7gPuyk991eFdQzL3WqyCnGegZHtbpcdQ
PZkoqQ+pZEtpIAmEwNMougW5mgA2rKjevx3Yn7K6IMHGwihJD6nzvlCmQpD+5igo0Drq+1hOrUji
qXEHIXZ+npQrv43DXBf9WM17ewrWHu+jK8LNEjsN8R6sCfq10RnUwri37Ejf/uS37eoqXr6b3u0M
8xWH/31VyAKfSl/NGErc8Hyaf1EMPgnI07V/5TEE18KLheRsu47ZOn22pkvt8/cLMLnHrRxgwRXy
Xz8nbG0s7FqSshxHgsG5ahOpttjUoLbT/4W6KiF6/86CHzunk1sku7hE1hLMejSa4X0STmwn6Uxv
5SBfQkclB91Sh2Y4daXSlZtuxAwW+qHE+dQXVaMShD/wV3PsBNIpsoDsT2YX3bWY4hbq
`protect end_protected
