--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
XhMLKAOiuQgtaD7xC6vD4UKedNtpxM7j3FDzc21WDYN4kBByOxaJAS1kP1k+DbzgoC9CZewXoa9C
6SvdY8ZyjvvA1jd3o3Z5fqzE4LGqA0ssNr6O1IQwkrzOP7Dq9BQ2UFATCR2v3CMsmKBmS+Ms06EL
EyFH6ObPcoYUnVCLcUN9RfdSilp6wXXV+ClsF8OC4PebNVIBmH800N5vujj24N2eHKP0ucp6plpB
dwDl9hQFyDCC7pKFxhlnxIw29mvS/1At1251GrvZM85JoRSGnFFv2G0yefP+VoHggVCWuQ1GQGFn
IH2o7PGK/kaAQZ8nHCDauZTI/Gzgo05E2L+sew==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="mETCq3Vx58pYrkvLhEnNm1zEPqSmc1osSkDaDVHss9Q="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
eJNsLCfqtJSQ8tD1WL4U2dN76L8WZeo+KcOYuXaA/dGAKUe9Pr2vG+IvfUC6a88FvyAj9fGjUwvm
51jL/cYT8Jd38EzbD2TXN99Dp+r2xYqfj5FVn6x1+z9SBBTFNLnu2b1EHRPv7kO2LyQ1m6Z2/Eea
FvOBd8UToKwhqEFPXa0VoqduDsVpY/U4CkaiTa0JT5nicl/tuJH2g0Noa9ylfDYMLSof9Hm7CdnZ
8GKcrU2J78Wmtr/jg1NKlj7Uj7Y7wVjIHG9LrVcwlirwnsCvIEl4QAaV1ALYgp0qamIza1thNTeS
m+Rxx82RlJIkXl2sngp3FHaeN65WF99/jAUuCQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="UUEBkX9jvx9sulLLlO8zmQ1WTT4HWHm3FNpWD51QjuA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2544)
`protect data_block
qJXirlgzXtFEmd9muoubU3ZKpz1STpvb/bc1eIzVBSk0Sp94oIP6OpKlzvdtmRJv/y4JuODa1AV0
b3bNg3m+ZjWQHZPZLi3lGjleyaihW62iGJbGXWmsy9ZYetz0MTwTX1LJXgAnujr/5k+peQ9X9iCG
5th8Ju6MfeVmTchZOYjZhhKUq5aSylQcuEJ9i/5pmCo4OhYhP2duHg/LLX0O3zEPMjwen/jr8QEU
WKupeTdqOCJ2YnocDD+ohLW/4nGwbjMHKtYZwx1cfioc75YR1yvS7AfkSY7dBv7YYvy0lRm2gVni
KGAfnovM372l0onHliXpsY5uwl3bPH+38UjjXeGgYTq064IGlRNjooxrVjFbnxWguKXY85hWSa7y
NKMmOk5T2GON3H2JNYzWYVONfbgJV2x1ppY50bjHh6WY7XWLY4W+R4xB8tbBNOJjtTtdQ+sVfhCQ
DTSW+cymuIesaMS9lvOYbBej8JpPQrhs4HPrefZAVLTf8Msb143XX9ZoylYrO22BJiVgzYWE+t+o
syIudtMRPOtaFWxAizjWQ2ZMZ/S9s4ycy0512/AJqivtRnTYziZByFmznfuBKsmgW4TMeZukUHs4
in6K4HGMsLMGPkETeRur9BPzgMgm02NDeN25BmILM7PsygACU17htwkG0CzZWzictkiSWn5uuvC6
Vai9Vnmh+ZzYQXsSvyxBY9kKcxgcD289nXueAg83+eF3RL6zythB/dVUjUAsslGct5nYJi5X3FOB
ChSESYWha66rNt01zzwdQAKuYtlt/AuCI8PG8u+IdihffLFj1gA7gueGxglUBNoETKQl5MDurlzP
a+pPv7bu0ExDh5D2ORKRlpm5CRNxA6SnY6yC4/IcUz7PEbuSL2qmocoaEIHWlow1ZbmsTs3CE0L/
vMh3uIXIUoXtpMtq2T8u1okD1w4838dTDlTR0gizvkb9eHuJvAcjv9WRFq6RE1MYHXl0yOCviYzn
qpMHd9Tivij6bKfTGGaCBKDlZTgw6FMQeDnFihue2RpazhQ+fQkpAmtAbd1cut/FkKqeqLY7dGVJ
AkrcvXXUvQqbGU2sq59CmHkbaY46iFkrXKZTIdq4anU1q1Pmewg+MZVfjDnjPQrStnXU0uYKzC8K
OhK2Dt2U3oa8lsjzjzPWvb1QC699FCt8DPQYIzuMGv5zBDDOPu0Hvqz5ZWbsliuOPhCocwbt8Jfc
txYdfdSekVpAod61tSINyCCecS+yc/mgUFi5xOw7MI/oFEBmqob82opokarOz+wEeHVAYyQ84DNY
l9NrgupDsvRik6tV0xarruhfY3Ib52oiraj7HAy1g3dr70wrTg0etF4gnyZQ8cUj95zpWKAgJsSl
HHGyks/CqRwES1mZcBvK4ph2dMcO6sxZlKhjLG2x9Nz/8AkLBGWNNzqxcgCZzM1PIH6nUdlqqLyo
UnlP/sOd1dM45E+ha7MzmXRL2PZuDGPL1yGrKlWZpY0Shv/vE64TuR/aI34uip1lz2RmcJQ4xpRn
/qE7vKZj7HTmCN1Itbsr4WulE1UepB5o4U6TDtchaZhdmQtp1X1pIdeTn121MIHpjfEXB5hFMJGp
MRQxXXzPkKcZk09/zeHf66UewEeG+EHuqkh4GuT7K7UDcIr1iCkANwQR4Xgl2mOmmEE0Zqa+qOWo
9BjphMFseolQycZaYBnMlxcCepbGOg7UgA64snw5cKM/ZWMVMG515N//do/66QniIpmMuPXYDysw
uhI/tJiHZ6cGQAspL29s/uYvB1UHPNFEU8O5VL6HQflK3P/lmz515WoMCgQThmkwBhWwJ+LdXRx5
MkfwUgkqwN5X8uyCsKG3r7Emi+nBvvW+7P6L4BiXag+88CBsJOhKm0e9IKko06LghaQr+HXvfy3A
OPQ2ISNL493h9F47HO+AA1IsKlj/ubT+dCHzJiQQFTRZTyE1ViGGCbl7bpPTYx0LX39kAzBYFuXC
rLCUIArKcAD1pFykosAsezTi8fOx0OxT/j6y4ti/ZL5RIxtLImcThOzVY7nMVXBJu5QSzLY8STjc
0znJIXVGRopjvTQNS2lv4tua/DuOa99+wSgcZNfjBtAYr/wudkV3sdsdyvmmo7xugo3GDLwKjyBT
GMU6lCbWLl0OEyJrdFmp9SURgd6ksn/o9UOLaJI5nqBrDJS7E7yrv5di8XeBPTFc+vwH4HfbYPMa
GstOORRiHASbxjpxvNfZj4O/XK7YgkZfYn1udaX//Xt+Ml94Wf0Z3hS+HA4NQw833nwCrumqLK4W
wAMQHazQ9v/mycV1kgiueQ2iLcHWL0arArGudkx1k/KJnGpE6E3pYHoYr7arQTBzfBPZNW8Vd9F+
EH4noEDuz+uDWHh2i1PCU3l/MkkbJ3xn6sMT6dyC93kDOBoyjdQNU8b2Oouw74y1tD8fBsY4Vfzh
1Mar0W8jP4qlj7MfPWu8Yj6D9imn7E8wMFA2zApasmAzwg90Fr+Fl2hNnQfjXNnVVfGHGgOw1a3a
pXyirdfW1g3w6afgCkx+AM7bOLIZj7C90LRZIU0u8j101NbD75M7GWTqow554rqLTatiWgsZ83tS
/p4Fb0L5Y8t92dseajWGWP+ZvinNeQPOt2YqbfrTTsXgk82j5NNbzOkt3mW5e5d4jnb8oCnVx989
i3FIeeurnSLFuiSK3fQkrZJ99fQh7TLid9ltR1DHjSlmLuSjkA1oyHicDyBdJg1mtQZ73Y0n6Kwh
KnzuHpuEO3CRIs50KnPX/Y1fiQlM4O4THIzCcwVdvQZGVZxFcuMbrYMQkvoH91RXeGlCTN3JYRlr
UBSiBQDmqhJ2Hkz4MB7j1dXqzYJ/rBG16WL5Cxru+ghELpvOtEosbWjuICM0nxEpX/ig2SMptuoT
p4c0zqDSlBsmXKtpoxlXrsH0htlP/FvBYHvasYzzB7ZMj/E438l36hdvuoSFB0Q7GODWGAdYghgw
rOzmDc3bVFFAjMBCbMKGW+rklVhvWhUexE5JOC2pdh5depcwaDjyBMTBaMvZfSN4pLUCCX1WSZgY
PRsncbgo4njnBuCk4vUBAfb0hbc5Gw08qXS+VlJ7lRxR8twmHy/dLDL1mak/k4MOcuj7SaloeVKg
rmV0zEw1uiY2zvc8bPkikYw23YxwdAhoB/G4/bKopL9pfZwmSvA5XDXQPcg1pWZbyhF0vapVBXS9
0TeFYdv5eteFhL45avetHtq8Hr3LDMkbozTRE7DqjEoco7CMoyfVxrCPml3waWcp2T1sv6fVDRzV
/hNy161EzSSLpHlC6M5veoeil+AEEH8wfhVS4mOwhshjGwLWbXFV5f5SNbwatGTvJmQlfw679ZjB
v2TMe3DlDsSCJIVfCL0rVQuANm/CL7Fp4j6cwVKkg+zvvJKp
`protect end_protected
