--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Y2wTrxkbL0gyyhmVnoSGcn9UIteQRXgwLRI1LusapwCJ48nA32Tb0/EH3rmfRA6OOgCOX6T7J2tk
RjOD/g2knTK0ZjCYjsyo+5VJkrPzvWvVS9L/BgeJXY55pBQhkg7vQuH5UX1Z2zf+8MxVUExKMl1N
KntUS0U+S7fZ9bNAMqi07++a10/zWeWSk1HQ7EQ/Ypy3tI0japV7c6OM+xkxXxw2SmVNlvmluzih
Zl9Ya9r69/PMbqaJd35Ugp/DAJveOdqCFONan/XiSLofqZE9qQznfxhuzR4UN+RY4gvV6e4LAv92
WqumfSjLol91XOuG/ziTzXdwMulLHVh+/gbCUw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="B5SjFSI8RKDTlvDEC13wg6GH7fjtDtqikaRqs1R6DWw="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
DoIxvcPsui8bdHbaOUnkXAjxpCL6MAdDdNsXUVVwNF4wpIxZ7t8f96QV22zAkXS45U1IagwUfINM
/HiSNLpHbNNozNlczUbjBGH3tVghMK+pQkHSrv5J02UG618fK3be5tUQ9BRRVRp87bWdI6o+O86h
NU15vUkD4zwtmnc1Az1EqiEyt7yrr/FR44g1ClUOxkAZIzUfVVoS2rBbpz8E54804okVaet1r7y9
Zw0IX9lc5ooV24I90Jb5AyEKgYGKn8WgTRapK1hcgT4uBvgk96Vmd9pVV3rRlQhbn+FQ/tb7c2ny
TEFJWcdJbaE4AiywNmXqtCBk8j2aKq/A0zKMGw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="siN/10gRnNzECI+6cM5aBtUAbC91qPltjVTQ+6o/jVE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5616)
`protect data_block
uvOVtzn36VKjvkqjfSA1qrPA5cjMygluxPwpVkzbIbvqperbQP5bJtoXCwLoY2CefGJtRhj7Xpxx
cLIsTxmqhseVp7kwTR71dgUrigfvqDj+z6nYuIFzoJzbsRD7qpaSzWgNnUbIB6NPvqSZqX48pKzB
EuOdnZv9mgGhntw6HzhpfmnLTlP5UvDRNcX9OHfIGjttq7/1it+XKpXdFvkrfbx7pDY8mo51S0Ih
c9/Y5LEMSuBUOHbYqYxTnCInvYLGbXUj5YfLeBHhK+jqmi3IAjbYYK+YtCVivgX75qGLP3tLk/5c
7/M+Uc9nzEgqZCNFbAo8i+1x9jreI1H+fEg/wpIQJ5eW2fuvjROSAoiWpyIG/iIaMSxrsa+4wAWs
G3O/8kaArO3IVhuW65MI9HiDIxjTXtq39V98gjW7J2c4m9dNkrC2eaLd/+Yd6HXLZzB3wHqMDs0Z
djZ/u90xQPK5VqeXFPstGj1F3Mxi96giH68hYakYhABiZM6ZJofvYHXlKLWebbgEf3znPFrKXsUZ
LbvqeId2ObXAicenE9eDrd/cPGDGiW5CJqoBQwDtHRIJuPTX0RpnrfpF/r5jQOMU9utAtM+tdvno
rHNY4/2nV6d+sgZou0ryS2FqaHrQsVpvEPGbUnfQU90WjlHnlw8HgnNxGdBwOCVbmSmcEABK42Ym
keOPnT4CWiaUeFVf4tyRYX7bjKxcDBk+oeyNhWcmoxlP8OqmRnmmj+6pNcyaXeiXu1IVoV4Fv/CS
gchRgFki4+lEXG9/EPCQxbAdWw9oeew3tOBqy1IA/FLl/laD5EP17If1JEn+8IJpWRzjpLw8dDRV
Qtj29EZt3ym7mseJqDxk68Z/TPwPqLKUD1mFU2MDmesAC04155lzEKh/Mg0zGy/F2mEzzp3TGKM0
AG7nbWvsSATf6m6Y0LBDEYJFk+fLgjY76EUNj5FU9RF3SRyo26wBpmokXLfWMQKabLCGE5FWQGek
wTV8XrPMXd8GqIVtLdD9UPCxde5NhuJprXg0MTAmYTwhK4vjZBCgB0pEEbR4szy8gcMTN832k91q
aJfOARrljXCsyRv5SJFv9T9fiTDBxNHB6Cg3+qSlEQ3u5XEqo86nFGjaRNKdzqdnqfQNCSLxCcHp
IgasBSa3j7WsCj4eeeK0/AnA9qGShOWUhcHA9PNQ6REOHGezNStpk4CX1inf3nU199X6HH/5tgDm
5hk9EY2dtXE4V/o5Gp4kwpcqG0gd3YkLgY4tyPbsuSQq5sVa7fPnkRbTKVObD7RJnHKTlBEBF1bE
fM4up5az5pyk1vIVkmml8j6l3qG47dtfB5bdItZCTzdeUq7bkYN4Uce8dW+FjMUk2MOkzoNQeyjP
FZS8J3ZHOw2ENyY9sm4ykZimMH/XXW1HBKoKv2+DCxXc3mVLzFoXTrne9qnu4kU9TLTga0OmoLjz
pp6+vsjkWwwe+Q9VXzdCFuOmzkDVFw+RDdx1lr0sOLpw4wlTaIoNqrxTLRnwNeGAtVWnmxWdK3KA
AkfD0Nmv0WgvW6W3ftg0SfNFm328SZ3xF4vCNWE9zYH1GR+ocAVXZGVj+BTWsrM4Sa6JVfwWh1fN
+cD0sXEntxocZD+7WFW36s8FfaaF/dGWpfOVxD6cKYpm+qb3i1XNI9jmTEB1MlfidSvs8QMiT0/j
VRemeYBw1jcA5FUnnYv9+Jg1OAoE7AAqhXO4xiZQhx3+uAUgmYwTZUPe4QhVpKGz8+r5Yq3hSODJ
sBbMLYRQoLxF9bxOFLciTL4j9GyavIfYoUG6I0jIhaJ6sOoDsJKLpNdZdexVBZbA3hqoA86v//3d
0xftqOd2UtUJNlxbuhGQS2fIaLI9Y6ZLa1cMhUsmM8JtFJ7vpSEvyU4ez7ZsmNduKrnsbZav5Miz
5gbZlKOhH7xHJR8qHfOBpU2PAbe1FlPe1TKBCoiMRI6ySmiEQZCYnSzIwWM8Ulj5CwDyu2hK02UI
J+hMN9X36/3lZLbBZQeybUzElLhfmpErqrV6o1wQuboMwRLFZkk+FjNa64Vm9K+DJ1P8mPJ3KIdu
DKHl8QzB7Q/88TjOsXSNhlHecHmkr22IpvaMbHUtpTvIsIUrBq+usn3sGhIufVK29V8J2OKo6Jqu
znYOUUdk8VJ+XpjGr1PUex43G7w890yoriyOjR717UjsPrJBcPcm+uUg9TE7QXjDE2UZv2hC22+M
BTrh47YPiATNgUD2od8ktKLC7iL5zuaO3Nt6HunD+aSo3PdIwZ6kSMGo5b9e+stnWlfxHBvUV7cZ
MIsRP5L45bFyyazAa8eHJDAYDg+gLhN71THldjcPM93buIJH/HDnc822siwBulphdI3xiJWPIrXp
V/xEz8GpkeO39hqaenHfVwfYUAx0IudiIf43LzBzjHI3xqesGEAOk0Ba+pb7KV8XWS28mSkGNC3y
YWtsEr2EC2MyBOjqz2dvvrjfBqhlztiupDRxbzgFw6KpHk9eoD7C5xOLw/BJj7Iemy1r3O1otBl3
1gXfon4diQwOc00RxZBR12skJQznUIy0bgNUnqyW//fdn5L1BfE988p1lVY9dPWyVIKMubS47XdP
ixv8OWaxGLQPLDMz4jGL4qIUgVbGgXoVEr5qBlp7kBitFugcFE4rt3nP72iaOATvBNW5tmWLkmMe
bnl1RNL+wMSJXA4+/z9NlNlIPj0HmGSxYvwj8VOKf4sxzfz5DqaDOvepybRxmUwoPz2kU7AH94jq
3FjelChymGZVbIYRwxbSanRsBfgfVv5eqfk1LsWF3Gw1Kh/mYsJx9kuzyfn7y10vW98mPOwO/MCP
oCjUyOemYVA8BrZi7aLXoerMgb5DHnHe8xj7FpGEPdOx0vJV0chb5+YOwLUthMNrid/mcy1Ce/NN
qMNANwAeX4/G1ovnAe98ioXtNq8Ypol9TUHN72yAqyuv4DjPMC8nl26Qb77bffhF0miSVGDVnNBh
phc25YCO/4fmDV/U6D9EkhMLkNEKlPhFPDO4W0JZJdWQhXT9bQfMCPpriL3b7sRsVZ2eFIlz7wbC
EJh6LPjemvJvNVSfyV718QIoNin2OM93RN2DIrg8JumtWs/dt3ynlRF0vEkcpnPX9FYKApMFWr+y
1Kgmz5+09u8Sf90BqWTjv3uovgKCs1QGu5wje3FypXetAsuTOh/rpOkaTt+1mUmizJRIZXkUb8aH
4fpv7MLDnXP1MS8yMqNgNlAlqjIrLKeH+2x4Xjh08qIk9yv16/kiWyuKw+vUpNHSv2x3QMEtmTz9
UVBxHyZkH0Nvxxpkc5613SIGqK+5ZOXS/xJBwWotcANFQ1RlK/kUz5vqn6IPNqqRbTYqMJoKab+V
qHUcUauI3urmbBkJOki3BbLcuf2C4ZQzPmcArMeJTwxITxiRu7OWO8j/ji72CiWvLr4FEAAeZI0Z
rsUyOwN63i8RpbrHe2/VBCseGWVMNAMNsISQtJ3AlmsaxX4ucNLImQWZqbL7I4RLn9kOX06IBEmi
XqzLggLQZPGoL3AZdeYJo+KtjDtRE7Q9dOrB1iezJJYCdoBkvtbLk+3SSGziazim3kDc58BdQ8UC
pooO7E6umMV6CqVJQTGZZ9e+k2faM1yRFxR7Owsdbc1WXwJvvpPGf1fLUOT1RrEMQq36JFo3TTih
CVixBpaRY5d15tXuDLzldbim434uruvRoz9iCgh2IsEac8CDN8RnoX7w3aO0RsYrCgaqo8r72IBE
uRGcwxthvR941qCT5kcVrtKglrp4MqS1rOjkUOJeikDpNgJk5zONHfc32+5GQ8PqrVizEPGaAHKo
wbJv/e5JL4UFKZTTY7vE0pyReNmQl7wP4O8uPAQ/pR1TdSFKZUebnRMD8jyiVZpe/daijnRlbNg1
Qoldv4P53BQbYOLuW88dFAsSTZwmP2op3prWCkBnE/lylhF6z+hnI++Ma7p63Re3pllf9HrjIfnS
lDfbxtpi4d9qta+pPfnjKjrwYIV0igiTypsqwAXlzs5yoo5zOXuGboULWLRXzNKYRKsoGK9O7lXl
pQb/SpM7HOXTcu50Wtjd+DnlhiaHW+ftiAlm1djCZgviLkb5DEvzWVZhH8938cGSCJMldyHL1OkB
+DBDx/wHpnH36sbtXqt8cJCGmKzHFnjRAuQODjdy/K1ypD/Z41+V7DBSpZhm3EsnEfBiD35P4IV/
TAe9bqKVaNQhriN4BnFMpuQh3kzkcEfQWMvENjh/XY7XP5OM4jY/eji+Y7RfFA0VSGe6gxN8usnb
OfnYLo9Mrdatv6VMVFSlb+ScWovrzOkxCnAlQIdGSg2a0cZixSUHfM9+arfPoZIX0CngdZ6LbKVB
crT4C1rrHX14asb97k2k0H3slR0et1STOEPix8jPmkpkrFKVs3bzzeIiLHCVtWj0uZp8Ve/dhsKJ
ycob70JqE14oEFBlBDgBLa8monfcm/cSzsu6/sl+/1UCAqnjVMoTNJJyW/K3b1JYwt2E6wL9/vZ/
092sl3GDqPkpPX5aIhD5LoVkTMauQhSZf8vf7u4/1qVCczFnC/LS8Djb92Xs4V5awPe3oJ90KU5g
qR8yFYzzFAXPXHwq54ZLROo+9OVdlPtLkaTrMOLdAFtk83aKXlk2joWJggLSVj0lghywHFbMgseI
mONxm3hkS3uXaT72kwaPq0TypvRFPakXGxwB79BC1jdIVGloQ8QZaTy5WWEIMB4aWJHr2knyJNqY
+jSDQWgmodI1Qm8ZA/AS3hBrAEhszv1zUB4rxVD6zoMlsy5LTeftci9tSRxtL/FvnVqyjDSLOeJL
q0PhnxBphiB7OajgJieMUKSduIiQWbCzT5/hPS7qyRmFCPUDSnUD7loDevv1R/cyWeC1JbGIC42s
lPALTcmwUmKE8UBxzcZtHVB/aUdKAjLEDNrJ+Zwl1zm/X+AkQ22cVP2AYYTp3sADKi88MwXb3Ucg
Yws08/6+O9c2Jqzo4HYkBGgYJ5X2S7yS6EE3GPf+3Gafvd4llzzBQ2yPTTvX6KFX4bL6SBH7EQFp
xWewIXqTQ2Q8L5O1097GnfT/WyYxuFOeejlbaPpCg+EuNUbw0FiSvHcYYEBfA6tdX++nRhF8aT6V
e+nn1iRwhsxFsbnycO4cKMH7DYON56kY7EoktT3wsLs2sUQSLQPSIbgqBu9GIW0OHCKAlsjhgaUt
1jqI8f2UziyOXcxkKkJq9SCazt/gWFtcSdcIWSbXdVpwZVbGZ1Sjxrt0lpHb57cD77IDHXjT4LFW
1gsPNrK/kG8z1CsJ5yZjMA1JDQxxydG8SKQ+c2Zu+DwONiOKR/ytFxCENRrI05tpim0IOtoQR+sZ
WyqQgNh3Pk6En+TqyO8jMK9dEPH2vTgZ4NCw19OtxFqcuS3YFIo+FNAFRGt5CfONCo+r6/EWY+ZP
TQAZRF+P8OdH8SSUVQewfmYEnKV8pP/tand+XyNZAgB3aERJ5gbR7tNxRRBBQsI0fYWv8OoNfJjF
PhlFFBLzF+Yszr7zZ3ZHX0xHpmIxuVUVsJC54zhIeV4XnRueyW1qZPq5rmkNSram0wuvmY/SsuHS
zJVrTdcYuiCx1ugXNVJ8WcQJbTYpx2WiCFcpQYCcfdRc6mLlvkGvL7GzP/6FCJFm0iQAZFhTMFeZ
QHzMdd8e5N0gngriQviJQheJFCzMMmlMAvOuCc9BZMgEbKyCdpzGQu7eaOmmPR81odMKptnHaYQD
eFFfYaxsRA0feOzAs+erZLijzW0Xh+BzeiL2v2RiRqeOsmLM3NLLkfO7ceHhKRvSmUwmc4PYNd78
G2LAmmDivj6KXK3Lo0U4sG2N75iNOCrrsJOXDiyni/qD2KmPwbezKJyQBBUoLceYx6v/mq/N+onD
Jybf+htSZKtpOaPpF02of60jktdLVrmFX8mU4S7trhyYy+Q6OAzZH8Ikg8s2eyAUKPtTnxDtHfJD
Og7te41baotvLNkeJgukK1QQYrMqM75JvRH69mNQzHKx6wbWfrFyhfDhBDmTqCtfK65bg3llXu7t
nQ39fdCupZ0cs1wdLNBB60zKI+tzAVE0+gkcwTLmJvhohVIbqVkPYhg3k2UlEzf2fOvw3X/pcb3g
ATgBg2l01Oo/RhvpFFrYAQbdvZiVBB9faJseYoDdTKP0qb5wAxHxUURgpYKxYy5VISgkLr2FzFRN
lQzVUpW+TkwMCvKzWXI/SCbnM07G4L9RHt6ec1paJFnB/NmloSPCgJZMnF/N60bKrkAHvgeUqXs/
yit0ZxtXEXrfSek68vvhR0rtvWY1MsevI7pWkhbnCqIxgc6tKt7xeAZrueoYG72fvO1RunUwF56F
z6IDDyuGTPl60bEqXlnrQS4jtLHArgggU036WyOF0/M1+5xQkWepZWwYAXAG7erkrl3mDu1c9YLR
dOqk/sCcNxfEiNURfKPB8chqsYiwHSC0kiJIr5VmqYTlEWDaOpObfz7SnL9lMjkmJxCZqdtrRKkb
k0TpuuZvtIFKTiwmhbJEKAHspB02Yk+Tvikv4/oUQ9uEt1igNEFThr71pU33VUqeHrsWSQ3EBJuX
TFYKBP3eoaf+q5KzreXro9/4GMGTgVAwtPdi+dkWnyqyphqfbIp65dmec2sEdfKgUsh+ndjL/L0R
aa/3kFpEozYDFMqRNmfAsinc09CzXleMyDH8l2oVIuvT3JUkt0r2k8HxUiZG+t8be0Mqf7xOdunl
qOyxQXi3VmB8zqnVhJ0/ZTyN2zcoSQXokUwIf5e80P78RynrwkUjUonbdpY3i6Ldpw0VrmUnPxep
ZC5IX1dDNhcXkHX46qO3gu52qMt0yFsyD3P8G8Ckpgvj1C/BCY9OuZmJpvviCjQLvEwXAVltxfCg
PM8m5gWu0B8nZevunaSwa4OAp52Jg+cRfsU7NolLZJj02d4R0EqgPA3/0SNub2Rbxj67YMDpGsB3
eSFjHOpXhmOB9jOYksAEBvlhAvrEb8b1Bfbb2yeauYT8MaXPNnPqBgBihaivVAZ7eU4Jx7hqTvW6
WklN2LJEo7PZMu+LKJ+YCo5yY2J2YqKX3nBj4M5ybYyj6Q8lAvhiNxCkVygwILhcwHkUZa09JeSS
zLqzoEAsB8Z9LmpN77Ij1R0UkOrMuw87FFjX7pCTTxyVfkgKwZDWhVZKkeLvBk/TTBAXP+MtvCAu
r/QsoaZZa2lDkN3XE4dREjurP74tAIvfsj5RmM2dTZ5Q3hG2dX6ZRwU8dhkhkK1UYK0OP5djRLGH
QivWEUPPqW06qn6fHiNzt227cSa+ahKCaMdC17crQ2Hpp+ad+C2mQ+cC76MMi8W+mewaRGgVU0Ja
1+cfjR/Xjs69a19VFhXztBrMaBRcfZ7jGAcwkH+a9ggyLNozG58BZmhhZ+wFleNl2B9bgrG8Bk47
k7nbNGcD8/fzKpLqLHbfxO99Xk9xQV6qjX1g5K1vCN9eoj3AgoqFX7NzlME+KtTsCZGGiFmy803F
977DA8PoCXpAYYre7FV4uK1VcIS3pn2jDV+f5T81
`protect end_protected
