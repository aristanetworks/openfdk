--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
bLp5RswPe2/6LR7OFCrqTYXN//FaRqBd9Ah6cdZv555zV1avo+Uqozp/kJaE/xpWAXmPekP6Hkj7
SpZAqJEzbp3Pqt3vxK6aONBvId16Ggv4Q2vTWWxqIjm4pTHI6jrwWtwsts6EEPL4WK183x+Hmf/P
teYmqUs6PuDf2WSSMLVHyNb/YC4rAHX+nJgvOkWpSe0YwZadT1Zo+mcabwH3qR2LqMpn5v2dzQEf
jSZgjnW26vIm1woHfsGOoXAcMomHstJq33DWwXUFkAMOH/bfAybjNA59jbQiuFp1neirtf3hdJzy
IoYk5H7hWBpl+IWsrypv0EK2lWX9jaTC8JPD1Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="RuT5vljbGEkOOnmrs05wPIhxhcpkKK3xygFB2X8WsH8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
iuKcl51Bva77W5vAmm8Uq6ZvE0g2i5FNNWBVm/bLAnbfLJnTJGjTA1xEzj+Sj8cl3oQZelsbAJ/g
sKgLnes28+oFE7BfEjDKW9MqiXIieHOWa0qqxe/vFtP6ev8XrNvpEndjSuamybiGSCESyF0IoLcB
UB8k+SoLNc21hkFaLTx+2J+0wvQjqM7CklRfzQshHuM/1VCWnGMnhDEJZaiuUL8ldjGlzw2c7lQT
uNPKEX+aY/ymPM9ZsIhr9lQIg5n2Lp3Uhq5l92oNVp6MvFIqWcNrjxEi/Gh/uac7kNCAUDnJkWqA
Vo7fvFId+HnY/21a9O6ocsVYhwQNtUatBv9yaA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="OrSaPYTUKGnH3T9xQvx2knevM9+zvvFS7s0Rx5S7N+s="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4480)
`protect data_block
ssX5zJ32noRD3/Zo59yKUG7Q/2EJVIaZtkEZogEZdhBfaKkNRFc5ODnibgHe3MkAPQw9Bu5e7DpS
eUwCB9JRQBgZUb+qIgoHNcUfsx883nB0PpndLv+/TSF+qwZVuifE61co32ZSUlQAwLFzHmh8wLo0
XRNboBaD2TlMIBC9JPkbjEEAhFFj9/OKXaBYENzJU9FRKeEmVYLA5bi601b8nC8HADjxksnz4aP+
s0HFhI/r8uklQix0l7SOT1ur2laJkOWLh8LiKBWgSKFXfJBzXP4mxnW+Zz7g0/XhDnJT6LtuEJoD
nH1hiOp0fSVUgW1aeXaKXoXeqRceqtaNd3Npnobkj0p3o0pZS8zafiLmeSiN4z5gaoUioxWmpNLs
GOJAoceUg4bNZfcS3P1N8etmGUHZyi4DsxZzgAGXLiSy+zk96BGVxjhZJNb9HvdtJj4/+/jAwNL0
2CM5XsIpL51dzvI4ycuIqYOnfh9Z1GpF6hD43tqwN6X3P9RynDVe5abCQZNjo1XAsX72A24qUUmJ
nklFHMfbcXOz2nwGGeyk2r8LsfVFU7yEipPw7VJ/b1xDNTezXjO5s9fIowbOCicsVkm1dQFJCdmn
lp2cbNEZs6dSNOxzYMiFnYnui97QIJbffg6LOeMGgs8cnEMFdGdi5zk2zfHd6XCybA4hDDewc91d
PQ4Dog+J2ik0E09y3tuzn+RhRXLvzX9IT7Pzhi8u5JUfFBNzO59+xjA/h1E7T9oyXNECnpHTtEzL
TPyqo9jkwAHai32tdv+KPecPrtVT7Cu1k6uckUeF61QrMZPmSp8OcyzSnw2STOdsK2f9M5og3fIY
3HB4VHCeEdd7rOSCWPXrAtKRMRLKEaUPUmFXRQk3PX2OLA+OTxxlpBZI1+30NlpBV6C1DD5pSkCS
ToCjQvj4edrWr6weFuR6jKJFagckg04Ms5X5oMywtF1VMh3QpvgOWIQo7Prs8IP67UfiCXg04kiH
zdy8h3exiSn7xAClpFI7swuglEQNsGACtsTVLvmB000v2Ls/g18hEauXEFVFkHvbl6nkUyMWym0X
YD1G/b4YMvSBptovL6mTJ1scdZ00aec4kHx7z10dkUMrLlqdhPg3pjIOS/KA6nvA4YdSCovHN78B
lBgk/wwLux1LSk8gEYKAn4lslslfUhAGt+bddP8bPT98LwMilwPdNtVl+qAhG2Z+ELKqX9e6RCap
sym3BW5AJnJvdw4oL88W94Upw3ia9m5FMEKRJxeZkbJ43CPYwW2eIW8fONzLikXe73vyj/lp92au
2HnbULO+t1uPTNUfHhNa4SYSED8C/e3m0OHsuxAqTtCLZt7OnU5tghQCh3LopfsQFgZF+wlhT3lO
6+onzijJRdf1AR7G3j+njKoej2kHuQW+Tx8LUzDpav5dRo0hubu6I+p/Chdfbe8c9e1oDGrfSc3X
1XohA4GQwWci1kFUtzEO9HvBPS5NWXj8Esi4e8sL22phbHvYerbSWdWOgrM/RqCy4CRJ2ddrNm3o
T9jat6nJAdit8b475bO2QlCHrkeEdGaj8TYfNI2v5oXoVYrhbKFjiYQpEg4V3ANfDLkfr13Eic9R
5y17cVRzv4xzU09hmZ3Yjvk7F4eLgMcqKNpyNp6Ff73dK7/UFOtRmwhKiu3YkKj1zRHD0IxH68zB
C9XCGwFrCONcY9VTew88mS0JnIVezP9jVjeGPwystjRZoNZ5VF3kXBpOKXMV3EuCIcAyRXFaNzgh
/2BsROXIsaaQAvKyis0+GtJND3ABqCE+ZrYC2x7cCZYZxzVI76KT7oFJrGkYNyLHdMQX3BX9FpbZ
SZA0qWjOTHylYuXtn+WCK3J3J/Uy9hqKkqHfFX/MaKtHb+2SIdI9HW5UEmQ8edeEmLKiox5v/rXb
DlotQElrvCqdASqYMna4dtGeMsRUzbS8i/1SegnfvBRMU3LMFb2iYrNDSc/yEnYfy/vQzzJ/f7Wq
ayTwPZcd+hBP3c572WbqWeT/EWFQ6UawBkHy0jl0Nn9l1ZUKELsW708CvWzpEDG8k10HbgN/1vQK
nKO+0/pkWBKT3VOsNp+1hnqOBusVPhjGnU5GV1BvtWHc7HJDqgBti1iUI8kLFGaK/+S7QXN4GyGg
XOhe8o6dE+4VBbf3/AoroEyJhRxZPyVMiEguacht6FDmSv6X21hFTdOCV4UwoZbU3FDqQZly0FlD
80z2U/96a1DOrlgcYgrAZElhivRK1R4+OOVlWXEf9xTS4/hJj3NqkAwXb5XAKY0sIcz8r/ur8HJR
L6qyiWYTgQI3xtSwObbr/pd0RmB/PNNg7V9QmUXDtOSd+ztyNbne3rBZ1zRdv3c8WQC6nXnh0TY7
+Ei2pbZrdIQN5juT7OgWiK6ClDfyIRcD9B/U518OWPYOQpA8TsszoZP7/RlFGp8A7jwAv0ok1+vu
asvJf6u4gjly/q0TNPcrh3m5aiHdvOTiHTwcjOoqf2DBYzacAtcz1KgaZfPDK1hIGD9aogTPBW8N
qwUdjeG/7RmQi5FU7bPay0/KiRfQ4K9i41WjJGh/2wCVAd/BcmLwgiM6n3tPYRCXDJef/BVJHp3c
2SFlePR1uIv0mfd1g2PP4j13O4abSoGFhDKd1VKBvd1d8cgDpGiuJ0b6qjQmF/DHf9RvvckJg9LF
tA6hrq3CbG+tjDlofhbOQdMPRlfh/+8cfnQRMKnKGFBmDosX5qduQR7KsqpBhOPidbstdmIrrxFj
C4zZW/8tdjbXDh11yCrVBU/ho+XV5BMv1Nit91KHJzFRMqS/L2LTPm7JFmRBm9abowJ2BD7VbPSx
RbZRujyrO+wbwEdfvjiBGWaMU7eu+0G1bsfSUOHgSAT+cCiRseEsUGT4zAETTMwhu97IQoOIuknR
Bc2NnTG9qcCQGq2HK5zXf8n+Ok0CMS67p6AAUe5p6JoiQlKp+qXORHURsCtxxNiAJEkKOTgMi3pZ
iRFUhaT8WrPNsEEtY7BERwSymTJAR+bhKTsG/NR2L9UJNxVEV9aZutgT+RQUXTuNLpF98lJjP3Dy
q6ExRnm3x2D5hB14wOpZjhsjvqYsRWMzRSKvzKCUBa6OyvLeKHhzHomebxsaCdHyKrhg/dT/kx9s
kGTmIrr4ZlES9nnB7RzRyhYdGwHLZZcXE/1Uil0qM7vLn3okhzL9r9LY8saGt5BLmrCBvFe08dAt
+Con+PtiBqiRKUe4qJ3UiwcS1mwXxvJj7vQ7j85dcP6JogeA/1MPVuMzhys9oCpj+bkN+oX9C6dp
+gVemGHsgs/e4CHTdkvT4B7bfVAh+0fK7U6guYsZyU6hmHarm87vnuNcULvTvdOU97jXNnYXyjnS
rFkTCq4KbDuvMG10hANIfbTe6viApqJ6l1yVEV4gq9fwGoX34n7zS+nGEcl6G3dxpXNWkicFfDnJ
H0qiwwTp+roBD/HrFdzqkHtyZvIOMuNuQLLJexr6TrwlZjg3BLpDxvnIUsEp+oAvXikgtL23Pl0Z
8M5a8w29k9vTzvJlAvxkKAAUXUhHtzHpLPzWaK+taIn5+LxdENTuqwYKsDtQsjUUgaC398fAOF69
6ZbolHOon8+/71D+1CTRR5i1kBbz2sisuVyHwlkhRYHd3+gi9r1JWFX7F42zeDvPrX4RGgOJJx72
eoq6fCy1P6/HtY7pgHrHbnIhFvoS4Og/rCSTOKieEO7uqkkgRZiZ+TVYmNVyOMx6F8U9nuqsZlOQ
/9aPpjuXwfW60rrHJhcHqOWp5ZU+IIsIpbX/5Vhpc+4bMIiXaCLfdS/N1CirtO9mkNeeh3tj8qvW
FAuPyjsK5KsobCWDqpm2xdnScBBXNnTB+cJWGrQrivgAvxhq4rJ8DG6v3gQSgQSrGDkcoLZ/ikvu
fxk6QG6M0tGE/Ua6ZEOzA2cZY4SCzaSaeuE/Y8pBo4quWHTL9MKu0BTXkwCkUCjl4VH+e28CreAK
njCJfBtvTBRR3u6LvdMUmMoImQkK/dzlLFSrDwgGv+PWz3kBjZXmf44bOi+XWHQrYlQvP0F+028Q
aInXOkByzCt6VQtyZ/k8FNhQzLLlEwaC9i+lN8IFoKCMTinHLo3Hmj3R3QszlAxnwC5kRh/DniE7
AiNpB7rVPvsU0ZbFz6dmITxm83ieg8lxbJ9K74xuF/X68GBZwLg5B0YpNDaRQJhIajQRSrI6GxvP
VrxE30o6th8UpLp27bIt5URM9TPCfxtHDkolwXebGkEEwOyPgWKWgYgLXZPHD6eGNDuNbW2i4pC1
P7BA3CDszgDlRaWF+oKUP9RDfK0HQ59X/HnSK+C+DxObL+24dBQbP4VaaW31c9pkDU3A8V3tVNv/
apvjm40vKrxEl48lwK23WLxn4oVLkPk3yXq88+SuS/S+aa4UmXxEknxooB2qfGgvJ8H2VCRpYkUc
iIwTf+gm4klnqJEiKSydQuD19SvUvbSYTuHvPW2r/K1RHA1CKVVhjWHTPZ/C0ivBI5PHcLePsyoG
rlndR9vrW7+bCj7Qzbo7nR6lyfll6THV4wl0yzWi3UHeBdDWxwwOW13uNYMfrfQan4aVtILMZ60B
e8g+nee/bio0dyQIJPWMTG1XQ2lIF+FSCxwdyAJOEJehJe1ReRs+nC3UqHWfahW+HIxDeWOfQ2jb
hp1AyggUC98y5EqhXhkjknmOkQO0Oq0WLCiUc4QbCuHAQtBTltBgkeL83kxiv0iWSRYSKGzFQu4i
kW9KB2IZynfqdd7Ger5RKfjJARAgC5JJPNw+ni47CLCK4YAqsjDGOZSagjRaYweHwLqaYmYUqvru
yGgILV9BvsUzFl9mcCbElDb4hIOBwEYSdXDt8D/43aOrBuy6E2+qF3AfbmZuPVPxxTrB8JWp+Y+D
jtwOJrqz64MlFbRdE8lSzoBVTuN/Oz0S2KAOsoPwoGNpmN5zQlfUN3rFGVmiHbgpmmDPUUJbQxoW
or4lfGwSsisLMxJVreHGcupdxvHr0YUQm8/UKTeECxZYSo93WJSObRLgy5G2GiWm5T5hnZGjrowD
BcArmMSsOz1G87u8/Swt7RXHh3vdEnMfLhleGnm2bqzHr0j/UKHCTSSELp1bbMa2WnUA1eHpZKMx
VjSRyw/DsgqYW0FhjAoz/1PRsmNA9Jv6VclXgnswUrEIa7TmPevkMWBGDdRH83ppukaRJLbaZ/SI
5/UbF67FEDRZQWRl3LAB9BoZF9yhEaNO1TxdkTJXcqXHaA3qfGpAWXjAEMz5WbF/USouqfuMg+xh
BSilfak3LU6gMf2xcdGUxDnIt3vCju8q0AabWgY1YaaxCfFtClNCh6uuUhdCiiXCzOOOlBC7jhdF
nomUX07uoDXqBaAM5464usCBhEq5e3oMwaBKp9ldqgMYNmyocSInTqVn4HSp+YDCv4zB3FgVUtVM
4IruE+FmNwZ3T0mFT1xUtsfrYQgky5tfem+RAJgZ1bUBJ2kuXNsAMwKlSZ8LoS5kjvvSWJWaRzjo
ZpqDEPNU9NkCEpRSK/M/yIaHfF3I2nKw9QB6Iqv33mLlAIbCYhUfGtTr6XlzUHPueZ/v4D12/TyL
tMHrufQdD57dinmTIy+RGUmcMq50WA/TQPYNQwtBBXw19ltC9drNNxI6dBtkdAQJP9/noZgBGJRs
LQudZdCK9eeuUpDkFEhq5Mc6QmkP4C1CYW+quKmJsN0d8IQkFHTv3BDtQEGZKlOKJG0oeTg22whi
3/4LZKtksUQZuPYQjWcxa999wUKXlRroLtQfpD2kxjSQoORhobf0vJ0fwN/bGhAqL+Sagt0iZe1a
fUK9boO2rC/LMpMAcZD0uVDLIXnuGN7s9RRvCIbMI+lJrLNgulVt5URLHRJwmi5IyFaQiWg8o51Q
8Ax8rln/6tkfunRGTllB8pLDlimEcNgxv0B6YorkXkB2XU7NwoanXEcQNlZjD1WhfRkQe2h82OCB
woZMtF4G0WBFNx05p3xcq50XYEEIhwNZ6OUW3WwZz1FivQ==
`protect end_protected
