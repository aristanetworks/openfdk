--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
djjDvQrwho313Ct6UVeAkfLpUA9hls0rL0plq3WfJruQNJ1Q7/ir5kLLZWP/TiplRGPAAhNbk8QB
6Qq2a6MgeV9VNYBpi+kC7ctNAhbQN20VAwvAjYjR6KwvByfnuqaTL+5UWkVKnHF+DH+5ORn44Jj6
RRYzHD48b/9a5qi0GMGd2fBqn/HeXO92DM32kmScXZUHcCe2ZwS6ot2IiYWkojDl5HCNkXPwk6gU
iMXg9yoXPuXT/iUqxu0LtviHp9DgyWZZWerU84dm6DP/daNz5M3I7rx+lVLH5r53IdXdf6Vd82xV
cPZ7ykvYB/EL8DBjT5upTM6CdAru+MEhV/cBNw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="1kwQ7bg54WNRfsoElggQLoknEfJDE3bD90gG+1zrFas="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
BNrbD5/ei10otM3SwTcRB4++wgqHzU+NcCCnvLU8010fWj87i9OUu+Y425D11A5jrrFPst/VDmCL
RYb+E2CXkbxsdxP0xkBLgdF+U6jMf7bFU0lC+WZZjGkYbZCICGON/QgiX5G0SnB41FLxfBk64Ppt
7gijX+bp9v3QMCSWk4tyR0V2XOHYBPNINteclGb0tHy34WfCDuL6c71/beqzfzd/O7rBTDSWBH8Q
RuCZA0V2eSaq0B6rHH6oz/fydHvauzrva5H2gss3sGJlAadrUxT4WhelFcWyPgdh5MigzpSUkJLh
UXSBNEz0vb/nZDVUe0BUHjHshAPbihz8jiKjkQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="UI4ZvahSF6vzxdOGZ2NFSFccq4MEwNRBFdgAGLDI7R8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7632)
`protect data_block
nfaGfEP55FIRTMmmN4CAFDIaMMfMuT9KILwwJS8TTWlvaFbiHhHvVJcF/udkA6x7hcAA0XoX1QV2
enuIRgi43LsT593+jnftsImf0GfYSIwJnfY0+mJUaDStQDv2VDRsuFxJu6PAmiEYODAbVwxYwC4N
SMzotMUcnZx1fMe48G0dmsbtnU6oRRlGJCFXcaCsjS0QDeI+yDfhtlkxXBQwp56c4l+WBOgQBHbd
5USXbdV4gZhloY++Lg8aTSlowHT2ZW+kZKYPsOtvCcZPvVtNHEHT1G2MMG9wobSqAf2klN3881hc
bYu0dZn4xCGelmFSgpDH3yRB598BgE21WatmGYVvt/57dlOT59s4F61wyTNNTTVkMGH2xOvOZhs3
sdbcbwdaHdne2OmzaIfUsEpo5JF6nGhy2C4k/Cs8xD7qm5iaAkqIxfWNYJnKJpdBwLmNp/KnH8q9
qWJFzACY8jXEYHvtcHxPG0szaOPQ+gSwC9PwKD+/36HmKI0geboOjR06l3jTF0qw+0sqmD72Yf94
Hss6mVn786ITjKUwFFp6feGcgWOUxilxi9gijREDvBXiPdNHkF/rFC4msMky4+cHhsag1gYr+VF6
CgbVy49GG4YkEahHSET3zlwkVhwAZUCechq/KPEfYhsqvnxl8bcAgCariRnxzqtvr6Xz24tq7y+8
vm4KAUEwRdgg0HCru0ceaPAYRw/a+QvwlqAQw/sGgFEVWOLbSAv1Xmsr/W7UUGyt2DR1k9FNmQX2
E1guTixjR9sD8F1bt0D6pv9qdFcuDAq9xz2ZcGKgPhUd40lqRtDG/+eyTDgzPQOeMWp/PVqb3DTK
c5J0cbeMmkKHp5VIX/SjLM1J9btdeU0isE4g9Qa0SeJJnCYs4McgT8+QyQCSpcYHC36/xyqqAkYb
0lPbAbJMl8bA7meSayrjehRQdWh70SZ6AEK5HZUPYrHHhQcg3Nhg6KPKNfTWWGRiqvaaA/hMo/F5
5f3amNkGPAhkqWbHubt4lH6TYlnvXjrXiH6J6MeIovzewkxEWP6rr4n08TbIaienG6eabs6wCRWR
Ah0LMKcMB8jFWZpasFlHkgZ1V+z5c57a4fR+sA8d1v4Z6HFwt6aQCQ+ZYSF5vshqjR5QydvEB00H
01Y71b/nunsCOGnidcELnngC1DMO39wWiIH/oFfIjx/N0BfSUGvbrkDkQPGoTELu4ocsxFvW7yvE
41WI1icyJIjTask44zCOWT0spN3mH6MYQASfcmKvcPEtoYGFg3CWVhZy9M6yoJzErTpodu+oFrmW
PRTgqAiQqsvELWBWBYWXQTDQ0eoINYM4xIkTvgQTaIBnhHOGEmhre+1TGMmobeNjhOBiaKdCNc8P
fp1H9sYNxo1UI8shnikgVs0VME7Gv7s8+gUU4qryTkdcMpOTS5BZe9r8AWj45epnh5ZoT9woh5p8
66puOXuzmbAoB39MipyH+qyNF+4T1UX1+T78AdpzLyJaDKL3LpVHTKE30wrbShVfjenyC6QF9XuI
79WeI4jt0fML3QGrcyRcZ+kIwzLm4l2daO6aFBDIDOPzHuyuSSI69/kYwZeBEZRVY/SbnAk8nh3C
a7bVcx5uAVi6/qMyhuYS2R7ghCW82MRZ9YS3V1iLnyZq17J4GQWEJr7r42Kf53zepPqv6O7pw6Rp
UXn6ImlxjAIyFK3uQRHBJBUuQs4VxWcebj9wrPXKAeXzByKuqG4W+8yrvHNUYD0q4Rv3rH+8S2Ho
TAQLShW02CtPFFR54MI1RcVJXFf2DGBjnGTcTZwLryMcrIkjfDmKULQ/X0albJEObxdhkKMMrp6K
4kDZyJr6U1ohdTCsdg+lp0jDC+q2SMpyx28Y4mgjhUAgeqEC6FaH6U/PZAsaud2pwLyyTPRaDFqS
SPm7gsds3PTTUE3l+IWw/KUoJGgGCAfkBtikqnseZ4zhs3kP67Ip8ZWSYkKm2RM779wRu4quQ297
TKGoK1gChqghnAqM0YByDKKRvk/Az2SsYnOaqKoJ3+Wu3cdaVBtq8sktWkjjuusYIkPdb4GfO+rI
eKEVoDGwU45m5BuYCml0cLP8I9UU7+XnmxGzuVbv2tXaKRK/1E0QA1F4sS46xYDyz6/tPjdpraDs
1ZcRktrX4/4kgl/r/zlgrf7O3OlrQQPQ/oMlAXn5iu6Ez2Iw1bgoiqPKBktJq1qHnSS5pYhMw7bf
we+wlA7DF+9U1nyQlX/jnOjvz7kQe/H30BygulLxEzfsaV5fO5s56sgh7rFAt4EnIcSzmdK3fost
a22AvAQxlNSL8n9KI7l9FxDpkQvHIjNICGWSppOgID3vjYQoYKPmTd6NPlkt4UCcYBOimnE9Rkk0
GC51e0Cqvp2Vvuklx1WAtxoflD888svz4eo9Yv41YWLG98BPWUBYidk0ab0wjw7EMFSDG//oUtwz
LJYDy8MztJ6eLL7zQqKcHO9HNf4GHnjoy0tF1lUXJTYFmgMFGUVv+K4kZN+FPQdTCmTMJ2dN5anD
6MCMHM/VkFScWZIkffAZn+/pPW01kUXS93weVHm/OOP91n38FsxA4cz+0sljyoBQCebtKAp/p1ft
QyOxiiooBEwQtMFQ2VugaEK/pR8/5CJbrBaoF+B95AoXmNFRQcyZtXzneESmmuL/hqOaPVych4gz
i9RPjYnJvw0GqwHMm/6FWO4f82dQk66sOvOug72d0Rxo5IEfRhmKtqcw64c/gBbHcQHQmOOeTtTn
oCIATkk2ahJ6v299Ig2+NL8dnPTzYBBYvxJsWCCCftANBmhogayUCDFsH0eMZRDIk6Bg/NqMv3kG
fsomzo2X65inMdlQg2b5ZN7jx2nyI8k/ngPZc3tDxRQdPFP53wlW0G1m5GrRtpPT7Jyc8wae/6F7
g5vgEVql+ZhkYzvLDAyk5L08rJoBh1jaCTiCbteCCk+Fn/TgtPeYjW6yiddOXHaxX7NQF7yNYnUe
M1NBtIbvpG4RxkLpC29v/w2y235JmeIiRAM1jlcXtckSBc9Z/hhJf95ThdXHWMaA0fv7HufPMuDD
FW+M8crQoVY/fh4219f8edxZRZAw2cm7KB26zgj1VUq1sf5f+XJZC6ZD2h0lhfwqHOFFd61nM7Kp
hM/icJgDMOi2aWem3wjM/YgnvD9QPxFLiLoEfT5mWOZ6jjtMJlc/+bTGFmxTGSCS17gAO5uaXIjv
EQTElpHtlUlqBvszxF2wnGZ3dC+hicJ9wt1xWP7MHbW8ifYTrsVyQS2hiRzEZWL7ui9mI6Qs/oif
oUk/kaV9fzWOlpi1wqTIRDzwB7yQq+vFoEQ5JIUSmeo4OmN2cAwWBOqKLt/G65MdxLeYt9eCsB56
agRj9qc1S6YWTbEiNpqu+GILJW21GOxgtInGt2WjyV40iw4xaNx7upqOeISnc0ui/PakAHBToPn+
Hz6ZIngm4F98ynpbMk/51aqRX7XF/tiFy+R42YUNLklYRQAYlDJIvi+vt2sdoHZpoBcDVmFD7R3R
Y8iMmjmr0HpF3JYUP4oyoeg8AwvmvwMbIdeAQeyAyuo0pBgkzHaDKzCnZ3n7N/kQYmrPBU9IZKHS
fExidCQvHvRQ1jjsws1PwupVbh8Fnv479179KfFnf4c9sEz5iFsf6CvvKWqoMmGftWECBUIbDzaL
5C0+8Rr5AZptWRN4d/jGqzU+6aqNEtPGgEfy0PXNmxQprHMYDBCiMbzgmzA1P+Xtyp3Vetbd95OF
P3OmPQZvq8T3/Fbbdsuk3ciQsqxGIv8+2jReMMKAnJryd1qIq5WrB9cI0xKrfPIdnbWeu9Qmt7cY
o5t41zFi37sgCGXTcfdDAzqXRcKfiyCGswbtfQ9Z7XqTrJqIbiOcJpUUiJFdZWgjyLqAKwwjWZHF
/dPpqt1qAYocypr+RHOVSlk2vlppUzlwJ1Cj1AdZoPWyWCqHmbZHdMJaomX0tWr4ami7gWVXlgUx
h/kOcNBLzttcfm5CVK1Fl8V2RD2hBS4NKnLn7zKWzdb3yLpH+N0VrrI3/+DieVvhRBxZsNsO2CD2
Trp9fqzIRV2kcYekhWRvuM1gU73cD+GYeWQsTNprQmyXRsM3NPx87K9YO4jZz9DHjTjRAxPk45EQ
ET1zuHjyyCG4nc9SWH6j5lpYDjcY0N3CYafKnQO5/NsKQqPrLVccXjdmV0q3PNAMxx5gYtX2CdBU
UvwZ1C8yXux7oMKhElFt6LIL5Io+mnYOZLaInl29s0DA0D+TE39JvAnJXAih8ZXe6AqupTgNB6A2
d/IwnJpIxJPAHNmDa/1fADGRslFWbdMJxGqGAw+G6SXVi8ZJkzqOKdG8jgN4yMCAFkiTScm9Rwp1
ATIz+aNI9+apZ1oaXtLuLv93WSZVgKm83EZCfIKXaeg5NJISwFj3z/jfqGtRcfXs91uinV3XLM0Z
dxz2qPoLdQUSbT5CkUwFlAlGH7I0P6iDPsuUGq6k4puSIIIWwJmeEkpBRM2IyV6okitJ3H70a0fV
Qm/3s7b/Cg97tFwmRVFhRyJenr+h07sRDipfGvcTcMfzg6AC5P307EQSSWcMy1Ns1nlB+xG8QMO2
6+SxlO8QA9A2umbdvoWUUBYzgRIPuexG807SJ4eVtlBrjUvuIjMloDB+EEK5ZXh/o2fU0JyGjRjn
+qU1WDTuTCCYPnbedKOhsdEWhVc4A8dyJPQrBCI8N9Rvdirw36pJzG6A1nOieXI7c7renSyKrsPU
6K/Wexft3TwjV7ODVJn2GYA4TEMBhM6I3pF2KgPrSP4sg2WxqugZj7ecslciBt/ePcnCAyKjbZO7
sIUMh5P2JjEu5P330eoLz0mFsKzMuFDGqQcjb22WSMSD9V5oDAkegrCkqbHv3qPIhpiqmht9Z9BN
eWyjhh25uZnZvnzWWjUmA10DP8voe/dJ6L7cbSiGYECFO93cRA0Rj0YW/2kTox/xlXp4bWscmX8Y
rIpPqFmIvIKeBDMf0c6wemG/IYcbb+0dl23wLf8RUolhilTsu84BTmzi4e1LlRav7auIqzi0gjoO
/KAjJ/qXcJeAU+kgWMgfqifgjZw3k0Y2jPqSnGmwIwUwe44E3PfSddpFgmdoP8RQJ140onzIDLHM
CMBPw5DLhKju+xaVEQf/ixTSlVEO99XGf3zwe+Gahp5TkVgH/oMnomO8Hk/1uTKWoOTg/mY9EXdM
i3Jv0P+c2o5xDnKjuKt2GktsiYGYoOGz+9+4pi/j7st2bOL86UOkiinnWUGi6QG/f5xuH/6umea5
tQnPYK8nupgM2FUutNqFHhuzyg3SQ/Lqb4i24xffJ4HLSNHlmDcGGwwDIgZJS7KuJI9gu9BwBnW7
wobjA6WvqmebkmG838P8hJ1Q1wGt4g2foriAYONK/THR2nC9SBn611vH0cdDbLXD4RbGFVvOA1PO
YZoMCzu60vl3URyB5Uc9FbNpzJfXjoeKa7Ah186Rlfb4axEUxfcc+gkrCUfuAkS8nmPK0z7Cwwbg
T4s7TMOhJlECvPaaH/1AA/5EI0RmCLolttkHEmB/wc7YX9GRnLV/YiE4M01lJhRX7yBmdYB7VLLr
64oK1CvHTVcB13RoFFIdAFV32cCn0clbPzClwLDNNKLcylSpeMr6WFZmKdFtcaONTCS1LOcyTJi9
Z2aA/TLj70LPHbdm3TevEqoqlta2zOwnn7iJapGwJcYkiu8jrcPoQJh2cWfAplUhXpt3sdOrIC8z
pL/zCVaEF7kYYXgbVcFhkBCf30i9GrbhPkAhMveNgpU2bYlNzP265vlA6sy+bCtRBEkCBJsB4zzK
qgnAAY/u8qwZ3ctmZzUcpmGdjYtE2cCfhR15+cLjFGWPRkNEEgcPUFCmum88uBjx8kJl3mIsPu2v
2YYkSzyNpUcOGPhhZejMcwDpgBbPcKncp3UmmyEvUnaSLYMrKgqcSUfl8H85rdh27SctT2GQ279B
5PssdXb0U72YEY8BNKlc/ADGk52D7aVdBfws2wIa0ttTz00A0Mqwa1TiG3h5Qu3jg65ks6y7QsOi
7iGDtRQMwsWtW2ttgU7Wlj/LTFvOyxxXW3aWUbRELAOEAh5BqzPPIDSmYotbuE9wvxorfnflc4eJ
K7AL+CgyyFnmUKgB3bl4wdr7/3auguYLjLVp6pIyGmAGZJHRrZ1mo7i0hosqKxVLRpNnXbU/b54r
upiCYBfYpxS7EwrFHQLvxgxY9pGcmQxsuMbdXQNuRPORbj5PKFuuZNHCaZDdm/ANRoAKSTC8q/uj
iAG6QbkOID0dSPK3UYZw+7ZH4BYCDeLpsWR07v20t6zRdz2/rZ4kc50irNbWsZC4+OY+/K5AnU+c
XbrieSpbG4tSHbmM8C9fgIB0Cd+k6PLujo4o5/CafUZgonjh5u0cm3U3ndisRO9rm/DJQynQutZu
aR13WUn0Zh+9AXNhaE0tjPdW7HbpEnInalq6xhdy+FGC2H1Ovu04nqXb0cAM99/acqns6GsTi9g8
spYmnpz+mf2USQOGhx3haVldCVZb56K55lYMafM4eXVVfggm0neMgEgsoa5pjRMDp7mHbiYHeWHg
g8lorzVbOUMd+IuI9PHO9/oQkQ43gkfocm4NISYI84vVJvyP/u49gdEFIzG2fU7Y+AR6c5Eogr4H
QBtkpawxCj/u4h3oFZg3lbHwbA2Kg44zMPSynLgm5IVtlSiHUtWoCdO4fvlqmG8NHktcQjx+gdMu
L0eR83BQevl9gIsoO7w6GwyH1WKOLr+FuRSlX015CbQo5DKLjZ55CbNEA3LV+ScgOJiveyszbHu6
ht/OWHm1NdGc3pyZyfJnHW2BsgUR2Uvm5tUaerHNaxsoeSZ4TO22tcUmjCTEkJ4iaFxQMm5+HaqO
xNkr62t4AhqiozAtsEkB+L7vTZST8B0sVBb9zGWopgAgBsQ0cquy2oWY64iY1FU+ypkr+BvOev2g
AO+3CiEuE/lV9qIBSB78//jNt9vfir8EWd84sGDBQ4cNN5pKvH+3EPXuBzsS+9T/A4L6snrGsFrH
kW5gBZIngiZOb33gx3khUk6EfYZS07kXUanzeb1reo3+LdGd+oDyc4NXmYaVnso1lhZGE8/Yd9kI
ihWrOg7yZLNX10BkhgZrMzfLQsF4E8aJikicDNgMfrsXFoQJYhEabZn6FX26hCASmCFn6F0mzWBN
Ate54HUftCo8QxHfrwKblA7thP9Nz+ObQmiMTYH3swI0JRCCSMEeb0dz9g0VIn5dvCG7MmDSfTnf
q+FSrB/DWJNcRXXwJGTBKIGFGZuFX9cOP2Kmqv4ehFSXNXUlY7woVteMHYWdcIfETPs/aKS7C1P6
GySjqDtArrWmy+qfg4+bqLdRELs7OPwrW2lhJsm9ta039MKiG6tk/F5VOVh2UYQtW9yeNRERWU1b
U83ldO1P51kgoC0aIB/are44u/nd2HrsvvlF5HKZ6KhNSpzdSWFEu/Xcgu8UZHGPRqLNvi+6ZrPe
tIjlXw9NE4ZKabuFGMxmw4SPG4sw/uaQQZWzK8DUl3evj+1K/5TTwjGHzRVvrn+L8IW1PLdnjdPN
Tktr/02eZjjCK9pTNTxcYbawT+X3eqFcroYHCxXQcYoVdjnxLecJw3CGMx4622iwSX4uXzy8qpuX
sdmTzrs2bAvJcJRUz9qMC6rZZIoRxK8B28shvgTXlXDNsgKUk+JOErl+kmhmg4Jau2JSmcKPshl/
1tbpJbuUHsMZMVgsN6OZI73CtM+FkfMfxSUxtnYzI+ZV+6YN/CONivQviuaQDeN7db+SncK0AWQr
96+8AK5Cf6ouGORStUyxU/auD22uBdFDzaB2H7VXMFdhWPHrZyo+r3AikkAidmY3z4dABpVx37Gc
ZyE4M+JZQ/0mKLRQJTad6lgpgQiAbyo1wcTUcjli+6yc3FZDCTIBkLW5ku+/VZlZRFNBIhO6L7wo
3tNmPyueSuHReKL3hMUwWuDYCUJ4pJXMIDvlg8hlIJZsVZKW/MQkBHbp1TvpUoq1dYXZuD6G2t07
NvwS16S0apaXnk+PAC6b55Xjy0rED+2M1XRyTVIZ61LkvyKvhYEcSgkD2UPCq9Od3iTsEUsC8tXi
3GkHLLSMz0aqPgtC0yrwAmVkDa/6gmVF4qCjetenz5cOGcHVqZLe9dW0ifIoPR89GRSzoLyxNV62
EduCE37MFEGcrAeH3IcGEo9aFpqpJFbGTZUewW6rnvwzhhBKfe0Wr86wSxeTpyYjEAlxCz4Bxvl3
QxhWfW3E8ABkfg0p+3ZXKodbVndnZ7Y7/NpZHJk6LWzCN+E5nrv9eCNtfcEmjMe2R//n0CmMe+ro
APprCKpQoCIrElEw34XUm0+Ig31w6sAP1WoNz4zv/g5So3oXfwyMdyzmyoYuAGvPgV99Nn6JV9t3
hX9QYnHm0cq9nNzeuXXv2Q+bGiFyoad/8hqZmIOHp/1CW/plBxNgIMJBAne7BJYu2IPDkVtK5+Ug
ZQ/dzx0+6wQlWdNgqtAoAUnHvZPw7el1aGPpW02+2cGSHPi+D2pG9SKP0gS1uIfObd1ux0wnuNdS
6LfXSMGRno+xyhLFHQrnCfxOVVeMyeBy0iejY0LKRLMDjIGwejgClROnSjIxvKvTCuvk1f0Tnmde
h3aMo00s46hWKW4qH2rvpJQ9KOfCJmD1FNq02+F/VtN0LsAiC7p2VG33DQ3H5PSm5+b9/kCtPYKV
9vYNNSyZNZL8hiR4RJlxATzRvoOREP8nibbvgEqCLPjgdlF2J1/pwPq9mGvHEUlglRJnYKSJKi6i
oTulDGu8QCoefHsKpW70TJczLOwv0cx3PLYct9oD8GaCWjSGSUzYr71Agti9zjXQyEKA2rnelyVF
wkhZwVFWGzbL6p1rs3I4FDaDepMHzrI1co26UoduuH3OYCeaJmOlIcarmM4VyLLtALHdfjOmYcBQ
/JXBpxUs75ymN0UqabogWPoJksvJQErvgLYmHRDij4TV/U5Q/758iO+vGzxYtqsQMSQh/ElFtqUs
w+AWSJ0kA9PjAl755/3JfFoTqZ8xETI15WoWEFEYeWHLnTQybsgJuPdEDprDWuPh+xzGlOpbQzB6
EyYQn3yqhGLJ9iLzol6y9SlDJvJY80bAwZeKE+ZkYxwcM6HjIlemCWUf9mZKnm72pduAzxjB2iOT
XCWtzR5g1P8RZAslKvy4OE2C2p7MuAhn07xFIedlHBKzaAaYg6a3YTfCGqxsIWHGU4XAr1LYyQ38
gxFX2sDaDIM8bYgQ4mfpZ4G4vgGVqja0L1GN7mr6We3mRb3/YARtSfaJP3lgi6NRkezAncsapUQZ
mtyBt4K4S8Mbl2nsjRww2Wyx5leGVpYNoGLvTW27nb0Rwc+c1GGwP5DACGH/6LKLKxOc7+Jo2wx5
C+K9ceFqsgDQOTAdC0uIjVEtJll0AURyE4KwpdSHsxy7LSWvYGrKGRF5oLWGJHtKJJT+qAhQGk1y
wPKzMA+QuTdXhnx26eOoTR4aJa999kSvubdFj3qT/U6FS2o+cAwPlXHCZ2HHUM9VKPx3JBXxXfQH
L8NDtnScdDxWj0P9dLh1bXhswyxirQq6AkvV1GrQXPHFY642Z6ebP7nZFbTScveQHjs1WBbEoWVc
BlslM1jL58mAI37FWbSJde74U0LARGU5KlyoiRqqp2GFU1QHKx7c2F2Pzc8QVtSixHDzoO7lBYo9
5ciixnSsVT2Rreg5pAs32dYNjilvxPQi0mGSnZAdT7sqGaPxeVh8bizKq9dYtkRiTI3rFn/w6Atg
UYKrInI/KyRhjdRXNGXDx4bMTMB3+uW+8OV+P9ug5G1z1ngULKIKaLPlKk3bB2+NTcDE5WchmrCR
JWEUfIUaA7wKu5KgufzyBnk50Czuya2otnH6TvP4zlEyPTwCam7yGoPa166RRfj6hkTkBmB69ZNh
D81gb0Z+sULO7IsyGIwegoPAgmuaVMs2qTbrJ7zdMnWZcTXOXJD+yWZGoWBihgJmCm623f/It5bi
behGqlbYVxZoov1F40VjcvL38wq8YZ8KJIg3eEINwXH77KqyINFPU5xg/pV/jpiwMZKt5CgCQLW/
z6/uDpSXrGKwYsHLShpBvKeLpkIssWprgepISx/9LyNhvFtqsEAZEbf/hp2YO/eVRywQurvuCwda
H41MQvbCP27cgFm2jwp1zIdBi//vMmcIXZolEeGyk26gDkDkANrAwc2es4DGYfrnd6Gg
`protect end_protected
