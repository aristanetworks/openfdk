--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
FplIdnP0YpJHVbhctathqgy4lFCsfciM3Jfdi7X6hrMrySzsba4pGleG7CGafUPOz7f8mO4oAlRY
nrr2wAAV4RxeWRlls8eg8SIa2bZrijaVaZ6knv2Wkg8I9PFm710btRHQaMeR7Xwbe5JBHYKSf9QJ
mw4+JNFqD/ZPacxkzhfPQPVxQAXMQeGfMj32dHDxa+ydPM/De2ptEKnS/PPdrt6IubXTFazGsG8n
awctPL0t0v4A8N/S4tPeFK7hYsXAUrLx3eN9Vc6uZRe7ed2uPI7BMRGjEf4nwnOBI9aDS9kNvdZV
eiQOjM8Kmk32mh0vGzP//ohlqEmkPJP87eivtw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="2En0EXURcavZqsKoArO8K5Eyo9guSzY2+XKWHKX7pQI="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
A2ohwqitaso8qnA6jl+naDTtWRGohv+LM1DWLLcAeZrA8wmMqwJrtHmVayumNF2iBZlvEOtAiZG3
VSkmNqRQwZ2p69EwpJ8ulG1nRdwb5lOmmd36jRlPSCVAnEsI/dAtM2pPeWIgBw21mTJGJX5/bmOd
Xmz6vnJXSGAudQT5bLis/Uvd3kpOwi+Qj1yO59JN8WsGSyF0NhoF9sYVtUt20aWJ3kSOzGwRqKT4
9OPow6vtFLiRGDC2y5qpDZB6OxSgp7L80RkQHQYQ1r1Let9ukVXFSpAGaFtq7Sl56C3P7nJHuZsV
bmB7nv4Pl2XFyRx9HiBYy60trYkqtm43yUn/nQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="TkJNpgt+Wp7+9dE07TuMJWgtEY49bymNeDySGTRqnc0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2080)
`protect data_block
feUY084nEGn4QF4hOnCeiJEzeyhfocOKuxLnqfFBCF/qLcPjBV91FIxbeVWR9GYua9OULfoJX8fa
YzcQRGhCw85QU4ei2F3/nEC8LUEun4NJEHdoTqJ6lkWA9cARPK7V+UBfGWDNH9Zhhb6Fn976t8cD
lFt4tqsVProhfitmIboSiDMLOoc/QRtQYLgDVh0+CoEqN5Ab0bGh5YSDWt3DdVAzYOt9zKKLoG6g
ryrxO+j18v3DJMy3+K5zGk+Qyqg2kS0G+zq4IpLMnhvFve92NjE8TyghV7R73RWSX1kl4wPN+oHR
oGUK0JGjqgAm1oAmmlLxYhBMpWnr1lp7KH/hy91iFMhXMV5MCEqZYEwTFfRKoa2zg6ldTZvzqI0U
LtUSYG/unTyPL4d9ygi0HWhc7ypw83JGINaPjeQqI9t1cwNBMhACip0ymZ+s+3bK2n3zMwyBX5Cm
Z7uKX7WOmgwW+ilFhBSVfHRe4Rqt2OjWr6ZwgctwKOIUOx4CzfUSC88J/6Z0nuCPju5FSVOCViJh
fPXLpDHhl/DupzV6plDLy5tfhpNcdCEAAZ5HLbI1aS5OXk06VLJHobfP6lHHd4NfPGL1gSt+hoiB
u1+jpoQRMuuvZXBa9MGHodokH5jX2YKQSAZzAt2l4sUU5kwhD5deDlA6+xoirnLXOLXFtXZhAjpg
4OqM3nv0SfsRJh0fPyQWehoR7ZaS70LtEZt1icFy5eFe6P6uH+tWn6EFrI+Pu4zKBsbEsj5tuoM+
6vNKOUkTtNxd4xgdh5lQCYJ2nOfsUpgHbfBfljHSVeQEV3TrBOEeLq+t+y6rMDfqwhAzIp4KN/im
Y7hWnXgoy//sLsDxqXH+6v1PMfCeVPZECYJ41kGPy6JcAtjDu/bhUrnHspl/W9JxzBTlTnCyRMr3
vAijZcm5ikuqA9JC1l0+JfttEmUAEh2G42UgBzabdkMb148CUDhhvBzaDXKHY8HGJmNfyTKaMf9I
5WQlYmlm0EEXcyr4a2VFxESXolkEBBxjMRE3838lXkc99D62b5C6oHxrA2ceIU6bJFwxPJbhwTGL
OdP+J7FGrdmdE1wbfaUwFYarRdvANzz2HLajK+VfvhcPMOyu/bLKcpRJh5papFXARNYuz+zKqUQi
oEIva9fx7TgSyDBvRk4LOf9yKJsf6lyERroZFhgL2z4WQs3pjX+aJCdCGEmC6RUJXVc61EmDqI6X
bYmV3zBcJKcrb2abzgI2l09sGdUjadpwdyEnGOI465e2CL5U6tsNbYEHm2rzH7Cn4WcuK5m+t6kR
MWOUYjy+DTEbdl43DSEUBGwvuQeEW2x59XGg9bWBgZAY0eeQdnHz96AdG+ya0gLygsyINcq4FdD0
ugwNuKhAWbSiCDGVSr9Z59U5ULvRIVEEAiMWixhyRNeV4YJldcT3j1EH8ecobxWts7QpjWwENZpB
Iuz2mgHH12eQ9F/yezR75mfB8zXH3+mGSwUnZcStmFLwr2DvY2UOSAQNzL3mUTcrwZ2JHX6wdKcW
/yQpf7CWJEoxsjrWCY/dco5oQ5YrtqgRqVA+DXZuOadx3ouq8pQlSEg6poik2xVsJZPntodFEXZS
y7Agq/EtY9JEtLLOOjUWVvdJv9+wlPGsSKuqFA9/rmRKVW7DiLjfx2jEBc0YUWtdZrWuTT69xLpe
9yxuUXH3nHJk9xWlngqob9SEcljovoEOB3LIe9LrPIw4V/ePCTL/KGqrE/QZeIPG+/E3sh+meity
UPTAz1gaImSWahJaxQT5lj9/FAbAOwi5lmSeH91+jLukti2LqERO7GOjCRFyS0/B9KwlRciE36bO
w1ygqhjnxWmF2SjeP8e1xSkBj5bDvzj2WqUf8zP3ugz/6RgVyYHzP3uTb9HDdECSAiXuJwTkVXBq
J7SJbsgCoaYo8u1xfU68uSxXQrvAOouy5a/bERPvPet+P0mp6LBK9rpCABEHs8ifLw9qUwHFHqyX
MQCqlITgN/tyz3TdYbe6ckH4SErCdYS3yZ46bRDeCh614pxuYet02kEhX4c4LEYuObGikBX+ICZj
XfyclG+nKYEsvsOrzqqoVGlwfiwjbcwL9fpyA5qUz9jI6WGg+KXG0r8wA9CKbdibOJprJRp83F1s
mHeGZXM7RBhrUoHe8Cl18BBbQqlyujzya6Gl4EyDDLWaDnX04h6WIyxJ7PxsAJwlc583SJwAiGFP
TJ/+VgT5ncxVSeLUGNqllsfEgbozi4UQXQVvMbeGVck9WzGgiLr44WZtG+qnsVFxK4wgM+nrwt8x
G6BptMOVYCjSIe7fd9Q1rb7zIyJv5CEW1HXDxhRc5uJZUH/DrnOamY8ki438L2adfnN6xlT2aAmK
CSxY0HcCnXgwmiSlKFjIZZ2zu3qIl2wJspVeaa8LsLTCGouYFcs295fzh3WTS4av1wcROIYyIhFf
nMSesqIKqyRbrp48o2KZC5f6Sp5Ng6cE8Um0lCA6QvqDwsm5lJNH9hop9ekDedRRgG2GLJpD7QAe
sSNWJInjXnJfJ2amLKf4uzZl7rnpQgytOEi+unR+EIXUzxNcwLwtrcQxViJBTEtrHJKa0oh9xunD
1pDjLx5YmGzvKrgE9P5uX2Wfu98/tWP5UbwgIjL2H2koQ5x7GCbIl5yo0YIY80dffWo7rdqxHIJQ
mZBUpQwkuk+aR2EI6eM+HLRKALgLXcbLNdiw0/J3ShmchrDhCYbx6oOdirfEhegZ+j7tyaHvJ+PJ
KBFbBBGmqamvRr1axF/92nKd9ams3tPGK/s3mQ==
`protect end_protected
