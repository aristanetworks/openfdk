--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
E05HeF2Hqfu/k508AmJHCIy4Ubnrs+u/skMHs81YYHTuaXoVLarMBe1gHorgsZ90K/Wi1gkBJwl0
cRmAx2bfb896ZTjv4vtAqtWlnN8wYsXPDBIH/2Y/Y1+ZDD4hu1JdoEz/ZbD27p+sNa+46xw+K13t
LadDg/xgex/nAJdKmY7XAE9pW6hVxW73kfQjv3H0cRw7dB1179e2rXz2x5MWA5VFHBR8U9JWA5I4
icVxBGKIy3L/x2dw+uGdvyz+k2JFz/y6x0LfZzqGJfSeQ2CPL5tapFGPI2FssZXB7Xzv3g1i3sYH
YRUii6Y62UvwcLBzf5A/AaSB4ezOuegUrQqgzA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="gK1K6vxtpyFMxklNBxPfA+xwkw1VDxY5Ck1jWegRNtw="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
eL+OZDfNfqjYc+MjEUPP5qm8qcpTQZxIDysTbfn/OwQF7n2jbP3VI9XrYo6Sc4Lagm3TFglwINJm
k6KBhGsaNb+/gXPCaT09gIJ99H7ALKu9ENzvAEkKBxssP9171R+Tvs0TqeOydb5POVE/w8O1jy6b
UFY5gY6WChZYuRgHxjGgfYNMF9wM/smKvxi5DCBo0D7d/hwnTEvfDA8sTPjruHiYpkaEZnCvvcUr
a5coLacikBOXi3Lb5KRgcnh4VlNwzTdKLCg+ZrrdUGDBxsRSkA7p8B6/prHalPhXq+D5tVg5WxVQ
yR0rli0ZSlfA9+LJ6XFu45hJSx2M5Mygn4GUFQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Tn/dIWD3JvYfWBwa+pJrwYlaBF/M2VP7yYDw4TTBfRU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15504)
`protect data_block
HqQMe5VD183HqtKh1N3+jt7UlfQFyZoBc98sJgZZVjbOW/5ctP2pyByRFb0FjOQE9ZFbKnDmipxV
yh3zfVabth0dH/UF+750QOMQfkRTfW8OaSkyLDnOyHX/RtmJCktBq6HqV2KXHaf7+/7uSb0wQEhh
bVfJzuuGlsGtm7RadaMWvmrSuPXdrCBVufRv5umdThy/DGj6/U0epPVrM3gGOwT6bRCSfT/lVvlL
bzqcq7r6nfiS3KLgD1ianrZ6IXv+PFvkfeSjExeI5HPiewLb63bRWfmazTmcU6uiiuWU0b6mb6EL
5D2MaIBFX3/NCHscECaOSbJpxOv8VY4tOmeykoRy3PhviiANVdcF5EXO6v3CfZXuZ8Jd5QidlVR6
K68jjS7KCk/VcCiyRyfZasSiMYyf6JY7u+RnujOPezeL2JEEleiO8lwGXxKiHrW1H/k7Zz4FTQ4c
gFlMFE3JEa4d4pu7HQdRd9l/VTp+Cs6zJgCGOdGlX/cv7uKhvM28uOrxPi1FZoYqfKhqg+Ci04B+
3HbeVB9oxHL2YZH6Q6w+w97PmZbf88R7lSPkZ8inzmTovy6NRao2ixy7j2ci2vreCqbrCg+rN4TO
PWEHX1DyWgqTvkuoeBK7y4n2lnx5VbSkZTci7ybjHSc+GNWJRjWJJcvAA6kbx0Pb6pezs1HdRpOZ
9keikJj9XwGIQxbf+WqWcfUyi3sfn2C7i/Vzox4ByrWvoYDk9VDf7wFRClRaWyPrR8ij9eNPxEpW
ABz/XEurEahHFQHcfW1LsDXVUTHLoEm7O0rY2zOU/jYXDQyWIfAW2OSOe0nuqWXu8DJPVXfF4DGw
dPVyjSjhLn0UodC5IoQthMw0TfZpqfRdl7FfLQc65FTKbJLo9gq3jDblMh+5OzfrwSoGytPwMeKG
QMMlHU0ozfu5NdPMXrMqb2ad0G+1aJlQY+WEkd8r6X3C/EemRcFKinpEQJ3v0QqEJG6dWRV8ZA7j
XdgMYfjVbaWCzqwNG01sTgcFEF3wepCM/sO9EthC7Ro7sK2XJRmzSKA8oREcynkDxrnMzor7pBZi
HhuTlVYKQ2WQCHPaSPA+s04WltqEV1mxsYxO02oUAUI+Cp4aOlnZDH4xb8zIhFr7N6gn6LZHq0oh
vD+4oc/QFmYs0pRCPE9bFOQ5weRQ8rezeLbZimyq9KMKRWc+DC2QTIZHrtr3LmeViKKnxPLamhwB
+J2NhjOferPvH+AyFa0AzfNL73dzNdvu+tgTmcvG2He3ABxqzgtqg9rSixPugyZdsLdCnJXeF7h6
fYGLAfvcUxbbfPUn7MUopPS+QTy5jA/kDGajtBwn1RLjiOJ9dBMfedaVBxtdG2UGPkfPbukdTyS6
LtIKLWKa2SwjYegpvxth1HAKTiZVw1uF/5KYHSutg4necgC1FWMoW/tPqpQ7nBxK+TKy0tftx1yy
kGqBv8O9e/IcFsVthfAucvlzmj1Avjld1tdeiYI0CMhiFDXjYiPCGqwkFQeE1rnJaDZClpSWOD9l
VGqb8QEOSlX7BDZrhewh8rtkbe8LPJBVx+vibfs8iVnZm1GN87dINfU+C+I7a78LAkfNS4H4xQ+p
+6ZsJBmgVtg7cAuO9KhRFiD/pn7P8q5oYqp9xI7kTsMAGrhSYLbKhGa8/ZFkQsoBaZAJv0Cg7l23
3JxY72uSBT9zA5LF3qpkVcYqI1RXjQG+XJdl8K0B9MraeBFxpCygn2VhDxbMU1nms85Rm/krHLZh
ALyIVu82m+dya1McIjK/Hvao0hayvAJCq9nGmQXDtyDAk0C8/hTFtbrQqQRN/gzEleJ+r8hwzGXf
qpGUhJcFZz8+87WREsb5c1R6NGded7QEAYJDDP33HRJc1UOHUAp5/CYUH+6EUHnR8oA77dhdCUyl
HFV7d4joKTqvdEStv6+GdJY2/13hi+KBPrdUDVEZF+gZuI6gvEreWvKDqmBgLKeMbvCOVAFR8Md5
AtuCb/1MOJdkNP7jmC9eCIruhsK83Tf2zWA2p/2SfEKz+g8jRaagUahd2ymEbwIqhdP+goHPKKVp
6IniECGXkRf0zSw/KvYzYuD1KKIQUuA3n2GUtC+8plJuyzBNgUuuE/JVW5HyXWkmvSaUOd4b9ThZ
QCZog0SIxGbl/yjO7dQ3w9pOXc3z2ZAqEQwZ3a/whRDMmFoMCTvzsjvOHKprtub8R4pVc21A6r+s
b/QThwJQ/z6brZyQUygQh/EcsNXnUPHGULPmXQpgffKZbXkOr0yDJfHhTc0qoQ4UrTFu2k5ScRDa
KTDDA72XAH3C0oMcfKE7kI8oknbVjbrEMoYTcTJn+0kDZy/aFfSFDn8+TgS8CI0gl1e/ZLrxRujx
gmjdiuOsmGEFy2dFuWt6iUvzOUkcsrT99en9J1/qChpv8RoNYLJH52fjkVP5WX4czWabskGEtvx4
IkwCSEGoQYEuCcPAQBaSffwlG7Rxvs80WG+47WkCEtGJ5+6suNIaRgLfXLfjT/pW/INR8ymNqwyW
PQBnIb0cPhR2bo/ZOK1aYwGKujTen9y4Zjg3HZuFe0Ib0WouGwue1dfUqlYqRnKsCFHqIG223tXM
MS5B9+U6tiEWrKMFj7Oo0mm2TPRMb7HYcIGj2CfG2hTkciS8a/gPAieRGOBVoAMZbqEBF+pdNWJw
hwbZkR7e1t3CZf3q/O74vRoyZmc669nmE0zOH+ihw4QO7lkssTzgywcEST8FEh3YXcr/cIliLQ3Z
rfSVwHZwJNh/m//88S3qT9/8NHTSoLg5pRl3vtoLRBE2xpbUnuFCaFkte3vYd+hvImpGOApSqHzs
dxr5Jq4r4N2qMtlGPjNelsUlqUaJq6r2HXPaUVckoP+yVWLXJOBCn1G6QW4fHMqLnYdPyqUohb1C
XwVHVk3FQOFFbsd/ryfkx9PnXMQVBGrZUKQNbBzgie6XftYrP0Xkqe8ebI6se/RTTw7AFLgi+v5K
yiY+fjYyWhmZMMV/KBOo+0Q6bXOfVoGpPZjtpqMVrAOpmyh5mjkTnnuQP9IYoHCsI1KqR/GmChWE
MiDoGJhPI8YUy/GlL+y3v6A00B3bxRY50cjHETpOra+HajEiOz2Z3j613vsmHsulMOV3LgJsZZ6I
Ke1qgpimPhu+px7WJwMRJfYd6U+QUClPBflCRLEebYSnerzInm2R2L8SVsF9GRocIlaUYjEK/a/K
1/k/PkASzJ/cWq7le+LzPU0NH07NE3+x86U8hRpzCvJ7+AmPiafob6Ejw2ZFZgY31kxQ1fw8GTyL
IGpmHqsVj2yX9U9WnywIMyUw9J7e0NOlo1eGlY3JYMSRBfqMQkXpRfNKNsh4+T/MKCiuahtWSq3B
R9DM45bqWw8770H+tUZjhY16V9Zafi1WakSS8wxrrBF+/TYzPiNBqJ9TPEp8Iz5fPKYJr0QN0G2y
f6JvO2xzWhBlJ5Idr8tLqGE+1Royium+QDmNGNI+t0CthlJrxTyC563fyZdAn7eG/yX4G7JClILu
2Owyw9/SeQWoNpZ0bmQDEjxdXfHKTRWE94mfSVcSPUGoTal3tzy0LGCGg0utzfpOGWG0MkpnU6QM
/viaUnRSOJ4CHfcfLFlOYQmHAXnkdh78NzbvQtdznhTMV+qmSwj6wCww3sGftt+S0XILEK1bE//8
JpxBKvFQM5+n9YVCoLXonqkTpAGllmENWzywsF4Y7q+oiHd+mQmYILQWc6AEO2JYnUaq86yVHAr3
fz7MaOJNGylEz+YdtNato9rnmEPgHzux1lw0049JTNfHpzvWpON7E2FH/uvdG5GXinpFPK0e81RO
KvlcrWAOfkyw44lNThIJ/XG62qiZkbEZRTWMJqhBbqXK7kab58a5rh2c1Npxq3kNEAfGXbYTADUD
7KBDHFnGHgFgNsUgEzttMBtgSYD+wtzC/0sjGd7YVO+WPGrpissow0c29L46w2ohJfV5ejkl9SZL
gyfXjIOS8ZaRf7hVlA+dRdG1GbD5yd8YMXtxMGXpv+7okzSRiPk15v0mJ4TC05is6SsHLp47P5pe
/Nx06TuGonTsBxtv3CETi4dzadnxDMue9TfNjuHGiotgoPltMdXC5n/4Ted6J+feSW6dRQhQoBFl
7ZG2lvruFCcRqdelz++Ao6sITCBHWNx2lh5yB3569MvVjr0M7F86N3/CEqPgCvfGu5xxwfJ/dvAa
awe4Vxvq93BVvG/VUESJsAJTjxhcN/6+wYrz8c9CB7FY3MPjn2JXJ5AEIMoa9Yj7QHHI3VtByR0i
cikp8o1NRbCG2hpF2ileVjVjR2WD7YX3NC0S0ZerQFIwzHKUnlqbwMegFrWYuSBGB/zxGVgEqZ5f
zZZvIAXJ6Yny55pq+iBPmMNx6UR2b/Q2RE6GbMxPEkUf9nIuSvFwd+v+rBnnz2pNuFPd8FEluAuL
nkz/wrswY/v/o/Tye+qMcbnD8JdmpCeI9PbYkF7BTM8rwn+HBDU9D2afGbBBC1/sF0mL/U3xcGmO
Nn819trKSVZ8M7MSFWzxLj04qQa4UqofcLQ1GZPvqljq4w5E1uz1Qkfg191eHlsLwN5kcll3Yxb6
k2MslgMv3oZGLsBvA8gVPXpyLNrTusbxnrFPf7hO+KSXWQS2TyC4na/ZoW8vWlDOkyQuZeoMO6Vi
IOXJFQz+6BTocZFbZKsDCXLCMFw9amKLUydsricW2MpRNBsyNmGKOxSjevuSZTcsdcfgPsO1W9ae
yTvsx0xliVVEMCTGjn1awc/yqTmjv+wWC+9dFq9jp+ZKyGF8oIwfAlyTvKBT5QpnJvVL1TRBkL/6
0tgKU4rNXo4AwoAFlLjaO0K/gxDyvnvvBuV9ciKOUnAGbr/FSOFzsIjOOouNMDhobMwD7LPsCCEa
GAxm7v2te1K8uGRyh/Ecmu5mCpE390igR288tHmCzT0Q+AKq36yddSIveRNIICaDF58HrWPTcfxY
0kwMjwI4W8LeHxnTpIpnzTWSNDiy5onFPPBcWyXpg0U8SF4Qe9dbq0VypRczBvge7BLzKOcI4tcl
KbawLUAhmIxZNcSiUHm4jxKSn+JdKc50eQGjS2iTavU9tY1t834LSHJD2guJIWsCcyXugyB7jnz8
uCN2Q+vFBOSyc0Im5aXLFZ8sB4f5NV+ggYI8YZOLISVc4VDBIFGm0kCiYXaHrERrEKBnBm3FiTsi
sFDyOBsZNlSn5QEATiZ81xG7Vg7M8Pkj//PDNPor6osdVTLHh+dPTj0L+FIQ8Tlu7ES1djAWBY3I
8hd6E1VfvDGYwUOgtvWR83fIjcOfbRNfoC1mFi2fMMPe6MXgS5iExfNWUvWWbdj4eDPqjHjErxNM
ms7O2arKVKa9UKJ16i8jESOTG+VOEIAAot6PrdP5J3qOJYvKUDem7qB0ULpCdB55AS3GHaw8fvgk
7JFQtyAMl13D5bCFHnI5sepMduBGQzbUpZRNQd48AIh0kRnyoXiYujH1uVSAPW3vOjJ+cVPOdlRS
FR5R0imrnnd3wRkkIL+6RAdlJ1oYBDhwCrD5EF72mlxCuS8COpk7wFqJ2ppF+Uof8i7fcahdWQ25
BjCzxFn3IvlSrjeJWaOpD0YUUq7mzGKkSEH+NrITuyKoVCODFLwgc/1H4UD/i4PeBbIxk1ws4ViE
DUMzUZ+2xbkm9REjZhaunebpfPvLvwZqTXo7e/FZk2rerh0ir7uMw6ypewgj/U7jfdETMoroAie8
RwPcfrBaX8K3uB0xoAc8jll9hIVBx8UAn8gPZi1srMZAw7QNsUN7DojvNS12NDlFQ5unNcL0Xbv0
IdX/Z08YO5m0OxDop3cZLP8mjPgzXY/vMATUdkIadyj1HMhwt+8Ii3bNCflSucCNp30oWtLP2MbZ
DFtRmS6BTY/ksLChSHJH2DEHDxnXQEQ9TC+7VM9ASbvwnTfMKkBU5GDso1+P6XKoP6IkwgP8EsWi
6++z/9XbJqRoYvTie1/3b/0pleAbdi9YUnNv+FUJqK4uvWqSih+3MW+sS8R/mnNbJEBaRFA91Kx+
dG41giKUKp1mzDLcOFjVeXbhIO+8yWCnRLLK2sQdx3RDo769FGjAtD+HiwDL5iwpLEaPbOX6VVkw
CPgJzKTtHsVkZPTqKfYUkwY/cqSCcZQx1UgJfCHQZBSRgC2rYDZR3/t8WcU+fR+aYZmzbvcsZ91h
63mSx/wO1upOEOouKLq4jGgJSpJ6Kw5IrqpjjbmTCk6Uogiv74FHH7nIwcnwDDyr9ZX9RaxP77XU
SXJveOOjz/kR4RCVFoOC8adNSjZi+GOPYAfdbPjAtoBooR+mHzMDhkrs5v+JKlBbCSVhUz/kJds/
heXbHUZyU+0LH6iuEXM3w9+15aqPjWfOZs3EvKgiM/hXwWnLAVG2JUq4AlKwOwAsZhmh0gfXcbbf
sPHSacyhtoLqr+x8M+XhCJqObZNa9IR1w0yXSHDx1uuZqcE/UUIf35qJk3IAxuqN8br0kagBDb1Y
w0BSfDALOy2Qc8D0RXbPZP8jgnj1myYDiZMjBFcHnTGjNdZ0dtDGGkMaUe8wouzNzHPpZpGJ+R6I
d9yFEOPhr/+7epksbFwAQYl+OgOO2rYIbCCyKa7efFk6fuGowkY7n714H/qswiR5AOUIVUy5Ki63
eEVsx/z6B1RAuUlblKb5wYWAtgd035UjdhELBgtutvLe8hRE1dZ/y8uX6E0UoDDqvqRDqADNyhnN
wldLl55W0jDAu0yV4YKcN+jztR/ag+j4U6GuiEQA+YrTry8rwZp8HZEj+2JBtWsyu3Mr1cRE57bX
lKZ7B/s+n0i+flw1kPbZFDJCrf58G9CE8OLrXuW5Df7CxzmsqtsVUHgYwKdo+5+SVlMuA7cyfQk5
TdvX3TcihZpXHg4+yN2M8xXcjaJhH7XslmrJxxl7vdyaksCnHoKTlSdSgBeHpu1g10+bIb65/sxf
Ov3IOG5s4YOPcRaKIFGUrsIE72lRnznOJxi0adlXiOF9AbjggKTGT98I8Z72FetxQ0+ci08rGMc7
l6+R3aifil8YILX3LUCe5PjXemVJymXeRRbBHK5wrkld8k9AD/RwU7nobZYtLQfxEyHKeH0BWPwq
F7yOg0Aru23t6EnxNAlSb9HykE1rHF9A/YCdnZSfEIo+0WqUb0BDfKzWBBC0vY+iMRma5o0dNRKN
G9A9TjD0e3XqD26cbplKmG0UT1eAs5Y7XaAwMwJFbXfUCKZNhj9lAhIrJgRinNC65R4yrZuC2skQ
3Ok8VVAw7qHtUrL8gk3XbdyBQzxwwM1PFMewasSY0eRPD91Ab7i4wV9c0Q3mIaLMgZKlj/zGNfAC
Tdq/mWXrJOfL0vsZPtr/PksQG8e0qu1AzOtVvt7WNDrq9RKsCeBmkgZT5s+CeZZESvTX7mCAjQ3N
1N0/4wL+1jc8D9CfHOwZxRHcILTOLEiaM9HALV/ZTLoqpjBpWrrMPd8n/UZ2UGoKv/mOhxUvSnSw
dESywGWy41DxlTfrcN+T2Xz5DZiJ7lF9h/wONXP61Hw65NuoiBzETOEertdRwEcjZRHOvdmlOEON
Ck2RPAGtj9/vMSfoTycp8ENnzOon0sRRwOWVkLyj9tmwFaWpFC/rykKfo1ZNu5TyNapr/frmfv59
qzweGHfuAE+UpTaE6PHBa49LQhzC5tfIpWX/IxhJpTSYnMtFvgWkZl59jXlX3cvAcVsPGgJ2/0m6
QTKRldVUXMnC9WRyxHqoZYEerEapD0PglwLkZA5zJW/kTxSmrjANSVQqWcKshwf+ViZ2mdStPpop
nXGJ2TpMFTGwO0g1WRGTSgAMljceR80dK37ATyWboVwd9UdUhARQjCgag1AuO0wBON8YbAudhzpc
jcCs97hSKZbWc08bC3Mlwb9EVP+TnPLjExqAG9a1Zbb35oldY9BqR/jXStLkQvQF+hz5nvzIE50l
eB+MqBqrsIutWXkEuLmLzK/w9JN3pXVAqZd4/jFF2E1w9iN3p/LtHLWAyIDOmuN5T8gH8k/Fwb+5
evd1G4oLLIub8Qai5MQtKKCjUQMcB+tThmq8agoBmJzHKD8+3Y16DnUFmydXu+KXsdPMQgM8qee0
BFEw8ByUAjj0ewO3/Xi5z2k/g7ijiUhyQ2IFniiUITqDfIpOVql6lpeBcAB0c43rLu4L2xfRFiO8
osYU9vHd6taIw3a9rKDqBgVFbF5tYpNnazQEI5Idb7C5MAbMgmCDneQk2fVfBs6Te0Mx/7KPN1UK
tE1dVleMJrbs8MibSx6FQoUwx80FdiObdm5xb6cELf1U+Pcf2CL9RWUpxfrhtOm1JViSz7sa46or
Xz5x8vv0cIMEoXMC/YcM36s60xK+fyIRpxMaotVhqAah6zq0X5cln6oPPq/pM27KRrCEJVXZVmAM
K3jykCPMiUeXzPLEGOV8LBoPDf+lx0S7dZBUd5q6ZKdq0x6B4Jd865d/UevrAjaEGGYAK/36Kc+I
uhfkIQcCJQFEWU7SicPnVRERjZVyJQNTl5GMS9SNs8Oaar/wvAHiFtzrAzPkcC01z/jWiIFVntp3
8O9JzMjHM1nN/CaAu2pvApLLg0btyoGce31ajjhrbqf53c3odtfDUwWrXSQfy168Nc5VWqHQDEyA
d5IwE/fyHKF2US7Q2LEqZIaTBJlW43ZqSIGYA0xjUe9KFLkdvozL6qQyNRJ3W9hdUNt+QKWGtXy0
BsE0hYfjMJ4xIG9fZ8n4nIygJVcLkd5WquaY3GWUHxunUncoSOXIYtv7gt9rnlI+Xpsba692w+jJ
hbXuaN7jiKy0fDF3MLLSpBjXZbkPnaYMgPoFObxoW5eEnTsIXRb9dOnyRWAHCxyUYtULAcQMav5y
xie8QeBN3jqNbdTi0QF9TyZ3+HMq230uQeDPvgt4Z0hp8vJ0iIK1jOxWhalgfq0HTg0osc6BZqeR
7uwOXMCH9aJb2sgjwBZhVOPcEzUXrgPXczGDMJLAffcLB6cyWQ0tz+1Hz1d++xNhJdNF+cd8LONC
owqSzyko80zWMh0BnLwT02lVmpcdqGgLa4gQ2XaUbYX3Y2gD6N6vVY1LO6h5NhVekg3i0ye1WvJ5
1Oj+22bZmQlZPzEBDdBNefYO7WdM9kcfmlXAI4O3rrZ3x5MT8y8OkbDFKad9jAGGDvkM+UDEFnPq
BBWk5z40E0TYLXFHEIT2Q1mQs/lMH0ir0TzOCXDRrqail8SVz0Djjgsy8NegQC8O8TF3bM2+20m7
6QkzZSTxmz2d1QS9CoHk1wBjptwsZzWgCZ/5Ngi60EZMv+8RiOdqYaT2oeK6gHLvUZKLYBhGo0M3
rSnTeg0TLRDfVbkzHcupjX3HvpvpGIe8hWZ0uuoaz3tOH5tZlazhfoX9ugpk0rHEGOpa70xR26Cq
slWjpQ4UyW62OpKcJLCW132ghxhkMscBw1W6DjpGMOtW+g8S0+sVEfRxm3z3L1NMWmwhJO5ixG8f
g285NrJ2EEj++BkbdUYH/blJLK+7QvY0Mt/GCO5se1mgZ41UFDD33RqjSiPYTuzvpiynOLVLXQIW
suH4rw5YuMZ5u5SIfpq/9VPjCb3vd3CCki/YfRzf4p2FcxHmd+q0+ltgANtYGzIQfpB4ETfpJWAY
TeyljIqEscd0wJEu/UYOke9XPV6zbBUyhGjqvyHelGJ0dyQpm7KDl084ep2J2GPFeRrnkmHxnXYd
nQkmSv+arjILRmQk9r18Y84OLC0WObZSC11yDwWx2qM3vjq88LbwxumUUM78q2+8DUMklwqArpoB
yIdf8sWRGQDoBSlFg2iyx4V6C+pxophQLFAdtcXlR6c+XE6HgeaOlypSMofKDt40DV9HKFZa31sX
roRonWx4ZVVOk5ygpQffU85sNDo1svHzMn/GRsIrbKcKVHy2qbNqYy5hgj7dVl0O02nOhnvnMCsU
yMtesIG0U4o9Rsa97ZnzrUbScW2YyPvtZS7v3F1FfHpkc+pOWROFopQSe+HsWwdCrNBX3W7p+k//
gVxsuq71MY77bPhtPokW9xpwIl+FAPVIUVcLeXhnhyjfYojODmr/hqP0JW0Oz5iokJDsaMGPOhBP
XFEX37munQ36ZCQbwwyA/OMn14SpXUQ5WYFwNT77EWbOzNakRkpJfYHb6fRjSTZJP9PDTVSFHX+2
mbholRlHI+76qg+qKYmMRg68alriWlE16DADhxE1qeLCuUjWjLHcCAL5idQ4qAq3YQr674F9yCOP
lX620/ncnCnaiOdZ9w+RvB9BKISEoZZdbHuIf7tJXgNG0eaZLQ9says3I9egllATZZBPRyzhxY76
vKH4msZmthrmGsE8Cu7S3WrUFdsRW8uf7TxpFl9gpKNGn4DISncG7gzh8+ws4dJUx62ZV6wGaQph
K+jm8rZ6id00ild9r4EPN3LgYjXuHm4ybq/dIcNw0hmaB31/b6BeNW0PsfKtLz95Vbz8kI4NluG5
flpyfj8zbODtqZF7e2DCQb0TKabbTQbZCVSBsbpgvh6OxHIDBsAINIXpVijr46RdrYLwzrMwjZRf
FKVGwxEOFuiIAPt80Y1xYk7HpFPOvf/wFDfAjGrhspdb9SRvCwk5wZnukHVkKClcRzb866UxoNjh
enSr+yYgUvOG77JaeZ49av6rG+YxEnOZOf9opc+tqhxT3uDIYA7379y3diHUDvFopwsqrvWsK6cB
/5EhoGxhDuZwVce2PUtf0LzpCYBp5P5f1s9rQs8q6Os9LzBcC/Vo5KhOTnfX0iffeRbV6DFlTm1E
5hBPKaYIKjH92CT5PdITNakHseIUJ3rAiwxoWxvW1l0qMlcfJCpYMiJFkY6z6NI7hkaVzPxUqWgG
VgonCGR/o+oz48ulx9QebYaGokgiHiXUzMEXkuYE7zxjrOcJvuI9lr9Fc4LDEjEH6pAiTU3FTJNp
FMl8ivyCjsAi7lk6CQKGEwqAcRy9Bf+LW7M0OnMDuFBuH95/yKXgdEBlxk28EY3De46A3H5+96Fj
9JatZcr5cKdmKh99HgfIF62HKoQpVhcYbkAhaNp5eUjl6jmRsDalUy1gChUGvfJ2CKl4pWEni6fg
vCdvzXPqsBJGvqD13C3X4l6gbwRhWWzm8ph6QXBRXiCR4GhEhtL5O9YcpzvDb6B25+szxHiJ0FjL
5oeSt2Wud51IUrIT62U1I9ZYAhaWL/UmQHyNjkJtaHxAOMbFNmxPAjBqUUKPji1cKGhrj2UuvsIK
XQ9C1v+/T1F2FD5YDqyvJZ4kFjk69kM5mp9BIHGrgksmY556vuFwApqURIzhk/sgDDiOWZA23vbP
nEm59UaBdYU2lxOkUkc7v/QQ67JAIK2/ZfQqwpQ5v4J1Ql2uXfnuGJeT+N/QRTa79OVJD6qIArLU
XOxcfI8gORvW+94o0JCicb5nJ6Ocy6c3eUQTlyhPqlkNcY4tuZ0IALnN2fEUlSIuxtSpUi2E+vtb
hZXf+GcfZT9JBnrk/Z0MA0f1eoehy+0OQWeZPDN4kCkE10sIaY5gnVk5sF7IIYdETlEOaVoWNq/e
k3QZLR+00T0sgXE1oSab5I+/AMb4eKQKzXNI4mZuGP9oIeNb5fnvb80SvHaE4cpC++Kbb4JzN1su
D4HpfJu7QfkkZP2Zd2A5MyfV6de5UjPTsBV+Cw9lwEcI6nyDMQLWu1Yme3LBoaWZqj2+ibQmapw1
/LtkiT/3EXFhtQdcoMfQAVOdr9t3YrdyDIfLmfwa1wPaVEibxFfebmqhR8JYg4ATqjAiGamHoaO9
0435xpQOo9UXwQdIQfOumTDXUzAlnaeNlIUpNm2cgKdc7ISxjRwEWOzKN/UQLPkXND8VwJgNMz1m
b6eaK+JNTKSAinDtNiwXLLqJxeYhHX9eiMTZZt4X+s3cRu5olPYTre+yb20dRXixh3Mc76QrmIzP
8fLWtjPzh3xYgEEt6gLW93VWKr0h5GxPJ4NFgBftxEr/N8OqDkA2Z0DQJE2Wo+4ZI0rGx4alPEUw
Td8g7jbmFlhyOh3PjqtAsWsZ2gqYX2m99HiW7bDJICBji5QC6hZxOVP6I/rL0yEso/J2XS4y5ggd
lQ0PE+D3nKI9htH9O4MI9+QRStfVKS0Tgn4izQp43okmsfK6g3fvsJpH55E1iLaVcjeOXwih0jXq
LofjZ2WtBMtwuGSFBPK/aXbhro7X5Zi8ofpl/c8Hv7pYR86Nj3yf94qC7v7GEuYwiG7DTm7CK0mY
o25mq+9uk1JIbLWRt+lm2ol+st9Xa20P/XAVMPySNotDzDCHYMgoKfpaQxe90dt6CwhJ4jcFjIXI
ngqkETwrYHwwQCiW0lsXGjgSUmE7e8H3V/K0W0mWijBYgrgopMgt61upz8jYGxDcd3VvMKllJzJP
RBTAmphC6ViAlluwxKMHcEL9oMZYnEkPOiKTaWC0W5lht7E5ad4r2KbCqqmTOMDhlcYJFKOZhWDJ
gDM6N1SuUCxUNirMYDqUba5cqr85mYOloFljrEx7k5y2izrwZKygwzhW/Y0qpH/Ke09HXDTAw6/C
dHAXGbwPl0cofASYQi82SZ4Qlk0Bkgg8FQ+neRn+0BrnpIzke2+aXaur++umfkOecltVkw+TR9gW
Ky+CGbQHic6sklDLuM+z/ZrLPC3luTn3DziLTGRrf26E/SFg1NqW9n0pg/Nntv7ToBVy5DYc0Ouo
GPmfZg1ArlgiIQwjr/ugUkEZIATJ+hyqJnjxlOkHVqv/ciWTh86F4IK8RK2gCMNUJ+cj+kWZ3FL+
Ay79LmUIDFOZdKeIwdXOVVBGmZr1S5SKU5my5YvRIqYI+5uvCwO5xjdQtm7kup1GIEfLnvKlbrim
B57K/7tF+W/oEFGSCgyVHdJnNLpT9VxX32kB14QNLTMwkmErnXswbODqGX0/ZtpFqrXOiEnTKn9Z
Bw/BE3m3tDOe+bWo6+Rzu0PBFzkrIiIpLaO3HpQleYH5XOsC5ljESokSmVDRBapcXqYpda8HLoCf
fiWFEAqSzl/IQ7dd/szQQysLoQOJXqVwe0nb+jOsVrge280EMtg9DEwp9nu8E1UKDC0Fkfq/lk9h
vhSUrG0J6Xs0vn5PoSdR+B/NkogYOazTJQx/dX5ihcT6XD32oVl7Ba9hgBauo/SwKjzD/iEOXU+i
jXXhl6GPRuK+6bLbkpwvbHra91YeAkdUAaoSQZtie0pdTaWs9HL1uKm0Gny+kWe4EhE14G1+E6Fu
eAp8bjWoGNX+6XAjdvBih0Mck7TLklyq+BvD+N8egn4ScWQ5UtnNGyipTn4iluPE16hvsWxDzA8u
VS7McRvB33wMaQCDqNL/9GPoiNCxxopm44gV2A+tWpyed2oCFtDsWEZie2jMOgjPMo6MyYu8Xwe2
n+rGfhJTMUVEGsQVEdALd+/M3ySNPqfizYcCidROJ5bis2M79LVbeq+hSpAI/CvZTRkJhsMAPlmf
6ptdOTtxykPLEYEvL2JUW1nG/x09WZfUlBKIIaPj6OaJnsiVvgcT+xlCBv25wBhjHw+63cUIEyS+
J5VWOY5MwI4+O21PIVu5qy7NCco/uo3a6/veUqDUURfXNnA4J3HDeD7z4pI9Z3f0v9g9Qj6w8Rn3
GiN9TNtc+Ia/cf2YfM+wG3l+Hbl0R68EkXRyYl+y8fSGx03IV7EdUbCTKRfSzPK/n2aPYidiIzEK
OgeuAeUsTiJgDQZ3ZRssH1Loj2GjWmtCh5xvlzfpe3O52C7aKfllgyjYruPZxO3V8bPRaWWPFSF4
7+6EHVk9ouYbyTpmymyCzPjTVtWX/zIQ7oanfwvKyWdhN6QyvomEOVhuUkS66PdvuNLQ6VzGn9RL
gHXmwEdu2FSiQzgU5S3ZBKfAhjkRxCWaHf9Zo7bOlYSuLUwGdaqUHxKlLtw5SkwnRAOw5Ty61ttr
ZivqAIXjzrTDRxZJsj7O9k260+sRuP53ItCfc1hNBiJOIy7LPHtkaIw2zqV/ibEJirH/T17jmNCR
9OkOsd0pywmuZFflr0q0kvP8+oC4XxnZ4SLh+hCii8f4P+wIF5dEotilAuzHftZVAUBLoaSwKjOm
M8vnXSwPlb89XFyZAmXCafnGL9WT6gX2Wmg99srXfebOjX+pwA7tIY/38qRDF9jJWi3XZA5U4hyM
OLi/m2MCxQBLKOPGV0ZFGd7g6Ghi4wmWdT5MjsfEr2Z/J9cNCS9GnochpS5Y4NZJ9VPqmJOqikDq
VXLI48KydHiXU1/3C1e5dmUWrGRw/9QT9zC/HEq++447sgGOjtpUbwEmUKAECEoF1KT6iiIPC2fI
mWZT8Ve888jlsD1v2HREMp5ysigim3uXNWFpDrBPCTdnz92V8Y8r+m0uhzQOp00lwpsUGc44J1JH
BbleNuA01wHmHwFsaxakHFyKByu3m1bw7FAhh8FxYIhz9PfvbItdlyNND5hMYc2jvxX6BoMziK5h
DBZpzVUJr4pFpAwJa9pSi6B5ZkTil0zIRoCdvGozW1F+S+fPwg9Yzmmw2fQWtLLvU35BzgEeABEU
HxERHvQks2RQD3lmKr1ZSL+m1CSrBvF4uXoIq4FVEVGJNz5NTFeBv1WpyLeFqvErm3COn6EY7NFV
SJD5RriiU6rSE26VuPMrbK439S4NtMtlrInHyCI/xpd91PgMXyBDNyUJenrOb84/HAjWW4O+5c2T
6HUvJoGgpkTOp8a1133SpzF5RcSinVGjWF0LBv7VvBeKIeKtg5yvvH2b10FAozfbbaQvnanSvA3c
11/luXtsCavgYsY1ECA1B+P0k7y/RhLGfrYGOqOFAoMmwgrtP4CfbxLcsdP12sc0Y1SItR686Qif
AZlG2hbXrALtcWfrfr9/hK5CsxC0J2KhdWplk32Y3PpLeZQdsaxCLZ5X3YdwSE7lB1606nGccpA8
KDaqB53yBApEE87CxyHIw3+esa4JquuFC2IXuv7AUWBdsibyKeHAMpOLgxVck+ZgKoDu+nyDIuHW
H/Wmt6LskappbeUYd/XrKZvrBi7pveXOkWGqpLyVJvmMoensmmnINrFcukIPKDQ3SGQFx6rCZCIa
MJOQ81jZN1uwue4jrShLuJKehqzRGDLlBLUSVOXHdfsVqKkYnCwAkQ8Z8vrAMfgno67lDNIbje7N
sAmiMGVpz6Vn0dqpWwQskz1i65FJwoY/OoE+DCNfFuU2R7me6g6qEsERBYgPK+7D97OuEw8V2YLq
dwLN+Ws2XKIEiqrp0H28cD78eIaOfgQ02Rw82Wqh/0mOoKYjv6jjHtqI9aIcotCsFnkFH9XAsovn
Bq2gBoFGxc+1LfYJG3kcC9LLSRNXOVFCFDvFVLGp5AMiuLQMYOChWO+HSfxI87BeOI1EeJJUWM3K
bRrXIP7p5QZmcHstncu/fGnw9mFI4VIjjx27oHiFZmZ1KVdghbR7ag4sjmR2bQ7ISQtJO/6BMmaU
cwL6/Zvqla4POiOjJQTTNf91HvwrPa9mGCGVNFnYPoIOjMXes2awNU3WhGyTWFtX76n33v1xg59/
lX77J94frl3yHPS3ipNPxXIhkgh47pUcaHvgOSVV8pyH2skxMnSTqAx1/n5KRlIYIFTHYr+dUusN
wDF3y1HKeAHNL48UW8nytAMYYMnkTbwCZl+6GaKIFTtr5/pcfPNt3hzDPnF6U/cM4qBJk+K0Y8lG
Cll4qZ/1QTezU8F5c4KsDsTApSGf5gmiW43Rti4R/5xHngm3NruSPPwmQguxhNp4fCXoIBIqcs+A
K99GRPgCDWPiOUTESv2mvFkauWnrW+EXdQ5D232gjq/f9nLaZC8rwKx097Vc5fDoZk3EbB7TD8H0
PRid59jY5aFF+njOZ+PtmNxMsZv2lp5ED34z8NigsKHRxSJBkm5mjmCBCtdnrDkUIZ9hSOlk2+L/
QhI2mxxqfM8XsGoWek0CPa8Wp0iBm7cRlsFg8FaDcmxCOloPWAKsklhmUZaa4T8k24FhL9W25kU7
9GnoMKqqSFioqDg73+txW6hTgbafCW2i0pBqXDFcxq7QsDWg7djhrGjRffPvAzhaYeNVyXKcULv5
lOYs5oLIkYk1Uf3npMcYdvA5yUgHETE13GUQgYK9MTRuUjlUQ6vrCGnZRhlvbn2IMbW9Kap9mCxr
q/QBE6G4e1I2Scp5a4CdtSCVJjFHwr1stYkyhkRUfzsghaDmA8DPL89EpOMS6CDYaGT993FNBi0Y
SPiYehmFXx9gaJ3nMrQZKYyK5o6AmtfHIiOHNadgpwbwFNtxjc70kixQpUMCFP8mATZleRlLKOK+
5mGHgFn/l0XjvIbzHwH23wnu/9glELgKP/Kx493jo9ALtPH+iuD5tWTqNIQ/HG3L68VQETm8qAuq
rHCKZ/Xv0Sycw8He0S5rQ5Ot8WBA6CQEQi85f6HSCvxnfogYir4DlxaY/YddRGW1AVU5ED2iiSYd
HNO6Ha2MNpg+2tHG3pmxHULdCgWcnSAybOJ5Jdd/EPYbRCM2zpnFyIA4fzeT6+9+kIaz0YtrpTRz
4zIOcAQm2YR9V3Qajwgpzr8v0ymIjGUPdps0lNQzfqcOIEXNtsyoLqM4HIgYzRRNQ4Aa48rP9l4x
FfaGtRCj+9y5i8Elk/zYml7wOiAvm+YNCbQ3YalkJ1Rk5DXXR1jwqNBD1o/BQB87q6ITT8Pf0fRk
71mSvyQxhI9ibeuNv9D2I9wli4LBxog/Ryps31MaM7RayUqqgpKBPOQtgi4fvVke1yQEqq6/r/83
WkWodNIYNXe1vJjwGmQGI5KHhwCGxXaasvu7G79nR3nTOk16k8l/HPt1p13shdBkHlbxp8XqX56+
zF2SGEPEzQkU5D/YMp1NV1vl5iGt/049COPs0qWtrdG87BcpoaSV1fJ4kpcv3H1BF298gr7I+4em
1sAIEHqANAHm79niu6AIE7Sr78DuMAj3hCpWQMrJE2MUz33aJ6+1LOweTDVcwjRIJKDVOpc7pKNW
IafPNO9eGSXc+fkkKcRyDqEnIdvVC5GnZiSu32OlvQ4EfmBzWvSXEblVOdQfIJztrZ49dV57TzOk
SXydJnIc0tpPltJ1ou64ktOpp56cnIOlHvzNDrBlh2yXx5A+4iYB7BxTa8n0kL9MuDvDXPzkI9tB
Uk+0GhIlCm3orx+k/lXJhmLiilJFpGPk71QKUFY3PyVT27LV9hNQwWhA3Zb8p4mUdOmKZwBjzrdV
w/hKXQsIAuiu/DSA00uDbNVvjFrOjqtXdcw6D00Rqmn4MwT+zGcdBAnR98uk/NvMkGRYw76VpuoK
N75zzVVpVNX9pYtRQ+1WzfMhEtOd1I7ROyQNgPSZmVHNOiB8L9qAkqLzOT2v9KPnhzqKYCz/HHrL
u8CKNq/WeCqSBjDEXf0us9Em3KpT0x5xAZit8rAmohs+lude3Jp/8j6GRHWrYKF6W4JNp/yRN0S4
RmlPjQgUekbQYF13SzLVfkLppcBUh733myM3CpKoI8Lx/NUkc+2v+TLcPM8OutPIdRkrZh8oUKW5
E/472fiLFJ0uag8/vjjDc5CKSJ3xzLHvxzd8W3BPsa2ni8oZjlgnzqgZt7+M770gpTRpqYFc+WaZ
HF0CZ6epGV9bYc/rB384HuOtj8vZYx/FYr+WuSCUTpfyTHZdVLaSZQdjR680YzgO1UiSHv4ITDJG
EpKmlj5jaNXOKyygbQgiri9wvsI07QMN2gBuZhk5BTCJ4iZOJQ8bdX8rXbqHMvgmTtIPzd90MMIR
kBhWyVLln7VuU2IpqmTlgFt3QZSiUSQKai322RmvuUkxls5dt72C2eeGvlLaWCbUQxhMC5+JtP/t
i853K34sCu/TbqgDNGQMxMcqdVZXlqyuEElvUG53JZADuj4j0hg2TOTV00oxQVHXSIhNhSvNjyhn
LUVpnolBlnf4/VlrIGAEWQZDHtBLDn+w2v54+IbxSu/PnoTaxsRQOBiId6fJ6p9DDvjOlsa7KCbi
E7ioaEDfI4k1KWrc81YI8Z7ZM09BFmQCwfMSonuWY/iIPUTFu8MT4Jzbuz4qhv5PHEf3DJBWTv8N
pvNuNVqsYT8Bk4wmwlkacUdRiNm9kX8GZCXgTtsAdL0WjX4/MG69KaVT/FPR1D+avyYKzY4mFsEa
P/ZIIeGd/qPV7FEtIAy7X/CwcT62H2CE5AbTSrhivkq5Qxkh3LN6+j9Sm9sfD6RmgAKql1tM91vI
Hl0XE4cSIcJiGz2hGwCwDCN+nnYwofLNBjaIZHP0IFspiKSV9h2AbvKu+xeufvUQi9LE7tQME8BR
Ynoa8Hl+hnOYEGFaq5WsykRt0Y/HeXJDOgIWM0fxIcHetPoBcO0uqgULDcl/M9/CmDRlsKryGeyj
INbFeImTM5RI1dW1OZ1eVUaR3WiSWx7TGas2tj8DPPiyZB9crGbzJQgMYixcf6WlAovLYvVNpJcX
wMWSsFwNX5Sa2CuqVUNssFhPfPs8jcsQ86g8x9i3YwYwxLnJDLq9VGz6Aofnj/lp7hNvmZcOW8Rk
/4KqrFpz28lTjSZ/WVpgeaiUwWqxhnaNfn8D/DZucCMovh6mC9ewI37tOWBo1uk1ytEK72GVaidQ
h5xvFjMEt4Mjz6scgwCxDvGZUg+mnwQH/3SZcUn9qQH5uwXwANSuKrJdBwoT7YCixDAWZRH5IIJ8
uCaXYEPc7A1fjYlu335vPforTG9XWk5jYQlkg0SAFzncG+8WAN1vV5FG2uo/PmKATvpYCcelZCxG
xKlmaywUgJaXuCmzb9gLnltRkKkZT9Pfmq9S1hUn0pcD2iRxa2IacoLj5CW65+6hnwVRfEdh4Q4O
yQMLUemYRMbwEU2JUEH6OfrhWfu7vFlNfDFaIVyUKwm6DgNc80IipSFiig8Bwh7hwrFn7quo0PTi
0mWvhOxe8BtHMX6KGRwPvIXTqpVvmetBHs1ZdESIPMcW8rDWvMW5HOVW8TyFjZFDMRA7wNpX2cZ0
8bSof/A5iyeyp2jKYHLhYbSmWmcLfr7jstWbl528TWRFFVw+7LVkkzPNNAqb6wASypFNPyx20i3j
PM1B0t2YuVrckksVYjwhq8AxmqipS5eh5P4V3b7Riq2tt7t6QiyNJQx+RVxvd5uT7cGrAe+YCgE4
AZdNlM5GPE6L7E/qQaRM1ZebxBuFE5xiV8Zs/kYfkr6kHruIiA8pvnuDesJIEN8eKLiaX0wnOT4a
qY+XCrJapMRpfV9jM1hSILTuKDW5lCQ/sk/fRbArT4OZIRSzca3yPF1peT548ygQGvDdkQSGDEvx
WT+lmORtXiq90D2yYdTSIW1T4LnFWFA48uImbKY8rZevZ4SHWsIJuAI008Kg+eNPyrdaT3abdvqq
XCNnX9han0fBq39UXyZxoqudBYPPiJJPnnoHXRFFvAyeSxvRN1g4HOK00NGB9WJHDuXkp7dFePtH
DW4Rr2HVhWdIht4EDdm/+bOYU4Mz4HibITSd2OGgNPPRf/67ol6iwy5kEm7EbqVwgpDG5RCCKwvq
pPKNXiQFrAg1ENkgX+YqKOd2AtGA+tTxuwmBRTAN96HUsbC1pdKYKLMEtvNbI2XuhtvSBFrFsD4q
/VEIrqTWMfCEVeyUPtDfhCEG5euKtUNhlwX9KpDXwIqSY2dZlOOlpTEWMgoBKPB1nxOqcsrSWMHn
w3fpjd3T4dkQWgLU0pT9oOFp0l8ZYggPQw893+WXPi8m2E5Ku3DTrxqfHxHXPnUHrazwf/n1X/Ur
BYIzDJshTpefNgaSzbL++d6oyuVOc64Gd6ACtTw+I0GZ2mErE1NsK8tqT16wUMGcg4ZnsUa7jALp
PyB9Ddbzv+W3qtzWENaQhBnOevZ56QBNx91tgd5S3YpmkU9wIyl664AiY3fAnMwz9hArkdEp0mV+
9YDJNUcpO8WY8J7aAI0TTMHr7bXAWC2U9vJWx1et6gtlmIaE34zsuUtDwRFZo3lVRuDUqcRNwa3O
D9FIxWXQfgRwIlnYQHENN+5V8rbf89GAXKAHOOKwGY0s/emcmMbKxCnN/Y71hIXG5kyWNK9uYea2
TCWSms3nR3Z8zb7X276RH6LKtq+NvnkXJZChufeJ+Ts6dgcd0fPWygCwx5MLROUIbVXpVzepBFOY
dxMNn9sH+O3BskRBBf3lney54DnwG3N1Iaka1LGMm4yKXEnw9YKRIBzlBv8mHgWuxbxreN9dSgZI
EiWiUBabbJ7Ugl2VKEJB9NWJaaYhgY452iMXaFRZVDK+pDohuXZvJfpvkhOTmE+dI5VtYZbILyAm
xiCEkJqOldnft/siyh1PDVC5uwMsJ2DkujQ9sy9CWqROF+z3qBcPsEde5mYrN1NkjUuzDZ9ye9dv
XyuCRly7ynftw3gCiHGGsEaJxEYkS+wMlOMoRdqVXH7EZ9BLG58QN+r9tSWm/yJ1gWn0EH59ZxDf
prP+MP5a+RWxql6O1I/HEoogBZnbe2K9AWF1gvG+UjThEa1FA40YWEn1pLZ9MRVEhLClALg29Rah
tm3xntpg67BVSNblZHmXyl6ffVCXU0PpvFxwuQlcWGV/mpwp0194zhKwUGMIOFGyl6YP9avms1Pm
iGjsm5Q2fHsj1tvQXl+Y8eX79PjLdI/37nvnmRGR4riY4uiMZfkoP97QKCmFS/FRycRHvin1qfpc
SJqVM/ExgZj5ft17pTq1H0U54rXWgbNqHO6ZN35byANb+ASOTnngWdAfcRpo7c0+0CL5MtWuIVk7
9Pflf4hgn/jiJKDK+8f3tMBQtY/vLxao0Bvxr9EHqYSk3M+K1MioU9KY0i8/JpVf1jC2IDGdGycC
`protect end_protected
