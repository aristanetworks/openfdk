--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
I6Dmg8KTINen9ILipqutoy2/Sob6H4EnQnJMz5b0go0gZKmKuSAMr36Ri203JTkhu1P3OUUSoSeP
A6kIf9RrPj9f02rxs/VBuU2iqUgFq/rGq7dUIGhQizNh1yUtKXSzMKlAv8XE4eCnqBLSRurwZh8X
r0uFIbGkRD8R9i9vGRtivK3+0BC8xYANiiBY7a9cCxEJfLMCavPpQurBjPUspwICwolVvkVAzI37
6Y9IK40F8NEncehST1c/BGtEx18fXV6BWQipANC/xHR+4M9mYRvP2WnePRZDsLC+S3t3EQewDaM8
b+ewB97Xej1JInT7ynRdXHDxZJvJkP6xEwDOjw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="iUyDwII4a93zKZRsNprqQLeNDWXp4N9gs6WF9Y2b4n8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
K1pgWp0Q8FRVoRcPM87JSrK2pwJX2EMwP1tgXNymeHFXGpOaaN5VQrofRd0dlElLW5k2UplSSVes
wUAEu64FPxlWDA1uyYbuJg+G9kyWEJ95Lq4MUVvXu84tCndDH50UT+yx+42PJtEZzmWxXvNvO1XU
U9bpKO708nW4pqNvDiS3S7CMEFZAsXd0JY9JNMzwQ8zk3XIjfNPI2Vv0W1/c810Go95APnHtolA8
tLOd9E2tKazXdRkNSgFiXUzPmTWkzcsJsAStbXURMvq3kEslD0SO7TbZY5eQ5VxDf+0lOTD4jCc4
+FQqepCtgFXwx/nhOCKgDYGXcW96Pm2vtbsPhw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="iWgrE6MP+2h1/kXufh6Gg+0JbjCO25ELEef+SV48hw0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12816)
`protect data_block
No8G7wSZHUmgMar1v/KFtFREloXWzvD+RO14Wo9tfLAajH0jEL9YeFS3oyS+ILX/usT0qEriPJBI
nRFcbHXG3W8hdW3J13NeTjFhbApZWZJ0BbvhRubw4/a8Y/qz9lkoI+gLNjgW8opnoXwTLagnSlmM
5Ta44C+l7mqb6VIupinPHQG6R9h4eHmVngMbPGYqx0+vgsigk1A9oXsUBGA1J36sdA+qkxTLmAfp
3vW3mgAXlMhP1TaUpRaDqc9sfDX97Fqqye1tkTc8cQlVO302c8FlxRuWyutiR9kXXpqTyd7W2u6Z
CcovATd4ii7AnUfopnBlUsRv+1ZB7ThlRvGYzoQzzSLK8Z66xLb0wkRBR1q94kktSVAVNa9lMxMH
RbQmwDSM+/zEhvhEro1hFcf4yglk820y0yZtxX69k6I0H+DVHB+Ie333ppmVV+7Kk23CT+Bdptwq
qAIgkD7Xjz6q84Ud+Av9Bx38OoVJvje2EUOXlsieYC8fNq/QtXrXg6WxfXIPwatKmFXBaD8VdQ/i
ZZCdkqAFxm7/788dV46nLUUC0Z938rkanM6zBPJyCbI2EuTSylud7zhcpv9rkHhR4CXXu7SR1u2Q
bw93LUfFDH9dy3G+8Matbpb6Jrpy6XMzdZKeRL0ptraUa7x1l3pRSbiUavXP3bdk++p321I5uRs0
DN4p75qzRZM0nv9AACK+noh5DmW6KCxggRAxZabOX7j+FS5+3yQm1QngF4dkS6vUDcDXDI4cLrSM
DYw4Qj8ccYUGg3zW2zYtnhfNx6yimHZ45MhDXnp1fslHR9/93RCZnMffJ5ftg4WHrtDFKJSE+eFU
oVjhLruKjTyrxVwazIiLfLe6eU6Sa39BGMhT1RWa3zZSlTJUUXq/jDqOW1wcNmHqsH9L36earx76
WYYAPNeob9Vzz1QMQAqDlkt3Jx1Soj0rRVNCXgAua6eX3nkYxKCU5OwYhC+Y44T5ozy1RToMAE44
pyyjBK5abjmNra88fqkYgx8oIaVr6I7OC5KThAtmxhIGpI0u7uwaw5qNsk1Kw6nfS88KODgt5v+u
OFaTKstB+yBdlIpNkXz0bgHO28mDRubLrIpcgUSC7Cscm79gPMO3eEM/08nCKwaaZFnS4KFKFM61
8WJN2LBoo5l7RKqRxYfIYGD0yqBseUgtksst1hcMj+vTUJLNcAMxP0BpSQCt9ZRyOdR36ody3Ysd
SrgxONh2sAs9fpkdfjbms/tw+TEmSn8VE8MkNzPC93vRTRSBmCHsXp7oI8CamRQbbDmItD6W8NHO
D1SI2uvK6rsiZMNhW1kAHoKFO3faSHliElSquxk/Clr6pW1vrkWiOK1lPShZraptyBSPkGtcV01b
98gkveMU2LwsjkSHELwddgf33yGwTRi1/iqpbuA9cMu8xqrA+o91FIowq5m4edqosGSW/Wv9VECZ
/uSviULYhpISEy6tecNBENlMiG9A55K0Rxpt8wRF0WA8rY7KKnKFDvlLWjYnZhgwOnpQlKafEX1K
4sIwAkVH1PN0gBBnNf1BLFCOBic63Z1qi/UznXrWso6Qc1E/ZZ1Y4MOlFA5yuUtTTSsJ3I2NHcVT
VRz3YFQkvFdzO/K8uGnyd/VTNjmaClRwBQ1g6jK1IZwlN5YFn1+KOlHjw2ZprIL/arJfzTPBdi0j
YPee2nWW4rwFkG7QWpPYgjUectrqO7ryGA7A7f7pnrfG4uVSt2kJ1n/EZbr3AF0eXZtFTo/TFvp8
6Ngi6cutnsqpbTAjgfL1j4+UQ8NCPLviUJkTR8RmbmUot9oBFt8RbPyGnQIst0PveeRo1r3lOoeC
fRaRr0qeNK/MJuDH94uDsej60ItSEc+OCLOFAz0dvr+rvwPomzRmseB2vkbEZEK+ElPhn4oAXBU/
6BFg+1sJa/bWruDXwjvLJjIFcgAeQlJJNul/BhtPV3Yog7IXxgJqIuGLIzpsYtMfTixcXNYE6uZ+
c08Efd0l+FkBrOD4JhZtTLrGTUed0mwZoPhulr8kHO6/1rFz/rZ79gmrJCLAQgIMSHwIpBEFamqD
ImLbGnWyAkyhCtyeoW/YKl7T/EAQVi2RkL8T74MevwWYD1lxQ6s+KGIB5EqrQfPBHQEe9TWHvFGh
4EJGgdvO6XnsTtQ7fjOaw4kwiRj1MQ4MyX9jzNEpNdeaH2bQtb68BIWBDFXGaDm5AzNKhP0KpWNv
N21UK4FLqK72ux62WkvZ8kSZPJ2LxFwo62FOWtPEsf28g2iBtIWhO7pncn1x7WTEIdUoSGRPHSwW
2y9t04l6XlaKeORdjqk3qn2ERwJNqX9nxpLGRV1hQru16nstiTKMT0dTOuocNJjlFj1MUnOSpqYN
9bh/qjqAJBrp2XYBrQVkgG9mXeNS2tIF8Rc0XKMYMRx/4ErtvX11no8zu8Eu2Wi4eB9eS85rmcgM
Rpanagd3muO0YWkNNAbh9PoBSBKWdSFdQO1ZHjpOHineV4rN0Fsl4eHWIfK7xydo655vfA8FU959
sO9+kUvBWKzhtDmOvLnAcK5lNzGf1Knm+2DxVokUrKK+kaWO5gJPPgTt866CPo2KastHLhvHWN4o
bWLp+T6HcY+BxuKPE6NplfXuvrb4NZAiUH48/e7atyYe/5ljfaPdwXkcrN1n9OjW0D1+eHIdHQ94
q4ogOTyc2oEZV9WhwtJPMwra9/Erv6HmLJQZ2hMpeVnIR8DyEV2t+RWFqZ8OvfVMJItoTsIzDm2k
ZpY9rA3j9Kut7PVDFHb5WN1f1WiosylWtd6QX7TWnp6fXUhxRkB2UAmaWMJEmmTTZJGuBr57YyUc
OjOsyfyHwGUKqLuk6NuoTsgmTvyrdxSYIjIwnJOD5gOmR1e/QV+XT19vRop3uqiLJWopCAGs47UX
qCs4EWOLOfFzqdNx1YT/t5IoYCuxoxqWi7K7s2G0RBjTAzEw1Z1oIBQVpMVVg1ka4Yx1BiOpc2hd
ATj4mY8A0kGomJWWhiq+ImU8wvR8kTmPfiq2HvF8DIsJgzHt6B2QBcT3/+PVplL8Jyd6iYh46/8u
AJ+/q2bJDTOPcOMxs1wjKKtQrxHlDQt3ABC/dG75ReO6cOR2kRKFFrRjLHwezX0lBuYbsOe1PNaT
tfhv7q0xdzq2/UqxZyV3Ud/2yp8hwwlowkK4VOxMYZR35cWiaX8zhOjeUEqnfkX7dNsBx0IVaPYL
6XMxZXQRwyosY4Z50kZVg7G0OJyRGb4jSIk9aI+9/b0Bvr5prg+WB6Hu4NHOnqTYCOIUrh+g5RvH
mxwpIyIp0ImX623gOF6Il9O+9X5RTKygVjCmKjKf+d2ff/kpJ+L7blWymcCZAKnB1l2Vgzo32D5Y
09XHqPvbZ0nHJl52QK7VC+Q8QqEJ/5kYCGIwKkBsx9IQZLe9j/o8vDyWKx5nxRobmqaT/d59V6zx
7Q0FEw9u0GBUR87fypZORmQXBqrcGl6o1qzy9lcfQiwqMONMvmclnBwRU8vUc3Gae1cT1svfwZC9
wdSdTUlkM+ufpDgzIjxzejrQxznLrbxd3fQk3Z8WD3Pa4JtdOT55IaF+BvTa4jFJBj7uSRZwPj9V
lM4gSNjLfUu7ipMFb3a+mKypO1ogAlalYASiMURW7VxLcTgA8LBT5DUNPwlkdDScjPFeRqB9U2Nm
0bxl7l1tUKpwXUhvzcMN4KoQTdwYE23xBnePeOPp6fJTaXg/lFYbGn5xWqLXX5b8YRPvSWxdySzq
OM0DctEM2LBrtZjWasANYkEhrKLrJzC/5f4a5j1SZ97fosKjdo3cC+vzR/JlmIzQi7Uv8lOlMFhW
jommjS/ekpEy5guQTIi3H/7yNe01VVuJ35R0o//EQak090k1Ap2Rb/zYPd+Mo7BIuqC5ASjB/AgF
DqXSipTjNedfSbI2jaozQhloBqeRCvb5N1/lFJmxAFbLl41Wm4zJTR+645M2Wx0NCXn3HQJUR6Cn
FlM9KHawjjgazCtG8GeWHGqDVso5NuSe2x9NoQwV33j8+2zU9c1T8vfL7cibwZDss3NURh96aTi/
gHj3t4DXECObn2pV5HGsS1tqwWKV8QzsbUvZQfog6AsGCvDRz+ZRbiJ2gOaf81kyF+L6bjC//zIu
XmZ6gDB7xCi10PzKZmjxVkNyb6m43MzcWiujnMKEnoYaZ4XWnV7iOPCvoSIXjj/issKHWSDWF8s6
69tOzQzaWR09aQGncpKdKYWDKA4tDIzQhVxVziswiagLLFIj7bEEVr16maSoYrJGOjWrLyIIRgBI
G2RkZPQ4uP5dsOmQTFhv27X6jZ9duN+ZGmFdiXaWXp0ka92kyW9aBqJnRNi6A/N2GGzJ4m6x6Whd
3fkzp1maSqwcG3DXfn1iESwOJVdru7JYmfCycnDmqqk4Hql4txEZgfja/ubJU8Tz7KvWuh/PZbjN
xDy5kPEEx7plVqLlrn4mBEyQK7n14PTX5Xw+5hof6m4Tm/TjDvTA6AExSK/XbCSyvJ3E7ZQB7ygd
zygZCv3Htq83UsliyLm1C4dTof1luj+PyVytciPUiPZC5vZnpmpeyJql7NV+CAlM2DzsuzckSXeY
M8vVbLCUC6LItSDYZJsWCjmx+383Ey/tN/wmun6jDv2i8k8/I6c34OE+bzuJEIUs1bsjQGKlbhsH
DZmXkfqF0as3sngp5/lfuHAaQSEFtxh7u4m9urUYZUZPjjBKcZ+b5ewlCbRaDp5FVjt3cUMXGPtK
J8wVTgCrHWhSr44EDd+lA8h7vOeO+OcDpzLHIMCAELr86XV8RWWKkJ8FyAsJMH2/J+sNyiEFE1lw
8w4T+XD6uNwf9f5e+9ep729/WOGd1z1Af42elYty8/HhK63GU9dGaN4GQY+C6LWHM5T/pzEp9aqu
3j7CRXoKXn8f1XcESb2nXMKDC+AGjUdFYwksEKTU+VH5kiErgEkcdarL3Y80WeA9iUcZ6uM/pQqC
gxIKIfBySoKzh0yj70ZCT0X2LpFQApzt1qBJV9cRc+UtCJFjz5Zf4BNXXmBI7s1AMyxS8ioyOf+Y
IDXicenS3/5Hi7BkwJl0uQMFE2Byt/fzQL5HKcmONa//SuMO22RGFUgoDqd+puhg5fyLqN1WKqrE
QRRbGPiSiDOxO0k7LwWI4qE44II7V0psX9f1+586Z5RgjSFfvBqbtGWCqa/15B4uZY7DosErZcB1
43zKmGNgh+7qXsgBxTDSaZae0tKSGZWftCPmgKt1Z4AYzvXXqCasQInQHibD/oAxg55sIgA7UvT4
XHhfJ5HRn3j4UxNfMo0xdNZhg1YSHjFLTcnC8HuL6FWeR01xfx12PUdUYT4USuLyKACzepmWjuGu
v7e1EBKfa5UCfT6n/Dhm0yYb90gU+4FvhnmD2XKAdrshO1J97YfogGMNJhFfNgtzzIKUD/RCj0bF
HmsJKAFluG3G4xEOmau3kbKnEfeXgOvHm1Hurlz1wLqrOB+fhkPKq0RHo5Vh6gQ/iOYDaEqugn0O
9HSMt+to+GjE2GaakL2CXp/8niP8wAVIlC0UEMkaKQLuAjsAzXw2/TG3d3EIa73mon8l0tGDkfRX
YXIv2njIBYtdf/o+pcC7l2dA0d2M1+ScFcYyL4H0KKmVgtLuQJ6nxvZH8zG3sugeKY/qVd2pb26O
qLob+V3bqd7YMm5ErlYvdYQ8p6Wy4RyJ2rlGk6biHGImK0TEuW6QQVIkPZ8yxoYsRoRy335J/Un/
vm+54T+uknWjkY3kA5fvDop2XRbxIBkYE1JlCtMDb1r5qWKjBcfP/ax9fsz6U80rs/ylIt06Yvlk
GVFPY+UoqjLEyTsOI6A53Q5GdxYSGu4j9PcFquzqVC8JS1HOV32Hr7GjP67CcuvSqVzXyuvQJSoh
bJrfEORzsry1zz5xdCBJvoebnOne17j4eXSmoyKy0uuPPJc6KsixMe/yTb33T93I45tBnk8x0osh
XnTPWx/sdtWDlvmgr/AhM0vIybNe6bCtoK95PRK5/nMazD0Qv7ApOtCum6bX/RKFtdsLeLuUdhlK
3HDNp8RtpUdwB93Ehj+xmcvRZWx4wmSrtwbzgfi6AFWqq73KsWpJUuSTThtxxlF8wuN/oZEWV5yL
Lryz/Pv3C8piOUpCaHjNYn953r4R01TdXCgRBlGo/cMRJoGA7lmqYTz7SQ00rJOhRZPTKBrDestJ
tM4Gf+jVbw1O0tmbAcwfDsQqkiRzMxj6Qemve9BcV+oJvnKt89/onx+ZEUaX3P8r9oL2cgafYVcA
k4JhFNffNhgaUmlF+OPnRxw2C89rjPdkVxjUXH91I7zgLisJAxK74fpwlA9apaHMNqdDQIIK8E3M
rpuLhaFPih1KzHcxjAkgn1ZW7p1gd2YDc4/ygoIpvTwbiggG4yWlxEDmIPbfi5vq4104+VgaZyww
TrbuzIJVFS8wtuYWvHAUKDl48FI1fDfEBrcMOO53kyeOvC7Nk048fyzZPrzwRnt1gvugGSOBrv7f
05U89Ws82bpbLOi7lvDoWCqvNh+iXlr0iv3ppH3qxAlvc+J5zbHqY4L2uEKTkTmGy9/VDA4jfDo3
cQmUhenI9/GxyIagdKTxXOtpjl3F0UzTGYnst6tUXAP1mnX/SswrJVGp5hgZ/L1lw37d2l1XBJpG
Y1UhxNTk1Xf4enDEIiVDSgWs0rwzu86TG5Pn/WsIPiNqGVEIOhPEAnVw9eSZqHU8O7BazzIPh0p6
pz+1ep22xuDTDEqd8ALF251cSRbi64KdjXLckCnBU/AmtmTBv/rGlHVT6iq6G/Y/YNpR4l6x7ZWR
fVoMiwSrrUV+TTc+qmSibpALy5kqbEd4xOhNFNNpf2I6n+oI28Wbhd4yXqWTqzR7l7nV24f7BJ3X
eUiIxjX21vwKX7b5Fr5GtLSFwWqWtv3IiX/cbZSnbzKcuUHuq1oRxyH+kC2SDzuKViwZXsBH4202
GDHe+2pHZPKOagoptJ2i3YLY0e8TiQKfmpwcOdt9o9u25MkW8Q5xUT4/dz5Btkgj9LbDH612bKxx
tvcHxzYA7epAMaRRC+AhI+b1NgUFsC2jIQAbrNMnZ5UOIxWE4CrjgpFM4HYA3sVAnGG1SBuOYhEW
O8T+lKo0W2EIKOn5gxR16xO0kHkCail4PtkW4YxqF4rgI47/54VvGSzvWHMCufPBpdRruztBRGal
ACMkkt6ZbQqS2FDvhfXfvsj0e12m/Ek8UD+w8ycbGvr4nCx+dmzfOHUOH7VIrjYLnKdL3uEL+VkG
I6FNavyy8K7/241HF3ykTzQXOTljE6DB35HYahrZfmkMqQQifiP4IuLHv4j038cqYo95LMpgmGKr
jhLBcm1hTx3i4/8AX5gXMuQ7Ku71Lm6ZPoHSs599Xx9vkdiEImrbbYuHDivDeal2DLE+kLMEdyEt
DaGOXrneGGbRgRu8NqU37XqOupiFo9thmOpjOTQdtZeibdDl67SpXfUUDSnfOG3dM/fwFMDsdXnX
Yaa1nbWuZw0ZJ3oYwrRk7ahefgheZcV8rOyS+kHj5YDimDyV8YP6wPFQnqrzmkn0ubPETdPUAkSK
tkVgJCqKb/locSb4wyij3SwUIK6W/D6EZ0AJHxGYKoz9FEo2M3VKk7elEG7aRTCyYxz6XaRBchLB
jkx0mwLnqdDrHbzb4km8rFqgvoLq6Yk7ZNr90DTEIFu4paDeCNdpU7IyVduNeUS6ll1Za7IRYby2
1F13EtPee9pqTeNcPGSd7Aw8XKGCDgxl12vVZ4F/C5LYcMOtDAZQPmFrRtZCr4em7dukIIp2ihzj
qcGxp434+LuTd5x6zAi6foXra+CX1C0uhtPbVe/fvPK0JhxIWpT+eA9WTpbCfNZ3ADIqJyxmzOiO
busWZT6ZZskikQCjjBKxARLrKSLDNw/N19I86RNjbRmygR8s0F0J+hhYpg9QO1JvfFkAOxLtd0Yo
K0ZEd9noY0JdoQaR2lo+gaXI8Q20GmrYSB+GvnxCtn2K7lyJrf8ndl6B2HFp+4Hv+3xI5iBTiH4a
klqP7Y+ELA49e2iIwEmtZX9hTEGx+QYeANx7IlxI6HuNMElLTg4rlnNszkv9BZDOjlwm0yr5rC0T
zs+Dkx4vK6LS1/VwoOtzS+QrobwxjvwKD78vGoO0FG8l0Jj2QRJsSrCxw+AJvQj+qpVTzuejI/9X
vlAxrzCXCGBgvvGLlnkGqLtb74HvMB61zKIVKCBKpyTyLp5emtBNT2wZkHWJ90D3vETEMQOtZB5u
6T9SViwVAgSR5TnNIITn7spjCpyoPX3EFrvJPGpedf2TjR/DJjmuE4Odytz32vHwHoCo/xhLKY55
b87LZ6fkyJ9wYzTiiJt/WCrlQ+lIHy8HdlFpP+suxWowjVB+e6gYv3sYSJY1NrKheLJRWIGCkd6I
tiDcQXMFAcfZUVq5+In7KKHMc2GNY4DS5Yk4kPSpF+Ck3xh5T+ULMe0JJF9EwQDvc1CVBH+56tTh
eC8ziuD6izaxwbioGe+3X2p7qcEDDxui5QD3uCtvKWj5rWAvQ0LBvwhWvedZS9ZCp/+ZvnhDEMZo
OBGglxq1q40diEM9FVljfxVYSg0roZZt8IwlKFEYjAxQCoz0VuE5pgLasfhwVn0cMm6g70RpA6jg
KVD9SDK+UDadEuVpzG0HUjS2FjPJ8AEW97IFXaJ+NoRxIEjrF2TPo/Zn6m6gnzgsSBAb+1biZEEu
uOz+lHIgCYbLHyZ9zK71v+vrEmt+kISrPENl4Hsv+lcBzxDNLccyGA9Jx1kszr1XkHJjYFp3TNhb
jxdH5aS6l+HSkIvfsyTyKh+siKl8H9z8W6gwidsX/AkzIulvkxvEZVWTolYCvRAMnLFNIzqAsVIR
np8sZ87mysGlQfwghx8pNyoNbLGSWUQeQUqARDAHjVjmmkFEWVIOzvEkSOyp8bp0htQXRZZbVxYP
6ep/BCrNSsSYHiHtANHsFUrBpkmhyj6CYcGicG2LT8gO+zYit70eOUFnB9j50E6bZgvHvumNcUMS
4l56fnqp5fhsw1bU4gZTC70sSXg2LGkYfPzrfpGa4lgMhLJKsOzI/lsc1WgieRPC3bZFwNavF9/g
3ws6/wZMhlmDPpSi3c26hN3CnOEa3B8/aLhlUOJGET+tufghXGADt5RqkDy5AWgaxTqXH/qcd4WD
+VXQogv36Bt22TpgK/HuTuyiZ5DeOsgFyJOjFxZptE5K5hKKFnioq4bgTMfG/JsKN6Zp71JnOkOz
AmIsJduURfWcd2l1JnPfSsU1yogVw1NcneNJdHSZiw4eeBOhpyAqm+KKtyX7eIy25KbcefDP4FHi
xxNWoLK4ex6tDM0a0QR9kjv7fMaQKWmGmO9u+d0v/g+n4ZjDgvePoIXgHcZfZ4mtt8zekjad3UTM
QSDMtu/Qw/ySuMGEWF/PSN+6DAwgatBqHU4Em+pP3T2iSCfMb3THkjjwbtEUduT9Zb5+rStMjTv3
ezw1wVIgqaK55NfsHUro9CQREaI9gEisRB3kRqQBnmhfyLgiTWnZv6gZTMjdDOyy34uIWSY/7fp/
z00Y/1TRrARKpH3JVcvVmcY6f+9HbvOvoQfoFKblRp+YUaGtrGNIaFqryp+LxSMH2j6zSnGGmWgp
Mohq9VhW43UUzeuTJABx+xeFEwBnMwYS7u0BprSSPmA26RIpybsCdou43BXttpSCQrKzIJrsXZhK
uHWk4b+hyyXVsWliP5edu3hsJcUsN5oMgH3nG38Qiq9mqKvdSbu+hqnPWTdOYkZSxtxEs3w4NWVA
QtzOKlWxDgJwsBULA4cLnMAyaGx3vV34FFuDPb/RVXTOA0UphF/ZAfGy5XzHmlgtDRU195GGcCM4
szqE9zENRMXGK/AxNR4nHSY080p4N/60mJPJg7/SbkP/Exl4AsdkRV9QC1qFLO/q7WKRXzQXVjiz
G6r8nvfki9EPvgL7ZIWkz7FN3K7EO1C/2lRzMZnOT6j5OVyl8cuN37rKa0vQSSEcRVh4swFsaStG
tZEUai2XrSiUiTQRSeM+N/3vFUGxRH6joqm7S0iYARPiVjpHvQvta3ymZZggmTkYrj+gWZXfYis6
2IHEnzYdiMBdjWXsu9M1b2a592oRjLHXAF293ufAMh21FKnppVRVVZ8QdO8v3ZVv3bHbOW3E7Kd8
JwARQM+2SPjaSebamFOGFHhmpRJj1hgPm2QuIPTZPl3pwugjIT9D8eu1yjVESDUUqdKv1120hCQ/
oTOlHpSwMmxAZEqgLfQE4u6pjoy9jnxP68FbUUZeKGXX7dR8E3n4cxyxwbN5oXX+N3zD44nHEtgh
sleIoS+scxsD9rgawfbKawqQRmJEeKCvMZyGVI2L+fSVR/dwMyvMPr2XMplHGfP9XnNhIDqOsGBn
7C+QIqBtgVQ51qExNqe/uzRsF5j21UtifVXLHCn2txLO6WLVrwN2Zjq/Cwd2Bt1KRlAo2HLE72e6
C1VFYU2GdZPbBcg4Wfvx97bukzD6SUQHkjC6sS8nQXopcnd/0IkkzWR2MGeAuwM1uI6cs2WtnkGi
jcubOkXhKvKPPZgSsQfRyHSFZEQMaUQfdFPZeZXPlXD1Z+5pMaGHvhv8gpQ6rJRK3R3D+4fcJKpl
XF8lmjBCa0IJAvfYqXmk2n3Etx+LjD6okefgM2xT8TBjqP8dwbh/GU1vPVlue8LgrPp/g3ivHYp+
PNr72dN8QDLDFVUI+oRcF55dGWtxM3ggWt+ZL3swlzpd4d/oF+X6GtKzssoDUfEm43WJP4U7jgWr
OK7uDmmQ120FAAztycFeQ9GYRbLauWLyrm4jFEmtpedsxA24jEjBuuowwz5w69mXHlq2qtRt6JqS
ktgyRezK5tPW1Zuo1fblCx8+pOUB66Ycwtx2eBgBn0QakbAWLWgawwFXfhrImdVJ9ZdR5MVWzOTp
6SB4X334ZcpB0xWt3cwOZVXE4uZAvth969EfUwKs/LXefnA7zQt8oKqlp/VS/fZvNedzHCbQceel
RIfwvlVlqWu5NqHULEow1RnlJEp6tkYcIw4kd8A1f70ZTdq1RsL00rgUSGDiquNZn0lSlWEbpoBl
YyDnTuUMwuka97pcURqo6AX3LFqbHe4BkHpGgMJHo13forXPGkdkFQUC131LB+twGo6QZ1Qb7CoN
uqra2cuKquhO2mmLvRK4IVB1SgInDPpW4U3ZG6mJz7xn4HWfxoiJZp2nHm+Nc+fF7kz9DpBE3IWC
EqCdzBVcv0EFwAcmEbsKIpNUyaZlLWF7w2li6pYEYGNgpjCHCZDdyp/xX0MZoiBuTFhdpfaiwVUs
Ihibq+ywek/LhO+KD93hRHwAWioE/QLIZKmtqMfcMyUrAUSgaPBWJziInQRBUlod1Gz2HbJXa1D/
X0gjGFLllE+e2Z65qnqdd1oG5vvLHwicz1kBJO+Gya89OROT8ygMXa1qc5mNe9zd8+zPEE5ahrTj
+l5xqTQVIYJtoxLlFYUCWksw/oYniOplm4a3UZbUQG5M8jF7VsXHlZiR2OOXHdKj5gPoKwqc/Wty
V3X3NfNVdCbqXizrcBRNKCOw0NPLefFjHnHRlYxRBzhM3tIRaehhi4BM2qwwt6WxcdnjWqcl4cq1
13TssgjmNauF0PY27lqCKNtzQo88njPhG/sGBCmzMDaCVk6dl0tFlUpGIDJQyxO2tYz+nbreNcpr
b6g+u8vtu6VWPFN6YkLXnUNsPgedh/6BC5xXtDSyhm/V1eGu5EuAnSopVxNAn/+TaX48mmTeczeF
qhFOhfE0iii5cbMsdSRBZfKajMWyUkIPbVIw3rYnUdywUAMSQrRBjH4OtqqNsVbq84uwQgzmWRxs
CWwUYN++wyqdP83acmnRM3lLPcdwF9FaE+iAP1sFsMqBS0qs6yJDFmbVLsmycCXW44PpWf1SNg5G
gz4HiCECHQzGVWmB3BI5qW/MsmoFv7IHqY4j0KAypwJ7leCOyQzUaVQsNVEIkgWFDv6iGoYySQg1
1Z6VTxPWrZ7uAfl0OKNAEBhzkp89HdGTb/apVIMo114IvZA9KlL1v9OkyCkDJp1qdXdxp8gM3DdA
0VOdpSIBqc2prLUIohDhR/FsC2k31OY36++IpRU86LVXnev1zn7UFrWLJAMg/iaoz8cpp8n5hiH3
HbpgIzd+sxe2uVWXj1yOIO8uRIbHC4XJd7ropGWk2Yc+JrRRWEMBCx9aadRYTASXXX6mhzSB2WM9
sVOGlfIl/BtXc4K94x2713N7E52NWkpUOLPDr2D2JnWP4K4UgMbvMxffnV8l8h3lpT7+4vFZc001
FAlPnUOt3wOL0TCrAuDDHO1L7yuU3lLmPOekQCESmmUkgl0I9RcUezVPfGzdDyilMj3zL+eWdnDD
+VMu34m8fHapiFptHq3lQ96BjVhVzv6b/UWdINQeD6e+/2ldW/0ngQHC2IB3ZmX4HFyl8atw/6EH
MkNPSfx5Sy94VgLMO8epffBC7XcmYc4rrfIHhbiMuLfN1j16I/SM6eMTIfmQJxey5lLrgk11phE5
ARekshQouQDJ7Rv2V+B3k0deuta+FzmpGfKko6ZJ9VipO9DgHau416XsO8edN2sHQNqh1ml7i4wG
E5GGuVurpNp90lipH6R7nIQazN+lKlZxj4KeVma6XK466FvEdAX9mKhG/6HjGECGs1nhTLNBvEey
RTKFeYwChZ/3oWAaNhIT79V4Cn0Qi/QOX1eTt3w82yWCg/dZZgI7QhJhfCwsahIMG14yXgQrd7g0
NacSeygKdINgMWG54D3tfnDgRX7sbKxhIrRrpp+XuFIXXVZKkC5nURMubCVudZDbE2xVXFJF0HOX
mdg0pXnTDxIb8tr6ymDEM3ogE2S4eISgbj4cXeYPnEg5ENmfqPaXul4zv6hodQqLIG1uKhHCxPK8
27dFYhh7WG8oBdmxJYl3L1WcyAleEikWml5zkfSt59CZLGMdDqJ+YMOVeDXlTA887GJ0f3xrDIXS
5QytT2t2jrqY+it1WCG/nX99DxTP9+veGeqYK0JOGJFOHdLFEOdss5AoMgBC660dXZH3jDtqnSmK
19fbHogdAiSUL0sTVCXa+uBRAZiP4HJ+bHRh8aA6tr6fwz+EyWyFrxhxqMDuV7bz5zY0wB3C7moZ
7RWLtIP6wTtpz93/C13GdXOv9SDI+Me/MXOSzDVj5mIw5hymbeu+muJxjuPUDoUQv8CLGDz/a6lM
GZHG/hymG2UHiZPrtVOv5AqXtQaQyRQJBv9PP4KqsbzQddFkK0l4Dm4Mg6ssg9ll5zdtN/LBu78c
jrp2/HeijyBtRigwuYd2KnbWoG01OU0sy48S/d5asHwaG4nPmQ6PKTevxxOD5eGKHedoZBMapXB4
DnvZIpqU2563OqX5xsjVbECVfS11iuOsoY7xLWMOGLbww4gGLw3FC2rUlTsBt8DNOZQCRObYXZXb
4KjtftSxTxXJiUDc3KP6VUFsdOqVzOQ+jm+La3rJTdS+YyCEZLivfKsFezZIAA4G9GPqflvKh2Jd
qbgTDbmfD0B/hRDJOMB6fkbDrwIc5fATYVjgC7zNeSz0H7LB5f0mPcomSriA0VXFy7qbjGsvmBmw
g9DydmyXGx6KzISMbeOpTu585K5Ar2AGB1Axer/7qg6ff6g8g5MmEeTKGih+dY1CppZ5KVkEtOFv
Bi0uagbPnjE0t5si9Sh9Hr2I167XJDNECXNT4VRoD5WbR7Lzi/S8SAkqBmX3HIBYOGJBXpy/Ybz2
eRKHNNoq5gJ9Cxv6ZvjkYi5/zkwSGf4W3hX5vQha/QssJCbXMq5Wz8L5bcMnkWlOBqQcrUOZET6O
DUXnMqFuzMWudNR8aEAm5c5aBWSty4iI7/f2n0DLFZ7/XY8dAnNKiwEwNbdTXAirkWPj0RUIZ11Q
t5znzsnP5gfOrBzVkvC5qJQqnmfEwja6Wj7SXSL5RHiAzCc21QpsgwKBQgdJ+Ji+OUba4vGzekOi
2YbXv4Ex0dJSPdKdzrX4j3uREui1EHnp37Be6wU3MjAcTVJQ+5+KqoJOIRtKbP6wU9crHczgK+4F
fZfCOeS/pa/Aqs11o2IFv4mNfG1rJmRSse3BFUy/D13+FdO2/tzWryedv63WAfn6m9bi1YdZn02U
8XcnqAfmSoJBOc1S6WLicJtkalyIfH7Vv1aOyUwK+hG5QTGKk0aUFv5JV4C3lAXnsnH76PIJyrCO
9e05MP3jkCUBWqvKFIu3ZqL+Slnmek41SV8f1ZQODNBUwDgLaoIya9LdyhKeWPFWG7TQ0cTEg0ET
/hPtpPBnQ48v2PafK5j0+XFol7RIqIIEBVgmE8Q25pJMAGrxMgYcultLPdwh5KDZ+sQr9nSRFUlg
Oa65oF8h64EM/+bbNlLGWiaU3HBFDAreMZrQU+Zo+KQ8jSoQPpfOolFHTi6VlYaOaQGVZBZ49qR6
zgMglVwgTNnYHE/evwYtTvuXf6BXhHDtEzzfnk8Z/1yIv4zBVp/qpZkrjOqpcL6drDt9o1Jwn6wy
1rnG3kog5ryM1YEEja1NDFgkf9tXYbXt67rZtlXm7hxUDfa8sI1GBSKooWbZdkOsOaYL+CAuSrVy
6ABadJuWPQg+JsVRoTXI6X4YN06BHoH25Kf7n/NyY9ZibZX4XUGF7sBWfBVOOdLzx20Kyv5jyECY
gIf8rjUQ9f82NUL5jda3AXCouOHq9avPVnGUfHI8TkgqcemJDQJNAM716PjAX2Sq36N2O5QfYrNm
yeqy4flsNOnVdCuJIZ4G+1gfewv2fHTXqs6xPqwj3CRdoLbNFzY5xhxyNDn5Pw5jdev10QvSeQmb
9VNze73u1guIGYTzRZ9UmNh0kxSpHlNhhZyuAnhnY+Vgns+k1SpdAz6gYTLb+wS1nCHwwgNkAncb
UmvyKbEXDE6nuF6ZIx300/29e1dzWRr2oqEJ1/6co9TGTU03FIRJxVRF003RY/TYy9XKuMGicQIu
jhBJj/T/lN9zdUdox/N/6J7F83omZ0Q6Yf0hZ5WkYJpfLsXPvzEj2qN2CyLeAkdO81AyTlzFBmej
+xMoPFfLZ2UPjsRgt9CzWyzsgtYdygKOOBTM3UvSOhkscKy38jAHWAqqhJAxeUHuSQDzZiCUY8qQ
DFU4HKq772iHIqgCpt4ZFOrB7d1JeTk5oc7OBEzDIufrMVzxreMrCdTORExzlF7lOYfJS8gdihUx
JAA8QdMHB6ixAfKGJvequmF40KAH6enYWadGQglKpSO6xTVTeMrRT+xTqY/dhZguLP7i94IEfa0U
J+nicJTKyLN3HJs1PL/A1reKhcYLxpy5r3jpUo+q8lBNlGoiReApziioNxYHjw+rNYwdaASK0vSf
JRw+KfwBfn1NdbwF+TIPfZSnM5NAtJJrso29lUuQbc2AklPYMr422ZwT96Go5L9skEpf3ZzMZHan
BJMROck6X1b79kceatpJhqYJybZpR1Xu/JDP4qPz9l/Jy8YiAcx7QdvVklobdJRemvlZnAFpccMQ
90HnVDniVbxmeuP6m4oU17Gv+6m893bmOUJnMbvv8YtHlS7wXd42mk+7Gd0b3TQ8EqNrLhqDnDpP
FYoJ8hoP3fd2ecOwFs/f0QvY/D/eWtuNgQVl1zWOyc5cCMuZzvwPFPjMkowzBleRmnce3K942rBg
A0btarwjQL68ruF8JlvpFfkt1AH88qoIyNl2wF8eF9ZO5CcFUsZRmDCLj7Hdl33phufnTB7jId4h
ImGSwzNqCg/Px3iavvsmuntEFznIduNnMAaKc/3bTw+z3SilXvlcHZ5vAlFE0VfPnqmIJn/9S5fg
vMZaA97J2KsMrJlErsoysbUPETqTBwqeKY1FBSVadt5/Y2GpoME03YQTU9MA21kj5kcCfiht89KR
FahMPG8YGlGDb5iYdraItXmVEWyIo7cFqy1G5edYxcWqqkj2qpyz6eT+OXvUSjY1RTgdqEf+OSfd
se8SBIEcklJDMb0t8YXBdfn0nyxNO1VAgUGuxlNALgQhf5RZeLsKYg3JVAajFCMxCEtQk2qPNzQR
1bD6XlWpTrDWWfU0YvnGvv4H66bFnxdmbACZdoFcWBqPMsOg3GunQwyLGC/R9v+WoGe24f+GkJM6
b2wk6/FzBO9LEaIDpv9XHw7zZYD0hxkxjYYRjuwqy2ry3CCtenlJPA/rwG+KfjgDaknB7rw+xEIa
bZ/HkLW9Nsc9mD78akrJpnrdnxSIZr5HXAlPwjaHkcrDOtDTU4/eZc/IjNvZyjS67Xwe2bLGHdUJ
8e+YDckB72UI9dNtlJWVfrxs72kg3bxWqrVbuz7+Wdz2ttvWbAqb9cVu3Umq7QnmjR1B7kR0fHbU
9+utgZx7VvOP6jDG06Ry+z9dE3Wl/CIBUNHuqk7NqhaiHuG7OlfxPDb9pzed/s1rMYzsSERDT5Ck
Gj0OCnOSku/60vGLTzGKshL1TcyrsEThwWy0BWwNMmlJct79NJVxj8VTV1zxngBnh9QYbo3HpyLb
d1w8JW80KMW2TDbwiIMDwMTHKelT6hczXW2nfuDyDftQ0zJAgaTGfYnoymBMmrOBlJHK07TvGszw
1abv0UfPWNqYuz0ArPpGNjERIP7JGh83MUoKPrtPgW0+un04WhDXhw9OG9PAa+FU+PIVk3W3TjVi
okR+M5VWBJZY0V28+n87fDlARismEBMjyL3ILW6uxmWGQ/X10c/BmjCnXl4wWw2pHGoDtkXejn6n
7INRVRo7zzXNCobCO6pN4jHuuNmhW9qTNjQL/FMqN08/DHArGSe1dmxMQCuUtE7ajYhzLiXeE9Gg
zejWrlQC2hjE0Hw/4SzXOnEOT8Ix3Q62GR5GBf4MrsKmLuIb7NM2AwRj2k+Lsz9bYcqlPaeXj3VU
+SQTMY19dx1npQ7J1IvHL0gjDBXeheAORQdpW+UC/GQa5htTpEuOtjywRQj8M0Wh57MRKGp8vxw+
RMg4AGoajz9rilVaakrzpAMVtpBcPS7WLj+KtVg6zzjJvlu5D0hTUX+0hGL6tZevlKkU3tKY8Vya
pHVmsPljc0rGzdDpcdvwscp/0qYKZcqOxUfkz+rFYSkS64c/gfar5lS0hjZ9k+lCvPYS6cWjV8az
3+JeTGJCpGBHKMTnZ8XbNqfwjEzPStRGrQ2/Gr24eKqnWvEeBjcda/eH7XpsYTeC
`protect end_protected
