--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
actPGY2JkxIKVKIcPDLMmMXFyGbH9gHo6XEO6qaRXVltRHPwrXFD5eRXtpnFpDk0LCuMBnBtrqV+
lLomG7PRO37JqJW6mf0C4xOeXPRRh0cwVoQZZjc8CM1qpP/ASCqGqiqFnT2V623AwHrS74iRI0c+
rgHJegDepxeXEamCtpHj6kJRjEC46P6NrMZ3oWsr5+W4edaTae+GEtMto/MdAbyclgjWnKxutONf
pQpNM5MLej6tcnYALh/IYQWSPsDtGOzx4mN8wMbInfpNBo0MPyzKj5u6EariqqZROAhfLAqRfxcn
gOczP2bodOz6RbSml25iL3YdgOmES7YnKx/f5g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="mh5z9O0OXGE96dGzVCZV4CSHt1QNY+GCZbx7cU85syc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
e207wu1zcPI8x8BQXaiSmEUP63DdshF+/Qs+vR+miVapNqqS/NQ/cT5LKIR3zAWHG5UNqFB2cEf0
zuSljU7xwlCgvQajTmoOcZKkxtu8pQU8pJ3mTksp44KEwGL5mM51Nf0QPKRWgCBeiPY/lgzMq72K
Ea0ftHUu9cRWXuiecYAkjJu1+/lizkM5MeA9SRrxBRm8n++uBJp2k3GxGiKuZhWhs9Nc1wARgYPT
dVwyaLavlAkQDziZV4ybsWhh4QpamDvwAdHFhE/WZ9Q+AvlAx/yc/h7z/X2J3Z6qmRvtTCvDzoI6
k6cTgH1oq0h/aq45mjny5oOZbLjNf8rq7gOywg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Mc292dZXqdZ+ofKiyOGp2qX8Qq3lIos7s2vRYe4KwMs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13888)
`protect data_block
Mktho+/m4lw9XRVicYdkVi6TUP59kZEJF8tMTTSQCr1lt7ePuhLr07ewDkROKrwU1IX7FFqp65Va
DNFvWftd9yfPj5Vq24qIcAdD4NvmLUgkvE0sWLgXlYX+GYhjoFuwWcTrQf1dHzaFrqq+hyQaTZjf
aU1gmYaB0mA9xOWlSusVfYVVOwetLalchVL0xkorWYKAa8+/eV478cbXHnyCQX53KT7hteEHyTWI
ovUZ6FmRAnvmK5xHsaiJoDfvSRRmv0Q535W5LbC4Jah0iJS0nJUc/SUqVssOUraj1JRFD+IqIS6k
jxCdkqYTeWkAJyMj25z3YV7646gPY0MdCdi3sF+FAWQRlJmxmoK0EPhYltOfHyMhi9DJVAGNLw/4
nn/pKbzHg9+SHpI54SNc5bV6aZ/wyUfydkqgKXMyv7/nfDCjXjswK0hNdbVAEc0nG/n5NX3BFw3y
kuIsTvl3ZT3lKdkxi0D+XrEDmAHbQXbDdzFqxf6fDLKKL2C6tBLyQhc/PbIG43AQIC+0qysER8v5
o4CulGeHdgyGx2qPk1tCf0Z3WHHYKl1XFbd1jS674erwkkGqZSVguCBO9iI7kDr3Q4F9KOR7lomX
fMktnpj4F4fmYP8HSfASZmYU3yqb/ArKihbJmPiFNa+V1Fy8fVzRrkeGO/Y32hHCbP2sIQfru2j5
NLdcZz/TBNGeWz/DcCO3WLUA5q0rJgJlwv2mEFUyKkxcW4HvZvdfTRJAGkp1k6LisSuMou2TxJBX
Otw+/uDhKJ08bVJGrvFQkS6AzAD2/N0DHO4l4sxweQF+8356gJ0Z45R9olo81CKM2PiBqZgvJs+8
L1h95NBxdv23r492nG/6+Jxusr8fPqFoP+0d2+FSJoCDIXI/CtuN7uhtv+rtgdXOJGaFHtPWOU7z
P8WkG5RTl0fUMiN/wTQTEZz/pYZod7feowwcgkOP0t076c5bq/7LZFJ3naqx4boSIqsCijlHJw7g
SD89BiXvS4qweeY/Zy9qcXmKbyOqSiYgl8tlMq93CkU4lnqxYGMCc7CpISjnQhg3IrihTvD7jL+b
I36EH8BGf4Kgj7/aocwsdZA42nHuYRgjjyKu6FTfi1kvGN64+I4yulaC0gKF235E6prOdRhCo/jj
/qxHSPx0sK5vze6YmIdbLdWWbJCDGaqGjqFdocwqPikBCtcp9eV4pDDhVKPsFdBiFoFp3nG+VNrU
YKkitmV0IE0DquBPeqUM55NmPn5KXdYWWLU6sesTHXmNlDSHaUX4JASmO0sI+7qMfuspaNG3sMCO
BBytjnMn7R7x6JDRXP0ZPQbNq7HlXs/6tJRfKc+MGUt/MCtkbKlSt9JvpoO7A/wp0L0/Qi08pfDJ
LZYKGIH7DZq+P/J32BSxFrg2UORXXlGHAkKzxDPh0T8MoZQnfJUEC+oG8HbEeDGmMy3C1XusJh4j
krgBM0rBis6HKrElyU/49XSSXSlO3KLBfqhxKokEFIBlgfUny2oNXfu/GBjPj0vOQfqHYjt/RPp6
D1SG2gKSOT1MdiikXdGMOxChcjPsyzSOAomoVeOpW77t7PBVfPcfDA69M6HGgtRVJI8UT+yX/0bF
klNf25OjSAAdC/QNSDGU+9H9M8PQjcYza1QY9ONNApP/MkTnaVXEhw7BqrkUyqBS1Nr+iRc0w2fw
oBXvxtUtxBJk+fw/eMnlW0TmDDrIxPpPswXM4+2XJXHD6YnEqs4lsB+y/4/jbcOck6ZByxgt1isG
skQPWDf2vC17W/XMg/aHoLLZEysMJ6mZgrglsKJ48R2hDaGXgeRMIVsNZaaLWOYTznM0IyRJoQQ1
QRhW8re/ZLhEvMXbvCrthdny8KvtTWmhpdbk01EZjtkymKO+GmpI3ux675TSAi5Cqj6OdyZjmaJC
iVlRmZdADRAecnswcaW7+sDRMnSJKmitXFjo2R1VY7ERt9uDtY3CMXWce7dYxxjV2ZCRvafSLv2G
urE6lT4Ep4EeskpZxlY/+b9TSnPHSf2+l0Mc0ba3+aTSZJc6oNYOslT+gypKRW3rsFFYUReGylDZ
PVzMRkV3jmGjHvwFBESuKly756NOajVp0RHRZm/F/VWF4E2ZDMqEdAastZQHM4CG5XwHZOy4nwaX
ddySFfYncb8knXZwDCjTkPsGDU3Va0rIo+29KhZoHdgMEdsz2nS9y7xAgLqq7OnOaeJ3l/IyKWPg
1OwNYMHdzqCFA7D7lLhNayxxlLPfJuQ1jIJMA2iLoU406X+92Ahfkf920NaLTtnGaE70/SpjveI0
jwYZDFPDem0hKDCZHgbi/qT/cc+ejg5hjdhRC0cgcBqJTqQfmjX6uyGpJgpLlH5jxy1oClrvmmsb
qa2oKR5bBs7of16Q1t/QLV1Ihv8RhLZe5n5y9gb/eAsmj19MuUSH+TMy21JxKDBIky3uF4gCX/5y
blmvbLNB4dthUM2IqOBbyum2ZZ4tSCL6OmwbbyDu955gU0qDLn7ebLNABREDVMBpH1SyLRarYDek
cQFVC4tHI71kaV9SpBwpUsX+vyga5EvIpq4k1hv+Mvny6kLdfP6CPwX+lb2s2XqRwLWSRZhcN5B4
gXdYxWSpdMl1l1qXMnStjktBCRWvs9mo/0Jf1ZwhR8voRcJAVE5T7fOWeXL5b3dWReEZ+eStzeVD
A7u3FxFkTtj/9flYdXII5k83CthGSZXzEnwI3U9USWmYY6p8ONwPsFIUq5l3j6m8rGZ8qGiRGXXn
2JxFXE/cu5/IncNS4+FdRq5xXo619sjZE7tuGQC09bYL4COPO9Td9VHbac64lHF/Qx0aPbpqY0gd
VNtOfH+thRh63/elADhNM5XvUJdB/pLeuSCEPvW2xth6XpgbvOlZAZAGzdrmmcIT0RqV5VU12+Yg
UJ3zLibrPkbMcLBOyUNMM4yXGNMSI+4wHPKktfSw9ER0BzN2VY2crBM3EqvBxWCf01lQ9wQO73dZ
XSAlNlq0LEPmasz16ZsYTninOd0jAymRiS2TD4+NB/UMC6NlKimBRazzHv1afJT7acU2RSWOwZu/
2GgoraUn/ub/qa1BX888DOuzpeQgh6FV/YgwQH9RX+mPyAkCBbawvQHoadBU1fPdH8lbN2zTT22F
4k8PNFrYOVFg3o4DSk1gE5B9EULsnUnNCmDS5qkUgK+qNQPZlaXHphyPRQuhWT3aojFmRHHNhKZ1
04dRcQ4OjUaX05pDC+RTMjw0KLQS59rtQypRRFD/iwZkxXMtjXZI4etQChS+cZiP9jJEp0Ph0YJ9
qCGfelncYdK+Hcfk1z9ZYXbbpiB9Vj5Lt7kHAu/HMDZ/0NNWvnbdTlG/LANUFVuWrgO4ur021ox0
qUnBpCeqzQ/ChG/vNtZJUKFWWZi9jaGUrmiZ0xi2njV3fRltwLPqFTORVqIlH39LwPqMfYLD0F2u
A8HEt3onzT23nivHp858+8CIzr3W+5YQnwFZQfOWv/G8Dr8JSIO9fkwMN4atBbX4xos3e3c3vnvc
O0iYSZRzH6cNdSap7J8xyzp/HZUwoPEZIUSLVGHrEAU8xlSzyT/BPkKoQCAFn848R+ypnUg2yLMp
lx+cTznk+rFMY/4+FTIQBZUsEmjKy+m0UbnicZwdqvc2o5zC/hbsUGXveP2BBLFePDUtH3FA6DaS
RGMGNrZLwq/+RYrKh+Zssv2zAUInoLE595U9Fh6xc+6PLPclBtVOp+HjRW/SrLwA3iet8CVxY9lF
BO6FiyRuJflsugpfUaM9oBwSYJnxT8XovJbg+ib6veszOGTuoGfnKdv05OO0Bx3GWUbf0mQsAgCc
WSnFdBCwtDgDbn+5+ZdIdhcjirD3jsfYl6qSWcNyzfR57y+a2pZbh4HD72v6bJX9n3gpTrOeMbwQ
feSz5h0YdXWj9MEH0gPNsLEN8fYsRH4Nm4FFuBVmZwQanZPMTz845t6bbuTb4vpxRNA3R5xYsm0Y
LpHNmXEidBWsYcWzpLQpMZHlEBrSZXDx4TcBS88yV6wS0y5B+oirCwSl4HLUQyu+oWNkxY2YGXf0
EV7FPpWPV2pZ8enY2ueSt4TvGsA/0tSdWQyhnCpKUa7cTByfUI0MLCZSduELMiGwoxFMSUR0UKsu
1Bt7LTJTEwwZNJ4g0SXRbxI+eJVKN7Zn/PwY9jSaGt+FM/w4GpDp43N508b1KKAm00RMG54tlI4R
AJwgA4hRMcW7F5lwxlCda7Lcmf8nO+F7SNtws6Zxvaf5OWrF5RFKtilT6TsoxqjWNhumtlYHB1bl
YsYaNLXwUnhMhzZI5AeBUH5J24gEoNriYXNAuaY3grlOrCKcBZH6rTzilX66d+pCcBySEoy6WEVQ
8NaGZWqUlaOnVbjvQkU5XoMYxqTaYTVATFTW1D9TVzF4tSFN1N0uW7ck0da96SlsIJa+7gS0Ztto
cQoIEZdbSAMvGioBJfJXNlMPeFoIIXtmPfnZlo5sFc9moDFAg5v1SbTC4NXH8E3Koo+dlRmmWs+X
Yp3Mjm3yE1cmQBUCVp3oj1McRPPSWmxJX6a/fQugCMUYfjhD2A/LocmA2ckhiWH+t5kZDEIAmLoT
+SC5/9dY+Xq4n7xAz5/yQg3j7iaLN773blOtPXBXNPNS7vmb/JfO8I50ivH89sXCCreK63W1H174
VXLIYy9WYvJVdBMYX/tSYeXTmIK5P+35zPD2GVfIQvz+ry1cN+jVwGG/6M1ArQquU2HV18XJq02h
B5kUc8eTPBjTxo3cjxS1w4dGfafgMHiwfkeszqmU+IEHbeDcqM6pIkmEOLVu8hO2h4ZPO8X3LWTh
PmN2XItkTtEZMHfKTLF4YCNAsG3Iv8W0HdnmbEzVGwqFoH2zpIBg4q6fVt/4fZU9JkWOUUx/M8D4
ifUw7HiFRR+MXL+tgX1oc5ph9db7kQaxrtMyjYEgRtegA/qD6jCRIMxOpYNkZbxz2+B+XmM/VLoP
vc47HzfQboTWsmOE4ivs7rKyXvVU9tTZxtD8ajgWtNd0NpuFSqzlDS+Kxcenx/8bpZXss7XnH2Mz
iGEY/5wphOmrNgHK2Ew2G+1LX+dWNOMTVeert+70u9Tf0t1XDwIDTJ6l7HQ50uSLt2nV9xZQ1R+w
3fJ/S56ox61O3i/mfQCueIvLD5l0iA23uoJ57uYyRvWq+cYagysv52rTporYC21aMNyo2jeQaB0B
A1GwmnjxKFB6zbmiuQ2OQM0w2zJH4sUPCJLwF9wI/tuQheATVwBpkn16fCAW20XDs0kikDf2xkkh
gD7RFvjU6xbu8wa6I/qblNYHuPeD84Turzhliupqd659wgKiShSrbwkTPLpZG8LbqjfCWcwo8on1
kBB/X8oJy/HMisfmeOf33AR8urllWtgIXCR3vmSfD9PV1m8iPXpeZBDDM/R/7UwjAMgzcXFcrfEV
ITOTJM9zIUway/1KdU9wMVlWyaWOxMBL7bOeQmA1tzAacZl5cBDTNv0a2SbMAz1zcFpRMFaaCTpW
vuw6O9PIaTWHQAwoLpdF/FpMlTMndM/lDFtF4/oci2b65EVhz8IgwxC41hpj2BhAhN6nY1dreeSI
zgpkpVg4IS4wF5EbDPKzNlTEQ+yI8ZTrpbQX6PKl4/a3WOjZJ2KLLa1H2vXNr7PKQM5BnQQLuf2s
Ps60bLdNBA4KV+8DmHZlI3+oqzkjJsK0/PvLfaTExSUgszW/b/X2Hsg5IAbEona8NWzHdp5xWepw
1v7O+593gfFEtQ8C6189RLHP7jgOZhKsx2kXpa0HOQMq4+4mIbXWvv3DXuuRD67WzSo+3BhsrIsn
4yCPx1yD5kulKf1ojX0M2Ky9GveGuG/lbZq89CIi+OR3FUhROZdXSM5g2ORU5UmOzqczlccmYwM2
rwP2x9KdmWoqr2k8e7ePK0xmMV1TjpLc4lTyi319TOUWcqZIne/j/N1BfyR5RInzZF8q0Yx8kQLM
OP1rDD7TutTsx24rxC+QNawbCxE90Av0/XcewSiiCbCF9F/OK4jAiumJhOaDaPp5kzoexijHW+H1
GnPbDXEJA9QlwLU9kcaWkG8spQ/y8lMYxfDfbq1MBWG6fjyMP47N8bfvU0Hes0RJxEnH/cZIn95t
XmoIulCGdPIgMDILTOuCQOCSmsB03PaBqRRNDJi95Hk27tDdKqLbeG6uaozVr04FMxYzuUf5UNkO
5JFwEUSIauwSNOH5+EWsYC84BaURu0lBJBK46gGh2LUdERqC7l9hkQigeGfO2OJdPQO644wWKIQ/
S6YtzwhJUDdTeJfG0iycCwkyWZDjIK0SfLvpFQLtPS7lohSCBoIv3xbeQKn6x6jRg48mEDFD+Xl4
97eCVYfEWKzoakt6YOLc3KWJg4uWQPbsqU9bjHrAv2v3d68rM5qBLaJkCWd+bvZMvQEcvIhvyQu/
CS2LAR2rkJnzkPYB23RBQsxXbJGdryIueSBCXMks03X/mzrwJ5pn/f6/zXoJYmHeh+zPtSkGO9XY
cMpcfdINXno0SAeDdXdEQVsoTA+uM7pULegKPWAAgYl2XpfjzYAoF6wbMKsAzQon5UpTJBH9twm9
T97ieNkcLBJH56uAS41b8pq4PbtrQxSxN8oHj/y512ucYtCOHHxRdTkgZYD/4E0KzVzy9K4x2772
Ltdwnv4fO5EwoyJp7xt8YGOCJj8LLKyfZlOp0FYWUtgtexkgzZ2LWucwO1sv721d911U/yvxM9Ew
oBHYmNIsCnQRc6oHsn5FtZ1A4DbGTy1r264wzE00D1biqWUPivRHaWkh8cT0Z8UXf2FWNS7c+1uA
Xg9F+QKEkCmkntJs1Cx9GCJg93oNSf6+0tPd5MD6LvuCoeGkezU8lWZ83ixiC8v1I/oRgrLOjLli
Vb2tCKcZE5sn7/WaCKRjLAcvAXfgH908RtXHzrBhrmsuXQG98zC4mA18BsYJ72B5rwpxhvuUop3w
9a1lYo0AZTojrFq3fJuYVM1epjE2bx9anyIhLrA2CftuX3jW1hAuSwThEwWP2uO0Gs3r82CeZWEn
adVpQWdQA7ukQpC7pZWpis4BOwDfVNQ8b9xr6NMpCDWkYnSWtMYJbNIbNuvFa6LGXLnnSHJ06WjY
yzVDxXEqWOmGTwEu49PXq0zmWVyG6KmfBsEZ8ZxhUbTIcZ/+K/m35hhYNNYxOQVlXWyULMUkG2Vp
vXhdH19Hz46xfd2ZpsByd6nGlyJc5owG8JxT1ShJEP2D9/BudVfjsTM0IxBWEvGAkvh11ZvPIVVM
bE/iR3SRie02HkjbQRB7kCdldaX97hn8GT5phGwt5vT9oSb+RM54XKMqWlCWHdK9jiGUlNTFq2U0
x5OvAs+cVvsXqiaSnu16BzzqBjZ4P0gQ56eccWbjMhlR+5FlFEKRqKtG0YO0+Qp8dBoXtNBRtaG0
UYytXKRX35oHxLPPTGcEBVRBvi9LkjA+4x7mghkpKgQUrqkzVDZTd5wieLqVcxp/PttVXBA/iDDD
7OP61SILIkDgOfimAXs4uFnk9PCEPRvN2LkWEPbUBw203h7rGz0Ui7/uHuvotsCO/970rSfd/TJS
Dc6AGFTybwUiTWPVoSMeZ7n9mU6dFzshkTMhTDDQc2ZTMdlyhlvjyWLEB59Of+5sjCnYhXjIRPuK
n3K9c3UcFKAJRadWlBlIxCtUbPYS20fJr/+FWIuoBS6Zm19OOdDk1kyoduJFOAy8Zvk5ifHLi4MF
LqAe46V+tdLnAEBGS6g77LL9d45VwM8WYn7JmlTAbiEySbz3RwCgOa0xfHeFu2+CjdJvIWBdLJcN
Wo+flbcv/EAP3Obj+DCFG1cSATNL86BsYV+4HPqJo5vb7pgoLZxuXL78Fb6Kiuaw/RHttVGsjnOv
fTw3H/LTjg63HsKFe5HoHVSBcCZ9xzy9oILNvnvZxWbk/JfRyK7lxQ+SnfOaT9GxNQE+WmsCN2LI
2rvo6ecGq27RJmqlNJTuNfBPUjOF36zdtD3VOKVTq9lfyH4E6tSVM3lsLfLwAH7hPHugiQj1cR5e
PiYGBo2TDQjjXJ+/qZQZbhw3O7Ja4i081FazvlM3YWJotIq3rEJV/ZU5uQX94UqK6hQspL7Je74R
xaiSdHQTMBTm88QqENUj89ezHisK7Ecb1+7vN8jIO/keZhBXuaLz7+pU2LKFGFAgCamAnK3nJAjh
8a+4Y94u7qUHwiVlXChtquRBgL4bbzPqqgI986Q6IZtALrTBrZBv02e8Nml2x9oEkQ2ftqpJ1oB/
e/NjyKh0AmvKgurVxlkVpVp0/Uj3BonEpZiC3VWCcXjbh5DU8U0iRQNEhgPKEyCwYq7VFMtH+ksY
hRg7ZF8JI7Hnnm58mFrVeo7/OFaOv9NlbNxk9h+mNlKHxC3B2ndDRy2Xlxf3NKKRTKxVKrjf+f1g
yKmUqnWnut6QVszyL8FhflSRmOEDgcKBYVpfi4tJOkw/E9OaxABL/a51HEop7OYhjRkk9touZh4H
Gto4pbv8c89SSvg293SNoQ8gSsD8w0VQo4qOGXaC9j1YmGCwOhoQdwP8TYs7noZU83IrB+W2oLin
V+OhGb79RDp8X5pMlb8Myq95xxl890z4h5BG9HXeXkHQ4PQ02YmZ78Ch6uSTPWhTZ2dhHpo6Fzh4
Mrswp1bm0KMln/rwXNoux9/xNKQyZB1y+yAIRdysB3OWMv9GP/bwlOcgkpRXHMizBaGaJQFc/Uan
19SQIfG3yv7MHOKkCciEQ0NxLIXYI5/WlHmFCX2PbFPmBEWXbgzToYPx+uFoDlbeLwYjK1w3zAcR
a4559sbp9hZno/UtW4lDSKHxWnbuI1mTeQhauXwR0apv8u3v0Xj3t1PDz5pvyUriVV1IreAxBS5D
vC6B+o2NACFnHvaXfejw2zp1mCwwAXJhdzHAor3cT6eqQLd2T7QHJMdW/WBnZv6CNkRjoaLZe+o0
VttDhD7+Q9Gsi+KdYU6eVQl3FUFRjOBUk5DgzK/QHcf2YJcm7iBalTNuG9mCVo6UB7jyXHnIRba7
dGCvSTQ2kZvGlk5gk0BUFCTEs5ygJrgFs/GUEMzi7PSGtXr6vAATg9VWRmBRv7AVRZI4UP52Q6xM
z7qK1SEP5xDb9mppRQTf9y/1aSn5yKafVWgSQTJjy282AEHND1qPHD3k3YpfT+9eJIz44aprKpAS
0yQO5uKwD8gYjE9IXfmH9RTwAgZUJ6b9S0HURo9OnpFvUCQA/FZqOe48xRMflLcRmWjNhTwYCEmb
I6p0r0N4BeKr+UEMZm7SOA/Ouo0gWP8QsUvb+2FDHYGiy3mjsc1tqQVEd9HniRTN79TpfKvojOeY
rqbuo53y+SnDM68LSn/db8oHbAvME8NhhZvorLbdGhV/KwwSLmllJBY8bw2b/dMgIEJ3HCRrxBtB
R3uVOAAp2JefNK61RzbO1er7fydFrKQeGdz8lrP+4i+9s2o3gBjX0a8y8yKizWYMbtEkMbI66QA8
3fzsy2qoiOayCPRsypvpemASpKXU7+0PJbNVy5wWjYMlIlgEpxBJpM2+YJJJ5AJgEDgKGM3RBeKK
cbp3mpgrlJUWXOZcbczd1GVDT4lbMnawT65FB/+IyW/cE71RZxYPDHNJVc6n+kN5v+IpxrmW33Fr
DD7YqRXt6+uztVuH7wjS8iAzIodIHeS2RzEUWQ+bRlgQeeshpjN9sh/Yk3T+B4QOzmPc5ohv9Ox3
vGmjS3f23dwVfcvr1X4kdHagOKuVxIkpQn3XxB+5XCxACWwG/onWvyh2Udyhm0RZ8PCUiDnrn+61
k4se08HngWqOP21On0wkrLq6nR23PkQGNIf2ydbyL2yeL3hY89Z8RQ0c772UmKmeItcYuzKWJpyc
5strrgKUJLxkYzz1WHmxTiqehAYSDkfcK0pyidXuaaq45Y3DNgf95RjqV7wLaiZ5T5fGaeSKQEqj
nnLgePEE/V09nf1uVYBH6hK6dv0+PrI0brLLEoASTuRV+Iz5hJK2uziNIQBkV+hV6KPVBQr7SuVc
T9LeHxRxv8oyCFyFV3LbGLD8y7yk3gDUuIbtsat9qcFMcLN8M0cT/dZAZJAvA1tfZ6IfD1utSl+t
aE6GmiNtc5mWfl4+/b3tT9I80v/4/ZVEvZRh2pvEXtATrX8LjtYbcVrQ+0cATyCD65hVDIgKTtB6
GuIMd/NZO+OPonSsa13MjvvntOakml1sh7zvWrxmSR2l4wSRhV7SE8XCjtMj5zHkt15TD1UGTb7i
KBsPBOjRc/zDnmW92VyCocZmjfKzyPX6flE9rlGLOssKTI7G9Uzaf2KhaUHAlSrZ9mrhUiMCIhkp
igwg4gAPbKVCaJafMW7jcRk7LoxenXYbi4SwG0YJGIAGS2QRC/EsTNDrs4LY1NhH1MmMGTlaJtzh
WOuynD5sIhKdm9sii+6HKqJjr/kVXbV7Jj3Gf9MNByHAeaWSI+DBiTfwGmmvTQMj8HN0Q4Gg8oE7
WeE462iM+I/mNoqspOXjrld4fSEHc8uu7/8x25pPRkOt4DMNTqyf3urmylkfcxlNcCkJQQRTjg68
Yh078R7C5g+Jqly2UxGkkqpQ5zADqNCPaZ+eLKXeMJZFbvrulDyTWw15zd2fDIRtvjvFeitYSIc3
no9BrFRmptwRfP51mKadAhCQqqwycdD9BuMbpZKzCYUvnUTjbRDt/tMiTSL9o1GaLF8+RzLnfOfB
mHWU9PhOemCq7X4DGkDq9/z16e4I7oz8eEZ2iw0D0ffD5jA49BC1ykdA7etiTn1NdDlKfcX1tfLT
B4+IZtrUjy2vNlOHNlcm0c58/GCQ7B8MpGVb779774BP+g1lhNSApbyOz3xUfPKHtDeSzpP+4Wxr
XUxDTZNH5WUbHMj7I0tJCaVwJ5srYCG1qXVQV91OUinH5EudAAly3PSYeKtVscx9LyQ5scusgcR2
XgrVjblbfVVisIMMfciVqgeezu099V/vL1b2Qarg8AXJLj5bBEkXZId5rFvPVtY74Dv+FZDjZ/Sj
07b+if4zGF69CnCC6/Be9vXH5TT2hlgp28WD+YFV6xCkXiNBE401OKcr3V/nupm1bUQpr1wps34X
paq/pK1rja2WgrQQqff7BRW3i3OZ70VaBp0Jg5BOpzWzigAtLjgF0pO1+Lvhxxurt82KbzNw0k11
w2VNOpCHLAiDYuWCG+wqR9ZJHS3sVFJVO1a7Gduc1BzTKPntbzV8b5a8TCs9Xmd9G8syFvvS7cKm
p7F57AhLGmcaLfYRJvsLcdCpwUB96QzbXaOnRcuMmd3MjKT33GlIuPIfBBgA+PzmCHEEHG2dyzd0
Xe6nGu7zNHCpSjY7FFD6drTGRgj7Qk7kmgrhusgIEHryIMRrY7Pb95Hb3UaBmu8o87FvtVeriVAG
OIavU/FVRgqLqY649FS0k/3GOG5pkIFvhQ2kYD6cpZjjDMJjREwyoxW7bGZpqM/mr+gnkGcstvOU
/qSXt9JVGUo4LFGZvrgBQmL+u+qzIGYtZBBCd3N8OGSDmpTCCTDjEe0pASV0mpZb6EaRYrGKqfFh
74tAlvPRGerfQtxjU0jnYIkKAjqFfWOPd4gsSdWgeB5xUCWinaeouRoR9de3VHEpeUV+fVOJ3ogd
tt0QSrQyXf5JhaNPiKDTYjV8A9Zy/PZU5wJkZSyUMniiybryE+xAAoryXqJi2cxvXt/819sv9hot
U23G5YwdcwPnYbekkwU6hMJxWf/yO0tJZGmX0oDU/N2CENtw6fLIW3A/A7Ui75v6eOWD+A1cfeS8
ANIuuq7X1+O7Rdrd3ystmE8PGmhS8Lw6AVtXjTxPU06TZKs7WH4KJDUrtapWK2AKboKTY22gSase
i7891rP6PTJZ+YBG1Aaa+5HywG9rveFtdH3q6rK5gIsODFaNmrDLike+Hu+pFLbjsWhfvQvjDLp1
4r1sBxJeRsSOhLTr9VnC+DtYZDtcbENX5uqBhK1DwSGbTb2FLbyNdZeyrr9tkSGEeFtHBgGN3kGf
O1ISPVjVXXGVNmXcLKAXchqQ3lovhwn0+3IGcZHGXMDEeCznTe6mwZpeNusnrVcg5N4U4UlUu5Rf
hL31E8EMPBcz0UKmnX9oGg13baIjnVHnRo7MkAp1Rk40JBjdZ5AaytbNt6udpbwTwTwqChffJ2P8
Eo6IZTHkXoazLy0knEF/JQzd0vRdP8UmFcav7zVQr+wF5I44H0+yW00Li6xg2tkbUfYJBAVru9mj
ki9T7anFlfCyp57dN4GJyYBG4db6HpC+V1fxbLoxi89ecB0aBQTx8xEDClDZJHxJwh2nkyhu/MSE
Wa5r73XmRhhqcMftSkDj0Ichx1BKxSfqbPW7ErlFw3kNTs4mByv6nFMlDyBeC3SQIZhWJzVplAaJ
Z4seWoxbr8Nxy+4/FEL0y2FMIAvz/pe4Hayu0uMWmNq+Wq1gth5iQU0OfPdHpqcEBAVCJkSI2dgw
0sPLpG8KAF+8CpdVkYnHSsubCdQSBduu/w9bnzPz7YuZMhuVeNX5vnYoY5UKI9O65DVdaOy3uL/e
600juuZtei6eVVXFotaYzsEw2Yd52BFmJ1YlyKBoRue1NHg7ztnpNHyw4zJhNLFXG+uRs+L21/oV
5UTB6kH/vm1p4oSD3glqkjcXuLoSN8s1YPDLLijxetNHl9viWEiSAP60iout38abNL1AQO287nUq
h3tFX/SjhaQWfKUjNGhhqNjt3WOOLh3Nol3OpUjDBeiXk8kjtCQNjmmkS1O4D10//mYmSBTBWaA8
rtdSYt0grO5FJUls1OkK9g9GNkAtYkdIw9izxbtduB6xBhDwzc/wuUOBlpnuPQgO08SvPhXb5y+3
MN+6c/cxs24O6qBoYe5wNR27SQtfpNlKzQ9hCcuRhD2XxLMnCPmccHTqQZW3dshiIK8bL8ARDIFU
B9qZ+KNzgTaG89XpHoBZWyYUvd5WxjDNfNXhYrKl0Iv48DXxl4HLdMZjVvdUf3rpgKeyHu7Hc4fg
6jYH8dlTmS6K/4QijG8/0vUZG6jrFDXGGAj3xveW3/VjHGHQfPhSlWgJ5Pxa1LxC30Jj6y+ClsyJ
2a32dQvcW5XqyAb3TQ2O91zsIDcM4LMLu0le0/JrbAawMsCjBTTfRw6gs2wTv3fe4nSQWMGxAphX
ZvkbTObKmm90eTGK+zKKryOujN6ihVOoI2f5/HUsuJv7tttk2XvIiBo+ji9H8IsrDLMl07pK2DsI
z89mKQxp24+UnLep3U8Lql3arfmyrxt2t8WKCGtJLoJzORiSDJSvjEacpxExgsrU08DCXEhyfYFz
QWv0kTLozOkMpAfVf0jOVKlJUA6+cfTsG0TBHbgShfFwm9dm9V6e+zcj3cuQyI/GllW1mCWgKeoF
FsJA69oul+VtqDSoqg8hi0+mIaNST/8EMitx6NONb3YpptdGDrUMNq8ntTGuB48qGoyPE0QHO45d
T/9jwA/wgXjXE5I3dj+mjEYCa2h/cYEUWj8s2kMJw/CLoYtyZHHMQRgw4Yrowt3l3F3AnLd3lIEt
XL/r8sTnm6+2thz7kSQUau/PGhSawHfL73gHJvmkVI4hDe2wT2fjqsNc6LI9zUcOdT4+Fap8eKXm
AOcuvMgr7P7CeT/l1M88jifc4xEh7KmVoJ5ifa44OBOsaWoGif/qqjhskg3zUHk7N3RzlZ/rVxzb
R/gRB3Prh8+/MdgMGnusMnI1qFG/9zzWHE3/5YBJem7Ebqg92nsNqc/JYpQbZiRNp01EKbppcCLm
+ByYT1Eesf3r3qjlLEi5fK0UZbnLImV9rZVuKLze4YqUGoYbse3M+AUg7RiFnYyP4EP/xefZcqsO
qcVWnKsTLsDQY99TcVCQ7ZRN+e0sVNhHddaw6AEO0/GcNvaUl5Bxwli2D4Ae7vBzCTAz0q+IXnk7
rmbXM44rUx3/H9rEHuw9IefGOBqeYlVcYzxhRV32lJjDtsZRp9+xUB6CWT3GOAgPXRTBigRqXwa6
0vM4FT0lK6peqruInJwUOXvV1pOGx91xRUTenywfiCULnfokCj4f8c7jWQkPGvaCD6XFZnw2v28j
XGRFkkWIqQmz9HxCgi0I3xtkvrtrWntzsTbYE23zeo10CLXA/YmS/PB1fL//k3BWA2SQrq82WBy1
iEI6H8/TOlP+oheiboWav9yGhy3Cqm5jp++tgleTlQJt6+GAaV886WLnkgkykDgnnz+B5hJjJO6d
i8L37hDSjUd9fnheWmkosnY9XFyp93Wv6IatEojMpNzysBlmgtSQ2e6Q3P2P96CMuXEqR/1U+lN9
OKsQweRXZ6LznMlRygGInuiOKTR4wVlY3+OkHA0gKGxr09+ms+PfoFUUrQTZKRQLxqU/6OFKGFE0
RjGqtYS2uG4MZ0Q6ef6nBod2ihB3wo8uFBbzv65CzD80SjPwaClfvWsEMGGGogNBN8cneQSQMBBK
FoIhi1CvWGudlqejAk6vEHBgEOMe21Ji2u8OVZCllJeeW6ZrYEX5f82tAR2R2gFESdfhmBoX+jqb
J0IbbYXboFIRHefTdU0jj02PgP3ceVMAzz/TqVysfDvsZm0BTn9o/+8Oi9eS/JMQhZOg9/trwm2X
biJPyMopoGgQfFsySf7WF2/u/TY5UEz1m2iLPa3c25ZFjO5hFL8hYlXLRlTucDjuwwSMmi6OCz0i
Lyzhf+JMxzm6snH/woJhYA4B5+N0rd1PY2vcTmqFK0KgTSK0fF1jiLFdSx93KK1sMFzShl7Z1dlO
v6M52ZrYu3Ukjwg1d5uIN5qvjTT2qfBZXugYrPAdmrg4Pl+kFxwt1iEtayjZNfhj/Mqa4KsTyVkx
WfSgaOn0Jje/t4wLl61X09EniJTB7/AUgyd1ObkaOYiN8OSpXG34e0AQfk4Yz4rKleRfD9I8gWvL
cH6g/JTauqcFcJWjigKaNJsI6J8Pzzo1xb3agg9drgZn7XVYFgbk4nyTorrXZyNuyDVga+qAjZfo
WuAUJwCBrfXjrS6olnwHfst6greXkiOMhvtL3xJPrcON89NS4KI/gCWlPiHcioCR6uPrkJNrRyCT
V2iPXiwjcBT4+PsAt4Wdqr1Cc0hJqbQ2qpunsFkMlARSUWYYYcwUbqMWfbPvofvuE+ZBLyJQftf+
2mWOW/68O8rMnq4XSK6UsyJ7n+Uk8vwM3ElSYa45fj8NH11c+iVhPQ9apzxe2QUnYS1QW+Twt+Va
pIMeO+ncMIkstWdEZvVtZYRWqJlaV51ZWM+cvA5a+RgzudDlMMZeiHghTknn7f6cUbAguUfioaTx
gKrd2UCbvZJsZx9TfDFs/EM6F0hiyCHrd0STmmgAy1FSawNG8rXftAz0hhtvH5lWjOuuxd4P9lGU
oimQq/D/JHQUagvY9JgQXAOzKQr/MzOwSN8saymOCqaw/Y0aSvqGjKmzkZugO7UB4r8AV/25vRTW
fDu2PLyUmgA5ohQiYMlUCpQT8rTiPPTGw22Mb7seahg30ob6qSXd1DaOc9fBLTvj5emQH9FT0dPC
vPU2/mLRDjTPDqUtDLp52nMkMIKQjgDsirlPxjm3ymDuz28m7YAR+3xDom1XMivI5RIUCP3HZkut
8VPVmDmrdfZG7GsX9AWzsWz9d0NKd37g6rd7vnSXYi1y40X4z1bvUKGGsqay4wvrc4UPPKS3c2Ne
8RjY9sfbVHoL9oVxlDnTAAtuPuwoqVkOQo9FVHe9GkTsWIAo6dI99EUREmfRabKmIm98swIr/ztV
3ZBHvsDBO/uEUyxGB1m6o0iaUDSNp9m6C5He5QCEXRxeA1ZoSgl8uB8JWAshODUWsf4Bzbb1MtiI
aRQBDt7gorH1AfySaGXm19C82+3nUjTy+pSbki1b7RQp1xLmJPx4V/7FnCl1MnY+a8Aa6xYbcRbX
ZaAL+bkvh3oSawu2my1096C0cKr1vfKd+GEEAGQuSE4BTVdeIPHHTMweGo1tyQTnMz2gem6j3W0q
VT8MrYKJUf9bT29ucLSzbVATd3r2pMGtn8ILHV460uGlYHYG/KgQ1p4LrVAWa0qrti7u9jvxjK98
mYTvR6W5rCN0huofU33qxrJUuA6/AjvC2f9UT8/mFsdTl/s2urAeRLDBjjxH/RVqNSJFC23P2kHx
vHFPFXv953mLeGbwEqTiwvwu+wvx0qSgGM3ggl3Ao1dj5jDChVFsaplbQ7mxz6RTct9QAZQ26G6p
22/9AsHAm4dQQcBEfusGHCUTp7bRCtcSWEWlON4xR7cwnmzmoCFPP9A3PYv+tPATmxBHZ28SonXj
o0A5hqLoecRsdZtiurpPMUX2QBUoy6hoMdYTQlP40hj2Gsj9BvcEPxl3ZwNdUjbS3coDx7rJUzd8
L6Xo32F2RboFFwd4Bah+BmSDxtCt/7Vf9rdzWtqFWVQn0/eqIAAayc8P2UEL7AmKL9pVrYn2HpFs
awmlP5RE/elFeGwFllZNyOiB9YX+t8eXqlbgF90fCsfIpVTwDy8g0jlcYzUJ3u0WgLEnmtBl5SoX
ys7iY4pZSmKGfFWz+5uBUsg5DukfTLUKmx9e6Kg7pieW8tJbY4ztIR/jTsumRQYg9CqSOeiNpb9c
7dA8+W68/nEK0taB1LQje9vh3sOuqJw5FAJihm23yNd2Kc2CpkZE4/ewLq8Gvd8QNtNWLqKvoazr
T1AgC0yO/jk6vKwVC6DEsrUwRA6vbRKVyERPNBvSOzK7UbwWvcGtEQ9umzx40psJNv2W2nGpsbA6
xSR61Ec0WPUM5Ksi0+k5MUdr0D7dn6pCWgnS/DNGe9IisIPYAx3HHvQsHC6qPG/JPnJj9tJSy52F
oaQBflW2Tf7vszK3FD4+9aVWVcEfMms5Ha9kJab5i8Kp3BW76eOsZqgeK8rbwVjA9dp8wrsySMI2
pJ1/JDBptc0YY0vrw5iV3EEz6lmjDIYfenWxxcPeu+TUw9Jmil0Vc6WijWI/3Qs674FshKVmax9M
DuEAdFN6+Rqo/WX0m1rVfsPYYWaDHH/sMPCAH0PoleRpIUZjZjWWj2kA2MfCMf/2vSYxKofQgfVM
b4bb6aH1tVGz5Ly3cgiIZA5nh97d14v5W/kO+ZxqUx3ENyD489UpoaNN6O+36VtTuqSMZps1QL4Z
FjJJUSkWoWmnrGecrOQ4VSXXaMjXq2NKaLYJaiQLH3DxFo6YxjLxsLXXqOL9pqnSB4OdWzBAUi7X
0wYC8q61KGn9ULN+4Kx7WT+Jh4rUDWIFDa7tXCQcZkcnODIv7rvzQuhHu2r/q2ai3i3rCTZPIdxL
PEzbaO98kk9A1EUA4FRL57RlEA2q4njIyimCUaxH5davLW0JJXfKiMpUJ8qdDTF7URANbOwwo0R8
9Hj0saGoN+OrX2GHqZzCZJ3/g3HdqnW89Z9ZH6PFpqhMml0MgVYjsERYpZR9t/d8boFpmqpX47IW
ElSP8t1DXifUK5w9Hy8/8DTSbyxshbMvgy8wn3WFY2KWkJjUyrzqrtuJf8yCnzRwniNb3hRrnkMX
GJ8s171fSFZO2Fx+91mNY4FrfemMdHk+7qIiWmD3PpbUqtJIJmeh7CqwB6I7LGzLS/eMxGBfAzpO
qgiSSO+ZPnbA4adtkDtgGrjAXZXEoz9fNMznWrko5Onic4YocKmFd6JMHfJ/F3CEKlAOtKWkO4Vr
j5gYE0Ki0+vAoFw6PphBD4HOYUqOYyC5fu/adOA9JP2HuBczflNIptvHSM+cKWQ9iebpoAHSPOpP
wOImTSuhV0yzBdachOZBzj5dslrfHjDpjmVJ/FaMEQMC5T4tSp3fcpRrVftYSWJjEXHB0eQmrx8+
Wg6utoV9jfvs9Yku+w1aNnYpmsmch7GP9LoPKPgpyHbzo8K4oAA0WXsNDjzO1H21k8wV3g/s++1q
kNqllV6x1xnkD988+5+Frhd/YBnNNZ0W2yRE+aWXWHbtl/tUCWi4+gPSbt6BHDYZ+PdgsTueNa7z
GoNKdELFmgTbRYjuaiUIEK2fAEgnNNjGw6ADKd7z0W6VVdhPQMnTOfSjlBUmu2Yb0ntAznItYjNy
ag+iYFiQRdulbrQgLPwvCYNkMSuZZJH/Kj6hklW4L5ql/WqQcya9d6wh3Jp0PPEf/m6wSDsRji6k
Dr4wRzxKlPhGPXrmM5lmkvox0qD35fxCjL8OLcfmo2lHkWxcrdwdyOk4jcMhww/uE4wgax4oA/mu
hS+PNRGEAftfWaw+nvZVbkktGtLx2+iPInC+9XWbIeaw9B8cVyJyub+CGv/LnJHOkiOf6rHf1b/6
e8N0RTLefUsQ5qhmg7XWXYLXOKKkgxK0iXUT8ED78O5cM5aR7P6gFspVLlRbM1vAdn9FkrV+0Hw0
aGwgda21jCaoNfzMm7c9GK6fhIYjf8ZNzG5yXsL86tTpQ5pY/rXaIgxWa/zfM2RB6+omEiAhqcvO
Tu7uRdhzG683CAyhIav7iMQLTg0Zyf+rTJ9iMxqDg1V4KqthvkIJwRfSPTRJe3gSGVzHWnyFHo13
dDQpKupoXfj03bKAd9dHDDibNzUaFslafY/fDYBAI0YgT4RLp7vGyv+Y+2Hj5t3nMqtJ8NMHgF4h
MJ4kLzAP7spn/UBKS5DL7bNY7pEcsVp9NL4H1ysmYjK2iA+CDw==
`protect end_protected
