--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
N/kbSTgHKtK5Org88a4mJwUMvIjCH0OH9M7eA4BewzLCQgSqtsAgTIdPFTBK537L1TTMEirqjScI
5AYFKraynjJ4cXBZJrgOYfV/KFQ7CtGYsZhnqIYGssyMigUozoQQnX66myo79RK+fmWEmKpfTeL5
izBfKWmzE8vtsIF9z8Ow5rvqKkCxHgswxtVFMp9Ecw0hO4Z/0tQu48TRAklisnrLCtyoslwrgz3Q
DPfHUTzAO7DKbchU7rG01nWgRoGLkBUkxpIG+if3clMcBpigh9LR0drti0yuiSG4r4KLGoYud2B5
Aao8lbW2/04i71Q3loq3ShpTQVWli8R1V9ToPQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="GrSdw49vOCzI1wOheShYxJ3hYc3NaAYo4z9flEiVF4g="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
ijOO62p7MkyN/7aCt+l7+6KQ73jmqXk9vXgU9M6uvR7mjYgMZ0LC/0r/1p2XgTsqlvK+27k7iWcc
BG6DgU/TCUgVmTMrgXnZA5VuC/Xqb6FgxuqI4P2sAQsy003JU575YW0SUdCkBpvoWAG0Rs7G3nYh
ItSocKVm8NuzQlCAHOtHPZDlwGZyprVXcc5W1BA4NXwwrkRigkAdhvJAJdBA/EuEsD2wI5sGiz1R
fsvRntvl06yvAZPk3Z25EQdywQ3DDpN8HW/XYXnH5zgbgVm4nTkROO8Foz1PA/nSaOZD908r6fzo
mYcYMkb2HAl3CQBTyW/HbQMjO3SXRzZKeslkWQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="XNQivE/ppnUVR7cZgPLY3mSzTyA4H4jLk8dti/Usa3Q="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10384)
`protect data_block
wo4BTwKjBYaQ/dsL2EAuJRoccd/Vp1vcQorfUvGElgG0A+bKEMFNDYUe4T/Dlv3E5fIUtnvgPoKM
BkNf0721n5dj9jkboiZU2VzVblHcJgkW1CDI0klFJDhQShkmq6E4O46uWRSepSTNFm9RffzpBPzw
4Uupb8p06z+2iUUP/yPDBv/M3TPhQ+RL3G2eoLpq/aeooFmqRkIPOoJk8sBfULITUQHtakSxlnGY
GkFcliGoCEEdi9IXvNmAkIEKShJCqfjPqg7npX91yhb10EcFXKQpEqLrPBF07lqmkl+/+X+MVVsG
1Symtq3B+us8xTpAMzO617t7T8ol0AGt+rXJJ32MqIqIhVkbUlIh/lOEaIH8tBJjacLKIg3wJZn7
fc9Znc1xTblFNgbpJT8twuZfzN9CRQmGwpQ5HLblPqCTkr4emg02BnHL5s1LjkDbZL5ohc7/C70V
kWVq0GkOoPwwJqm20z9K2nm2NdZHOFx0saGD8Pmg0vgPcXVj+q2eFW/b1FoDws8iYkjzzlRlWn0V
h8TcG+3hqo18VXhCG2CVkV4ncEClh2aKoHK1T4FKZDcLc1o9Ix/MwUUrIrnVhHLXx0KEAWvjEgcW
78TGoIZE2GA9Esajoifc0s61cK9CbQoiV5btSNeBs7fD76XWcBSLmMlbxfOdfZ5kpc2jf+W4F8ZH
TXZhheS2a4UZWN3dALR13lmwylSUvrVSMFLGQnQ4EiKExCqMliW4mJe0QAQa2EjjFPrvOi9JMgDH
LW1qg2vo95FfC7BfaVdKsVw73+KtovjUoTeA70o03qDLHRV1xp9lpMoM0p9bV0eYeMyDhEEzGi+9
JiukB1mjHTUE6P6nikxvRoqKb1vaPdU4HD5dPpJcVTmxa47P0U6QwaXs9a9nhOgVGYjNXL7gd8WQ
L9rTA+hkcX1dK/X4yNyQwAHI4OKDTEdzWCW133a76Xh/PHp9tnjMce5O500vEZAKgilEI1WqxHgT
a6sOpDK8QG7qxFt7n/Imto+MQXMZx9IUA2r0Y1OIfJcj4I28fnPi0gEWc+g+RwhRn/D7dnqEIgu5
QYOnFCWH0HGAHF+TiQJWgk+oltTAarI+y5u5+GwG5IL0wiF5cABsrRmOKlYBfSZVyUfSvirN5bGS
Y/S8OB7GlQW1lPy0JO3g9vUG1L4e+1/ZmX33KWT7izvKHms2Pqr79N4aK3sEYMWJVPK5xZnZg8P+
DrpezfU7YZ0hWzcIZgrre2bEvyZzDopWtpjATe2vIhzgE0C62+cgSiyqhgBa/+u1BCys2ipMYEmf
Hm87SOHpb9/2hpvLCoiA9HtoX2KMGumUTIg9fN/7GtxXsp+4mao72JVZHsm6lFV2cxPL5WvUqaxe
ld0BxiGcgBeOkkxtXfX8C+qv+J5GmGhkb6N6M3sADyQqerDbIiCYPU8di8XKQAqP/CWee9nWNtr2
5fvfLLpwH6I9Mu3bChliitfkNKxlc3rBBFarsr24Dc4Tn6VHptlxjg0gNYrq2bQNZrF1poB8mL1J
pTye5+8ULsOxQs8M9HjzsV99rMMB6u/xtPrC5onN4LZ+mK2sdAZ/vONZmTVWWMMT+A9PDwFuMujK
+xoKseWFOtBpHrz1zRMV6s8G13dYpO1dQRojB/PbQDj1d7PUUDxaYcNg9ns5NISBRhvBHdR8CTwb
SW8O5o78BKcVkOrILi01XnmXBe7lrJsMDGuGM5uqQxPN/34VVWhdNyNgkWDXbjKXjhd80c07HzYY
pQ6zwkOBNtweG5TmSoKPwWgwg0aVANsoH2UUvQG85nxC5a9hvUwQPyJ6XpNx+Wr2bayMNejnn+Ge
rWDoPsRiTHEAG+D4eLdTIgkuHJt35uIygZXKnZYVcnS1R/uPk/h32E0FMELv02Qmu430zsv4MiTr
cJgXytTiOVJrgxX81HVPgr1vPYcVAvW89fThL2Sxj0K3cXuuDTiKOXZrMSs0ZfFuBoAX4RoPWwID
kZcafnNS8JH44H8zsJQs741L2uxRNF0K8U1N0kOs5pSj3auFCqOP5pAZ+UC2/mpi5EwINKlMgrrN
x1G2StZ9v9WlGKkNsi/5DzzkxEdYtXUkjx2q//7rczc2/yytmcar4J56p4iPwk78Xe6z43G89bXj
mUSkECN1at0bYdTrluziXZ1lusSlLDSfI0mHseDEWhyV9TIBH7b+V59g1EPZiyd6tr1Z9+K5zGEh
4d/lMuyHm8sIAH8dz/0OudRt3opT+E4jvGVeaGPKVizzmEIeN+gTU5QZJnNjW7DQ6L2pEI/6NRZ2
e1Pihh+Z9AYZd0t67WG6xVMyyV9SSyLpKNCw/CaDgJQAey2qBrXK0GrXgYcrgHoWKI0HswQK/tL1
J1nQBoOAFvOFvoltujOS659UKUBoFKmF+XcKP/R8bqyybHd5s4BkhCt7X6d5a0PcxiNrOQRQCQQ1
9cALKbr9H/Ky88+HftQoJ870UVcXTi6cz1PXQ5pwO8qy7HQ+puAaSOfDBwJIXqV4cb1yZcUIepgJ
sL6DzxfYCSyCgm5eHAhfUKCUEuxrFt8LzyvWY3BO7LlO9iABs9ysIzofG8tANYVylNUJgy0ExjkL
i0l7hP6sLM+cIfrpU1k9VvA6pZZo/dD0rYR8wTBHOai+qXxNk87be4ZoOh9oZWk1XYqmPyfKSF2P
wtl4JgatootyufaQLeHF+d13JwsVPbOdrVT24ZSV5mbHeagTgr9mmqfdvVToamgtRy4l43dLcD5N
e+hJWiGMlDHKYbIikeOp7OU8+1uLpqgrjp6B6xAZumNNXcnre9w6R/7evHLnvebwE4u8GsErIh1l
TE9p+074b7nk7W385fRL4zUtQ44u1OtTWWMOWrIjKVD1V0vSLgnFgmOZA4dAgbntlLomG9SfMGv2
hV/ioB/qpOtEHZW2rSDDYBUs4uNwSbJOqGJ7QRQcumHpGeyexQ0uQVfYt9JZWPpAqHjeS6/z9jj2
Cb1C1om9WL6Jk55gx/nlIsACOStBUh5M1sh+fRLZffOesdxuq9cF5tuQntUijDTLFoY1jaAOrxZu
XK6kbUzhAkJ9YAzOJjOoHMF07YAbIo3a67yQ1SOi+dokT5Ud+YEqkxN7XMgMu6xK/LmIH6Hw0soL
S7dHiB6RSK2El3oP0QzpkpypigVb1+DZaBHF/gdbQkZUQQCQXc80/qzRVpQ6Hd0+rb+GAQyviJXx
vAubwTqy3pBKQ65ZCNIBg73NQeyGUyvX+DMU1I8CBqHAj9FYDLXbqdRHnetB1qzebNn8c+IN6Ega
ugBkafJCh2NodRdYuPt4iKjpsnhodixXn26LH4da1GDwJXFKHysjyo+S5UB/n0mfAf+FuQwKeamW
kmnL25zSBy9o0GngSy5Pb1qg1P8bqiQXQdiOAcktQ8elNjCNNfMviTZbdjPzo1Zq23SRT5ezUB56
BdJzwtkwSGqedvPqcNXO7mbJBHPeU4FJ+9EzjcXGHWGrURnBfVj2hJAgFmi2M4hxWdzqYtRqjWUc
Oxqdws8zLxaLpYrtVjR9X6LxYkyJjTz0GiO/w9KOQ4WUtfDdy0TUKjsoyXzwewYLUgm6B5u2zVNu
rf25jESWHy+Hcs6KOXwRDh62Vd+4WTBhqFmz59BUHrJ+bQLHAWo8zmr88FooFobxnmTPEh8C9dvv
hx7YyDtIMpqdXFo389UhUX+1aDxi4yBCTdy1uFUkL1ZvsF+NXZqaiT1OoPHuEpmjGbfdPrgHuMH2
SuHmtbvyBb5S/Xp4m7Z8oSmGLkdhJtQj/RNqLpLVB4AlzLbIAsxl92SnJ0J9gdkAUmD4gy/wCKx1
PZ6D+zK9XgTSHcZTbwsiXGh/keYVKyuDqMWxuCvRGX9NYoL489sxIJwQu2aTGw3OREz2bQETMJgO
xwaJclRa/iED+yteLD2QTCgg721hEYHto4RZB4W7JFVVzedKRySZm/ti52MjWd5TcxtxoCX+cScd
RH0oAc74aiOCCnX0foWCejSQkRln5xNFU2/OyL9b969o1ZuZ/Np8YlTNMnxjQLQ5ZZGQeLRbY2E6
nXN4ZlJuvfmULCr5ruV1Y7UVpsuD1Thhs037h2iSKCam8zMFegd1mpVjlP00QxEhpzj/ltvlpdun
pAYlFrHMtyLS0C6PNxEaqUgXYai+DHdsFF5i5WM6ZNnHsaukk4C3Dvw9bMpePch7ygUCJHtNvOrB
ITbayRLH8t76xhKPsz9s77DZ9c9szdKETx8bEmh9Tyz64/+31djjLR8jifg0IvZJIo10jzea8bSb
CqqdSboaL5BrsTCC3O0Bj99yVxMnI6ljRip92reHjpkfpwUZCbS9eKbhTjlKnykcZUYp2GEUzbdg
Za2BK/xAZR6ncWJ1S/4Gp3pFdPvFrnS4sXnrwCYQjCSY2fh+Hw8z3NgdFPcySDP8MoUnpV4aFkVv
hpivE7AGI2UGCGe/gi4iTzimZJ9IF/1GgAxqbyDEjPXsMyipGoAz4vjNd3k21voeTN7W6m27xPTH
JFCcSUSQsgGX5oamh0+wEc7qYeYiGP2X5OBZFt9/oUdQf7j5OaqNQ4S5XWg2DHG49VdpL8C0J+V/
rVJ36tCAsyBwZzGRrUWDULLmM17AQ5BRd6rCEZ5evu9vGTHQlqaY85/a/x2vR9uyc4xDbEKtdphb
wd1lfrQAz8BI0iJWpd1P+jWF80pY1iBkJvxL/wwG7a7n89bUVGRuiyUeYw2x2A+hMbkkd8+HGKsI
6D+b1/RO/Duiih3lbBqaPh/W/RrCJ8DMIiV8pgjAWynmYsnVZF6sxFzpQC7lb4Dkh+aOER7ibiVW
+BY2VwEdzPNu4XNh3MRKJaaZoIAbXXAxWr08cAJ8KZiuFlSbdHYUnQ4VV44i+v/Sxcgp+8VHW37b
6daZWbK9sloEMmMxOGyw/DyCeKUP/6Rq0LvslvsNV4PxkpGkHtATH46WvxX2qZUJ0Bb9ivndDIFO
Zu96skMKguhngR05cTxjSdV5b5zxqm7OX6foT3M5AUGdxOYct5LtAlNfHYAdGRk7wUz32RRD8ZAM
5dV8/RRuM8gotIEWn4n3vdsd4bMGiKVskJl3Z1WTtOmDgSZkTO5N6o32T8anpU39adxF9258Nerc
4794iz93+JBZLuJUFarbE7LhXE3aGCz/h8eAJc5WoAK+Z07V1Vwctp14+Jcm655mz4mY8QbZuw99
IHmk7lyTnZM8VpgNVF9W4V0PKmy3D6eY1wYLTsF+kjZ7SI1R+ikp+ESZTBlMsW+jZvZKfn+TFlsi
Al0zkcvIkFM1Gw0r6JPdbuhZRQTO+WRo2Po4pHiw4PXgO/aF0IZe4vTag6v8txbkvHDSUXM0ivtm
9deC4SsalxQ0ExuEHMd0z+pfWrvukBOxgK+xbtMh+URHQtOg1g7otvXT32hGVgFGUZXhSQVEbZoW
M6ZFL9HoOLvJd6tabobrXsGRSB9IOTBKoXGK3EVh0xgWQe8O0ZXODhkHl2Kuwz9ZYiPOKEO3k7Ms
+Y54ikbjgPwQW4gMELDfuun18m1q5AO91suotl/KL9HLADlEwVR+s3uHm4uxXrrtZbxxJ00BDse3
98U3I7SI2Sl5lx4uM6gA0XghMMLNPwTTBSW2pxd0yyiwifRwMfOWS/fuhOQPi/vAUyk0QeVXGeFL
Sk6t/1sRBlYVC/hicKC0B5b4vlGdG5cfx139/Pv5jgUbRZyRyjdfwauvaaLFB47BNbCspv9NShQV
rsw6vnDMCpzsCgL/yujpbl5HFdTcb6k0rSZiKXta6D7LipFXbva4yzqyIYSZeu5H6JSSTmscoSPn
FJ559Wn3Lgp90BWp2tDAMza81DA9L5dG9tTE2eDFDS/DShq2pGkGtFMloTYuCT3BHqEa4yqq1i69
vuElxvoHGylmB/6L0eUzSqqFa+qeFi1u+lM/bMUv3R+c54nyegRE3/+6it1enECQY43Xp1i8KSX8
sahM2A0ndPa7kYRA1WqqVz3V45xJwaWRAgnUVyw/haKODwTsUCDmtvyAkfXy6roKHqzp2MthZxA/
16kCOpUxwtuw6CamhsaPGhVbG39B3EVqbDa25JbClaKD2QgqN33PoGomh1ATX8jri56iYoVUOL+0
10IVOijPxmKXVg/HIFf80pc/LF8bktfbkOc9rW+q3w0WPLE6HWkhtH6QtIOMjOjD8b0PpAIoADtX
DYsYM5pvo0IXtDpY+Qegr6+f2+SE4yEV9rrroI6KyVflr3Gin2GBiqTQ0A7cClf/w++a5RKaNAEe
emQch3MgN5kLUjcdZw9k5hwXKdOmPtfiXQkmRtJes4EOUx9zOpmQQKJjcy32ujirPwCAjj+vfi12
O8NMoAN2nytCBrsXyI5edba8tL2fHOzPTcd69yxKd7I82QM5LbXVHhL5cao4ttW725iMzGEf+nJc
JFZxpstPWJma12Rti+gCHjfDZh5nAkN1w0wvqerxInv+IKQlRXYomEw7sKl84B/yvMQZX5+qpYZo
AtQmbq3YSwrNhVcHT+0Mph0jbEG11dgaeJS7aZzsJzREGZHlrcAriWCSFJLbgZ0xPkBgW3oUd3UV
/oXjTZsicgeq2ielxkI0JXa0OlVXlg4UDcSXvgKjxmDAfhXCtfVjnFawPIUVjvG8b8nQTwvFZMjZ
EA9TXIG3xFXC1QM6uMnsFcp4vZOdJ7LZXBHdzvIPBh9btIpmcallWllZ0Ms7naa6z5PgHFmt6fHz
8wWLTKhn7mPA0ZhyJd4du4wC94S5AjZjD5QeAdC0/hgvj0dESPEHG2FxD+SJkAlzugPmw4r5K85z
Cjv0PoN+maNM7eee4PftK1lc/DE4QYfYhiZonLR694IYAbVsjjVoY40KQSUjkBki+CEr4cgR2WaK
BXLqXTNlthKuHdoeybs4ULCNi0xTmS9YVqSdgx2kruQLFUh2/4RR621JF1hpRYuL9FfIJfEKyaLD
HjnSQcb3pd90RzuwjONnCgvjzotm23tyzLCYTu3MPNIPxrzI1yk42FtRoRtv2BHpzs0C2hgnFft4
WVoyfRITa1xYFKkjBaqMkaXelWA4YPKnhRtgSkF4hXhD3Agd2to4Hvqd1jMNZ+RwBcW08jQCiI9v
yGf9dF6qYySYA6UBfEDwQrGK96LftG+gciQ4ZjnUc0zAEB/7oCFwlDa2rCnuulbzmtMrXc3HhzGX
NdYqA5CsUV1CCXxoQGuT8OgcHqQRCg5wU02kSkFVKIUxPpc+h4D2BNIYaThfyezwCkxAn9TwN4jE
ZMJxLsGj8e18h0rX4u+UQsiJRGeVxOlXxJPucI7v5g6lAWTCW06rlg+okWBQX/ViTDicvgJVw8Pl
pGFYvIeQ228QeVH5IFUdprKNnWYiZ6M5PqB+qBoKg1qSoJSNDG7HShq5twX69wUDciSngoFgBHYE
xxXWkcK2E1OZpzf2fBxZ8eo4ILWc1lrTXrwPSMtZ/uLwq46TKLYMXoKkLEtlof6sHksEGKYzxb89
Sq3uUnAnMw36UIhnwLiNLG55IWmcUcivY3A/fYC3IbflwvMfTKM4v9p8bG6ysSHqoBIhaldICKf/
fh7LkcX4bdDLylWjte59/IRK27ImnVOHrQfOX1lSPdj5bb92+4IZ73d3Xc7KsvKEqXAZTbjx/Mbp
b0j/QE3dyzQYlCnqZVFIWOBFM1EqNztoANb5APStmjTAAEUGv8gobr/Tb+aeeXwVUtpej5Ar1isu
PPjEUtGuFOmHlcUSGCLVe8h9/z/fD9Mtdgcs4tuJNg2GLJcC1LA8I+Ru5GWoCVpHqzkMOiop09q8
jQ1kVmw54Vhi/jvqcKhfBFZSLSfnDu1F+HyPRyJbEkQ9jbLT/c8oPGQditUwuSISbuE8iO30LwgG
W98W5Mfm9H3INceV5qHV4zqAa0Xt8PCqWB5yh9yjOt7y9EQcw2mojc5f+tWegWRH6aLTiQ8Aj3JS
8u/F5umwvZIUCEH/KARIbGx4qKYOhd0D56yK99BxFHYpSzCfdyRkQm5YNTuRZcVmvmPB0YZL12Fy
EpmeE28MWNJt7bR3nfEI0moTO7HwaCiwBGploMZ9rIp4CGcOLG7SvOsfwlLQqlkC5oo+++88MR8c
PlkeT78/Y7vFWzUVOIohHoyU9hTP/bo9nvYsgo+JRj6u59o4pIvHiecxSX7yJhzYl4SzscUfIx0n
v8/9fBj8Oxxu7etfbU39QvntbX+aOqJma30MP+/37O4OHnXp7HrZCxT4TaQ/a/YMMFdWkp8bbuSV
YeinTeI0Y86ESDffOiQAbpaUw0flfbtg2CAwfD+08amalCJtfgwlOD0S8Y280azFKm8BMFTzg8oK
zTx1sYKgfcNU5N9gVESMSutVY/R9BwwkGCI6G1sEzOhv4b2PeZaGCAHc74YeDX/5jU5DFd0dM/BQ
IH4DZIMKZF1QCjsLRxF8zxS4xA92NyETtJvDjROJ8grcQDOOSpMHYBP6ZMZMuQ3bGyI/Yc3B286D
SecuylTNaNdPwrocdxezCyWF5ltxH7hFT1R7t/LDy7mdoVUkVC0Eqw/73u2kx+MGyxuqu07cS6Mx
1KNS2N1W9b5ukZk9QFVddYy3Rms3YZoGHjhSMscZZA7Q0mNd8DjT/BTxZNoexjpbwa3y+BqYPyHt
1fysHQYK8IshX2hW25lRDP5Oizy2N57qPwWJdHWJafkvIqnQh9Jfu2DXeI4uoVdH3FOLB+ijQvxc
lklxvcTfVDsOpzSY6YTkQIeJTAro9o/0YgjXbUfbetpRd1Z4BCLRRpN2OCZwBgUpcj/rfbk1IFOx
6cbc6FwKx//roX9w/mNJesOZiLaBfvhsP6J1SOeYP5zFssHLDjKLBAlUnTUHmlXcgYq8mnStTM5e
qKeMyn1iZ6jOibuuIIaCDQ2nQgZcsm6SiVXFHRSpRDll/F2ejS+jASFuX2pTfcA15CqAVJzGJXT7
zQmZDS6t4ugfw8rYjGtUD00aYMn332HktcAPDR6nLh4OM3UbDv4OPWXwNq9UeKx/2AYn5RnObbmq
dEon52b4Sd79Sf032KFmvE5kVMSIqx+GDpaONOaCdQRn5wiNHkzIX1cfJ4bjNMHVZaIW3TLRDita
aqOwYElApzJL/bi6RuETjzk0B+Tx8Q6Ml4CTTXjqHSTWWEoI9ddo3AjVLhxWLpoXWVx5HcLFOqgJ
AHO69J3scEnGP/oYcyznH94lEs0xYCU1x5sD1Wy4RZj4JD6LOU4pyu5vkPIgW/plrnNUwR9JhShp
vcYdqNDDWRhbW02j2HL2xPAea058QwnReYvo5O2w2DSjVD6EDHyIo3k67cl5YeI7sKilpN8kGaYX
dSf6PHZQeDthvkhnwE70dEnaII2oSgz4o8URoRJQlYK9xLXX1B51Q+o6Nc8qjgcRPc54RJsKTgrn
BjSuOT5BZeR6La3TmnO+9C3wCLmAPx4cKNLrCf9AZFmRBpfHqJAKqB5cpfu8zI8MhlW1a4gLZ8QX
tYykXoN9vEag/gMcJM1mpWf7jo06Y1eH57L/FhJt8A7q2SKn9ef5g5+6kttVPvX06wECplTN/fnO
p1LckyYhYVFpz4r/ErqHI8LmVnaydokgMa+6BAt83CraPRHVfOIzG8Cn/jn91tscNIbps9rWVX0a
1J5S8N0bbIhSwaXkr4kBHxyGCSNr/BMg8/yFALXbkHT/jnQWmYEnTZy++AGX/nfE8iM0+Nrrnke3
KnPiYhJBHvnOG4iy49n6udldNu6l0vivsESuEOoqLZ9DrpOmlI4zlE9S9eGBN1CTh/W8aHiHd6nW
d9gSPgNtv9m+6zNU7m6q5zhdMlopzWHkGXlG0Wtk7yQEpVDt09j8d+y7OVRGOL0ON3H2EQrA+YCL
sOCKgM4PJsmCxz5vL2RULKONO4CjR1d94EXSKiZXyEdIZkd63epX1sQROR4wFx8Do640p/VAayNG
BQi77HScmkQkzRdxvEjhXxiUj66LRLXk2wDXs0bPWh77Fq2Np8uh2b3qajVwdBhQahSnqV4NAW3k
V9MSvuyqgoirq9WzeB9TJ0nQzS4IfH47FPjl0HNvVPyYEj4OvDnvfmiYT6wQ3n7px0HRn/bdFoMs
qeRcOgxxou8LiINdgLB3hjE+B8XXf8iHvFu9U2k07loTXqGS0nGbXwQui9h49V20T3a/H0C4Q8VU
Xwt9BvHVagzePwIJeKJDAJ2bW2+wFbixLcL9p2Ys3n/S17skiF0DnA4bNllCsNGTSTVLStKHaS8H
GbPWNI2yWysuqpFg2yxomS0k3YSn6e+Rk9EE/SAjTkSmPPigGC4n3pXd9k/qqUzd1PZSmtrPzKND
STQVAg9W/jyjx5TiSiT8mrCEbJZ09Nsyv/tQvqf/X/p83zM+1C/MSv42mRKor6pV/qCUSX5sdCwz
IRnxFMwMBxB8yYsRPejidM1YoSiMh6kZZVe27nqCm+Mndntb47HaO+D4Wy6TUYyyM/yVpNgtukW5
FMgI/wdsLcDy3aSmG0u1xsYZa7cKesv69DgtIB7b8vISvs/dr0dTahRlftuikwxbVJKHWSly1Py9
3LxwpJO8wL5z4pe6OUt0AxtilmmR6d5Mv4Yy1MEaxzyo5xHWj88vpnizIyCvWxUynzD+b/cZNk47
l8GfI6B/F8JdQNbmQjrewYTlHe5s6EZtz5VRcM1aLSof31Wh8kyCxeUJMjo5wA2xwlCfimrpUWTt
mDtsl0vwNk6CxOVbzA9D7zEO/YIDeobciH6QouMvpTunYmuPQCf4lc2sAsptaRwesTC2H/d12gAX
CxMQTlJBWP139ttFRUXcRwHycOgVVudobTLNo6+93LW53T88LIRDcRODEISG9/cs0C6oI5Mcz4YM
2fnQKnWozSJM8iueZDOLqisTlbvmBNI0lp96MAaeZi2qpF47wCw+1TsmtbW1q9Iqch0JKQ7XqBre
nicU7dNhM0KAxI8FgE9KYlNPtvGLV2aza3WWHWRNdvr8wKcaqcxGgZDM04t6mT4fcymS3TtYO/62
4LZP+vANEd/4OEnU02XPSAm0v9UwkF2S3JwqYhijJqVXkeFl5J43I0OEDBAIj5fCzEaRHleVbs28
R1iDpZydmvnKwh7BWHjsi53eLvzM2oqnqflQw77RQkasGf9jlyeDUYZPQyKE9izFYDtrUo7/qWSH
OLWUHifa1RSw+S4eNPV3RVfGXZIBcQXr0lEkmS+768cuYJbtJnDC86aRFVKo3AdsUjYbfOGmKVTA
Gr6iV0E27YvyAqmcZ5iXOnXIeL+EElKSfgocMceqNSC4GBvLAlcd5iicqdgcVcK6RUaem/jL3hGs
4Boi4QWnR6JFa7l8TqFQhEHF1tXzCp5YdethsIgTqtvJH8dd6dxS5udnrAHGrI0fYuPQwYSHI7Cq
i2N7TYg+RovOjbow6LR8x4wPUTod0e8xdkMH7HCou9V0QnnFwUlixFhdH5MN6Li2TMNCJXI0pell
Ert+xe2Mb8Jafz5qhu1n9EKEnYDhBbfb5ONYUXq+roJHlBqAj8bEDCI8IYOFDDrArSNJ3WTgshw9
ApXP5LKFTV40nCAWbNvX023mR72GUCRAhawGVpJ3yvLq1YvHc3CQYxpxtPYp01qpXggYLvUTZSNk
/TN3Q9sZFBBMaf0oHZIlKtSEoQvuYIy2PLyV8K/ulf3H6hLzQZsadFVesI2oTIR80g/SNLLFxurq
WbD89mtrLqbg/gDvPLZjO+hNjRV9SClHO2rR3SNmpbMFW/OKw0j0JBp6AnQmPplNiyooqj9TvjJr
/ysvdedku+J60RN57RQms+pn0Hee+tenjf0Fj0wW7QP8zCWBLkDBK6BbWulTGQ2JWs/zHpF5uhTD
qAQHR1Ge+YdLFwWyOxt5ZlUNvSEtSZEv6sNchg6tuGWQZtm8b62LUGaKjY2x0UBjCqWwIElYPws6
zbotM5Yb/lXWf3X77UloqEuImkte9/D13D8PhhZqpyMWQIv5rTgtyzSA0XXy41U85ZVFxS5mzF9m
NN3RnV+QSOFAUnSN5j2i3CaqVd97bEs/UE9W/suPbZhwm7Kwu6eorlO4eKJJsx7+ygDT+6TfczCJ
C59xsZ6hV5I4GImMIaoK57mjAlv3mw9Wwd7jYB0krcnetd/mD7oVxKDllPbsCGJGDn5mgmUZVmxe
HkVQQcm/POPi7XMFcMOb9baHR6jORYrZLhOtYALZCpXNOlaqB5HmJ3UEZTMhxU6ob4mdbHLe1xQN
07JDK+rILhYpTTiCd+8z9XSmR+KXgVXFbzkLvlIw+WQ/HmrglAyT4xUxGb4f9AN7HS9NKsNyyVKw
krHPkBx2CgNUKHomt36wIxblgZeAiGzqqUMGYKS07OXDLNYxcSLqns8Ueii9Ny9apQn3X/EK7f3T
x+sPq/4H9rIY+R3dpKus+gb+WFwlDxP6PoYPXjM+aFrgxNwSH1GmtE0fKzIL3lyVKvlVCm6p818X
Ebucq77XPUOpILWehjonevCfMExMQCZqOTRHdAwXLKh8a7q2XN6hKRFWLIx7gOUOj/luLoD5eFHZ
SdIN8Zl5vkRTQ5jSHJzLh5OSYHAve8LDPNJ6n3CAS9mUzohPfXLYUpgHaCcY7jHVR5dlRT2s8qr0
aegnK6qTzEBLD9G6ogwq2hCzqLqvyQyF9yHhS0DQ5XitaXlmvSK9NI/WqP5gx3b8Dmaq9V917Moh
h3h2Ni/pO5zySIuy8o3zVwspASAg52RsON6zAcQ8Izp9D/4+YjlC8YPdMSxJYewK+bQkW3BivbEU
5QZo/GY28Cx9fnY5sYtEx3teo+DWJN8x12Afovsh+8ZkNXx0fGXbJdjD6xwgmSHBaBM84Y28ygcn
31KDMe5TtTbu/MhZ+iHV7mg6HUYrrjZHW4Ep58RwPLctMaWO/jFqRDCO0LURTC+4gxs6t3iB1vxV
8p5jl72y+J9qyoUw6e+3/X5jTfXw0fegndz4zePR5jOEeEtsz96Ut9cAQkuaXa4rYnSEdeiIe0L5
zzkTQq9h/pWXP8u9BkJspB1r8ui4+pl7/M5ticuyDD+2LR9TsUwrkLjsgzWKc4SuOswgTTYL7DpY
4CWW54pbtEMCqyoOr7N583lFud8nEsViNEGbfk/3TtlsMfb6GJ096hUtMKbHoTYduxv6UV2kIpp+
XAt1tYDMuk6k5m4ZTY9OitiKCLr706CzWiqMtwyLxGx2ihnVW3bswHYzO0MZ50BR8dOL+yNkSwLl
5nLbc23u150y61ozWo75BDRTNDl+mj+AEesimzXHfN0lssxFcI1yjpMe9+pJXdhcZ2oQG7wWj2F+
0/0iYzvICyFNu7eXwWFx9jtHW/xA5SiZUG1ikpAcMjq4pzXVCP6SLgdlAZlC9TcX28bNkjcJ/Qld
ABwVyGgdn8WyaTWFw3mcApzGESSWi2++npFysg/Vu4kD4OzswlcP9zBe0rzsyCV8W7Aq3ugYLVvv
ugxw/t3HONkc3XltYZuUITncaeSrj5yAAlQyOTDeJEdsqmzG2iFE4pyFy1fMCGUp6KIPbspwYJUp
6V4rG1ZQjvpDCpeaoVmAiMbM0iaTLYPbl41ThmTalgI6vf7akxp5gXOCnlhAtVTflfZCQfVNmeA/
v+oL4/3YsQSgwxSX+L4PapsdKQSj8ceKda61Y6wh3VCvSxKv6eB64qpJiLdTN7fFQj1ReHYaGKr6
KuIjg32kSKi7AwLxdhLWf55IFzw9Kg9Q2x92OxQPJ7YXgenTig9omHAJum+WYIIrvGe/xwRy8Hby
7lrVakT6t7djDGPjsGVJ7+RhBUjx+1aFLczopxOYacV8KLeSnWHYe6HiVUysIUX+u7QhAZM7+W05
mBd9+NqjXmtZsei+nRGhJINUXkwWM26oo0SlbA1pvgivIogb252tyvA/uaGmYegOoXLv+Mhzo78a
XruswS4yN08Exw==
`protect end_protected
