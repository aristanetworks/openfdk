--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
YqXwpzoKNpQxhugogMr83JwQFKlBtYcHohHRX2VnRWUeNi6t/ZgOHdA9fPDqM8was4UMgCkVGUYO
l3Td2gbW7SQt1aRH4BHQ9Mv7UOR5BHcKL2NQQ8amuEIgp+2GIykA0VTFAdJ47hItnyxri674bd6j
kibtEKJH+Fk6KUFsgMCQ0xZIjlItT7XeZXubIznRYM4dsp4/AT4vYgJeXCi4cGN8/4hkJknXwU5M
WTI51ok0uV0vX33dsfdAz9AWAv0P4/L70d4VoXVNRRyEc2DL5a983KJvR56mAtD2wQ9znDS4ZsX5
ehC7eAD6tOghcUmo2LPbIfmL97yPw+4aYlg+Ng==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="pB33JlV6pDvtsWbqfjoouxZrjohcH16ZDSmGRl3nHIw="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
MYRF24SG850WN1IcWbB+Y9bUH1jBiDEXjFqELEv9CiHvYOQvu5q/AW3SIMdGHJlOjUd8ED/nXOxB
cHAJ89JLvCFuYUhYqDR3Fdi5WeeKsjMP8ZhaWbBx0g2LCsjTRWKICo5tZYLr8iCc+NnmPOFAHSkM
Liq0vSWfODtepaZJYBs1r7vvlhEiys/yvp0yMMqezcotj5Xlylcn0FftZHO8tKgKXNR1fwYRjMMn
eYGPnWl/CfhsLqZf2btcw6HT6kIx8orOyiKvKmHhLaHUjT8Kfwi93bpU5YjA2bTfFPOuEbcipLFr
A4slauh6+i2B19b753YTJhIRyFYj3lv7ba7bnQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Op1Z+x4RkkG1Qy6Gu2t413iVWs3II0LcpKOgc5OxsD0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19552)
`protect data_block
sfsWb166DGEJdyS+/k8tPFWS4S/8s6j30iPhxfqskYupxX2TCxtpo4245NoUmRRrZlxsg7H9CZzk
qCNex6eAqScygm8Xg4E47R/snXS6++2v1T4f79EsxNrb5Wp00oq2OOF4SnQcI3fVA1QO3URPiG5+
irf9oA7kLnze0VE2o1rFlRDbcQ0H9Nu7ADQx9y93skXzn/UY9Nb+vrAm0V9CVig/FM4i2igVAkY7
hpEl6ZCMeyMnQ6aDKckGYaIxmkQOcg/DicygumkkjPTNVVVC6Lo9RkxbkXKyqFLiCKvKe0EPA4JZ
xlLDisg1A3QCNn2Co5W0hzSvyyLz7KKGGhAQZdSjH/DjyKCrTxr7FlhgfUlFG5leit3/PYmawbia
cKMv+G61/+MWQi+irWPhtQG/0DTci3P9dVJInBo8+rNOQm3fd2dg+MBVTtZnQ9JiS0w+4aNLULeX
XQOkE83ZCVDONnEZc+HhN1sQ8onMvR4v/6+vf075ygV3aYQPQFrbLq3aTT1xGvm5Ef4XmmaQGV+6
VMeE3uXL4tLC0IBL0Z4gkcATO+LPa6iVSh7kyXS7iE8xvqWaK10s41CdW50epCNQHdjZ38j1QJRI
pU5kQ2bJy3Vf5zuCTEJaEVS061I1XVPN9lqlgzja+C5wjIwvxEuEaYBj1uDNPeK8a+po6i0AAWS/
dE5VmzcYEIZD8KeCbTtTOvNLB234FmkMew4tErcUgUdiQUq8XIA+q/kx591j1xxE38kh1D87EtyR
1vrGUBZlkdbd3psROyIMUbzF++2iHhkd7uYh68/qCnN3GoCxBBpxiTcFpSzktyfbPyYFG1WpOTWn
SSBLb6pRHCQrifO3AQtFVYEJ39v4eHCUWg/TePMJ+NsYDaNa+llDOvUF9mIbhkAfSXIwzcsBJ765
1x+QGS5ScYeEdHw/E9pUrjoR+mNiAplxl66mQ0s8j/k4wCPrBNs6w15A9lvNV7HT4WVmP5748DJK
xfKOyAk9ri1bG6h86T57nY1FkkrOsp9FXul2GJxXi3npwLOHxm3SyLcFzIUiyZFCQ/jgw4L3jaQO
Z7Ffnr5Z9d36YJ5CuOnTJFz/bO1Yvqr8mXF1d5Ti0phIosCAAh50cVh2qUbSYOlbRmYvKfABjcA6
jdOw1FBZAJIXmFqm9GdA588dkDmqag2VMsoU9Pem0n3MVByT0sP+ihT7d0MXKt8G5UoCrJuMk77B
VwdT1ZLKwKpVWPKEIAEICn7Us59M/V7pebzajys0bCa7iETMfYpmAXp0zfkb5wY83yIa/0uBl7vN
Z2bfJe4AEt5tmuGzqCO7VEKHRUjnDNNfJq1betTOT0lpNBEVY9oWHBppXlhhjEHf4OX+7D8XQPM0
9C2QPs3Elci/ENkJBx52b21t0rycBFPSXDBTRMw2Xx51KdoprYc+t0UcUs4+sc2av3If0WDyokxw
ZqHTyZVup3VpHHG/o6c3KAQk4fglge5DAfIEy/9pA4R8SLpcHzXr1mDwYipKDV8zBzojt8TUcMnX
naqgmFPhfsjIet3IMk1Kx70RzXvnewtjn8CvJ0+4qEqK9Z0OyNo40SD4UWH0M1BmCcZHn0InBwTd
qEIx7jGH10KLgG+EJsDw9z1W7C7FHk2GiR1C1HOna3yeLf+Wty9LTrnmmSA+AOxmu7jsDNMqluQI
F5YnYme/WF7O4nMv7fesSabS6tu7SiXaXQwGmBr1ScWGQLgAO5j0bjoS5E6lbYyVOpAU/pFKk2D3
dLu5HpK+oqKTZ6l8x61flJFVo8YlFzefc8Y0/GP58iOL/sGKRU2K30cO9VN0TWKlGJ+nkfJc+HZw
AS3Zw9RTEWXOCBOyDnm595xFWJ4azPJcRBB8RPg5irTe9wRYLaLy3UG2GeM6cC0abKfwQnmZcooB
3ajGae0g1xfOKALpr5CvWCVq0vw9LTp8hCA4RkdH7AfRK0XH9iowTnYGiCtA+T5fwUuGqQe2KTqP
PTCBXX2G6hdf4Ry8BzJn0xpzj99Xn8O58bbsKyt7MMwnWu/yF9VJouxscY9aDek7CLnPIgmOzrbu
pc8LK4LkWtECS6Vled1hpF4nvquCpvrHYl+fWTahJRsJnB7GWYwM7Ode7+vW0W7T3khvV0SHGxkv
fDwjddPa4cykOgDHgnkBBmi0spFZpDCCVRNoc9UchvLGh5Rkv+/xeEX/qqfd3Nkxa9G/+RPv3EMD
K2CHVeqWK+O+llxR1jpyvezLG1P/yC1Q2/pj+5dsqNGPW7zTORUVQzZrRt8QPLYNnsQkwe2nGcyX
a0m6UjR/ul3gzuy3b3HdGC7p06D5Gh5W0vHM5M7OWsxR56gQZZa5z99TP0zcZ1YzWcOZ1jkCciJC
DvdJtgGsBqqHoMNqpSLjXV+mePBFRu9iewMjA99D7YsQz11rYK1Wvc5RcCn3oONGcxZYVsKodwrm
kd2z+Unqr8FMuDvxk3xpuSE/ImOEu6wY+MzMQ7+L7X8V+Ar9xjuKej7CHpijxoZLrFU3pF2a8pNF
TkuKEDHWo/Ne2pbfqGee7ibjMcgaUGvpliAUcj4mcw8IYrg8+hKW2hL0HCQyAq4NRycEDHhWeJDp
IDmDONfoU5IRWAJohPnKzB0tT+S5N8I+fhdUbh7hfy3mQeCHesdCUqJqsVC5uqUnjtSG2n3TowOi
qlTaTUsOT9Nt0uI3n25MWzgrqmgvqFhqfCc65Fx6E0VyxGOzRxkJwXp97rK5eqCY4yubAP6SToyW
HGcCx0hmYN/oDwVRm4b/vapzeNnnlxHilSW90K3K6+WwKDuGS6UG4+C52a/lMtzvKJGnxAQBma9p
OA6b12ByrmIQAY9fawG4z0AC7SXcO5iiWL1ffwa16MoLGa+EZfub/4883bT5pIUsakG0jwnogMCe
PUZ3lssJKl7c8H1TYMi7yJvbfEp6A3MNadp0CJnccI39SFOAOfyb6BconTZeAs5gV8qEejg6lrqV
7TgtNVfkBR0BcEO2Nx98xGAGL0E7B10RwBDPJrNsvPZk5RvPBvkyNuUu2V/5CYPttd9hKZfOV+gX
RJ4lcBXQs5FS/wEAZ5mPgIl8v2LzmlZNEVlSI/CAmeW+r73ejFaIu6ySJw7XPpNILQqf+NDDqsHH
5KD90LSpXXaPhuugI4YojOxZHjt2k3XuqqcAMBoVfDba7gnkJwHhArVe/xdOtZ+qDrdLLYcNyBM1
VGe3HTwJYYZ8sPs6kGsFKB0zeeP+3Eg/TfZtYUg0ud5ErhK+vRUC/9LZDCt2FhaknVnEGRU/GOf2
3xf4XXHH58hPQpcufFcSTdu/aOs6AbBGwLF8nlf76L2MnaKBRTMxRrS6pkxU02v+8GvXtxaoo1ck
318xSPORZ0ovDBY70VJIkwdzKEWHhik3WkYHhMH4Jhx2GfU3mWmislnVpTEk2+jr1YhDQe+6nC83
cPKf3LCy7O5StBFH3cil2w3rGwfvctVUvRywGI/N1JoeaqlTk6PvqPhgSeuXK5zEiRYYAvi4Ym/9
JemruDEBqIkXig+cRoqTG5yLgaFamPAS4Rvl75xd50vUaBFQyV7Eawq/bxp0J0EwIY48Kbi4E1uh
1smiCBmAVcc5+Ie7ppELWhEvCYk0POX6mDiLnPaRzgiccQMNKFkRSLrG9sTS3nobhWYKu2xwT2Gl
cVE21PYUw1dG2oXLsoFzBQxq/EAzggy5HJuqMQtfQ9DBO/D86b6NemmoA7UgOeiyMjAxQtxxZ5RF
dL8L9+LmbR9fUOnPdyuaJM9m3xJZGclWDngz0O9vWiXSo5WOkyL0h3i+OGZUlxWFIjcNrKl3/51L
IDqQ7d/Myk7Yu8GAu2SN6ldqhGULIo3m/dzVEBPR6bQhaPyghF7aSFThko2OrAx71eaxEaULBPSM
Rk6RktFN7GaSDaUCHojto93bwqGJ36icxhYPoKmPFvCk0jn1530Oz5xORsl93A8RIYc5Nk6xDbbV
NNOwe6ANN2dr35+wAGxex3aGpnuNG4c46iF3oWxe0jBx3i+e9yqaMgJCNtLLP4q/uTcbtUsv4dtK
6GAbjkG2HakGkWO59FRzI/le+CADAW6/4Bb6DQeSROJIXvz7TxwlPC9cDPpR6gi341DZrM6bWvMx
s+5/TUSsdb/y3sXk2GQBtEjyK2x+DPpsOrDtgkWz8AmwB8a3A5z5WzloaZWQpCmcPsCSjquRO0Wc
w6SfxGBPjxuNxbKP25hM0nJNg92lITytb5bHlRDjZR2/UEvQ2Iw8YFBK96DsJDSnYKCyZ9W7ViK0
c7Wv5MS5FdmQs9bsOqpF63TxmT8L1xpKgB+QbViP4S9gUI/eFX2yBi2jnve0Ckfi/2BgWl1MRk84
oBANqE/mHJdDM3wzfS/HoUNWvZg++/3Nj975HY4SDoSaRRGRtUiJAiHEWbzKIs1wj6xs9CoHf66c
Rt7JM+ZDHcsmwcqt/XAgzjdZNSo4voFbkqSGsA3U4z7KgDvSpi8F+0puW6RssrpdcpJdwBXrUSmy
xuNyV1Mn1ooiz+M9h0ZocEteCyAiKqMBUp1ziU1QV44azAyYPJkHT6LqbYDHS7Z0HX5b6/fUCeXH
jZYy4MxMr1MqfsVBe2l5iHmFSuUvY+/CaY36pgFJapDUZVzf0CdH6JAHHxqdC+iPG6qbS4NTmIlX
7xLDJ3/F2xWBoC9rBo2dcOe9RMApAphUl+3lBxInqzdPluiSgqsgd0PT/GXGK4+vZjMhYYFcwfSu
6BG8fx8GRuU5Zcc1WkHmGaazpXgOw437Ecy1sKOlR+oFN9IvrD43cKe62QorZuSRUKF2mLbhxt5k
6NAHvCJvyORjwIvdwc1JcUhU/gJcoP9cu6GX/b0h87LP5dcY3m87DWL/nr8A77vfyrOUSnYOj/Fk
nQ8WV0ffl4lLICkTVymw9hd0I2llu8JhsZAPCyu0a2ZVfrCUL1M29DSlSQSB0udaKwzpNEWuqPqc
+QuE18o++jEn8ntsYhqIz2VLff+oLBc1QJwALNWTDQtOQv50vyVXPMlkC+Qe0aOt3hS+xkHuWOye
TRRv3roI5RAF/j9w+ag1pVI4zC/HwkaIYvyZXJzXdsWaBy9GqBZJvhQWu7bbmQCrp38Jl3J7Llta
G+bzt1aQySAV25gNhWQC9bCzPm6S192OfvWqUHrNcadFSrFPKRdZpIcCeAIW1LULCdydH7TLPhnz
npkmwVv0DFfxWT/tOuhDxUb0gIEVykhznXwOSBS8xdDAdqRIs6rsPRDgXaP4+Swxw8keLP9aoyyo
X52rjAbGIJ6sxzss8CzAieUkXDJ0ZpYXdTOJp0mafq2iMimlUf3VygmvL4V1/OZngHDlHyOZc2UP
vfZKm2llgk/7j1gG6yBzoNidhJuA9hZqH9QFiq5SMJv7KNM2vq89I1Wit+NmVOCKvoq+bpgjiNNp
D++puXBLSoYq5MiI22edeIr+dGpqNu/pPgcM1I2qc7+Qo4J2Apdex2sDlNwT/3q1KIAPllhvKUJO
BTzKT2HzRGUHw6x1HoJdoItKG0PLaOjq7vnQyA+2YDg0MNSUrl07E8RTBIWIF7hTreqLm/kzGt71
kT3QvQSQwhgD5k20Yu+eft0+MsFRyCgxuFhTPO9Eqbt7b+VOElMg1WhrBbIk+Scw+RuuEQzjqxOG
V1PItcqDr7CTHr8lg0+0OENTQ+QsbIyVO5s87RvKexA2RYdnvnPy+ItfdhIRISBpI5xaacLCJ950
ggZHNE/QXZgVyT76PuuUCPXXJMtPk2bIOcxkpt8miNoh3qXzRtprxEfUOlKNK+T4FPb/08SVIXHj
6sTi1IVUr+7zBHLe56PpeRw+3n+m+cQSTohYqwEodWVJtAMMcb8kM2jWjPM+FJo5GSqC22ep0OYd
ty+DdNrvI40wYLG+9ZbZ8EShF0dZcfaHgsjLDS9GwRGc45FLKCHADybi4A0oHsI8zH0f6MEj/SU6
DndEshrwyReGsFO+FwNfn+Nq+XGXhpTvq1FuepticE2GAWv6ZxJXoDwcLyndWPTYZxxBAVbzttKJ
MLcYjKHPjKkSfBjUo39r34ABpSG5BgMQ5dBhGx33FWM/0MVwIvNp62kpXur9H6Enpv+U06fmmzfP
WSCI5qiXYmmgc6BYGxsbWMGgJtcAfPownvNZ5McD9HczWmOMyihFHWebUnA+ie+w3i2o7M9CACXg
M9tGM09Aahex4StAbHdhaokmzPyAdpXhka1Cfdz9uQppuN/b9XGBW3mTlEks6CaX+o1pwYi+FFPf
BspHn+XizjZvIuqoTEh7iQc8nSTxQeL1ejlOuewxkeiIEYl4CZyo3CPKdX87dHEaD0ziMfgKuLhN
1b8IGrcVGIuDkMosQ8YDJXa4kdcGmQxVFPcvlJ55uQvOPcerCk/tilABIMFVx6/Ideq/w2kkFy1t
DCRMbwewWuchSch/QtxR0ttrVl/FkfDg726Od0zn+mcnoqE7VxcEUAIpnjN01huMf0Is87x+rurC
EDTOE6Gp72EVb9hp+4BW+mbx5bq9mML2QnMck96T03Ctg+0n7Wi4CWdvrJU51I2Ewx2WlFtWhTne
VJjs40g3CIEdrcxpeZe9uOKuwD9IAqEU9qzjcd/8HvY88VQStw2j95BRAUZnfW8nf0BkLUPDHhhl
Gp0o2VqbyGcG/CO2yBAz3nTymvuBoA9CHPpGgmxbOEsKkUswK6qqiDANGF2T0KmP/rcvudKtk/sR
wlHSj5uXsVUD/cDa97CQn0MUBGL1W2bhj68KsiR1ntOpkHSebBTOqfWmygyKANe5WgOvJkMDoIwx
8is27tTO8pPGOsgnGN9XtMr1/Hj2FVdaKE4gPeY4PUUsUyY2esW4v225W8AOeXo6/H6pgepNW1Cw
Z0O7+qZk2uKCepp25+DvQGFPUpBFfOyGk5Sl7WQX91TpF1hKsB4HKyGgRNdjDivoh0lFbDWsveOz
jZ8Il54jA0Z8QwmDbri8LG4YChR/GYzcWurPQyl6IL6EXJU+NsqEFbclew7ZqEtTk8mv7KW3KHVm
ZXXGbrcX6dS82XYWCv148e0NWr3i6nph9FSRlL0okI+UygJKui9dZSejHGOOcLquD8Y7CmuJ9atW
Knp3mby+2Zd6PparVAR+QCN3ihv6hKRXnHywJK8BoXwB5oYm2ahFMofa1mkGxIAc6n6V7ENgcgFM
91WETb4BOifQflcg2FuMuyRbmUD3IBTP3g97zLnS5ko+41IoAOPEnVQsPX0HBuPvC2468MTyMGJ7
gHNU+6PH1HYPHS8wGIeK9bssHNPCM8gPhk2dUdodeQ7djlhvEewi7AEingr87th3yP+z1bY+4ZtJ
Xzf9Niri4/dpJV4Rwjm6VBAUB+1dAg8wPMbS1mvncFApCzrYI/0ZuCvkkOTPxN7pMD6/bYq3PYcU
0qiu3UwZ8zQleFkRQlaPD7C+JRjpdB4bh3VMqzJGDiijT7IHOdcUT4wI6hIQXtin3rU4PtJUsEt1
0n6T/PJPGOKvr+KPspurHVmbZbGnEM0FUVZl9Keu61oH1nCoSWgvIsnxNtSapSqCGN1fMcQSNRJd
GpqU+YDYueOIYX/qWyY92IDIDhBkFWQcnLDSIsE3VqoR0W4yBP2x886U372BGz6p+6TNmQCW/4k2
Rjm4YT1iw1uU3FFbJ3ZWOnI3M7PLHJCbB4sE4dheoaR25Q7jiCg6v9PsH9h2FObaJCJrz9jTr5Ke
61CaAR/i47pxdgPtQObZwQSYd1hIBUsc7S9O52LjD4mkc911YuoaMVBSvwrE9PTrcrHRf9pDqod8
vc3Kx78XoyFEaxe6k37PaKlO/Y8QkVlSAAjvCbdRmJ8TFHalgVuIqmhGPonFnR0sILhUkwJrZZPt
hPZUFxqjLoSNB6pBeU9uuLlcUuEDafgPSJJmQk5uFA46UzpktojP/1XKBTMUED93Qlq0HeXRHJZu
5O7gjbh64tGtqNWJb2zs7x3MXeC+RH0z0Gn6ncKYlJmu4OaaAA/Hk6L3RV7ABcNF0E20GZIB+1ix
CYdgbVeqdk1B8uI3YIbhJuPnIhCKqngSLj/gBnqTTOu5mN63lkxal3uyC8BMlRxixlIZ55vde8eX
Xrs1TgtZ6dgAmWgppPdKAKMCsDM28Aje/1FioMM24RwpiFsSvWRLhkJXMohPQ3VsGOwhlAuhG08v
W+dO8pS19Y5uX17DxbW0ms5zNJRCtSJ0DFeJGaVb73Z2jk6U+FQxLqYzNeH8Mt2sYGoEwBHU47/1
xtAO0BFmD+JMkwPHbjRdIcPGGkat7jlbDA4vtDC8gvz0Od+xjH3ylLHR0IJOE91AZWp3aE59nXdU
FxGfvW47mHa1DVxmihu94Gc+7UYAifAo0BurQUsdQiWcenkV2jGWQXOpmitzyCJrCbqPvfu6pXKJ
QNV50k0GKbawuIQQxpHgk8yqO1lfTwkKR168VWuYrRyyKcmywEeJHyjlTBJhJnlWh+kjp3oCUgWI
Pewxzpnoy5zSukWvd7/HkF3MOfYeKXjLtSV068pl3B7jqq2i+9jb7VC/mSh/NVXLeMTUMCU7xAnZ
D6p243+91wBk13nb2wHtXnse/KZAcjhuspLZuEJ6MR3CQu28ohJaUJIKzhsv0sfVY+u6AvBZh/Wf
WDXtzlWEDaoBE6JsAvT5sfXJGP+hstv7cV46ooA4W1dKhGTqyII/Qp4Veq7pZtT2yBDfvW3A0Phs
IUX3NVwHt1Ih6c44NJvpB4OMn5kQYXL+DJl6ySdeFR39M3cS9y+waURXFHs5bpzfX9VusU9BNQVg
aJwmlt5VfbHevdEtYEhg1g64Xv7E2Jc/Gq9i4+v9fdlTbw5BsPcGtebI6SYE3yIQ7MXHMOceq7TA
P+Is/HPITACf7/6SDPsyUe8B7LkFyfpib4SbP45cGCAblVR2p9M9OdPfcQZUXefTVpGKlPgRBfN/
WkfqmDGeFgrqLU/jBTAdCd0CSCmfqDRvEBb9hxVALrAoVgZjGZzIFUiEWhVpTghRdfMJW7Ikr/z6
Jh82ByY8AKj0GwKt9J+zk/pz+LGJ82z6GI7z6yw4CNyWAHkrcftT/chl+a5VBgwDfl7Brpb2VZ41
34Xf7qVOBzBkfSmPRch83++GWrjDf1KbMNL9djkQ2oh9q2GHx92ODclCA1VjbZypH1wPXzUbu8AL
ORqLCAkjhhOvLrZXovB1LavYcb+825pz+iJE5CrQhx9J/HKQWCL3G6kIKQkXBDArownQKjhjdPG2
h91LkcWHQTRAHm/PKRAooT3NehBe/7S7l8s/7Dr6BdVtEJwbRUWPnq10CgMiO+mTzTngBi9RtDDU
xvkQs7NTIZ/dzsZ5fOETJfZeRor45uQlYrS42/SlskFupj1lLwMJJ4l2L3vi7eXPZVi1scfdvqmN
05C8UIB4fev7pDXNwiys+LbHGnznltGgrGyy6Z3Z+DmE+hoVyQpJwQQKas2+TLFDAN2U2b7tYSZd
UCsJi7XXNIZGBRFYbCBnr89oCbGiutwQR3Dg4ihIOKe0sPrFz+WOkQLQ6C9COSvh5WmY1vsg3Cx5
BFoIt95KF3vw9pndNCUNV+MnA1Cjc7fvZdsXOtuu0ksEHmESX8hGB2dhaBm7ALaOQU2iQu7RM13W
ZHfeEGxNsfWDBF1JIH12IJEvlAdA0zp+WEI+OtHdgmtob3wOwFAzynsrF1c8PW0L6jzlAsjKE0bq
K9EffBc7W0oBHRvk5VfX8NLsvQ3My42PJTFe1ke4fQ2zMaKI6Wv09uJ9aQJwETSeMps1z6Vpos2O
DOWF0g/Rb/JEwyQZqi2etilBDGnTuxrRJfEOj/Iey7qYydsYePIhV+ZnT4tpS5Fk8qdfGJPTrDPL
Y5xcEeGo5jvZiCkmGXKU/of91+ZbDKuCegeF4GHiq8GLp6nXSsKr9PAOYLzpcBqx0XLKLX2uHddH
VaIg6vA2iCv+pXd0xpjTKvIGvBHMYKj58zzyT65v5/Ift2g/jQQql53zRAic2YOLKQhLYVlmu1nk
z2OADSFjcL1b8CsXZeyjXgYgJvQjfbI+rO9cgmryTDU5je5fiSQ1zxDflTGSChtpomnfWjEPZlXw
0Xi/lHelkk2H7NxHQsIqWIfZcFnHKQCarpIbyBla/11642U2Tq5EtdUuKMwDpEFAFxjMBYEi5sxe
Az8lANHV6BqiVMVuXJ3vN20Xski5eCBYPpImXXtFQZQ3hPt73R1R2qCcozL/O7YGYSD9oCQt32fU
kuBTVshyfrcay8DTFE1myDx9wli0OVTzQbK5Xs+3AHvx/5vQfyMkSESAH5DzYzwDIlJvkqlfCDD7
s5U+fYb6CIeljcTBjrgnAmE3I8FLn7eLhgBweSm6ecXEgNGV/F3Dfuh0WtlsCdhFpKZvA74eo3FM
YY0IHQcruLLqdfpxKQ/53h6qujN1wKQ0bEM5a5/pDTYTHDZmM+wFhiErwSfP4kDaKI5lO9r7kSw5
eBdarT8IG3V1DiwMouFRo39Wsc2fLctPLjaVpzsy0VQQWsfRvSRZrSBMOflev2lLVWgaFZ9b9szf
mybYMVmCmnzi2dYHagEmWVDYg5jiteSW+Q7neQkMllbOAy5WwqJXyM62Hzmv40jvSP6aOtMVqJaO
kQVVJKHMkAx3RuYnp8xrl/kqbvAPHgey1ahM96LStrNL/PhVhubFa9Au/hMMp9i+bDz6RMdmNm4b
iCuwbhggZSVwkHOXr2/mhf7pXkv7l1ca11kh21eiM4mGX4KjSMVurXvej8dqgg53TnjU2eM2+VFZ
mQjgbElrr7yAkzjjGinuVV89v0MgZjlDCsFnZNV6VqkrRj+kVLuBH/JTu8b7Zksu8Eqxo0NplP87
WEsQY9r0Ii+TVrVbF4/KptOVKT9FDgb0n2UtHS+fgSAYsmc3sF0c1CjX/c07LHxrCj00Lf5fBY5u
4ISJugoRNnk7vUp5MpTt88ZNqb76Jbyz+BChNEwcOXXuvMeLxtfE0+Zx2qnnvqIEAEDBxPE4/dNr
UmKkBFJX+hkwes6aT9Ors54iDydrOhjSDMkrHdbUxSCj9GibRljRhvdmYP+mczH6ZrzxKkSB5NgM
/gDX2rqf6i/HdUhoQmW20lzHKpo7Kmr8nCcZODhohK1eLbSGdVTudgYX8PXhLojQxjB2suuUegDn
K4L4l3Ji5UTCD9U+3sN33PeSLbK0/5i5mZPH0r15/k8VZm/naRZ65htnNKpecEctMGxhV8JSp2LT
lXeFBwxxcgkxY/5l0XOloRcTXOxrsf4RWsfmT6IJpx3Yy8fqAj4HJN3aSawt7LP1bHRcxRchM6aN
Uy97cGMlZ9HwGUN8COzCmJzeaPECInvWlwGwB84SxHFJNQGMNWIvQD9LFtlglHj67AOF0e4FKrg7
rQ5z00hw5GoemlDZ29I/vt9joKhDoi3eFRPDw5sE2yoyIODxtsqsWH+vTTXfsj/JCiHoSw4s6jK3
1zHBaJfA4MYUQE1bLogqxZVUbgTNwupn2Lr6YhkQulpf+6/oZT3zJaz/MlxOj1hiT5q1LM3Nm2ab
K7HZSlxlOGzTSPTE7MmbVC2vUUTwx4eaNrv5WtgCQX2SPcNT58KwKFfPC9ef0w7UhKqTGlqpFEVx
TatpiGu88rAAi7hrOXyOfG7QcnKwz/4wzSq3C1oz12Rb25B2jn4AI32/40s8zMY5ciypuf4i6+xU
14HAY216r5ODe+hfOIP2U2sdJrKhfv/PWQ1OAx+D6V3SIzlbHXQ6/jQIvgscljWHQU2kdm6ox2Oq
/7+Udcm3gGc8xkdMKp1+QfXgZpSTy5RS2WVPQSATIJc0Dy7i5AkP/mvwgFjzVNhwf6aecwlycbYg
sC35bhaLtEGG9tOPFfr3gBVSwb3wGYrNhlTh0tp95bfZijXc/Gn+dLd9TKVauL84mN8UCQHwfuUW
vypymwbhoM+9kDltgY6/2BdlZA1Hs+4mi4g8qDxX2ZG8KWYYYJbq0za7WZJzdx/9LQxuM04JSm31
gqSbMPgH4cPT3OTYsZWxeQGMJoDT93JEyv2OIQp/pfhLmHfTrtV5BpDKz3xdRhwKmu9RoHKlQAuT
Zfo6VqEUpIzYykNf2ReyBqBdRGQmgx92odMsT9JBlhPKUfZEQrp9aW5E3EpKBEZCp7Rv56KHU8bk
HMnY+wWnR9AAPLb0GEhuMs/7CVHplCaX0Fs+Q4nuvmf1hYUCyTX7pxcjuf3vd6xzuGs+YGKcvdHI
c8p2+94ioYV0wn4v5Jj37mEKFtBSTFm9BrEGWPVP2l+8SCnlZx5MV2EcvJsZYgPZQynwGLLAqNJ6
znMwnE8Ta7DmlAoenHjEWwPDWmUR6D+egKcEim7o6Nh+eNamLbPxxxRMS0rrpVwxUc0Yqm7xRD6H
ALGoxmSpK67OXlgl+5VBw2Fopls4rDlqMj8gFbBEacVyFUNY9UN5OJfxB5MBT/Wx5M6NbceH3XTN
42NoPfRUlpmwrgZUadu/k+PBR7biuE+auxXJU9JmXnJeJAPJPktNKFORPuK0Al17ETE46lQLKSEf
TBQVtQ2iOyHZxkwRd4LXTT6ZSaiH4TSLan3/X1jb7OteCw/EvDRO/+aHHUnUGLnBBhLQtHaTl+Pj
h+CuN0FXIIF/7T7beO3PoxLKkQttupJSt8xPDDVxq3HMAEjqgJU817eSk6q2ABAdnV7M5VlJJJtc
/icegVxPXPHxICjL+8jMLRi8bLk/RxoUjhhRMechLkT0DH8RGUwO5Nq4lr8nSrJUb/p1dKfM4zPz
gSwFMkcjnQeICn8GFt+wveLNZy3TjSTCU0011Yi1yqpfdwaGyvpeAJAko6E0mF6Jt7lDKcvBCtO6
Kkd20Kjk/guEO/LRyy23H/Xkj3T8VP0cgjLGNNbJuHjDeT6rIBrRS1NtjCF2ccx2wK4YEED4RF83
09qmyAc+BEv+mnKfXvFc7Azi2V8YK7Lc0H9CoyCYujvZlX4Bp4sAGl7qBp07AfSPxtRpACP3qPCp
/HF4PM3mIvg+YRpF+Yhmsy8+xX08rjtBUAAmnlnc/7jzp1Oixt8kvolR4bOp0KAx1iTVYgjn5YQH
T0Izodj3rRRza0nhLOE8FAC9n1HIiS6egNV82+1zRJK4u7sJpBPfkU1s5nRprepugK6oVSJvN070
VK1qyDqdnqcOpSOFuKGO9SmrqU01djEz2jhNIsWtwUbliQhrnEypYedbZPJ01pmqN4hhpiIUOjBV
rlHf2gk1dhFjQfb10ZXDKkWl9YLhNRu2Y0mTjCejfFMpCgcWUAlErYrV1Z3f/4jaNZ2GfsiyLxp/
c3VUYViyJLu7uhXpF6a4JxqgxSfwr1Xbq/yigzv4BldFcQTa/6GwBdVh+R+77/L1g+qMXyyRYyJu
WOWOMqdIZUDU8kKGdqbvz/qb+w2HFKKr+RMem5oZsi7Giir+SkNgOyV/mgRbnbS6WSBUk3bNSXbp
oFd9VHJYVvBgfH84q/xObujaCBebjrKK1BiFYAi8c0Rjvy/NtoorENbLCj8PElw0TQlM/2ngS6ak
8DL0r5zGmzd1L55uTQE+Jp5qT5v2jEqkgzmh9ObOIP+d2yEjGzfhCMznAMkQxuG8UzghudgtY6OK
FJhm/Kj0ujjBAw1nJsJUcv4euM+GDZkGs95cZobUp1slLRGBoSZPP4TvmZf7bd0BvZxWUoXdViTv
H+GrynmiKW7gOl90zi4yZxWeic60CrdPwI86LOmo9s1LIaV8ENZjsOwEt+mi0D5znundP/EnQdU6
eOyXIGOo4JbrwXBFxG4E6ajeNKhPrb3LL9D/29NuYNpD5oqALgE5GLbNWP3I6x8CBA2qIhGRgKYn
94lvqUO5dvRK/BDNGTg5vOFF7FO3sncOlMC8UlOe8G0b7X3Gkpk23VPN7xb/u8JSbVBeAi+2gttF
5MLRtunUfjAw/KVMnDqKArgtFkolrEzWU5mYYgw4EErhdRaCOq9UQ8V4L0N3fC6OOw6YlK/8XMgm
OtDTPV+xUN2aAfb2VKFKyn5YAXgL25jBnnCklQNclbYS3W9WFbjOxCiOmwQ5VDt+GqkMknO8phza
2KAt+yGY2NcOtm7fLWxKAhP2v1D9Q8+ezEf245Hcfla05h6phTmpCe8eOs+GC9Ju22LNWeQ4Ttvw
a/++C9tRjO6v0dsUgat2Ob/dUot6HVU6FESQTuB8N0agOS+PYwpcwiEI8RRZvvLVSWdVtkV/WRhV
j2nC6EIBDiAKx3Jb1POM7EyKnntPk1Y2LReJfgf4Fos5Bw7teXjB6Mte765SNVz/GNSAs2mARJc4
2CJp6eTvIwf8S3Mad3HLOj1VZDWK/lfYhpBSVhWVzLgwNecoWfTHBYZTGFmtpIGEEEELwzlp7j5l
iBgYR6MsTufUodEWqH3Ehqf0kDfxU3HKj+EXZVthB9HoUp9ZVeLDWKK+faohYaoTdHPD9hmdtqac
ZMg/8yB5zSBVO+gPCKFFUR54Z1iSIRs2ZGXRKPXQKe46KVrr6IXdecxZzj3I7KDbEgJBm6OR72Sn
7X9WCam04hqZeAMspDP6FfEnqwbv0a9vyGSqYk7aSno96qmnyYVbPJWIRZgYGiFh2S5teVjpgiSz
bw0Cwlc9f12BPJqMpEQlOqw6n4aIX41C/aFKjGI62cuAXToM4YiTJK/uD4I9BKhVbWI+dcCC7foH
kIofTsnbtLsdVpOD2ASx4H3r7RK0WMDBjPJ5hyeq5l1XuWWZzb5In5KnxXrIRlbhZkNJfAzojXMH
PzDlbWAYsDBbs3Mf5upvIv8i1T3BcLUWe571sU8vYAnl6ssWYzJJgubYsZomANC5kUWwfHeHP6Vu
Vcss57b2XU96AOTWUv4qU16EOxVwF2QNX11f8LH7B5vG3PS9qLuW/UMbI6v2QEGVdvnZcUNlo5Rd
r5C8YJ5uPPHS19c+S3Z8vItuS53c9e73UmjBfzQxT9ciEtKHj889CZ71jHlaL1YUJcz69g6YkehP
IQqjxQJvlevv7eTt6RQvKRnMut3bpFNjP3ucVW82038uxaQ8LPeBdTV5CyQPY4tczi7kJxMhS53S
mVR1LR0Ux0X7IGqNOZQ6yrUx6cvGeSFajXCLE07u5qxjdzNihvOrw6DELSzNvAFEDJr3jsTJkmjQ
ZpnBm32V7p+2L8zpcxa/iUUL4bBqV/tfF755VMEKqycs5J4Q09GBFM7v7RxE6dedTEzP2xIYoNGR
E3lO7Qk9/xu/CAGpZM3FGl1LJ24/qQmCPO7HMz/zHLxGZTMsD5DaFY68vKQg/o3U+/VbwXkWrblQ
EN/Hnuhh+0O6/Q5u7aP4o105eoWHMjU1RzajVScJRLLvg5Hwfg6RLe2nOfzEdQTpBV17Qki1VhVb
FK6UoMo8HthEb7AHq85ips9h2OYLUZayeINVvJOl39WEDtwgYynGowgOSn4Fa2BRrjqIX4WqaOXE
+pMIYAva8BH4f8hoTrbyWQ7k1zq1W2Ez53e3vQ4/VXxeZei3uuUmDS+2LwnTMLrOvJtHXOvAbHyA
qif5s5jXVduuo4wGTUyVJvXDFJACa4O21DGEJgi2zImDwvwdK3vcwbH4Ir/2LzXqjgyqDHRrhmEp
sVZlTpBZNsF7tzZ2T5lm63+gbQgoDoPXkBBmPymq9N15eqxHrjZ4UXd3KyvMAuyNO0HtmNY0q4Gp
yEbUzvyvOYH6srdTxPTHmZvSn/f2fnyrr3vJsP1RxjhnPPA4YypSF/rHiU2hg2sTBsbVpKFgWref
q9EirtvLNePdW7UoT1MJBM2O08Bj5C2KpgL/F79sfo0Bqhj0TOz5sC27ZerMJD5m60rzg2MvTkxO
PH11Wv8ZH8xpmtxpPCdS7T35Bi8cvZ0wlyflIFazkOBr3GgxKK+RLQic8f+JzAdK2Q3UudFlwKxw
09WxidRBUrp4/42+1LQ3X9Z32epUGrVTpq+e2Lnd9nFH7if+Yeu6ErnNDalQdTClIf0PlV8Vszwb
A6k23/wrD9wYK1pwz3J+6WbO5kf+Y9rch2x6NDUujaXaV+J9iXLmnTcZRUtJA+GysRyCP5MZiER2
ibez96FeKNDWfh7C9nvGbUrrxgLJJGCFlh57d6MPMsS1Qo8qhsgBncMlDMk7wVolKX4IKNZRX4LU
DhPVsBIy39Gg3e+DaNSJrSiMvJT0vO68NVI+5tf+pndYqOeRzzKzX431n64KvDcpT1cHQO8N/Ian
v1HnAZOeI67vaWwWi+43FIshsYXTrjdNtAzeObO84LxpbsW4NywSBG9nQW0LQIdnJYMpelvbADT0
dBQtO1Bk0q8aSTtu0xG+LKijG4uFnyDpkxkuRWQJB1t62GV+cTGYSOdf40Up+fAYfWv4yxb8N3M9
hgzhjLYtqQJsZCcbjMbIxzOc73R63kTkybeZLocyk728MfgyCn72SDyvSZImEqtPUxVVZlVPj49o
wljL3+28IYakVBKqxNp2TaYt7gpT7engzvplBuPZK3ZUOlXvF43ztGRLt3zHQf/jq6pvQTOLDoly
Hh4+z3UxY8HibzBR9c4abNrKdplFH3q6MxQ6m6pjcFBjmx2VJVMQ4tZNlnRGMHat9vQ0HZlZRlXb
gJH6Wia01LV4UOEMAwiULnlX29fJtdgSdj2tEZ6k5aO7rlh+nyrKN4itUEJGM3vggVa5kKdk4KDQ
tw4/Qz+OacVdc0Doo7kNrqOjVNLeZZUO7TUptsBoQDyIXrvHlT9U8JkgHY12jpw/Ct2Bz7Gc2YkR
Ggw8P+fep3hTPswrApODf671WWFOQaLaF+oPfTF5wLAzBKQZq2R5CPkwYtBorHNXq1qE7v0cKbYv
BinMvrBTmW2ek2U5bjtLKHH/eMGCyIDG6a7Ze2A4rV5mURbSf7NE+ukpxAvzJZkxCB4r82neWE+u
fQB1P+xysALlMs23z7BljnmYLKccdEeK/8vi1+yhQ5XE7UTcYesmtyu9p9dJiO0JpVX9I8arAKCM
Fc6WSwcPTdZwct0FhOak7KwTsDFlcWbENgEyoveGMxXXoeICpHvBAXiOOAyewrQ3We60J860Cr9d
Dbn5wVEmX75H3UrTLIDiGh6qtZGl1oG7hwkEFXze1RVMUDUBlko8z66eGx1NnZBv/+Gp/NMfDMF8
873LRtd7bmpPKhtbppEWGijlKP5n023ut1J+xdTesviUYQZVMCyzLBiMXWcr9H9xAORxp5GZd7xr
BJ6K46YKQvBjyOz5Dhmsap8FcmrjtOZkK0o55MoSHBtYCT7ZDWQEKZWiJpYCJQwXcSVUvFwDnYuz
OoN5KrY6WBaKpQfrcmebug6820kagP5YVXHtC0m+m4IlOdK9AQC0dpbDvZsK5B8mdq9wUJAXY4zc
dcOb3uQcAJUuGsoeqeL0B/QMNKxVmiESBo9bdxIvF0XykYg/VsNC7LyRyL0V5gqgE10asY9qbTPd
i/YmXUFlXO6vceVKrz6djEFl6J1cVf3SsGeL2V8T9ZUNBuUm1G5Ka175ELMLwW7p14I6YfrB6A79
Y2Kq5NWsB0uVSMEoVAiZz2gQtmbAvoiyTb9Plsu+5OweJ/kAJx8o9oCBUbJRFDrmzf8b0bQp6QlC
daiu2XS7PJ4xRKkdE1G/876ZS+iZ3VOktyLdH80Z3rKuhPP9NUbmh3H/PgVBSMeHP8tPGtPLMBs2
EThUl4CBy5xlQ3WIU1MEY7W3XljlGZI62fLgVMaMv3PM4991tU5GGoBhan8K/KaIBrTLRAnWPWHx
di/i9hMWvrpy28VOhyAE8GvrofFvtqvBf2YM0LV2bFGseY3Ga0p24zr2V78ibSBgRVHzRlLldQCR
fk7FgNCiiZhcBHgf/9xmwYaqvCZcxANhDRxGdSzemIdxC57bGOoxRupAz4pRBFCa2mh2ERmrU1iE
BUv3aXf4PIv1sOw16KCzdz9Cqe5RXcKVYulYdhXZDsO3ibAMvw121QKIXWc9s1kxczybvN96Ai09
Vp1+xupgb3RK7s4HO6CkZoYx0TrXfgegRSNlJyAwl00PSFhVt7gAyP1zldvGH6KQii4aDbOpOXf+
ZgfhaEfTBU/hCSlakxSdOC4BS/Wy2zlK/iJGoB8xJn8oC2HLrqizBp9i7OZ5oKkkvq0wRBeePAtK
hPumsbnlWJL+J+fSTjem4Fe/BrtS3QHGSw8+zht/eFcQWvgWXOO4YbLaVMPwPAN/0gTQTtqI3Gl8
5uK5KU7NWdb9LqCgcQc9er1XEbj7DW2f+Y5nonPYMYNiOE0CvTKw59NZ588rbJklGaH6rs7i16ed
yDSTaCwYin7zwIP4/v3dLIqqF+MZwGOMZwKS0k5SFrLJNgamlCTGGcUnp53ZmMUdTxdj9Np5R91h
0Er1s6MtW1ou7z5exuG0V7rx86drUw/ExCE/r64RvF1aFLB/UavoVdKfCJ4n1SmPtB6XDZtp14z1
MYKDyP0miZ2oRzTiEQC9Jc2dsQNkAQb6V5ZCmuckOlDVMoGodTu3oD3vbs11dy0BIlFzKi0rwSiJ
M2yFhwnUuP9IX4uZb/RN7xmmrNWTlB+ap/5Lkdv2tPdYlEthkIh6kIgmLiDMo/HgIwi9PwevNf8+
DeLwPmNSTefyCPkjN8/dqqXAc6wvkzsAK7rTT+BxQ4S5Uy8cMrYtZRlNllUdWR6swIl/PStVzBYI
v090vVElu/ap1p9crl0+XgvYWt9smQ2tQA6bMGEqNW8KJ3RSVZ8/ZsWzBpvg/F/uy1tMl5IUyAlA
gr5IAQSIHgdveh3FqhDztlbFp4xT12xh1tfRKSm3laCckI0tSVrdomSsRnueSjDDkWRaXC4WzTnP
mVCHDoIJtOtw7XE3nBVhMUVtVQ578Irr0kgZ5QCq4wmtqTiQEJwmrjkZUOF9OHKowwhuvslyDTTL
aJK9oN7WeFw3tcYz1ruydi62yAYZvrP156RijYVapNSK2t+lKGkUyIUIZPipAxEl2DDslQmmQQs2
vCJA+R+uKfujAm89vUljqoW4HcV4lJ/aUx49OtfvV+gLE9N1PpYpElMlmOZFlMSxiQvgtHwrJWfH
vEVpzZEPTIPEe+l+cKLQOd3i3pEG6Hlu6guhT9FXFkPDY0p47mwTc7AA/ysrfCKA1e4ZiQAj97+r
Euz0h7btcYwopTTlcLy4wE7g2mUMTeTP52rMosm04qQBNIVSfdwhPXPGBXBWnkwU8UyIdlGkprk5
ybzHUPo2sVBPK7/HuyvK1hSPwgEBo8H1GcJ14gMEZrK61eyROwq2GhsbbvaakjUS949LvSbxN1Ye
K63lpDsdGdMwSs65rGpWTaPb7YTXdo9hWTl9SdMeXELQPWoiKMLIGTRQ0c4VgKc6GuunGRWhOhiC
5aUPteaAjQEZC6ce2i66A6/QIJSo/P8TDk4UHzInu4DuLVn1BYFrmGyX1L1egP7B4/7L+gUsMFTI
emGwqWV4XCGXkPD4Xaj8HZ5F0Td5zR93rBndhHxLcQfg9kSrIVsFOlMvflQqV2TsHuynBEYg8hS2
RQ2HXl030wZyEcC8KA/kZ3Hw2/cYV8vV95MHe6X5gixPu2NokNYRZ+je9hBgs3lGFvjZ4AEz1mUH
xuwJOjmNsrOs9AXWgPbMXLHQj+GrKLx+bG5bOBtBbEQQla3jqCpnj5rE+p/bC3xTDwRdec5lFGrs
/h5PvrnVuxEbQbNBGPIqv3lmjsjc0IhfnNlUd4gu70bSTySLGG/Ok8CPrMuEKMJfqitJQQDqHU6W
HuV+6JLH0aji251NCeFnst2K727iDBRTLGuBirAwoU/BIUQvOSVlf1cbtaoGZJQjIo1Scj1LJiXa
A1X9h/bVkhhLZVLr8JqRVBpN2uG2n8+b4D69Byh9Nt/0oZ7tL+NzaF5vjOfDX1amwgNr+MR3x6Qg
HGZ2vTiYF0D/caJzLq6rFhQShGf6PrwFFmYz+e+5d+TRTJ48iVjz00pB9ROej5lkRtFa96Fl0krN
5uPXEKuX3hM8h/89IDv8JaeG06aOVcNFrU4EI9QJmQI/SH/ItbpbHiLP7J/41L1+0nhz0q2uWjvA
+pRAtP25lvxdy5sJZJBznVnrZFxESLLEJeRCCCbmbQFx9Qx2gCBUnd0ldPIPVSUsIEh0PS3+rx2m
oFIEHXOuGb+gIAaZ7UZTfSUVET36zLiwGdLrd8qjcK4/Wc/nwyZ7mJ+zZFNwTL4yl4Qqq8uIjxcX
x47Fhl/yFd6xarJitE0guvxIVlYtQA4hKfatxDYim8pqe1aJijgWwdGPUsks+Ub0b5J53VRaMdbt
Iv6tWRM5OcloqHUMJo9FC3N2jj217JOC2tlmFae3Gw3AwR380uIfB25N4lU/Ej8TQky49QUuV3cb
nzsHRanFUOqd44KbFzOsXrMCjygnfJrYed79Z3jTSkNErfRaVQh1vvNDADrTGwfYv2dc4w4YQ6pl
Xj8lWT1xrm4UvmqPT1dmLCOypBvlkKLpj8Oj0vttDautYpsfMEkT4BQ6vE32SW6pyIocJMNYJoE6
sLX8u8MW93J1sV3h1aMQKwZfdx9yeqUH+mMkRdPlan1BSyl4toCFRmhU+jYMlbXlMbzJPGxFQ5Hm
Xm9tt+KdXh5z2eEx6Y4hLSQP2XIBeErDBB+znQRA+2eRXRdB5o1djJpThAFAixHo9ZrC28xjaWUT
FhFUg4Ku79MKFjngm9bFcKzBrqYefifFbtcYjgvH3DTpZMFg4h/B8D8zi1vEV1XRcvifrE2sbptR
tJ0X3d+3Rz2aY4S9DOLterf0iFqPRJefoLq1EM0kGmvZaY3o0NRNiV2kXQ7Q3BzJjx7ex7hn/Vkv
vZdr9nABpDpYEo4gfao7S+oZ3AhVClWFuioXEV/eQmiESTBzNKT4kihrgQ9tKPWHj68B0fVBy34s
ZRkElNSDQHc5xHaJrwiV5djZfQLoaWz2cXq9C99oPE9HGZ1EFoplh4VDV46CmlcWH3hgM/9YYkUo
NyxksnZF2ihJgNqOhtW4d5naHYeUKYCAkQRbH+hV3gLy44FBAFRNJ3fHOvFUWeIAD8UJ9j3SqyES
7p2bssF5obJNXJ6T3eCnjHXY7JxIkP11vdYuT+abgRAqGg2fMgHjLW5LyrTFXyhMYfBMoPGQc4Q/
sweqsF37f/6K/KshtTItHuXxdSSZDNCOLTHB02il/LkJWGcaq6O9AzzI6uwDaNwmYD2IYvZX6iHz
PzBf/wvrzHIYmpH982mriw5iN1hOTjRm/5DouJ8E6rv0smb+Iq9bQIjvTC+IZSHS2ZIBnS1Y0g/7
iHaymfAiRUD1t9R0NaQBbSckKbV73DtTvYQY0OXV0jy5HN9/BDbxDW5rtVVDmBvu9+YpaMzcTfv3
wpduxDEiysHt4u0TnfR0NAi0XDWLqSQhZC2URtRJPikvkKs/D1/0tfF2A/yx87Y/QKYBbSrPQ4Ym
XmCq6EIOESV7Kq0d5vvP8n/F/GH+vZSMmNAPpm5TJgUbYbJ3tspvwE/XpjjmsD+dLhNn7zsi/7yP
6m211dSqUIfJx/Ck6e0+mVLPG3v3neI2Pbd+AkCSg02dHSEugN8F7R993j1X0XzTW/YOVmtaOgsh
ej4/J7fEUv1caUKFlpxN+fUc3/zW02QY18zh8LPcKIpPWoI8mL+lvde1cBv/sQOwP9alwhNJ2USZ
dcCXe8tDMQrkzNTz63DkSpT+BDy6HvZJY2zLNzIMpINYY7d8Jk1yjZSoURRjlEiIYzzuRHG4/E8G
4Tc37EuzjtSmoEIH+3dR5tD2JFWZ5A9wuW+wypPrXmXMXhPE8aL+X4nd1CnVFobPomX2CaGNEAB7
b0PXHDhUHz3VOvsv3s/iLZ1t+2Rss3j7DlyoTzx6PGtd9XfwyhDCk11Ist5T8wRmiV6aE08agi3C
PJnJNGCAMZp8mPcq6IdX5U2rC0qdOPPJb4+JVY7KBpmTD4Z1wE8uHQp43w6BcfDlqdgQphfdCijV
zYm8McUNb0hdh26RGO99pZ+hs+yh3DGgRvV+iphwCcaJA2c3ur9vhwjZ6bnVoa48WpE2F7OY0Zhs
ZqzrFJam2k8/vrK6Q4a51Ob2yZOuBeEM9cJYFBCaAoAhGQeClLr4FxL5riYM4luEEMoiQu0+DSgl
OjLalxgMraZTVGe0Anc11xj4RgZurv09RgAUROVVK7m3oamUEVHNAl7IEVwesGoO54T4TIMSlxuE
lX/d8LsI8+SOkaU5Byg/NTb8ScbECt5R8dcHwM/O4LWJ5dKvC18mVgoMJDeOES+y99qrtMM6Fg81
w7mm9Ua3tgRbYmh5Sxbfk1Mc8nYETUzRDX7So0U+waso7qUZIjBPX02p8EX7S6snTU2Jbt+Op0kx
FWpOMKMHC3DN94EyBBkgpLcisJUkm70+4wlORoxcKWBFDzJCWy04WAYNyoECQ6Gw69KL5r3e+kXK
/wJmih1vuBXsmwq8nEW/cbUWphtob07+edvpaEPlgUe3B1owY++P+EZXGevdlOIKIEZqP4sSiyXo
L9T1lUbeuQ7AoKqY0Q5wMt0u2wMnGsRcZEnCHlOeehceYt2IUzvs29Hn1f323JPdpCXgGoMDkbK2
Bw00O6jo5UtQsWPhCrCV2tvm48ozHi98us4bbOXA+/h7yzOAZZsoCq1xKTF/ITiQcO5KaX3cJjTM
mvyvG/YqcvzTBdwvaC/kzdFVR5+8oanSHzvGXcwRNTwwhXklgEA2/KK8Iq6I8NrdUS/GVY8pSOCz
x9oShXw88tp/SM27/CyXs0B8ZBN+oJ0DXYatEqk2U4Ri44wc/r4PxlwFopUi3H08Dk2U9AIT/DR2
ilA7HVDvcR2gXGCghHO9gaFFM0vdRA2+x34ceqfkonhmzxLKrx7h5Sr3Bw/OGJt5a/cQlVLKNREI
L4fHVb6OzxqOo6BBGNZd6+u1kWBrxyfDGsYwInx2H2X7H5ZDj1pDbI8x14S9J7VXVtsje4BQA0JJ
+2KIUt7FimqeVxsWPtaoFVt0/ZaayjgKIWHsT1Ncq2zT6g6AreGbxAHwjiZ9eCAnMMfuQuLgYtzO
aWNzYBtXmM1gSowNSYxwAZnYT9MHYybBh/a9sGKvJo/5feyC1b7YQUdvRajryd6hVWgneGPr4mln
ApyCIjMEYgZls1VqVMUL2wTBPT2IYiwhZA9tA3YXXq3yNIFsKTCu0K0vKsm5+JaLibbKwJ8Vbypd
lDpGHwdQrxwoEYjDoiEt/y7KwEUPw7il3tkLxeDsCEF+2GDC0WVCoPxby1ynr0ObDeHqyFcOS/hf
tZ6MILdNhE1UxTsAVJdrCiFDIqMoNnAfksvZB9clXA/zQVk6My7hiyLdqgy7mVPVkfdQlbEfM+MU
T19irrTX6cxplzRmiJYcUoCrW6vt9xoa4onQ/2Dp0eiL6Jlj/JSsRgbbIgKh3jh2Ln7XnEqINXqb
KkmoPt7284SsjPy+9Qj81SGMAgG2Af0DFSwqKVS0LzB7Dc+VPT7s8T0DVAb8ahl1D+MygZookfKY
fllKyzlkb7DIR4RoDubrWiabTBs4G3gh4dTbz9jI+x4e4LjGxBEwUYm+GI1OhXHHbYmPg0Y+kUWF
XSxyArXEdwHCIB781Bsmb146WBg+x6A01KnMYFtoO5UMRGQXqRtBYZzr9USa4PBFXQxsVLzIRpP7
WzpvQDtqEpNvUiI6wZnRaigNxZNzD20pYb64xi7tWSZZz6RXQEpkkLjlU50v7j46NO3aqZsuxR02
iFaEect2bTv5bnrd0CzJ/kqOQ3zVViRfQ9ISPKgS476eXB8mvqs5z7KlDayA0G+kL/Y/DzT45Bkw
t+Ukx2o410SChoPdedQMUxJSwV17Lsubjy24N23G2E6+nIo9mga93VNu8HOWNzawbnParCjVllKh
J5dJXaAPjlf/6JixWiM7wv0V1SJSSOw+wNvCR8Wj5naJR6Mu14qpwXMF8s8gjDQFYDHPMhLOulcV
aLAgCw0kXVIQvEbO9x+POpyySSeQgoxDla3yViiMeghVZMtw474pfYHIhnou+vdO8Fp9KoUrlX0n
uXsN+dvxfckdFhXtyYX21ADElxwbIu6C3g0sVBLB2qqi5Kmlcof5F/eMxJ9dVjKvjg+ADdqsPwfJ
u3YYEI5uZMQoAcUSdxUKdS1xbLAxcTYHaFG/1fAZw1D09VXF2dRjlCaehmDraktf9Xi+8y0Y+tH2
ZR0iBTYQYjB+N+bE4c45S2p1O1Wpj3PlSiEVToO8toHPWSpFsyc9GBmo8PBKMwMZ3nUBgwusHc44
sXgYkm5N2FLBbyFxHQT+dtiRYfT1Al25W4AMt9Ukhx1J376gdosvg+E/ujqIB4DH2yUEoUfniqGs
eNPSWKw/XtaNAraUSp7A7x9kZdbFXV5wHDBmjRWN1iLWYjkXyju367ZiEY+rJxwei0+3AN0Fh65s
JCyg3gPbMm/LJJmC0m00lyWGcSXr0D+ldQaRxxMejzxho04FyYGCyXyv99Wf1bRdel8t2a6zR280
SIuxB9fss2fcSdtfss1WpuztgRTOq59iv2tPpnBc6RLKnbOkATJ+4aeJcc5X6X/PEzf3b+LRfx01
+67zoYUfeh7Z+0PR0cHSVYd8WjlOzYCznjGTmVv0AV4Dt1M0I/Dc+sB+e8y7+Mvxvfzw+rEIs5Ab
dA8wxzdk4Q52BFoHsdbjbjY9POGUiI2GmVA8zlgeUZbqji1qI0bM5Pa7IIvJfM+Soq84ms8q5Wt0
OZwoLL3VwAQq2MsTMmXu0cIWy1qvlyyqgfUeqE+dMIkfE9w0YHER2Ca6fa8+kS+V+D7jsM+RVsUc
4NC/vCZbXVnvWaJvOMJUj9M9CFittnTUKwSaYmK3miHIvrGml+nG7Kw+n/Ev6g8RNGAZxbtPPc+S
4BgMC6wS6Z5c+rjfa+FyzDdPwxgPHnvSKFjk6cFejeGoUPhUUaT3hUtRYhAbRFtILET8zT604vRC
qPhhpld7KtqUKAhlJy6hXqjWgkVzryiU0BG4vlt+dBi1wPkhiHwpUIjmBLpUfkr5YOvKZmUCVNMN
MJPwoznwo4yFtcrNWjRT8tsjKS+bFNvAFwqjcyih1iD19wKUdrS68qwyXD2ewyGRoW2xVJypNj9K
GrsZ3FZierdaWkiXuZ/nreC8z/FjW8QiYMQ030q3KHzxbXr71qffpD6m51PTJz59PHTPMcUID2lC
QvAhSN80/8+Gmp8usXpQ1fS3M9F3nH5g8LypnPXlQ9EpaDrAH+w4bT6LD2h6aaPvzoThSDrZgHEZ
00jt9gQMqPoRfKc+8a5YfNQEQrBmwqg7YUNPe+MF2CJOIuL1UZShAS7U5kx/j5fyDZit5iYK2AZS
GV/nis5tes5H95BcI7F1LbgnN0O5usSLCLm+/nXqoctB2UrheGlhgFsHkGRiJsOXE8q6mpOiW0cA
fUxFhvN3OO4WO7ycO8ark2rSgoB0gpjbKpCl9AnA+6yhM+CBklCIvEHgWLZSLdvlodz7MMQeEx8t
Ferus8Lj4Xv5EJ/mzn6ke1OWgi65YUuMMpDLyE/MIbEhYGpKZIeEGOBOin9zNQK+a2292PJ9KYU+
XCf66XmpmcnANEsN6MiPzw6hq6IhIb0sfDf8yLirFe7pdRgauB7/eYCHV+OtKDrB1MkGgyy82UiY
eWeqB+mmrfdfUm4IS5TU6ts57M/73ZGFUAL9XhSHfOOxP9VIFSPYPh4fbyaXdzjoS4UKK8rYsb7r
bJl0GPa89DnTfM0x9F56jJwMZa4W0Xrgn+f20xcDc8KNxsdOicUGcn5TwXBDCX2eCuDKPFSkNVgY
TcJR9fz+KWmTWjuOC+I9HoVRRjOZhowjDCHwrCyPbVpbXWlVxqiljNaDsEb7S2Lrez9cAd2tgbCK
yTZ98OEZsMlPGws8+NHA0dfS9fQE+fUcAyXqcEsIL40U1ZJ78DO5XZVyEmCm6mbVkM1z2RiK9TI8
xQ6MoouhkcgCiE64BUO5udUeZ+oCaACQDbhiNt3eOvaiJNIBd6ve4o5RQJm3fm0JHDVwWgyEWePP
Atbtliyxlremu51C1VWOi8r9U5BHhc2qSpAYcY0slD7q38zu2rfY4w/oUFHEnva3XEhqyb61ueFl
j0qODbMhEHyb5Fz0+vDB/jDpv3lmk2WnmIPI0cb0MBA/dKLgFWmfV76sVNtrzcymhzcALUgIA1Sc
lBMYYUU7S1DMZIN4brEJTOxpvfRaV2omx+xl+gDUvxqaet7EVewTxmTUAU2svLuCY6t/aInz7agN
Vw==
`protect end_protected
