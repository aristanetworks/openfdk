--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
M8PIfetDhd6qove+lyGX+Gt9CqtNvjOsLHgxud0N3rGjG5pzdpJ+IXkiaaIbTSKqBZCAoZ59g0Fe
+r09KWfaDY4QgMn9sVUTzT9VhHFBh719vHKk+dzOKHr2dS8rKumEzTXQueeh57EaYpmUaiJ1Ntty
Mr2e5K/kImbsJnhhDQJMpvEgeteApo7c3A+s3VTo8oSxPxAa5zLL3zwFGA3w5Aob1Zn6i8U3UFfG
G/kmsY5rnKdFFBERegFb3ZPSpkz0c7NgjJj9ulb3oicMRQ6NmXYyoTEXOVW5wvvhgYeCpH+X+3eC
gHEqswmFqj00Ir0gSAoqOuaC8iWfAn6XlJRRKg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="koV+z9gJ6UkwrfeRyATv0mkPFfFIk1OekOpnJ+aFCng="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
jDuu2h5jMoui2k35gpxek0335ZU0SJX4pUFrWSwiyitqR9AHds5SudgTh3lknT21uPIrDA9Yrg0n
2F1ueiFJVVhC83zZhXrS1LdN9xAhLEB8CJ/fUzFftoqI2wce9uhUY8koSZCgTEtIa93mfk+H71GT
mrDGvxAH/pLyAu+cYW2RoMTgbAhbeO90cG8TW6wH54kjdPJGBRdopH9ZJMfU0D8OMjJrr4YvWqzR
HUhw0LGIYc8xHKRUEpxANnc2mV+KAK8N5EDPtHTMh9npOtPaHUybgnOa9lBy9va5wYbi0IXG1TH5
3xVYnNdgiQOcdCIbhMt0ZCt/gRjOqo/9jT4Okw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="rze+MSt4/xCmojoZOo4qMkTZ1UfC3OjxQd8p1qV+PQI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14800)
`protect data_block
pr86MQ1sGg6ijaboidq5IMU9sKb1r9CJXKDXDsATfR+4HlTOzJoN9QlSBf+O3Vv0kMBLxei3WPX0
eI1heyeCaWWR6y8pMRTtiJwUlo8qTxQhgV3+/gXr1kuatMqD8YVeTWccmyUYgdQeQj/gzl25ySE7
HC49DeK4JFwYtLV7AvFvzz9Xe0b5NF2j+rhhlr4njRBmT5puxUvLUcKex42NGjPKUsiV5Xt6bJwQ
7fGxYDaS/PRGZfaMdt5OBIGmykJ7YQD2PE2U0x+Z1EGz3AMckfzw5P9XMFR2dMDlYRNLEp+pqsWq
Z35TSFak+SHJ7lrdgmOSbqneK1RKEcDuDKDGrsSWPX8QPEVz33V8Sz+oAm1b5y14H8gtAbt2gVIq
lu0QA9pW8xtm/wcFJkqHMr522tth4yyGr7tZnGCeD2IVYgJvcL7QIa2uDG5CkxTHZRP+82wvPIrf
DRVlsEVxV8f1wjoxYcVQcg+Vd444SY2OFeTMDEwjmLRi/0/sU3Rk9Yl7VYA99XQB4UhbZp1wIqFO
OuQi0+buyTpD/SqkwxY1LV/Kphs1Z4LhhBwvLVz2kU1Tb/CVbBBXl8jkwxxHrv5uu7/6oBarCHkb
OPEy+p9Cq6sBRWFZhfTnQDAh9rDEiTeWiJix8ekQdBTTlMXqH4GVQWBZ6b5J0ja/R4i2NMZj2pxY
Bffl9U/NHoKiEE/kOvZ+wtjDRZdYbKcrZFeRD6/UvIT22M/QUyfaNUfEy1FfDZedlCYS2Ileg9dM
x75dbc1Gmf8IMjVpCjDtz6j8T3kWsjB6m5k+Rmqcrb+4Y1QonMSKGGJu/qV4kLRm9oukfE1P4cjP
A3rqCTkZUgkP2WVfWp27ggt4a+GI7/XxsjagQXEALx+iCmowF4Pu4MOrb9vxg8MjyDbIq+oa9leh
jVDuuHpsfDhZmjdi27UaSqPqIM9sRNoAmkViL6w1t6N/l7EM6ic5pVwpxxIP2qCL0L0GYEATmOd0
FWGUhoXCoIKPG5XXVaBZw0fzPoR/MnHI2O9FKSBeddmXAj2yUhLEtjXJyyqeKFg9l38C6+mzDjP6
+JuU+6fpqJTYraaH5yRDQM/wgpqfKUvwODi890vTQZwNaypnI2dfU+fq7JBgDNy9pz6QIBNmZBMc
BgEFhQMarXFtZxeCQhVLOyugWcK8mKEy7LjJx3iLEum4YjJtfr4kbZoeLNMcFwJ85YeZNdErqhJj
gr2guMIcT6z641L8FvNhGD9Bi7btTrn6ROTmhcrV6jN6XjPSJXWIup2VqyMreyHvO8njwlM86BYD
QmjCKb0LrvnmHfV1/jw5x57TFR7kMe3N7+t4RTaXmCUYCA7wKFkpWBCwzgD1Nb4CoSdpp96CDZU8
lnEvCFrk+akAYmNZY8V2URLaE/1AomyUAG/wpjYEKaB8DaYYyg29dEgX8j+e7c6VA8XrQmmWsGBI
zgjcwP+u1bM4wyHl145bSvMU4IjVf/SWKPC2uKju3VjP/T2aMAHdlDVS4+SZAqZeUPFwLZF5Zq+s
Nzj/lfp95fX+1bzwUxfS+VJVXevqShXonGtYIIuqXOe2TXhuHolu3i34uC4WhVfJBB0BDuCe2VJY
P25UTEw4594VcJk0LrnP35G3P9xnKg6DB9BgmrtZLlURs7HqTOEV3p6BPSScbfKcpfAQfxpWGJDr
EPbng8lVyCmAoRP7E7OcyVP2Ur7vAArOL7vxwYHAP2SVEtGvNTjCXMLM0plD/tRhSdkiB5galKkL
HkRliuC0hLm7GrHFJ16PvPEKytIlKN5ftTHsgh/X+q5RHhWuFwm+wa+O+QmN6hKYI/ZSk7Hm0xcz
eJXKuScTss970c3JX7J/Yly9jN6kLGznHCzTZ30/IS8Mvx1wCnw/4d/hOmMtdwipF/g4UM2wpCal
dBvZ3XqsNe9LMpelflp/iPBJBnk30p+oGkx55TOIp6vTSWIN0KCbTGs4pKIWElnIpGDqif2cAFzX
4MYt8EgxP43gfaQNHJ3BIC5+jRUYVJRjsvGfjlNc8dBtvzKQcQvldBHYVfjUaeBFTc2mQw+zFEx+
KLHgisMhumHjcdHGK/E7S3bGTydLyjiO9NF8B7mo1TYCQGE5q46ELelraqpQzIaH9Mp2KngrgT94
Kq6H7LInDPM3CkU7L8kuzPj7LijOSUqp5x3Sj2usYud2mEWt8h9yh1dmqn1rCP6s8t7Qh6JorX2c
6SF0Rmf4wWHBt8GBswYosFXzX2PF6syPaFfMB8Y4EFEo78zWf4hMtSCeuKZPgjGQrW2YOfTyIi/H
Cz6/Ur/tEppkApkjJpEiDX4eH5dGaLYfL+xIVMbxuRxn4ru5+7a8qAEFXOnslFAX043ib3j1EcON
zBWHjD1HDaPWli7VhjXCw5JTUL9dYtxh0zqWNtCjLSKyWvObxCIsD0soRufR+mXGMPcGSpPQnzVc
40dvdEep4PrQD/eRpoWjCGdBb4U3YD/NaKWx3PT1/0mGUBe3ByXqLdAqFsTJJRsneh9KUa8OAJrf
yNSROzE0hdSe3BpX/BTrnKBGIkeAUNBRMOXMqB74f6U+vaqnF7DA8g+DrXiy0h14t1lKPKScfsOC
nPJ4EfM3vZ6w2w4XgWT2HFTWehIkn2W3xK8gIlL+YLp7xi/4J076JjW9pi4qNa0+uzYLzcJHD0mU
8AYWo2PIlwppSx1CQvF3BknmRkgVbEMzmj6VwJIuDnXxfnVENuzoYUc0n+MhsAu06CFEUjx3LTkm
ackdfiPJxm5T5IjEWGPTlDZOeJJL+qSiddbwCHsrPr4SjkYs0yyduLlmiTOdWPen7dwA+p8YksHV
eAxNUTfRdSHbhLs7tawEK/GfK8lZ9xOkWHlwwRsLWzD1wsKoxrvfC0Suu0WqWOisWv69w82pdJYW
KStzcalyg23QxlGz/+CYH6E/D67V5lkppuo06PGNTJS7Nt519CFF5ES0omX9o4y0q11VZQDCzZpw
UZXK+CkHNPf9MOicP12MmwF8C0zjgtDJFeQOEySv+XHCDZ+VfdVGL3Yw73uxanwmHKVaqtPUDNc3
Gr5iAyn+b9V8EQxHUx/Zi2HG6Nj9vZEow1i95pDMQSKHrBLRkdLK0I7N3gc33jfhFDLceDFvM9qD
bQ6p4dis5hVNN3Ndt/fBCl1hk25Uk64DfHZ622+OZu2m8E7rVNn94mobDsbk051bT8w8QIIZr7Un
4SJavXUytfRzqCSmAP++7G+oe1Q4x2bjCzuDHj/gVZwlqO4hcWcOk49Q/eoSMelU1ZII6Ey1yYTW
GWM16YxqLVmRoszTZguXXuigYBdZ/0t42pv+nwJtNicvJ9oZnqSKJi3ZHKtl86OMDH7RlHNA702V
ti14u8ee9g3m6VdvTmj7B8GXq2pBW4cNGtdfVHT8v2eX0LvGNFnjGzm1NQQotjw9VGV5S8OVpmIO
t5o4z70lBjibbnfeI8MRavTQ+aTr9BOz1J6joYDfwvBWDYGuEzd+5XmKb+VaC5cgI5MUf4BVe2dI
457H0jnzhWD4AnRqMEQ92JWdsaBlUZH2Hu+bQQBj/lFoXr7zubphxU+yHHogpiOhyVfwcDCELe8y
vbWFhtkj2x/AjLWWEMJfC4mNvp3dgp+gNmmOQRNP1bGNAhD2cHMy4YByEUe0uh8b4N8g+H5tkKR4
6TTkMSyILpDUQUGKOUgPa0d4qMl6015g7XXasdZrHi/99mizl22bXzkXJ6/LKZBFvxoIe6sf+duE
7zGK8Um1E5DA2vphZvfVS5nlnU9Jgq2UF+X4/Z5bawdHlYygzqD6SrCS5eXebX1x3WrLJ9Zfc1Fb
WzMUZkf3Z9lXztLl/CRdxvfm+991+GMecr75y59MrwY5CaMr22sfg6tyhp/RQTLVMajkAv68/De3
c08ADFMnMOJNbHZfJQxfpz7KOSP1oHc4pqKjgMCrnZkNvFEmXYuYBbjCp9EhymdC5UgefyECZdOY
or9L3dowFTUzVFlPRqgrO5NYhxEdPtYjgVFG/XzRxNjGaF2oU8tO/PHUtRd/HYoEpPof8CPNDJOj
eEIUxZvOofPl05lKHJNTahP3BSGRiJiJu44PRSkigcM9dLUfGMNgGc1yjsNBeMDmcSgneIPHgkU8
9TkAcoZ8sZWvSMOE5zmFCQCVqzbLnIOrnKWrqjxgPZkYdlI/UK0RJfpBjqHWtHotOU/QcYAxAf/Q
kRh+7v1FvKpu4ndpFM7EZ7GH+JRYAcdGfs3te9oCOsue+I9hF8tC/qnG4caWTqZKMczZCK4Q49M0
fse7oVEh4PHbEdYcBvmjgk8dubWPKbLyeckJwgJ8cDdWXrH9aXfXvt8ovHAUrC6s1NjrnLHq6yZ4
99lqJFJqVZ32rOfev05Pk01DVupJ9Z70plfcI5CHConQyKm7VKyu7sOmQli+u8CuwixR5XGoPHXG
dcJFzhW7iukpQ7WqkorZNOevG/e0fEUe0IBUQk7xDG599GXJEpWb8GeDLQ3jPHI+6aajIS1kFV0H
/zJCK7xL+PNuYNRyIlhuEY9q9K2tdaNAsx97F7WHNy9ri057pi/zkAbrV9xMMkh69fDB9sfUIQ7C
mN0JJyNloACmumudf/dLizC/yq3nNNsiNdVlIv5xQuAu4PxyI7T12MFYTMoQx1zpF1QJASAaiCfC
XyMMFriB2qSj5bhtLzuu+EH7XIo5kPDSTdMrXoTHzTmcvb1SkBY3pf6UPhnTx7G1l+iS8OPKpI+q
SUCrHbhGILi8uk5JEpGPSxfcRO0pQoCbVWjkdQ0TFk2vUy1/RM1sJT48jwo1McMI9YnpeLIZcxmo
g+ce9clRd9qa9dz078j9mYyghiTq4uiD7EA4HpEXRYbVqHdLzTvtl/hdwlNGIUCKu5VcUY0iQvia
KEgy4kFArtZui21be/2Vnu8Rwb3CAr7u82+g0zdKk0Fqz1wqQ6BJ81Jo31lJ2DSyjY7JR88IHH2+
aysYb7H2oAdaG2Ih2gI2h/tqRo8/2hMQpnp1vzIjDYRCkQlEyjSGIZktJBOOw03Xu0QTzgXjE+dR
WTxPWZ1KHreuIsCL2deKTV0AM8OfY8J8af0Zdubw7beqGm/d155uiwNB0RhefhGjnx3xANpsi0a8
B8lRc+a/S+4cUcnHDtLwcNlPh7wB2NZ63AaDGlpCfZXSkh1ovLLti7uvskY/aHGFWiENp64a072J
oPMDaJ1KgqXwctWkx70SLiiwZWhgwyuPj0XCECDO2LD79Wha+ytwIYxOt3stLOg8u/adNns2QJeo
IBkBgb4U8T/wz/ICmTFO69W3+mfoh2ogzM36ISBPYwCDkF+rJ07TdsWIH2kA+valNZNZ05F99bHp
s1rT8gXwwnxwJXOKyDJdAlhOyrcku4JiURqd9UVvVLBHW//2gA6fn+wqReM1p8TrSuBWtV2LlXbD
VTh/9s8VlwaierDmydCASdeLiLsf/mvZMWyjS2vN/VDoFtuxXhwaX0dJ+MyCCMN0f/quMv4pojqe
U7HhtxU5pSwsVEsk8OZzgN1w9qoudrKhY/riTB5W7Jjx/1lCVaBpbaYJBPWr19cJrDMDAZB0EflB
UlCImErbR1Rysc2n1edMGorsJEcbbchfACDkRVQWIOQieXGTrSEvXGjgUMfO4fXUTVt4HobNlcyN
8fmsPhVeBFYzP4T11fdGP6oMLBIcgQdkrfs4VZ9VUIIxGJxqKA6QqD8PoqzZS2rQg53JufLdTahN
RNqclSaWWs0HU5C0YbJ5BVm4XVqjdISPit4mynpryJWoKFpczRJL8My/t4siu9VpbWJB/9Ajt46X
c5QWCzUZzcyvbGpK9pOpRvp6uQ9HwBVdBr0WSViwQPk95KXhXbIq6ax0SiXfXiaPg2KSAeXbs5Qj
qZcPs3eke4YeclCO8g+t63cLVFSTAb8IDALQd9WA5OVT+JKyBorPimi6QOP0WnLKxtGPktVn/JPP
hjGp+4sSB98Dz0Q9hKR8zo8gicDssBuWsjNcm67hrqiuxyGuB0HSnnMoss70uhn+k+XfNuiaMj3b
Y9uCepwclZ7goaYj8cDitQrjmrAuJ8cb5Z8eAYbE/2kDVLnKMNY7PzcXdnIQDs5RZHWxg20i0/wj
OihJk1mGLbIqCnSnaYiNWfqwGGz00CjKZf2jGigrLRMVWAwXApVLZURqt+loCfNt6dvoGG4nktwX
ds1at+QsvUYIFer3FRCjJuA8JYOFe6eCA76lL6LRpKVzTdbbAW9NR1j1kBZSUo4sycdCT/KhngbK
J2l4H/nj4nLMtPwUduJSKxP5mgYAR6941jQ7sPIVs4RlqWIbijE/IKzCDfhZReomTqCbCMlL90Lj
gUsbVSifLOB1xq4k/2UKvP/Y7Q3fXD9z6fWcxd6WHAo1TAiIxNOwRoHj948tb6drhR4achYtmLau
miboZzS8u/8kfX6HFuPfjXQatKyXfhVoZ6HqbFQL+McXcefO/vy9KKETV9t4LtI9qvN39NJDMJjR
nEZGOe1UChKMv5ihV5iUYqAtOyT1vCP0eWogdL785z9WUKNoXtPwyOcQYBnhm+JNuRrUrJJjqVL4
S/RmOyGLnXtKEI08zDuzSfK2QTRYcqF5ylidGi6FmAJsbO4GgNmcVKUoVDTM/d0z7eMeFII9xP1S
sdDrsJyxLgS0Xw+Rv5HEz5LOmND2DwoJTDi3TllcB+qs/fglm4sl6za7/xqRcPq/1apVRCWXLQpp
kt1EyndkyVByDWWgGWeO/kksqDiH+ZeoaUTKJO/qR2MHj7aGmMcK/Rhhmn8QjUItv/dwaovqjuul
TldnhdgsOXECHXenUlZqd86tAScnMW1ceVx+hK59eapekapVgkmcEAFMyokHgpPG9Tl0sqE77CjQ
67/7yuXi8Jj9s/Ve7/sx5zD9jdTUULiSNc7VW6UjRwpVxIn1dsZjTX3zc5+q5YhF6nbLk9A0/50e
WJx8udKjLSqDHeH9rsJUWmUDMbAfgsKbfB6aRKIIfur0yD25/Ecp3UvlG39qc/wN55/8pboWUemx
oaLaQ3xYtq/IUtC6xAEk0PpuSU+9Tm5WT/AHgo+zQ36b5pXmpJgd5uB/+nyhWqtuI+g5z6rsjIQV
3cKlNMV9VuPO0ASe5f0bzYUosDNbRFyNqU9eDM5W8uHSQrhmIZHgwdCDy77AkMJ8GH073bx918gL
mbdCaY/X/QGcj7UN+Q9v7rFhnxxA5tksrSWQY6oM3uh1P+FQLM7QyaDKmdC8mRLvpECXTFTDuT9z
e2tpo1RvuS3TtHLjIw6XwFkPciSSy4pz1+7mxeIh3A6fB08i4mmhvA1MRFDb0YpFfHvi4z2j9NxX
lkzihCIgqxOIiWvfOSjjnrFDtkrEzotNsV4s6TcjtnSc92MmPWoDmbt/cgLmB+oKuqwZWYlCMjvx
gnVNBlxr3wQcvLzM/6JJNYPaAFkZU5iPslheYD307cqlq+nimAoEsIcUFqkjRp6/sERTSnRfFCsa
Qu2EvGabxKznvhQc1CP0zaI4PBaet9rruy1NuVf2TJ70vzaqCRHHImil8OyTD9GXRMlDjIMS0WQx
uOJeDL6c5PN/I239MNN/2TJiWkwGfxkfxOdvccbDzuGjMKgW1e95JoEHCJ+Nlm+sOpys11M0Xk+R
ZApyfM60vhTtScgU6wjlBhow8EYHZ+QgZ0jPIR1WIngRCL3WzeGwP37a0WfordZc4GYYgaPqdCN1
pJtokiEQCdj6RQRbJ0vHkRMlsu/I3A2sIhJLs1Zw9xKeFW69PjebGUUC67gBUNpLfhYXxvien6UL
N5KMULZOeGM/0IV4pLfn1lrnIOtOQhqaYRt4r2CXjTw/XE5CA+RKfhwQDGiXkyEoKYiQaJ3YpPr7
znkxPSE3eCVuhv1Hj0nlexGA+mD+s0tJTL4djEp/vatcOzopPY8/lY9C/2Z2jB3egbIXW3One1zf
1BJm9dNCslfVmBuCjGw7QKV4iwIVbhSEDibUrUBCYMVNeeV7dL2d+F+JFQL9n45AYKzgOSR1BQQM
CRo0jDnEO3B3ytXTZFc24zjlPhD5oG8NEI9ra3ajrgfp4P5hggXaCarimXzppXBuwUU9dufYSbq6
LkmDj6MDDPCc52ho690xReZsNOy+1CV9y5o/U0/Ic+2Ca400xz5RJ7ubU9nFRov3S4tjyfhSNgJO
RA1t6Yk8A+t+4e7fpb49KeugIGfxSSwKaVr3fPdFTBvptoeeLwNFcngwuj9zSKvFzsgaWuIZK1i3
rqo23KgqhKQG/jxMMpqBj8RNosH9yeQetwvAw8kRy3U7JTSXEuGgMlpnwTd8uqttFuHkqomSwuNU
n9tFATZHsBtAo2mU4whmpXIkIxGBO14ssGrPqMrXzjBFcLruAdfjHoHsIDJazATOjDzm1wlxj7IV
RMeqqO4GUQMWgLTwCZn9ibodF8pD7sK7Uz00IjFsN6QBp81ByNm3MHwqUGi09m5V5uUJVhluJM5p
rcdhkeEqWYeCOzSKGKno7YbOIWVPrZageAO6uh8TuiYhY49AgSvzuUpIyZUa+OvXCHhHQmPxUyM8
HtgGcIHxcQjGq0smC41XqNIm/Z6IiaZvNkq/MuiBmVkaoP4oJvyCDnXOo3oROjlJY6r9Sv7tX7Af
mydCootoyyNROs2ZYHPLj24rOxWTOocD4jZCUAetCSRcqccGaVduOskciGMnBVHQaq+uKFZyJ3wK
aY7SUut+Yy++dlTErxrxmkAktWPuJ4vaQNMvnZAcsmKi4LuSqpLlr2SxRPUlWuWW6XU3lkPacIES
F5waVwB4XOWV07PHKwhajpI8peCc9DM5n7mcB+MibAj/dRLnKxyYJuziB7s7NUcN5IVaM9oI/Txf
vVCYosI2LfAVv8HvdmzpwgKtk5PGZ21d7cHqZ+j4I6j4iSfqX1Auriy5LSLxDilWV0vvVtX6VZKY
Y/HcnXNpLcJV7LAQy1LlqAftyYIPxREis4/goyVtPn4OuZhdDBlxit8xPkiluZ/Uo4v44bro+Nja
QQo/aHcZWv66mly2yC+noV61wOwsJuIQFv3DuWT6QJpZBA+Nd34mhyibHV5dfFKadFonsDpXTcLf
r4GQ50xck55iUMP0OO3nySHX47ZxUl6OA9KMwRLTdDoB+2BvScWw5jsXUP7bUnPhWKd9Vy1mNlP2
3C+ES8YiUg8NYU3w4GkSxrxoJJLzMhhPXS33s0jKcoKyu3OIOwtH8/nyltM4utPYFEvmo//hzGfz
hTGbZ9UqYUGMIRp1iEtRn54Dt99YzYD74uBMsKVtgg58nuyZzkBq5zTnCn7KGd/bYzS1AWVzkXA2
ApTGLedjoqJbmITt+Ev4idwTRUf9opL85SiJxV4SPpI4OyvbbEc+IaljLuIPm2fK8JehHR/29Edg
wwPwFcAQ66LHKlkDNO1sHWhuO/mNcvjSqfUC0rZXzuMW5PuvER/BLvv3ULjBR3r1Q78YfBPIm3iW
/v0MrDdDiq4vuAQdPlijeRRPvE78VBN9AZqJwhSFgdbBmU0CnE45llwlVQbJp0soKdowHUnryuDp
SXcI2DgpmN2s/z9SVJdrJWg5WhwEIUqoFBU/cUZ3RWlkQY+vSqXxJn9pk09D3uGVe4YT/HfSAijn
B/SmzyBJ3jeNngDEMy5vVm2s89xmxpXXSwTBpKYnYgTFLgLYFP7sf4WFGjIRFgR2XU3MBwvdqnA8
BJbgW+5k6W50k2RHKP3hzffv0eh3xmg0ZbBtw1S2XNDMkfj020l83BOgYBmffqZTDKKJXzhQH8zi
Ro5hQzlft5utqKj0GBbZv8mM5al3mK0Cm3szBe7QdrN8Y8OudiWwGXzXTT1TraPHqXxzYByg35zd
VdUWnE+OgCDW/aNohgcY7mMoGqEUuzlHqcDWa6K8wp44hdLXUKhewSza0lAYJRuU12wUxWxrhxR1
/GJupfxBiquFJKLolTxKvlEP4MDddcBxseDqBvRXY7RzZuVQ2AnpXTlE2/zCToPcBnFhOSllpFGT
m3z8/yPrqkLjAbJyvXn3/L9HD6MgwOHc5X15rHaSjcII507BKVL+Hu2bV3Pybf995cDOP0DdQx/D
r7q7B6cMIk5rHN/osJYFBJ8vowW0q4hT92wYNrmZYJ+pbsfAwowzS3gEhutyZ00D/r4l9kJIqy2b
SGL1X1CbHU57zHrVOYGAhbnqSIUBfovdYNLAn8Vom+Ld8xsQs/9ipE9lvdaaYtUq1C4DfAt7yQU+
id5UmuPu32+3BttM/pa9PB+YkUCYGxUr4kFIc5CxUuBjnvg5kwVZbRGmiyIeASVyfLvA+VgTXBzZ
aznfLoEXkCkcrKLf+LmQnslvJ+vCTWNZJek5cW/bygaCt5L4vqionD7tHcMX5y9MX1+rS3PIFpCg
akSAq1qDhraPMiCWSh2jE5TLRTakQ/0Gq/FQVVUSfCwWGqvQc11+AGjZJWmE6x5jOO5Mn9iSU7gR
7xBSkfCbsZmSmfMhFt6E6sAyufDi75KoIjERsfLIu4bIPOAmARA1yK6B7jirfk8g74iw7Fy9HZLF
gre0EmSAJ3benT5E2Y6r3HEfSsslfyq+W0PyfVaddMPSWRbB+aJaJdcNYCPmfzmU4qWhui+yAgxJ
qSYKemiV5sNN3NIEle++7jDUGNVH1/LVFT5D1+vQX6+dagkttlG9NzMPfusvr1L+aP12QYfUNuW2
9qW7y7iPNHUso5flGEYpTYwK6xRSHvfXFrExz40Do9mukI1KzjLYz87H2DKehRd2q/CbuA8mGCBJ
fFkQNJR+pSCiO3AjF1FITFmR2Vz1lHGPYBgiNyEvMNzb6YVwi6GxFNZZ/aYkGfC9Zj9OnHohdt4m
W7Zy2J7QRkp5jiLsuyUBfm20JkmS9xdY4lAaMRWgz0FAIABeyJDXvzjg1wdvhFpk4tV6rIzs5W7c
oAkEYwusAqglEDoz8kbwSvhpWeOnVDa7/i9o8n2ULqzlNFf4FYkPq/wMusjbor11NwjUglPiWnG3
Db8fLu1gEUk69NK/eHjUi4NLIY36EBstyYmpQqIoR1s6Y6LCgJaHUFSAKXPtapjRhUWFxZb7BkST
4Giic09M87IM/sfytRM03Np+GvV2DU039rnbFKqzo0zz11kI92rl5xm5gptFmgS6jJbmOOH5fi5A
PLfM9F9vrVG1VnUuKVNvYG0TsRvuXSDeGHdmIszNbeKVvf6Aw7SSq6KzklAdXI0aQ3ZRIRew7LAy
CoLBVL9C+MIi5jTEAfDDx3NlE/vcVEgxRYz4O+RERjXNs2O4fa3BYgnju5hnn+Tl8ZsIbFkCiiHS
uzk2raafQVZjAitejKQ/PPN52ni+miSt34RBcAud9PoZfQhIIjM2qupD6ChBQr9iQH0nVZqbksC7
igAY2etBy+zbNnR895U12MCyDRHl1TKoaaQ7hLyQRnCfsknTRo0AtsLcglpwl5R3UR+9ysTJUIyx
ujMS4rvzseg9W2OiR4OFNm3o9XRoCbrsnRWW7w/ODVtqLpqtSnFgpMdcciTtrGROK1653TdRhEMi
mkkiB2ooe0L7fmYWwk68wDR0+86rraMwTxMdApBPJLb6ap4izWOSnBsNsbG7uoc2ujGnfYCN6or3
0MovZ5Ymai/ORzr28K0KKIPhTQaKwOEDwYr6hKVhHoybt2ICeBYOcLR8bsgf4gkdt+YShRX0F1et
8aS9gd7a/lvkxysOlkL7D8sp65SxSofptQgEZneDlVrWq/F0Z5g2zi06LUEpGQZZf0saVgUlnBsj
imfX7Fp650j1b5R95XewtreiBH8RFhkioOfO4OXtdeEZeSZk6sic+4GKUvdEsysV9SiJzIJglyge
eRSxMWem/+sFXjgZa0fzneYa+5MB2RPeb37mqzINyIkTZ9ashV7V8alcUiICZIYawXvY1aJAAPGX
rvWv+qAeuNHFbSQeSCDe0Lh5M7xiRCajRyhPbrK8XW9JB6kEp3RYGPdjEOhHID/ToNdto/HxOsYb
QxYeaWpiSs9GpmGGonV7SSYKB1XOOXwPMS1YDguRj8B57ZtM3Oh3csztaHVALv4GyidVO9kNPrPT
81TVopvE7VqEy6h5nXLaUYtqNymrS4Rg4if2VsvAf2gKHbiMh7A8tzBgyq1JxpYGFKS+lZ0TBjHW
QUhlsbYhWqFGFDk241uAVM2bDpGUVIVSojm4UZay5BcZZH62iTtmoXN6HFIzgK0gKjjaeFzrvmco
U/GzyMRzv0l5Rbi6PCDele3ZJJ+OFq5x4xnqgBKODhDFkdzZYDJiBV/pJSDSp95uYvwPQNWdn92w
oTq1Lq1s+qQROQWN0y3GS/MewGMIduAtUgrNolFBqMNZ5O9VRecL4vgjbPY+0Ys170P7Ysno4XBB
1EnywiYdFXH577tdWy2lrfzevPIJZ3vkariY/HAPE5+0Yv0rxkbsuM/RTqw3Dk7QJUDC0JjxOQxg
qomJlrEZbOP1+12BF1MaxdPld1kaRqlHgxjHIJ2QVz9vufjvXduZyfpyjuyvIjXUM2VO88AHvCes
peJHpJFvoTVexn8r2yRAax1Q/spBfX0i1CsEj94PJhPVvT3etPInytqwZ46npzC9WF41irH4n+UH
gJY1dD103zJota91b09g4Bn92Qyq+iw2nSLsynLEem/L49NhBfN6zAsURQQnGMEHQrBBwkOd+CTp
wofI8gxO188S1W1VGJehC5lj1vE9EtOmTJwYitidczZLD1iipTFs03BqQxInx/rajqlVMV1ohVqg
DzFAdVt4zhnw98NSvk9sH8ZsOiIpeocsArWdpocpvHzp1XQ0umHclfHUOux7vis3vxHp1FP4Tznk
7PwkWejx1trTVbcUCEYKwEZqvLxUHqXuq229V3mBcAiZF3bafJkfan+1/u3VXa4FAIvQ0qaVVGRO
kP+J3KoIykyStJRTtXYPsOXaqbVztPiLojmTjdmzlei8lhoX9LizjQS/kMV+5KtGlt82epZj8y76
clXhe0mjNeXnMkR7u9psg/r3HPgif+Od6LZWeye7a89OkR5NWcb+vowk4z+m49rTJ7sZz+1uxmS5
9qqepcuZRL3hTvMhgyAAUTg7vcGzes1QV7l6agABG3+6i9sMGSDXYM0em3MfMIIXbLz1KkG8V8s9
4hi4XvwcqhFe0NmhKHiranVY0ae9iKJJASZ0OqC6lIuxMb5EvlsR26Kt8XDchNqfNDLUf1meX9pD
1rirfQy/OkjgyMS1r0IP6+QHK8X0fyw7SrWpGyRotzokzGAl4Z+qdrfrT3Xcy4eOuaBVSsW+CHhB
V14YHYq5+FDqyUjnTvLN32TKPTfjRLK7902yImUFMuZ7MY38H+nNaz+QiJCJfyPVO/3DsTBxKEy4
RdEGohlgrU3w8zLbqmRyBeER5x0eqeEbBPmQxBkpaE5YcU6Vr1dPwgVkzSqBO/MWtTSF6m0VCNFi
DEcpEEhT2CRkCLPvDHr0ioLy7XuJF1AZzwPn50UrDeIHFFDzSIiUEx279sgZgc8R4KbIz5iYhzmW
S+6VvYFRFV4Rn+RA7nA3Jgp1SVuLJ8Dl9sIL9NWeGm4TIKk+6ZoTN/A2Oj1MDLXY9e1aVjrH8Dpu
K++rk6Zp4rasFiog9HezWQU5ijB0r3bRUjKC7BYbKzoEWTF61eNeCy9PaxjpBABivmPe7EbfQJmt
yoZiCG4hBI5jT9RL1ziVjusxCgjZl71tilsYHoEv7bMPuhM1atDfXoQ6DqPdA/Asmsz3plWwB0k4
VWYP71mxhl+PpE+CdI06DFZjsaxNvS+WK3YU8p7j0cZgHSBsK0OoKZmlEicFaM7UmZD5nUlGeYCm
vPpT+GnB8gFuHzIb2kYU7zZwRbtJWT7iMWEQrOdCDd2mkYQ33RAy76XgZRvYRNwCupY9jF7yZ44w
cUQd26aI1M5W36xYJxmx1HG19wPac/emHuqO73I/ECLXPAIqSfkvZ/iPYZkF63x/gSrs/Jpd2tOW
6DfXrI3eBoqIPdAddfgNm4v+h1wcimiyMFG8cxjmVh/TcTKExVRTrQPZxV2cyA41kDWwTJeoL0Gd
cWS1X0Kjjp3HizDG61esP04p+b7T1IRwbTiJkLYnCrDsLf3WW4u33sbKgBgRxUhWRUHuYyQg5gK4
PR9wyhe/k5FUH/1fWhB7DvzzDetkQ8QvX4eNWd521BxYapLVQ4RT+Wi1JmRNDWioXjVQKppE+20r
APGy7MvJZk7kF1iWi68JiVllF8ymzG/iZ/8GR/VPvSDoI0gTHkBZ2G9apbIMj7IHDd0jBXeT4LQH
j1WpEC1lfwrsuHbFfz2v928Yl6zk0qPCNJuDRMRqFRI5Y0OuAIU9uzxbenETS2E71Hv54dhymXzY
w6X+zWc6Qmg/lkxzmgFgxDb6UPMowNIeRkpFVu5vBzGPFhYVzqe4vB/y4EKGLbmzcMsNoHePQeFD
T+ojRC0ml8i5deiFN24LnHKbs4UEBVlO7UECCZ1ZpumMg7bK5mp9A5grnUL7BgryiAn2TbK1VEDK
IvF7dcL1oFwKVyq65NhIIIC/7M9OE25uzxFZW2S0uc1KqCuOMa3xDKG+S/J+Ql0Z3c8yzsajTS0d
Wvc5gi0cQ/wtoK7Bs7lJVk/lJ9UoMuDY7Q9AOV5/DTXsDcFWCVi3YW48/CgMx/U9iC/kikF2fZHv
3waG6sK1+70IEOIrTkWyRA/2ePQoY4vzEouw+NboCWXcX1f3Kguyelp4aDQSL8OLVgVaW7Lk+HlC
k4XhfU1xdtjp/4km60ffsYKYCOwpHVi5Hbz9cjDJPombfoJfTFSa2EN6a4dO3m3oYaMOchZMZ7K3
4joUPL6YT5EVwM/Ln2ctvdqhUBSpnmGCIoJFvNWxgFisV2eDYkE+rVbwYhKJZHCoizH1R2hWK5mV
MXPE+FMJTh4lwKzZM+YWcNtKfWsSTDLS74+pjqZBUmrTigoeCh9wsKgxoYZCkDAOZRXfBE374oJ1
TlMb7aAV/RChZZ2DSzmdKQA88d6H9POO4DiVZ8JmORW2jFCMweCHTwxz0JAt7f9B6yEDhhPG5twM
Qp4PIvVE2F8NfC8pENA2QznR7yxGmMV3M0BX1Z9miEjPP+LggpaUXG6vQEuMcyX/HJxKRx3RsQ2m
oERJvxsg3HZbtp9SH1a3Rjzc2m8otz6hKB8hNAKiTzafGKcr50wm53WAxlaLfcCUeE/dBjtObMpC
G9aOe7pPDb5quCu/lP0ymys5zGCw9m0s2uDspJ6alDunqCoXpnywbyQVLNW2DEk63ErEXrMM2ZYH
1bpBg2MxoJ8UslixQi83NU8brLGG3DYTYwyHQfTSZ9wYgo1Xl8NvvlK/oXDisZLRQ+Z7/JVFCdmA
LF4+nRPEqahRRKcobdOeLw4tF4jzZMfSZKR7s9QQGsxCUh+OF0gs0QH4fJ26sAy5Q7JJC+6wou1k
0+1OYekjZF4Lspc5uObC/+HrqoQPDEvOq3EUPQF/58m5y3QHou6+jhZ0jN88dJ/qAt8CQx4es/qY
Oht8yE56Lr6BUGj4BBMtHNS9wr6RftuDJjevLSWzI9cCgoliYlOySdbL3s7AFM9uuiXGh5nZiz6A
gjI6mXHb9MLUFXAVntpHgh1LfFtKJkxFdKaNgXisbqrUOPrburflClIHsXmYmZ82RspBYS99fDpf
rYb9HTmnmcJTaOmbnAyD+GOfR/5IOLfsfjORRvrUxYeu8TTIjWtCyW88CIpoTGoWGnuRJ2n1fJ3K
7pMgHZNzIQT9J4YWtz/7/1NBpRbqv7xixzo9wWw8fpG4Lgn3aith1bSFMHFiwjgonDsy5MiBOa3j
rYZHp8twTgcUtWcCkeKC9fBdWUlwvqjuGKBmjhbNoWo52XsEa83p9GuELQZ4YMSkKJz/BxG6IFPl
GeMxy7V23Uh/4meLEfHAAxlkrMK/ZYPfERsi5aEyPALibQu8RNEm8ppJ2oMWUiFh92jwBF8C+dQZ
9N9cITvFT+6KFhtlA7XKM3gexp2wcuNX8C+PMZfXOmATk/egNCt0F4wvJMVSVjC7mijqr7IzcrKK
68+JP9PMGBpI9du8Dgy9XttGrz4tukknyqy/5sjxF6uHsdvW4wxrgxPemUjM/nUlRyt2cO5hL6YP
6Vow5/oL+l9uXwMFFtZEC4G4choB4TQpiBunRCEhPKg4AguPgAqU84ryTZ93RCzPy+eNwe3n+4y9
oR12uaCb4JBfti3+ktxhG+crXERsrlvGlGl46lOytManZxAkmeXmwgoSHd4J3UUgOmy/al+E9BTF
qaKQgFltO2VdZM0RfyaVE95BmKTFFt3VH7seWeRThs7oD/dXBCO8jP82xiA6RiQO3oHQlScZuRQE
MnDnaphHYf2s7A63KpwfO8XiqiV7LNGHovF/a31cLv1IT6yfz9/zbpI/CIR3meuOrv0gAnKcZX5d
XuRp8Q+mYKW5i7Y3gxNDOoRQj7bed/PDe3DCh4E6zrPQaoLzOo+MtYazZhALK10Y6/rlclSoYi9y
TcleOuRKzfRHE9cSOqEoKaxh0wR3y1C1Dyt2020GKbQPE23O7jaIAlgoj+spBldNnAw9Okwrb6Hj
2ghYXpxPKRM95iDtp53oFez4q+rt0FBhV5TrLpB0lwRraYGghzWkP1sdDG2MmOjJHEjpGwegosnf
Xw1AEP2P93Cfd0t6FXEZv20a7s6mGuxq3lGDZ3FyekiDpWvpUe1bTMochmS8zwTPs5kCxccKUOK6
+Ku6WmIoRx/o1XD6awrOoGPIDAi23lxnyZZNxNCbHvv5sCm2N5B98t5i2zXYklBX7OnYEJniq+pj
qZ30GVv9MS38Kjwq8G2kHeNBzqXCMrr0vrmNtrjqCd1X/xtEZx85wkxQMZzJhr9H9Yl4bhE0V0BE
z8mh1sw7PhCB9YNDpZWLxxYchHE8i3b/y6kkRuRumHrZhahJupCRYhtGEqLloApp84gii6TI5bc0
uvlHWfZ+rlELaslJQb4brYAloiaWyEoFdAAaC2CKyiRlrmCn/m0oY4xntr08Sk0BtHXS9ui4Pamn
1+J6epzVU8qqz55cWGFSkANnBygmDRjsYNKrkBYAuIDVmKzQksZmYaxl7tJVklLlCwHl1UxO40y4
/bbiHKzvMO3flgCYZXfdQHs/qp3vKSINWA+69YNS41oY7UoJ2cmv0zvGfrym2K3Crrk9xDQJQ4eE
6ZxmB78LMvA9+YaKjYQceoAGukcpKqGATEkPTF5+bpRMn4YXcECdBIdWC8F+9Jw2hwln7x6sjVxm
1teQdaTNHcXVyeBEqAWRrAJRY64IZsZ6tdWhoU1O1ESIz4CVeQnQaJVf7lOWNUqHYur4sht1zS/l
hYjlLJElq5GZiXZGFfQcVJi8PWGD1EErOWENT4edLX5HpmAlWG8dl9ai200ouDB17EFc//iZwE3p
s6YH2JNSTioDV/UmzExm7AT9SlzvhfQxCI/4we2jiI5F6l+RCKI4uoKEB+NYnVlqmVyniERGOLz6
MHufyi64q9iTl1F9ToYRx727VWNs3nZSHaA7mFiF1Q5LXyWjXfovFa54RdNZLWm7ySvh/EZaYC3x
lqKULabQJWLiVhv1pBZxKHpEoDiJjfI5SS2ifIQXGjk3vSb7nK+dyQAB6ZwerMU5xgKV00thOXJb
TSbjxt1jagAeoBgR7Qrs1OrS1gQpm70SeThSlzuKMrMa/n6n26Wvo2CoufaT3KZVF4xRXlgFtAEG
t/z0fMxiz1Tv+W0/Qqp8DndkZeK1FNISX9IambKAuurxFlXO5bua9YAXw5L6BaEjhsn/wmvw6zEw
+qCurdHL+k3vdx/7S1oIrZLlaQ6L+apeojHObmGhTRcmEniJa1N/voIZxnKUIa+PzcX/glJhoOpG
LGSU05gQ8FEGQgXfJWW6QKNgeCjOzlI7z4jEKChEKmfc5qvzwcPSwqkzhbM//37DpbON+zWEoDkU
fPhjVd7RYlvlt3nmrW4mReRly/jwHwaiZWP3ZlNT1qFVS2/P1nwIbT7nuqFU/4IkImM+4/+vnDHZ
u48iB3WS48ydvTZOgd1G4RqF1Xkv+v0Hid4SKjfd04ZWawA+DebmHCzyB3kOrcukZKWkGQAmdi76
CnOsYaaL0yqJ0lkIz/KYCIThs5C2qfSLb4pKPsKVqSga4bn4cwqJnGoY5XGq8BK/ou2P4Zeup8Ff
smlCIJL1rVyHfS6J29tpZBihJkh72BJsJlPlX2XuBWsrX+o0saktxn3/vhYYM5iOn4oXRiWUXg6d
Ig3LhiVl6k+L/n/mIhvN4BNRYYChso8zbbEX37pDyECbHhownupO/t3aV2jrNRxSSnROgiFedEXz
yfpzYhD1ll5VxnCM2rilnm6x5/uWXMBLMtZgig34+nfQEZmVg8znBTNKylZ6sCcs5vuOwMifDux8
353UXepxrrngiP/zkeLJQU3YL9sa5T6QGp+VgA0E+cJFKhH+uA+SpdNk6pjfDMce9gXneVxZFz/O
YmZM9mfrxBMJbag88FFQf+lPQe3qhgncJbGoT0Rkx47XPYDLaQD7WmkfpFPepWsK97EbnGMRvaAR
HLg2BaXrKfhlqezsbo3rsGFCSazjQJKlZFeU47Ak5miHU3s3m9eQi5E0j8tJz6t4fAoVmYj4qiaI
oWlp08+aL3d2nOEoeuP6O28jKmU7s8Fca/veiaI2DDIl/LFNAYEb94LVhDRgLSyUijV7ieBORZbF
yD+f8KKMu9DyOcRkLJLplSOqfWWplMQcNUNJRjx3S7HE3yPXuBRt5bdoqfuM1lyUjTmq1cICzGwQ
ajejdeGgSWV42MnvaU3uyHDwXFzOjjsVkgOJ4xsEhAqAC+cVcYybvS4qIIBms88eB1wOpgK34eOe
tOsjqhuNcf/Oojf5h8gxWRpjWKC1r+EzbYlh8gWOasY5CfSiVyun19pXXUgrA9K3H5RwusYjD3Sk
XBG20uwqR+4Ib3ujVKeoiYmkdBajGWHXjSd6tY1VoFJeMGCZlsof0Yxzr/RKKnvOUEr23qEtgC00
+N/QFb6F4FA9rsBGmCjpw43P2wyHrRsasZ954D57YH6IkhP0Hn29S3yED5HO+Rwu9BFVwSOK9jJv
aW3IrXYUEKJtVLya+mysAJudBdaGAOoiVnyGnFcV9JrI5YHqdP+sEUgOr3SzCqXmEfj9jpTB7jLc
F2zEHh4cVE7y6DguwWFf44WbKY0Nc8FdfxJTjmbhRIWNVMEmM630Wohor0iPcaFFKdtB5C8h/r1c
iORv1OLyPlXsTjn15V6BYCWvQoDUgsEtyVkC8JmH7uSu8hylBAbU0/kGFKhqDlT0DFWIz7q/wJ82
9QBiT0hiMKLUaEMo/iYPGAM97gsrtJ0qjuKD08QLMNmE0XdK29pUW7UnJXGcRF+pY+IghcsL9+ex
0GoKMnqdL3pOLKnnQ4vs8misPNsH/Nl63a3NIUyQusGLYa6x5mn/uS9B4Yv3+jNHE1UVVLcfbR/w
tsug9c6C8AEzHHWyp8uIoAgZunTmAH5IOReoyYrgsKVP7vltozpr2aI2V4c5iuS4fvvTZ8NNHxbY
PeKfTf9jrd8eDQNrEEw88OxatOv4ZhBnnQuLsAx7QGn0eGoGtklOhY/P6vw73EYi200YaugkeXtO
jWSG+JQV/THyHtck9ybUmkOfeRoinD+t3yb7Y5wyVP+Acdqeyg75XcEKiwcIFZuYWimEkyNBkajK
KnHNdl8kRJEpLa/r+qxTY2yB2HIXC9/XgwO84DotXiLbPNXzRFLtlIHwICtYgCdsyhdq5xncgOmX
bgZSHImOzH9n1syFIkDEL6gqswG5Xd/Eli4uRfDlKiVdsF2qFg==
`protect end_protected
