--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
nYtD5Tajg1SLLJYSHw359TD+6sPpE7V6q/c1actGDqGsRMqLhICcJ7hhv2ZEYWHOegotKQdcgGgz
fXH0cHcu8WV4EWa/daexD93ofDNIMVQIJONo0I4srWw2cV1VhYh6P+QteeWBRQSLv6Xg3jFQgLbH
xKBaPV5UNeGSk/VyJOB+Ty9PnpiJySYq5m6v/pO7pLnOw82m6YhAyBN6IYt6QMJF+72DKiFQmA9s
jWtmuVt7b0aaa1UkvvUmgrdoCPxng1Od8CBgM3ArqkNWNpTASuHmgJGhkjzjA8QkBWXN7rvOVEtB
lEXq7CyHjJiqHBVsG9hDpz2cnlgxD10OCszxQg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="udWaM0PfAP+xYdIKKj2Aubkl79VryOxzV0lo+G2XCJo="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
lxUTpq/j0dp6weh8pRdwMzTT/BWY+P0IxzgNfhnL5YuhZ9bWxw0HZ3fHpXSKNOm7J0nU7YRyBwyD
qawXf+etVt6joaJzP8If7ofecqOHq9vU4QGJa0GWWbxD4QaFkwyg/c2sDvWOqVIHKG+Y7trWQSH+
UFFvoeNpyihE6be3ya8JW6eBtxPGBrZwRq8L+RRWlsVjDReAXdiyPfxsthISEDawNKvnNKIekJbG
A7cJ+FdwGp2+/GxZ+UF13SbIKkIsckas2XdgDagcBn/d57SkpByo2vsXhqEmngtceQkpF4dWZTmJ
NhFFFfF1GwJEFJ5vUj0I8TakIFgCCszcWd2f5A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="oRD2PguochBUfyjJh+BvVFGkyvu/FTfPU8fgl00ILqA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2512)
`protect data_block
oErw/XPw//SSMC1DfLeQ2dvt+Ag4qRqASgdcmJM1T2BCVtSH99wxtu50UAVMhAQWACb9qVkv/VJm
F/kYprFHL5/83R591JZOpo7sNIuQ9rXcLO4MTMokfFfn3d8txWzXR4OJR6IQKzkodv9xpk119dM9
A7YqUakwHldQ5TjftoN7coWQnvO5Q83F3yypmQCfVCF2hV23QMHR05OL22sKgud4Y1xhNZUUb8sn
Tm2vdX8DnvNa9QtXGk+n8zbnVe31BtulQpt4w0qkc6rPSRTCmJuW7llKTglcYYgLsy1VVSsZ8hPE
zeyO6G9aTXtv3/v34wcNmcXQeILFr4dtgFjCLaohwF4nL1xg3+8YInYaPppUUq2lIx8jNQtbfE8e
/0w5FsIW7SJjXQOXtc0aNPXFX9Rllc6xS9kN0YtXW8Q3ijoaunmfnWB3DUs5xJgv8831rmw2g7aw
hYMwN/3KEtHotyCdyngEGsh9MfG60vcuQmTb2xiMvujO1Ep3v8b34iQKd0D5HC9HHRLVIk45sSfx
GUwo2rjMUbFW/zsuygVGoZaYZSvsz5Yy6hOgf+8sxxaVdl8vRC1VxmBuFyrC7VBqRlGGEO7g7rEq
29p3lcr747SftlHxOKMXY4jKYkYYghzAVECTxrBIZLMYmATog4Q5g/UqGxQdrtu7516zh7T6yCeB
a2rF3tmf47kSM7m4lV2Ou0A1BpH8jwEcxnxadXAkf8Zf7ItxR0dWthQ4YlVef65oK9k6D0BU41zg
jAxmGFRhVMN71pqtC9tDA6LGOT76juMFjdUEkFVD0vMS0s3foROHUM2iVfUaC2ushkX5TazI2NXu
CctqPmMaepoWAexphopsDuSMhqvbWQdwTBD1dxYNATmU7V4HVXr9Jfp2R+OaLLNLf42v8y3W2Gxx
beV8jE2EfzoNN9DF54AtlR3ZszaxZkTryBF9Juqp1tuzP0/wrx+ndCMyF0VLYh/hwxaX4ODI8DrM
h9aiMXhtbDbeasJ6jqK36zuciVTFdOUyuli6wfMxOmd9/dHVC86oE+id5T7CjBgTdI47xC8qSw4L
bF4B/NeVuB+oWKDLUg99oPxLSeqM070VNBiqjFhAAq1C+yKHE+wyNkgJ4PHLKBPJRL8Try6dLS5Y
1SETKKUGIyGwKzxK78wH6PoRIbS082UXDeeXRGLcJd2J7qh88utljqiIdvK4JdybsSba2hK0KK4B
jVMKw5FIIU7glrkvTAfPABatrWDwczvLbz88CkyCcFDdKXdrFlqC4W4ccj3vs3dneAUH3b1+QuiB
rStIEQ2Dk4Cnv4vtLp1SR5vIQa3fYUkxjhSsnpFXaYHjGD8CzK8NY9G7G8gpxz5hloz52sg63sVR
8dNNhQcOPAX+pq/nd5UmY0T1zYV8GoQtJ2WQLhEj9oZHtzYDpikUe/YEgKb1R/YsY6d6isk3WuFm
rBP05zLlQZiW4lkLzDcSmYqvrIdsQ0s7JyDqapqUVOHQ6bBF86z01Ahjv7UKlUeWQZN0IcRfU6xE
xBYJydv1FLte3rg4zER1VX1DYi+SMDFYs3YsChvn4VpD4fJKs+7gBHjlXxKl2mPA9vsAf0vPuNgd
jFGGP+QCd4oS6cON+24tqv9PMIz7dv8OpgV6U5zEW2K+o06dR0HN5BihhlvplQ2eO0S2c6QK0PrQ
T2ghiGGKj2nMx6o/+uj0WWovo4GOd/e7xBBFOL1EsvIn/XLwYrtw4GcFCv/pbd1+iQpuHgP17OzS
VLHUUAa6K619HS+0/51V5lzQ45TYOOxFsh8UN/Z5z7oxXJLQ/vM9xA13/qtb1A+5lduQwHO2TlHR
vgry9WJ77K9lYy2xLvoEllDchNRyYtzY7ZIo3Y9+44wGLAOn9W/Gh8glHUs7OAlv+4jqamqMNMz4
29hjGocNyyISw1END5qSgRWAOEKUNFdJDpvP1sFm6ZC7PEZsM8OI0ROJnefaEtz2xI/lXh+tVkZ1
qqPNolg1gRuncVzrlyz2IfDm6yiKKgKps0eAeMWv9vWCEaucZpnx5Ww2yuDHfJwDfMZEeIbsSgga
O2tP8obv73PmBFIsICknaEq+aIEJplp7NQNoXlvMG4u1FIyKCWLXPOrnv5X05l3ipAzOafF4qMxq
MkgnCevCyKYpaJ4wD1NGtFtqgCVGP06QNcQPjaUhc08fWQi7HkA1EcDil2l0XpAAJM28uZ3xJxR7
9xsu+EV/5dNl1l60P8fff0+6K9G6NGIQUC7mIBRRZXhbGhB7usAeKL4gvjSWu8ahARJnAx9EMxNa
UuO+fqNczRLTNuYkOPWD+w3eSM7whgj1WGK+uHZIZPr4HFrpTAhCf2FyWobEjz8UvneZX3VXa1Jx
VKypvFCmUGteuGVoizwesD6Igz38kqkJqmF6z311gig23IhUMpN79z3EDfNrFyhiVaGuth5JluQ+
V3jf2Ndck0/ZPTuytvI5nj1NSQ1cuFIbJT/pA1G4cgBB1ChMdb3KVD/U9685lqaGgsWVxQbSRucI
JUdq+XG9EnaPvl7cu2Nyxyo05wYpJdXkF9B/0m1ZYcUgHX337bFhHxdeKAWEPlR1n4/5RVXrrinp
U/JjvwvvEWQR9zeX3nkPTzM47xQqIt9pHbH5RT4pTBvaO9e1U0mxAjwKOVfJTyCruqxjOwRQxl3H
LgTfBh5TejpZXA9cDzNgzDNk0+s5OvBe6yHOQYjA31xQpa/5ok0ai2hu7m/by3OSRQo6GMKDGcuP
pkoRDvRweMbCechAfZOObAjQ/d/Ur3bcz52+iHT5gQZoJIhujDgVyeK2M7VE901+Kd2krJc7M3Vg
2yUudJWnBuEQSXIkgt/R5SSHa4IqtZc4U2eBdciLJl1kmGE3/mrzyK3nB3FUOJrqCPnPKnXtN2Oe
aonblJKlsztpYspsStYqdXDfiS9jz7JvzT9JdHDnVEk+81Qx7AIjQFgGyHabbhmZ9k63iBR/CYpM
28ePSA7wn2FWveaXTi7A/6mKRFMIx3GY/hwFOG3zRe01QJn3xjH3/ehuKj6RiKsiP2jLyLTi2fTq
oKapRNCmVLWTywiL85sWpJmNTUFQ2iv1pmuZbRtPGRxXQK8ZRRdKJO44rcCEl40jQoAOGqatYLOr
duF6NmDdSa8+XA//nXsPFRVtLS5PghcqqRHbXsU1DHgGiryI1iXn2Vjo4avSwlLliVTnOATTkEV4
udey+u4+REdFUCCsVhftlYbCifh5h7kilbYrMDeO06q0pFx3Sxa7OouqV5KzveYOmkEF0CUy5cmK
+ZkGpYSkMLlZkUaLAg+L7wQPS66bT9D2FjI/i8bni45giWFAFGoov5bzv3bk3IAXhCbWnFGJA0kI
rn52AA==
`protect end_protected
