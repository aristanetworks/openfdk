--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Q682WDsxJeax6h1paoiGhx17CwKtRGxy9Yy8lUxaCd/CjNEfPa/ZoY544HLcmjXrqJlO2IMzCfKR
edPhc9EIFZ8RhTEEbJP1kzkVgWFl3KlDbhkQAwX/R1xmxTdnVCC4w9eaEPccHmwReMDPtWfsdDhV
hGCKInM8OlSDpalw2SSRLVbV+7W2QlnMaFLxmX6FuEWH3PuLtCOJr4kDZfBbY8Beaoi7jkiuLTCB
8tWk6TxyomJH3mNG70lcjPlfEJcx99c9RnCHDjWUJiTJDHFsk7Bu9AJVQVPJkJy53bKr3hrJorZ4
RqODZbamqv8qffCGYD2V6W1jL1DVbN2ncj9Qvg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="QxIIl7dhN+/XU8ZoRu7yDAxwCTxJDToYP49Qi0aef9I="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
mvLc+zL+gK99cH5uNw2X+3GxWdUNHPPT/3BlZW7L73ZFZMlMVKPzbWrqt+aDc9h0A2EdSdkCFqT1
98yrHTHY3AE9PWpfRAulKKHZfI+WUuSJhO1dOmT2o3RDMuVKm64ruO5RaMb5+3w+aaDzm7726ev7
9+ZzMOj0g6lZTKXGQigEDJ58Yv8vUw2tbgbS+BS8TjtuAv1IkZmjB6UWUJvjZxUXbv00AGY7brpR
o3plF96dp08NWPBETzNqql2CBVFBFrXqKBSAcJ5VVaShxtrWdG0QJqs5SfYdoVU5YeuqW3d6yjhw
WgJuAH+rSiCraVh4M3wfFOdWLExiCdOn4Jjdeg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="zm1DcnXdkwWf9zHk9hLO3B5o0DjaRpAnHfp5SW0Ggxk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2656)
`protect data_block
ZIIYd7Z50CUGnl6wNNSJvIh42V8S8oObDK8qDPPkVG+PFp4pLudJMq5UBGR82u6PdjL3KRXutB3z
A7szLpd3sK/RoXV8dgS4fYRXnWHQ6qmxAlhCoOD55+cMFA4V7hFCJVpdS0DRWMNjEyOFgEbP993k
x8/GWtjKIA2cpkLZzY2/rikC23/12ftIdEs03VuNwL4Sh7EaeQ8daziUO4RuES0unwSX4Q6tW/tO
szV6TwSPumt+zYY3U0JjJqVL8dLKBH0qTtB9oV+Jw8UzwA7C2mBjec9CBkxYS8Vz4ydDBUbDmJUm
fqWBbXXZx7aeJBVQDGoKw3vgc0viheNvFbGoY8bgGWAVUohhHy+fz3oLNMkxGGme9Q79+Ldp9ad2
5ljb72M5XCbzncl6AY/3JUsgfN/Oxu232GDJvJ0YRDAbLih74oPTPBRjnJELK3AwPHbmRM2WaQs4
rjTxNICmrVIRy3p5mRoIli4y0B3bQz5Q2AxvzWF2MppB8oWYseqzwLYvuohJELoVNKLe1yG+5T4+
Y0SF/Gh0GnOvwYH6r130nRXCNvVOz1tMwrYZ2vo3c6/fFnDKLc3m2RQixTpvC8kKCIoi5MEF8+Ib
/4G/YoPINvJFJz5o11byqVdU0OzJBbEA9t4/+q+N4+Y2zFYTFgRCJX68CtpE6mchY4ijhOrYloko
yMIfwf98NTTjCssZ0mmx0e7iZ7z11Iun4WmVRXKh+5MxCot4tatWTuheyfjllfgsyU2JgRMcl/b1
kHyng2DRl1EcX2+Lnr6BYE+jVMcd9SSPdwHllaWAfuC8osD1LHoHkQ8jV8ilIsDiGxhkg+u+nFlf
/f7CCGcfTJsYPex/vuompdHiSchcdIiSGHxcc/36FGhIlXjPoFInOoI/1XKsG/OqptLoNxO6uDew
QrQfGG6lPIjdopGjNgYJN2O2YePW85RJ73TEn12vDyEiP7b869qBkVDLcVmOmgnCPwW6Xr/2aFHw
VQosylbhuBSjJHsMHBoCILvYykPOBsUlu4ijQdwbWjcJ0EwVaWYNzgphj+kv9bmQqsq1C0rGWTyM
BGBbR7AkkKuit8twTnkMGUtpnOt3kgPt7d2uqpuP5ro7bMPeKx8LdvQaSLfICqXNUQXxJsjpPoI1
QO/zC66l3EJ5x9qLBSLvPLM0IkGEbuOeQoDxzXEuNELSFN3bdBL3++QOAYl5J3pzx0s+/EHdgi7t
sPowSuNMFVBlZL6a5BL1BEz/4WmXyIIjGWtwsnMeVYbnbYsCf0RBdCEV+OEu3toibGAuaxrJDgi9
USkBQGfOd17enBrUH3gyISy04ua8cBA1pV3SyuIMj5TxzOjtqp7K/AFRrrmzSVFF/Up+ESIOO/tw
pBifk9ZZJMWcpy0dUNaak9N2nMyXrc/hBqWk7epgip3iagKsgJptPcrL7Yv2IuRHq3mWdHVlgLqG
XC1gtFXiqySMMxdrypaUzy8N6Pom0WeHffEe3zSH7K9sDV8OG7y5OohcEpcM/z4OFUM/g87rM7oL
QF8qTWvbPxOssWMNQJ6EvRx4q9g2awgWmCj4DnzL/AaVx9Qv/cePnG+mmOkcByCduzjkfOJOH4sT
npIY5EwdDv3awEO1vPg9L597nPYtw96kOCqYZ2NZZLvPMle/KpjEDffhrDviZhtaae4JoLZ49/Y4
M2NEBGGUOwNRVQyQQKMlpIkoaRwBOsk4T4vueHCKuwTRj7ZutkXFNkI6xQU7sez9d363WACHBmGt
IQ7sSWcF1rVNnNFxbwY6+HXg/nCN4HnGvN+AKvFYf+4nYLvFzQgvUhO18HScBIWNqkqPRHYn0tYD
xuuMKm0uBFfUv5ttljM+vlb51aonn7I+spNifoJxf+PROmT8DCmcdl4P0V/s+/sKjCiGiT8JS4K7
ChGUKMTncEmJuTtu3qsLOVOWIr3IPMYKdFLEMy375kUV9W9VhhAcNOigal9tu5/gCfhw8ajw2wkV
59ty3mBbZB2YuxnuDHFPMvzCCVYaXLJjqCdBFgStkq73Od915hZWk3brw9e4OIOP+t31U2Nm+lNd
zVKhw6PZhQGEg+qO6/0LIZ5rnfCmBGMz0FDTlK/04ZLKvcKAe4qZuQiaCQi+ntj5q9H7l2NWLLLp
kLR+cf1QyWS6E/q0/sUrHz2beWWKlKdG/dz4darqWdqjwwfOSC39IxtIyoSuZllIVq6HNEIbRCBd
z2/YI2RdqY/iLgExpbJVJF0aTh8C90oWEq6bHTFqykCHhZ6Qav/05/bQnCL+FKxtlXG/xEBzgPOb
Q4LndtNYGZKGns0EDRXiwfMz9Nf1hXZ7cNqrBO8sCM6azDADMjXMp3H7ZrFL1zO4rQAlg7g/70Sq
3zeuphjne6bb41slM6BwCXV+XG3bUdFJUIUOeD97B2EPKt2jzQUdasMrXSROZgbIEp5HEEAjxF9E
Ie8n6PNXvhpJNNCw4f0swCNUTyEx4VuwuHan2rh4NVbm0AJB6RGayv1q4Uameo6Gl8DM7TyKqvgF
wqOvpTTonkAMPRz8iiWSANS8Z42Bd53uR6dDaO3ArgN8JPg/rs9hwE+Li8AjJuLsyoyxIhjuKD4k
mfY6Pf+Gbe7EKpm78GhyiQH580afwR86aPB0+NGalioo7te5ebJDBCuo6hnS3Ku+T7Wlg77l1RaX
Q3mIx6rMNSTJZ1CJHofzn05GsjMFsjiuPa4fWQMO6un0/UFSLIoznRewUedpiWOKsvGwbahJ2aSM
nERVCGEu1ukDvRFAJ1VFhTNjXHDpNnrLpRcunXBYDluWCtF8ikCtHsVMIjAuhvCIdQvzS41UX0kk
qo26I7dv9ybu+TTo4A+nqiRndbKbx7fxG3R17ijSVLVH4E0VzdQe5p9Et/vIYGQWNTqny/fBemCa
RoXYs8jXiGsMsy3b7sqTA08ViN0Jo+SAKzjwDPQiIVJO0tf/oeGb3R0/7SmPJJZ5EH4gsQGdOThz
gST054ho3HYHoBEOakBbeIHC5cEurf90tpeVpUyGQrkUX5lw23LyCSTvFDGG/kTmoJOHN4Kv2e1w
/zX3zI8F4LCpqazkQwl/LZHTX1xtz/2V1fo0ADXdV92CypT3R+d+aGh9gkD12PxpZKK+tU0PHm89
6/jvqlDBGGlotz/xn1ZX5J269ltA7ncDb1zwWjd9Owgw0CBZzsoNwrjg+XPLc6oNeGZlYlY3zUH8
azA7T+5qJwLXvEbTXuPD8M9uDV/10WE7dZHCoL7w8Tt5FgErxXpRHW8+UnrPz8/H0N9qWOUE5Uvk
cTxD0qovQ6Vm4D/2BAAV1QdGQvTh7Cjgxw19BirVWXz+wGB2a+6Z6kTWiXFqCpscjGz6cY7JLX6w
GUTETpDkeX4rdrjaOW6m36mEJBrX18cYnlo5WE5z0aoJ5/Vly4q2IXPD4hF8wEYR5cXOwjO5kYPM
MSD+0spTqHDMgIelt8JRfNGD4y+c/Vg6lq20PE0Uj/Gbl67rQkDON1sxpoLESjmFxQZw9hRS0rlX
5a8lafxmGsezhOcOtbdZwORSbcE66bHMV7xBJ5qj8K4gvg==
`protect end_protected
