--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
UozIQRE/bmrDaQ7rTI2lv4OjY8c5V1T+24zKadX/tvy9HisXgMEl/vw7GD1nWZwNGsDx9MsIrp5D
QLw8RURd0k0XNj1tV2uH8grgkiu0/YfkU0co51gx4UeeUqY/6dKGuar33GMTAHhcwZMbq6lxxFZP
lZKuM+oiCBQdtfybmtmQTJSIQEUs6yikPfwlWfP2zzka0GnGX8HUamZ7SFlrEIho/B/grvqASIrE
Y306ko7s9xJY7Z96n6aD3c9Yqeb3V4jaUBNnAcPJtGO+CJ5iLYRu2v3q94HKyIktf87Lw8x6SLmL
ZYBWyhIwS9e+yP1RZS9YTknUOCR0HPa8iT5r+A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="bvRb/HE25CD9SW8Vek47v1O3xOEOAItt11A0tUgdafQ="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
ejLjbxOnNvp7Vjctw+RnFCXWEal9h06pn5W55wJ87zppxlmTeIVVDw7Ho4wqureSvH1J5YZij1s6
bPp+ythOmBOngiuBQpUBU1zhPy55Pd2EiwZ66VXrXWKi+bD1KJd8LXDnBO5danTuAQliX/ss6sWU
fCsPGJyJ403rn/o91/kzqJL+ABugB5C1JEL5uQjOVjmtCl8Vb9HPkwvlWHDaOlp91a9PApGSmZ61
UXoubLzdS7AObVxBvHeSCnzvQzjt5LlRI9CNfJEcLr7edzzWFQHfw7DTAtgBoklVlpLVHGjplqSb
Yv2WzHNJgYGAsij6yUhcki1mddjU/keT9eEFDw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="i60v2mOns65a3xXQLYV+GV663/mcJqTjmpAjzSIDZ7c="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34720)
`protect data_block
3txvKM74lhcmY5PCABbzRZ66BIo1NUOcdgBXfI+ITBXl1YoIVfKK30h7rrLjmsqI9ZvGpCqyZxBD
lEQ2DNdNGeb/kT3es2S2X31wQycTCKxLPzdWwftVU4kvaCVXekAjMJNVbKKJcoNIZLD+FFJ1iBrE
R/NgWwW1hMKzBq9p4VS8YnaPSF24sUQTxkZInTmD5qC2aonV607NN//P/OoLP5UVro2D8IWohQSp
ChU3zktAF4ZioH05UI8XPx2JMATquqNv7OE8XHApTZRD0UQCpweIyDJhB2IkNeTYnkbxOcEFXXfV
p/d6nuY6JXaKMS5Vf5jgBTuwCOMytEUnLQFtcdQQKxGv+AoBmrEDFpu0reaZ5negFqswALs1HyHH
Tp9sagYkISmGFzKg9MoQMkn1TB5Q4UqqMi3P4GuiSK6g4XoO/u5fEc/ViAHWv8Ptb//PAu04jobB
/aKpxLJng9emAK2XoB1nuiPjz5wSh8PvsCqDtV6WFMy5qwmm+Trm3LH7FgOOzFnDXD9v2CK8JAOs
bIZMeC8YaF7vqpCI4Uzkdrjxup1mJc+DSZnBEzPcZwyZW6j+Y9K/CynJpquW3lXyte9zK+PzRI/h
Y8sIxdxmlvxv2GrgdONRt/x1tQAqymXNJp2yRqmeOQPOtriChNcAWzhaSzY5f6qvvqtxa+MwLOWl
5trln/d2DSvNCS/PjRFwkhrNyVW1PWIjGmhH36qrnegUrtc/gHRQ1eFHZwVvu/a4j39RhnujyTaR
VrfkXucw7h+bWEAkH40ltJY3F5d5awexjRlC0bz/V5gGwTumpS8xsl0ifnSySC+ukvCn4VKpS9+K
cK+ONZOiHgYbcPRu0iYL9/JNmp1NtS/aJLWOZzS2kpUJe2KZmpsqh0COjTwjOTEMCq9RXqLf0gDe
pXqqgTMqUsfXg9W74rXMA+qdfbFbVCoZP/gC0cj+V9lOzArsJf1fz0DmuzllmtlWzvPflBtjRY6W
Gi8qz98ZaQIiTWW2pmgHE1trwQKyzUVexNUZdErHjT31NDeCd+4QN9Zp/xFa9KjOBA183RglaLYK
mnbOLOmghUG8+RW52GoeHV1QqAEM8Fl5AvUveC1e5EyyKle8oLWTXJQbKjZxk9QjM6M+K7UuFKBj
6cbEEDeoK8P+idmDnyWKtN2wCGUR0z0gl+5+kI2t9Idncjq3hNRlrkM7FpIlN8qmzKCh3udTqbNM
p5NEUss1SbZrgdwL9C5cc0XYa5DaiLLKyhkCYTq6/V8JN0LGf0NrRFCI1i7auwJjL7VYesXU6xrS
mVZuWagjE8zIxiFbqGaQacoNj/2CNJKXqTqCnbKY8FrR5tRhKsYT2e0Qs9iQy5asBJzi8RRhRcm6
8rwiv2PbY2xZUCc7dUcQxKjJr33jIQuQ2tehW0xigFKJfxZdEgl38jUg3b0v1Z6ZO0hQ7O/+9y63
fEjeIoHcALm6W7LlCqTYgHPiA91MUcHD4hVtGGyXaQimrd+VGoay0ZCnzME2c7mE22bWDKXI77tZ
eGLrlUMS2oJWfHn4mRK2eb3NjmTVy7LiIAh0u2/6dn3HdkYvsxTFBD50N/3dciXnwHzdaPBWS5Tn
CJsy0p02ZrKmkdYlaSc+oWMCge0w1c2RtWYEimGOmy2dwBzbHvqDGmo35qLZAHM8tTQemV4VkoQ7
HZJ1E8n2Hillo7do6lBx089CEcqNYkkBOvGAZd/aUecm3g+/nbMgiDvpwHV5MtW8GZUsNjQOPobX
kMEvRu38Hrb/l+QjjYNKQeg7mqQFSGwwBROLSDf6xv0IEpybLRIdgPivt34wvrDIl5+H+AxOedSR
sW+PICVVEVlPkofcUOg/wtYC31s9SO8Zun+bHgtw+sEjh1br7XDaY/ouXp9HHwGE7an2McHWUYaU
7oK1GRdneYdUB9mSgyRnyctsHLiDu2H6RuKVJTedWMQdnAUbkADOnAs2XagRzzoWY9qi+8mZE8ow
nkX93cm4s3533mQyD1dVflzoMfxyfPBmpyzi97zDq2ryGqA5zNJ8I8O20z7ERzpz9Ac+rsX1qjio
+++Ksyx8PKeWTfKS/b9XhlCxKsV0btRL+zuNt3fhJ0XJjfvvpTrZIoC45PQXlwtpEGsRVBfgtfb0
K31sJAx79gTkZDwuidluWdI/FVkybbTshCd+svv0MRAMbBYjMzL1eQRiME67LgPVm18f0Mp5yGWB
xtxL94r4g/A0gErWbCzOTPa2bMPhwgsUjyJsOw64eoDBGq1bB4FAOzgtljHmwarMbfAe83d3k/io
SJjuT5QykMXapAhgnSXgQyJAoMH4LP03ze/LAaFOVrysAAiRiQUhEeiK0H3gdKRZVU061VzRfbx5
FRzdBk2VNWvN4DnI8bDKNA17PwxqR6+CkzzN0NuizmYsOQPqHMP4J3pGonwFvNY29hTIypLx0nQ0
Q4s24OJvnH7BVCKeNuygNBBIE9dBofrMnNOX9YaEyUHqDhFvepNil3+/nSnw6weifcySAQPuGcHf
6uql7s6Bd+1G+ebrRDx+1wY48PfO2l7WoYgpafxRFlViA/KQluKIkU4KfGycZASstKR5lIvQ9Nkk
XntQ6c7pcV+LTVpeRKgXtH/dwGLuIP5Xoy4mDgvOv+Emrf5EEOIitmowMykn3cNDP3vobhvii6VR
5BnxkYxBEgsyKH97P4ixyitoASESKEAv7P5iBU+QbPDOBigVMxHEvXA/wUECTe0ao8hjF8/MpFXA
ZFkvGVpXku3nS9SSzsaM0wfD2CE/kCmiE63PVOiRKFqFNnsJnQ0DupmswUaGU3m1wKgaoqjJPxkS
Ge8ysJ9n7QIAAkc2zbAwBnxY+hB11/iW1ielT3QeSlOV7NcH8cIn5PGDyxuKxm7SD9je8rHekKlV
bn8wmKqgMsO1AWSXRD7tCe3Az+OBWwcpZsJNegF+LNfSSwRATOhyyjcBib9AHEFS5vBcrljGCecr
xYP4KfXlUc67pdfBOzA6w6ihocH43N0G671KBVpeTRfE1zylZc8b77ZGRfe0yPr5XSZWZtpAdf7J
QmKdtTWunGB9bZMl+3RiqBMcR77vmgn9vKyGGQbTbGySxPTX4XpMNyvhWktVn1zZpJfLLe2OCWC6
QhAA2m9LW0UFIghLbO1U2wNHfmkLN2dFNe1k//y+FtpdlX7YpKug1U68nOhEzRmDJF3Tw9vM6rVW
1WaFzH+SnUwe2QWZW96EjvjGA0TP69CwvF+SbC4trsoZ7OePPDzyO+s62gOgKst3Dbq+VY1sYmtt
xJFnBkx2KQzEaLUUP5fPofhUJBi+9xKXD8lEsuL80Jpgx4s7Et4LPzsoOdKiY93Nhf7Zi13nL76B
HAJeqN1LtFDc+6qi4BECYzepSPo9k3U6/b/uJgqba8PeLFh9RDhkohWvqEH/pnPJxTv+VOSessRi
E1wnbrJKPT6T2+0wQ2z12DjolvwVIvvZimo6S88VDcMzcfI8vH7+d9aogDcwnQz2nz+bTdbNW37E
FBVE1Ya5/WBEWFlkJdMQCWaObmGB5dgdWE0sq61oUvEHoKgOfEHJB4h9ItW3+lElegX07yb1tZfD
iit3U84rcK+IYvnSwLAAnTKS5rgsteUqsBbFCKmD9ssGO6+gX/ad0QRFweSsB6N0N19B0EtNXrmP
z1Y56bU3X0utjAXcjH43nFbjTM+g11qGW3za9MxJMULM3e/hg7ef+lLJndKlSIpRzHZlgcmAluo9
LgOMOCOP8SCktW3eiCcGvguQmhcAjxIv5Xw/YkWVs0LIdk0tE2At7EXlWlgKPHQkXm3BLtbTXO34
DNZSeqqw+EO4g/zJqlHOboA7AnYpwI+me8gu6hAzb/qme5b42UKRZZws18wJq92YN20CMJ6sEZcA
CuKnqQS85yNLMFfKV7OSVEr4MdsDb5VmKx5DE2ZqWEqPCtkRy3OPawbYnxSexrKrDrcVQIhFiGCG
ecFA1/yVHXSVUGy36JGm5tBTkLww3ouhq8+sh7wbpPtDnpsOmXdhJ0UDnwdU54dEKodUsDwKIajC
o5U8dSaw56L54yE3hI8v9XIOxBRfwme/xlYqBP1iAARfrvFyg8ki/ARleABwFQyt7cTNKWSnbMtg
YZNXUYm9+aeuaVKB4SllWiIvKKA8lQCJTdoHnWjsgRAQwY+pHoW2kQrP7iFy2ImhgnENXe+DdKij
OS6PrvCH0xQ/zVraZZTvdQOSVn2RmgnWkluKgmNYLxxYLqpZfjuBtNPf7yWN+eg0++/UQ2aGT1je
NYKVj/9Y1B6tWylnGl6wbVOhM/0eAFSWzdmy9NTRdOrmAoj3z1tYmnMxo2jyamTjdAijNRbbS09E
QlR4rV1GGZ/h4IwUqYWPbT0NT9nl/9qW19qqr+Q+B94FvJ4BJLTIE7RLWoYmfhtzF7Gt0mfQ9PN9
ur+8VfqyVoiTElgcSbH2XaZQ8JmRUyq5p3ZytD6Vv8f0+atOmIxoi+r+3K7yAnVDZ9XlACZKzzlP
Fo5tn8Dedg25XybH5TkUvZoKj4MRTHm467P1hOwr+ZqIzMzckE+gpESbn9uXTLb/9M9qC+DUFPml
tilwNksLX6b75sfmX5kby3lEelgNrDUc0idGKYe5/w0cbAomxaF3gmS5O15e9FWfB59kZ/653bMW
xDKQGaK0vnQtqMRRF0u7913Ja8syoYN9PuS7OWiwO84KcFepII0PMSQZjzhcCzFafAcF570cx4o1
6ubRZImSDI2oN/G6FZR92JbucV0XXASFhwJL+6+jr6IJ2YPc8FuQyQdIaZeMFMYj+JeQ2hDeP+eZ
shHTDBfpuuUSi65vt+BWhdhhc8BVSw/nmibdWoYTlron/+7MJeg0lEZCtchmf/jB3cO2vx2dDdJj
pC2AbPDQMxYm1avBU2ffZrqoSFj+D9uVWMdusD7tz3yd78XYYOYvVpNWEw6c3nIAQQBUOB0XPBv2
eFbLnrZcrNIb2906HU0F5tTXvfxwzBke1kbqITqXkvzVgOJKrjvpP93g9qICTw+c3n2ZjjPrxzjw
9hk4/DPSkzZsGpJ+Em4FypSzdN4SfsKcjNM3MdLSgLzHPQwiiSDpezzVS4RlUmy/ouMTd6wmO5y9
HNR+lyhwh2XlffCQFo0EGz7f9DeVFgO8m9qaSRd75SY5Y5f7Qh2z4u2NUZd+1xgNWcAvEKhFfDVa
5iuG/IQwRDN6u5nn5EQuvmK/pPOnBSQnPKsGTKfjPQhHT1ctquIh5t6UHgVBbzfE/kRvTe9rk9c+
kKTXr3wW2yj3R/elNZawNzTCyuw8nCmy9+2VpMFKR0qaal02MF4T6RCMvSdFSw8uDLL3U2XN0vu8
YHR/ArK/eA6t5vRw8BUgLybGvFp7JsAogROko0z0SWBlzVGncdxqWa/d/PuomrUa2jcz0MNZzn80
b3WHPUhorStese7tebWScevLEqgwFVSFnLibEF5pXw5H/LZSlViukFlTDF/7gsHDXJJzmZGbvtgr
MYRg7RiHsOV744gxr4XNRSYAYWe1n24QQlnXSctBkVes4C1DhjUx+BJMnz7XfUS7ZePXIOWCY3ue
kbhXlP8Ip9/hA+dIZMq1OMQQcp1zYxGQmgxTe4teTPAgxhgIZI43x9jCZqRw8TkPYzb0F0NpgUoK
3W4X3JHRu6bz8esV501q5JJIGd1SIoW8Qoo7ITwaBm1WMaLIUy8oFyoPrsPYEUHR8lLTNiqAYWkn
zQdoUjF1hbhFHNcqbWBd7cGYobxJ8AxpszQyAUzDevHABdTZLudxPeGJyh5jPgcQPiE7wz/uXVWL
DORwOyxK4rTLWA9kcKnJt8G9W1byQtLSlXB1uJl+VF7c6GSLPt88NQqfLzBuSqfypm72jVFvp8Il
/UudnBEJYLeSZ0LeLJv7FC68EY5LZSy+LMnyGsRp5VCMP5Uq2bnWOBtFeM/LIpafhwcK1vGR0sKQ
SRKrtJNHR3pp+L2f0mM51rAfDk+N9DjXrOaDmiiO8OZQ2/MLqqRnReG1/+OheHMO15vs/j/rVtuv
iTaUJkcMWgJq40u5c+jY/usdGo6m4kf2NdZOSM/XEYkUk5ZW5t1VMaDx+j0+bWIdfh2b9GYSK/NJ
EXMFONn3yongSrHT0pc7akaNt76No4SoE7N7fi2wRCCQOLcGEnckv4JM/dV0P1Nacnq1Y7kvsMrZ
/CqF3YChrCXca27MdGTY1RXI/c7PYMPhJKyEDsiD6OQeFZrk+iA0rBxQ6/DVv/ZnYYkLBggkCkK7
zgic+F7UemDI1l5S07OGIYlND1xSBhhK9OhGmMQ4YJOKElHLXYqQqFq55xDqTGiR3rOUXJr0WzB1
55fuEFY2bT/d7iCprhCs9sk+UZheLEVgbx0nrCtMSTbJdK3x19rjNe58X36RTMtsQqZkFTvHyj4f
ypGkP9UdTCuN9QPiAo0NAX8R+3Pe5caRRe1yOrRx91G0l4V92dVFf4Wv1fLRhG5kL4qO+HizfXyG
CABlC7TT8zA+2/E+HmMrLqY5arEc2sm8SLyHW24mFnZFRE/doxD1Pi1z8ihMduabEsX69lYPlETE
vBeC5g2wCmYFVqlTKLh2QI4a2ofodHUg/hzV/t426vt7Df4pWTiQa2sc/i7YrPf45rsbKxMMzh/4
tSlVsinVVbCmSxB4E2dQgKO1ivQc32ZPHlYre4Xqc75G7ZHEo+RUV0ph5E6snAkmXyRp+/3syr3B
g7L/DhnbSIX1NruxlCCpQilW7eijHqEe3UY4rV/9yyOa/lDRZAaMolQ5KUvV+UiP9ilcuBW0/fNw
rFmBA7VDlo2NEBzzXZ8K0zgYLzpCed8YZizeM+nqOUlOvZbuvwM4CSPuFHB781vexxd+ldIaM9Yg
JJjFFQNH16pO+00VpaRYqLREpdtY3UwuP2HUzzsghQhhBt9U119L00cB6J0n5SFqO34fMoZ9tMjL
W/J962UVbn3PHg/1Q0qGGBww66b4XKFwXGz3dz3bMK9U5GmPijgZZST5RWvQseTWdp4MRfQ95WQr
Sy8k3vJ56PRePP8wnrQ1MsTfH4Um74Q9qa59SoJb1UuC8wb73JxgSDoeg2UiYSpyjxm3ucsXNEfC
Hy8i6cbNip1jRWKvk41Qaa3TsgswtRA4UINlMErOYa01/5Xem1A4ha4MEaWIOH0Muz66pUYAcJsx
OHFcDyylFrPtn7XyCFr62Y6W6Qk7/K8AP8yccT0mFG9Yu3NqD0udysyFAwd0FEArzIF8g7M8JEQ6
fW8w4Jnk5MruA307Ng0dN+Eh4fFCKhv9/Wy59aheQ2fIKZUuYfIMUGElGrF2ggS3E1enBr/nWHHk
a4jQjTwraAMwwpp7MePgGTu3WVOV5HXpqhLx1OuxciJuDXOCmnANXfV43eWTQImN/TAZBxUQaxa8
DND4tswMCIgnjBeaX2mtIa1oZ+/8hfaEUUfU+wtGVRgMiZCCIsLgW6QoEvQIVsEUCsxTErIrHIXn
7EmH9Uz2XYxhyeKu46MxoOkJ3jXWvQxathtADMOsoqDBX2G7ncCAgqm9jOhFxwEePHpagmpl/1Q6
BGiHQKoFlKksWxZZr3jpXJ7e1RhF3UN2HxcqxDii6mRBy33GqHJEopIMQbfNXjMcr+EqrV5bloI/
v4GsS8WSgyO9vu4EWbC148kP2MXDtHz0H489t1P9mH3SRnoK1PPoPDfjvcPa0pDSbc2L/jqbOzCk
fFI/L+50I3QoBm2WohDyzkDLRChwGyX3wWKyN15A61Rr2QHazBSPxgwZ4Zuv3lKlRkcx7zxB5yWZ
58KITU0rihhxdm0vnKIn4RZoyjCCkzNnZ8PTAHGKDZWf+Ojt8bkLUeKYF5k7/xYRWS0qHXmvEo0D
YYtCC2fs4j4wwPLMlq15W1DUHiFCA9wYEhygDJyJRmfxW+h4SxRurVWZCkgMA+SCQGgGB4eCOr2S
ExlKwe9rhoGZtQINq7Pi/XtAVuRnF3nOKncRpP9P7CcW3VE8dg54/kA1YLJ2Gi1aGVy44bo90w6N
5j1MlpE8I79FekHLSrqDw5BQASUwZC0eV9lNCmJyUgaeDoIh6stbY9WRzCWBuSf9SbfNEmFlkTH4
trHM8WUseiR8lioT4PZDwNNHTXQFxOBzhX//31zACl33WdZgqX+PALpCgKn3+o6QkZWMY5ZHE32h
s8jzO5Fsm65SZyCzZBndgWQLb3EAD5vEnjkcCwWgeau5ZBn+YdiUtcBwhx0jTDXPhjIw7p+QlnGA
PtMUtF3+d8kemMCunpK7jiprzrTPRNbF228uyuF2WXTyeqkWO+GTFxLMzfbS46F3RtUEwgxrkIuq
hPw0ArCTgG6JUBGD1eSTP59Gf1mEKao5J57mPjgdbgFz9rr7m1FiioYMenXCpd7NWizKY+x9nTNV
fa439EQ6zwI7Ep40Qyup5IiaG0khy6xBy+gGGE9nFJIyS21jNkh1M6fMRZMzkG4c7fdP9+1KFdgg
UuBhfhyBzhWL0gxogtNR/PvQCg3RrDSRaMMBsGnNO7p9aSy3F+Xu5PH8JcsNxYUkaTCPkH6l9AEY
Uwx28I15qEB55kaUk0+xsyzwcPXSjV6bg0ElPudn5pUnQFmIBYEHJik5fhylRW6WpbVMTLRci/eh
0i6MTRZ3FhcnBm8zErJXW8mAJpwxvK8RbGMSqgVqJKDqNL0gMdBGN3f8khieQkYHdIQ4rYAVVEUv
ZXZE04yHNQ07ZFgDwuO6jIF4GY8eR24o9VDwEpkqnydwjGJ1JDk6cbaT+qYo+USUmyeXObdlXMUY
WapT+k0BGuRIT9TOW1H6TROuqkWgRyRhx5br5z2GVi0+oGvwVti5R2jQBr+QSziQVG/vQQJaez+1
DH4e3w18R7ODMeKoJ6/Mcp6G0k+xifx6DR6Cy8SJBuZ+nfSjia0JuEjnmgalio0rrdPW0HZJBPHj
ZZrDjxWotSw/0jNCARXOVvxF/eFmWy+W1/7UvV/txdymy87P0yKaRa74yhwSOkFNopumqzMqoAwu
SeII0qquTI4ofFGWon8SVScdbGq6AIYKJpWqsp+MxxycQ91CtMQTk5M9uspqVn06i5sm4GE/r/PO
Mwc4rrgNejay1qUoY+mct9DGXnjfesze+FM63RPSbMyNVwbBoafFmyru2gX/iyFddOD6tmqJhsJt
GdrBA+MUUQmN1avjM22YtzeoKkbl6k5jfhNgJEaPJ+W9M+UdG/Aw0+4mR8fptZWJb0GeiBoSTdr7
vc6PJo/LGKhbzu8oMBFFNQmVGvn3mvTDMupPC8RVvSo4MZ7XrzXoSq2V1s0/OTK/69MwkYCZBkvs
cJZpH1ZlW46Oah4a27PndEAB6NuD8zKuhtvb1iDcKTILICzhAhk3/1Pkaeo2GkxocBINKHnv1naM
OW2HeoMPreNeBpHMe7g/tIiC9z50eHg21ySVluqyx7Bq3x3Q3bnkSbukQErRVMIA5FCWB+OzdSDw
YWJWs18yoAPKPNhvlj/X5Fl4jEsvlQWW4A2cFIhLQLqsGM1cV4VhofgZrGUmt0fwE7kE0HAXxmAr
kmFQkfHhklaPs6YqzoqNU1IOqLsFUSyBJ9+wHoSA97jfp/iKJP2XHE04wT0ZIJhninbNJQHCBATM
+2SgZjTvylqEJFBETf7wa4W6iR9zc2ZGaZwM0eM4sia+M8Wkes8wTRhohgrKKZ6IW391DN6v2xJC
9XYKdn/Se3L2XBVnE6vCISwce7P++jmGgNJ9C9ZSGe0n05gkFOWSauDXWktGMpPdfyPMqDzk/bvL
2p6HEmFnbuJQpFh7Be7UfBqc8+8wXNmTPAwVco+wXt7w1wzkLrErN0+gGu/mzXKK91ebH2uKLOol
mV41IJRzQ7dTccuE5ddsb6Hoq06UKUKdFn/BeaUSVasArrFJC4YQYNXuU+WAk4KZsxLEZQKFzKKG
N+DhLLqrvPzvP4DmcPDuuZX/pAjnuvWfqNRgQpYYxE5ZwswaarFFvCg8CZxE9uMaMCPbyoCpfuBX
OciiO+bxaitW9X8OldRRypZ5cNm5oPFdgWOuaQpxJiubkeqM1XGNF/XVMB0z5cn2Y1+PDjCVdSiI
vnvE8gfIxp699FM2d+2WHJoYLsdt2cRWLbt4TBM7yttIGoi5VI63jfavdz3qWaiGGXVjIsUk3o0E
j4eWnJHQ7zKDHU4/83R1HEn3CdHuH9kSS0wPNY7rimyp6Z/UWxnO/7Gr0UOIUXqR/fPeF/KOhft9
ld3k9CYhiMISJR+mXeW+g8p4BwfkQue+P3AKo0/3IJD5lLSGTzC9MkiGjNl+QKKM11knHWjtj4Dh
xIqI69Nxh/3sovhouRI8ad+bMDjTz0KFBxn2PtHff/VYrgOfwpRIQzc8NkDf/6YTv2fva7c3YXkH
ltzolkqM6tWbBgjzaziNK95yaRqNGoulzfRktOMsGYsAmv+/28eoxMt10MV64+MTlVN5eO8G+TY8
6qz3jH13ynfIDD3p/S88bRizCcyqDJhOm5IE6otI2pXwSThNl1VFKX6YXslsCRgKnAxVKd7v+W1k
ApImGoQ8kbopIUX30+58GMuOWw+7DlupgPHehByt58C6miGgPlBkY4DExveXLDXsAtTRQUxMOTVR
tImBHpowiP4aHnxZkQ+4v2Ps5fscmHvRIVCCAwyAz0FTbxSjZ5NSHDm5w5qaBuCL5DD0PqXXvsP7
eqPxvxrHwG/O/KHRqIonH3SNfyJwq+NMzekP+8k9P7OsOwuW74Sf/fSSCuKy6Rnd4rKAfMsJ5zT9
Y/Tl74x7eli/hBap1tHxE9l77c7c3hek4VhPzLCEL51O7Mh0qeDzCDyxeZdct6UDJqXTJFbM5Tdt
yvRUeS5DS2ekD+2x51MG9HuOFi7/IHhodbIRahSeT/crwJGWxvK1NzKsmSZwe6MKRfIDHFlzlcon
gi533wYe2zJK+sxi1gnbam0N/9dnMts1IjMsiJez7ZrucjoIUD4cl6/evo7hmwp+f21ULS48L2wL
w9O53uC+6px5oJJF1YRoop2PV77vz4D3vLNa7m7AAKgMW9aM0t1rHLBJSlH3wpIHrhREbLAhZJMB
iRKP2pzYPLFX5Bld7r/cTdlScvkR+WMC1PUCESuz+HrY3gcDxpdPK+ZvhOJiEV5bnehwl6epeK3p
9v94ONNX4e0QX6n5QxYyFkxELRemkkpPTbAewxw0RRbruoCH09lH+EtRh715ZZGb9xM5H4AMFelO
b0zhtXQAKUpX/bX8Gbqy1bO5ypQEn9mOUbltLhRxyD7UF7rPxGQdhUQiT6qzAwQmh6suQueooxjE
ggd4quyF+wLLHcPTYVVUuyF70wPhNyTXXHUF0OkNbslVD2AreFa8XncWsss4dLw9F6Qw/eIhSAR/
yGQBndzbHyQS8UAv5H2U9J3UpqURrMKb3HDZy5uLAV2wcr1Nnyc33ghzQX67uM1gflc50DKMeJxJ
j7rCl7m5owL3WVn+B7rMOQDAr0uH8NjPmlWASPTwNfQTpr+oCRRuc1X7JhD8CNuKX3I8EfnEaTsH
iMOMvzSrzfrsxSAFsfTvZvv5fpLMMse08GEygR8YA13tzvEUFLSHc9221AisUhreE9p252JUDyxT
UQsctSX8G5TebHQZEeK2Sv2ajY5NIxpsMHtLvJiic6FC577kVAoWQ+BBDz0S/Uw+27HDZ8zDQS7n
dL3X41y1z+y0aoCxzGNvxFmhzJgF+msoCuc29UZf4lMAcFqHYjEV2b00vrSusc1IoMzIAd89vBaH
BdDzOBgd94YMaguc05/7bh86Z74mkyXE/gzHkc70/04Eqztasrl3WeciZUK4MP/gRTVaxRyQzCKQ
PMsJorIRHBAWKSHLZJAiC2Ulw5s9U0h6BGQfX4Gd54jZuerGDNti2AuCKabWm2wTL5ZA7MtLtOfk
sjWPygnGivCIuwAB6WIYWhHofo/nxkXkUUgIQglYTQF7tRVkRNMbya1Y4U4KxCA06jjXym9RbnmW
Ek9CiEmU/NhMshF3IzAiETKXlyltOYVvIkTMrZ5LXo+CK9iGfiUdgOjT5l1BApU/2kT3muzio0xf
+NwhvP2KX6OmZ0oHTUcJd0HcY05sJWijak8v6J3I1ymWrt6CCWZ0B7LxXfIbFoOquHQDhfVV52Ij
ls5PGbSz96zAfdVlK59fIusCur35+snTmKzKkHIGRsgEXbgI94Oz2s6fmLPlvGjkTdTQLOKIat7D
RpJkV0PRv5yIt47MyVMKQ1hGMPZYpvCwYibiEE1bhANh1KV1Vei/4oApLO1v/MlDmGtwn5J/LYmc
0M6/aOLZ6/JMDNAR316iHNr74bJUg0L8DhrBNCK4c+vKPmytVHVVP1Gt7zszR8MrxT+tCkDIPr5i
tJg5PfwGEz/Fj+HZzgAqqwz1zomZIBsP/PFhqKlx+zP+VNWz0kz2bZUn85hDe+KEKyqZmkpQJ9x8
BLVqH8UF7T0voh5RnMVKxraytRMQqV8j4ByVpccRhMxtfmPxm8QWL5tHfp8X64++p6AAcx0/aXpA
nD+eruPhYHrqsZ9+wUZvy/ua/K8oWO50horQ6PL1Z0unmx8zgjAqiyCjMxHGS115lJsuwYHlZGO3
/zKOp9t4NVovgdrcNuJ+ctMSaAVVArYoPGNG8ElnVK6Er5m1qD/PI9huAb5pC8sOl/X25bnokK20
WdI+nGgeQyBvqNxpR0WDd9RRJESV8Kb3eoWkUw6XU0YtX9JRzT9BBdH/M4yWnZGMGv8leXznanRJ
36y7rViLfZ3KDAXURFCWoX86VmUGByOjiNooViZ7hms3hO4DRoEehykwe8038LCK4xeFUEozH3GV
qJsouMBHoxp+qb8p2iNmDOdRpecwYPyrdTzJx6PuaFvnBi/LEdkXOOtKYYTHBFm018dcM99vpu0A
JaRLiXO8XdxHJ+g+6WTt4cesnT1FgiHGaJzJAyO5g3Cavg0npRI13IoLiyBBkVSgrND5KRPFJFIh
iK6K5TBTu8Iw/FR/dpV0llfBHc1hBIQcy2Fj+bJ3/Tn5Likcb1ZUqzB4LG7vztKxMGrwODVjbUl+
O8E5jw1hnxCEn8H8buQ726gzR/uGnE40P93g0ZI9khdc4i9c+em5ehyHl6eg9v8S1TMtpA5VPHfL
U5dCAgr36uyRbAuBFtjzZkmkHgSaX9BEB1WgUA0g7lopN7X7lN2CVa37G5T0US2gJ4quK8O+ou8I
pueUGwK/ixoXdnabI4eoYYpwisVMbWjCoAmOPOX6tN3DBsV6filAr9CkCzrAS1aLkcqsGTr9biwZ
u/w2lB26YhnNLi0fvH44Z45AEPLf1qFV4JJWVbQ539v2JTfa7ps6jPoaGLrxcBs13dF7QWO1HUb9
yMgSP4ObLD5F1v1cDbUKkIiwFPZR8u2scCYo89tP4jdDDqRmWFPlreh+uYN/VsL81Jysor7XOjKi
FG2lZPHxvo/1p9i4Ixjwta41uvkBIKWcH6bO9ck5zOnZwjy79NIGYQ23ahnfuSc7+s0QEZJNPjZK
00ccm2lxBxPsASlI4urud9XamIlnP01nXCqvGHkPZK8LNgt9eUdavqB/vb4S6KJ814EgpMLyNAtM
HvGQVgynDNEo2vLXhEcgo3XhUFiNQKmO5HhY8W72rspFYjKWcvNTyOrNYWPlFwopbvXg5ZObbWr+
qDP4VrDCV9bVclgQUnTYXitJeytMAQw6rerBaZTP8gwBs6mZJGrPwc5cCPcs5hySZoGPxT3CvK18
Ulw6SztMNmFVoYxsmhaW2KP28hCYFpISMnPj8YZDVUy2biMFBB9Me76+bB52B2OX4V3qU0VqHk6z
pGd5ylNJI+HUoAM9JGZDuUyqi1tmCXDnvWIlyaa7XvdTulaP85jdT0M1xpjniMHxPMwDL2O+odns
yorGI41xwEaW1aFM7CL1YICMxpm3LT4zV5G/2usx5bwlCauXu9z9BA1eBHjGWQEGO3oQ+HnEF/FE
+Zn6lFXvbLej3dNZxuEWUb3B2i5FygnCPZBZbDRv/8esEWKTqGrxToIKa1pPKJRGaCyCrTX9U1c8
8cyDEX5ciuVvx75I9sz3vN3DQgoYeoEbapOxRYErSN9bF/j1eO6ysqVvPcX5AtihyDw40eg6xmsI
xjKhllG7LiqIAwell6Ye7vRZqrOrh/AQ8deQcb/AKyhF2g7xzM311ik6I5GvQys/8UwKKa90nQPB
ay2c7DUQclpBBXhx6F2w6aeE2KGfHnY6QKWfX8CNDb6zC8zoarts0lW/8V/Mjo+Jf92LZril4w2e
rNXnubjrFAco8CbSilmWEmbAR/LWKTzpiem8skJaw6fvci1tGKWHlCWRubz/llmNBRdlSZVeUYn2
w5h3AoImeY1dBY7+aV2ziXbGSlXhOD/xMk8m0Izg39k9tHe0kxroU7pGkP1ozqwWpmqcDWllGOSa
wKLbJ2rgE8DveZBZzpmbWCt82BIUqGlDK4pabluWXHJWq95IVdOOliyGjennvfRfiKnU+zZLLr2a
Yrgas6tp+l9Wec9Lk4IV3T7DLf6UAyXqp2s/dOYJVO/cAHKGRpo1Cm04fdddA2g7etN6q4s5C1f8
g5K0r3fK8TwH0qVg/gd/PXTOD1WFlXBSoE+7TV+6xobUenTo0Hty8Hhw0DN3Ormc2315+lzRtOd7
wqAF8Kk83E+Sa5cqZ96n84POILmTYea3XvjDkfIIan1nLUo0koEHScgLUhgnZ9b5d234KobFJNat
cH69WycyM+T+jpF9U1FlGYKEb491+BJIF17KbUGPrRriXMLiRuN140YIIMw4DQMNv3IC0u08sQET
CbiMXNrCGo7aiGlCXbrMSLmJCoY49P5sOGdS/YnfpVnM1Bd71qrk7nWQ0LPUErfEoyvCq0ZXwt/3
qRCIAHelOCV1u/zG+ywqNUTonMyGC7pdf9dEXAFSSmw2l8oEMGXwf3TBtGuG+93NN0GoMhqwiF+F
EZA9/VaTNK96fkqBpQrzDUhM/hPjwl8prKkOzlKtShbfg0B/19FAU0Ul61tKzcWoaxI1qweAQhUj
qIhj9HiKEF/daZrFjoCEO0rYCbEMFqlA2ezC5sOXGotTcxDGJgA9hkxrxJPa0da+ZQFf1fT9EQJt
jb2jSTujm8iQhaczVn4gaCCZXLcoR64M09jHe/DDMSevwHW/gljTYw2keqIbNsbuwqtzTH2ZL1Q2
yCMoKyJTdpbPTNiQiFyPu3wtKIuL4WKCoAtR+fWVED3CsL+3KQW1+tkINl6g9yC2U1RjqdAlzJ8q
NpedKNQhvmy7FmmPorSSCEEmzdiWGBH+LGJd/1k6SmbmC7rEw3ptoBkTvIRtXkdDsYzFhsUK1k1t
01G/DzIUFXt0rRrqH9NG7ka+BN/wLvo2xB8BnDTBo2sYDc08hodEuKZCoi/O29d5K5qnzx1q9e8I
NqhuHrs6quxx9Dbf4E7WEob26IOrBS8kQFFmIOgJYDMerX8Rly51Ri3JamzYZ/27c5e1djEZ29/S
Zl78cpsxA3MamteX+9KWC79TuUxxUxehHoDHTfzKYXLaGQMDjnioBmC4bVUgKKl0ccDlTcH2oOWO
GKjCMjt4Nh73THY7+geFuidNrNN7Hav1akIS9x1UfPm/MfSeGkgLYphCGHM8sYGLTp0/GQ6cS+mP
6UMoU0yLXa7snkUq0hbMqo8C9KOFgszfdO1VdOr8M6C//YSofbt0oEhEDjOAS09MCcz4Wnvoy2ij
pbttXnkAErRAMkohhn7seW18AymqP+3nU58ifqEIZaCrFvr8Ntn3bX8zfwoVgO110bpM2rL7vNgX
zwHA2OnSeuEi85Y9P2St5FOqjgB39CMX47tX8tak9O/H+/THIZ9/5SNtz1QuMJI/dk8WQSBxTmKv
6mXUz/zhzZE6L+rlcFWCQD/5a0P7eDT2bMY0b6v/4TVRYJ9oye5JuVvL3mmaSAOzYiKgz2hBvHBN
JiLVn8PSabv4NsF3r+j54fLsI9fxzUE1oABQv+PzsLt8CecCU5xu/ZDMSf1hrRladCL85IGoJg2h
ZedBwZzCHsjr7/q/XPiIyw0OZTSukogzM1YUA82OExYH37miXwR3Mk2t8rpawto594D/IOnztXV/
euRJBUfrvbHWNO7ThmEecCyVSGLQhlBA/24CufplE2wb4KnTqaMlPfqQIzzi5ooI9IOpdTsnNeKD
hF206qI043YgtGJDDIUOhL1Y0DL75SBQtNIDIVyTMAPHiJhjy5JO1DOXYelVtbG0nEs4CgLSbYV4
QQgf/xZhOBl0ynVcaq3a+kPJS+PdzUMZKq9vv0oKImnLIbaQlObhmNiFMMEXuoDFH3k3und/4RgT
M6dSp8iE1aTRrjHF4WWlCs2yjBGMHbjxXIxJpf6oVQRT0EgH6gWaMeiSRVgFd6r1ZK1865gkvnoc
pNSPtoUQ7xS3NLJYRix3gEUmwNsCyA5JVw/RNZrIAk1/KW3yjvuuD4hBn8KBTyJ67i0v5O6csk7N
NNcs1CIb2UFdhnBcjv/NT/oHkvPXKDKmdy8Naco+RiUBIlx1sEodKzFI1/O69Dpvscr9tniJq7eM
jzZTrABinMBWt0tU4twbh74GJk9qd8gVMihlGkx4ZJHctM5LtCKrlwBuRPiT0Dc4dpufo6c/b0FV
Z6ix1v+aMk1PJf/hhi7khnRHZQnhWeDL9up8fl/zCLy233qkhd8hHTfR/9Vqhiy6GJInHmtO+58S
PK6ewDYbvlY+zW8cWoORKpW6hw5ojdRXwDIgbGAKk4Idx4eJwV2+qrOh+cyrzFetsKLgKOf6z81W
ONK0IJKWJk/+64vw3GWTvTWa13wuVD/hlWC4UP8i9aRAXOKEV9UNM7pbDQjoUmIubhigSz+8IG2E
jUBlPINGv3tIjhjq7Iee/i8iNXqtHPaV5DVHL5mPY60Dam3/yWL9dy6DhHg2VoBYLA2UNswWVJfU
XFCGO//FscNH3NgZ4wYHs5o34Gx1ftisFR1mGhSBIc2VjlPSBllHxB/tW/LulTpZ61ouKXSL33VW
B1PK9mnON9Wq/Rq/HaNrLqdPXWzb072G/7p4XUz8DBtcvV2cnRn+fiTsvRvAHCPAlKev9exepujA
KiiZrFy0G5htHIQh7A2R9sBNSak0ojl4+ZcFDnKvyOppPYP+bTHCjOEdv2pJeXayG1OYJt2ftuUD
ExL5Nb+Hj8RMXXfeEZsXuk78cggzn6kgE6Ssgghg8I/EZ4FBqKQYUZpB0mNIxg184MCXQPX5/egT
mf+Fz49Hx+44Atv4mqOGQR7h9TOnvtDSdN4T2KEgXz9ycsmU/B/qXDww42Jx7cdlVC+vrVnGHNDt
+64OcDr9QXKKnNddkQMVCJoUO04QBemUKW410iIRqY0Z97x3tByFmLKoQhUOgxMT1DAxLq1I9/Oy
1xEq5ZAxEpvXA3mxcNeN6ZXxqPmjsD341K0BXWckc+9aYSsYpssKyN0lPvosI/YxLZDJohFsevuE
SAi4IW1ytLVO8wmSsAafomDtNCmPmgEfV2lc5wUmNpoaeWZpYAEF6DE4NIYidTzV48tlRSyM/SzC
IpqWo/XTQ95vdh7RlMMtoUsfmsFpNX/i/yOuTui1EE8+uirORqXbnsg1WohFTps9B/5em/xOiDPJ
ZSHX4CjM/qWH2g3DobxRxE20G5kwhGs7Ri6/ZBz3XYKM+SfZj0yTlGnernUw8+FoM8IkukAyfzp3
2XFyDpgif6ZnDHYWXESI9jvk3aUEsoz1sfOJFCTYxPDmmO3IThNteVqAgVs4GxA2JC4KEtWAjvsR
D/95M9eHqEKnoMVJZVnlLz2UIGLxQalZsR26plL443qb2j9lPz1OY22wGWzp6Hr64Q8SdV8J7qLS
C0B4+0o9uBaNN0A4DUMf7fq/qnllDWfr9/8A46zjSqXVXvPL5G4w4wzm97j++hdB8AAxvPUvZ5Og
29N/f/XeruGyyBwdJhhhTw9/d7btvLnLGrbV9G264nL8AeS3IH4y6ssNEw6ogvuxtNSR2Ywu0kHN
aedAUzTqOOJifxiEEGH1VzJDthfs8bO3eo/RnNxLMoRBRiQG+ZRIJlkruJTFlW5+yQKsElpoeFbB
NN1vnZSpImUnS1F1SjEbwouQ4JFaFpJVuEjm1ioAVdi/nDXcO9ORbKB0MtakgIiiiDL97Ny9JIDw
0xDEBJPzUmlHtym1XHzjwKUCV5dj7Na8QQP5PiPAwlu+sg73N7tLH3ufzQiZJRShWVwd+18fwBXa
CYG0vkVSI2Yc6GGX4gifXdXuH2jGEoGyg4yRkQa2TgukGrvKjO6wsopjlJpznLLrSR4GvFdjZJ+W
QW1C/xajvT3Da4bfblp79LsUjip+bJgaXBBtFIpc/aGTnzd/fyr2OZxo/rE3xn06AE5xg/0VyYBI
yM5db4x9o+581oyuzTprZ1DRjDadgceVj4UFDM3OiAbwkGZcV0e8i7jBMVzXZoiU5B8lSxqLM6hc
+knmjW2nYIFxK5pAQ/3tM+MrEr+pVE8fPbElsWF+08H2n/E1OYQ3N08umCrc3Y5SOF5wqS5+LY7F
a3nug1y5NCnf8RGkX+qJTXCz7JIj31SaEIOL9APubjVhTtv2onzlhxcAYgMTIsonOsJTty0F14SB
P8BR0KHTVISzRrcvP9XfjlM6lC4r8q+oUT/jG/WarhyK8UByxY698/t/4a6khYB3czhyXKdDNMAw
unLe9HKWh9GQw4LeNQpprMxjejlffiWvH9+0MNTJOWeCVIU6HKClv7K0ImuWuT4lZf1cEOViPpuO
EK69/SRbcqoqb9oZZzzkiqz9/mm3EwD4HxaTmhfIBeh7dNpUekqgHbRprpnhO5FMPsjaw30fSz1+
zvJxdqZ7Erwf3cyVh5GPQ3HWQRXK4X4qHL03990YUi6sII5NEKNGINj1Y7Hb98T/ja9CUg0cOi8o
Cr3SsCSMrja1+YhC6vP5HWCRw22koiB0q9f9EGjSmTUF9O1u9xqsQduDBNe5ObQpgvOUe8QiDPeu
4H+5QlGO3J5+77g01b2/H1PG2tk4LJG5L5R4lU02LUuUzvCmG/I4LyJHXjxEENgQHmJCS5H88Byy
bNrAVVbvD2MR3m9+MQcxXDU/LKCNxJ34iSUvCpxOE9HUyyuUZTCE/VpvcOrEXr9kqt2z9kasKm3N
HiGnwZ81qKaP4ookdPWkl03mHnv+QZ60Q46Ob65VdB8h+GdE+cOKlhlm/W1KvoCpHyd/xQh7gns2
rx9uwOXVhWT5oq86NokleANHQoqLh35x/NNRkCQMjW2/XYdg2lYI9DNJ4LJ5yihETwVPeF/EtXYs
VoR71CTWA5yiYeATefVmuPXprDBEvwDW2VuZ53dvK7MF52BNzW2KPEZnTkEGMtoYQWbRxRp2nrEb
OUh368zpCEQNVOg1ezKDMdQpRh9qgm4O0pgpsYJudDJPFR5pV0InlacMFpw1nSnarAYMtUaT4Iy8
LtExQNY84KKJYEsOdguR5HnNCVpEVNAFAwlTUiUb72rhE1Mhih3gi1Xn3inOFfgvo6PsPLHxVBQ+
ry6qeXHDCj/LE48cO7AgjLwduRXewGxFq4hFoSWFbjBK/zHlSoN+L3/3mMq0I51/vg3pNuDG0QX6
5TlDoMqjBDHC3m1JH/DRrD/POmppVPNoQkIaz1GiMaoqQZbjIzH841co04RhscFgJPIUiCqpttu1
LL698I4D761T4qAYNtlwa+4r8+NxzKSVvcXVWw04GAEo50wQ/TXLQaxuDQtuphegdx1BON6SZxrp
lfWx4/YF0Q1MGuHgkA+mrEhmSNJPEjlyLH+A09PgYyxA3hqGi5iE9g2QiAG4tamHUF6Ncd0rzrZr
ael5V5wkresliuM9+NsUPIRd7gfOgY75SLMEzebFLfDhWv+IbIOyjfTNkRalEhEl8fI1cfRDI6lf
xDq8KU4fl9yLcrYmSGr3DUR/TeLvRicCgdyf9qSZSpWVoWPCnYJfrJLZ8viQO8T8Su5NeiVEGZA0
9LBf2sYwCIvqGQqCEIgNFPVIygfsyGK2UvDd+46ERb+yj2wu/3hlSg9MMjWo+3BIjaKetPLwgkMJ
PBwrTc1KCJGcRpPUHj+vXdECYB2Ke0FlkLJtDY0Q/OhhkKDpVBm7zuTzBZ8rCi214l6A/1/bO6xe
EBnff5FwhEf+/I8+vwgPdWIlZBNGT/kRXjl21q5G5z8SDzVi/MXIMhLxtwh021j5fFkpRt44FlDd
Z91/5b1yZA5ZofDd8CBOBYhm5TEND4XMd/wkS3sI1svq8mBpMNXPhF1xO6hSf5RUXoyxpNosrdrD
30xkjdyu3Qz6/5uiruPehBNk0gwtCEQSXR2NDXsnlaLGxPdvjcvRfDIR1nDOxNUbDHfOMfv568Rc
kt7aa6ltW0Mapf75+DUXD1oqu4R1tiiwBvIkQ3O2h4QLEleH6ltoA1UveOKQ211FG5lJit1DRC/p
lb3lKotxwUZF8aSGxMxH5KkJ5B8ufu/SLSjjpqc9gRjErJBxDBxI6YNoXlDpEU3mfYqMUEPMtQ94
tApwKmdIwJWlN/ZeO36Nj4fc3LqKOFJi+GTwXQBU3zR9TWo2zf95+iL0qJUKrQuFcK7+uAxIv+Z1
SPbmPzA7s/v3iE62h/jtqDlM7m/+RQtdg10yA1qZW9LDCEsUbWOQHIPgQlt0GXiMAbpIeUYYW5rN
drQ4UO/KCDt/er/bUa6ITCpk24OrW0+qA205MxQXXSbmTMVEQqMXVyYENXg+Frzhvp6i36Shjtr2
2kmrLobNAjGAwR6q9NimgCMOE/R06ttkVRwuIRUZ5uS8YbZfp85ZhS37eamgZto1VjrTi9/1Oa30
B9QQPaJ56hM7PA6zj9nqvc9+k4fBoi2hAKXO+1cVRTscK0QFc4LpGgOtsdt64rQhqwFFqnankFEw
hVWWDULKQcP+RNWSu09SX5ScnMj2xrWSUhTIT/OlScaQndy0kUXaTyAfX08y86bFvlSC6URw+HtT
zDe6a387oAtfzxd1xEIy9TfLwcckJsmY9+HROvlXz5zVTT9mW/F57m/ng5uao5f6u77FBm528RIA
+vFuuHF/jL+8MuAMSH97bdGZWye52eMEZ+8fevzk/bpSGIvnpbc4D993VfYstjgT2yMNZdN8Bvab
eJ7gnicD+5iIQg7aJ1Unp7sGBoUCY0k+8q10iWyBJu9qbh5jvy+15P4ciQUo8O6/CRUKjmJO7DxI
UhzxdBoKL8CvGNPQmmxh4xNL3z3dyWVyq4B5pOCd/qtGlqpY59TPMRLs8m/SGX3zfyfvV9qhrOYC
Ddycy7qz9F5i+jfa3qufMn9m5Ia3Eejop4aN3zLHrfGbLLJCWWYSDc7FvdtMiStPNXze7rS1qwm6
az76F52ZjgAspZZEaTvy0Goantt+CsuT+CWQpsndXAum9rZ9JVI6aHWeh8lFrojyFmnxqd0+57o8
RmFbDKc1PEH4I6iS+TBJIbTcX02L5j5UOlx/Fc2PzlYK5b6n8e8ylPvxps0zX1/cqOUlAoGoYT8M
9e1QyACYF7yz/9r0bPqOoQlT1uOLjP2Z+vye/zeE9RTNqF0priDtReXHnr3wJ4eOPwdwv5tNBt/8
1NbgwnBFnd1zvxtQOLeeAzaAs6oi/3uS8crtrL/AoxaIWfxn57fCaWLDiw2lJObG4N62pvASpmzW
kCTvPQv99tr7BKM7A4V5wvowRMbc6R313r3lblo4bPS3Jm9IWE2jny8thxshJcdVIWIy+VWvywZW
hKxYl90EB2A/ceZ/ULlxsbK40HDkem8cVr+gVqKbppuDWTfm2TbnYloyLcTicv6fgstfuVPcBiNw
KcO6lAyF5ib0zNl5sHOegbiKUNq06IwDq2g137EnFPRyb4048il35ii3Bl1qnigU3YYeyo0qhdBt
lXnpJR1JkAkfAHKQr9EaWNGP7Rx323bA4AZUAU2gEy5QKpgTYgVBuuXFWf2iWiQcDyyW58ItmoIg
GHvf8B1xiiXcf2VF071BLpEA5K+uZGTTsHfoAcV2ovqu4yADTDLKk8VAbB3Egphi5D8M6zjafzv5
tQTmNKywJzaE3EdZKta3ni0Agss1D+xXa3a4/rcdE1UMTevac5GrmdwM6bCl6IQQnBKy4VlxpkFO
x7lR8Up62yhNse9kv+mwYaASZlmzqSMhF/4oK13yXFmZUMfkTDfSO54HKpP5IAMjWbxvDjmzo3J3
CqKpq2+wRJCdw5L9yqeqHkhXPwv/1L6/LdxI/hKEb0zyqN+6mYRAhBTUbjVQvPLJIEYK0cvXoi6u
KZ7xjAXcFoA8yLXvdd3Qm8UkhwNvld37UdnAImZ+Okwc5Ur6G7u0LcHPFE1Xv1debkrTlbxzFA4W
ocwl6WOlQ3RXzUUtlJGufGVr2ODsE8zF6vYaB4HN8OdryLrvrT0t+P3UXD3iv2Th37pe5qbk7jmh
ECbOspXguw+1rkVV1stmAx9uqGcD0BAKCuW5u82y7Q5N9oQySjpDFIV4UMb9tVpxJ6nCMdycG+I8
jPuzALTie9eFggQtlkuknInazI4m302KuQc2pgxO6+W3oNYZhTPqVLmYb/kWs9mzAjaW/9XANrTl
gpUZc2wuM34sePWWCP04Yzyp+1jkzcntsB+HVUFwTrzT3foD8YSfjlg8s8kwKOkJGIeBzzsEx/9J
J0xwtDAmr1tp84/X2h51tyxpeXgQh3wyAp9hEarV7LNC6n2/6PmjPDJZeh4wnUbpOoVLXS4vpFrZ
R9fPdlbBgFKqrnPnSg4/UK5mDNhz/MEiiADaweieoYZBBY4Q699CGVHWzH5PL+uQMhWSw951Xwv2
rhEuXEwsSzbrv+pNV2IJr+V8Hb5vnOsCyA4ksipx05v44YA714E3BJX8JUUXn/6Gku4+wqmx9zef
0yTzuL9PBQwVhFfSm3ppBZp165dlnFCh8ixyWJ6pjHX/vphfI2bVCYTOWMvHI4+C9+Mt3Y52c/zx
AR+bIBLtac9aDNVJ7nET31RteD5p5hcpDqUdBj+5xBT8VIo9G5BpMyRClv3hRZTyk7ugi3IcZ2J9
YQ9ZAwlC+dw0VhlQsMVuBDXZ0Y833Dx0Sw72kS7Gvlv9vVN4LZ9LUOPOoLdTsw1ZjB3krotaD+qQ
Ewwpt9YHjvqVQTJLs1YienpS76I2dNOOI5xAxjxVRxScBXSC0aD/BQJPyDeXMG9qe7CbAV6xb/Md
+SARcnxINdWHKK2dQgQcjhmJmH1P3YLjJMswn9dkFYAd/uJOi+LzgFkv7aAQT3mAgEq+EiMTcm18
bxq8c85vQ6CJkWWfnd9vFDGe3zwUW+BJThQmH/0MXqgaGln5PB9WbaTBA/yb9U+MBYeChkVmM8H6
WZR07g2LJkRLFIqjWtYXGalcojgoujuwG4nqtUjF6ymY3Q+49Jl5pJ5MY6wR1KjTZMDXg452HHBF
MN/KTlP5hF42pKVDWv5y+KIhMJRqAXm2IGnq3hxuP1wwVsXQA33ClY7t/jfloH8e4wjiujdqXO+f
8NCldcg5JZAPiqwvFM05zZvKlg3FYmRzuUj8y9K6HN74NjVpc9UGPwvrfrdJ1qcEr+9J2qEDLW76
VtJL2B7o1sWBHfc78GMR1nrg5fTjgvCnJoTgX4WCRypQv6gZdTCm6fKbMPKx4eCu/E3/Daxfr0Kz
oKwlGu5Bzou1WfQa/H6Ev5dtYxAy50h+/11u12KvteIlajCOdSAtXwfOdNvXk+MyVbqhmyFR9aCY
hfo7PO3Spxg1apVq2BBV93aUUWrxk84NivniQXJwD9gn/A4uBIDi1e0YkKYKBVj8krwKpxYepvcV
hv/l71czS3Rk/08JX5WPwfzFSOgQCiLQKj9ha1n111TdtaixpubKne4dqdlXuwljxG6VfYqGGhKU
twcVJCYWQtYSw5GAjM0Vg9S3NPSoMU+UTTKxUmaToPg9ov+BszkwGWTgAMzyvu4MGTzszEgIPg0L
bkYOv3xBzPuiRs0ZYBFG5neUPxBNG5waPPb79ed8LfiduKx8/9NMFR8h9UtFSkWLwDKhIxQ6Ev4R
+jyHgnS7H0C3dLVChbm+OIPfK2FgJ1NMzG/KxEdMBodvL+b1R08TNnCktNejeG48ZSLfbO3WXtuB
oUkwB5yyOGDUOTkDyBxNpX+bk+/PAAFaUAEHm68uJqXtsDxIAJAoCyIN9tyoxD1SmFkjxaHd106t
NVMKBlUjOuxbDRB2DCJMByVkOm3GE0wt74Vw6DCNVSAWbhxS4IXIR1rVVk3zMW5hxprBSLlm+Izz
dxV4SagRSKgiqI5YMn2s9KqX32teYH425rdvg4u6SHZva4af5ba6Lj8gcq0e9wF7X6kReJLAkI2S
vS9HvnSCdsWn9wis1gosxzKjexSmrQ6OJflYaU2KqoLk/wbQF2aJvSImi6k2KdqOijDDBXRnj4ys
auhoV851bC+luTxL2OoQ4msEoBTfQsQ+KblBbODszE2ghu9myusd65o2aioto4u0Uk1H3FE4vNf2
utY149ms6JuGjgnrENMs/6p10UyNT2cvmbeFuGlwdvTieCE/iOpBnxUwlxSXTuQzSIBkFhcsUcm4
cwje+npqm/4oWlVfgQcEDlN+1/YpXIq0UlEkULsyxgaPlxswQOcOcWwCRpfmBya+jdtj9lYXJx0n
QBJeVoJO5BPBAn+BxD51XLFdPOgbNCTFnLUvC+WnzpXLsiQuIYAmPJZw6jbodHYsTXdyJ5X3EbM+
Wou47dS9VBRVTwZkGRcoPYfaf6eaL2qt4+ieJReD6xL9D+t93Caw2mqehcuzLqKzuT5PlqGT9z7d
SR5sEf6Xp8EM8jFQPtVP4pCjXhX4X8ks3+nPEoIfF+WMgM2gztcLp6OXC+m8YMnsLLLRxvPJQnZN
GDoxY+pbiYFlZtn5oQQzdp8N545yrkVhwJmPWFE3J1xW/86dLJb77HDpS3CUOzpgXZMdPyFYtcSY
Cf3mGKmPq5y+kSIRKYPuUJXMaj0lq7TBgkAuZkaU5m9w5CsNG6X2cxXF+4I8ErSsNMPoJzGabGRJ
zZt4Pmjy1t/Emvd49QqK0yV+34+GBTPHhX80UPQ5KQP5ROxCs8d1NnjY/jKOR+9a7q6spDi1ZkaJ
c9/caTm+tSIrPGRUTUdy06MbWArlpvCUxBpwB4/L5TEImxBkOjw0x5xE9lIZzEEEP5KSAZGrDomV
EeB9v0dHBOcobXfOm6QXlpdrgj9ypImnXVcQELF+o1soTqoOM3pKiHF/41Zr33k6sF9OgmG8wHkK
0BERrvEbMrSU1wO02xoDO7+b9RIulCBKdGWHNXnExc+DllqqlDDBrM9FudyMHnv7XPHbxHwZ1tB2
n9uemMXnSwCgeHh30rgQWGslcYsnj5iX0CRBy6/2nMkYFOQsWGIu4aGtsicJIq6sRNjLPwRjE7wI
IY2uv+o2fYhCudrOsVEi/yzTu9233z0v//mC7nB6yrueP6smdvgNhbOTJMwxlwqzGRETFZeydhmv
lT8kjCE9sZ8n4Ay/H7UlOoF7AXeMsauHfAjqWeu3+Fv8pYJI8921IPJ7FVlgba0n9UqCLPgYRDVp
A6z00DTrWq+c4CMe8FUqTH97YzyunBQgmuCZ0C9Jy6ArHCn9evxq78rfmQTNzR0vnzwVUKCba7/m
AULMOaPnyGF0d6S4LzvNkZ0Vglo0JVjcLJq9PxVCJFh6y+TwRZ22L1QEko7mqAylY5FjVtpnHfWI
cPDFhoZjK6UQLwkINDulPK4jgK/0F7YYrdEV6u5ibtmfqXjooim3FLLe1dShaOdXusBK47G4dSle
ZllEE8mhQPzbESSszDHeQt9cWF/7Hmr5gIVOFf5r7/ey2proGnyKz2tSrNyoZZyditt+QtsV971Z
BnOJo9GYbkIWMWIqPMtX7qBeBTs4lSyk/upuDPyheUMi7b+m3hhgeVtIz8sYJ2uzoBJCih2QoLm+
7gbfRcf4i3ifvZX1r9p90ByyZF5R+KXgy79fKp5tze0wWV1fk391kQEiNLD6ohSg6clOKVOBbrTD
ahdZJf+EMrQ3koX8kHqPpw6uiKMA0u3GPlHuMElqdl2t+BoftPEvxlcXf4WGOiwwtn3Bx0dRlJ0g
fEnZrIjD3jH5VjrU7DZkMP3z3RC6M+TkM4QIJ+NJKHIkSsnf3sbsnLjVcfCZ1577mmKPOgo1+T8N
AHMEZR8+Cc84lDWn9gUHT2QyDAG/F1AJpdfpMx4Uk0OC42Fvu058PqnaCpf9Zb1gj25Dkk8GZWOb
feivfsOgq/YfOB9a7QtiOD8+q8EGMzaAv5qR4p4ofufX2JHfZWOkhSRgzKrBCbf76VxutYT35nGz
H9OYpiIZnB+lHLC/mwgolN9RqoapDAjx0AUR+G4cu2zH5i4SDW/mm75YtCQ6rImq0Nbbnf69X0NX
AJ/y9whzwbKeiSLmqQYQyPzTPMTCA2UodCN77WXfNXaPRpSBMl+YltOpSHLjZKQIgHC45KtAIIdQ
JHMLc3Xr2GVW4COt97jgYEHfVkZnAeBY64jMHPSwbu6DyVv0qps5ldxwyahcjbT9wS/eOADBOmbv
57HEVXfC1gbrclJEGfejlnNzYnx6EHdpryj5aiBVFg4Zq+wjfAUEhcUNIJ7WGhS1zwwUDh6fVYXv
lbpKPS76EUJibhuQw3MNTzW7BiPilEFkN6K3uSTecQZiwbnv7UOtt+e1H0gunsvGWQDHUEZCWR+I
NHv+II9zq9+ibYx7aAcR0BptMDZcz1LEpI08ByU6eKgLq438Rtw6haYitbFXmvkeXxX4QUt7ah7P
mnrs0g+KzWCvkNV67dVpq35asygwjj0W4uO7Ylh6XULm3TuBvIhi7xXFVldRrT1Z/bIwRlb7gHUO
IKXFAh5nLnXvv2oYcMg79MWdRd8cHgwMBb7dgOz0d05laNvGq9PGdBXIjGEzqNeFXQb3hX6aAaNG
ZuQO7BgLv5ibtNgAB8mMwUzai9keVvRGIB0rw4VXHqHDvXjrAKNzOt8sPDE0iW4nTxM7lZ+s5mbU
3GTRpUSU3R/j8LxFoKHYiaBcPBdrQNzrvqBLasxqTTU2hwpnR6sKfqBwobaenPUEzG498Rh22fn+
luBmY+UFPGspHDTgX6FiDXoOXSUIlKT45wUkOapR6CoqYeirom/v6loFbE+kE9Rici1adslsqbuY
jDcGBBAI5V5Pbo3gNWgeSGTUgqPCyMb6x7XBQphTniIfK0tcd6WfUcnxhEXvNapyCzVQJVXaXRKC
dvoOM3F1oik2N05z7Y8ahPvwWbzeEiJiyqjzzr9E66TjxZcnW53yJXg6Z5HT1vo6Ufg+w1Z9P5P0
dxTA0T4a4QI6ByKsJbBiYzMcpd82JJ5d1CcuLovsTXjtGNauNQLyNledtyOi/7IsxpoTePC1j83n
5rJPNQrzcB3lCZVokEGoJiN5X0u+JlrYjCdj2rqnWXFlQkJ7oYtPmZsVUoNTpQ+f37uIdooreKbl
gIw0Z4MYD0y0f1OCrVk4LreWaHRylF0gBSb32ZxSG7HUz0P3jTJPUjRN9XJb1uyrAvJwlyOHCr09
khrfUdw/pEXlXTYKyoI5OIQpfLwLjic7qWXACmIXm+lmCdoufxP5COD4oNeRbohP1h01VO8jpfhq
EfJxxYSeAJaY53HDXAbYwsZ6E53ieMi1l5tn08IHb+s2xHjy+/1XRXz9vBuQ6saI6Vgrm0+sa5N/
YMc+Jj1pyEPSGv7DvDyllKWOh6WJxJsh0DVS7WOCkklH29G/cCZtXKSKsBKKOrE19jglBuegKAaD
65xpaLjtVpVBHSxjlgUmKhRw2+kqLjhJc5HUgUsiTlQRi/9CseWPyFvzFNWS88RKZ2gZU+9HVfYA
vLB1+1INaI8t81wHYw9DJ9rmARrUFjbkFyAZhQsF5nuOy4UUUwVfOV4tGpGTm37xwt1lOlm47LTe
39LvtUp8k3g6j5rAPs9vSs46v2IGuqpTXyciawopiIMS/RpIRBIijZZ021p7JKYwh9BafevfWBOo
TFF2V8jjhf3BLkdJDxb2Y0qFqhrb0+WmTo8t/s00+P0MVisPZ1XXVwtSzUzRe2OJFZjpvHqOCuqZ
EHpxDzWCsmE5PqJvmZn1Vt0W0ETJXqohQ2Zr1ZcrpR8/E6DfnzfOVX6EqQ1h2QTPLgu73Pq6s78h
yXbwm+b4ZzV182t3iaNIfD/ozmyb2tkHwug8JLKQQ6lqsCc1KDvDKuX+xvC/yVy5GDTYMvSpRGDV
Ewa+Ztl9asjw9ow8ho2aHrxVkK6ZAJCS2o6MDlSZHHJE918H3hzejehU1i68JWvaoI9SrnKUiSbT
NULw7Hb7CieY4lGzcR8zbG7Bjh9jip/m5OPnMR/DzJpCUd06z/3sUZvax3XLjbRouHYqA5xxiJ+1
RPzCllq4MCjCbtt3WHaGe8izcldBsXrSn/cxyTiXb/cxqToZmaKDgu3iDrTIwiH58Llf6H24ukgk
CbGm2eqjXVu6LJJK+6iT9oR/Y46qG2nJCQeUWz1DqEUvjIVo6CFDYjPaICtT8qNS8r9yeH5jY/iS
na5Zuq9qdSpoEPxYgdgQ+nNqVZ3wowvB6tG9F7AghWnUYjbRdzCU6/OVj4c01bqNX/ZisLPJhdGe
q/l9ioByOrof01SxmKDs8MAapkdpo6bsDUzABWnnHYYdFxtjHTic+syAY5O8bHJNl/KkXxmaMGMd
wZ64vDP3W+8Ekjs+WYLzDCKbFNIkXJM9XwnGPMC0h8KBvJDFCYlmE9KJ50FE2dUJXcLAppGglv9Q
Tp1YXxCwrlHqaitrZlGENEVemZc/O1PXgGYEYWyaYQE4cCyDcIBDbxWceE06donaOHV01lY9lX9w
CFTkjuGTUCx8KfrSfBSqysNzl9bg2GPo1kiLeU3bXdlEqRvRpkziRhY9yOrm4iF40wZ8LLuEAtIC
ODjYhmPOLq8yLXr/TiyVOhU8Ex9kCC5jEry9rETmowIMqX6bcQf64/iTpnJ5+wMOWSNXB4DpuwLE
MS+Wp6Tpu14PCX6DaQcPO2SvU5JPVTM9juAAk0NJMpRVXdkl51jhPk7Eq/6ry+jgaj2MKlr6eZ6G
/gsu5DYWbwGvjrMlhDijxKRaBUONpsgsfI3XD7+9KVvgl8Zb/G1FwIHedxisnLegv5689V1ClPyg
DysepxvIH21G3Pox+o3upmLNER5hWXXAK/nwIBKkJD2HT9/HZ3PKKwM+x2jT8yi601VmMLK026l/
9SwumwOB5RTEHMbjiQqHvsB/NP1NybYw1kiR0oEGo2aDMETzSFO2O0VpvmNE4U/pszsZhMRgNvm4
XAnaet2jrn2tN9PFF5h/dxfGh3nF6BuBdFMjR/9Ol6qDXdEfs4sQwCY89KtFfq2yj2ZTUhaYRbKF
U7pDLUwaLjWC/f76qfWyqz8KCSzqGYqBH5cc7MvpVHXC27IN1XVrQ9xfv8W2h78ktugSrtsgq0a6
xzN1qmTRhJLsIM0p7XVEcvmHku9aXcyMZZBXowWS5CBNOLbaUXCh7trG/PbEpEi5x63UcFxS+L/L
D1L6l5xPAYdRtob8qRLvBs5xktuVylnGnmsnSabhX9wXBknDD3KvHnFm0GXgRa4rs29PutrsC2En
Vouc8SLeQPJEN2FXYl3Jnmxv5v2xhb2bV+0y14GWUFyVFa5lDNdimevjWlGkW+9GRBEaxNum0hRA
SsOruGvZfFP/sOKDkAXB70O0nIhK7MTc3qOTJgWTbLdDjdoxDrMDtF2Ev4yVve0pfPbxXSoY9MnU
3yZv1uZS6QdwDw8sh1iGoOTBm5K8HQ60NmCd3J2tRtV6v5r2Dod1Sy9+xe69o2VPA0b8fasLQyN+
07bHbEWWvOAPH3t00vjw/mi97q53j17EhcN2lZUirTANKxDn45qLxlFLl6Axm1LEfl8cs+yfo7gN
p7NCKjzhSQnXtfOSYUe9rqF6SDslOmikfqFr+E8WNvHrODJy4HNgvwybaPBvnSZMewE1JGtNeH5V
xoX0Am2LDpO1C79wiXKeOcAMlfQ3vvjp+LNHXkXOABIy2b451sQN//y3nQhtU6Z5VfvUHLMJ4Fhc
9lczbb+IWVZnFs1mINK4f0/hF1GSjI9rkiry3wzcUJarXmg6USRIRccFz162T4v4T9+WRg0s8OcY
VSM7U1t0yAEeOBYEfIuTdMFdHhz4cXPQSTU8+TEzM2fTy4w7dj2QAT5Zs6BH4SiIxXTMFYW0fXhg
4Dv6HRUiIXMdP6zBZ93fa64AM77ciYogRuuJhwQc0Nd8UyZBEVxcSm/NW9EbqmyNL6Fdn8riJs1t
DW/SisvqwoKYQoESO4PhqTiopsTjwVPnOavAp2NIsbCcezbOPO0Y6Age134gKHtjHFIcCRThrwss
v4qKayZP5viCLVaUZrrtU+GF4yn8mbjfkq+CfYyumnk5jVpaqmHupahDbYoRU9UkSFwacjKkpd5Z
6D+/inastpHjUmHyuUAVX0QhAbOTSGNc0kqiA24jtui8YlXjmmgi/3lH0FzbWlEk9hsDi8Cr4QMz
XL/4nMsB78tC3gm7x6ML0Lr1O7qW85g6gz7Y9ZbiVkh+Ol3wwpYgmBZ75ljwJ9RKftnVJqLHXbvX
XQiKxhc2Ww8GFIySnwDzHDp8DK7bUbOD6rsM5w5/XUbF+FRT0s3daUsa7jVNP05W04jOTPLH7pE+
3BV91IqEGjoxOwkdqQUabMOD4VhCA1lWTV3swplHVInBclSsJr5AmF5+mrgWmyDOt1eIVGj9Zt3N
6O4p5MhXJdrD6aUCOuWphndHDJcAB3gR9tGYhv5JwmGsS8s+TCaB0ccq25C/jk2E5+GTJYRIwz9K
1s061aZq04ptfLZ87A5U4j01RszmFTo8A2PWnkFWk2Zlh8OgPplFuLVNfBtMM8l2/7WAYCFVmdQ1
BbCovFzw3LRP4VuKc7D7JAclv/7j4K890B1JJRXz66KEEGX7p5olZep227ajN4tebuV+ONNfPLuo
QG1u6T/Xu1UFHiBN5haiDykfmWfj1a6sVfViIflm80dSe3+9St+8CSHgY8BNJ6juq982r4qHU3MB
+IMMChcCgAiWtpUQ0+VuRwlGOxAk7SViICeUs00lDW4fKW0e4nleijHJxAMyZFdWuWiQ1w1GCbcY
UtXe/6gKsZkWgHkNiih5LvHX3VDxNpnRUUGepng2pynM82iz3eBx4Bj+KjqjVZquBZJBRFh+2/Yq
rK/cP5O18HD+zJVXqipSAT0rs2WZqarwa5SstrLoVHAgT7j4MJEbSSDZZi7g+hfnP2/w6yJYgbG1
Fe4FLWR+2T1vGaqWOFGwlLOyAj2/7ZeUM3ME8i4TyjwZhptec2W+j87F+Bn91Im4R7+WZO4xJzdg
/0WdakKsmcUS4DOlDAsfdT9KfCDUxzZZYoVXxb/Tfdczd0N+KTtT3TYn7n33NEPFp9TwQMsyxPLv
XnRI5SsVLIxW/InzbGZu7GF3q+I89TKKyfQEatbsIprxoa56mmVr6Vj+sCbJhEeoz++WQcQ9A3l5
h0ng1GKAUEaw/nUV9p2r4odAgsAmvII7cYvLda+V9TsdbIj/1yxKThK58X8RUCagDqxxW9PBIe2q
V0+zu1jJxNS8w16Jcjq5Olu+rhin669dIMPzWS0tPvbmmCljh1Ch+/1RMv+Y8TgxjJd34hpXgdNJ
sv3Tl4ElDakF/3DSUOHZcCeZrXjDdiKDFN95QcvhaDwCEJNqXscx6FHdtg1wm3AUkrqiHDT6QS4u
nhXGqwMXzGAM9KAEJ3SIr8z7wbqyzj2ocBisjXAyt/Fn1JwiXh+lO1CLzjAWJhsupE+jeNr6SyVd
A1JZ4IzeAAMNb38orZb2ZDkQbsU/IsvgwwKNQceVeJmCbZMO08VQcyGBDN4bjz5T4Vk6Oj2q/rv5
gDX6kX/5V4QNSyo8bp3HGZowGKFdmeL6DvvL+qlGaS2wi4qyhEI52IrVFu+PbozILiAI9Y6SMnDY
EYbpR4Kzy4K81Ye97C3NSTdfACJK1FzJ94JAvbean58eQZqn422MqqyhF4izuekAJUfdicNOAS19
EuWGa0GHj6GlOzFYZiGd+uNjkXT0e8u/1+3yPY+m97V8my4VAgqe8t1mT2Fhr1H25Uy+S2jJCmQi
io6Yq2YoRGOdISg/gsRK+sbReBb3g3ititsr1h7U9wUNtMf3/lhSGR87z0fvLaZ4zw3vmiAmzQew
KgdP6DZpkjCXqCiI6mX4ZJnqhOrOGI+rJo0PcOKlPfoytyVREyQ7tQ3J9QZ2t3TCbOOMqO3k94AT
xJvUI20r51OnmtajUw1TMtQWmFwRZjepMEbvp0n9vRu9f544js6MG0PsZqudiLpG0CKd1AP9UmgD
qToTBuApaUB+GGmkD23JRCdfqMgQxX+OggJ8dUUypT4iqsbtGJkiz7Q5X86dTLWJCr5P+KfF4zQL
rNi2hTU8DSLfgP3JHeESWJqibFeVNYCULJr0p32LpSOYiiv3yi7GhCMhMtdilR0B48iSdpmtj2bK
9IqnKXsvDTJ/vgGakScpsoqXgvurqzyIQtoFyPRgQZlHVx/nft60Y9j1Yt5OGS86p2mx7JyHlPRc
86V0XgqG3nifSYqkHlcIPHin9hmSMJgNjuUjuwe7uVRzn1OZdduJaimbNIjMBypXjJaCpUMpz209
d3nuna0jKMxhDt9zZ9nJSRlTFzZbS4bnjw1EPlRPAN+oHbKkUJVwNxz9S8YusDkd+uxHhxdD093s
QXsUPefeLGQbv/kYhKMKCQ1KXx2QRfSKLHenqEFn7k9NtBuelDKkvUYLvPeqQSGpm+pjkaaXaJql
fFIPovirjv8Cas4yoCphp15TJrVlJcgspHuL1BmbO3/pWgz+smaA/BCo3p9nKytvbWwYsPHBcXi8
kKbn4siwMcCl59aU2mdMD1/BO1WhrCpIbY4fjCG/qRVtRWGHzKAPQDtEpK2YSiHiLPtFZIjZQJh0
ljw5IPshrKUNzE+hYOJvtcI9YFVuYzrpEPr8crhOcfwObQNRvk02NLP7EzWE7SsGgHt1s5CxioND
ZSag+UpU6ddju6oKcL0SLru5d/MEtmBWA9KfBOErRd1qhnv54LtSsKnWaSLI75AsO0ZADdiBbiml
BKXjqFjKGRdctj00Lo089dabdzocfO+lS2uwaUGuqDlSd4a7DVBJTTcizRnDXYaStgDiHK1EOew+
4MTyWxBlVH5NGIkmy40kmzcOjb3h28deHOJr4HwhbAfyDHGEEWRNJkP3b5yeki4bE/FZSac5XtGc
JK3zvDXLkZhSLenPKJqzwuFExZAgoy9cP9nqXBfiVEVja7kVh/t4bKnqFL7GtAD44PjofHyQ8gsb
ynNw9+7YzgmltVwJG27Jb0ZdI1000IgGbQpvBLlr/wX6Vb3rdSkJ9NAf/f3gW/A6FRaHq0nf1+jD
tPUjjjkOmFp42msz7CxyeJSYeGR/94agVkdGzJlHx0pVNVrl5sbivelgWOqBxT4oeeM+tXZV0VzI
cH1/Lq27qCLNqEtoo9nj3CmZW05Jviz9Z9XXQ4VK4yMtoeM9Ip/EO+SWhrv9OmNMVcbsOqzNSI0T
WuF4GzwBG0A7R+R7IT0q08yCCkcmnB3y3P1TdH4zfOc2woIdCK+l/LzhIxUOKV6ifg9h2RFFKzKt
4+AwjPkvR2WSY7sTu91qR4MgT8+AXyaclzUiWtu77uVNMcO79TA7InHgGR6FvNxmbX1IP1JOU9hD
PtkgvyAtY4n6dR9DusTAe2fVcq2Z6TCDiXJblTjS7LI9cWzwo+p0lZTKO0jJqvuPoSHRt4r+RiAy
m0yt12AUNjPwDRajGJL8z1/eD0TsYRhFJxd5CTyM/qfIF5A47gIWUt9ZpfW/xAO1xnVE2zL1++9W
mPCpweDQ32EzbAw5rEfv4+ZsiaB+58eBRWiNN0PRUYzrNohcMbv3d6CzfnTHjBVVQdU3OPkr4lXs
j5IOTOCIOwuRK1SrVsC9rwZt2B/J+4QBO2CEhljXi5sz9WeMQdaYQgKsuSW8l16oAIZwMkwjet1W
bVWkMYkY7JmFuh5Wras3LWs7Oyg+QNwQh6s8BnH7B0nEDdljrPWeg0ywzNdaBa5gXka4PV0Gs2z8
fOoN11JqG8AyIWU1aC5W/Xyr6lOUFVRp5NyvilC85JZSFoYN4gcPYPaL2A4jtUKTpe1slBxSIjvf
ulX2jC/VMabHcqVZr7ZHGvTHba4Jx+ln6XbUL+P7Y0DqG4uPgp0jP1xDwUFBEn53hJBucHzGNk0b
wSswY/BlEiMVDOvb15TfFQGiuRBAn34ulzKofdgCklPOx34tWAhv2hY0H2aI3nDKX/EjCrDjFv6w
AwBFamN+8ZBwFEUgo4M0i2RBMcU2WHL8jAYLZXrC4jooN/3gMNxBHrDHMjzUh3BuXjcmnhbPry9O
xFH4jMcYFmBwgvMnKhPpIkL9KfILpNgKcDzeYIqtQR8kpl+MrYXqWUsZqV0AEZpApzkp+r3nRd6c
b3De56zCXMoTk8Yhys7lso4GdP39I7aP5M5+XCfSC8od3xUIk9ld0UPjFJUrNTssaN06djdO9D7y
cAHpkCR2Ugj/69a+Ued0ksqOqsw9iKAq2hXVPkwPdtsc7cVamDcB6Zrq32IARNEU9h1R33lfhMpA
DYEALwVt8jG5piSJC7HATwmtRTGolTCazDKUaIwOWvXa9b7EB4JvOUDJrZaGV04ia7GDV5Z9O1eO
d6A2nuWvNyuLqLIY5d1DAuML43j0Y817Ufgma040YkyQRShDnhgNZ6RfBfU+UTJpthxwEcFOCCuy
Av/xxLi7m2Ow6abnbZBkAIlrx9V501DijUTXYRYPnLMsbYnvKCY558BnqZfvDYlWp46etvFm5Ehg
tRhGxdeTnTmnCqg3sQmemRIP7dHkTbitN4eJE/Jot2IP6DtFZvRoFNoCTwLr6sOznT645Dx5BeqV
qXGFYIAYtoHphbDdCURyD7p9K0ttMm10XINHm+LrA+h8PJ8Y8fHSVfeHWY09uB5bw83PUevmCLQ3
F7qc5P/uourdHHFS9n/0R0vX051YA9N6t4ZKYnRpiz0ivQORXizUyHvq8AFAW7DSmz3l4arr5XAr
NAWmovmUne8+y7h5x6Wrf/Ewa4vQdD6uN/ihsmN6EvI/+MsI+0fH5GUXIqoTo8CPvMMY9ljr4bM8
Dfu/YlyAVMBieSP14gMeWbtYWtbCtighxL6iWTcnzzrzW9ZQGLz422ZM6cQ5W6u30vmZe/y33RwT
e1VQaukZo/hNfSDexPYEg79j9NoNINwN0usp89toJR88s9PV8X8vWnJijzeHv5bl8eWIOJj8J8PW
fAlIMPq0wLmhN3MRpHFjkQtlLeGwsBF7qKSlJZT7SGpSR4N+zmDPJOdLLkzBUDxHQAUeb7l7SVqm
UPuS/j8QEVnCR3QqLnFHLVLtH1tWvQb0kRvGfUa6sVKK1fsT/ThtrqcR9PtAu3k5TejgXxwxxe3a
Mn9BEz9iN3EB8oSgQayaFh6WDN8RC/AFTSJMrJhUKf58EU27TiJN7CzfxvY851mrJWsXFaKoS5O9
McjQyxpz8YXN5yHb+xNsnbTuG45EKvsXDxAqzkCCyToY/72OpuveSTtrsjQEC7W2Mfd8NRyk/642
zSicZ3O5/PkQCLnywOUM/vZbwx4ChEusvFdrC1rkkq/n6BPeWLZFEXqzDSEbwBywt3ozo05v5yo0
wiE+QX+876JVAAowaRv6odV33Y9b2LF6V+dp5vakxEGoK/xUS6jliCII+D/yS93XrWDL8XsLcqna
YQhqCyio/6lqh5N7LV6P/oKvqCpa+LYw10nEPFIqA735uI0fSzV8HQzMW2Dd2KAunkYM7VG6Qf4f
OJ1+xYyA6fF5hU1BEM0eQ5Y0Wd9kB5HZhiF9tV7vYC0t4vp1DY55r1CkK92xxuGvwz0QypCRe6tC
UN1c9jLB+j32jCMGU8m+1qF7bZbZjVav9u4qwzBrcPLxZZXCNoIAlgXA29WWDJVIY9KqHo5d3/Ti
xOCOAzwctqtNWHdNLaXXrYLsI4ZMqYCpQUqzyEwGT1DtMOt/M1mRXWaXo9R5OkGgZoGYCKtqYSB+
byMzGhTkzZhbK/mfyD+gDIssIiKDdeSwLd6OnkyjfqzjCbQ8nopmxrozR803whpe/0mHyXfdoVt5
ZlyBNjznVQv9bWTJS9csYLJXeI9tUVYCTwptYTDy9umbQimOw/1q8cQd4GMGshhF1JoVCA9kbgJ9
8T2rMB75Q2wHzyBHccOzeLuwPbhhpmKqW0kcEJL1lFT3quwvhyNz/1Bhd6ABoVAH/4in9A1RNPa2
FROrb+GJ65lc95gyBAdU594PyrQsCNkPr+kZAO/WFGKaSdT1TLmABuILnHdCWuw+GRNXfK5kbq8Z
FqeamkT6QHRFC3m5bkTCXpVwpOV5V44S0E3qct5gnDwEK5bWTgzZCeq2aeJHXgtGLXLc4xtW0l7D
CMu1j/KXNnsvWtURj1SgWU9wabYJgXLTJHXJBZh00A5rEBxB802bI4Bs+xLZlk43uv2fqa6nI2Bm
pyBE/Jrnpwx9PvXgHJwg3gRRNoquF3Olu5YnwblBiiG676N6dNVSmxIy+IHxfFjN/M1uDfOdjvca
RXiLZwst7BU9YbZDWxDbjlbs9sTSSXQBF76J0e9Mdq4zlVc0c8KPMQmZ3Aa63IaDKJjCPMvktT8u
h35eR3YNg9K7R9NI3Yn4bAS9wXb7m0XUhgXFu6qD/bnEWh3zz+GJykIpZH/5zawdyyPLfEOT2gPE
w8VZtK5uBZF0yDo+k9UNruB1/3RngY/lQDWG8rtv52Qt5Eqp/DlmgAi+YBzeBexChKWrmwtZ6n7X
yGZqe/PvQKegaE7wbHtzZLf+BpI090hrmHoSxugDxiepwzXrxtKlBQT7Tk6VMG6Iu0XIrCDwOiqm
1H/xlkge0D7xH73ofIvipO6+cbsJY7ONgDCc/h9i7SYDqnm1WMuC/XQ4OPRDSMgT1+MVEBxnIYhO
wrE21jlGYihswApWTZARc8Mr6UrF6f841InYrhiOC3QZ94mi+YZuqO1tmQCZwqq9BKjepn6e3hR6
yOPufflufnsoErRQB8LqiMHeCaHIXpEsElYsjZFtLH3v0iUEs9eGNVuCmvg92/N2mUlzp87qf51r
+Vq/A8POw3UlGU1IdRDE5HTxH+of4gbfGtxMwLspFmOTlHvHaqPFDMptBjQdJQP+hr/5mqS1BAES
osBW62Uidn1mS0Ygam7HOIB92uaI/VilK7aTV5MBeopYsiqJPjK91OFghsfa0hgpoDa/SWkOx/vZ
whYmze8vM3mkLUoAo4SIAADjrIo1gSyEAcFD6yugJXFt5ooY9egMczfa7NJsPPqTzgfRXCC2UCPi
7Dfejf8qdR5JQCG3SOnzQijSER5XMoqFLBeVd485+AneRExhzBLryOxEuxukLZyARKDhk0daYYzn
3UvDlRwc/xdRer+LaxpH3VpJ0SGMuII2k9DmNpZox6lmfWe0lVp7/Rd1urph2xRpiiAsl3LufISa
E7VuO9zWp2RBwnrxvDnP6Evke/wgka9YX4zs51hr9bCPanT+SYvz4UDS240GSgUANLlVrZcp6J+u
fPsxWG+aao1FWFGPGKvILBKopZ0mvSTytrHJ/qRHRxCkXaHOBW4OCfqVXXlxmu+szrt41b6e2XHh
B31fg8vi50M/5M+J+msIixz/ZL+QcpJGXOBkwzN0gibsR6TJcXqQiCBTVDXBGCu3i/dIqhuxR0dY
MFxythoujV7jN8oWptOQMbnhLr1GK/ea0pc3KFt0qOvfuX3MvOoc9xllHmNzRM7y8mAwWsw1D7+F
WkSYi5LseVCTwXuL0dULAtfTw77NIeuWjQVi3HmGqnMt2ck97kfTLhtURFtUVOgu+zUKNLj1i4rM
Rdg5cIKfIcF3sB6dSz9Ess2cshIlXs1kMGCtiXlKWQrQbrKS9vmxXJ/WddO/Dt/bhvBJxQaIUYFU
jaWE50mTVs3Ng5vTUF1nSw3+iKerk+HqpXsWsgL/S/nz9Ln3a18l47I+EzpkEX8Ax6HBskP3xYgj
JaD+p2VDjocl3FKFpaoIH72qldQopsAJPRHzrHz6ZvLfgLc/Y86Bo6K7i03O++7HHhu57j0GLaeB
5hUS97SHp1mBkSBNddcrDvAyogw+wKkLvuoJHqOYGmE0K+T3GTej6p6PGVQLBBKKQR/CtCDuVFv8
J6IHlYCaAv/yeYjRXCD0COmPgT5FSrgMjtMFVc5uv40DuKCWZI8saJa1soLw3EcSoJEPEOj2/U0K
AsKqrs3MXO8bvxGB1yi0mx1lDHqqnROuFy5KKGkUeYUon+A7v/Y4QxKHEejcoczNNNR8wC63/IAq
KccEFHzp0CG5Jat3N9b334038iFg4BTtWR52J4LEU4/VJWpL79rdZi5IVeMTJQqLpOSX4+n1VAr7
qG70OpQFUruFo8m0zo4nHcILhaWh4nLgq7ftxFblpYS9TgjpAbn+z/LX6FBGipcLnyTDz/RXt1/P
RzNS1cdNkgq4agG3UwwN8kbuZSVFf4PAQ6n0g4/lKIf6Sl5xpIvHjGiMkiKCIN7kCH6aS/qUX15j
U+RZgbkaN2/g174CxMfGEmlna53U9vMWc0KYlFWr23rhoxTzvWeZ3Pm2IgmDM9umpaLgGOXR1w4Q
MC2RMdPcZZe9/Lt+kBH6lTxGvKp/2e83Z3aWW4DVovAKua67Blk83DeTsOLYVHXUMpAbvbpNNOfH
eZM687dQZBHOePTQ8Uo0uSztuxL8N3MJYMzp+J05UVY/FTDjBFcJNf32OqyMRfQHifB+Jzfmaer1
IdxdyA+R1Bs4W4LdHBp5H57IO/OxLQXQaBfvZ/odn5LA20A7S342kidAYxnQLh/mbcJsvTdF8WqR
VVZpk8Q99VIcoCgnWQkzNNtsJRS1866VTQqLEHyMO8NAqufdrbn2ngKRMJMgYW+YRpLuF0N6RLb0
zdzIXAGZPXs/Z3ADydJCdM+8jaOpxFol3J1a9VEaO1wXGuxeHbZPoJ9CK4fBJLY9bihQPxQ989dX
icjFrOI8q0oAd+BfUUpNCQ5Ydm7r8fC23zoNXkSZ5RH3zUri/fD4eoWPY2cEKTJLIyGpmTY1vKE4
08ytLzFdIvMqp2+Jb42O+p0cK07U8OGCGl+x51+VUTFEWdHj2/XfzosTDmH2wDYHNmY3mtfGSwC8
oUcajMtDrFHXvAfx01xuEr3HRNyGUmVyhhxyo7u5buScN4fT0lPeOMVHyelSAjmjFITDXnuGkbrN
SHRDEAnkBlN4zo2kiV7VKrQiYCAUAWF+wqEt2eOaIrdIAEHRjJMtoYUd1mCyncg1sFsR+J7Bwc6O
uaEZvphG6AC068yBJzAZqZIqejGHGdmryKlGkoVE3nABGVCnEqLf2hfzvZjJG0YctVuf4IORATmZ
XvBv5OwXz9bo8Ym1ezjNzNa/HLzDo0eFzScU9g/NhhcJ6KpAW75nVllB+KFulxxeZJKID6qb2y70
k9gxiMPX5Fs2HjjxcvEfmOYdr+hwyw5Y/gfQ3nTR2Al1LVuJ3VSVzJqYWMM6fXA+eP3V5ODWRQYM
7EfMcG59BKSGk2RDbOVmfp/oUrHfOQBphzaO2jcAUN/sJednAzw0IQIQhVDnZfLKulhXPOpdrYvd
a9T/RVSU0qf76abHMyf0CA0NgDBByZYjI2qGQ2z9y1k88b292tMc8U7TvX+O97jg5l73PHIOHxMg
OaN5C7rb6ACFWFutzvSCOsSugpD86bugsBAtMFRZy5DUcrNW5CwpstG1cX/BpBU+Yg0BeSmq/AO9
rzhs++ylhlbbnNJr5KBQTbp0ohd8KxSDDRKIcN0/6FAznAWrFRlgkDlPi4P8aBCmKuRmCGyyzDiq
NO23Rg3VblKEod3EsjHHfixu0osCfK9gyHZGEeuKsBvWAdjlwPPM1WFAXLUE35QbyflJqi2vAxDq
epwGxdVMs5UtWJ09qdPWyOx4syqvlB995fPmzQUccxpAvKIM1UD6ZJ+eIYqtCGFnUhngswo1fAya
KJIo252EhujXTdV0+lSit+aU9IxXCl8ENvR5wSo/9vNotegS9Ui5EajCelw0sSHsPJdwklCDfDp4
lPV2Nitqa0MVATlcXh+Kyyr3NnmKDo+QUMbh1/f6a8iU7HmEuk6cw4ll24ed8xx1ev5o1vKrOQ+q
d4xKPdxTKFiDGtlqAx7gk15bvbyKnh+3NfND8cTgPjW+8vl9z0igMYqyUMg708nXaSBbJdo+wdia
Jl2BmWZ3HtIfi/TdywyTxAkdWeVeuM5rd0v5HWh0mVoLu8cZS3UyIjuvjPs9hP1INP44mLFJCQfz
sbf0C6K8WYDMaBWvolGMt29L3mwMwF4g0LisfYehBdshsNgynWxKnPwxNgcjQppJLbotm4sS5xuj
qi8iaxejhNHXEO3nS3VHA5FhcPZ+KC/fatAhoB/qQbVkUq0O2xUi6GpFBU1+BIay+oR0stjS+hD4
2TSifEtRADq5lieKkCFe9LsqwRYKnwhHi8bPlUtmojqGyg8W4CjszCTsXWbG4mmFsPSRlIseImww
dgclddaGIKwEZzjDzYgcW0vX1Ofn2U+yf0ydb9KOuIog5fYKBS+1LyDzbHO8p6VvIIiZ5enVYNEH
6ehlzStiM0zYTB5SrFr45fQXqPXp1J0XUn6TEAnTrZ56Q7HeToIh2yLibWLCbLSjSGjTkk/aWjja
TuFV/PpGUUduWi+Z2/SPfLaRGGY4abqOdI+DM0GWUQSLr5zwu0ZhBioZcsOSHI8eARpSj15P+95e
Lvqu8KpQ0P0iptgExMRMggLt75Se7bshaUaXgWVpwrrWfir0aDFqbvoI6FdnUtffRwpExJOBAutc
WROim+0hOOMHiiFzkpJJeJgh8vUWeNKj/z1HEHY3QdrTg2NOrgrBW6uuIaPSjLdylIjYas0s5P+U
HK4076k66GUlt6HyaK4uJ5JiThPgEXTGuyVaYVYvpkOfOi7+DuHjRlmb425JDIyWJxpxkrIBD52q
XYfs+Zuc4f15kN7D7N53S2ozDjzxtdsOExYv9Ef6VuSTFzD8eGF4hrtcoW0pqHn+i7QZR2sxILo7
Te7W9lHBKIF4TcTPv59lXISsE9UYRt5jZ3x2jX8Qtw/Rgtjs/ZTUFAc6CxjMyrQS9a5mEXJnY1jt
0ZbVSRupIMZ5DYQrrkVoezaJvYB7mp+TtmgQ+vAYgGTQGiCc5CyjdQgv9blPtfSFc6D1h94c9/sd
0N0MGF1RAvq2BKTjW2OTpbEMhHbPo1Wa27PhiXTBhlxj2o8n365z9AZ3ZRP7rOFhxRqHz3BWGOrF
7KFKb1GK2Pzog97m+7Y6tsD8HpRFefxspzfBaATtDp32OLKSfBK0I/lx/Df8/gWQyFYH0WIC3cpu
ZYqxKFL8pWY9dUZtMxBCECZjaSsuuJ0CU9a6vQ7bOVad1pyTikRsNfz/8X8MeeAeKBoVpdrhym4H
53/q1g/1KA5Kfo8nQcjWKTQaIjvJtnQIHc5Z0Tfv3qFALBT0LYnlssN3rKNUnmN+65fkpZDCqHft
TgUUDEK61ZFhkebJnrd4sirvMF7DAgyDneAMsXVSHnwqfsxqmvFPwK8eN6/jfjplb60TF9BnOBzP
LhXm7Q/drDnU5PrJVDe843phNG3W8YzHWak23HyvXZhsnKWb5bPfVwhlXKy34bIXV04/oJda8jad
zmFUUrUGsbCVKDSCyhWMS+GQGdk3dTYewz8P+REOLbRMsJOxGuaKGf8svzgL2PFNcxz0eDmSSg9l
H4U/rklTr5+yjtk3rNoajFGNwMf2SX/c2gl005DYnD7kRDeKmQ8rv7FjDgv7qmReZjKw9IQrTs+3
k9VKZIg22Q6nX4Qy0W+eXGVaGz+3e4bYbwILiOVUBHpj2Dx+DdlvVZInfPNyIv8W5aNv6j+tKnVS
uHaYgtZr+dAzjcChnvYTzfQ5z8855pkN9o0ar3cWStiPeV+FG713Ln4945fExdwRkZub48UKlUDD
xerbwJD54EBh1DFXoWCGKXTuFT5CX2shVRLMmSZ69oUIgTyO23P9Vx4zXMGoLzmTQDyg09V6SvDJ
ZZ4R9iFMLxQtBt8/EDjghzLObaUXk+7TI2yNgE7IYB3aAkBZG2F1lRtPHTYPKg0rY0iA8790sphT
4NsmV3i5wciXW/H+0pdbVQcCgbrjj2/GNJgKf09TA3GTPtqBw2mddmdF/1qBGC0XQasiDU0dLdiO
jzma51InNA8Md2erTlJVfun/F+ZBfU09Po9H9XggDxKDk/hTlZNI/ZQoMXetD0fkL6PVOWhLdNCH
HXrsA+/4BBXDN2SmeVym9aT3jEgHBIRn7XCDTlP80hZwhCp5nHcuckJ0bTGGRA2WFxu/NHjNNF9v
0DrQoII3OUs3sc+s5Eb5RGU5pszRATcOAzPuUQ9eJk/noQBIKXKY6yn8UGMzGUWUrI9Sm73ajsQs
Fui9YKUV6x1mH79MNGxNNK+eStOuW5dTpJwLAvfZhXwNyj4sgfxPvWDnPuC2zvyzcAfFnS/GrG9/
eTTDn7y1uSCL9HmTU4J+upwL4XPnGkc5O1Psp0Rq5dy1tARaAT5+kFK1sXQjBL8T8L1MV70iFxwS
i5jx7Tx8VvRIVeUfDnEqMwQeCgsUdydpz8vQCMW1WV9XVfDxdaMCPsNCFfn0nKsU7Tah+xfnXjkL
RClXGUaJQuNq46rdtkb2AksVl4mtOHBY11g0Os9fAmEq/55FuThsfgYuo5lFoURqG/bE+k/wDzfN
kKzI/hX+NtsFTSRDs7Leihc1JNyHCetVBD9EZ3hnMI3nXJiJBRDhFmGJdOOtU5EuON0io4/1awbn
UWgzDtp0J9u1FJx720RYGI4M/cSGQB1YzgVoDMF70FN5uTl8sQmHqeZDgvY9+Zkr+m9+1OcFHTM4
u5NlJXTIiyBlVSzTFoWSVFuc9yDMNCoMYYAgRm0veiJLiCBarBSVztBrAmhlPtgFAE8GiHEAShxD
JgD5SJiY1aGcCK09/WkeT7+lZr8JMo52J+KsTJRg+YSpY/7pCc1TPweES3K3cPieVxd5xfdUTVbn
qmrlcy4+DgEPIRaOcBkPsYBnBvE/4PUTlFihKELmk4NKyxpnw6ZzzvWTko6805N3lbrkFUS12/Jz
5apXd6LCgrwSmIz58rbr88S46yFQMhpcy6mC9f72kvNbjuJUtG68S12AViHjKBJhv0wWTrs+8Ydd
qwRHMiSoNGnP3vvfvyGZXfFdYk/efRyE0KLgF4w9Rn1PNRm8DZE2U+KSgyV8+vyfmmPQEh9f3MaL
W3N7sM5IQnxjZddhfNYQoa1EtyvfWbD1xrMuV6YjR18VyKN9dGP1kCjuRD/PTTS84gSO2MSl4nbk
6iSsj8d6nJbfy9hCGz0+TtQ/BhEb6nsKAddObLaXTZHE+VQsI4V5c4y3S3e1Q0hGghzT9f+uMC4h
C3XMqYVb1m0YfvfnVMuBEGI0k62xTjwG7LKxpUNf3vSku0j9PkW8DiQ78YWM5If8wbXBne/Wvoo4
ZJqWbyOZeVhohTtMEfDt6yfCCCrmqt8zBPgXtz3DxJcyjOGBlbGDS/owBpzh9vet67JV7GVMpMip
S9JJztFrK5aUQW04sDvXKp60X038s/E59c1JKNfOeBcfFQ92mSDVTU6T+n1VdF/TEqsMswYeeHpj
WbMiK/gy7sWXli1peKhVUEwDqTlDVL8wA4XLf7Aw8mXs/K94SeiF/mhi2wBYCMZfyzV3nZUuhc69
PmbI88hU/Lo0SojUlm+Zo8B0RaCq22Y6mwhTK0NQENbJHkl99NzLgueV/6G2PwtWyJZjr8ULnBbx
shUv6b9pgZqKNsJ0/rMpJZsvipxJiwhfb3i7lvUrGR6agPbuG36pG4g7HECiBfzLZZzEBGgVN8Cc
aDrVLbNjmfAzUkzH9zOb74/ISr0kPc4vMBCCEE6DsRzPre9ZuQwwAwYiD3Rsyj6gFiQUmxbV+WGQ
c+8KAuS6VK9fi2rZj7/2EMY8tG/d1xahFisJ04kQxwx3zeMgLewNlsfVNEbLHI47iRaKa4XigHhY
/03+TXnxoBrmo2rfUVd1/3nzbo3gPGwVu1q+j/NB1moAlYqgNm0Fj0fQAmJFGccVnkdF/PwBYYHO
9bDlWcscSSqg9xDqQ8CglYh8FXBBf9kNPTHpKXDNm9wnEDG0Cl+Y41ZpIG1dZ5RKLN3quW1LBL9T
Y6wiu5fKfnyX9j4BTe0h3WFBuIEzLL5QycGP67QzimEa/nFbzkc2Kz3bD5KbfchfcN44hJv88sXy
aEURZL1E9PHU89F8YGQdoKy09t4L/Wh0G69bn06/PuI5D1etvKzyeQFvoqtXaeH0GqU2AGXOoUyd
kKnuZjbMy2NhmZ5QjEnDvT0DdcuKT+4cVqXVIo8QGUx8C5q6ETSBGCk/CA8QeZXaUcG8kqkqpV6c
CSTrF32I4ZBP2QywTNSyOmLjDc7eD2Dm3DNjLlzB9Nl/3aj+3n3KzPTF6Xb1Vutg+UDvn/0eqsvy
uZXIxBiHZsEFjQ329TZGDwPJ7aZ8qAxSltN7yOxPOE2DEwLcZpvOQFcrzv125yLGzG81Z6EnEtN2
tPldfJdnPEYZCJsOqS2f45/OdAZ9da0hRfPAZN1eeCbQaKfjiqXwRDqrcedW6dbaPYMAGkvcfu2X
FacRjIb80VF8wvoqtr/vzIe3raCFdqXaz3an04xv1LhvpgiBbjQbeY8eSJlgGRltx3y9+XGAETdH
u9/CHx8fRrDqKRWGDJMnw85oRIRVEE3A1JyJiy2k2vyV7NjMDQErkNYzFTIztkoXtCoUx/UbCpw3
+4ti0dDG4+0DjkLu6XgEHGh0r6zmzs3KxB8VlNMv0lnFD/lGESUP+ZTZMPe3k2F+WRvnK41MAFjI
FY1vdLUY4FkmULHbmp2SnIEWDx7O81AQdDzyEtrFeVp9Vvho3W3LAuNh5YqI0Y7Ig9RzT3FJCEfk
mWKViqLsjyycIFk5BMbKeZO7JiFPNWLh4xKVKjICYAw20O38F4zuUlooNaP1nbgbYOuLcc9INFCu
Kh9ilXuH9VpnkxLcQ9/hNLq7p1dMi3jazFJwNYXGtZepMKVxOnS2BbB596OatvVsNOHeZOLl456E
WxzLw1h4nw2mD98DM2MpTEjxlc8vEvhY7MUjp9huWMKG3OmcdWYbhF+lVFR1V2ELm77i0mc4Sw7i
Fd3KJS1ZNQyglVzOFT9pFM4ugVEDz2yW3IWY3M2Kj5i22lnU8WDfi1yI6tHWPHJjkWAq2OsSQ47j
UW518gMOnhuMCNPVGx4Tf0jnTLn5GhacZ8Fqk2/neIhJ7jYQ+JSypquLebDWdhUqXPpUh0ooDM9i
67K2/ndzKvW0zZI7h7v099W7f3iumVjPvKk/ctwqwKHtYu4YtCC9igU4prGwBETdyrLV+OAEhOdX
qgAS2GGcVPjmkRk0rN2iJmHg/H/BDYGvtBgbYgSmxAvHTTjebGjd1FaQMFIi/et9scHw5NV4vmXm
cpcmT9Sj5yQDi2mvUt0t8XryhAfeGBk7pfpK6qf+/2q0NMbMbyxh1XjZamPutgIMJJoEGlv7109j
bGABO4j0Fe9qjQDtYXLehhoRZpN0sXlEiHCFSjlMp6zwPEOKjrqi8xmuXEQhJIGRScWYURHuzbmp
dXCQzzGpQKQKsxvhm07mv/V0NOWu/3zfk+7retXzXSutCO++IjqNzzF02LCtnWZP0zrmmuOvodE2
//jvoHcrV2sy+5TEQKTV3OKfv0/GVv7F1InjMnr0rhJy1iLKcOs9rXGzDAuZh0i5XkeKFWWCfolQ
P4wfzZpOVsa1WeX0bfSICqzDtzmZhTa97JUaMR8V858zVs0U2r3+XS1ReOwW0bMeRcqoBZMIuLeF
/hh2+flAAIo0eNKiO3Ivd1l9Sztz1rYzGZiBu/4cjEOdXVAsjiUkKh9hAYcxf2GGklgoLUI7ABDh
b3I/BCbeZ+WuI7YELl+b7Agr7TOl2pdJcHrrlw8Ugrsb/+vDQC7/9/ZSO+WkM+MX6g2CoPrVBSt3
837ID2mAn8g8OHIcloYradkpChNkMUeUyZlf03QGyrZK2zocQPWhc9CZ0rOUVKOgGqBluz8KLsXu
huoyfIXgWuyK8vJkLdKlz7vIRnP1/GnVSiD7nygsHRpMW+HyZpvxJ+9wl+T0edeeqI7/pHM20A+e
Q6I7I3NKNGdSJJ1x2FSkhQw//UfrlAGZjGWucaiRqZViBjBZgDfi+MZKDG91c2ZYSKEm1fSgnRQn
0IjMl1kBqH90dk1uKlwlajx5Yq0ypkO16mmoH2pCt6bFmRCRpEKm7MFWdN32aMTP2n6yOmjGiFfc
pI3OoDMqU3Razlj/F0Bsw59NAr6TTFP5FauxfgGW661rzfF41QpHI/LbASuUT9s99Na04fy/3euy
ipg+kZogOw==
`protect end_protected
