--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
oR18mZAiBsbEzoQ0y6QbkVJqqqCWUIPUSwYqf3T1goPwiflNjN2V/iSToz2DorEm3AH8drcUQBub
9BM9rpF1YwxtLm6lkjIuGAdmHr4lOqbfKrZSBOPci6ME2OVHAdOnlPmBbO8h7UFEmWSZghe+LKaQ
QwF/UIkmvFY9YQWH8LfjCpziI0omtHOZwRXaRDlMm8bl1OTEC6Cs14iikv7cmKPsQcFZI/bFazNv
uHxMkeqmQrsG3/G32L7cVOugkk9TVKxvWh3PLEcKjz2vfZmfm9rpxD89ptvSE/GxCLpYJIzumiXH
wFoTLCzg8LAAS1XF/vYY0ijZaA4Jzg594PZ8cQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="w0TgLZdjltXQozEGi5cjPia0oa121AIhlyX5vRWeNZQ="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
hegMEhY/SGnh1FvvlXpFGLQYV2jfvVPcivWtv5YcB8cgBsPknNvRDWAkHT+ergTWwfpnPy/mwGN6
XIJ7F5oGYn7kRgkJ7qICJIJd9onASslhBTx5GgfS4bmDAomJHLxiRVuhKQeOwrsqkG5UdswxuYw/
sOzXLBzqcbWQmrK3WKgRgQ5pl8ug/NbdHC8w5WCFhrwqCuCWCLbjWDcgsC7qNe6cMtG7y1bPQFi5
Y2c5bdOJsNDBpbjr8FEfp8py49YbXlVK5bWqcJCe+vdXECRUUjBTgjdxaqDC7tV/rm/cPmbjYm3J
nn1zBGpRDP7lUDzd589tlGiUeDRnlmI6LQKY6A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="E72V1OCIkhowZOP6KXqlFwJj/U/aDIbu0zbUkz7O0Z8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4016)
`protect data_block
yl9mv6DF4AJXgsdmNe4hzlfDQFnbjuVvHo6jPeyZWHFbLaNTTsjN2Xg1th8Tf8Q+/RlH6U8qGAF1
uwomc9gVWJucDxEFTXrPW74OGQobRk2j5MpSn3Bsw0m6upNI2A4ShclSclfged/uqk/CCT9L1m3y
HDFXbzuBcv9ncppDyUkVlg7FqwOoMjlcMG89smRhQuhplOzMu6mQSTRzD4ywzyZoNnsMRwTnwbGg
PZRJ/3kxUv8QEwAS5XQyoUwe5DINkrWSNf0pBVVt+/3PQwvXJ4wKeA/6dAuSAdTv+wvDHur8SXKI
baRxdLJqSxfa88PdpF2FloY19UBSOt2EPA0c6osXqU0P3nL/I4Domvrkl2mFdSB76uquAngQLH/h
FWjWISdqj498vaEWGtkFCQd2+3IOrLsPe8VUvg8BLjQ8tiFeXbgOqWoIv2yLyT55ykwI+CV+ze7I
8jQ1jXfm/tpJidz+0dTjaoH7lekI8S93hLfkRoPE91HtTxpNZgNbDHDAzZLu5mbeCBUkbF3OuHCL
mo+Hm2dEVgCMj3mGUwl/LUIknJndayfVdf45+uvC6hsgdHaMJjY92pxD+NQ5xcmQ7E2eulwduhMb
fQNV3MhDiEBPo27xIYBAquHyNQzefQ4KMllfIqGiUipTceXss0zGCYlADdNlzo6RzjdnFK4KRePE
q6aYo9Jeuh8CtGJ0GjjngPA1KwiqMk77bUYQGiiLpKZOgfeOJnnLKE5dtAYrzzOdCh17a9LrOl49
ut2H41AzAFXTVZLYc+ttbyu5vFvoJHaO7FANo8DDuJE+P6h8aEOHubOEG9j4nkKUFhi38tYrXXTP
1sjndgwKLynw/4NwsT3ezLCw3TiHPDGImvn2TC4t4cG2/SHEDPp/4ZFlvtFzyO5p3HTJ91TXhn8W
+hTUfCPZNiaXkVCsblEW3CsdvF8naRicBH8kbfd6UNYgrWrpsEKzL1txvXDMcPfGFosAnEeF5SKT
8a3fB4GDG0Sm2YHtrcYNpjhaQ+V/hQMNudOROq2x0YqQWnuX6qwRJPaFsfNkkUIliVeNLSwXqOhG
4DG7Htk/la/ymUcM+v6lN7gowmVkcD3DE7PLGGY6Ny9Yu4ZVoGtJVDkdq3w0iQgBn/yUKU5JNg5C
WUm63QOthkukQ+NWvKvzggNZuJaebZQUwE647BuL6fHKb31m2Vg5KEufocwicBMUNioVUSO67dOu
5BqwdmdAjLekziwhSP77G/b8OuwEsQRvTrJnYD5eqvWzgw41TDu0SdtIj1G8DR36A/CV36tNnbiD
9d9czoGf7Cu5Ppdon66py398R5uQK1Tb9cglgsG9zdW77XfjPT2NHXjCsH1qPYfO2F7O+Bl+E8vR
HE3tOvSZkhdc5TmICsK6R5rPoVNjMQicDVBT5ZP3pDk/XBdbivB+cIi3+4fRzAf99BBVddV0V09u
kNN6KyEJ91Sk4bKDJEje0KgkZ+jWhF8fpphd+I94oxycJBOcNyDoZVtUShao/5+N/P4k1AfqJl6j
gSINjVClCPm9XtPGorbh+eHsxwqLbq2srwqHO291R3K6am6Ss1FfC5BQqzPQ/cCMfjKHJ+EbCOxU
tczhj7hlTCWU9n1tjpuGtCL4caVzRJUUnwDMo7fPjYFyWuNbVG18Yrk2YL4aEWKl3tAjUWwAFaQs
q2QDbYAJIev9PTjSkj/+bn5UzoPs9geyuTsKFxDUbOSqILn7XZ6/BO99elXWK+C1KX09i9Iu71ZX
lUQjGL573yC+Q75i+Y4Oc+gECAmqtJwWfKDJvUu4qxRY7cNPCHlIIwqVPBjYn1BYI3XGHCTWXkGQ
6cpr3nwZk2CNOOmnR+hrCr2xNlr+jVhs5apWUvC/UNaEJp6bhC9aDtVLGEPDd4HaMtYbiPsB6bmw
GiND8NIA0afG41ZAy3YsJjEvAe4RERwwys/HClU7SFMRu6UkHe+cEchq+j0UHfMknGDEtEGqMILA
cwcdt14dzc8GFNjUyxnRBIwdv8NR6sdnalrr6WG1sJZCejV5V2GneT94GRjFUYdztJpmvi+eAYnN
7MEMGkNmwsqH22Qhb3KBtWGqurPZzC4471QhrGnBOFR+rjKw2s88uWpBYdLsLct2K5venc90+Eta
bXYGtnZFIKnObdl5oMR/LrLF7zmr1oFnylaV2yCjA/M85I/dv/0oIcPYqXlNQEDAum8XuT3TbEsv
Np4bRK2D4qRilPRU/rQZsseFnuFmGuXezsZ8632laXTCedQNDoYq91cSZCRd50mTgaiRjCt4rg17
8ap7uiUtDO9A24LunlLyNxy5oGIqNyxMwCZxiZqUWtzguPy2wEdK6F8n8ppCQlCf49euBUCNcWgl
jAwVKUF7RDl/kcfw2vOIrbQue6mqLD1nD/oF3+JubajVXpyqMFN3g2BEcGmLjop+Ld1NdRaz54/4
bu3QgL+/SbA03/FZBZGvpLvSe9hZ38riBhPwZMpec+hDQZWq1VVdZk2kqrY/7a4yQrcoSresZg4l
UO73pL2LUz9z1Pn0+IwNd22Y9p/gFjUYQ3xegfJ3FBAXoreTwnGqR6rcQrrAQ1bxqD2bz+u/nkNT
oej4Vx3QbEMhFDFHFjfzJntBaPhuR4/lvVkuQSK0S6KT/qGeCM6vv7HZra4OVRt3mVngskYxHM3k
czfsMmJwn0nDP8wlOcdFPN3iuPwPFRxuB9wGWTYgpzH4NTTUHIsxJ4FCAlB1ZJAsLhk5K/wAMGh3
wLmxJWIEBexqPiwElsMsDJcqQ3fE9rgQ12SUsCUYdCe9bQThb+PT2B/YRf/CdmpUABRflxfjRzc1
LbZ3Pe/7HD7A5uMLd9FG3YBfo2HQ37GOJfVi7X7EH6KrjwjBHSIajZmr+9Sd3SfBSV1Deux7w4rF
GmlCo7dPv4iMZ4VSexqN0eKlZN3d/ux1JPeEISfCW+YU2fdAO/b/2L+0Tn3dLiQw3bgaUIOokqV+
NoAP2xQQgQbW06PCIhwL6n9xX4OfB5pAT1HYvrz0CzX8E4NW9Aor4rkre9MYDTpkzLazYPCVBsxN
quckKWZHCxfCbdmWWDLSKFpl99qgyPn4eedn0HaJryynfNQS7Aua6a6OM2QpacBwefTvSWKAmvMf
bGNqtRnOcS1hy30uAAW+SEb075gvp6QUDsiJrwhZPgpbUjbpoxPB/DnnSFdg7+GWDLAjThoTW7BZ
Wm0UuyIRaiHMaZk8tM6molP0wmFJnFnOY2I1mZfoTQykzEM6QdE6vZkjT7bGnANzBMIG2OuDyVek
CrE8XoYgdNThGcEmilAIY8LLLJAYfk90e0Oo06b1QIr8EpejeBfLsF86LBfAQ0B/jqfY5G8NH3CR
RFsPEvlqKEzEpGXKckviFJkQNL9BAToLwxsgrrKStwyJZDETcIAqHGgUacLnNQ+QpA79PgPX72AF
qQKc069y76nwMv1jeAdaFkja89PTuMJdRHEpEWVJGXHBD32b7FpAjghoVpwN+1sVPtnuvZkxtWg2
J2MMA73lki1NAAaxHKua5Db2WjXtvMMCk1D7gdiCReIIx/6gG5H7MyS3zAcE/XK/xHd27+gT2akc
hX4YyNnIGEebZdfq1nDgXoLvCusggUkJPwUKkolhk6QkPh2okp4xJdTPakZirio8+gbJ6MFkIt5M
TJgu0cI4tHNxCP7xcwjFuXkU4Wp03OwqGh8j4f7PDj9cB1o6kYhaigm8xdBHepKQ0PYLGVs1j9JZ
Hwkru1bF8aa1eXPkuuXVPL0H9XTPR4WGlRjoWaPlLbzxbKVqI61NJMWmJGf/2SQpxGYrW93nKMmu
+8cJ49cfiItEP6YxtxY5dTUH4hmneV4SKj7jPqnFV/QSRm3AgzZ0GZQDyc2KhdfK2uZMEVh4tSB7
dx2iGyUuKdplqrStWHtWWTsSRwK53Psw8pw+QLFHnVK5cNw4oH8z4heY7u8SpD9QUcdOjQ5W7i+a
IeYUz1pbNHsk8ugYNg8RHXlC+jq7hge2plXqYFWSE6/wMS9sP6lVSYNcBT4M8D55q1vT7mkb5HsP
e/fNCymDClhOvUDDd/wwT0gwfVdacCaNROk1MEr7NHEhQ746AlcVtYCH06Typv2GfHiOHxi55t0+
uDWeKtObfDIDZfoIhybmcCHmJdTaK2+gt+EmgbCLwEulvPLRpnoo+umlejT+llfXjjENA2bryR86
2HyM5LGBoI76oxm9mLenOu727f17w2bL11FpaFZcVUI9ffQUbi/ZkxqWv2uv43UE2rryG0S0BVlu
fxUwx9WWEG90X+cBHy9jTC1J9ewjAyjuiiIi05wCl8EW7WZwiSbmucXCkQeg5shpVOOeLr6klmBw
szD/8Fb3sB5vMvECZYM2X5NnbGXbnVER88r2x0uFdOJw/tw+KGn5zb8jQgs+KWokq/dWssrBLL3k
TWcsHRbH1c37HgAgVZrZVvzDCgrxmmPrwILP+2A6hP/a1X7u6Cx90o5xmawkgKIyadCtTEyk9Izn
j1tg37iv4//dqZwCH2BKl+E97pwlkdcIgUawozKIV/GPSzm3Nmspjwi2CiV1tELHVIghmHu2ybvX
jNSnKHO7msFmM9hCjN6jTIhSu5BacaN8Yw2QaL+0Z8i0Hw1bIzrWxBN2MGdwWarw+gVL8gLgma+5
r68Q1IZ133FgcvC09Io0gaPMJIx2yxGvbFSi0YMz16PgCixyHFUREqgfiO4mCvAq5XSRBf/sujgi
9BSO4PIAeYGejw7b71vXFXZneBOuMFZoyhk9VWMs0SGnB9P+DfMOGIekS0jC5TGNgwYrNxHi8Hne
56zHuM+gOpEVj3xGFQcfql8O5SLnultDRGD8spyX9CxPvuEBaA2F7rU3rNki0h17vwSP1GbAY7Op
coofoMYA4d+iS65D+gQ6QEJKomjDtsZ4YV5Tmj3628oemaxjHMUjvRyb8PCvUkhxb4sDIa2BgSAZ
r3yNyG8Y3O0jyKM4DMplIPKJOl8T92iyJ5PVs2t+A2c6/c8tIcGUSLuTab4mUBTiTdOQaENSQJ2W
sUaaoClE9Ry35jwvyu9Yrm8nVK6j9agyD3CdfNwlxjMgGHikm2/W/xia/+hTsCSCYnRCAnTidjGn
nOIY1sjJTzpsb/LaNpJUTquPXrtq6Wq1hrsql+8UrwsLwRcs+QZZ+wid9bhBmEGZ6Wi8JliRWkRh
XzHFPLyu+1SDNwnDXOw2eHkRk8yebkockk9nUgBfQymH+6D9FflvxKo+cFoQ9lreHouQ5M0AUMfl
k/GR+XdHUPLuI1xr7kGGpK/z4+vnPu7TVGyjZ1bWZUWz5V3N74o8R/Z87B6LtHYP9aCpqCe65Pke
fkNuExwqFc31tmrArhAiz4SIA55nP1mcF68=
`protect end_protected
