--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
NH3aR6/SyTsEP4VawYxfbDGo1x5cW6/vW0DGs6kBcEqLToKJBhgS22lmFDIf3Kz9juj2ZOYyP/Nd
1u9XV+DyeXMRvTb+FFC3HgYil1AmOpjvTeePev3WYIEgOFQU09RUQVa+tyfCp7r4+2V/nzcO///5
hEF1YLx82Fxq2faZurFuwUNePns+3CrvnHFTBF9ztJ3/KhNWGPND52K7F1s4/lHmER7SuFdjBJuH
9W2Nkdz/SHqIhffj/DqeH6DyRBzPXvJLfgk5s2MMntPhSCLs50FVtsoQP46YddvpQm41BHUicoMW
xQjUMbr9rqLcYALbCdZ0j02oSdCjeZcDiK0mhg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="O2lxh5dPCBAEvRgYtH3MeaRT9LoHq87+zKw+oqWd9RE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
EJdmQAcBKdbIhCviGfMEixn1SH5jxp8oW/wRMAHa+BB4x/GBXcPpbVpQpLk1ALJytOM9zpQ1l4tT
HeHMGptSlmPfhu3x/3C9fjgINXFEnZGKg25fVcaX85GQFi6uRYwbYYhiZjyyOF9YZoZrKwtQzas2
fMhnRmy7+FYAUDUdEA0XYGL1oNuN4x4W7SznHDU3zQXdklHLV4ll/WbZ3z7DYQkxA+utMZqal6jT
XN+CJlLuOpixV94zCMn8mSQXgH+Z+aRLhwNPHE7iAwJIdoXLflO28xTJXfdcOF+3pXuRWA/uf3rW
Drn43qOnXh4KNgiP/80VdN9wjfwsHRgP1vZ1sQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="GbE8g7GymTqp6+WE/RYqJswsADnk8T/TfwunpjGfqyg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2512)
`protect data_block
hvhORLURDI+GEvJxBw5exDAxMFVC/3gVO2QCiyZxU51P9giC+kXQLxYbJyfhtUqXIkgUHlJpTFw3
FrtAI9ESbMdYLaiQTWUk+wRvnxUDyONept6RIh37m9vPWPtMx1FKPOyDYiOjxLCsk1v6T7py3cf+
/KDtcMGc547xe2JivIEwYZzq7a7TXQtzSuN+P9sc+Jc+WY0n6cdFc1MlrDoz1teQ+ao/qZl+EYkv
wGIjDWQIBn/DwbbU9DiylpAcYbScdTrtYBZXTKb37CjsIjemBSK9VDY51qMl7uHi7xbjAfmO4VeW
sj6f6Zk/A1g32dz9r8ma0+ZY6DxGhiRtRR4FvgLGNUDWN0cb/rGWt50ykKqT/GlR5EADbgLV+QC0
AtFAd9FAvh2rEprVvWwlnwF1rh2BeAZ56gRrnAHLjPbSYqEg8ZdSmDgSjAccjTEiNFHXSFR3L9nW
sJglYNsv6/PZzQkfRZ6sAQvyR62ho6Mu9GLifQ7qdL6P4R5ObawjR8yXiX7Jcb2UpamNmYfA0uHB
1UgM7uAFRhKcx6fRWDyvnKk5FgGfYREsOsrHQzWTSaK+kUZpiBqEdiLaigIAr9di90pAmi3l+3/Q
IwYJm+vjVEBnb0KJsfA83xUAr2+4hU4gr5EjKKpH13sD5VVu8FiYnkhvVet8FJJDVIJ/wCaIjyUI
ItwUna9LLAF98Tkuy1RwgXbVE9ynU3JjMDdpLZG08OOgpiXOqvIOva/hhemogQBv2UK3LWhyMXm8
xu4nKSSf2EKq9Er38pXUtlb/AWs0V/8s5qChhXzyVjTM8wSvTWSIc0eR0pEg5NUL+kZG+e41Xz0p
cs17whvcpoaVZLZD/apIZcXvy41d2m/DZZ9LibL9mNIfT9vzbhQsf+oaBBt0RjJBNRlEYP9RIlmW
S2HVaLLFwyK5pyfFc2QVOqcX3r93vBqk+6GT9XIfj9xqqH8m5N2aj05bnbFSvbORsitxniLJin3x
0rnVmASCIEY0OCtzGGxJt1nOG4VSAojpa2y/jh/zvZ1IAD1emAQjLUT5+6vuT51Dg+SEVwhUKJcc
44HFqzxIR2H7h9SCC31lqx/uONlqNuoaEXOFrHfBNYxklwl7eH8+8yVHE6G7mBd+tAaVCzLoYngW
/mBYOVn1UKMRlOMIJHIdzI1nzOWF8alT2S6cAZFg7aYOEMRnKiOv4iIkrvoAOMlOWfNkQV1YaCMM
aAJ0x/s8dwT0BgC5Ms8w5XV8xRQTQ0oXvOJVihOLH6u8Qd/mOdeBgLOuzAnorqZ20tMxNITyXRz6
tv2Lg6Y2SH0N9FEGWfhH7PPrkh9lmbCZ4c/GEjsmXPSz01dtSllz1zyRjPnvQSSbDBBJ7WG3SYJO
rPEV0n/0MSlgqCm/bdv4tyG9Ascrvt7mrougSd4LX6jAoVpUCheNNzEFpAIhis73gOe0qP2T1EaP
Pf3t+LuBU6ZOZi1yfQIfpgMOeXM1w4VYsveU7r3DTf/0SIId9zxQxY0PVGVy+vpS2SNgTZd3yUrZ
xKBVjU9qRD63uGczd4DKnky8Yi7Usyzfag7Jg+7Hsd+OKCmsdhzisY37G1O+pq3CSlkrMJzKw9Wx
JnAFrS8tmL/0NVdL7x953QHK09BOXI1mrbKmQyw3LNyO/DFnnDGRY+C65z6iEY8wgC+UbFjqrojV
mPX04X+HlBMxHoEk6+GIWQPdamAIti9quAGsxazm3+k0tqeks8bQS1brmfL55SavJn2PaE6S5twD
VHLf1e275ursyDUBOYOtET3Zvfr9DtR5y5D1eFghbVSSDJlI2FDxGfDYDgkCStTTUCBq9JEaOFQz
KnCFrMi+VFkzB2KiyQrIOl48TrrMy6ML9NN8DFsxibxKfVDTZuR100zhwNhrKX12eCnm6L+7PSl/
EQhoetpvfFEXS9k2cPpCOzd+RaJIIDgCehE207u0pAQ1R2QtWW7hLDB8YM7Qo5hKZlMAudT2WOXf
SuQMLjljCVhXb8PWl9RavEXMRp+qEfM4MU4ETAPc9aQJ4uYXbYk4GLIKRXs6b5hzq7wJhTuLGj0y
p5mM0WAvxy/YcQi2EF32SJVUzPqxUAHipQR1mtfr7WbhxxMhNqUhHUaDJwobxK6WyLCIk5fhl+nL
mugoc7D9cIatoQmj+JETZPzRuL/RPOy+GUIgaQSbh6yr0BLi5y3GZWykDRWhj7Pbdn4XM/0XNFoa
bMAlDfIhbXCYBl1+x8CVSjdqoAp21BFJzzrUHj1BbEwZLz76+Ko+j7y5YGWgqrqQNJnGshVyc2XA
1nnODx66gj9dw/5G94AOHWqOj4u8UhB747+KLgKMITbMIzbmRBoqsTamx2ZUhVqDTVdc/86T5UR4
+BkBGFsuhbGbIr2ix3zcSV6ZD9NLyxU1ya9USpqJZTeqHFFDIEk7zB0xLIn5sTuKLLR02mbxTy0s
jlIOyWyF0p7j4vddk0YlyOx0NkG36b/6WJ+x+N+nq/oImmAx4BxqCuFNET+Tc1/RMPy1Edow5k4e
zq/yXcakE7l8Epxs91JBPLcRuaF3YYkxIfsmnCwk98t0f889BJN51o2CggjneD8T9Ky2PNXPABTh
EPIVNkc8b6hFbyEOY2r9YlyQqNMT0/AK8YVS04tL7xWc0Qexx1KwJ/gdO9KCg8NJ9gWdKVzpmhi9
qKhFbZEnhd6a8UEIDN1i2Emm6Js557pcNhDrhOiNjQcUM/JlstCMTLuzIc/qXzk3HabPeivMq5b0
Xlh+qKYEKdw8oWCPqyTxDHKUWKhHlMMpzfv6knPwc3R5Z65chG7XS5b4kXpNkGMwsYy814KtbQxh
cxwJt9TmIlm7tV+0FLbwZ7BUqwLOm2D1rg/fhpOiyQ/seELkAgILxRDHVGBdJPieFXaYHZV15r6I
7djOOdeEUvid80oqKgBp2LGrl6lrRXespzfFmG+2bBhIhBEWqZcpJbHNZTYqJGY1XxrzKPBL2ILF
zNp7U0hYak2TLYrtNeSmPlmxlqK2vSH7JgKFw/sNLixsCLgGrceAuWqlCQQyf/kZ1hnJYh/KWfhV
gB/eNA6r1oiYIauSrN9SosD3hkG00MGWamBhon/XG3AKD5N7avcPypiBL3SIvs+vg1IQyxk1ZOjC
8k1UDyHI40vkrIK1H5X7q4Rv+0i89YGqmDsFvETTqi3Ta7NT0dw9qim50B48lZ9cRY+9uYUs8Qby
fx21v+SFpo9IIOX8HPm6K0M8h6BffoHlDQrvXWm5R9cNjGHiMJPfsumeD+uS/X+ruQGr929c6ZAC
TyAS0+cZSKAH4K9tu1iSMMZEGIfkb5bGpAWknrxKl8lBqYBE8fRWRpqXO2myjJL9WxCXwojQJbx4
LL30iw==
`protect end_protected
