--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
aRkN7IKmRxAfAyL6FBN+1C0z95hH4qoHN5Aj6OI8NqkTq/7ZBe4lqCNZhA35yZT1P2Drp4XIHVNv
smpjkcZviPGmOV0yeMxE5OEarYW9EH12rsimiEHwyGHkNTi0fwizEnjbhIa/q8TeY5Ehc36HABnq
Ae+B/DLlp8zHrNIauHJKNcjmGjbM3tQ4uqYRBndRN53+oYsfpJv1CHzUz3Ux+hWH8y20sbLJ3Xab
lbK6rluszUZgoa6xQc9/m9cbgYiNZgVqwuf54WuAoIXRtXLjHOorELXEZKyWFs3GTxah2SFnEaR0
bfXpqkuGZo396Ku8NlB/cfGLgWTfs2veBOL8gQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="M6bbGXfPFITLr/wEzZGZMWgj3bU2ZPMhfEwAa65/5dk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
So3DPFt30aO4b1DAeCZ7IATW/QzydN+qVyxPapKC8h8ZLXEGaQipqLj9xezPfam+TKd7oh3edpLT
yf122l7gHdNzZqr61SRM9tr+vNj2xzywQYoAdfj2f3SItnSGLMbFhsViv634Wmc3aQL5f0wyr2aL
PI4qHFdYS/gSiHe1cCZkMpcW0IaLzX6B385le0NUf0G5YJ/1W8J8syoRgxs/dNgoK3TkyprCHrfO
49bcfdTFPonBSGAX4qTHVQzPGfT0ImA5VmcCV8IspOV9IBVu7l9Ul9WdlDzblVGSPu2ACRf9ZhDS
6msaetDyIlU133pwrZcLn9tOISQQhjmUx6Z7UA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="tQzb8X9PpcdGNq2lWYmb+T4uMacubm8tXbaQbxMmLlw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14320)
`protect data_block
9yeQ06OVZ8vpgWAzLQCoqGpdHXy4WaxMJMfVl/U6QTcMzMAF0XknNSXvqEwessu7BimgX3YgGdOS
xoW0fEDTELgWIoRL6Lut6zuUyqVFildKzLfwfmEsN/6FRQI8wdc6jImN+aypPoK8KP2Fcc5qqOSk
ZqOiP/12Y08rz9u12+0tJ8grHTGgBROopA0ijw4qMoKwXyLVF0rDJGmFvy74g1xDWWuKQkGQ71j7
4ipv98U9PkaLX1JRKw9GVOhqZJ007MXeKdrru8w8V/daoMIjlW/aQRnO6MSJGHzQAaINonxqqRDi
WDRl/4DEW+Q8jlYddnlqeKF1MH2nvUoUjfbU8VEsiAbmDAnCWe5v4kpDV9nr2hlWIZ5mL81jjrId
JLjZA7ssfSzneWxRUX1mAx9cLgex1k+0NlvbbLNQw4aPB5X4j9At7e+23+nH5IcS9fpf5XnQBUG9
tte/TQ5b0e/sAtxpbtUIgPHyEYX+6gCtbOHjTswEyUgdX79D/wKXRKXRq04eIQbzy1tauTmN0LHX
PjVc8StLngjJw7HEkFuGSR9YglK+kqESQkgfs7ks2hXBEZoeXG2U2qMAxFn7t6LmgFu3OiitvAqB
f6FxQMafBe9iidMRGrRuqyLCRIMUqXEzsCk4MtEllzDuO25kMjFlHUO5GEswUCFmX7lDNwZ7w/Cz
vilkVedHIPXZZFd9H02xF4IVBVbvaBlSS+FeEVO0Zqe3kQQbx4+Os6BKAYgQF0Kz/9TU8ruG+qO3
8c9/dbXk5VQEQ5ieMFpniN910tnDiisfvH3kbwAdjNlBto5y+B8ZScZnla0G+yQJysRGTtlBSJ50
1pvW4lgZRQdH6HP4ImkVX8fjsJI9MMStzonu+KuEEaZBSP1bCsK6Z4Y8Wq7OOUOIvb60hcukdNbL
nu7Cvo+aeQMFVneGbNQm0m4QoT7NKNpiAD/egusvZbxEFEi54WKbsrtOj4U+mhiEd5ywl0dWfFpC
RCf0rUg2i3hRA1QTleux7Ev45Z9VcnYMLn1wlE5sCqJEDd/8xKG5emjl80fHHgfR7Dv4m7as80uX
gPaKIvnWbvWSECRNMaDswxOub3H2RXsoLbOfNkvV7tk6nQnpsbAoZo4jx6sUosUJmx8nXc0daqmO
+dVnuHADwdxmG1UhRX8mO6Ww01gEZPeHFuNsuY2mQxb8ogpw1WlFXVVind3BDzt0zS1XH09udqZf
8xb7N98Mza/fYnY/XDpvSPcc2XnpZyp+ScRplEGsH4N26M632aTrQfwtH+jyqAv9xwHffx79OuPT
m0gXPRZf/gtYdtQiyYgrEmLL9H8HpxZ1bcrBwHQxDVNnT03OLu0oZokEM8Sy0xaffodcDzL1NTsL
xivE59ZW86yUU53KoHyTvNzOapnKSntWwQ6IvRJ3K2bPFQp2iDw2tORXfn8aZ70vQXqzGNYHNXaG
JjnReszjGnVV2+tOq4dmnvn2vUOSbVljGgnr+MiAFpXQZv/g04n/vk0GWn2eD1MasNZ2U13chiXV
osb29FeCXruypjuQ00yXTIXyzWo8rur9ib4qJUI/b7af7sc0coyDagpq6lX43JkilF0x7D7FoU4k
0Lh/0xJkuhQHSeVVIO6UlR03zxwf7LX7pZxINy94rIv1Z4PwNX1r35PuM8LHsPwo/tw4GZ6Hf8Gu
QZRmSgzkXuA2F55AteC/PD5TcJQNtkDOrX3T3c8AwU/TE1+Ohsl8YLPGk5DFdcF9ypjlmIGfLFbO
cbB9OYXr3Y+XF2mIdlFCvVWsGFFBa0H3fiUdvak9jm1O/4HrxNqjaJRItM2ooBwfIUqH7jw6zaPy
yL8Ny3WS0Wblt0wivTNly3E2YsjWKzi1W9wU6ly6GFUPXDHvW4SRQPNxPHItMYQn+0XZxirnTXZq
VAPENQtq5CJHDyd/jnF9VxQ7cETSvtJ4vf3LvPerw8LHsRShHTMkFqyEHWN4cQQtICEjoRPPKhMb
k33vUbYWc5PdXkjedbAEUSKcmSNWxOOdOS5O18SfC9ynQehLKuhRiSECoWeZWt/KNU0GUBbhxeSx
1dZYL/YwX1cbNLqHCCpdZviHPbh4Iq1sT6AwWb7Fys9sKm+ZnYX0PUx/YhuCbbSQyWU7q9cO1QrY
cFbrNvPYZsmGLgjgY4rijJbggILDQcGHks8SHB4Mwb815h052gt4n9NzgFIDztfjdD29I304t9W3
VTiui6Mpe91e57Rw67fSugXPSg6KbXBv8EXhO+Rv/uv/DOGEc/66ietCZsNmqep65PJ6DepZVzbM
faon/MN87AZqHUevmhN9UmH+KCDrkJYyeNKfDTjdpqsDOdu08TyrK+GALx0L5Zu+NYnxxFiIPwbW
dXySdOkFDAy9C7E+xHKSCSfuHBsPkpYdVmml+YSZYjcrSdsW677WEsUqguiBt5OSVeSSYnKM/Zg7
2tItv3V7wvpnk42+ASP0X8BLt9zIK0NayAn4GN5Mt8WusEf2DbTl9E06//8ckx8oFYdXSipQ/kE+
0+QUoD8BWv4q3NJusbGl0vyjoByOQY3TWjFchZ1fH+scQWEl7bdrcFUy2dSp+ii+lnyzRpiXCPq9
1JbcN9ZZnwZznvpCroRQgKw1dt/BDoNRshHPql7Cm7dTt+j/ZFduFo5c291og6KHsPmsxQtoRc3W
XpKIODq/i2sZ26TmznbEFoNJBLhvo49XwzYiGcFAFRwSeC1skx91+DVC8rRbNDExTiQJGSlmzbTs
jM+21p/Ss0d7ypwituM9siCatCdvyjnBvAVKjQP76jK4+aA4TVebRXBJXmg75MP6zphvEnyBfsgY
TCth5RJ2t9x+LoUWitLqpmi5/W2FHO3T0t5yDp4JjKUAlnMHUwJnGtdEHmDadMl89KdSTlHe5k0u
mFveLx26dwqv3DZMPVQ+Hb2r+MME+s1V26d1xvF3AZkV8Ug11Ayk2KBobWPWp1goVxnAZq1jvzTW
q4VeBTryOkysvy0xvluj8Ka14ZetUYT/PlDXpL9NWety51gx5IG6cwV+lYz2Ji98ARXqteUyNvGh
LOaYcyCCJPpJvy/ZZtJsUWzW172LcwSV62g5qeTmS0GSfnq5jcaOPcW0eRRIZauJK+CgyoCl0oTT
ImqSOXt5PR/5zkjckJ4BK8+R+BDR92+ktz/iKSwQ50ocUYl8yUiItEQfgF8T2TI9tx/mChsrLADc
Xd4YXn5qraGIz4fp+XGvvF/PJD7tX7T4VGOr0e8PKrdedk+UmR6YEQ+UYpeaRyeLaxZuVuZz6/+R
+j73huVnOTk4uYCQsAYzJ+K4AuC5eQLUoWWkLN1juGgfRDcBxS0ecksrYku8QPloWnsTyRKUsp6O
XG7XW71koX+a5SZxhdJjKD5Dh6GEnwJCZrzSSTMSbYl2iZTcYtvFXGbo+D7JLNf1pZ8mY9Raeq7v
vaPHUa7YBM/qHLRlsSpMFxkX2TYpSfjtqh4H9JTJt9o+KrUN7hr1q7Bo8EC/KZhIN2RW7/XsQtra
8/uFfITsnMNBk+/ERIDeY/7P6r7FA0wFTlYoBcVuo5BJFRnXQdpsad+NoggYT/jFINWCZdQEd3UJ
nvlYsf1+2Sx8NVrHhVrTVrLzfi2kl889KBNCeOvUvcrKCxsu3EMGLa78AziEHw5u1hJyDudHEgk5
c8ZEmW44bOVp+l7lDM1mpGOvBPYxk8s+aW8L+aZy/RC3BXxNH1Y59L2WKQbAQ84QLvYv8VQ+/1id
1JqSmWo54EN5lkwHG2jicmdS4TZqLa7UXKisTva83HDmU68HTfaN4Ee1IHcEZgyOwpwOX2oK1oZg
tT9zei8JaOgXsM6WE/M49Mfe55VhzYoqDyYBS9Bzv6ikjZS541OPxdrAhxbyrxH1EzhyfrncVqzf
7+sJh3fRgepxK+MYGIMMK926w7rZ0fMLpUFDX8qE4w8y5sIh9ETBd+Np95fXhLgr6PY1RTlbSEeB
IWupav2/jGYjMIv3UZMZxrvY6F0vh1I8woX+WSm7xOkbOJJslrtQi28j/+sLV9HmQ5FV4qlImbGF
hXFomLF0x654B2ONPD7ze3DJgJ84GrDhCwQwUCkPyug+Sou2QCNG5dWE9+OUTbU/2lJbqY1QDZV3
LeJ4bscjyeqwC4XBp6EkLY2nb2MNXve7h7L9NVGr/2QLZfH6UGj5+VFEeBG30NYXGtPT13gQJzf1
m968I3QfA/eEy0/Yitqfq+glpcqVtF7D+0+z6RI98hJxEs6x6felXA8wL6Ow0UCw6/3B41nQ0ReG
twGvUCDBmkv/5HACNBmiwFkLnTGR8+l2bXBqE5PQR1PI9MYiJK6i0QV4ONkAo8WQ4UZjBdMwsOzo
APyo8YjOjimZ4O4QYvV/0KVqe0vEmUaQZ3lkoIxIsTyArjjDFW9/L90JWAql0iYkCJRh4FQhYkkP
vSuM9oEwtqPQ9SVxQN7B3jcLLG4Tdrf4a3wfOAhP3vqZlyO1Trp1YRVTedUkyzzVU0BYXP0A/zUj
qYsdXVo5VGJcPMvhlMqyet0jWbSCufEkiE68xP48pztVoP9aw7SVHSX3hLqG8aoLkgBbBStuS9Au
ftkxScBI76G3Q/sDVBEENw3yvDm/2rx1D1nBjv28VMRyqFUX+mtsxHYoGpPSEUQirhfmZ2gjtNQL
ih3CTmsdEsQCZy7JROOX8kqO4GD4OKvKPVbypFMXTKAmLzG/mkrVA6xfPioSChPwTGVrAg3evCEb
YsxBUviPxhX5c00KfP2GEYCN3h/tlnehMt154hwCvfYxj893dEaNJwewxoke0tqG+hhR6QqourES
iepG9PeItJqw70RL/YFzl/MIaI6Y3Ize2mXrNROPBmTYT3KGl0zil9qKPdP8ZVE8E1v4PXrK2Rkb
KGwiXrmAdyJoR6gXBXFGGiH+lRbBasthMLABQ40mRPrcoEUZP/vfOrLR6YmEUSZPuNAzETObTavJ
KYFBx5tOdxZsatMB0a6BJr48R3XVsJZ2WNoASBgxmhAFOVocsDQhBSY9oRJoL8bgdu7i/3l4FoO+
c005auTuljA3litLjM0OprQCLRw3TqdtKHrdFUvfvX9fNW2hUZfFvcNvybuR4UFBE0X7dbzUI5rt
ztbEfFwQsS8QzHXFkuTmb+A1PqFaM9k9Gb9B5R+QoRUOjus7ZvtF6IeshV2DElqSj3KO8WX1lo/T
ZUYkwPU+l90DsfpKdsbqrWqyJPHyNZKBLY71hf8dVgNp4Y5CpOnaEQs6nhrGxdCeFPa2scpSaA8K
83ayODeehvKEGCbJwjDiALfyduLE8WOKDtZCQIppA89rS/ccz3xsdBMSZ3NeAz4IuyJ5lZCEdnF+
ajSM0Xu0T35PdcrO+mmNLYCUAJbeaGWPV7g4FElTz/bgMKUEn4ul19Th7NYgxqdSj0qTPmmzKzy9
79OVc0ABimf1Y4EO1JLmBPkYrDx3O5qjeJu2BOIKk9aBCnolZ826usgGqsycT8w1TEx/5NyMe/UK
h53VrdhRP/8OeWap5NAf5Dnms2AkDSnBRYrvJp9Y91KUgqxBAct/gdODSLULD5KfzuO/tZqe91qB
uaHLtIoAJEN6yDo5MmvPf6c7KbrHKo8WHQ9mycD3d1PhLJwajnyp7yC4nD+BPTDihSC4xDEnnT/9
accA4O2xuwjVUAFncrGSx7GAf+P2c10uxXJtO3Zzytesb2uYYIGzTjejW5e2c30EMKO5JCT9hgTG
QSDIliU3LKcN03iF8HVmWqZD9zMS7D7OZ+nld4tXqwIdqh2hb93ykb/qewvZq1tj4a6PmKcVL2Zp
oUGUOmf7ctwKyNSecQSqqqTOcXOwPkoXvlO4UzgL7CZ447NidX6PgVXoulTDGJRlDOqipyesli/X
vbw2pXoThgAIberN6d6k8ZjaWVLlL44eUToY7YI9coSNyBOfksrHJdEBgAnHvK9G4qzpga3aUwhf
hDyOFQY9OfUZNla94flcyn/YjN4CYnMrlxB9TONBcJzIIgFyFuLeEVp2VrHpYmgTLsNkIwQuhpDZ
hGqvXrpnGMqpbl0x8Dv4Ynic7c8aMR4H/RSwXedadZbrCyNgUNIGu/Ca4maf9w04CWdSXhfJK+r1
c/oIhKLrQKETBXPUzRnd5JgYKREJgfP2XsNsemGd67M6jUr+XLb/xjAej6hLgeQHGJpcDFUaSXVJ
sXpSFQ5glznMGWdS2o92aOzNI81XPC54vmP58M2HBFb575eBKoOdUERITql9yzyzfRbe9CETlwQz
qsKZLD/zg3Szq8UTZlP3+wIXC0MN+QeIU3vJfN4YwG1Gyca1QGQfhGNIPn2SLQ99IHXdpgBm1/Q0
pGj9ANs8TIys/CywKouP3BCiO8RkKBO2J181EN9yzHI48wvYjPwrzNpvZt6j5EAEijiiw2dx2lew
kbCwrfvcrC2FEeRPOMkQDkYr+bX0DUWkgcPMzFiHVfpjoKb7AP5jsby9/mzkLsi4hGHbeoJ4OeBy
ZR1eoYQVEbgHDfulhDPO5gAWYHOLBT1HxfIaIV0QEz8RFXEgnuX4a3rgsJEpSkUQ0Y+kX8QnTTiV
r7vJigGeDtfdLQW8SOQ7pGVbKeKMahtpeVgz6/zKnILEHQWV3SprDv/6D9T2M5HqdQkDKz13ILmQ
IKmDS7gEyOakPjIF1CIxq4f1j5d1nu48Ng5i84/cgUlmu3P/UgAAo0xBoiTQ3rfSjCq3FFimuksz
yDtO7Yxa+HYmTgu9Y6JXjTUPuNfej+OXGnWq9sI9ljNneYtiD53D2TlihYU2sYpax1gmDdQKiZ+y
y3p9/lcIKqtAaRv2wg/NXA4QmdttTe00uwi3jdG9RPridE8APkQARxaXXehzSKLcH0mps0btPCvr
zAyieqkUa3vANtOCVI4LCuX9DHHd1pXHgLVuw+HLyKkpKStvl79JeXm/aY1fva+xCwcXTnsAoTIU
Hw12sxJ8iQkYltzHzDKTyWPTxpqD2cmUa7gc3pNtZniupncuCAmYv0zaRfD5eXQ9kyboso5gf+et
IUV+IvXh9lQf0VvnHgEw1Q5D0V/6VT5wnZUS56kiEsl2qc1ZVGvg+jfJQpFa7aT9nX+MczpgKE7O
vItWXpsD3Gsmg9J1vk0EoPX6cg2sKMC/4QN5VBq0DId8CLWF2zL4lkp+C8wTCbF6ME6+Otwa1+Ym
Nwbca3iz52vShpCQ0uhGPes+wHLZCrMwY5JciMcI7GOTxqUavwR3WirW6rK7u0D3PsrSb4MUbe4L
gsdUbKc1xO0N6DGOneV9RaG21wJdTw50p21GvLYApO/qfxXwXHfb1YhyfaP8UnlYc5gXkoIDW45o
chm0lpkTthZVM4Pam89W2YedHLOo7G1Ap847V1TKJ3/7jzm2fC/Oax3BW5+CwHRM+BJFHdsnuC+i
hPBVLGUw7yHUADIQ8WcJO3wtKdsVFJWMVJk3uMcN1zNQrH50dICd83CFw82QLXlO8AL2WX3xW6UE
C12YT6/7HKfWyB6yRUSZaJeIwAygz15LP5/1OQ6L3ceL5CoK6EYlCexMveSWSQMtXkXYNLiDcML9
Ya+FLbUZZ6KtDa/hzsPPKnX2uyiMe2ZVnP33r3gHHt2npwZjJF5KkEeDtlQU06OVfrdbh/UI0Z7r
atnjNqTTSwGD4w0s/GGmY6BNxOSYBSM1QgzWw8M0zcVV5rsej4UzRDOf2vAz4RCtEdP6vcxUW5Ny
gsL2C5RBPdfyW4hn3bjx5pDgFAL7ap9fogB7OLuPSAo4DvcCJxzOGbU5eTEJFFpzcgiA63Lf49Sp
mCFVDNQQGEzS2MIHtADCK6x5YLX1u9sJ9op4yPdZ2oQsVL5C2nW8XloS7aFR6f41hhF5WrNeTZ/g
eHJslIe8sVXwoZEBiKFeO/LX5U7G4ZkkxxdLJ8e9FLEVdW9u2I8i8cUfzc153Q8GFtvIVPH0t2Pt
gFiSqO3T1CwNrZzHMUj2ZJ/qi92C/UBsjS6iKZfoVhntbyl4tzfJrczGjywKekIrpxL2A67DZK09
gFGK2riF/kINrjcoQn1Apg1wxyvdO4L9Rd3wF8dgZHMCY8LvIJRHR2rgrWnhUEhvpJRBAR5KZTqX
z2e/SpDh7RbACCUXvR4GvCb5d5BSqAAZAbU1QFh+losYeCxZ/xNPQsdPOYCwJXLVZ8whZm0vTCAL
6Y2KSSQE7A87GQrZ6Xfzw7WXC/q31TsiEk2hgOPW8SS62dBBSu6T+qwsKFDaBw663bQJ1brNJff1
4Dpm6T0BiWTaxJrLZX8KrL0P0Kpsg79m59v9j3N/DknCT0jmVHr6QTH18eNpZOvZe0X67mNjsQrg
FGjQhi9C5gHnpkuLgqX9WE4FsKCJXqmkj8GFaqsVyUb5LjV3amP6Yp6rolgrPNTgodHf5x8HiqSI
6ibDrRqi8DHBuKAyHIdBlcw/pwWkUL2W8PqX6lQvSIRg0HaCJNznQD5HuDccZ6x+xKO6YboiuiDZ
w03wwZMducBeIRxaFxRMDk4WNwgv/zxWNvv08TxGIUE08ALg5rLgXwLRpBqftVkQOUiU9GwdRfmE
EOtSQHttOn4tohAJzIESmtYNTOzf8FvXy1QKtT2HbUsVOIUwDbJMbW0VwFEHiqmgMrN1RCf5ii+/
ZD2dO3WwpsTpaOtxumnrFlu+Yv+8JX9WpmOvebL5k0HsDWCtO7ShqYc9RwMhJwDdOK4XBwWTAmpC
w23XCgTrFPpjwSgqQKkM2BiF5hztjszgcFT032olIqwsvho75BjoI1mu9BHyzzO1rERvYkt6Ib1c
+L0Ie2b1tsWPHio5kf/VMnEGzm2ivB7meKUi9GXlWhiirtMhQpztt74hy5S77z4CidkP5i3JU7Rz
aEiaHe0PP0yLlo455BERidQ8RRp7MYUsQVBnz+RvSYPACfmoSQzTPUvbPzNk3UFJ5ZxyoQwx3j0Q
NdKCfjXO+ceYyT1QDFJ4sv8QrMKYwgiRL5uB25EXL66j35OZmHu5btiL+9iF7/dX5ThQQDeQCGkx
l2k4lrRz3QLlGqkw8XCcn70ezeKvf1bsHQLAi31PzPPWD7vG5tx9bEnheMlrEsNIqU7c7kGqN3Jm
rYKgfMl2BLDuc4cUV96zdXgojsb0y1GfgB1XgHAie6ssTIK46Q/+VxejziqI4jihcqz4XkfaUdAu
dXkB5YySRT6BN414z0zPwZzNavFzmHyqNrxmCPHl6FqWOKATwY5FmobYoNtufJ+0ggcv+KJDgGJr
FrDx+6+9UkxCaIrn4aj7wpCSRZqGatBSr4tbdNWSxMBy5t/WnOZouTwtcwAUa1ADxLUUECZ/Qynj
ABkgOyxfokjDtBrULmKSIYC6HgkpFfgr3FQ+Kwe1C9lfuCcUv31BhBHEN5qx4vNZF9rHkV1yK1MG
rVeNEaYrNYiU4v3RUHSuRoZzhPEnZTavCXCLFzovaS8ht8bQs1bvpLDx1fbtFbkHdiTGIpPFphRz
SARo29GyZAxFktLTvhOJfOjknWmFp777ReIfjlM++4XZ4vGaElqktMD/Q3hfKudN3/6yzb/yCPN7
tECfd4PfytkPHjGsCwGP8YMqdFVmkGwh2EgxoD4FeKSo3aeGv3CutxQUcif1a0ifagDDuOpmFsIg
3Z2J4rF32jXZRFTFnGh9/SNiGoBBWbOWs+ge3+kE8AKEZacN/NHzvojJ4slEdKosZ9ix9BQg2dtP
qpgcXHpiaxZRtHGGKRIhN2XiMR3LphS1FuR8SETZJSB7r69D/nCQmOuc6r/OwhuPj0t5T9/rWdXp
AKkw7HGzoMsXI2NfOsPYKElTWMlWw1JlqI8EjyKgrWupCHJP8Y4sO+YWQ3+VaPQbB4/ByAZXH3fw
Hu/3qcu7XcvHEEHmocg0TLDf98bhBXN4fZBpo0Kp7NchI1IaPFmRSpIFM6Z4wiWOf4rmcnqo1tNy
np50Fxyx9fLZgJDrNBn2SadDjQCL9E2M7WLn5WHlb94MyGzoVHyGPUXzIvjymXGyx4P5XedAcN2e
SvJo0x/DAmjQ+R2W7Y9eDKvs+x2SsDuOVnLpp79Trt+LW5z5xm2uXacpIStU9Iv00nwLRC37iXFu
R4asB2wiVCivUa0wf48sWGhvbPzVQPVRTURgoPNhwswTYOUiy3GXdpt8Z0euu/avttXuX6xIOPsF
Lt4ups6k/PoCy6nkzsD4MG4Ar5vzb72PeyPnQCT5TzS3a4r40HW80Lkr7gLabdTfgkvd0KN+72md
vw4JnZ06xlGUy8lNS96sY6AuOPt5t+O6pOmQHk2gtJ6vKlQm6es34lxBu2N1pKmw85Bh+AIrANub
mn6KGRRswx5D9qVBqsdBd+VNrBbiXDZkNwqWn4/Vymf88aUE254ReRLNxNCwpQMNaZ8FoTH9PF9m
XJS1dELOOjuYqxYQF1zpDTQ43DRMwvWnPayIgS7GeomUzodedgTaEIOvarph44BnW7cFSj8cKnwW
7+8ohLjVFVutmcDdPHmb1kdKj8XGXx0NKNc2fqz8Dyw7DDldOsRiJfCkbPiduPjs9Fjib4d8oguC
F+Cfvee5LYemeraSAMQSq0J2tvr+Dhi2VeiFdHmRmFqulccQ8XqpNwIqT3VOw16Dh4hSrqAvehPe
F/eY7JhmO3La1/1ngsTa9LWbL3aLq91hdMvZFWf4TqgAbKdyJGvB4soI3yzzYARlF7JoyAzQQjop
Ovxb4JzAvdCxROmyUu5ZrOy8aHTEL+8hU4Ga80gH5KZKyn8u5CwzzmLhfNwMqfTDqqKZH5IdMnTD
aIXWYGHuMpYViylGR0iO4ql6ESSVRdCIPB3rgg0rV0L+golKcepzg34QK6RXWhmoc9C6XT940iQf
zSInv4VYskde9WrhEvX9ooS5db8/XdMVbuOaicKkEAux8U0ST5YfeduK4qdGwv6zAKYaz2Jmxei7
wAGfqSDfm0Wywn30tVJRgligfeF4Lyn5Mq5XWEUcSNKD1KpoGRFtJs9jYsiydQtoXEFn7WZ4QIiZ
Z6lO0LsxjmjUACi7YhgMSfRQ21irDHov7J9pui5pJnSn2KBv8tV2YXUxG4J3JcmAYYMgvFm7MQJF
kSjhNYJt9CwDdK5CAw30hU2zT5F9WCykLqNBZejSOZ06/R06MIu3qVctFgG3SWeDOyyd2bX761SP
SGiW8GRnU5qyxoGAanEQy+Gcm6dzkdd11LE+xBUoql5L/SMxwzm8G9POFP2jNk7J2i8R9aIUtKfK
91/m/hj03C9siDZyTWPKVvh2Sm6LEbIH0eYTwkSHO1WtJXT9EKgQ7VwIplNq3bHQCt/VOypUxj35
/YGDqcibwesZ3eNUmJDwDtKGfOmg/hyOs+iF6Q66teXayKkNRj8VmUIGj5Sc35B6kw2UZdws07ra
uvN9zf82wg6UwoH0ScRVHgjmvc8x46tBFytzSO+c8z97DrWB6Zm7eD4gmcPIPFxlXPsuhHcsz8hP
YnAQvKSPzB5XA3hPCSszOya+407oH8jNckeIoQtMWD7VnTJed9gkheHHmttExHFsPSG/j5LS2jrd
UsXi1sUbxAuZiBkjSi+O9i9VUdAvwGGpXGS06Jeocs7VcCkXx8lIW5ElK4KHACQMHC8cg72bk0qy
cUaBwFUyx0FD44MEBH6/79LpNrv58af+JpdUG+srCLkCRPy4lnSgZ25QWq9JtS4Sc/mXgxli6vj+
oAmRck4KY2Vpwu0+iEH0OFszl+iVxFrh2KFCgJyZ4Q86FnYeZUcGc9uH4PciqWxq0vvmADxaFb1b
BWphjVcvcp25kOXoeTKYu/k8u0okL6lOkubMoDU9Ww/GzXnzVIxE2fjeJ4AHeNAjtYoVZi7CK/Xs
I4bCfiNWOlx3LpprWxEjYG6ndifTwEGJ+6/Ome18Wr4AFx1z1WgnpyxXWmAOyt9t6ZjJaKKVm2LA
EDWNCwieKOQ+bPKqUV/8oH7hiNCVuqt2jyCwSezr/7xTgoAgYgsOWXYuzx9//XyozOJCLwatb0ft
/soxtHyZT5Mqdj5bEoDAu8pZbkSjdzp5Pm8WQWRUsBK2CB1fkebUXE9mO4J1gIp6sFABdrEMChtr
esvlVVmaF9L8dQnGyuE8cSczAcZRbqIZM0mi7YzJ6ZReqfehYSfo4BDF2Es1WZR9owEDbsEh/A7v
xqtH4nexDeAH2ytI5IXbrqX36AKfIxyq82dSOTX8WRCzrqs1UdRxsQCEKZl30eHGGAIoQcB7QOIk
RKi694dxFre5oLUnh7r4f8LJAGXLvhTZPr3LGvbFvENKysb1HJ0RuInWhdox//jWBOyKRX9R6c2i
4G8y0GFDtjYQshIUEIeXt8SO5DpiEjqZkLe0PbfjpgD34IG3Gq7+jirc89Zq10FosJByzX/IlLiv
QeAumiQ12fg61pd3+fT90pCsPTMD+SQ2yK/CnbljHZBHDQbhYa/0pMnd6TGzrTsi1J4KKXyjK4nn
4lbtmoPW5LrzVP39kW8t4cW0/OTQwjW60UJqvTQ5v8ZF/LR97lcMRmVFXd32rt2RCmF+4RibJ/x4
d4PzrXgI4eybBktxVtXcf2p2tbo0ocsmVXmOcQ3zAehl0ZKqIaJpc05VXvON0Fs/ouGJghtMqyi6
d36/VDQKIYbS249IaoltDNHnGuNN7EI3Hug2IecNH6H0DNFFxzfQ64oODcSFNXnpNmmoj6lgnx7c
GwDh3wKuAxioEXLewFWYfobSDtmfOZgNtXiTW6+V7GQEPa6HTpwShzFAvI0Nuq1gDpln1mCPd1XG
dTYZXomL/SIoyoMXH8Bw7R4pYUypKmWIUhu8i3SG+xOciRfTbp5kGGcWouZoFXlDMjsgj7r2Oq+Z
oPJOn9kLHIpCe2PJVHUp/um1Bl0EcSSLxFFjj75m1kUEB2rVTtZdobEIuGXo8Dyb8YRsq9NrkFXS
FML1t+HW8GT4nrocCCgixt/a5RJWEzGtuL/H+p0HfzLgPluQwcfp3wK0UGIDqGBx0Vn9Asqydpz+
X5d07Abem8Aj6MW7V6Ba9KMiTvC6lVe6SVMNyB411d9Xk666DiRHTLxwxXC9dpDo6OJ7AY6BIP8E
14TzjhVbLCpNf/RKw4WFcuelyfv/wY/FDFUsOsasENgUlsQcV5zOIiFVAyUCBB/ACfQ9UMnlctGo
PUV37QXkoiKOuQrTxnaymho+i7tA+tp1TzdFos0/trpaC2hS3TVHJAdJbpq/JdXtPYlypwN+XmFN
rVelaxKB/pveHt0GAvp4HQBWvGJQsdABKvndc6Q3j8LV2bIHJWl2vOan00eCfzd1tO/syj2KYD0g
1OhmdEeeSUwgXhb2s6+oydcyhYJEr9gWLkVCDI5Nw+hXijV3fU4Q97gjKpd/bULnRIxB4RINWP1I
+9R+PyS2TUwRIsqngqs5KyB5k2s2DsqDgGGCv0TQeLG2wvHsr7OQlpKcq40GWwLjXTE44SqvYcJT
GK2bX8qyqQiGWnOVXBOSKhINfbCyZZ0KeXTHZgSTbN+jVY82xShvSndCpDni4IWeItEF9B/Ikca5
N14FnoYMeqxXgBLi0PDZCzgAvgB4BYm/wN5tps7c71uYrLHhbP63IuwYN8+zKidjUBdgmPbcpPFh
CDb7oS+Pl85/csSNWltLiZ5YWrUHHWCYrguCBekJxElOMrxJmIGllF5rvAp/GNISb0Rz7uJW1ue5
kclet8RkWlhOcY8vNIKSNVXYnKBZ5Snp+Ek9GTk9+ZSyU2Uejx7WKwV06Dq0cXluqqcktS8f8sBI
jn9IH0WxuhYX1DzH8X1WOW+449sDcJN94h1JKwcQLl+7bfXjckD99Yj736o/RumeeOHYfwHSKpvq
8bBX5P/1ZkqDmqYCWV0xFw116tp77iuz2QnRpj0rr9OPWmP5NFdct6plmzTXwv4QOWjhc96S9YsI
qpHequIBE2nZ22zpI06nrlmh1pY04Ml0LbsmhndTCurEQhpIETKzyZuzR5sJG2dVRWztkkrlI8QC
EcHeQ6ooiql0UNTieXrqvhV2LZCTYaxezg+5oFVotnfNrXW9qPgvWDxQukqdj4BwMtuGbGKL0UcT
myeupQCwcmRwofUB4fWfLijXsSRtmBpTrDo9srk5bcn4FvC1B/Ihg00xz8lhi7exkm8XL3mjy09z
aziNu+mMoOKVi6exI0dWaE2GHWIR7H8QgiyR52qA7afEV5vrildQfrwe1qec4cqYowf1QJqi0yiw
ctlfY4kN/eLd0LxiMEUd/YYhZ/6Y2L7O6NlIi958/4o4zS+YC6/ktme5uf/u0p/pq+6oF2pxxI4T
OAgmkFXKkZY0ytD4O+E/E9T13kgHCz39idCTPXwTODWIFe36vXdUP9p3l+R+bw+I9ta7mh3Y15MX
rOCxOG407H03VSBJvMJTHs3mmaydl5MV9u/ZB+hQk4B5Y3KD7da/3MvfoOhdNAUW5pUQW7nIxB1p
voyWPACuX3XFxR7y1pMg37t3uNRN54ICu8HaYWTKyCfKn3r7wpc7TOLQcw6mrZfwmKr8n7RN7e4w
3iuH7YMmVEX+5vKi+xqPVeM8DrLRD954oFl1pbVKLJorLy0QhAJvoEyLjM5VePgz7RaGbMhQYI+K
Aaw/ywsKINZ8J+SzSIhGG7LThkJRa5yrL9odVJyxHeB52Ojx0q82YTMm5A22bB42uiACW48nm2/8
gMRp5TvUZ1sENzvJNcBLGShTKO1oeL77oRtXU9bhVG//zCC7lf3BGFhhjeumVFhy/vMeCL4pVIXQ
mftaEqTOz5RYvoiiRof2k1m7QDV95CyBSVr186ntE/dsV5UtUwRmlLbBCmbBG4gdS0OkLwiLMlLU
0xFmcxk7QHWJcd7+f/eEvwpzveS5MalXdX15NNEc+NYGhLwmYXqVz/C09fSQSReGrpn0HcJezFjc
++CqyYnnF4f3cUn1KE15JQRnAzZgN/yRD+2YuzUGMylyLJKKgyZN1aIugnO8Od/+FOD+V/w5Vsoi
A9TuTCeCOjEsuv9fiGwLXS4x1DL4+pHLfD/Haken73Srvnkeq1ghNXYTgI7WXJMrE77x2kIVKwpE
tVqrIr86OHXtYwArLFcIClh+70vAmHQgqF14E8bYtfM9ZOb1PVnjha9bkgNnso9aDuCdRyTQ7QhU
/UohxUXGoaInu1bULxWce8NpQ+9G3QcPt/2MCsi+BsmJpzF/QkYu6h5uCJQhielO67GxhNrhsfrz
9yjG1y3fyzOIkLzwC83q4jhOw/Wejr1oHPfLWz8s6iJKWq9QLiwWhZt3b3FIG5I7yoT/8O3GtghQ
pwVrgfolZvnAh7I1Q+wr6/hL1QEPXox3jYHjhziT4diunrjz+NOO66F53Zdys5qNecQ0o/zYzFny
safaFO9syJiFPqv+ATUFsiF/278hK1jrOK32UWIIs2uL03wvOKsyh+cO5d/W+cYC9mV/FYeHxGwU
ab0iFXsb8iK0t131ycYrFm8p1Pe7BiPksaNX8E2lbWKL6pfcSLk2iIr24nIJZd4oGYo2AGOTXEud
48lMaLZioyfwuWNJP3LgjVm0tZuNOMvyY3+66wGQ5EkkLesbSkUWHPhu7pLtqIfAX4BA5DRS/0D3
maQk/T4zxC4mf86vVORESg9fV22UkUHdLNrecqa9g2+yMrOmNgR8Yf8rDGBRHpyai3YZmOcmVU8o
9ZFP1iozpRggHuOqtv6ZVn31tFuBn1CtJ2IfCTeQPE+O4PkH4/umwjcM1lsWypw8HIGLnLXZVqIO
G4bdMDaaIIQ7nx7TF1SYCwU3aF+qhzb5e4aMAppBxTyzazkULw57gHJtobWLmjEIi5J1twhEPHGD
n7Yn+JjdB2e2HkOQG79Lz9ss9xo0e/1F7OR+HALS6cO7l2+wxPZzmo8f2yOblTGuPgunzz6S3ax3
LDtY8Zgsoyar+EzGN5LI2v3yTq9UM5p6/8uUBZKW+CQql5nrpp121wjVV+5qUn/0WUJkRI9++9KQ
nDvnP/5tkyTkaMcmcRaFQuecgZZYedZfRNJvGGT3zsa89a4xZx/tLeLmM0wSBI9tzOlLA4EVNHKm
5CcKjXG1FPTP2U0BzOGDsAg4Xw1vETK8CCgPcuAxNgeCIww8Y8GPmXDVaiESEGUSmYVUuyPmz1vl
s10mXhR6T0u1I4di82QZrRlT+GgIQyPWEKgsk7ES8yAe/2MgkrBetmS5OElrBUVJWhFdni5jUAxM
YEoPl8U+BdH9j7jahDxP5WNVASQXbWW80LuYn1xGDVwxxiBvN2VwNu/G1OE38ITOM3FBnUdjvNwc
0rwMv8/7kJYuANochXIcTbU8UVIecDN8VOmLmwIKXTGzDIdzzsvCDX1ZvzUSEfsoNKS0W5fBP4zW
+vwcUq4gNPwTS0QpTCdawWspr35UplJskx9lcu0vhouyqI3IGSXyIEWdcqCeWSXQI+0aYa9QgTkG
jtp0NomFo+4uJJ5YvaYJdAfxZPZ/WYKJS2JsRJhnE2kMlAA2AURPUs00GWNmjfVKE4lLwkTplY8s
anbeGXEtlEluJJhlQujc3BW6fNRVsGQzQ03mV+v01LayrmrzhYug16JmqI6jlk/Gjn/K3eUGsxmC
L4YH3gJ0Oh+kTw0kvosEhhKAnQv1MIyh+fbI6t2uVWI5RUWnNqJIFRv+6qfQeWQ83vhUW2BbD9X5
/fYBsMH/LlTf5j8/yupib4Bp4E4C0+DPjd9xyioawYighSmGjfX5WHUKLaqE/TPJ0BC4f/aqw7Vy
iwrE/UOJRCTQnU5XLoIyAIcWI/0yS+OHZvK2l5kscx6ywOvbjhneakKDDVw+6bxJGFF2dp4rNvnJ
voI6oDnNBhEfHkm82QGxGiRaoLqAWehLsXqKp//657YxfWkHoW2qXLPkWYGUoeb0Tja18sQfyBbk
K0C8Z6fxCl+bh/0TtgDbBfcBKF3pApbViXcWkSymCp00Dw7hOz6Ztzu93fJVJVSbI0FIh9/41/jj
ObzezFS641VOHRNE1tVhEWgZwL2b4ZDsYjekDBFUEGq5RZ0fDoZ5K4JEjNtqLRpl1jlQbmdNCJlX
lm2mNgWuJXVbp8rrG3L0yscvSEYGIoScRQaGKNrkrt8E+JrYDzaJnCLYkZejSiiNwMQTjet7gjXh
EcAg67g4dYJFJbFXYcafFNTtLMPGk4EQREYMFtWDwu0Kb/M/u944TqUvBNx8JbfgLLaDsmOzj0y2
GkzIkLTYjMk7WcVkmM8vUr8s5Nmk4nOalcqjsFJS5QIGx6pgXd/nwXHccNEcbBPultp4+Mf8Nv4m
M3il3v03jvajCCgMtYpSUaHKE+TyX/OpwF9QHxKouulOkfdQhNeOMVX4/hr6hj9+xEcRn5oB+b82
eAihUfzvEZyM/R7aazJtzzau+wQzyfv2KCggbBHLBhqyC/DdsUG1Agsn8EbG5oopL9/irOKWbPte
9dpMs+MBlYVuFueqdnQQuOjkJu63A/fHLJAcC9nHVRvLfgzEykYoLb/+UxPfr+P0PBKL7AtvUZ0e
vs1pipA7NIDy/QOX6ZAq9dQqxZW7eIN2V4mdLVChl2L5vmj0opaBo7PJXs8yMwwNBA8gnPoAYmyd
HlvwjdOuz91ka5jDkx0IL5nKCCKjysSTfDgzSuISkCdXspK/nMpx9tDsAabvRwExxTZmqj6WTKaC
Y8VoVQW+PL5FtF+DcVpbHAiZo83gKDH/I3EwcR7aZfElQQqAzPqELsu16aDf0yEe3YaaoSCNf7Qx
MbslSpYn46Vqxv3i8i+BfdO2G6+4oftjCauifY8ghX3FMS+R0l8eL32v5PPffGmWzve7ug3MfxI2
u9476NyP1mVwTTgDd48SJAxpHcuO1WQHkuA/fL3z/BwRWG78x+u5QiJpwHiIuivR8eD2SnsleG+W
EHPlruooHWWaF0zKL/S1OndkIp7ZijGtM+NWnoeQhxRePYA9ha79i8R3Si/EoD1HjyQgZKksTGcB
eFSBX3vZA+eYcy+Ip+sNyZYMlSWcnIqdEvZq7mZwCAkpKdi6oYP7VmQlXy1yo+6dyz9H7bOf5OSi
bo0kBjWZtCfVfntw4JAE6BmPkLzJkCYqq6zUmYp9CbTPZ74NMVd2F7dYf8Dg+FsomK7f2YTe6yWI
Bv4JTlorpdAl59FXaTuzQE4HrXje9fGJvCWT+dFWD+uYjQH3qwhk2rZI5x3T053IkDYyEOa3olRb
UMA8Erl/llxx5qaZ7qAXDPCxjPnZNHhz+Grt2K+ZSIJX1v919N2CIEiAEI4pGuyg3RU0WzpBdT7J
MkiQPMHRUWD/gEkI05w5J4oRHT4qxR/qHpcW27lmt0JW3hU5I3K2ZKNjnxsqmVkg3SQOxZ+0r12t
7nccuHJPUsnd/4TE7dDvGnoF2z1WdtLIb6yBRaQ5QUUvK9zvpnXfEi0RbpjEGoue89txSOevD4ZG
2q46dGgfHCLwJbrTw/6/f6SgoqD/3xsKsEKyf9C66lEkxJpayHg0DcUS1QTFiFJj75+2U3B6LuwQ
KimJaI8Zjcjp3TclQd27eIEDI9qDSXkKqzowvgKYLSBQCa1+bXLRYuFwC9/1iYfhMYed1Wrdi+Y1
PW5JlouX6lHXIBJLbZf006brPNlYTlRU/+oKlNJu0HnNTjVSk94UXu3uv8l3tuXX0OquRQP4iJiL
gaQKtVivba9LLcRKcq2M67eMUPVF3bj1r5UJkNY/S1X6DpijJn1CoOV8v3K7qqR6uiZZcaPQQBQ5
2d1mN1ZmJBPwiXJ2dRz2C1OryMVFJQx5JSQMNGR97Dbh/3qm0Y0uTXibx7b6bC8wd0U4ydIBi4RU
S4QgPYMnmx/zme3RSe8BZvfp2/KK053Zgm1z63u8xyyaZpiplDXSUcvRlN021piE9N+5Ss1l7Hpi
xX4j47GzutQZRR6IQE72RejouNLqDiF7w3p3Bz7CKoG1F6HSB5q/vv96XSRBG5c2qXJgp4lDfs04
W3/NYJCWBypUtFmPblU/BikpUnL5MTulSk3d8NBFVjzjbTlsqcHtePSPaAPl2JTgrKGsfn2RX765
GxdiWhgQEliufgyiP8La+9WzOBKkTdICfQk//CeVAoLi1ctVnKh7cDVsIaEfb2U7olIpM5DJzl3q
SM4WinQgXhMPO/pbP6kn5jODhM6jnPH1S4asvwvowp1QgxwoGEF+IRD0yzUj2IC+nJoKK8rQhxlM
Mv6HPTsDREcsibYVZQ==
`protect end_protected
