--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
JEpFZBmLWzx8kjxz4M5Zz5TKdj7dX/xyBOmhl0/fRdjbggg5jGVWlNeJlLEt7AkEvEq+59aiusec
9O/kDgGJRb+PfmEdwxP/uw/rTKkQg3sju2QR8uFQtratea9+L761vITidXmgu5TSrbhTzGrZ1wIT
QB5gbmUcFC9zP38YH6nlJC3IZvjB6rOw7+Yj9ImIKALRhclus5TnJvVcMAabRSXE/r6xGUsp4Fgr
FQ6rqynEb0CoUc72C1WdIFCwlbDuE+N0oxYtwJ59DHJopSQiC1hNSsEuBsdBoryd/qUYYu6ZQbpf
w3dsZPiH1KbmDM4XRVR5Es9gDdwgtTk86j3pVA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="XG2rgB/3JHwiVrs8vP3GhpsPvDw2V3fi8J+sI54nil8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
TKhOeDtAK6yt1wRqpXKsWJrcERC1ePmcwRh4DkqXCqzNehiv8xNn8Hbkqws6EclWF324VbOy7kJl
1C9+f6PtaKC7k1+/FdIhrZCYfPFz1Itkoq6iHsqJoVsNvgPr1kJXgw3M2y7XvJJ+VxKKJhAWR43R
4wEIgZdkvPrjEAg1C8/ae340bRRikI5Au4COmG1XtougVtQGrW9wszxMsdL4aK6i6OaYLwNMrJI/
Tx8CVW6fGmLynatzwP5E6SsZBoTFNrgwZAIymujOgwT1iuf/8Lzktv/qr1xyzNHOwn/P/OI2ZRA0
FBIjQzfwTmJ4VhU1uODHQ6INN3n663R4LZfZEw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="3sRdc7HSqMxPnlE4mMufaQqTyGlLbG+JclbDbi+UMMo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17888)
`protect data_block
CIYNv3TgypRPmQTzs1qEl+Vg6LN6Zn/Aekrfw5Mi88m8yDfi3neGb06YcPZtflBh7B6u8eI9JmW7
NPcFj1ohG1WBjb1olHSkbjn34sDFXb1IcyYwndSq/uIM5bMYqtC27q5TBTAxwciPatUkFKa97wFH
1a6KrWBtZ6UAVr/elejBkwyvNfjdNh9unKf9v7nggLFuz7Ell5Jw59VLyUBvpMTSr2fSkktaUDXQ
Pc4OQJUkY6UJACogkSL9s91Wf5+V6NfsV+ISpvI8ZEuW/KgnlIh0N686rzV/DPFTOjPl51EiFBAg
wwpFLXHzhNYmZQAMQ87lHc4KMoY9I8Hzbd9qm8fnw/EpCBxuV/4sFmCNao0FpH3nkp3pwNFGkXVl
7AykyX+y/Cu9VuGrWQXOnSEZFcNGcYbj1IFmq5GvszWJw6RPKcxolhAVMYU0T6yq6reei9dNVlL8
DlcmHm7++vT9BM8qTIalAykZX4ZZVxSSX7SU4Sm2mK4T1a374eDq4+ZL9o3vTed5Oqgt7hQwBgAs
O4rjvciujks7kYVYDcOdZovN0Ekf2YIJkmqEtRZmmDMyDQavtMHQE706DhIwpgqAZCt368Fk0/dO
o0A2pOO3uNzz70DuqYzym7HUQvsbL7W9XH76sc8lqOzudR1Rc3eII02jgGEFEv9BO1/coRJyLMx4
ayN26l0Xhx11PahC9uf9Z2yiPXMFhN183/4HT9EsHh5teW5Ay9gmXCpJYYfzlJiSfNY7Lonf7yjk
iCZTJbyEBiQFVkjcJviCGJxeLelIQE8SP3db77bwCaROLCN4KV8f2oiDr8W/DtZv6wT2vjyIEq/U
sy829jX/hxYzsAzk8vBoqEfBRZttJtsSj9yzecT1hyL4sp0w4fbzc+cvMKq6HxM18/F0EPu/oGlN
lraSdtcOLsbB5Hb9VlADpA2VytWCfGkpRD9JOoL4RYnX06QZFN1xMK4OhHXclfkm5mgR/U+gcS6i
uclgz1Vp+bW4cX6Kj8dumJ6Dnvtqjmr1BIgzjHVSjdcITiV9jn26iunWAQD2gfuhwhECuMf8SX5A
2vzKTp0QxGvIc4HN6nx5ogc66ZhCeX5gYUITXysDTbEKoYZZcj+D136YIvRrQle3IKkBvuM0tXzF
uhTqM+R3aUlFPHd+Xgp4iYy0nloFiAFiVxPGKv41Jd429XpRDOqhD/486Wn1itebpad700bhUi9K
D5s418Dxztv5g8XofONnN2iLFW/jeonvbW0xaHQTcexkz7en1/IO9NcUhEQhP4KzLfabvhsh7bv4
93y6HVbRPyA+SJUPmq1soXVwSFjMhF4GOH5Nfid1v8siH6TApfPBmdgeS2nMaa4+ryrkohGsi9wa
MUAGxUdMS2nJdTatMgE0xgbKzmarbCbEqmm+AKglO3kCJdj4/L4UTGZgQU3T7mzDVrdd+zPUyZ8r
Qcy2IdELCHsRFT+0yu1lDFMeVTc5DzWlET1XO4SVj53wlUL8dDiEW3LnM6HldilwTX4McYk+7TKe
aGQ43h3jmvPlgemBzH7sQW86jJM9XvA6cTUTSyxqmkvTwyrRfizmfiOnEIAjLsbz0AaxO/77Utfw
2bFJWS7b8AM551tc6m0/s+lTfJ4LrVzjpWZhPpq3GpAh5BNQSOBmZ4KbJWz2gbiVxygGBFM2B4js
4x/utF2Bi3u21RvjefXiTyPoBy8ZGqP6vQM1KCZlUDwuvsX/w+MrThNhRSYg0jtFjNbZpRKXODbD
V/oALV8C7s0npXOC5jCv++BsElrznieasyA1BvgEJgSJ4Ok8XKbxyHaRjx0qLtzDVN7Vw7P3e2VH
3OZAN7QrW8ysC8pmmMF70XnasKlTLBDspwqtfCjU2ZrbQpXGX98HeRN4QXfelg7Mn7GPqbM9Ocq9
AItzYBGNEnNjC2WVmJ7m7nw1+LqUIBFLZWWVsqZh1NcrhFacZTqVSubUlMWL6/qch0+DHR1QFelB
6iIijelo42FRj27wmqOtU2yYlsoEEZajic1K5ptQeBGt4RMcDrEupbHADl8sZVYkU1MqXjU3Uunc
jOTfR4ThTEPQ6v5ENXoScJbC/sasVPfsDsv9/gjk0k6X5HtGF1BnpWOii0sj4fQTGIOq7iVdzI9Z
gSNe1kCK45cj+YteQbTh3daaS3Jw5wW0DlN/AXWSBPsX3fD5YgI+rF1YKc51uLBpuae9KAXxDcRV
n00RzEURY+cR+6zRDmtsUN/J72joNVcNh/HGMl/HxCigRIDzWvtC8Vi6izao166TQKjemItFEtGb
vQXGOiTQg4C+zn7Zdq2p/nV+6MkIBet2fbf5byg4X22zxXVT/1aQykXYdO+UvCwC3mcf4V4fNkTa
fGhJdP2o2FWrRkduGO9jluuXYBu2M5wpSwV7YshQmskQmW27XgP5tF7oiqU+rnvZvWpbPPkr4x+h
siuPkY4mnMh0aTVRwpMlSYgi3JP5igOrB2z5paLJdRll4qBQKy19qNDs/E+RTEcnIjrX/oYTyzY7
hpofz8sIumzvLrmE1hTwArby+YXbG35jsBDP/JqH9d5fl4sYMQ3W6UsqTnOKpQjN9GJHekSELIHU
0u3iT05txTelDCY1a75Yd6K8kZt4q+KS1qSYvaxhH08xVhOaJVBigUKQwxkikhmlubWdesmDimFW
lOrXalO9oGOTT+68jEgxgPncK7Qw9S6BKkKMRMcuIJEUCw6GNyeF8LZbP2qZZmU9XcO8guX4hSoP
7PROjD2abcsfFX0JgaIIEjZeNuT/A75W7BCms16PSp7mTQkX/wjI97QY71rdP7VmOfSTgWlumYKe
wlrK5NQrkoqznE7KFrpGd9qSRgBRDdCxzQGz4Obyu54PIyCHaiRWhVwM3rk5mzrmx0sPlluTWAAg
omvPyaY0cQAjrwTIElF3OfpCLFx102s/aavi4mHfqDvCAuSfUMc2LoS6AzAVtmDeRbzEQYueiPgq
8CjqQ5P+Hpv6NQ/hb0FXkRc/EeauD+tpG8h3kuyRHeE05fXKcPDq6vUbsx+nOXN3CDVpIqTmcVNf
rdzaJeQVH8gk9o8YXvwb/UbFdWYzPlR6bt64DfGZ7FnHbS30QOJ8iL8rztztonZxYdiqjGdwruAv
mwxAEvev1TXe564rr8mUOFs15ZFTjN6IWJMR1bWl9yDExWu36VukMCPZ/gJ4uEcS3Zm55srfGBYw
gqSmcqeEKvTFgmN7GfnEF8UcSiXjyTCP5nyfPYPwYABVTz+ARwR25cqj7bmH7YbubhPDk0KTXB4c
OlJN/0cNSA/keZ6Y4Qxp1aPOjRM5tpVJjqOk5uGuQg4+KN5G2sYMzcjWGqFD9AK4u4J6LKcCrrNq
BfzBOPlQZ4XJz2vmriiZ/yeM7j7usUNdq3ty8ydVt0eJmkDeUeC70GworplOH3LfRtmxiuszy7Wp
QlhZE3wRKVrejfn5oRVw5OQpwFnRjmH6+lQnYhx0d1s6pj5Mx4iySoIprJTnMyDLstmCVqPrv1z/
mLveNdQu6FtOyZY7wzGV7KE/IFDljl38TTn/4cGDAOq1ba9XujvOSrmHYbbTt994cA6kRwd/2xo+
nq1ZpxhFn4F1L6TOR6auy6Cs8zLpDIyF+k99gSoXGdx/4VPEDyJab5NJd2jfGaiA3lHeWT0uRuKt
UtbH3j7FzFg5BuvSfKpc2H7Ff/kLjufizxRgk8zMIHB8uJBPH5ip0aTfgTNtxNvaKXL5fTrPOO0P
sEZfdtIhpEYZLxrpNnLfbQqllnPacTbn2C2E+PabnPIgWRG9+IJsB1jxu1QQGNY6lkc6ra8YWMBY
mwzHhFRpD6AzEgJDW4irQBXSVYWj/dkj2h1yqnlWAoyL362Ur64t+nU2Sz4WD5lfFtUHLL2jq61L
0NGW9uo0S5ebD0Kttd7ZGPuT2gZ5A48T4k0oOd3WlrRuEzVrxEpwdCIcdd8Scn3JLsqlf6cpCmoV
wttIiVMcW1Suh4uf7gi1OL6158+gta7I5UihX+tQJrDJRc7ij0YVHJjeZ5c4iQoHnV9GDBMOC+O1
BuJldAbJ+J4gYkrjjV1bRs0+n2/D/+fV+8VbaMP5rtSVzfPUs1wAWG9K+sl89Cj+a3CLXQqeOEgh
Z3R2TNBF42ly3VkfGxte5DGzFaDHyCtXAxf6zPwdwyK3eAYjlzJdKmAC/oG4lKSuuQT0shAaXXuD
DcUhfnou1M0kh0vhiwATGKzObUkqPVnu4xRXUQ0sCkLbb2GXHjtoY6mfa5HsdTu1QIPzh3ZDhUjF
Ay8S990ha2sAdv/bb+TpPQ77hZTMda6C12aABAz6EvSF0y/cmcrRsTrd8wwTgE9C0j23E4ncBoXn
o33BYbsMHTgv5lFzduk9iEWv/RiZ3syuBOuAnDvQ4kz5+qLShHzaTaZFFxMsJEmMuTlV7VyqWu25
WepQ3nyr1V3X7wwzLKLCmt92yvnqL67I7+2D1h2pSqWySv4aHOi3xvLuyK8g0WpzSAFg9pOCGYMO
pe6SOR+0snJQd/GHkJuq5Qad6rlOM6Fn+Rs6VgOdMtgP7gCb1R7yLPpeK0YhE+ASwrDA76nHUpFb
8PSa80lJsQdTNPKGgTYuE8pOVe9P1sK2tiFlsvIMVasyevyNiQhkSwtx+b5icReuvYOCbHAjMuUq
gyrW4ziI0cSxbK9jHunCWq2cgpcaIXhi4VYDLb/746kaHPr8LVZqrRgMXiBJQuYUW7KJHZqSdLLB
kW2/CdqlkyX3PRIIJ1kZw6R9oIw/llU5GZAKZd6TrRmX/pMOjfEPgxaLYtUD08v+K3hDrIwcMFL7
YDDuIQ04VsHCLVaKYrqFzdlLRF8jwYZg+e6OLcgLViKAZ4372qwsPFdRI6SiVLqsLUFXyMjSKIhx
jmXivRvTikelamBmUJG4LyCHizZCtE1O68nzjX46mGvYv2hGQWsWDhBBuQcHh8mxWRowvil4Obqr
jsFixJl5+6CC/YPp6J8QkCSwYBc2nHJHVHAwIJobChatKYtkq1OT6TBm+t+JiRT+23FhhEtX4EQI
3zkyQrJwVXdKJrsoiLjt25Uu1MVK34yXMM+kenTgAjd3wqxHhoS38DrFw33w1VlDC6IZ5qu46wdj
AC98BFYWIZse4opAegpU4jW7xkjTgnmy0tq4q+gKsvv0S2gqNXpr84+IHkt/eJYJ1jobTSVhHgY0
vqD77uZ81q981vzk0lnKYxqw6dLx7tBHe/FzPYJ8XpRw2tRweuwBRAVvvHDIWHuuc+mM9v3N99zk
vlk0pODCPTaeco5ksHy2Vq+PDYgM7bOj8FlF2M7YROyz62xCMmI+WUoEqDAXxy0cWbvNtX7b2AUF
bThz3V06HTeJV0bIjZMZ1AaTAoxHSj4I/G6/hIJ/O4vGa6rH1h+0uAGE9wskQ2roEkVeOh9wZLuq
SwHbqW2SUGnEGMbiA2/635plZopcuAGtw4OFVI711I8s60fgeVIuPgVAV5N4QPJje3uVmtsmLyi/
5SEikANwwuftMcKNyPhCVwylXSxDUdQYXYXRH+N0WGiBQd3o6fdqSL+gTUjDTCCyQX/KFkQ2RGyh
mvMxl/hbpHYGpxCCpN7F2pr1JwepyPzZUkl48erU33pWbxX5piTNJaEqj4o+T+NSAIsnKBP0o6dN
gBRAWZTz42887rjJnfUkT4L6idPFwNzjxB5VRsmDxMO9lluep9r5jhyP0yQykpIjzZAr6/s0Yho8
uaMAa7Q/xwQyBagz94Lwicx/isR4Q7uqLPIW9KYb3PUp9QRwzdquCKgzirNYYNpsc+YRXNacN6yq
4+0XmeOPpqr8gwK5W1qO5hqa826usfZemM429u6BwXR8oyiY87u88/GplNgj29m+eUM0//f+sedY
si3zIvLvRx3bvMyYxQ2EerfXmZES1eq1iK2CO1ePZr0hUu1vq+1oFZpLSBbK4b4Kv+tjTyO0c6if
4pMve/z4LyJ+4PkQEEEy8XMlBGStzMwBzlFdLJmaRelQdULz8iuGcrawMLcNIxltiuSCuk/Gc/JJ
o60IYppTg68eOZ9vj1xFDfC2c53jTnMti7835DllK3hiMzAzxSWIfA4k4CAtHq7xqJa+ZU6TGy8R
QPOXgMG3p+IdxEJ+2ZhqvNuIrQwohizOdZvd8P9WYyqocDmDshSLsOAqurw+1wZpBbVEzVeI67rz
5N1geZE/2iJm4XfDipBwNEWSm+tE4JxpOe4tpQH4pNP3VWk9Qnoa0dPERtVsjxS6EEMTKWklnS8l
4zkr8q3FtG/QkvRc/SDvxgVYqrlq+YU3DVz0uQRSH1iTCJY5IGpQy0QhwxvMUsfUYCZ14sCyt5Io
gxO22IGq6Q7SFKoZnUK+GiNZyjiARYRzJWmqwiaQr9CUmoH4TM+kdG6sOTQglIZR+q4pkCoRHrZx
mJo8wK7bP7vwehihwHiVi4AiB64CPFmCGw5IwvQWUB0W+yFiF/7t0F9T5nIFikVsNo/cKPlrRONU
AAYmwmW8LS4Ba+FPExBefAFU2FekErySTmZwsTvi0AFtboqJfAI6UcLQceCXD6Q4bI754Wncp2cn
bplxY6NMoYuIQLnQemNjJ9cV1Cnp1TGK3/6cRQYb8RIR8cVpSmrlCUscjxjPVFnWDpNDnWAW8U8v
rdTTcvMek6MjhAl9mm65JpcSTnh7r8nzE1t1JN4h0j5pZTatdfqc0qbmTRZgTNg9rr6Yn16FiUFH
mKuLqm+Y2PURK3PQHLaIDJPVNiO1XBQGoU/JvzQ3dZIcq5oyHw2nRj4/PiFblGrkE6+m9N+44ouB
tTbZEaqn47vORs6+JxjnbRX1v3/CcxtmbWYrAU52aun5Sb0MlbHbAYuyXhnN2HX7QGLiT5bvLLMX
hkBhCwyQDeMmfWwZZeUZvQBxsK1PCNO9cQ1ngXG1iNA3SHn6owBBjoMA4BjGE8MlJwfP1mWX8OXi
owzux3uXEjp2ISPEiwa3TcSizQruHcgYwOOwHRzdnMh8opI9MD6t7q8pYJKQCHeo2YbxNZtTdyNZ
wv9HIS7acXfqYB/W2egWhszLbJFi7ihB6/XADg87/zyHCs+0uXcBg0GJujpNcGgsp91p1OBvJVo0
lCkq5YeS91SpTvZZuqZm4yr24OucAoMI+2nM6ZSs4gLv9+SGm6cgLbToszb5TPzz1IDIR6As8Ha/
z8nbA2CZTglZmTbt1Y1dbjUYzpOXTlBnEmhGAsXrP+9t77A3EH6ZU7rrbmFnOKA5SNodKBjNeBdA
bYtTiVMJQhLV5ajkh4/FVKQzYZKGqjgm4ekZpfgpLay2qEgxm4iVOwR7Z6oArsVIPd8I9ATWVTmB
zVVuei3cqHDXf+M8HwFgOYFEslvRznMYYXUIr3pK6+KrvoZrsos+AVMidLsQrAmhg5NaBZQgkE6K
bvCWNdb6JmSOYa82kEMcpJb7KMs4TU+s2pJgqLCJXVx0ZSU1lE1vsr2bAAW5RvSONTXKvznMY3Ye
ac6qedgH1hyANjJlNyfHvNn1iSG6Ululem5gkmHRCEX5cAiqXzoKp8Tm+ThbKEo94K89jdBxuer+
8M3ERnrEU/Np6Qiq0lrY1V+4qyIkqGg9xdgxJf3HT4b+z8Hqpaams3E1FsSXlxUEJVyqwY1sf7VV
UdCk5iqAAco900uxcTASrN1nbk/frMofmolGM249nzTjyk8o35y+xIGIbm2ShtXf+Qoa2LBYG+2T
6vhE/r+NapHNVDRc4Ce0B08sRdd6zauY1DYDN91vwkt87QAuaNfiwOMC3ehgACj3vp+w3Dopddv/
RNmEHG3OIY/k5tmCH6Bl/4E9P2hlstXmegjoTme33vM1w3wwurFVREKGbglPwWyUxmOs4Qs2q+z1
YeV0UCDPatle47ChWbWlC/ndkOaKUdAy6KEt4XQ4ge6MPzulxDoWUnXyl2uXLNYKvxxXoedbuAtS
SJom4A3ZN2NVQzBB20y/o/XGPA909KjDUeBUM+9rGVo/fEEAaVe/LYkU6NLgpb5yQtyDR0i+LRrM
aPeyWQ4EoR/UKWPfHpQQ8eTSDkQqOxdC4GQwVsGLwYEUSrNwMALL2DbmnhNd6vZsTK6nAmfcJChs
wOKfy5OCyeQQa0BJXCvMvZXzcby27uKyTFS4i8IrV7wuUqOPQP3fQecoJXbhCHknXeyTwWYJFVwf
ksC+hrtbzxo3rez3IJTZ2QkbY9y/cuzG1CYcitF2zPc1cXCNV8NWQk3sHx8dcgHiHvZsP7h1U3de
/KZ2d5gTPPvn7vmji1HWGQjDTi/kbzi9gX5LFLJSPsj52NdM93y6JvT4jGXyZgd/fHZFF66+l7ay
6sQXpqVzAmK/8122dKJDFTnEtOva7m/MCc/uR7IwKXFw4fsOME+d2OSlADtZECV1biQhWhLYLusC
9ICbEIiXRVN3Erk8+GVWtfBsGFD4AuOrdnWIhco61e5zSz77v9gSRyG7bj17hKpeRtzr0zx9I2qf
Pn4ybcBTl3sPvrMASgMdpfwni579P8ax/NWmXigx1Gd2bgn4nWIT6OdObH0IGtyBd5wBpN8RKcYK
H0N9OXrJbOYw41elmW+F3vmQ1/xPghutw74/jArUlnwyxdcYNm1Q52lM+KxsjwLuYVneTIApF6NN
OazkRgfE3HCB+gBtA+i4tU8pKLIjNP+JuJShUZ8aB8i67KkjR8leXqDlFuWgKIzW7QP7mYNM6aka
u0x0q6iwNNPlgRqvXtBiZ6ahHUfpOiR/DNbliFlMvfjIpjcKuarH2fLSq68Fge7NffNHzdsV7175
h5oXmWiEQv0dxCI7U0u45SVa803qp+kP891igcEOgRUtfCWjf65Z8W5WTdU/KdwcIekUNBpDECV6
atNI4YQESRtM4uxMNWCrVcnalJAqs06kb2ixiuuhrskm/u8L2OsGRkyJIEG+Lb50mcChbNpZ8iK8
flSgfoHJzDESmNbqgfKGOP1nNndbm5W5/JgK/w7SodhUXjD+NKST887iW8ZXuRyVUqpYMUNx9Z8H
iybzEc7dR+xp4x0QuBAZ+G9ym3o/n5UPxvE1nmccl0OtVAhTV40KW2aWUhw3k7WK/B10sB8r8F96
EMcN7emFVN200bWHAik6EUPJi2IYTV+O4IAkOROdZl7aeYWpzgTfqC9jNDmBRSiazBrGe+IsRP7Y
4IkX/wh22PEuBsxADKORWCp3s7bGMSvIvhmeaOHrzda0l3fomMitcmFNCUqw8RDO/7u5RUnPEn4X
AprdsOuOc94IKmChFSf5Pbo6D0SLBRkufU/no5dx6Yc29/yPeGJyjrcdPrCAymCgEREAIHx4QRZa
RrtF1O8CD+8oiEwPRjzh1mwST58mIH+QJ40gY1KX63h9meLpq8XogkOwyFPiC8Eskufc+xIV2N4R
xJATmoTqSo8N2fhnduPcdyWlOBMfXhR0NEffNFvqlvgEFR4iJ89x+2Z57zYnFjurIutBcJYb9jJM
uCU+mRPktVmBFhUpFrn5M4JA7/6Zx0eZhwYbET/ZrLbxpWN2D4sa1t9uqB2bD0/3ZYWei4MUEWzf
NUYw7BqgZB4zPMcxlljZNkSVaCLDZh1ZcXiCbu49Usvr7LXo17bCWMs9DX6pAjv41WNDd4Ka5cDD
QxdZldQ7q7fmxxTZfg74XSlvFsMcMTdzRd+YurTMKSfQogiV6jMCoTDLFBuvSby8gvgEqIy5xP6L
r7jiTcH5yY8WnUbPf7+REus5mKCGVwZpnK1b74ML3hGU8BnjWhfty2OoLJJOsYTwV9lSM9ss47CM
KPhhzEOPw0SJntS8L/nex3oJcwNmqCDPUwwPjn6dMJIJg4oXRJMZHNubZN7gHJhYlOPO4u3JV5Lk
Y6zmJzj8fK0lbhLeck1Qy9fITGZc7FibQTqeCYy9oJSGth4IQPbdlmLKQmvZ585XSe/tR2c5MQd+
UOevx9DJGP7lbyXajC5DHKXXq8T2u3jQPlKiNPsj58Fv1Ucp3xw4LAiu6o31JW3rn6weNTdKEmDT
ACb2oOtDqheSuscFXiUC+ClPTtSPki6mHzr49w1WRulIxsiQlVaNfXmRd32hjIWHnfvTAoFCyvyl
MKSL8E7BpNcFzLTwKzl+1PtXrOKhBg5zCkqmwrHVlqbnajf8rdXGYLgEmXui83NYTzIBWnGpiBJm
RUqNDiM64S+0Rwll5eU+yneQBv6evGwKzEzGebWBYqAdYepRbndTGqBzjjr5/b11Kk9ChVJDiM49
jc6HYP6cdMEsrcamNLLlEeop4voZ8rIRP5lR2nD/ojF/j2RXK+Go74UM8WjkazBaPsVCJAFM6sw6
TA11DgKsAmuNOvv7AMqxicxUUzVmgAS7YXFq/yW8Kl0FDPaCgQuTpoDM25VpyauinGR6RcAA8Hhs
W0Tljg2uzhyrLPkdlzrcRn2GQD4wfQRjYb3kJNgw4LA2raalxsNv/wRHrMLI5041xCq3+lBKUqsM
Z7XrV7SIbgradkxrU0znzoUj0HmVIoAVyP+7/UC64cEPgCLVGCAu/k4ueKz8MsDmy/3IpSgcC/O3
kr1ib+MsHch8xoi/SduIfYWo21f+sqaiZX8qqoJn7ueoJSgoryv8Z2kHNWE/LfoEY7a3MUqOVqkO
CDUtYiDuDwNIY5Hz+a1XO2dEX/anFkWsOm6bdXDkvEpoAqtEAHDnbe362autvGGZQkWQBveMVwPU
lpsUnlXQE9ZvSszF5Qyb6Xw+bw5zhK0Iph0rd+L7ezwPQpoLTcr4fFn7n4kKGw9Y2210vM9azL+B
dyZts/Z8JWbhAh+kHGxx75mKXfpMsC6+mtb0T6SMmBSK2jhRwpELVd5GqfSxdaDbQcYJfT+Kevre
CdYp1b/xYO88Gi5rbbeXkXUfy256bI53sqp4kJi2hM0kqIOR51dn37/TTzPSRHhIco9TZy04sKQK
i7Fpq2MyzwVMWEemNHIzO0vGwVh+q9v8rdR08wpTvZuK/dyog8ns9ziXdyeS3HGA8v/TrQr5p7GG
swtKOnPtEGwAp96EmjKfoaaWg/msCvXwBxWcX25ULrEcH8F/QL/GOuHqdUkoCVAyJ9yhkO0ovud5
6hLW+9prkxRupo19XPLHW8gze6eOo7/JA+iUCNhVVXT5vIyqe+i7B97HF4u2Qys+bEDIUXGpe7q8
GUT7kK2ZhsYYzgGF7jSGa4js2DvgwG8M2Lgub7Cbe1p4cer6bIbqi+g3A9uCJ3KAysx5NUqPy4dP
N/ZqOd/1yYM+b5tO2aIKQUu638b1nAXXpJTB3TEDD4gZ+Ul75qSE5IarilZeUOUZUip9f5eeHFR2
C0czX4fGymoZvPBU4eY3QY4hp0V12w3O/Uhu72VJG8/HYGpjnjeKUGINhoFp3emlPbQjnFUGw/DV
vxIIylT4Vw2NjmvMTBs70Vx3GYkOCJUwk2ymXQP0lgcww2aewvWUDcPLpfm6vHybR3P0O1L01PsV
Fw57hDaI9XYOit5PKp5lVwEHye3NSHY6hmnLAtlGUYxVbV9+n8fCe8y/ago+Qyi7c8VbnLIpS1bw
tGp1i/1eGkhi2uCs0UhpahcPcf+40yzq9d6x1JyhBWhC4PwMWYd99FDGNEx6sb4hAxbLzygl8ZY/
YuNw3RNbONoH764cn623clh6h92jMLHyyRSb7Q5WLI51bHt98Zj3gbsYvrvTD5TakjAHC8VSIELo
xJM1ZeWN3VCRA5pP42ldbTQJ6/ZrQNlKTTbelGzcB7WP3XPf5FD2+RWEQV97mPLT0GTKoY3jVAv3
XrHW4sTXOKwunUoc6LE93GYXx43Odew2M20gVUpHYgJS4/T3Yk83q10oALTTcW3sWU7tc54PxgRr
etaKJy74GWFk/ZHZlRT/H0TLO2nm9edomJ/o6F7W3EWoA1mmSeEjjVpgXmeNONphJHD+7QaRLdkI
EFRhngxDwHuUq8X7BaEmr347FxMVoRbtL0uc1pvyMpJMiQwKSMnzmLDOR2GaODVDDQ+Hfg1Zzf8G
5pFAnWKEMnfnhUbnlQtxcdknXevafU6QD8mqM/AEPqJEjZL61MyLb4YRMR3j31StfogbolUCEu2p
XUsovoDD1Ew8+VyFy1noGn1o2CCgUeAW7zNItAkXcQ1STplSeeyPLx3UHFq2VNtLhqiTc3pGYh7O
y3RIFetbkVzDDREBeW+YCf/A9FYEm35F72z/YKJDq4nU6Nlgr3ddEJ0XknIYayAEWDDhFMAAJMl5
a86llfE9RbOEESGJU6J92UxTFIW+beazlYPkhnH09q76FExVezwJtYqgkj0EKroUJMfabaqfmG9q
Jx6FLSlNOqtLFLe6PLYZH8mkxbXF1izHC1QOGoNbA4JiCeS+TgtRJi907cEqJV12ZazCo9tw7jY6
fnFzUxO4B08JbVCQMCt17nX2j4LjsWy5/V4g1c+zCMGW59oAVw6mwmktWVaJivoZSNo0e1+CW0IQ
4IGb5x4v4IRHUHBKmSUFYFSbLfYei5pSzxIvuq7+IqMhKrWJxxKDhKo7YYQYtJaAznYiOM66oXe7
n2ZpBASRlCIs6kIWyWZXRfHWUiWmahBINO0FlW2XkOt8VhxKmbT3CpDDwukYdZoBscm96BNXour3
LrrT9/DGgHl0ENr9lgRFPARQ98aN2uc9FemKhSYxcCwqnd/x3f+N+lj/aintuqHLN+ZUOAikpN+l
vMWcJ88b7YMRjJ12pBiUMlv/vpFdZBwfBr7ZNlk06/4YLFt7r2l/aqCef2DAlpAqUIRE7KmeA77o
aRq3JKzoiZSkM9eQPz9FQaSK1jwCYESILq//fpm6fGPrchl5Ec88tIU2BdxaphaqSiucBlPshKcb
dBh0LPsDAOn1lIiFVAVWYDAOuXwulyoLBdtWuBFwa7XMcE3elINPzoRosv/N9v/FZHkLMgg741ge
PLlaknMevwPbWTmMgAjnDkGTrkFiJl+M7oi+U0rNwGBprpK57yWapVTjZpAFpbUHrb/IocHBfZBH
bRQ71GhbP+KLRKnO8IzTDTSbRR0ECk1/qB4OG+XKgvSVtGcAxge/LlEia1gJ99a+5O53VUyhM3UM
QjW1ARGy9fAuRvnbMDraDs3gOkHVjVdwv5l6DIz3CW8ZmBV1aASInNtyXt+ypfLTlvUQmdAH7AQU
+6qVJFxkkeHyw2Zn73Odao1SisBN1C4qGm7FGr1L2WaksUPNQOB+A3uI2yfVp7o8BZ6FMYY59I/n
JF/YH61XETdIrw41JXiiEmn09+Ay7FdLPpcnrnWdJ6e+VCrOoxIYlWZ5q29iXYzKG3QdBspUxAhx
Vpzo9nsoQPhH11UmbvlxHs3/VevrRveLQUu2gyffen1nJ3d82rjoRCeL7bmQiqUBOzzN9VUKXX6a
Mf4Ctq5+1RyKHKUv/RxM1QyfGs10H7uWh9eOVhIhdXkOMV+skeDP3X/N83BVOsleV7Rmsp9wE3aL
GupHLgNoWJtgm3iagaJA+Vt8Mg94cuHjCOsN+lAuS50Vj5qJQzpKls0Epbgib/Yu+t5dtWz14bg3
5nejUCJQNt/czmtM1f6JSdnmxq3Owwm0KU+bb+oRGn8MiKdgFqbpe0odYS4VqJAqmJK9LcsyTssu
p6sfNCIc8Gy8vUcJ5+LDGjuQBlXkHB9Aa/+LxAb/+ivL44eg4XLbthzAQ1VqfX8eP1apT+lC8J+v
xC5QElPufz4LmSAcg9fkUkjjFy6xMXQWbG0bKGJIOpvkdlJwpKkANGQ/Q0zeU6rd10RKwZqN6YKu
jpcGT9Fc0/seOv50t9ArEaWpvYEh3IYEwB0mn/JicfiqqDBh/vraRWv8QatYdVUPFZLOOg3cnW3V
phGV/LMc9ab3JMHqGzBiqGJt4s1QdgN6DS8VyxZy8jW4sMMA4M2QF+x5ZF99ZVVLFrVxjRxaIJAO
ufpH99E4y7pc0Nuw3mMkerpOQwllZaepQAeuLABvwVLCQnbhWNGpgu4QNyKyRJlR80T31boy6jL1
033xFxza+lJzRvbSH6/xKeY029T7l477o/7nBwJFp9vSCPcX3Tdd0rHOmA6w76Is7EPTgrm7eIBU
wEMgqDDnIjBhQH/QR5EZQFr4iCUmLVlmEVhKAh9H+dHSdnb/hpeEcBvB9YHtz91dLmllyQ6RmSeW
Qg44BoXIi97ax6ZzNBy/dCwEQb6D1ZJr7NYaAwB2kNEm4g/JlEBZsjIx+1q9TmIoaOgeVlAQemka
F9Y71jt7XsxRbzUI8nWHqXykXXNug9sSdPpn4/IpMNQLeYY6ds21ng/QeHizseY2UGUVXl3RbOSL
bPK0TzXFNqaXFqVVlBbbnyFANQ1mNab90NfSMoYZlLAeYxQ43QXJ0E5rI3LXGVEydw9Xa3GJrXxz
wTYMT7ds23BRz274rXq1JJl6hktGgaXLQKDnp6RexGnfdSOJHy4nFc3dyyvUmMM9L3v+UY1juQ5M
40YFCt+Mb1eENKMbit2+WHeGZt2d21MPnika5/Sl+potXAQviDPhRnNtf6QHs1AusFX55yfXFj2l
vSNJAoM4SzcNWCgqJrvxm8Ddj4cAH2AkzmXQ+3z8tuU5CFFYLbtPRPK1A+Vh/zMSsz5oajrY6yoF
avfl2TbkcUH4OMRhYDYE10g2NP7c77O8QwDpt5M55eNxfpN1kA/lTCGrflXYuQtc2bbmAQfurFhF
i/mcKrxXK5gJE44wJEwtCJcSta08diewdcsu6YQyMd0MWwNOd0MMEhXDiaGa70CXy4+gf5FXx7De
hUNQcyWJ43ttduZMzEToXKKHRT+wxN9duu6AHfZPUYiqM9wii1qYwHL05vdH30ziiUY9iNDcIr3e
8kcjA3HMP0sVVhNA9EaTjJ0Lb94hzKe/G/zUvn85m0cgP6cnb21UwimPyiYLiyCsGGr2xLxAZe+o
Na8ea+Z8DRzDMs/Xlz3JtwDAFVqv3FiCTUCG9rKmLr/iOBzO9Yj/0rUfh9x6WgAgEonR9cMpsVKD
bEcDPczcs0SNRnyxoHhqPsYFzqhQX1dz6bnElT3NdjKaTjp/YOI5xP6dMcKL7TmnIjBD+wT1fsCG
qYmSIDXF1UttmW9cws5+rnQ2CTGyoPB9Yp6MtVheHFEzpeNCo0U/M+c6b7vcTeHhUbl3N6ccu5up
J+qBj7IkGkuU+72fUknTcU38gNCX0JhA5VEL+Gzssj0uAu2536or8OFBcj+GYYwLPWn0d2fNG3Xm
2KsRlY6LtTqatTqzoDYrnBKB4FhEjrUK5eOhakjLBuGv3zs9SmUcNsVzNyiMX/zhma2hQdKayyuP
R6sFWOruLWMWChMoyYMgkiMKxHZk09f1GSphmiMnyJT90gYiYjd7eLzuVutF7UU9VyPkmmNoc0wO
dgz+DqGlZjNi+Q2Z8UH3kUzx0UirbGYuqYkuyi3TprF4Zdc4hOkCp1koWXmTutFIG38xJ7ClRxKl
FmJ1OLpESnIGXzK41codXIh0HZCdNo63HUPRgodqCo4LTz3V4TdLqvV7g499RUn8NQmwRTz69ZE0
CDHs+fcm44S1+l7vXQnWwwRgyCIheb8njVrhHpRQ9wDjceqYS1A/IDnZg4n0vVAOnywt7vhPyWoJ
S3f6dbKeesSmXVfnrvjVE4G0C+hqmZtJeoq5BFDViDKP8DeEZWlos0w1pxJxCzLyM0+cdME/4Ss6
/BPwZE/Eu290HvPIzndH95HMoPwVWrW2/5DQAARX+ZafC9DpCbhFhOzebDUjwNYub7gCBr8USK4s
Ne4Gq33QQJoqb5u05Oyo/gech6pAV+9HA4JX4O+tVLfiGBhHvdB2v8n5JGGFyhopIff02Mi3zfyA
pJ55SrJ3Kj7Lfn4XgPWzjdhAVprmMIcTciMgSEiOY1seRxVkaNO9AFiVUi3jGeGFsZFXLd/2+liu
sPZHQdyEqaQ27CX3n5wyddAOzz5WcBMvdAoRGXT3fUs3QObW43Ma9tfL9s6EwVDZIlkdzR0ZfZz7
8d+95tln3EWkW0ezsl138XacWrXVnleluq4RO/ZM0RFg07XeE2ub8/sJoqfJvPrKltc1sVpqcXKl
/o7/+lD4/icjoMrT6JWj89U37LqyH5Sclps6YCZ2JaApSCfPan01BPypwGaSAf7EOiqYRJgtMHHo
TkcqyfmvVmaTfIkq17BTM/Wo+djlmS42r7DhdtSnkbl+O6OrTLEpmXacJVYCvj3LpN4VqTVHg+BB
ntnP7saCxg531Aw5aeqBHLIM2ydpgFO9EKDtnCbm5kuFsRzn3bUvLdfMJqGD6F6bUmfuNmwfM+9F
u0UQDQgzx9VvK+UbHML1u2UMR0LT+Slb+AHO99I62AdJ3Nfu0IMENCl68VLbILua52Y5H1TzRbpj
Zg2fowr1ZZPpakF3cYNlKIDRupcprI1JcJcP8bSdoOrka5YD09i180rITBe/QC3h65tDZReCn+A4
UtyO+rBSqmAL+lq2hwFUB1O9h1gYVlwayMt7Xnb83QuAblXW7X+57CFhnbuIE9sleb0gqjmE1ugD
pLOpfOfzGFLPC/FcrWUHwb5ySYbzWSH6CllOIBeGlZ5MTn3E9fyuDWPck1il0gLxk/RMANnGRhLU
TmR4WzTliQLo5Epfojs+1MA6STTk8npj+aO13puHzcVMR5hvb9vGUoJEYYtKbViVWL6m1Edwe/xu
+3jqAt0SFXr3w/WsFlMJYqwCeZ+86goUXLAK839OJ5UTIK83p9U1tPKmqr46htv4R32ZdYZjdKJT
Q3Wf4mlsep00pKd0cVI6cirI7JYOvMEJss/+gZQJhZ5uM0oGqSVkVqqlp4D1LxFGjqO4t9P326sA
dNQCujaHVQo8EBwzgCH9wJbSYWwZT1NBSOaayW4mJuw4PRN6BGgAzhoIHL340O7EtdXFaUeI94VT
9esYb+uO8CehH/5hMtMLAu2AHPg+7ueR49rlI29UOYUZqVS504ya2S4NbiDEsnhE9a0xUQ4fwJpa
PJjmVewJ8xxLZWlvETaMUvip1FktOq0/u4gl96voGtSgMVsCNAX+m6VxXpQxX6/zNcqy7T2rH4hA
PIX/g/s9p8XM3qx7Um8gr3FdzWvrNITmOIos4+9K7IvpmXl/Ul/nNloqpQi+lsXNX+TMuGqSw7TJ
E/DejXKKJvXSkzHs4p1Pfj0ZEXTaorVWoYoo7VGMVZ5IzVU3RAhsO0oO5VmV45HraTL+WN2PRLO5
s6TunVt4GZ9V8jayI3KRJADiQJnu/SeRYBnxfw/J9UGVL1VVHbsoPHEg2PKQkdfVx5uze+BIFAB6
D/j2S5xGTZUbmZmNZrPew5OcQ25olnKGfNH1duP41f8lHxWbqRV0C0LURGJfYx2sw4SvjmpD4FNs
Mq4qPkt83D+wmTwOvycBCHILkz0FT00FCUkSwS3CNB375qyjQx3Aoh11i5LusPpRwQC5uc4gTPue
4eUbT/xlt91VStcUoNXesS2KChhGLOXNfKlUO/TSJjM9qs0Yu1tRzWFhqIR2S2497rZu8i3CA0Pz
PfQRCVOojdCSCiCUqt6N1UZXXEdwdRdADVvjiXme7Fwl5/Oam2n8SYyJOYhJrXn1gQyu/2ybm+Le
WRq8xEMAkZ3LOe3pASgQlWS6c7esKRvYDBGpV4M0gm1GM0AGNxrwfBX12b/BsnUU94PA0wSTU8UI
hKZESFaSlw7JFDMrnrPq6gP1M88UTsSxvTmHuqg45mZbsJX6e/fHCR36Ej3yy3Dqv4Y2TOJH8eJI
A9fiYLat+MUWc5EPRK+t9YD1b27xuTD8J/l1bcswB3/CELpsajdthoXZdkLX7R5Gv0x6s1g9h2uR
5HgeykXOHRYNcDRJW0UunaVTVo0ButQPKFp8TAcltvH+5jdnHP6i8uedbxPXci13uPqKL/2blqAR
SYa7NyRf1by1ws+p7rxdjcobHbokq0xE4XBo2w660j63beArX5gZREJyhvUIbWlDRWBHbeXHreI0
vd7PWEbVb4VXBgaRANvgXHNzPL+8uQtJSWDzReQs1ySAK1R3ethM/aIJ+KDeiYFu9fEdY2xt72cW
oPq2nQj3zyHERyjVhQmuq8Hk8uA24PgNReoQlxUm3x5djI2JZ/p5/3d/yg4aV8NELM/JYC8pFrYw
gN9XJE4/JSEi9hy0895C1l7WmiCv8EPnqxLrVJlLE8gPZwlNcBWv/qO4/Q9Pw5vaAQux60YYuMbk
rds6RF/LHr+ReJh5ph7LYWOxlNX1E5VEWhhsM6524P1wuDWEYJiZljRZzWNs10eiUgl/oM847V6W
jfrkqu+42fn2lJFmpfjobFRayMpGngDMLIrbBuZUoSMhxKpHpCr1hH7bGk8c8UmVOvY879+EDymE
exTTPiH+kvyf3v9q/+6nC7ZXACU2LzQ06nsSfjYfbvKdDmER9Jmzwj6ycbmL312J/RKgAPH1aWY3
LoWPv70CpAfrOxVyMgK/hoTGo5Drb0Kyyt8lZLOOhznLWZxSq9gI9wBN6xpyMwcGgnmBZlgUBimq
xy/Ygm3/vUPPY00oLGMrwIZ0rEcW8xxisXp2KRqhk910y+6oFOLw7YJi0iXzdyhSn3zx3XdpZlxf
1Z+SSoZRkm8BeilWih9n6Rw1sjVZGZLJY2mLbaTIOWpZwFGm/KYPkrHBgYe06A7kA8OBS4HJJdac
jG0szhzIkcCS7+1QQKaEp1U6k2sTxyVaa69wfnOUcQT82OEYiMLgMCjz9tXzX2ib4WPM5h5B30Ue
YR94+dCRm2tGAWsbl9MQP7YoF5evhkc53Ea66LB+U52P+gD5Z4GXv0kG88o2ZYhd6JIGqZy5mebO
xJ3g0+MrX3W+wGWffhcLlss/7IMcaYVzuc+nKe/k3wfNhdnU80sikBZttuxdXZW+IrB4ZGRdZzNe
YJF4pUMKD9a0oeuunGuiAvmRheQSpO+InoxE6S8ZXBT/JnoZ5Fm5h/x0Lo0auC+xoPCGLvI2/0fo
BfNR3ht9jfTq1+WHfciLmLrgM3TwqSo2Uq85mMgw1bInLXu5L7xeNPHVUz6I2J7Dn1DqU6h+w1K4
nty1YjyQLRxwWak5TeNW+MGsAD1OWYczBvFotmtI0mAShRT03qnN4qFdtaqu4EQg1kKMC586fLXX
wl3uJPfecIQtvOb8zKLZTO5X0AxKu9V30bgmV4ZGvnjaXzkZk72vGKRogabcSCW2Z2q42vWtW4mi
caIvF9q1+0O7JKmbEPsciZ0Do7+tnPZ2vYyrqu/TivxqA/I/CSH+K03Plp7efxgDtbKyBgQ4tywx
gfIw4swoOUDq7Z3+dBLBHTSIOKvx0uH4EaTyjsxRSTPHYu0SeHhbzVB5DC1+jg3qMf3umoF718FZ
XPf1rZ3T0if3FB7x6yo0Cgw4ya8HKxOle8wqLlybkLLRiPN1HWTZEKJ+38tm4SrQqfcVCTtXzL9n
ZGuIDH7FOknMiVXweHKnIPldxCSFCMmmqC1IiTCR7aVX599kE9g5Z8Kvvy080H7E7ekfMJ7XH55a
SHdjbSkrm1Kc6JA+6kME/k5vQa8DsPN20tom62QX7hnMYZDPtKAcujDI4iBtNthGiMxx006mY6PW
B4Sqzc1O/3AR+ocZ2cH9Bm9fDmCtuQ1Onqxe1E8gd/h6QkJWqgvgaoMmdCLye3vtRNFiN3vHThbS
biRwaZj5mKEuoP9KuxFDEZYrJ3JTLL6lv1oivu+QqW0wWwAzeDs4Vd4yJJsqzKP/1ApRYOkUNduA
9WhVlQFStbQsz/r2ltwwyCGapFrPS1//6YXCtmg/A7afFSgOcCMQpNkq5M3lu/Stu0LgK1j1WJ0B
MR6fWp8JQyrRCQP1Vc3iFLftoYM9Zl/gXVVd2kOj9VmXR8bFCq5fxlRhct250s2NTgZ1vAOBUkF5
5oIQzUc/s7ClX2DJuV4N/QtVEJH9BpkRNQy0U4MMuv5+HNlGyKEHoF+Ted4yRuxWkPSD+YWXR20B
pcSA4Q+bR7PTzB0Jh5CVI8UZlnFZ99s3AtfPpXBhGMsyPCQGHK/ZnAeP94khHvt+HPGKom57bcbP
mVnIh9g3pGOUEa79AAdIdao3WjDA45HlpljggNznC2XjcT0mBjYpJki1N8qxBB2+iZXvqHs8q1e5
X4ADXnoqatr59anT5c33fRAtsvsGn2b4YZUYpVswiMkaRmlK4bDKivlTBSKpLBkDW2a2eaPAKac0
SucErnpVmM9u+BgBBw2KOOGr2uUvHVEhh0SbhyzUmRAShgwFbJQ8exsB3SqllfP52aKCzzGVRRs1
YU1tyOOPfSrt2zJuIfh+CRXnVBb5dUJs/AsmwVsYxY2+yXoWp5ErLDEOekbSLrF7YOhyp8IZJU5r
JtYcHQ4N5Az5BQpxrqV/mzLjrbQyU+EGADoZlhtooCvsknVtgigl/mN7ZyCm93v42PA4iCeo7UO9
2AUPyzaa1BmCmaXd6XmLplSHYGLTxDP7gCfsk82gLKcHFf8plrGoC5HrzGecR74P6yTwRNARZT08
IUlpS478TB5zy9yB+/aVH7y9BzYDayUug6igoOSF+poLp1d1mKJDFUl6zSWHVaUmxWgdSb0qITbD
nCQ+VuEwQxJl5qeqsb61yPOVQvkzAqc1q3bhbsvLJjrArXElAV2JfXT1IjAsYew9/3Lfe9ug2AIH
gNFTgE5BLVmC36zT2IAVIzXR9Pn+e7tylQPDVxwdAqNQoAEyUEQ5u3VWS1nWvEvDUw71DnzjgK+D
ei2FpQwX0hWqdYCZa4P3GFFkSQpgc2J4CFYm9Q1SRKficNRGhpDVQ5++VbUcgEROvmeYbJNQ8Xhh
rUTyIspEVMBnRZYtFngcT41zK1Li7KtYGvMGYj1dj3DdBHYKcNYr5WBWr4RvrO9yOJ4reGaO+DuS
oSsa4l+MzK9knyhlX0qaZoh6j9A90DPQfs6Lu512oHBYoDcIi8Qb1+uAubCo32Vom4+OpRCSNniH
ShFa9ioOSI4s2OXmdlXhmFJkpoNb+B3Yoaz6QbS6DLBIpyB8b100Jb+l/U9Hh6KeNn3Q6dz1WPcC
4PQHS4O2yygrx8g7BJR5um9ytiiuonLKOL/p1F3uo/X7c/NDNGU7wfnkQwDFkxXw9qmAIfL1xIAQ
4bTW0j53zgJotGU72ZoA8r7NCCNYhMQz4a0s3ruX1Coms1ABv/9TReJQlZj7+JrnsAHT22Cdwzu2
/zEEpmpjDWTuxzC1J1x0fxS26npcdm9M+fPNCaF52fTtavJ/qyEJ3/A0THojK1dnQwB3w/VwnTb8
wGMvnebfw0fitCmBQVDWSKP+8hVC2myjYohk1VQkRvsMeXgHUVDNCrhMJCawW6VjDfzguWYmGlcC
ufrjt/msPctGApdiWR6T44M85Qs031yPMpKesrdVhMMGbAuBJWPvD52cLDY/GP8iyPUsucb9qnOv
eSNRXEMnVhGRjRJJQUtfvewNHpgy1I/TnsD1ErW2nau44LcykzfvLCDKV6YL9D63VDZ/J4egqbQX
g5+UHeXyw19nwxCE0kI1l5ybr/qjKBXCD93cUwFStVV7w0WyCBBRQSNwh7j+Py0K2yR7eD4NXsEV
1Z90MagS/Md6SANbuBRV0q9a4rqQqkdgK9tzgiyCMu00Siv1DJ8S4CkdicC0OtFM7pgJUxsAioAH
YkkjR1G032mwQ+ZWiLOFzRwkR+o141J83a0WeZtrN7MAAXOl/FuG75bFLNHtI9F4166MBZYQK8Gl
pGtStxsuVGIyzUZF9icbul+NsVNKucxSwI+wMKZWIRIvFcodo1ArpHpR6Ycg49ASguf6O3TR+umJ
jeIb1BPwz+1w7EYA3uR+m7aj6iHWCQKMjIDITrzVb4ptPzkVAo8wIwgFEQ+TLh6zQAPkTTkB/0kq
egWPMRP9xnjppIbkZBwQiFYDzMC8JCjJREbMrZxhKVa71UdUx7jw9icRU6DTMd/KlGXvL6IcFGgO
HqnucVs0TFzSFERNetCisOI5wxpO/5W51qeiTJQwGaxh/Oc7aQylau5nNp98lFVmU/guQx4+Ew0L
qCaImRyMdadzhV9BmDZ7XKzq14UBp6yR+URm2sh77TZf9OEL+GPl21/yb7Wnox71msb06/DDA3wH
LCs8N3x5l7AHAZjnhmtCovYhu/sboJ2ed6TLkESpsfjKMU9x/tEAzD+v7dRBkwfAdgxmbj10GIoK
BBzBZGl3/vd12uR+k08KpjJEqS/9syeZ582j/Uhnh6kUHi7bih3K1ZGEP4J6CgAIhEOENkjjhf+H
l6oT9qQbJdly3CbnB+NjXkUPvFrzWf+QL83mOc5Jmcck2mwWuR3vhhXssmQiRmOfCr0na9E47jnk
X+w9EEtv+f+3YhQbywvWpeGboQVkBFMWKTmKOLvz0DyVnxOULejNEx90TjpQc7s47Iq5Esh/u1l/
BH+Pgcgik2dcJ5v8BZx4bGkjDV/XxsKXpT2efMBD6xibIg/FHp/8NhkokhmeQDJOeofi7GJRa0z7
Z3CV39QPv5b1puuKOTYcOykB7CKpfmCi9cn/+7e/mfiOICAgKS521EFyV7s34w6kTF+1fTLQmMjp
lomugAcsnJW5gf6IgUI6MzEg/lfqgQ7jO/rAHBwiwo/0NLACrB2KN1wmvDEnn1zS8nuEqkL6OOor
CFRIq79wDZ10nMDIPx6cz7fojfyLcbOm0MKD7vId1Dtv1E4fEUHzNIoSHcMGvr4OTnJ9cgioS7/f
RSvOCgZPeNwVSyBfEgmpBcitxXctDvSUI85+B8/UcSzLJcE/B8oNCwAXzfXUUrg9z+aQRJZJnGyq
1V6x7lPrKHLIjOZsT/wdWZD8oAg9GxtY8R1fI634zqiRIQtjZ7+0rk3Mrjwez9tfnQwWkj/ofdV3
7Y/ad7xZUX1NAqDMua3REmggQndl/XCV9dftuxASXDwNFt/xm23/3d3wi6drQBY0s+f+DssBYFFh
C2b4hqPLxm/8yEXLF9FwJjpEm/mJZ8aF/OghE2uT/KCRPoi1gpq1EtI9v4wZPIaldZ/58OAK/ERm
BVeTz4KHUnodNFdq4EnVu2Z9/1/wuj+bQnMyylC5qO6+Gr8v4YAMnIeqEo/Bfa26YeXHRkJnppxF
yGEeIhAnvA/a7IBU05IDNfLkOVOMJs0WoVtCennzW/j8N9raLzVYYyNC7kQwmogCq1+SDPrIZruT
c6cxRFUJmOLX9+BjC0UBCYz6aHxHaMQMbZ6tuEHR7f596oMKYmOkwsv2tOrCe2IDp0+oQRp7muVQ
BVBDEzXzKOTRlKFdcZs5C0qvIFkfPpq9v0m4rlNgPR76PbUBPt7BUIIICOyrGYNAMS11Rsqhns7j
R7I6TWub7qgVlII4e/tQU3CBV9H9wXZnRkYUuz2OzNXUNMVrgc7hISRlCRDyvJS7Xeos9gOB+FmV
nsmuhMOnFZT3Ep8EfEnJl1pAeFsyU3q1GG5AnkXqKOCRvJsxJlHPWUuh7ONQdZaawG3B9tAEh+mv
2iu1CziOWXNpDCk1gzIzRk1IR8mwJRkuNIaAs7nwHo5AGDUKvBgj8HGU7pskz8JWCv8V0oy4R4gh
nMaYzXqkaBL/OUzT4xc0rjyhr5dLwAC1nmJ2uIuAjmVg5JCa/VAuz2CRKVEUBCgczFFu+L4oP/UA
Ia764SO7XiWUentxpyn1VmGSdyYx2gMT5ehxbDU7n7qnjhICSYH/hHxQcHtAZGzgsvzwDa2C8MYa
QJoX7v4A0qpREubQoPO+PV5fWLKB5Cqbno86b6hYeRxAB/MfWtQfZfxMsnOOcJmNrzNbkR4NhM8T
hCg21WJu9mKpfspnjuo70CScsMUzLyKGDXu9vf1RoJng5qkpRHfuJYPOGLtQs8Xrk8/GLFTbFbK1
3pVLUR7fmxgBZ2sSZ5n6PJ0M6rTNEplXF1+qsxXkemo8Hna2NqjxCv5SYXppcsUugJFCs8lEb8D+
xpbWb1I/Qy5sU/mqGPNeWoiFf8Rxzy7NcVD/EzHBbIAlCeNbMG2giD6JAfx4+pA=
`protect end_protected
