--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
h5h6D2j8fWqOH9HzXGIPOw39KKYO7QfH2tjASSg29HcTOTc5WuJzfw018PXdgxyVKNSmk0Ad0dec
6ipwXJejXdWraur5hvzhu1CarMNHqeHbmhdMcusyhGtUVxkvxAUx1WGQOcSnU5ocgeumDqowjRyk
fKv2Wa1S4s3Qhb9aIJcHiq0nUTnIEm1v7Lh6gfchxVnIeygqzd+Do36x7xo34j9LJitA+WszPi41
lRbKZVDmdWOq+QBR6TWf40SalAsXt75bGtnYzo7TUNQxedfv3T3MNCXXX34/pOM0UQe9T0vqHHx3
n2GcRgNpCc9/1sHQB+ijSeiXvyJeIMZZrGx+vA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="IBzWvdDG8bdZPyjLD2RL/ajIHtXPUsBSpRdA85penME="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
njArL20vsi8+W12MNRjqB4NXQgYai22LHVeW9ohM7CZVvR5kKQIHsM1X+hcDEx9TvosDS5kqk/to
zllM9Ah8v5/lb33A184DamD5moVdPXVp1I7ykAeFxCjwBQ7D+X/pqiYNXOMYd1fN+gFqUq7iwpTI
kbSkUC6xX5LeusdyLTZbxNE7h6GmrXo49MkCYItE583M0GxGw0OztGLZRPl8lCjhyxcAzDtRda6t
A5ly1JrdWUFOcxG+Dc5YryGZrxcZx+BDwODXwY+Gwbi3yAUUuXK91LMbqPqu8uSK1gtMVvLkH1zh
U2sylszjxNwmwiLhPQaHhfIpcvqGhNZYsHtxQg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="ERwvSGJTnElQLw432fQy00XaOS5rJjKq3J4YtxrLhLw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19584)
`protect data_block
A5kwv4Nl+Yl9tnR8+37lIDNQhg+CRDd9LW8o4u0PQaWcSOOOyHtsM3DwWeg2EfQeum61vqWOH0Ve
In73nMswD87soJw8Q7sjiDCYEQ5sBXvVqzOfZi/h9QwToRwhrbkYc0Q71TbympxpoKbHe3GX+1fF
yyriJDVwVAvTXs/HYnR4zylW8zqMsdDy4GJeB/EFlYGi9X7sL1F2SOYtLSsX2D68J0WiBOVFMkXn
3ukN7vrdP9FatnE2twmTegHH6lmF3aZY/IAkOB0JuIT4Al7+UWTPPZTsR85jfCkahyQ/bjN7dq96
7Yu9yJUL5kEksABlJZ+HD0apccMV2qWn2GN5FQ/dL3k5fcnfiH6uvcD8R1FaV8xnmYDY7hfrtD93
mt/Y9dS3uAjI7J036Goka9jKgQyIVpcV2r2EX/lay86iordo+xvIqhvBTTe3wCa2OxMVlLPBEkCg
wQrtvYFQulNt2XPWVmBMmJX8G/UdIoCtMKEtXvT6Bot4twwJam7b2QAD+2+AvwJNixtJuKJezscb
wHwYfesT7+2zXTXTGzgdyXy4YmJ4Vw5CkFCBqk7UE7l54dlOOkA5dcddIoYbEgcmv/Le04MQbSEW
FgHTGrUcpnrhqQvexiquyG7olC0lFs+3HHvXkxuwzqE0HJRQQ00yeqFd0zDl1l1LOJQ1rB4t9kiZ
bwOggmIgphB0m0NQkc7YYgz95KSgeZBhE2Pr4GO6RsOmFh1D19U64WMbd12SCb1O17yqxrveMiZr
pWx1Dy5ZnnynxyxS+OqKebFxoshktTfd9BQS1AQmmLTGboiFBOHeZxlUeAGtdAflu99SOLmSw8L6
MLlBcughn8WRoT/Q+LLmp2OmY2eYWIlpUdWgiJ5Ah/YlkxqT0+8v82k7v8srPXbGyY3FZVvsXkta
OJyALboijgnVC9ybUNvM/Uai38o1wX/QAN3AhIuXDoE0ulZK+o9/7fO0sE0613fwdJpqpj7BpNhb
V0ukY4twmQ+v+e1ik/G2EtrhNWtVIfHPcf7TSc7LjqfkzYk/ZM/W/HmhwbPkcIhovWcu7rVmGT4q
VfhMPn9p8le+rxk+ol+I+KJu29WWp6Hjn45hquhr9M7ExDg+ei0D/A9PwUuW43vkBZ3LHgi4Q/pd
hIOsBpfKeb8D2J+CrS+N+q5Jd8vj/AGnnGSXTQtjreLmI+OQX3ocM5JcOe6dkPXvkFeUx6Wwy+zS
NfXpHCeNpLfSIsHGEp5Di+NRsXphDmY0p2MDpVj1LYou2PeNgV6F8+83shFcBjCC/aIv5DHNDYMx
UPvvdd/N7mK5SCN4I01LZ3bXlJyakDdX1dOWfZdmmMMU8Scj1zZZw5VENDinSg84lXjjkizBUBPY
i6Rk4odkd3T2piLVE53PWCQRpXkrXqe1JH1CIx5MwhubNXb9QGukYpoPRA/ies2LaIqmWpx7JTVl
8y0rI5dR9n7WBFEdyflgF/voh1DEZ1paO4brXxBSwW5019k7tMBPaHR5YquI7JMreQQ60WhOt0tC
/AbKEexrFNyiiv4/r/fI5RSsLBNAxfJl0fA8tujoB7rH7liI59vw84aWz0U9lF7utcat9ykOn7AX
97hA1EvYQ5NAuIy5t2HtudDD2X2AaAEH+P7qkbTdsPjzHNNwRKTxcwnDsub3ONGKVR6vxLhbNRRC
/3Ie+M6uA8kKxSbub5X1ASvZsp40BSPBA76YgCa5VnlCGVIIMEBIkx1tqJpF2uVtFxQhNt0o5Phn
rONCpFnfarP+ScxL7HbnRTBBw1nDE6VpQ5wPRGMOX7GBSVvOUro8gjS2kNHCw6FR9v01YalYEMn0
gP/N4Qxq/Ig8qRHL/Lvt6K7ZvfiV1PuTjdDtulAekmTUAZ0AcbA4sTbUZCNsknHqvEU1UXkoE+s3
adUHheW9iuPGuV3mPNjj1p2KFJlwOo1REFb1oqqLbtxvUJrREn8uWuDaT9DyLgSgsh8DosybEJ3V
OzpGRyi39DyR3aT8pxEmfdDqM1Ob7m3Lp7Y//sRwYMZCT8sk0GGnZaFY0Qx4X5ZO0yr+neXGX/3u
vG6fxik5J5C26+1CNo5djBKFXiZI5RQl79e6wxsdqHvCIAbFK5T2e4+ubLQZt8J3Q03/8C7uGinA
gquLKipFGznmnRst9zLdZsTwuR/cxcuWl0LyLGIcSundKY9ZoJMyUAMbGeg8je1vJ9IiwLE2H1Ww
GuhU5IKFil5NVI138NaT2kK5Ez5r8SYlN9g4TRtz6jxoqXW9hSOSFWNR+G8r4R4PiuCllWoUBk74
Airn/KUmmEQIqkvLyaqxXbMC6E0OSC52EmVPpynJQ276oT0Z9qiBc34Gd0tPMaGoYicVbxvGrJ6c
a7rfYHfLoX0NGukR2QdtfVMfYqOK2cYPOWxMxCkj7up04o0MxVnB06eVs3OrbzQkViLsH9kjcdHf
CFZFwf7UCabQvSSx1EUkbkKu5ZwNVzj9jE07mpZqLOGErPtxdtwcwJPiyzj/ZeRtJEiSctiLzL2t
G5OAVSe9rTs4CT3fs3alymtT4J+dL4Qp9112zJuWcqnmA4LdMdTpBZ/jaVcQ0dAnKMHRWZjvjqZW
oKM54dCpTuKr6YLidriIjYC4p2sA4uaygYb92ko98VpZ/QQxmCiDtIXC36Ys4h59QL63OdbEQmJr
k7pOH9vLiSU67gxKq3kETW587jfv0j808TaCprPDYBoeUgaY7YhcxwSjgJqF+SKdtZTq4YxjLpFa
buJOl6VU9Cb87fsrQsqCUUnHsEAw26TveEptA0Oiaa+OxbXQC1xmEc6TN4iRcUNtpM4iCcsyNw+9
fmDfHE2srfmf/3mfCa2Oh4054GT7nOWVxc3fDEQ6ZVDnI55ySu+A5F/icOiqSNnEOTSWinbXa2Tk
KR2mbdx5bXzA9yAnbAuEkDFoavlula3Ug9rnD7yx21iiF/7coxLevjewQQuh4AeDPcZD/BCGeg/P
ApLuX2q8Xhy6UMhx+qT8MMsVsFL3u+9iwrOJkHG+oD/8O+e9yalZ4AuobLAalIzB24bGbQzzsF+Y
nHspz16aQJXixT8bFpDPwWYX/02NtKIBkfA+aKRW93WHdX7A5qLwnW6b/q6kU+R2AOAhEgCnzQcJ
gSquhSJR2mwCmCOp3X4YSqjfaYZ9az93BeyX8OvTONTr0zYXzIUXF8Cj28kOtOW3OM1kxgeNR7kQ
9c94OzrGp7UEONNGYj5dJwQDmTozTLIsokFrV4zePJNVbJlQToyqxM3c2jNP5f7HiUlVueDVUREd
aIXyvNXDnqOHiN2YQYZ/1YEcPDVm7aGlykl9Lj1NPDLGK896kYJbW7QpA/JK+ipzMJGtqZAaDx/E
sN/8XcgA7jbOl4qITbEyejVaL/i7rgkUYtFLz8RfuhwSxSVdjC8OZdKP76I7+C1vf6kXpCpY/iN0
dY2iKgwXQmyNQZ2HWqXbTpOOZdjjMjTzFsLhvy7uYrR0gABP20abYcmth78dKU10cXDOPZUKiyJF
lwnLSYG/BNrcd7ijaj3eXjJD7GJlVxFpvIqKHOZ+NKBFAxAHk+J8KEFDUxTNDnBbl4iRItokdRG7
coX3oM0WSBLcj4eeKHxiX1Ae+n4Lowg5boZrKkwyIRNVkAm3sXgGMf9VFRsEMXu1rzH7cV0eqU+/
iT44rpSWbdtLmCVAeeWI5PITYOLGnfnfR0+xKMrTVFxwP+r9a/A4XKJv+iwzkkoBLp3ELPgshPhX
3DMpD249GlAyWRjFKhUGPJ7k01QUsH+3a47T0pcYcQozWlQSIsnMs5QbC1LkbABmGaGICv8BG3bS
2zVYt6VIBJqN4mXMPgX3Z5RSj7EYVaF40d1If8ViLYIrUt9eFK0zZ+elr2I1ufSPGDv0y4NqHLc2
H2RoJ3R6hIzwlbTLTVcb+MYMIzp5zn/qXNo1oxocB7iUq/nn1U+LsM6p0d0KBv3Bl1DY98UfeJsG
09jIi+Di0raPuCaFkMg24GhhBqR6V8wtQ9weLlJQ76jJZClphpvNd7O+vP0N2q9koKhdL3mOMgIV
Ch+4Ye20q+XcMk514qdEwVUKhpJ4QWiDBi+78FVLXDIIz5Q+Ercrx2SUQBsZEGRk7IujLnAvPwBh
zgVSm3VP9qt3xugIZiTezk17l7P0xHx/Tn4X8e1JMiSzo8PLCvzdkPw/iBPVQmMHOss9T6wkE1kB
BLr2hT3R3o0raXXdCTPFQgpmhZQnozYvHBmMgfUk7LQK/kU9S42N5N8tBrUsHgRgpNfGBxi76/lB
og7wTqN2IOePXJugZUvxr6HVPrWhyC6Qq0TpL2DPtgWNb2dHU8GiEnOJPf8ytyLMEpG1tqh8M088
oAfHwHt3xciVP8xF7kiDU3GzGyKP/6UMZ+ZPoXRLyXKOQrcQiY/vxVo9/Vb0WJTE/1ZjhhsY+sRV
s3sK1xbLWDVibe1bCU0zdHle7cQUFtQ+1HZpCdY727Y+Njs0GD+2mN5Zp/Ys00P2txWbIqBH6ZMD
WEbL+4GrbKRBDA+ohJwrzidcYkJm16Jf+2dZwA94O1eF1MJysrPEy06GIJKuasaP4TmB6ypKF44d
+3H5A8M8Tk24Qz+Tzbtv6mZ5oiiwkOmBabgxxpwhaDYGRdGIX6SyBRtFLL1mlmhUEwizWkwNp/MC
SwdTT0pdHQbh/Rb0hadCVf9be116tibSHCS5+6JGh/D+x8OOikB2XA874lnKoPtxvqJWIG55lP9N
FWNDyDukr+zbQsrrR9rHsx5aWpklD1/J+xZhugnpWSDgYMuJVKtPTYZmqbGYlmGvIsbMLLli5MZ5
L1dkgiviR5HtmqD2jJEpKNpFEYxjP/kw1K/maWPSUMkKeASvB5HM4NsoR18qeqZdDY3nfMWW5wGo
39NbEOtOIfWQ/f1LtSq5BFM0R6NCWwglYmywM7n8d51kRkBi8pdyabraNWwg7SMiSji0oSVxJjDx
l3jh6puyCWMLPN4eZ8i6vKelC0KJ0lwUbYeY6h1TGTgysvhWCo1EuplbrhHmUr5weh4usOjv1CCS
dB3SYWC0Ctc8oARXwwCdOTth1LzEMI+SsRzMue4bzu2Tvi9AW9W5wzjw78s1LyuoVPv/m42g+Z9C
XdgDXoDejDwUhTXxBoLM1Le6+wQYWigSD4+Y1ak+Vn1NSwSohE/8sXia4X9fcKYnsTp8TC/zLdzV
JNnQC2lVB74YBkliznfqZpsSg+KldwbfqtcXTRwXsnNgWcqAjiyNlhZexnw5jQxOMT5LaBbGUfki
70e3B9WmxAl/UT1KGHZ/Flww4Im8g0farUsww3A9VetnnmCtQGPp6oqb6y9o7yHWNXSZwed0Shtq
ao9fSRv+Gi8FnIN5Cza+az1Xj1cd/fZye+I1ylYu0yZA1UZDjSuu5fMQnMaqHAPk7FjGX1DzhpbS
3vSxmTEY0fIzs3SK1CWJVIewRO+C1Jt0QNyCwVG4Ru+WhBp48pHICDgatZapp+iR6vYqS5muWpAQ
orfQYszcs8blXfBCmHE/aor5zjmU0SmgXmgpLunoNV1W8ZaNNE33ItPxG8BF0zv12GPlJeuGYj4Q
GxaQLMR+yV2fSyHdViLgNPMqIeLFJaKsIrIE5r+NzlSZWOISEgIdk2jXSQlw9RZ6xSPVDQ4NgErB
b+xDar7cS57yYBSCnDHJitrHP1hWIYfU0hRZhzuPlLgludmFULY2bTU0YXIvCapIwr++n7xcFfSH
aDrpUErflPIp/bmw30deL98tngQBAFYK/dgaHPXs7++aJGQpMe75SGJ/StBlyTc6Yr3wc1HBJxZe
iBSnZ1OminyOWCaGvzotRAHFKVh02pcBbMgZATTMD7ZczXrl3je2EGVSt0quPQUG1OLLIBhjf3up
4SdwQfsMFp3dN99NtwsdrWuZFfJNAY90cVT4c1lrRbfb4bhqi39DZ4J6GhJwBvVWAhcTQ2j04zvC
T9fZzTLvhQi/h31BNTIEiAQXSfpXpL5dEJ9hHDDvO4bt3nKshB7nczyJak1CxkxtS2jAOqYAl0cp
Hv/AI4E5JjK2XG24fxmoS2PEC2Sg4eY9+oIWQIqNKcUUjuavHOtBmPziS3MBaZWusr97pCcq6wxn
BBYxSorHfhCXDRyD5Zl52vq4MleT5CBsv6QlkMj7+C30e1rU8ud3ZJ5/qjS63wDhIruAgHufRjHn
gViT1MHnJgH0NOI/d7Yap4jade0u+kK5HIZhl46/fYlGsi1yFMDNIEquLUVBjPzHHS5pOmR/FVjk
fG0ykwIpElaGYXRpfmLWxdAOr+c1dHAhQiO6ywBpMh8VZ2JhdK/ByFN7RsO3GAdUKgwptIJULpro
eI6jmR4AV0m3ZF+d3MxnDa+r3kwb6KZy29fGMNqlZWlTgfRsUxRvELogrUvxFQg5OtdRKuqAel7D
LB3eRSJOUqZiZ5ymt9n2UuIGX5ui1wnRT0VZOWFZY2Q3Uw00lU+HPgPNjuTUgp+5qz4rA0sQ7GPx
6TFFgr2+ygz05D9tN9UwKxBySFZDBCbyggZgfkqK9toTvoRKQ68S3Zvx2dZmQPBnrYpT2c1F2fHe
aENFaFHVEdKHN37eP4FM2tmW3rp1GlWKUix9qS675I85bjRCCKoxBStic+EMdG1rLtK2zH1c6lpr
3RWWEjsCAIUJJg4ylHRoEop8/+w2mkr8QKLU5heuLH20JswBRC5g41CeK6DNHPmDShmKs6FtWcDQ
kLld7IPD2J+aMiRQjnU3aC11ODK48vDmkSqbn+AwqfMWfU4jEiB/1nlLWrY+sgpNPqiLd9nNw74M
7BWrd69FFsM272lXN8Dt9W5ZD2I9gn83zCzq3X89XbW9nz3tC5V9sjCQOwKyF4NpuT2snT1MnmO1
FUsxRz/U40t+Rjrbw0sKBKx60oleNJS1UyyoqVD9ZWhtaqyTmeQleWqzIYuXOFXBIhzVNAwCkQ0B
ZORaSH3lN3G7eCSnWA39YyVDjvxHBLCzp5sgnCV9qne1T890QY52QdaJccss8EeTdLHhnMZk6CzH
L/jUH2Y/qJ33Re+7Aagf9iuj/cY+EdzKWaNPLtXvqKApK/69wrvCBi78gha8cGgZhQ7X8Vsa1Ewi
ZW8mKgb7i+qr9BwjUUTtxTG+/uem/QZ25XnCt7hMcxOcoXNuzdxoE9FmC7X8zI7phMbgSWnNzvvZ
uvODSgDwUmBZgTmhDBocP6zFfVwnF5WfLJOdum4buNw3c1BGpInk4gc5wpre8UAVR2A8B1tvm4M/
xr7+jinRtfbRwu7wnOqThdd54Vq+sG2N+D0Jej1cLiMce2L/Z6KJWnOjyx2NrQqLamRIfG4Ud1tE
9KI8828qI6mXCdu5OQoxAxofvYpj4Vr69U96ddFTJnQyM/l8x7EejB8xZwl24K9pQ/UDLhVztXoY
ykaUwc7zjqpjKPWNA18vGcHteC1G+3gMaVVVMbshPJA53GqdQbiLc4RsmL84HQN1SKIPfVIq/pqm
nkh+Sekrks7vaq0/20+ccVoGCj/Mau7AX5O0pkTN4aQZHY5ec+wZA6rfa9ocsqaxCX9HXVUj+84M
LPcHz+VHdroj7L3lQr/bjElaAwdc3m5DcYL/QLZQgDKpsV1GjROqMGK7HSmNrwVp/2AI/Qh+kCOS
M6xps6zedHGEl6E1ocwI2lqcvdjI4jOnTpZ0tw5gZJVbFptMQPy/ExIMwLn2I56z1DOZ82MkY6Gq
NgF79CWRVjFEuGkMj03KXQlMCMB2rucCvLb1GoNnMdRc6FQWuilxPIRqgYbaREvFM2dkzF54VEP3
MUkNWgwNrLDjAI5Kr/br4LGCVd/ThEHIacXz85EG7TlchSail5Q1VBMaTduUm+BXWQ0+8cER00Pf
Wtfcek1tl3Ma+LRIzSk/LXKi7ZrhmDAQWDzwnQCvDYSq6tXmIoT6P/ix9Ua+FgV1Kah1qis0dMlx
09RRKCXAh+0GGg/KCa090ZBI6bWKRrDzhy6zcYhnHz6vWtPpoLCrdi3viI/dUNwl8YPUHB9HfbMw
gJa3VlD1W9EeX/43PmkS2y73htN9z20Ar6Kb946uS9gBeuIxNipOAVpZauDqVWtkEFQFSea9fvvw
aXnjtF2vNOoCFue/S+PAJEkNrXI9zLFSMBRxiGucaaleiGKsucmU7y8ubwjuOIjbHA9cFwFbeIgo
HelIVfISSNyZmXubZJnU6GiTGiHm8skV4D7aXFBRGZyVUuAIFvREVNA8lvBZFw65P7NdXVx2JVrO
RQoz/mRciaZDmC+0qL+9oe23MUZC/Sqv6hTVraYPtQyF52ppt4CbvH8AVlKZfX2Ouh5ITKYAhgmf
0zAovS36TxgKaa7XFUbyLrFu2sHYhXMRbdFBWkVRdit0WBwVp1WTWUAQlpruunkwpywoiYp0F7PA
7hQs+cJD4+/sVpn2L1wl7Ax1nuKKfPvGH5uY/hc7S06kDBAv1uLrxsIE+iXbNrZ/PRtta3B4zCy7
9W2ttctWbMOdNBhzZfooDrCeo6/Axs8TGE93yl2vVJVJXW2UnExnOqqtm+Ff5sxLUA7P6J8WzE37
AywSrTM44Jtyybr7dCPbAI79ynAT+/moWCAt6qgcfD+sx309n7TgG9dW5myTn3ROT/X3fTIGkaOC
lp8mUpoBVor0GjywLiU4TFYUzOZllek1wMLx6WFlDGAVDUYuD/SgHS79b9pcfBnpeXAoKUPHqWc8
aktV0kRnW/7wnIz5WVtaeAYBvqVaWlHBDzZ67wvNyQLO0fqS1x4vqGcGbzm9v0/BIr9VisQI79xq
htEox6NKJCczsMG5dZBEX33bjGOALcZIRNi22ggt1BTy2WUMnT/dpbIKDA1ZavZ7ErkBUzQELfi8
cFrNczB1tqHqegpZ744hHRoBjCToXmsp42TNyNNzEi0CRhAtsNjdh+wHC///SfXJftwNx51ZRE9e
dYa+hp0CKdJESgk3T3vKMoxfxV3LmCZW97PjJx+js1dXj9Xw2E3pRJBlanf5LMQK9zCJ3B/YTLK0
26Bvt+LdDnrIIm2Gr7AzPhpYkKAUzdYsUhcsRKi2x56YivXU7T37tGsbBeqIv1QyhOoyr0+2rRhx
ghA1+c2oQvd1QhTufJasVd9vPNg9NolHbrD3Gpk3UpL9tJAMFw31MxtyD+QAumhhBKltVO6WNNPR
3LaQ9M9iaTH+R4xZZwxsbGIVqK+U3EBl0O5CjrMYnFHUsRp0eF40lsJjrYqEU26eqCr/Sa7Rt9tH
90KEPpvYY1XzXknFxWHR9x96580j+MQcgP0TD6wBpu0lia02XP/vu706KVDqkEp7D3Bv09HHxI5b
SLjsS0ibIWd55Bn+StUdks0CRcSby2N0C756pM1NfM+WGivuyOylbRWLZz+Lo7BjhmI/NqMN0Tvf
VNUWAuzEvNeowusly7frDKFhRO+S+Q1+XDVTaYZTS9Guii8yWKJZtSMUmvh7yPPuuYmxQKLrGPuM
ywmgDGDWNOv+ZpHfVbILzzMNEhJNY7zyQKH3otKdM5t4safbrHxmjbUUVD0H5mqwq8Fb3OivJVR4
40/aqVw39p7d5KwZPnjaJpJ0lyCRvRDjQkOPhZOTFliJLnkDD84hLtIaa4jA9nUneHTleyCJkvYa
2LaBUMccyh/J5QwfXRZnP5XgdcoyfHVp65utfj3L+6cJj9+22IlDJGF5rbXZfXfG8ZkqbcapasFu
a9kcAYc6gWzKPYs+Ku+muMGeEza+7IyaFkEmrPttQ+O5DPRZYKPoe4Fnx5abVGAdrGz/PUWaNQUf
x2xciNi530ZpmX2cmsPeSwsxIz54fdtnRgS+xMzmH1JBoHE4AtHuX3KxiN2t3sfAEf1gQVC0jw5j
MwkLRhbHumPGpR4DuEmqEsV19xuRc+0rDiKqZTMlW2Xzfnm0EvlYSI5ayfXfgBDoT+H+vv6llc4m
KOWiNlqYMCSId36gSlqFfXgYgMNW5k+9Ri88jXB5pjPwdl7TQDKMg9Fb7twr2IQxH4M90c2WZYUd
QBNW1HhcnDUgE/pJsd1XYX7UGTtqqpU3h4bTg+X/lbWjZs0Wn2pJxuHneXsQPVGrCwKMj0GHqkW1
l/ywwVJyWRwOFDPeq0G0JRDhED+/iq73vI55J17D/KInqQrscPt9FvDjDqczCXPi/2pkCp/DtgB7
q48aMYbb2jV7BxnjKQBRolV4NS9uch3Q3ypVOvoX+wwrgSm04661jo3AftMeQQ+GrTgnrDHxBAzE
85JoNeyyS52MBtVA+c+oe9gk910++flk9uEX6kRe2h4hibVq/PTGnKoI7ezllRCV90YA6XuU/I2O
t/bLIDTaB2ZVkq7lNxxDDJZHJxlo7gxJAzo/ylhq35Zfkl69S9CUvTBOdKx7SI9x68Or0qoNxcU/
glwXuGLLLdRyRlITxO40Hg1C+6tsr4XqQV+g/uJfx5Ljg+i30oMOCOqWiObPwA4PQEa7J3KONSXw
LBp+U/F6Uyi3/giEYwKGXEEL5fzROAM+EsLQOk3mXGgh/n3zRGyn/f98n4YHaY+Sjrjxx7xjBbFw
UehZCv+UZyHKRESvnsDmA4oY8FTAtcGtNcf+I5tAIFV+TPdCoT32cOQKAtSLT0JDM2/8X94mgA1U
eIkDzX5/x/HyGUYaLA50jEU3t7/FHEqToP35DzMvkjEDFsAQPBRthzG+rsvwSQtqpHfYrCwigTCd
X3y+wYN1W9KDXl5HUeOYU6gfjdbAEHPslQrr+Gjb1zCZFd25w0S5vWWHqXvT5s+xcYlylotpgPP0
AsOSMQn21/u53YS5phIbgs6lpDA81mQ4eFMTUGl9ElaRVQI1KCH0031CCRf+YBNLRwWoxNrl85xN
LITo2Tw/J6hWSP9cTblIxINuBhB00W1n6hqfSVO8bwJ44zHExVvcB9id7tNta6dz1gv8qDzhlujP
93DXvOLDIHtvvGUKOXx99vadwfq3IY/Xc85aK+F2c/KJ0pU/o3oUNi3CLqPNmbe4rzhxUBuy3AWY
RLnd2aZpfpL/6vWFIVPhbt5l1imQr7hDa/clnPGfFHf3HeBfdD1DImBPYdmXNsqlPQMp/nLOunEC
t2t/PoCmtDsSKR0wo4/PfQYdhfrkhBHSS+G89xMEwWgTdoPzX5GmofU6VriZtCBi76nE5V0Jgw/O
jezmHvK+sokrS9/eeEPyfuOIISU2LKKu+rpW0MA/K97cfk9UkP80crVG1HZEct0SjiJLz1Dw6DoT
Gb9bn3yv8my7KDDkk6r+e68HhnGz7G89ovrDcuiTE0OQYF8UMFZKy4wkTZy20ssUREr5M903cSpF
VQ02HpDkR5jTWsS/fFdGXM6Ocu0JFdvKhfcH6nEUAHEU1IsYg9ox5ftBZxRdpe/6ZdZJdHH4c5T+
7w9getfK2Rxczze/RRSCBP/JKeeJQvSF6MK8AR0QlKyZ4sq8QD7/i8DAvIrPey78Vsk89FO1oC6/
3gmTKD4OXCZ1zL7c2LKuU4VxrUdNmTdEhu/SyetQgStBIoRVmnHuB8ZEL5aAyO10YdnA3M/x07nK
tEtZd33m8qX0f2anl0ba187y6NmmLO4wk5DSvm5inBpx/4HqYgmd4xR8WLyHApXsH5t9EwNN9CTL
IUm8dp2RbTjsxjTpQ+rvHzdBGKWXgec3k7yWPWG2xtxMkbol2Vyq6f8ZYIpi6okDJxuaWGPwoXBR
jNUIziMhZowd6JK34+GZ93tAEsINEI1lCXeaqPk0sY4rDzJYTw6cApejKfoRUfg0XvuI9yqdJpzw
VPKrMl90Z7hRi6plV5pNdxVd6By3EzucLdwDTLg4pSJVrLt5bB0f649VQdbBaf8hUDGCCjZXuucl
g85rfjL5MpjkioMMnDxxbHMLgk053L63lrLAPBCqQDm3KWkte9N+x8FhB4n2kZNx1cjvUx2AGCax
2gd2mD2II/7Q1Pq9GMPvyPH3WZshBV2aK4ITjEeB/nA1wrDJ14JnTQ7fWaVTHdXA74cARn0u3Gpq
Yf3JkU06DjP6M9R+pZsvbz1HXD+fjEssV9vMC8S/847O5TXnXsP5WOwQ+E8XxIdCfRbbl9KGCyI/
o8aC61px9Tv0rd7KZB2zj8lJ/HKE/V4lMicQseso4pUM7RJ4I7+Ay9Jo6AB6ivcV2+1x1cXswPT6
DIfegVVHh2HKhxl8sAn326yhGrh9+0XlbGZepoLS7NT9xhhhebQvKVbLwCE5D1QDGOxaqBOX68oq
pSxuMfzRsuZTY7RHnU+23iUbLP/WSIxFlalcOpS5GnoVJm2lMXgL+aCK23qWZbXRoIf33dhuEERG
AcuqoCa7nDypnB5nD/J1jNj0/FdTaxo7XZIfxCswHYm4+r+zcz7iKf1ZER/I+0/YsYmKyZwF9h/D
FE7aNVNouHn3EPUUpWn+ThBMP9FULNicg9sPtgyFP/C+Xq4D278D7jZXkuBJAAgg/dvCehZTkqTl
wfaiAzTnrmmq2lhQJinsgOx5NpwT5K4spi7XkkIulwrF9C/jqv0UUdvowM1rdTyyM3PdtM3JWKh9
c4KMrSNZAnm87YNIR2SRolDajvtB2oLw1e1MMjTJlAIIG805t+Sz6DKV8ETxJ3v3MRg1TmN1Twwz
um+1qZfljebnGEZ4grQRQ1CPDq2EbzLG3hqCkTWN+MTuHBdgHN41grl3SS4uxfXobJM/APvKa9ID
85cHDLazcanjVPInkB1iIzMH9HoWJ3z66dvKoUrUFQHRw8oOujOZAo1olNujpQGQf0+etJbyBfRS
F8CyQ8nAWQVjSumdEmWM2LcwYN3K17JsXmBFGagj1VaJJqZaXhfdaSZxpCkUCgj4JG8MoPC1eOJC
K2NnjFDpKfo+i/ba5UocF07ouC7G6LmCkp5cd6adoOnrOpXWP7KjzXKUVt7xeg97r0J4NOMg9ICr
ZrgboOpOx1WnKHk5jMvtPqpb1GxQIwJk7k1hUDYjWRuz7rHO183be+4c2AjYcNNGeIa1ao4NNYId
xOVary077r4r9orYu5I9LozSTowQ6ZZoHONLDanM6hqqvEDiT1BS2Fr6nE5W5h/gGcskcF99FTo9
DwlJdSxqLJNBqTrs2Yd1P9gD6YIsNYvtGfwncmSQzUSGtx6qFnwLkVTwEJJmzJ3E/fUod90ELXTI
BFYUD7WZ5JiPeJ2rZNctzWnqD+HSMVvsGd5y44CoQv0Q7OTD5sT15aHvYCvnFRKZBTi8irMbmNnM
v8t6fSb10mpDV/H1xwb50XHBZGPTuZivAe/FxOzRRPn0MrQVErszakkwVC/Rmokff9KvwJ7An/Av
0CbottD5kOm0J4aNsoipqb1k/7vOEbNTmrx4Okv8ObFylHXrGCnQ+UMlXXaRvG+k7Sa+F0+/sp8Z
CYc31vSM/zp0ckKtSCXBbEI3BU7KTFI9KsiifARe+XFvfnJ5orhuG0IF6WPj4pR+p9jhHInt4S3Q
dbVnqeWsBDBfHJtXLBjuynigqsYkygkjI0a4EsyQXo5pHewDH5UHvEGrCorY+PZjStEhVn1jyrX9
HGXHvcImBvkAvlVRV/CYaDLS7rYs3X/jPHod3sBoiUMpJClF/Anx+MaKbpzOCKaUFwuBc+8CQ7Rd
kd+LvPbpavNE4q8ISBRm1OhZGOCyLpq3haUn1mk8+EfQmIBkBU7SuDCzoAMTmbJUybgooAxnkJam
AC1gKSWXim9lHe6+0w/aXhbToHGC4JPGPZdV3Mj2pAnw9sel1xGEn4XoMGExwJTAQzw7Z1UsePFQ
NHWkC8T8lKNt3ubyPzXXOrpmAlGqOgGx8Pc3XctUA1E8jpTGHbLQwZk5BS/ayFmY9CuEV+urCHe3
kr0sDOvZx12PY95hq+N40rL7butIjEDjwTM2+ltl4Ug3LpaZJK8FbHl13uGmR0JLL90SkKSjsbeQ
0U6jUp43E5BrwSeURa5OplM8zJ5fi/H/G5VgVKVW66wThugZeHhTRAYWTJq/yPq96aqjUQPlheOW
y4dlVayZuFNo8Px7tT1SUUberR+gIyPzYQ6MvKZm9NOrrJ1G7zlKVe6ab01BKGhLpNwFBtcwpUod
wtYWTPCpZCLd+k1IZuxNRxYkXfOw8NGJUTj3iWlzcrjEF+FxxSz1fJXt0n388K+IDBjVGu/MaBh2
FJp35j+AvPtObhksjH6TEQJIMusk33Y1t7PwtlP0UQ7P+IVUkK5DhaGL8gLNl8Il2DkgOi/Uizv/
yAjAG9imHnrbqPvDB4xS+cqVC7F6VlbpPEm6coIxmXjOZaLimvMK1mwLWxShf4SuLsjJDU9P8AJn
F/5i90qGUaPng+EhEnn9UXvUwPg2toUtxmePgwUpXAdDwzPWhcKMskEBOyE6bdjCI4jjfbQ6HTC3
3+EqwRa4ond7KjctxK/pMmchZ1VtqJbcJlzvQAgMJsMjxwBHsoioDSYeYb8faXXOtgrLrYNGsKyp
277b6LeESuZOLmgkdcl6J2J9Z4xYXDoVIdy3vkTtEfg772Zk03L2hKi/UBh3SesbvK0y8pgMvX5k
OHyORzP2nvv2i3EUlG1E9IO5MCFyYmL8WFEelJve+Bf7b6UGmLK0d2HzK3KacG+GYsYb0mLlVeyG
fiwIPy2AjjFgrK8SQTBfo1GTr9QmoTqsjuGHhTn3oKNwlaGjIS+Kpn9t8vc3oWnh1FYazKiE/fEg
TagYemWORsxM7IESx6WCeAgqHoqroaWD3diMXBUGuQAAJqg/ab5ruNVygr4AWfuYCZpOFvTiwZT1
rEQ/rFgb6Opz9DN6ToljaCxPU4v8/VjzCXdjfnjdd6FkdRFJLncrF8lts5W6fxLg4DjcnYPHm0Fh
2aPZZ9hXsKiiaj8LJGzVCSn70LNWS9S9d6sRThDpG5L53uhfhFx7fdfvmFFc/i9IfLWJTcqnf7Bf
OVaYu5TI1B0zcNtYyWOkRns8S7nflUEfDlWkyw9efpEKb0YAHiXtFIVnnWkQxWRjx/Jk8F+Jh3Nu
dV0UmU8V+li6FGhZycpjdpfgw41RBDlH0I9P38hP8eLPUTq5QTYHXzV7W1/eOyaULoiXW7QXM+bK
+Wj+UzHt4GSO5cHp1vwnq/HxBB7GA83iSQcsOhPK7LGMwMwXWFsDo3WWw/Yx984r1bbSHhOZ5/MK
tA2f/2y6oIOIMaAgIkD9J+cbpBFam3yoTyopVSp5O7KlzWEMe/q3broVb6Il9vOk4iVKfj9SLqvS
TNbpWB/DDfAN8yl3h3ISh4SXOZTMGwA0z6YDU4Oi14h0H8Keu3bOf1Ks+WDf/1jrdkbLCssY5UPP
olU72rkdxGI9/iaHJegfmqYmDRZLOMrn5XraslQ+Gl8UvO1FiVLIca+moLOLqC9eU5yM8jaGEo38
JCZ5tcIZSEbQlAhkqfIU1kmyGRFcCudVounWFtJiz1N8aFtseLiY8lcYADejsd6drcOFEBMe2rgd
ovIV0oeZVo9O1Q6wIkwr8P25lLkF4XdkyjjL2whKtwzLy7hSeKHAdppUYTJmS5QXftK+x0uwYBa/
LAZyvrn4hgftjqnY+7wvp5qOFFiR0CQ5Sz5/NTDP3G8A994vyIsxkls3c/x3bHWEjSX7LmuCGaEo
0495T+Ar1uaByAjJQUCD9KkAV/XUWBxZcRzHsOAnfiesbUN74saMrj0vD4JLR4GR63wh54Mnq8O1
5hpitkppV2Z8/vIhUssq6rqim5o+hMSZxKGkfDwbIOFkXd/MeNazJ6U0pFsCL7yTb1ONYxLb7x/l
r04P3ZZMQm3zUrkXamM21ZOx9dmW/KC9kZr/zv6mSaLNYFVONPdxWsoNAv35WKH7h+/XJBxYnxqM
kjzmCwed582WtJ6nBNrx3HRbRwB+59SlBgxTGRD2eHIgZj+p5iJUvurbNmnh5D2vkN0d9DSDkav1
V0ne/UHN90AZQoigKal35VYi8Wx50d6AFiQde5Qv1zlk52AxfbBfmHZpcXeb8GseJb6lvgSHNsib
30AdTIgECfsu8np5areIFt207o4H1a7SuOcicKs4kjz1EZ308GmPNmfRvUUkEnTFzwGxGRXNPCd9
NSs1bmtVBBqw/D7ThH62ffuZUNDpC197Tqj39ilAWxL43hejWa0VtWP/f4IlsDPuDkZGJiM1+/hZ
PXrszxq4f9p0HuUKgEEA99VPNsXqP/TijNtcsVA+uO/ifqWUNJe8FDvHzgWT1buWbkRvlE94yKch
yPTHOxy9Ef+ChJ1IbwauSYihozerQs8YKGJauh/wiP3evYQHWwLmhA9zcIKA/jMgoxnz342kxhyf
ttZ0LgAkCOBUUb707MozNhb9OtOfrPOxv37ClYhTyw1pWxe8GtXGy8V0i9HqV4sfCO/fmXCrfPsK
qSJeN0naGXh9nKaUV5iMatGeFvN9i072FL/gFScHfGy6WDy1fTRVU75NCIj8lBqqfNgXxTTPHQMD
jrI9lGF5IPmXrRhcZuqfU2hG9r3dG4wCv9SEDgsHp8jaGF2botjIDU8+QshV4j2lUpz1b4J5/ptd
tMhAevacT1n998prh9TkoRsDlSI634v8h6SV0OR05ZHGNPeR4jrHa3tP+a3/lo1O9apGTKzmBQXt
C5UbnR5XT8Hn3/3ztUi7sUBJhQB7RdpnNSowpebj+jimhifj45+yRLWtxDL2fUaFnNdahAKqzkhJ
+hG3CewwU9PzYdJlWw8dSAaZlaTcwWUG30pX0cOwn6HWpohBPsxLWD7mkuavYV8t8IxCl7Jxvnym
Jy6+y8DpP7W2xKYQeOlZc8mN+cvJQ5QF/GwovQdfZ5NEs0MdkJ14u0/x20TyICoLyaYysnFARhB7
mqLMu8yhHhA1vNkXBkpFvNQbckgPhtUguASH1wZdlKqRQ35GqWz+rFM+OtmyPbHIVGQ7bPoN6npC
LKsK+D0jIVGAAU6KXXyZAScLEKBKvpKlOjJkG8hVqoLhjTBIXiNwrB4/R/SAwmEfTg1HyN75N4Rh
5OnjIlON5gmKwWZevXr7+h50w9OH4zfC0+7WC2IQIQrRtKFbnX307IHPdCqBaRPNKMWwPlikaCtx
5LxXsTrHGqGlnD9KBMiEJDsU/8ZcLg+q6V0bWgqgdk+VInAe/2vkxO5Tv/4xcx6JRKPAdwCjkAnM
GgCoaqZEx24HDvcm7LPehzFsACLzhTPQBCwgsWvdne19+9y57poLuO2oN1e0QNG211bjW6oKMf0h
EMEDXmjIZmTTDECcEbAs8vGgU97m9QJzcU4sgMLQGPGqbHBTfQUIqu1vuJ0WYTdOadEwS44iR/C3
XqzGp8C3e/gDH8TFLt2eUesJhjtqPSixrprIqV3kPSFri0sv4vgWQczBd6JC0YAmLQT8Utv6977x
aEn7yrEcESAaCOhnW6N5pGNFSeEvaOOWwS7L/VfNRvWJA82LNsJnaAC9S9fJdhvll1tV43eM2Xb+
WNm/7ptC51pA45PQAni6QvoN0o43ihJ9EuvrgiNHiGPt+mUrEb68m8gepWiB+JOJG4IZKFZluY/+
XalgpGntGv3w9OQtUu2C6uus6FBN8AwBTCQemHpC8Qll/Y1Xc1i+St2OprscIzbnaH93bk/UaywF
xscONE2vfC3Q24cXT7csONHPd1NG8gtkchjR/m6snrdQ40pFhgxzX3bpk+So2Ra6LVChvdG9hgpJ
BG4+/0u6ZB1b8WIxb3dn7piarx+It9SyPtc8vT9tBdcCWax+H9c+u/Q6yedNbmrZ0L3srGIJIJ/h
6Vk19m+1IQu5YeBKrD3lxTsxgCft3nx30IdE+UmtAKTFQaNjWkdxI5oC3zTDbtsy1AnrKerM/dVp
iXIcwnz3YfmrwmxO4KdpHcytrI+cbmrFy2naxrUKJfGrdibqRlfR6+deE0/awiMbE7AZFH/1QVgO
Dz52Q2Pp1ZLDUACoAwUsK4pZ9uKW/mpQ00s48G31uCYKPJtqMhCmhUjG/WuF+PmCakkSOpDvy3/G
lBN9gHYITCi+ToxrxphvvhIxk27FgTPev+iMHQS/EQnKGVPFStwWLYQGPWztgyUJuLfhTmFl4I+S
Z+hf7rE1SFwVjItjg4llsWN+6y7/2UMTNZPW3oofCacn88vAklEr4bRLd/6Z+m0qJgNZRi26b0bs
K3qjdeZC3WXsNhVReDWVM2RxEMXkfmjyOp+Gxn5IQOVqV/tSd0S/l/MT4BK9rjQeuU/egYgxyUIM
mf4qti+pzu5g4++GZLTYJs2BaMIr89vGrIDIC/stf1PwAyuUs4wGwzNoafXM4l+fZTkGbyyYGcx8
YS0fwdAqYlXMOPlmAm3m0f+okAY/r8VGWgT09ldumJdP99uRqRAdgzbnGjtQru59SWBwg/JQ8jSh
y6HI6BTmuNpPLm5XdI1ykUhT/1mkAtpudkvAW1H9wR6MPRy3ziLzTTwGW+4fbOAdaNo0puspcbUq
a8mIYeysXjOuDGM15B9mIxgzB7tBx36nOGdvwaUWOZVbNqGsBkcPw5NsvXy3yjQCVpehTzk9qJVb
tNQGmY6zWzwKfmxM7uJt+ScpDQo/XtjoNMR2IrYWRKM3/H6UDZUT+6RNpuuxXwjzDwVen6I1h6ny
B5xI9u2cdMwu5O2BTHyaQov8T5bZdKRKxqiOdwBCw8ZE29fw91gVD2MPK5YVQo38ljrm2n+nO9ER
xE0pkY/iyjzXN2QXrS6YErFXQmS2E9VHaWTb1vCZTVrqKy1F+1lqtlE4dPrP5dZsHDu3lKJiZrRy
lIo1my9Rp4nXEhJQz7nDUrUgqjcL/gsdoeGY0YMXTvT+J6uCsxnDTFWggimlhyjO+A1pFLMqIKDR
Alw4ONckQAEKecv1daiMAXthF8BxCKr7zGGKMGDxVt8lJsHmIxICuMEf89bp8KEWOTo0+Llf6nEX
y7LGA0mrnAQaIrQS48eD0JUn6WoVUtY0ezV7LkDBcjPw1OLLIVZTGnRhxxd1qruYRd9INo8yHGAm
0tVKaopo73ZiWx3KCo3a2wQ+nGXmmsO5UFsccAxxnReAZ5cLn4+gBAgbwyL9BnPFSmdblha3e3X3
zHgtFSX9qK0oezWzeUAdj4VopwWZac2krnHwq53Mms0dlr77LjiGc+230n2r2p1wUQMvUkj/6IOQ
mZEz7fl+xaJIYcU8P2EogZJkTLqVsbmPddmZmaCmfMfGMF6Gky9BmsQ8wsABAZrZpfWJ96//E7Nx
eEXhICOmQzl4plfAc9rLN9gE6gk6vuMhX9OaE6+k81eTDag15R3mgYPNO3+R5GGMAsoJBBo9OZfh
FiD70WDmQYDr8fPTvcAPOWI2WJ9Hl1CgIb/ktA2eVsKaxeeUg/yYiUmeL8ujn1uVZ5SRAJ/oSNyW
BuXVCL+kBq2ILwOUBm0xOllt3FchJgu2HD5Ct6KGGxgfdOaS1T9peU4Tn6GFA88/Eqp3D39e8uzd
eqUQ50hOUd1sTMigM2d+ffCClGIA0iUc8PHkxDD+nuyzlcHCRtuKt6xSjfJMYXV34OF0KcIWjiF7
bhzpk3NYmqEYt5RN49K8apM/EsqtnGcFQQ4jydYVP3UdaviNZ3ciDyZwzDtTUMLkwVcc4A6yCYDr
9cCi3NvyzJL/TzGdbldqfgPmVaBjg1uBXlQhHz9VxyUrWIdb6fh9CtV1Lg2IUE8B9DyuSmBwA+We
a1zw1thKq2kMRq0m2zoHDCyyQnqzJ586KsptrGcqQyqeWOkV5c+I7aPE6FDSc0lxQnS8iHtvD7I9
dlwHWr5zRFKI6aPAOBDjoKO00uRpF6k7hHyZfVeB9U3FqI34kXPdqaJiGBx2+KOzmwgdm7KOwYKR
0m9Fv59nyLcW68FB5+8A1Pdvq2v8uZXdQUUNHj6cr4vGTCnBDURN+hsLGmMC1a+rNQBs3AgmH68T
cR12Q17bPs8kP0Xg0/c6TxYLKFxaAaoHuxliNvddRRvDpcGmDrWZOjvlWG97iwKlFa9JoQnJJDu0
zHoFSzMNmLMyan1gdhZog/Vel+WyUQVVpovAsQVV/20cw/NwkhaN7Rr4N56xB2w2uIiBW1mwPByt
2/HDPDjQswun59+yqAy5knclFDaxLNPHtMzTcQiB/PDo4NKptjluvGGZPUHQFIh+yHTCjg6IOfnA
dKCr3NSL+naqzMXuDch1TS9xgj+c+6+gacFp536a8asIJJ3uZJh+11ZZ47EpEsraJZ/in7wWQlh/
QEVcK5IGoNbez660cjUajrSdm+/reAEATedUF/elBzgaDyOX9UB/OTKpezxD/nOtd1QTZSuOo7+t
cn4KgwiHeJLryWqZilATEDKeqGqxmotqBeSiqeWnKgEmCWstIgzKwTPkm+J8eiHzauuWRxcms+KJ
+lgt+me35Zqogma6b/D4X4adcgLm9EXpICVmiBXTsTaW7hK+8hEbh9f5/anKx6tFOF0QokOS7tG2
x2UFFf42hyUDpD2onqzZ0oEp2ycxJ+QBxvRhLPtQJpl90gohROiopWl2mLWuNbD7kZ2dpASZ4jda
Sks3mTbrO3Un8Xbr2zevCBtr+7hSa3bIM7QzjHo+c4pO0pa4PnBIfh2yW9gUhex+dolaiPr8pvoD
14QFLf6Q9tpF1XoqX+tEuVKEpanls+YEyBkYBPFTKiUvO/Q3cocXYAqaxwZrYEFnvUVC+684KSQv
N3Y7CBoCOgF8ZCyEY91mAOFBpVqlnJH235fTlAGhaS6Dx9cExjq8MkujtrWgpkTdN7yKxDClNopZ
O84YwPtG33CXBPJRSJn5iCiRQNrsJgqI6x+8lIkiZYBlg27dBxjdwTjRZ+4v23CX3AQyWr2zT/Tn
s1pnDlSoE2o1CUAQHqrIwO6BueJ4axy2PNIZ1Qxh8jAQWevgnMiBTm6xISUBTqGj/S9mzKhV2Gy3
HOAofF1t2orG8O5PCuyW/6YgZO2Ky05BIpSdvTJQS4H/UUP9PC3wDmQCUgVpQ5o+pO4LQzfZwGCK
T4MBzRn7CE0cEkoiZdOWDwtRPUEwBl/36oDWIBYbc1BW/uxr30kPWdoGVpmexlQeMjiH4CMHaWHn
54Km3cQz0p3fdSa80qcguX7INVTBw4QwM6gtY/oip2qu3qQfaxtw+fovV5hnNa+vdecNy/n6odni
Y2Cr4jSgCEsHjq3r482r4NQe/SdmKmj6Of9syF6Ac8qFN0rF2+dTwPPw/mub6aQZuI3cf+yCqGDL
AMogErAeoubzttCF/wp8QV3sZC36cIKX99qDcHUeNkG1NnwsVP0rwjIobGBEwGtPqtwrAKnytJME
IQQGI/aZHQ2Yvvaje7DahsJgykyVh/dy0sPz/x3I4saH4n+hDtreGy9aWBvaUnFN0hN8H1rEa/QR
d7vPVOc6EDNMnErThjY0NCZe/hu/POkRAaYypQnDnEIdtSZEYH8Y5dWAY7+z6KwmZtJcboXXZNlR
SZK3bgYrK91+0C2gS9zCikSbhHT7ZAI7F/m+U4R8DrkHS4kYHQgV8Y6NF+OJkWm9rHUdkGaQjSUq
L1z+LKM8ytd3jP6I/mQTTHdudfw4WoHDZLXCK24nRU93KK5aJ74sDhzgqoJjDHQorg3aq+IyaGOE
zSoPc269O78a3PsY+zb84cESOlZ3OAd8jZOUVmlEHkPyNY4T0KEaAmlNadBzofrbxaYnuYHhi6b1
yfW+9oWqSJVVA94Lixod/n4EHcl1JkxL1CEoX7ccdYIAZoYwsrFTZ65WCZ2j75b2hqqDLkLrb84J
NrrOjwoxEoMGJZ3jisiVH6q+Ita9ZakA5h6BacAZSxQbT5mWyuDRc7xEwid5jWj3iC6jkcw3FLy9
oTK0l3ly+AMDEP5v49uJ3hwss/518D+KmUGm1ObWJDt549nrliMyt3LJ5nGLmuoY78qopNhVvpZ4
ILWpZ73FKkv2i4l9qPfMng23dch57bDVpytXVhVhh/XA09EynEKzEYccJp4zJH/8RXxaSGB/7Ai2
pfRDRjnCYZlrXCsmkoB6pX067R6JjF2RwwdpJghnjs5TaF6xjjeVH6ZCCiemGUY+WIuTDUysev3Z
G96pd7ix+5c+h4kfNR5DuLNVk0k6ctRRjytZAohz8AWjaK3WmnOILndJtsrI6fSBY1r1nANDGqfe
rCTutsRiJ+uHyg6m5IPwrIDIXwDqZY7IGHfqcEqhg3c01N4g9gW3bdfIYpnXspaBA19itnwL7S5S
UEgpkTNHE3Tsxg6LeiG73JrLFsRDWXbfxVnNff0qCGuy+FGSUBJfamGStWz/qq7p4niJGB68s0mR
TJCU1KBir+rj2qclV0Y8UWmAp7z/LyOfEIlaOBPokygFo9SR/Aud6n/jvSGXC6x/2UgT/h76nDeG
XthbNfNRouQ6DCHKtl3iUJ0XBlpQ+nG6fdbIhBYl2hRv2wABQf+0HDfIa0p45LGxUhp+N1A7IsIL
zTLUXBw1kxMp6Jb2kPgodZtSNxOMs/FZtRzDAfDkS6iEnUvLUVgOlOEmdkqtAz1TCW3vhSEuxFDK
v7IGzm3c12NJxFBTbgxeCtjixs/jL0oel/lNq8qptCsE97zzZk/5CeWoFdETSMG0M09k7DxLx1Uc
INKFHI19p2Ls7EuXQn/5KhXJxx0H1kUED++gAvMSjFN53tSuZlYA+tYHiJ3PvOIpMn5VTZLEx1HX
N9HvjYlnoKE4/FoYceaTQVpVqKdk/DhuLGKkXOVpwpwUxiPTh1f6zksPN32eAmdct2CTdSrlnOwi
dSoMI7HDKYzGE61nY5//p32p+Zf58nzuQrwlcHkHRsSTG8AddylJPrMBDjDNC8c9XSLGuiFA2qbF
SFLEZf4YwKmSUjhzlgSdvLyl0hEhEVFK/ZvMGVYOvPi62fHmTajrMoLUX7vBUljQFrPgr4MpwUhi
1I6FWkJLzsCjnp5FWyssRYdTDIGnglkg3D3F9fFaqbeM+yPGx+e9PxQ6OInBG2dmG2c6tzSLk6HT
dhjdcGGcVrgwkzhJetUs6xekaYkq3TiETQnk9zhJWPOqhPdJJW+AJlUfmWZ7O/4G2+JyiVWc9ZVI
C1R+nrAoIzsgTiO/3h+mI73N66vas3sgbH9rS4I5wlABOHCTB+XUgIuRMXvqrlJLf24J6ETWQ+iT
TpEGHkJ7lXxPWh0jwjC15uj9BpTxaUkYH3KIsk/vjMf0bQ1laPOSB75ErfGfliOoCUsjgW7x3oUr
KquYgqTARiH71vAMMerzlkxpQp4DtWysnb77l+62IarfVE0T5W5dQWjh6C1mxz/MHLZEGXrD1hT2
+UOzLfAJGQ54T7MiDCdkZC4DMlC5MPYyK/F9jhMcPuztrM2yUdRHB3X9WgWyutY/58TZlBu5REnV
kDQvlNJB/lSKZitCp4fqBZdPgVjn8rIZLIhGmvazAjhibv8T/na/TbjHVdGV50CRGG1Pmxwlq1WS
6e7YJ3TMLWaOel8ncLu0BQ7diaiAG6obK5IOBn6gWXH4psWBkJODSLL3TE7afgbxWPBxFzotWdsC
lHFvbA8iJq9bsRaQJEJ57CFh0bFrnw8b0vvHUq7bdNXHr/jEjvl4Z8GPOsll/zQ6WAelL5o+iqBi
/SZ7AmXw3CuYBex8JYWLDKaqWLRqFGuWMhBP7tFs/D5TGwoC6g9zahbnEcFlQNB5OrryFWxs+5qk
EDZIlnwhXZ9jdv9Ju+3qYD+6V9TUg3G02syaHZJlgpj8cNRCqhufjcoM3cevPxXH9bLCQCLNwkus
mUWsjqriDNW+kz5FO3asABCQeXJ8eCROxnhtFwGnv8db4Ls3GmbYPQTJrL1G5BTY52k9btM8/ckz
F2doy+AWFH3/x3fR68T67g9SnAroQG4sKyI2dJOm231+AH3WQMB9XzHzJcqBAbbj98Gw6An7VSSI
r04J5ZvOKSKoYinh5KJeWtsxY+3WUr+4S4N57kmDwXaHjr0WgTUqy6uU/rwgTiu4TrhbCfYL0+Iz
JkcFDMHJvE/kLAFdSrQG5UutPaSKRcNN9xZYPAFoShpevL6WGuZNdKhSNvJ3PQVlBCXZxF0E0kyz
B5mCJhoQTMvwnPijnv0z+tt9DjGevT5VMmYGhJYnegs1kCHXBzikXGfdmPfHw69K+tnt+8mElkEI
T3DIGMZt5oehC2dhg/wQMOP2C2SNoGIFMJZR5N4wP+DgFa4Ep3BtxxV+HMGIHlL2W59HbAGXT4wN
ye78lwmMuYo/FQRV3xv5va2ArIrmJgbTaGTKq3jGram5r2L7cntIh3dF93yjlL639ntp2XEBT68F
V+a+Wexjbe+gdHq+t3XMU3Ljboy9ku/vYOheSQF5T6JyYcHxuiOUwNjYpDdoZQ5W9D2UT0zjrO+3
HshRFFZur+7A+sGqQk3bfFJQ1mki9XpApjcNm0LhH3ldEatNBUwDgUc0Q5NzU1Tr9PpeubFjIEGQ
+AMLfm4LicBYI03G2vXhLFr3IEkeVWOy7HpFOwsrQDcXUo10siTHlPLnASu9tT5RxrkRimmggsMC
t6l90LVD7PCqDnscEljTE88umi3xPGC3gdBXmM37tAVY0LaNQ4YB1zTs/nV5iAlSSIbKu3jL8eqF
q6Ds870Ot1oBQQMu3YL8bD8pXOOZkAdMyyUKjDQzImixKp4n1/mFlAabeCOZLda6FzrzfyYd20Sl
sTGf25abQ4NM5WEgwK1dBbobUgERgGBe/A02TYaNv2bm3jVe7j89Gb2xlBPkw44wfK9JgwNzuzJj
1YMbH4b7kqWxj3UOP6EPLt3kqfxVeItI1fDNipU8GOU7+ATfsGsfPeZpGvdL0iLuWX/Ij/yHGH+2
A+GIsUDdhQ0JhtnSOXhsnMzbMa1vbXC/cUjQlchqUVq38NZLp4+0RpYY7QhqlFCY6BZ7/ALqdYox
aQSu9i8sST7EjRIOr6c5/gICw+kDdRJAWtkaGz0gZe3tj9Se9LPXMo/vSPBw5Jiw3IMqnsNsicc2
gQ6xaXcK3lQcP5rUD+ukck7s19hOnuQIAe1EjvczutfIaL2xerCtrGcNPuu7UXVzShsyNPECHhMX
FF21oKWUexIO3LDxd4RPmDa2WZw+rgtv1vCm461Lr+PnlLm0IkGvyL5m0kQM3MHUyWwfUqAGZYHj
cXQNZ5enaLhCTErAELphIuEIIS/t7YJRiObeaXRfr/nztS4vNb2ON3J0to6stiGXfUQTKyi4/LGO
n4Jj4CMPG/o4ylj7oW8vUW/wbXxTO9ECS4rq7ETXTMtnUe2wtJd0LxR5FvD3+/md8FC5te3G64mo
oD/Z1XEK9ZuFJZgp+45a06Eouj5BB8exWXyVs3LJVfKYw0xXD72qXAiSGqbwJj4cQu7aGE/1WMnL
asq3wnpa3o1AN/N6G6NO012GVTzabEMFTGCxTUtJxHTEOa+DVp6NXgmT/4Vme0uXTtjeyUVSdwPB
zWEW6I5gW7E4/NCVjf7HCC2j9oqXe7q3d3rkhkk0ogDxBYqe9sN7dQydvLqGgmnPFXVHu+k0LZ9+
MGW6+VEeD18Dq0qH0qEsVUVqcztpalM7YTMRo2d7kymADL0JHNd9BS+kBhECaIqHjn76USCgZLIT
w24z480iRLL1fgtcGOsOqn99JJ0o3pVNySOg6BA9zoJsbUI1bKut+qAhtH7uvmnCZWqLUa+Ly791
0XjwSsodyhDp1FgoVRfy4hlsKHO0n15GQYsUTaooj2eyVbn1qMvxWb6JRqONLPNHoi8Fc1F2qSW6
sm+HuXg8GfNVyLfmk698CnW/lwRy8s8eeehLhFOJImVcjN+gNm2a4nvAvNfytVEGLlwv+SQFOck0
sMbzoZkbWJhGdAoLMdMABA0C58LWiIjDvg1mOHhdeRzTlP7s+vbqLL1M7FRJHTEH/nDAqQrysY30
xTw17XdAgav/drV2TBRSdZUgg/Hz2aRaLJuv8i8T5IslG/XEUiX2UfxVnMKVVgFeo0XdQMyLRA/n
IPQYoe16XUuJVLBaAWmHgagoJI21e0R29TvfZyPJozDpj9xcTroN2BMBq+37wPYemgJt73GSN92k
uG5I3qwHceOfJrCuH/GlBmwHZMVmKxn7sth9oNFu1JcLoPJSnCmUDMFAZ0CDQhRn5hN1O5gcjBEJ
3s9QC9//K8mKYojRue6SffpU3+jxKp9Nci+8MdeQSQpRWi71CPdyJm+JDXistWn7eU3E78wXnZiv
2w7XifDsuqTF/76kULgR9URQKJE9jxuT2k13ONzXotK/lxauxa1TQDiwjB3zGr//EK5c81epa6CK
Poj3CG87qa5VLiXPPFUFA3zb9Zqoi4LGRQCxs3VIOa9s
`protect end_protected
