--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
PLdWelVQ9YErfAm0xiFg1EZxTrl7uSxvGnoWEm1DWWs6uWaRfRyEFWpkrHWf4nXm/Ds9mI2zWHEc
5ii2U9dPzBU/BtK/KwDI+DyZPXPQngjh/0MBPVAdEHPSfFiUd/t4SbyPmB4nUbHM2rkp1Y9ghycB
wjEVDWaoXw+gkc2s1310gJDWxAgVXrB5eTMOdI0c8fjpsYXRdCVwfCIPqS66KaczCnSVk44Ph7sj
2uBHAVc3SOXThxVHptllFOBCL4DIC3YdMd7JSYRU6ePePhMpup0Fbvebm6jXcGJ2GyuKwPOXL9MI
oe6ghDC+qNWDyJXa2DjY3hE1jjm6SydC4eEuEg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="5OSP+nwngzAOHuheMZkMAyT2vjterGqqLnDyv3zd2t4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
kLvBg389HBZmBLDAbq56NeDAzu4h9RNTUPoDYiZTAFAj2QIXyC8NggqVO03HiC5mXPGQj2UA7RHS
/uJ74ygIQ3eEsBytWBJUCHR/kmtSdxJ4fXdM2HWwSRaOZvezjxynCiqb8ylScOgACg/K3In9/jBS
SywT5ENPwOTi3j8wppaJbwSdy0F0RPqS5Fz/72tYZFgcwwrgw//stnG3ZX/5oCR/pna7MT4WJitU
qA0GDObzUHXgGYcw/YGQmKzdBVuFXd1uPPhwAtBbnBmxscfl/x63lh5hrc+Pykzwwbli8zZ2oOWX
skMQl5ANrqkhzHA9BL2c5gaVkuzd5TmIWVSwKg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="m71wh0hOHs/47Tvcfbdx42GP5l3DVDej4j5ngpRqJNw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34720)
`protect data_block
mIHQmoV1p/L6Ziy4UFsd6+153jAu520uOVDEeMGek93IwGwoZUd7gLNy//PXXl1xO967RoZyL5Cl
+YZfnTuxeAZUh9VuA5w3p6trr0wFKqpP5T0Wf3dNPkq62VcX54WNMFGoqYgtGgk+rK572BIG0KWy
RCJMBYrRQN8WrJUVtJh66JGtN/WCtsAJSvLQEbekuUduRVzLa82w8p+80eqOJdCAx4mknQVw+dqZ
Ij+rVqkGV/T9sIrUe3pa4MVulN8ok2vYj7FgKBXwWE3V9yxsD3s6dblyqblxxYjqaywoXwbD2elT
NxApgx+cAUxtphENKgnsl1iNMEXmswGzJC88hogxTC4o3oQudwwhj0xcNrcMyEXkzUjmCcMxyeIw
xeGsDeeJAKrNRcdg1TsVWG2zIMC+Dc/ZW/oGlAI6IsEdcqsEUq8elOBVoS64fI+nheqOltVHGeX5
bq5qP8R0UvRUFRGVc568cgNI7Fci3/ZaXZhXzOHzgtrCm1Ypd15HVU+IOXN8tv/fL0Ozp5uQBzy1
k9wXh2O6hsObVqTikReFb5cYX9Ifo87ozLRZNjDoP+8/aYoMMJU/6t5nEklxD1oy6Umd3Zq4lH+v
jniJ+shmMpEMoeKd4EyOWzACQ+I2EzJix61eqk8MADcYH9eCv9lbwktTy9SwndVxu5gbfJ5P6XIR
wPtjbFifaBgQsKJV8oZiPFCRL+xG5U5IuEVDNShCFfC52/3V+HHKZSf6fO0ZHHCrmGFzOcf1ucnK
PdnmFcglnoTfUJQ1dPe/ETLTLTw0xwyLdp3dmLrMj+3A4BlR6z3TyxaKsgkRxXEOGMgldZy0bU4M
EQ8nqizXIKcRFvuzAEOTfQW2jsEU842udhLqA6/OibubvubxOUseK8w5Upp6riyufIy8oQn3MEck
yk5clDNd5kuIJ6MzL31mes+C0seTT34TmPLo65APuXXuJNNOfDX2+miuPcUeHTRSYH7iyaI4M94N
a9FiqXUiwoe1DqHAjKvl18/gtiKL5b+M8xf+I9cJYyfQ1AUXRLmgmmbx7ofiOhfOKc/1wFsK4/SL
T7GVSZfAxOIks+jRViVmC7NHA4IQ/GwgyX5eD2LSqTDHV7I0EiD54eQxneKrKm/PN6n7jP/BSEpS
UE79FbrEA6RUTE3+ZrT11ZolvS/xURWhRzP1RsAX08tUZlRrgOQdH19GNnoiB6W/M8p8Co1+ad23
6YIQ6rsP7cTO++QM1nzn+ziGWCjlD43ZJshVM/dKJOJ5pbAGSLLDEKlZQeW8sbKSUXrwE5Dm6Oui
4ApJCptPWQTX0DQiJnE9CWvyUtfstOJmXcYg9nD6hre50/SlGzj/oTfWlUsNsRvc/PDYFZI586+S
kG2/vmoIbALHS0f7Ra+KliMKwuPepKeIMaI32jAHVZjsKy4hcnOF82LP5uWJR3nv9IWcK8pjgNGT
RenQ8g0vJ4kfzRvu9enE5h8+Cu8PqUAqAyDdj1d+n2NGWNSOkKmxRF60eP/V/sjkPLy0PXbg12n4
UgNeorje5Lr6IBl8Zm9Lv1ST4r4qXKA0el+bE/7Q4zf+qb6xx0Rbau7Q+7V37mksf8Zy0l/hNWn3
Oahoe3Ige3AVsy6xE6Lp1DyTCZhwcGUQoRXTz6B0H6lLWF1gEwuxg2Y3NPVhR63bzANh15GrHGt1
ESUwCneUOHPA3tKpJVfhilAmHBu6Y994HdqSBC8rq0y5vaynz56U8nQwUoBUDtvA24JXAQoaLn/w
LTIa8/hzdDoMLJzqJJulhzT2svsQGOYjXvwAXfFii/SgddPixh0NNeYUlkpu/z7csSaJ7eXETmND
FEfxn5wA7WeQgoo5AaAOI4jIxQ9IMDNDFw9ZngLoCrdLSjGhTJeq4vBZKZKrLoyZIog+iUxE2j2/
G+ZyAmiNmecXqRBtx+p9fED0LqfjWBifWpz5MQDYK9mVZUxqw3XQ6kKkvqacwTefsB/G5F4ITGOH
DQfMz6WarG+HLJo3GCFibwXe8HmLI4H54tn8W+vnIkY0hlBesNHN9pd9B4/B1/yaGU0XeVH1aUly
jCFbx/He5GVLgvqJbI0CR5BFYU96AyLonxSXdGDUn45VfeOaoY4kbXCmijz5nr4Z8neLBw3XEP3n
FeSJbixZqKDfCvQfhfl27aWMV9f3caOJOm9ta10Lj8r1tPa+B25iuxjEv44fQBrNCRO8LFpUX/yy
md5sVLEJ0HtJPcfF7WriMwBCZRfV56mphAYIKBV4RI6ehRcrEVv/HCRt4LD39e3DZfKnkqc0zsgA
PEfe85T2xnYfam9BwSvADjKICsMlza7EHghY04CyFMcmj8eSdIFZdINZeVLGZ/Pyt3JMB2NlCdpf
7yL2V7BGsKV0lQ7AqE8lpb9iKcOii6MRnJFs24lBI/rsSNUH7hGMlXi05ykQYu+pZqr/lirCPo6K
vfTtWNz7wpFCI4jaxXBOxbpWi/h+Crge13WOFF96o9ZX9902w9e3QljUTN2oHv/N2fgCCkZSFTEk
OMAnVboEEGMf5PuU+zfZrzviOjjl36apSubyN3M0SxevdEW8p2U1roiqQdhb9zBeRuvWqtW9WjZJ
1OTVM9PDR7KJYh6DBM4DrR3MuFGURc/ty0+I27fJ/UC5p5ovu4L4oMN9AXtwDH6BTQ6SF/xNuagK
V7vxNSNnqYk2U04s9lqqUG0eOvb1SwOKNxzz71ex4Lkn9Gsz1KgI+ZITYiQjhhT+aNOdF6T1CtQU
atlBecSnSATp9TskFvx8jCOCetww58MABTU3HIEEJDYo/DLsKShgeRC9L5H7RptyzKRLRE7NYi7b
DSkBKMi5LjGbmVYZmxjxdU7BPL9b55gdap3rnnXPiz/pJX/hmKpEbw5SH9C6zw+7gFBOS7Ntth4H
cRYJxSpYXEuuknyY48pezEJHNq5zknNy/Qo3UGWgQaCKBKtE4K3G4gwpqqJMjAavtNE85JF7jpVS
afvpsUFp1ZNJiCk+5ws3jLo/o9LZsEkXrhsXuRGL7iwrsNObeePy97jKDKRKj+G/mv0e1JOFw+o6
LWB5Xh0ep1G3LQUCOtNH30BYTse+fy7hVN/nb60HzwWQoeD71/3rZCsKUscyafymMkl76E1gwpJ5
7727jVHrAqwWoG9e2NBFXksSk0u+Dikt91dIlTECpY3Ena7+aGcaPf+Dz2PmsdcZBMRbFVbkY/o9
jOD+PY3DD5QDBDasdkONy9izAgh8t5MIylaDk5thmSvIiWtxvnsnNm3/H5obifg6E6sjwhD6+OsB
yFrjWLWeHHGulVQS8PRuLHa2yIdchR84NGOBXq/RNF6jdniqnlLQGsKkvYIvC9y+SJ66yENDSGYD
NiREZChXaMcJjnab7ScRgv7gVMJgAgwRHdx3K2S8mbWdV9E9k+k11gR+kfQPp9e8sd6dgZGHa4Oa
i+hqlXzbLySSdyMLG+qPcUfikS4nkw52K0Ug6DLgazyoTzpirKj4QO2kKfhm9X7eYKwYsAuSM2na
ZNBZaPZfAa0xdK04SkekcxCC/sSHTxK7IQP7odKDjvoNLYl97gPZaMuzp4AYEkICEc8X9X/rY7cJ
IxcKQJyOoqwtA4HaHplDB4D/PlJDFXnrUqJ1rtyx7ZNAcHWK2ZdFIQaoboM62NmxwiCOffnkOlyI
tJIpQA3n0JnV437mDDux0DrL9reunUYzqTlLausXFVrf7etdK84tJflRsgGnesOQ1JpzIdyjksJW
9o0nM+6n7eV8ajsiGIFuEgqXofhgtzyO5amcVKeU9+XNvlmLrWjAU0YSwAy3/mQKPnh3wkq4XEcT
GXSfGD+5LsAlNqxul9LLEMtHt0YO3I/16jDXt6WlfMaOWDQn6bMRAPFyfZj92qickZBTVyLA5QFH
fQsAyPRpZbU7hE1DFK5hUmqjq7RBsfxrB4v5e4UWT5lVTbJG01P562luUtVvWuJXsit4FYkYNNSm
NhvT7xqHR0lUZh1GMfOZzxu52ClC0/ftTt/kyh2DMNTOONTE4XXOSugmwn7nf83TGIJDt/w7Zm6L
+eqcMVeV0QqfJ5pOV8Ubl0sMKOgLeqwNiVagQuruyLCqyBwIUzAMMfRSz9oYVS66x96NXHX8ehGk
iTiW0R/hYeLuxNr7NBaFYxmBdKGD1qpJgFJF/7JHFL4DDmo3IinIJCAKSjVXbW/ahUMdGQn8EJ0L
yciNLQ19U31A/6IxrH+/y1hxr7URm0Ki/rCS9WMoAX7wumWF3f6ZXtmOW1ajkh99rYXK6X1dg5Ws
6PCXS4ERyIvYp4LQsU1uMxfe2Ky4VQ3/m9tyy1Nf7rdRwNH5f18LnWOOyMuivxNyLkopkcImfi0p
TmUuRvt+Ot2MPr+eoGl44ROcq3EBigsccJM2wpjKQeQYYEh55Wx7w5j0Zr/ZAeX9z3OD+rmC+eTj
V0SDGLaXL9VOXzJV4Bo4lMCQusaacopaFf/wEpvRmMJf5G+mKURwazNUHt/O2c3tBd8aBEVRDOPa
VwgR5EQy7LReYV9GHjxeyQ75gAnw7Awi9lWpour8z0L3iHQxsoLVewefPA8p5W/p6gmM6Tvi5aRQ
nhMsHxXBQdc8Vfj3qYH5X9WA7Tx4fsOzm9KtMjtgrNNakLXriQoIyW+w3q+rv9mPVrYaP9Mp7V6N
LFjdRROECbVVbC2bDDDVrPRkZnRH/ZfavG2doYoMTvGf4qFxgLXsSW+JYNwRTNvB4HHLYBCodd9Z
xL+nqryiHVuNvCJoqKL/vq2ZVo+OeE+g5JY8PCeBd8PqMElj+64U1/0wkcwFbgh9Rkyjq88OKGfz
VCkZnF/GHfVBEPIGQfBzNaNMxs/cm9DdqZuI268WBLSWkoclxxOiAe8PhmgeLz8qm5olaM04Ngz5
QOWho7vN7LZlWpskUhtrw1QUnMzY5mXvaByst6vf0I1Ss+/9Nr2AO1qLcBYGI1ryRLUhP37ZS0W8
usFQfsmuTO15jiiIdMZG68iL+f5aUp9tdTTzhnXvT5pqiyGDhlH9bA+LuVOaEWiU8q98Q840Xd2F
3aD5eyJwvc6kpxN8qjKY7rughEWXMsD6WbB8YE9lrIW1mxt+UNO/8evaCYo+gBgQhdbZyFcepFzs
LI7HQmtMFGL2Xo/iSe541Xo/Zn0gvIIxwXK3p7r83TDETPsSPSl8rNolNgxbaljiHx/MZAkc+m07
tUUKB85G+Ugk08cUXf21wr55PI46IZsiBGER9ECcSbj2ZmGn0SDwA0jbVuHeJ9vNpzmVkBPtGOKw
wOOqrbC8VsIc/kuWvg7NXWwvDGzmsETyOn8vSHZZIwujZWoqhJuIvqpJ7WeiKQR9op6hzTK9WydD
0bfvBWrHbik6sTRUmJw/951Qr/t+ciyUhIoCldiK1eS67u+T6E1udlgIijqR1t5yYvzVXV1JcXYr
JBHFAPqGuDVl86mewcrmufqghJT//eupPh5KdwJs7KYDkYam0TCufdvCBfssY21Zm9lNk/bBwPiW
kjE0H+JIbiwJCHdzxzyjWtU+qOjJ2DYLFonFP2TyQHbJKcoM5fjVB/r8yNk3pFrru45ZPHBgnR06
UhR+Mo8tNclG6ywuoLF/4S/6KVLgxfrs+yuPzkBssLgw2Gpgu0ll2oP6w05xmCzdwxqAtISu2TU6
KCXWQ8XXa0QaCt4zrnYE03wFxtH9dThweBSgPUu/mof3iw8zvkc+Tr1LZIFwz07nhdFfv5vfpBsc
MwZG6nPZmMs3zfhcRglg1CQ57QIS3vVzlbAkXL+SMJIzv2PpuW8uxyIf55Xx6eAkyo5NrK0ABNoC
7Tztr1zOfGroFn3Hn/maYw2u293Yo14vSxBRParum0M33RPcfapQj7KEtaPX7HzXjnEO+/l0zPTs
tfSe6KAyNipcE45OxVMMYCv7OXG9sKvVG9d1DqBA1IGKJUeGmHv8aUiCJscClnaN1JPpCTtylpLS
nlY4AiHqsXJ2/qdZkYGAdg4LFKfwRfcZR4qinQQdBoRoXgluCgmf5L5F6TnpQ/RuAs5Z3FC8jOp/
yYxi2k0Wd5C/ZXmOmJPTTif9T9QkXTL6LuzTY5+xOQ+T4rG3pcVZV9QdueHQugIB5sqgrg21UdO+
rOf07CZIT3yPbeOEE8jrt4p5kcvaeUVEBIywMo+WOuCvdAddlWnenvXdXXw8mtHgycG5w8y8TaiJ
s1OGhy4oX0e7fK5DoL7rb/bZSOyAR3ytu+tym2F/9eYiQt/nGolXU4zw9WAx1T5fFHiMw7hv0Nth
3j7fpYfQS87z1RZgRLJZlhRPWYuNqGoRaUNqUzrvbua4Rbg5TEu44g2+Bo+O9x3a3NGGCsgv2tI5
2kcnsT02Dhny1cMUWqKTlxTXiZfK8BNjOb18y5yVsOVUjoJyAX2dixSwBmqrXMrcjyqBgxyXWZ7Z
bGJ3R1beH8tV8P4AEux5n6szXBoAX3Ale5lFgIeyLvfyEBxdXoxfEKvuEhqQBdSfvKcaj2C8bSBJ
jw86uouhSC3eTYU/SPNoOVRL0QfQKkkuRWFkwmFmSrpZNDKVBrKifofeEdPgfgm62PrQECKf4q0n
4uawBQ6/SbBdAF9qE7fOtgIGjc1zZZyGorWkeLtB0BeqBhNTpKpboWsTGgA0eqgw6Qd3Pv6+91zQ
7acOcMnQA8OHsQKRT0Uis+Duo4G3jcLDbdfShoaQZ2eFa4xpaW2GkUytlGJytnToapi1ZpYD73bG
kc7u7QbPu5XM48MWsGNbxqZGfHE1JnIp0ufGhq7eSHzB5Bll+eq3Qg3qaxxFAZWnC+besxoiEW8V
F0VZdzY8QTi4YeDXsVulOVnErIip/HT4nDpBk9+I75cUcRmdgaw47IljhSj9yebBIrja9pFw/ZzB
IvLg2zE6U1QVXNwAcGZ5NU8V5RQMp4K/X1w+n5TyIlkIO8xHpvc7X9/gWPui1MnFS9ktJNUO3j1X
WjMZoPVFuIhJnHGYRS+TLPvzHyb/rZBjTq9qaNZrr+U5wvo1Z8eOe+UZB9C+7LEirSN/vFZ1yizT
aE3N6VPw7vKc0lX6ihCKeoazukGanPKfS4cEHE6FxqDDQBYUXDn++GsXnAgcm2uJjMEzlqPtWDYq
1OuH5db4hQ85xN13/+Ih8pV1dYbLDn1t2+K35CPV4UwTAaXSlhrl6lUmFSbca5UsTeyN+2xNRGRA
sLEXv4/wFCcehokorRGWw3IqUwIwQdzF55s0pr/NwmkmYkPG7XOSa5HVSpBs9pA07z5/s5fT8TSM
sPS0QdKCVUivB7zvwolQ4mFHNKurwTJJuQ0okiVFDPZjtwD50atrxkYQs/NNSG6DAd+/0jsyUV03
+b+Daa1slMMr/jLVCW2HPbnMmFKkfAkLMZc1OizF403moGU0IXt6nywRpiWpE1UmAmfleuYZaILe
AsFW6VF1cKqHUcCa2uT9nSlWWju5FkVXWiL1ZVhPBYXtxUn92SHVUP4+vlfEb7/sXTb2OsYXquYD
scVtY4sn88SalXn1sb31ik/2BuKr8SM0aa0Rw4jZwpK5pc9b4gpsMmw84Gdg22nSW++Z+attqyKQ
4nOzyr78tAeM58Mr4y9O4/hVrhQ6Feji+R64s+mr+X7amDfGAwt1jUFsiQpPg790T5M6ovLrzi4s
BN8jVZ/6GL/xJH6CRP4TdplCY661uR5ttRd1LPyF/gvPbbvRNjNoTy6HbSvcgt/SVBUXsEsFuXW4
ao5FMDwUBgOSTrUEEhuJ6PSQ4smmTiIguUZWsmUeMaL2Rr5etun0DvOcrINIxiOMjBhH8apbgPr8
zwObKDphTzWdauXhLIqCjBgX8BZFK2HTUZfwLdqQ9bkTyaUwlOk8z1U12b84hkIXZ1DPDSz+BYBc
GIEsWgqFQIk7hExBDX0+MbSkVneBCa9dGobd+aX4o4Bjas9rMs0IVAU24mskTvA5nGN8MHamJXSn
esIRsbLdOQgulkhVKAqAcr+qAS/CSGiOF5KSX6LRke/d/xMxgQCSaNUPB2Co3YDcyB/0lo+5WCpy
P5w2OuljX1SRY2PPtqbPKviZk42FIZqDAHgOzuhO2eD45BBwbzL/SulMpQYFC0E13S7WW5/s5Otc
QUEFdlfzyW06eGVcdcmBRx1CBHZYf5R/YSBXATIRln0/KlpzTxlD0FMOWeRxYktOm9Iq39xq0+vq
dPhs7mT7Q7w2ruOZdETFoQ0xjGEi/T5sXuDfxboqty77wX9KxsBvuTAWF071mquhzh0U06kRpjT7
66otjanPy0qLF4QkCgEhhjNQqqhDhRn6wer00PVIfXFBH6lZ0YffyBvSEv68AfjEOEXrQJWlYOoj
9qwSHA/cGo5ahfsdygCTmxuwRQjj7Z47r+3UVnD5GF9slXBwSQYiFHvgDl6nLAl6Of73IQGfpS9I
rsoRsX/b7T87ZHDojEPnjGstxtUW2aHJowZ27ArnXIhRLNQrs9+VmxFmV0a8bmUEUzVgzEeH3zyP
SZ/Cp2uM9XII5ztSKNwanOpNCkF7/xGTsBw/D/jcBXkiaomkCKjwDZf6foj8aCOQoo4cLRWXxtMP
odS3Zq+WveOljfpoCVsS7EGTkpNiRenHUZ8zny6E9SF6YZRdoBFQQa2+agtPaOcEgov3q9xpBJGh
QD3OKIPsB3D/sFempb2NRs+X9AHcMSmTf0d/dPhfMSopIOgxs6LvtRXSm9asldpJqbHhxe7lD7wO
MtMdOyqN5FHwmVgwhZewkZXNx+QAmOojExB23iHx2gEXba+r+td8N//BJk2LPMo66RX9KphDSejE
l8tsrpea8r/AzmsyStKnoQ8wIN7lcTPUcQjo6hEUvscRldtSHguZzATU30oGdeBuPotFN6Ck66Lr
yd9KMjQUEAEQvGqs1orRvikw9ssfj0Nx9pYpQEOuoY0sWhA64sKI7IYSBygUDxn9M8vGgRjBM//U
VQdVx/MXtqM5O7sZ8zeC0BapOmlVyZholOAu/IyUlsMrNaBGCRc5eMSqtPy8OXxVRkrQxAQJYXXd
QCH52ZgLVMcPmrpd+gfu9EIb0IBtWE69g5c4EMDxSdFq4+RX1CVhUG0dFBz1Ei65chDl2CDJBIYS
Rw64Qn0wjb2AiocL8z2PFev2BWoToGiicpBhVDrh7oYB0WC7MgYXN4i4zUm9LvAlTCy+1gXPS12n
0I5ZMx5Krfwgru5g+NSbJfRVtW4oq+euWW4fMygF5B7K8X4LXAN4clfcofJ64NH9qmkzDuA4Okgk
6lCmUoljDR/RW8ZkejJ5l5xwjPVdrRpDZrz+79zsVMDBzY1azgion0WYSzUbiIkfaDpvwNWhTONm
VSb2QSjT7v710bOfr0ah8JG/ZXliF6u9E9lCrBlbx2rYEmB/Cz6AG+WVW2BK6NQGMP5QxOX+5rKD
paw8Ynq2htyRB5Hpu9rJcJI97TNgGs6Mon59CP+p9ZBQaRxVI0YlArCRfSBZO+bF0cYS8dCsdZ6w
WxGtYiwnFKeNi5eYtpBvPqI7+zfMdhgv927ZWGbZGR/bK2iVHxAX+9rG0VAYgejzdqisxaRw1otd
D0ty7Qejh0a/dPQhgUCzRZbYoaXOaHo1yKAEy85LnqNQEB0QB7wBrlfXL5ZhtXaUwEC0EffUodGV
TsHegQ8AVhBUmvMsBShja+0GNnqHVuwOIPMofa6v+OJlvvpsv2fOEAm2B/YUcBJOshgIqUwfUCEI
IdMdrZf87H4FQxBqhQPdsKmDUgD7Lt1wDse8quBpPr+NLR26+gMHaV162XgN+wDM1fnLOnslAcIw
X9P1NB1dRUPXeTWkAJY95OknxJtUcrXdGUG9e0Sh7kxiy/QWVTv/E12UcSiC0Gr6BAmpMW/0hz1T
lmcUa81g2mn/dQHtUk9FzokcDLBJ0q/nRnQ1bOlmOTOShEb2V+/MyQS4WsWL6KZO1/ebsBFLoZSB
C3djT5t1py3CVOiVBBGeKP7zpx3gyYJaJrFBb0aPqBn+rL/c+ltPePzpYoWWsIrB4zOdIMNHcbDb
i5tSD7pv32bkxwAClLkVAbz1T/YdWPQoLgqn7dVLOdbcT4f/sLSGV7sb1JdGwOGh4RpEv6TDGE0U
WXVGHMcTdRo0LpxYAvkvoYUO/2FTNeX8l15ZO5ZZoiGwKALmrYR+NQ4Tm7APeCiahTz0nz5lcA85
SK9pE7AO9mN3cwhXoybGqT7xkc7gPRLOqcS83bVqMJjuU/lAUyTzRbLcHNFRmJAWeRqP2XMzgVk8
mkqPRTxqCjzh8V/HDDy3jxnWL8OfwjQI/BWK4IcYeE2oNaRFZ3F5DVBhwcJPTpgtX7iohwqADzuT
X5Jh8ROlzIGvuFhZFKuCFNve6tM2a3DaDUHbkg+7zqnA0qzysg6o7YcONv++eXuJjJ2q9sSlYOAr
x4gMs/30ZcFpY3CPYcMUi1AvRjstRRUW94Uxddla6kjDfxBtMvNvu3DR5n4GLhBTv93ojcASabYb
sFXRd9S5tGtq2AT3VyzNo8w3i/39ooDwscg8q3t26Ck9zbrElzYtHgzw8/V91w0mkjd9eQJ7mZdG
+Yj8OeuRqRHOjciyUgSZLgT8rTnPuz7IsMZj6hd4BneqUygMP0XWgTsTkXfzy7RnvFqbrvWZFJwC
nWAOZYxNke7UNIA1qhFNIpS0Jo6YPk6CqLPLnrnC4Zq4Rg6/CYhG65SzCMTIXun2ECg+Qn8s3E7x
gtMWUR+G2U03ajo2r9GOmH5bwbpjUWm2p5dMelB02XFDCYFAe+VYgs5grcwDAAudJrX5Z0U+NcqY
R8teYXytS5cEDZDD+cw3UuigWxPidWwKltx6fvgbJlcsuccZ1RfQxniy4NmVK8vblhfFI8fR1zvQ
9gsoo1c4NXOzgo7WD84GWoTwDz/mV+do/hoyfijuTSl0dOFKfRasuhHLKUFi5SO1JhLrisxVK4zS
qQtXdjtJbBFfJBdrW3Ak1nU7nk8uJtNjJFQGVK8KzAa+6uITcfgMZ9lrBBa2IE+JOQfm0kuBR8jw
sB0AzonN8Cq37mVbQ6os20oMB1vrd8/+bqqSgr6G7kqzaV5B4MiLKcNTId2rb6M9V+hckeb+Ulhu
9rA+zj3OmalL3ABvR9d66u1wK+InmeIWJt0X4qN9bfHxuobvaS3SoC+AoAOtZt8tmCRiFVDMzEr0
2VvVGvot7Q5e98RRUHTbR60WHANQy/PEKdV51cfE/88lC4eLUU8KinncnNQ6B61I60IpHx0DBaN0
jaU905K09Jew0C4ND0p4+TRoz2YAhzuAxyR0N+SEmi2f9s/zfCvB39f6qd1W/gRvFWA2qLRWdZyo
VgLn71bZq1pNi0i0YnUL6Ycg6TJ2NvQhPjQH2tPhHDE/t3/GjItfArGiohw9tX5Wuo2L1e4sw0fB
GX3Z8XTUgoNp8AdffbyuGHLpMYsgLByeyQIt6SDFSzPPtmiMqC/QbjzqhxyyAlwCkPuL6Z88UFgj
pyOIaLCNzD/qbjWl2EDuqYnkoxQp/sgAfI0uzLQfpP8DCyHI48IoqwCW8cEKmWbi7bxRoMGoAmBl
ofMP56wowSj8jakM0N/eUptreGkUcMa/ws3em0VWnE1mtzbbuhMdTXdaXL4EGe4z9w0kuW6f1lum
AWvLB0WyfL8AMT66bhLoE/nftZMSaOnjW6qCy+pO92J6p5M94S1gpxncKemsakTnFr5BNYCHSsU2
UZ2id0/hSrq+oGRGRj9ZxFsB3PhZR2FStSNiUzCtf/N08TLLHsTNIiQu3A5RMscODzTbzkqeHy5J
Thg3/wEF5VrHal6dVx3+UmBKNYSC0k7a8z9osbbdV1ixLHrDbK5I9os18bdrlpamyZMHmvUtpRjA
bB+mh48tbDaDJXFeN5Ar9lL0y+0GiPYiq25K/EJn08BZcK1HrmAUeILPZuinQa3Fwh5rie104lqi
TriGLzoLoUgdegkHTS7ZP6PBw5G8rcGHuHkx0tGErdMipeeVbQbcYlRijNwWFXgelLP3MOva5Zlh
dW+G9z2Qt7GDe47M0wWa6agOcw7RNfaYpOFMojpYjSu0IQDS6MkQlqGaSP4hBoDYZTKwZAFbShCu
NwShcqST7Ex09wFmgcu2av+55PNE5kY7cDascOaSX0M3+t3ot7rSXgJ5PlafSgIIqFgmQ9uj7xPN
ZVLVmGdCjhVfCF+pTOtItX7CfqJFD1FN6qb8wiDttQTOUmqPcYpTrelqFtHCgQina9tws7zbpiwn
GwvcQlLGw1XraqtkNL2SPNWz5FsIOlVYbj7xfq2IgTO2+06TpW1YOUsNBqn6axXjYuxiHrqhLweQ
ROlUikWM5gVcun4H0rYAc7IPwnBs3igaXxtW9IphAp0QRUKyb2Uz2moYznOvd+NTd+kDW8ldj14E
jcDiNHKyXRjeDDqCDR2slVeTqAjbCpb1Dq6ErPsa8hW4FXsfkXtMAIdpo5FMp+V6Vgb2RRhNbUny
gugYOteiwk6cr6jaRFV4O6yCboGmIMaEJYVExbkL8AeUx4a0L1BNLsXgf4EgoJmK60yA2ifnFx0H
itwW2rdWilvMpP4zR4i6Fun5plwo/ZdkzdlRJCEoLtzk/o5XEP5SZfYS43JJcotTyVH5T2RpTU8H
1rfOa9mxzmUlM5prSVKSiw+845Z05ExzyN0cNU6vBiml5YVhc4OldIGIEMc0kSPa6YJudzytmPC3
6kaTjcAsNyJvy397GaRrQIZZN78Ds2E1/2tzgglyfQznS2ypQdVjY60LPW7nhrwlfZmm0Pypi2ZU
2D7TwZejKEdaJOqNuJhHsWbvqqBK7UKxhop3mj4K92Lu5q5SmwXyvg90bUlswgNULX5x8kSrsvGx
jT2i9fnC6aXS1fSAIRhWtKWTREiXZqUEqmDiuiFia2mB4Uj11YLROASr6iBeAq50Hzy9Kve7MUVU
+v6F8dVdnfzElbHK0pHnfkiicTXiGMKRwa/XZRiqfJJdamErIMum2jrSBX50sNkvTou9XoL/HxJ0
xTzOtyy7QVh9qpLSkaLVxWf36lxrDreuyzlNYz5RNXbPlGVqmBPFxn+Anp8BdoEK5wjNadVH8lOL
dxKhlYaInbY0a1MqsB4eq3sk4RpQbsAc04HytN0i5jvab/5AAbvcf+R5f3jUJynPl2qnGutpE5Up
LRGL6NA/L0vDogoaUq7A7LPTZUSgtMBT0IatIsi3kDYz9sg32GWSUMBQi5GWy8wl/d5Ma0DQZ+SL
mshnPephNVgllfHgdJ4yPPW/uTnpwvGsJM8AysAdBXprCCDySBFH0Ly2xxZy4gw96nXVsO/bS4gx
UL2fL7weP9auPnuwoNxSPxne1P3faO6UVxaU2B/zrFpB1iZ+qWuiTesi1Chelwr4VGigqK7cv7lQ
MzyhSeMWQ0wbFXEHi9cGLZEwTcSQte1JTkNsDdhv+jSMCN0Lde8m/3NEdoNblX0wrF/w2NQBNadY
3Y50av8Y9dY7V7R+fJADb4MH/66/gXo4CflAwP0kdodq/b+Fos3AzOF9oc74IvfI1TGJhZtwRrXS
xmaZpEeaf4UICxsthjPBYLNd7tJg9JyjhIPtBtcJ2LVIxHOBMQK+IF5vQlckGwuENHxkTapgWQOR
V3MJvWP7akXup8/6R3ldvZx7ddcsRMq8Z8GgsXnOGAjSgBdEzuK8JY8ghf+kKyAS6ZbUCv7sTpdp
ONIZT+gA6pkqnTgq8BDF2edyFA/Q3Bvq0Sx7EeKm0PVUz3ChplDwJxQA3zVijIK89/QKN594hc7e
1bfZB8xV3CBizHhwmL1APgWvXaakH8B3yubJeuaFwVLd9RWmTE9Uk1RoLeKstE94TBW1ZISRlJFF
xm4vOGO6Aep9AXDB2+oWZIKOX/9M8ULrj0yj9vakj0ieM+BAlwoemmU3BAVX2M2JeJTgl6Z1q7h5
deZxGUq+8zcTEpaPhMvcvBQgEESyHhkrB+MNrZxwW88uFwHEvM095EZbO8d+PcxdvjganGEUH6cb
9wdLSRc7pj220G3eo3Fo+I2txFp9Q3dyB42hxVUHUL6TA/5YvIiIF1xBDA/b81iFgRDwOA0GQalC
7TFQJBGORES7g4YP/yUky1wiF4NBkhmRHDt/gQ+J4hS0Dm+Z41DaDKCkyb2R1Ck+5wTGzRdQjlTh
m6lyDyBwSPMLFt921SEOhsWP5wMfQDrw4W2uUZoHaTMsUhd5dxI+KuESyYDXzFhqyyy++/LY5kQ+
tXAegReLnSnYfKhPYwbshYxeySkE4mMI8aCgwK76hViEBTivLpsgaPpmmsWNlxtFIYDl9Hb0Ein1
ZomR2Yec+JpRq3Rczt1MmivVRoK/u2P0Eif3LPdiRaEliV6UCJvv3Q0i1anNzlm4TcV6eqSOpP0b
zwCBJsUJ+2Yhb/LKepXLWpnIYmqmVNTI8ktP9fmEZzPjrB1cg0VNbXLfUrLoRkVUA78R3XM25rBM
KmLi7lNxoPy8rqu/O+NMDWjw/buIciqVCDi/qqjBY1pzWiqysp1cSq5tgPYOt/U1EYu9sWBJaPjk
ROAPGs6qB69/MnSZXsHPquY69atH8boXA1cvyEENB8DJvrSW6dI6CLimoNgZ7g+A+myOXXGNlGcs
lEI61mrO+KO/y7LO0k+V/BrT1U7woke6qvm5gIIA0copjy4PMq57VrMfELHhe/lOQ3EVFtopB5QB
yHooW+NqM/wnrvPy5fM3OFjt2gNBSW3Q2Fy9yyKpdzM3dlUchFiskUcXUof3u6sSHa0d7p4w33+3
ZAoJ4Y621xgBMRxqHJ6mFItCrr9fRMte8XcT7qOjUgxVO5s6TWzBVqJFHRrffTxAB/heSZcjdIT/
YwzATaqVH+Z7pO0PlEtA1MAtNN5N6Jk+uW6bG24r/+l7TZn+MoXfI5xXFyQeBws3+M12Rt6JJVG9
XLNG2F6upu6rcch3zsbzQGluKHYYACltNLsiH7hWWc2Nn6ZciTTK10pZVCbYrBOe82fBTWmlCwk/
Ewm/nlICIwJrxqggQsogEcAYHu+dZzrf6p/NJpStYubW3mC3ScUQ6LcOzTsl7aExlbB/PSzLiv4W
z1s0SgRIfRmS1QWBqDdtkb3t52KftYUWLwRTfdL213UanfAeNNZ+iz8J19yyos8mMd9zoCmfyoC7
hbCqjQBEgNEwuzW04VgNhSrQ4baEdu+3CZJXvNICfUHBtEojNaV7l2KnP9XMR9UVocQLOZWZx/aS
uaetKalXYlJCvweFQsb9WEceplvS3fmcLw17iIQ/Zbpr/2tdquMhUroSQrUTTIUK7gh92YYqZBnX
xPpciDI763G23OjKrCJgX5oFUBcmsqhceyXp1bZil1cwxdwDw/x+UX8pUsb2kKiGLB/3tO4HoR5e
1ndb9NuwTe/fqkjYyWqworv1EJNMAR2+2cJcgYfw6A5Y6Sc5IHjFrgxT8Lf3Hl1dmMWazOkcN/bE
NU8+Tu3qMrhHQswPGoVdB/zUoEfEKHXhtVSfRbD8YWbKq260dN6i+I4HShKuXVVXXMuln23F72tr
tlKE7onuf+Z7fu3vvcLFIQ6jtJAg91gYu4N795gGy91L5KSMk+Cugo1dgOOEEhkAskMvDyMICclH
pKasNp02kMmeDS+MP/L10/whUSxfg0tcwwCQ8gT5Bw4MHYILkauhgpAIko4Vfi9Aum3V+UsAtrjv
r95+4+qm6fgw4iLupWXmsTz44W5q41p/axqn64WY7WXAe9ZL5Ao2hn47vYC9igZdADn6pBVZO2rH
jz6LYvB+MGyPdxFUlYOLbCKPgrZyzzKu+Nwbyuxqh0nzQL9F3VL5xYMjN+KwfhiFtXg7UfLHpD+d
PMmRrG2Bw1wSrBJFxiWn/d6Ggw51eGcepRsomMYdbcMJ+0MCDGE5RyxaNCOWX7b1mt1XCPYIhsOU
dv/dLEmkaFHtbdZ0hneDVu9t/SKmHUbWDqFhf7tWMwYhD7bB+aUprz9lDaOC4PRyWxQS0mpKyx2c
dRNzSI+95Fug+LtifDUYcJgnU0w7qmncs0A692XPcK8/fJDzq7NVwIUdDpJxY+V1ZNmZMfEtLhnO
+6HNof43UgqMGkCV4XrbHwkkKBCgOkYq39dZb60lK3LgEYRNTdL260CbuhMHiaFmyMQJ/NKM+Zfn
Xg4AelSjCiwNvBUNBkRceON64zTCh8ie/ygFyhf9+LVYAaZScz8shL8cxg6+r+bZr0AIEW7BHh49
7ddz6ATp0FKGE1AYNW/uUWujzHvkUz7dN60RF2eZVEPeqZIgfB1/wXlfx6wXklrRvTAooDY3+VRn
22cNUPv5iO+hmh+wL29duf7iHF7x9mBSUNLxS62F7ZwDQq4JwYD+tzSylfVpOScOejOIXZGIb2Jy
RHgkS0Ck/57miNne4NGvZWGcA6rhtxCt2keRMJKARHXCvVMSCDD2w9qVwpKSMcIjuT2JsqJJS3Mc
eDgq75M67ayeQF+z4asEMe0sk0rzSYIVBznV9VqVCTazpAZlLWEWlREmZ3J63cxuMBb/lsGkCUFW
Ii4wLKCq3l8d8yAQrmb4d397hml/xenI9uMniNGAb95IlS9vaKR/k8dM9ax8x9SjfqT5hcKulhYx
Q7MwBef+F9s97Kp+r8Pix0rIVKy4BAAvdrcRRW1PaoIy+u/q/QxUI7W884OkHJmi7lAAcxnSLCQ0
wVdzSlklPTdBym9vz0fE3gim1bvjRp4uu3MfVqs58PCR+t5CY6i9n8PV3CcH694+meivPd7vqffM
Co69UAVNDNcf/qnzluwtE5rS3XA8qMGVBNr9QsFSdfMOER7WEdttx9R3lh7r9HC82Xrr1CTH70at
QsS7YvEfSCWuyK1wXtBq9yBTa20EuIqHjX7b/mFJZ8dGbjxeZ0uX521LPQwbR7ue8zkthqA36RV9
eVALg2iWfJJA3hyxm4QPTngiVBzAYn6xRhOdumCnwcd8ZkIde7yZqs8h01Fk2mKbOzi721WG9HR7
qtF18pRb3ItG0Co/kp14UTp2k+a9NWw+hqnmXEpKg71vWOy3rFD9GslTtRfmgwLoDHridKRnMW6n
ECxgRubxDeKyDjP5zPO9ELhqTH9d9XhjSH3XMlHExo8hn+r9pPmK1tl/HIhZdRTzhBaFzcVZeP8E
wttz1Ca10GxyDTA4kc7u7AmsuCxd1LtTwnhonRaMGLSXcKsbauyJIFEGQIqfjD+Jbt1tLN0mn5fW
9OhhwEQIUmyCIivJdS/xtkuCkiOCEU0QdUg8P25/Ql0sY4ZQeuGKm899kQxeNonXK8KPu4QIhxmb
6pZsydAkcAikD9nVQUTQ0i8Ahju/qXRx16khWiHlbkm5nED1yQ8LedoiF8fZ0KnK/AVoABv8RLYZ
huKHdgFKSrq61QNOGI3wB1AAkkvzaaFlCIREDm1DjLhP61DGPHxOpAgN9aQeQ91kg486GMz1s1e7
jOaMzwQzqN4C13aodLdfgHCudRwMhHFRsbPC6xoLGGRK2MqXU2q1NYIGd2YhrGvSaiW7MGdP1XB2
L9v9kSVMJKXRFfH0gcSAvTzyRG6oq1Sw7O4Jdglnm10zMPlCLln+QeK6GE2Efz1xPK9TxPYL7Rwk
k+VuzNogn4Z1UeioDWzsN3yBEq1kCEaUJUedMXdobgyHUq6cZ4rHma5i4OLigKFepbOPhljG8Egm
x6iv4bcZQ15ML14YPOJ5WSWxFhxQDG6efNU4bC8O899o2euGRtxHjjuvhEjvAf62OGm2cDhlG/6U
s1Rvm0OBTiA9N+8B/OXZ2ou3M1Z1ojVAwUostEaSbkviebeuP89kMMVe0HzSaO04KMGABKMb4cHM
1oIZSqxLpGJyJZLFMi/DvhvueP401M2jb4tMYl9nyTAN/zmHRp23IRk9OGiMczVD342nWdw4pIWT
ctXc+ZAiefWh709hw3Icer4y/MpmkXnb7304pobHhqEuiUxXYt3weIFVL6mnB1Z7RBq9FoUVQIjS
IBksqlNAkt53Sj9gFoxDvmiVPa4lymzE1ZtFCHgIfGJ/n2x5VZGV5AaEfDZHxd02cZQ4Aeiby/pQ
qUY43A9B2+F2QLyGNivqMif1WVhWLjy7c2Z+eR0tUSUN+O+xJ/KsD350yxyND7AV8MITdPOOnlSx
RMYkxtTXRL3FmRSb/Q3AmzlzeqYR3syGp3AAM6eMq0KDQMRNMqak6cVwpU24lkAouKY/l3P9T3gI
T75dN5gW7epflTp1RWCBcnIcONjoQ4GU0WIGj4KwHQZT4fm2MdQm6Xkwpk2hMhq2MlMBZ3+B0pEG
+W7aosypVYpupTd/E9UwS/wsd3rFtNUTMamLWMsu4MbOSyzQq29lGUFvjN2Zpj/R9obCbZvebfR6
pXROLA1Qru5AClWGFNvDqkDw/U7z1ffgf5vqmAtwrqnLni1ABuCcg47i5hyN490jeQ/lfdM8693M
dth7XFqhMODxzIOtey4+xAcoQrqgd+bkf84hdBoHQf/e7gzQfjPSdoJSHR7w6tZuqztEyUVzPL9z
23sDDKjWLIwuBIeQ7khKgHtmgrLpZMZeXlaIACuiIbZk0P/gcW1VlgH+Wfv6iAM/ksqkka2F1Yi6
sOq3T4n7o56EHWLm03QL3ZH9J/F38dphjsbJLf/S5ar6pmy5VmyGJ3OKIRqNCkBS9+to078dm1uq
Om/YCFotS1nEOURqNyMMe/m9LSdPqjXzI9DowrQGrIOZBAwcZifJOH8Nd3owHnC37u2lTUCG5UeI
VbL6YnckqQQszdnfjrM/cOmTiye1kOV8IjQAD7sVktExFCkzt0MUO0XyKWu1wqfDsVdP/+O4BimI
piMdXcNY1lUSYnI/1fGGI9clrsLdj09zKR0qnF0h0skY0mGIXlBZn8JFfJTZjMGp6fF4QNcRY4IM
Y5NI6zl74Rg6ZWpFeTK6+42zwHwVj8gxc2T4ZLhlVsQfVfUeUO6bM2cm22LypKHSQ2MOxr8OsL0d
8aHvkrP/+d9NgR75XFkzWFj6CMNEBJl6GO43yjcXBxF4OB1mc8srriWg5MOl1qw2qYD+TZ7gS6Ow
pCPlTPsGUJCOEaGW+wU9477aA8M+x/gBy3U2O4h9iSxF/ahd45eVJ5v5zj/LVqV2uSE1okMuSmvo
TqFqmenA7oYMPJ14vda/scI2+AlWMY3ELIC/4PrM0PvVB/ujcdhTJ6BLXDKis3x30d4+GOKgg9k/
F/T1A+fWz3PNLi2O9+CHNAfAxtoAGGi6PsPsZlyzAhH3wCB0zFrJfh7YybTKwPjJ5ZFLPgw/vMqB
q2K7uXodfHxaa9K0Y2d+czCSnKaaBVjfVpVsY959t+4BtEQcvInygfCeLjtogIvfPybc8Ly8oMjS
bjt0/U1b6OEDc6MFHZfHJPJCZEk9ibecBPebv/leNxT5Y5DchOQqDLbKT+IfOo5pRTbsrmlTqvsq
iiMRDqEmX/2mmuLeFVl6+rj95fP8MbpiN5ZNZcWht5wtiBZRXvA2v+hpYn/pIj2hPAQy2Wz/3evL
vbe2yIi+MWVQpngl3ikyiBZA7sTFPHO0u2bFokQF2bO964UdF2dRbYPHcAR9uvNDk+RJFcbDLXk1
wmWbrkkvBJpBxA+HHrfCDEYEfEDyxtbX/+dYk2a17GD/8aX4yXs+FWKSmxYQ7LACzPRmwf/2SKsI
T/9Qdedp3LnLj0PiYPzmlU9sv6/RybMiEd1Z2aWM1HlLNtVu5/uiNxGmwTWIekeGrIVgPDjideId
Y1O6I3gkNOoKsy5P+2nG/QSLWbYcUMoHVM+NFjTZknvAK4RO8rUZ3VA19ahUbmooCHvt+NU4GbbJ
e3jmhfXX0hwuZns2WPTTNC35ygXmWNrjUMk5pT15omKbB75Gl4bmANUZjMJEMMZJjWJBSnFHcszw
sizO2zJW+I7XCh1vX+w1mLcT4oeObRxunz8XvHPX1eaNDCgS0lrlisZws8wfA3W3RQO6ucwA2TO6
EdoPXovdUx9xCGTM/0EfmD6aWJT3SJFNMcbovpcd+Dlju6b1YfArCY0J4+Cnxuzg1fUCfRnUa2wx
4Am5kWD9T4819jEMrE6ZIFMwkCq3a6h+6iaXJW8gIRmyUpl47saYKaaiDnSupl2rFC//n5KmaN6L
TdZEzwkX7ajWBXqiHaAFFBTKkAJ/NiiCio67okm2ObvthNNQeQg7/HOM9jplnUnwDvonIZXt7I+O
OcDuHOaycyyyx0Hj0ixOUBAgZzFOluFN7bb8f+HhfkrmSlfi0jUFTV/9ud5vFB0a/oYRHH/RSSvN
QfjHoUwxVl6cmxws0l5rxWYduwTCc19vJNDN1vvjSep0ryk/R9CIsAho4Fp1OwnnV5JG9/bJLbXh
nYt4lpmo1T5eQcKZig0RiSw0auTJs3QG7WjvXXzdjbdzuilXi6q8rxqSHUZnXgEEm92upVdAi6Y3
xkVszphh/P8C/KZJzwajzRNyJRp5La/EhqewNwjLFU/1Ua/eyMwZJW/GB0wFX/KVVRBPnHU8fJ3A
2pxJ40V7ZIlpsB/HOIa5Z3mEG2sK83Xw887y8S1xHwFJyS9tww+TUcydjDUAQT+pErtiLkyNqhbx
w3R6LGdGdvc8wbs+D3O80cKcsaW3sgldbNitSzhYNmoX6zm6hI0QVsOUqVC98w+LNCmdJLXX14Is
zmUkAi7SA9FWyd8qINebiUtIRjjTjDJXziPHc0LQNBXPyn9yAup1AAwDT63RkpgcU6VzvQSVGAmX
0WbTsC4pcDr7n1tu0HNer2rX8x0Ty69Wms74kjbXYW3rbjAEPLBfO8R70OIehki6jvFcPlvZ8+dS
LK+8CZlhTCQuMOOMhAUv0Exi4mTUd8PqrHrvhgwkzpnP9JXFLWiAJB49Cx+VvbQBnjGB8InnsDyp
WlAfBZLmIrikUA0UJN/Pyv5hpRBLaxcmH+xIJi9a28HmczeK6sURcv5WQfQt+JNrrIg8JkbhRQju
cTQPVR1HKdRKvhGVBRqpEIxTc4qkysEpEABnHQuIkjEIQpqvqhFDNlJrSAFDOVK3d/jpfUKhIQdQ
SiXblNMtNgzXNYFi7wmsiquDSyWsR6Po507IpBiqn7gJNTTsyIJOkzk/P4bJv8g4QZmwi2XKVm5/
ld9MPaYDJvOPj609NNJ4dmGeblwUslW905lriMRGmnxg2GUekY4t8iB9ImKcYOAblXjzekS7vTJf
scdUCmlvABtuNbzCey8i/U7rletjvzls8+N9qr1GxHKN7pmMYz4OoL5XQsBMPJ9nHwWn2tb8Bycx
/7WTIE8O08qI5tJaGvoJcmTpXkyz8IzmiWlTC5dkDF7UfQqOWQTCzYME8P/PfcIgtMnQHil5ixkT
yRf+bQmDfgI7wZVCn5pQEhXAwcgVb2Et7joLfbYtEU1oHcdxpOicp0jB4cLzh7nzhz4896Jc5EpI
kbrowKfyFb/1q6m68fBU3U/ZZL43DYBkVWv/x2UpEihpaZF6JuJ4FAY76Gb6nDLhBgTKywR1n5ML
sASJnyfl8gBdaAm2C1FdxsEhaarXar6pQKfsdP+J+gFYwZiJdJ1KpxdL8TgHaKQPZJPZB11MhA/1
5hXdlZZO7PnLUPcoXjuf1NOIpWvL+KJ+jJURJCl1CfqNG17S8SwA9ZYUSpWEzzSFVaCkr5ZZskci
laXdoWpJ6dPMM2kyBAZeDxvXXfuTrZ1O47CAU9ow0QhS4D9Dj4U/sFhhtFdKG0qVSLU5NMsMPM9+
/+VqfAmAd4s9fAzIGJOGww2we3y8dH5By29nmkVrY+Vd9v7cSvUWR4JS06uGRIiu9O4+8OYSTg8Q
pnFlOvOHNlZkFJAW6RnGm1ye+ND3tnklbu6hK13n6qWTi6A35W7WamIFeq7c/WBNKd9G7lXnbpZU
+aQI3MHVFsu7ayeMRpkKvIOltzrXJZNPcsMEj96Q6qs9niwJXJeJK6e3Byo8V9kBrXGF6CmAifDN
eboBLIw0fz83+kFyMr5OX95g5ZyuDkJSTXhC+oMo5Z8nArAMG1jlIfQGM1ZswaJ6T0yoOwsvXU/Y
iFwghNd0zHSR14n6YJHmDMPhoOsHUcHfAv1DJJTTgcM35jOF4H5xHYknk4Nhx3tkByfw9yMKD21b
+OA938Wax85hmHKXnWOA+Q0EIbwahvmkF26CcTWYuWQBULSGGExNxJneN/4AxnZCw5oCUr0e0ksz
k3jDRuFRi7RKCGR+glV/46n2kN39nmLjqStbCpQwg68W9RK3v0nMXqItZ7ghVcxbpUvGmTkrutZL
5MBlGSKZFFuQu/K+W3gagLJ08oE/fTOYusQ5fRDobEGO9oval6zVPoJ8J+3E0dVYRILVXrChzZy1
xZJX5WJFYMy/S7Z98rTWWUD5qKqx58c9tokdB4kSwF7qKQosThy//lWxprELwQcdMtt3XD0n/RyK
92pfk55kVxbPT/zLII/9Nix9BBwdMjlahH/yulJYPvA/zUgIX9MfDbtH3BbJ3xxkA3zU5GpLHnHO
LJnPMP2O7cXwVJmTULrZ1Up9sIKC9lTf3pC/JizuySV9UqCOOj5b4mTygRgm0Hc/9/dMPocPlSS/
sni61GNRt6ybn0pWh8AYqFRz3nqVFPeFNZqnSZmRa2mO0RhiKiCGutmoSGZNShGPUkRYe6RwXjov
oYugoL26q2OCcG62VJvp2wlGmejs7wzDMWxmQkkcyZjD+sTG0zzPEtZ2f9rBMDUC61dLB3HXz11u
hsDzsyYQQxBeZLdxZ6xltAXKpntR+B8pCafn38wovh/uqQvF9vSe0eXrr9M40LWpaxcJFCDMe5kR
PNknTEeUokzeipMTPwRBzkQ9/EA5vkMTJrrAyn69ICcHV3iXH9kimsHMA2ry625A43B40RRpvH00
b+NoJjL8sQMG/0uIhfSjSIZ3m3gREZk5EvcwyTktSytPVWA/MIB3o8B0ySIpGqyV3X/mRLLVeQ4Z
9Ii/GSRH1sjnzNGwZUZY5GgGNBtOBF8fRsB1gb0sBkNJI918Zu1pkF5s/qiYp7of87EBJPXFsEDS
CzD8Hzcifa9s+HtKN587+cpDO78o2EeCYUxEvfTSs/OqTokhJKPfW+wp7VZYp2GKArlj4o1+3t91
c7iUuK7JziYZ+no1gTRgCR0BXG+b5CVoZ2GYc2LpY/Efi+BapwDn1hfAx+rrLtMKbUfoOzEPGJ0x
Ha6mg61/q4/kwyotMMVZaSpGCslEaQZEo7Ul3Q1LnuSfaz21qlz6FX7PYnBwSsoFwwoYlIlBkymE
rtwHzTinjBuDNeYNOcaxYgvWyx2IHh2mQjNNXm8x7CmrPluEy4Bd9Ruz3YYa9VhuW7xob37/yr4B
6J0UV5/++33MDguUBZQgkQxzAs0CuKqqdczOdRt0HW7nXqSmJP/BEjAhF+zCW0Xx9IpRgAoPCBUh
dxzJeJkq3SOG0d9CoqTyEtqvRg1Oh6KDtZXVnB9Dfgj2wo26bNQH/B3Y0vJsvkpgokXEPOM+L+Nh
uVIXOg1uOES/vSEevwO6qboGEGAHkgYqnaBh0dHCax/FvWQeUROB7/NJf1u8znnlU5oDdizYiQ+8
wQvRnPRk0S7AS1feRJhhLiAvyi23ljvwaaXBtyDZ9gtgEqXyh21Ec6/MzlttDfufu1V5B0LyGZpB
19cLMgRlylmTChDyz6qiP7iWKYqXiRQJrKVR4TD814zzeSgAJOJJ2KiaoBoQmEzyGCaWW82e5BVt
OA4Vvi004DZAGbLrweQZaHA9rUt7WSmTkiJNqVZjlecgDObnlkuBazBVEX8kG3UGllSB7nZiR1iD
P7Z60iHWf2mRE7F4RScSM9ASXZlBvHvGkozVGGjIfBpC8nb6IAN1ncQnHvdkReyc+CcH46GxZBWY
iqjUH7WiNrIGF4wDOdwr4n35p8j+qqz8qHGdSH7886V0QntxxlaliPR7Im3iTVx9jqOmipatBuur
Zrc5nmI9Byhdzu+2DNHl10bzj9Megsi7c5oP+fZksQn9sAuLJkAg0MMGMk1+R2zOitDk2T3MH4Sw
/gD8NDdBDhC3zsB7j7S6pxKl54bEYkXbPX4dJhHqkOqP2YpRRVeTS1PGqh/yEySOgZYCJCdKcnEh
RzPEWhjpn6EdHcYr+xjiWeEAgXw4WRK9jBpafnnbqin8FXECwqM3eW4WNY7f/E/vudQJGbXdAUO3
yzzCSM4wHPHhsOCXRNrvJQqdqz4EjgC0AQwxoesgcIGbQ4dB7dbdPaBV9oaAAqbFC6ky1VEB7cbX
6xJ48b48qyqGo+lgGmmrPSeY+sfxw96vCoufS4InJrr5CPv9EkVttehzuJGs/qRavBqEKLhJ09gu
Wh0ubIakGiOFg6x2qGZCHWgAtLZkR+Yw7zK/KMTM1FRsa6GnEw6qOBIDL2YKpwYAcCN8J4a3+HRK
0LOqjTYMU4+Z1741bqpdcmwIZ1pbnsxbfxl/nnHc6b8iumy9NC/ZdgVNYfGtnG04B7S5eRk9/a6v
zitGSAXidPoI9ACt5cswFFg+dKFFHKaPw8gfMF1ylCACTTJc2zKKyfNn+bVYs4sJaconsZeePnbZ
veYyLMVQHHD8ZTy5xUW+cTbieyDuYHRL3Dgs/NKY6IXOtIYaKExIqsvb8QiWwvIHkwcdV3SsWLSx
04Z6kmPZQpVcS3WxPBfAuCqnqrD3Cy3rNvL24y7uYykF51UWCL7Kt7ggJpsPIhnN09s1aZW0NMer
8ubi2dnaRf4fx/0m92ND3ippUM3B/j59WdT+Rpf0Ck1zWjzz/lLSTqtAaBCq4oZ+OgfVxflZ4Ga8
EzRPayU9nrvmoRX7CSpSc5hTefW2kOQYdqRdeAUOMef/SO+t+88M1X9Mksd55m3aOwg6TLfUeS+A
wPlQuFx06+Ke2vbckpGM2d7t+Iyaca5O4q56ksMTBqSJmz4QY1e4sfUbgPMXYj/EIsxQmQiqgdAR
0SKV/SzCWddpOtnhdnH88xioWb7Nx9ksMaXK+BXd9Zg0Q4iP4Cy58oFYL8TMJgPPOl5voZ3m1eTx
ZTJ+i1EgBuT6a2edCvzjzuHuxnGWH0XG2aUOiXco5axXvifl8padLdkeGbhqw8cBJk7C1L321pvc
cyy+g+QFG+MCzZx4Z6HGNsB1S0QNeIq5adIGI/VYaEwfON0Vv7BtPCV2RSW+MUuJD2rqgAnW12/M
SfLFu66J3yu60ay+SLcDrWqxMA7dSbtzm54elqQc6fJhUkd/zOhOlEnHiPzjvUyl6IzVotOEmi/l
BN/vpGqB3pB90G4Qsl5W7ZNLvNCFlOFAJ0bcFxp0AuJVtVBLdMByFeJBzGeppPW9ONnr3EmPT3E6
qRzIA0imcHAdz7tOWqnbAlHwysIEW0mUOjyE36hVeMpuGLxk1DlOHvUepFu0cpmYq+8A73MuyGrD
pELMjDV9vw6704wdFKIBRotdTTtiEadXNVxlz3deJMHWOZPgYLXZQU2jVMbDZXaHMOwEq4i0t35B
yfQMaVFC7aDHd/lfLNm9sBCVpV0fUNQe4RXl7O0pXusTSRC67OI0nrwWdfVxCiOOTYJ8zuFmQcLx
jJFk3pneAxiL4SCrF3dMkS8IksbGv8CPklV3ehon+grri9qSIscTJRwYxi9xQ7ktO8H1pOHgq18Y
4mmFdBRfSbly2xEwC8+kimcq93zhmxMbzJFqjXfbrT00nIOublSkpadVcyl09+38wUfxx5H70A+S
mk6VvJEEJFFywDZ0rYKAqT5ZixVEIQf+1wrAdGg/vOwEp3hcvXIOdW18W6+cDUMCN6QodlmoViui
W1pnO7DcTgKU2/see//JfdwfRzpV7CwPQZo4WxATX8XIaajnbKEZrV4c/MW2f/7EEDRyGqHpghiJ
veGOKHKfenEYNnpA32CiZiVlV1QybFe+JgkL31oKHexRIWLn2O6Arfs85Ofmszwtp4sdzziqIFOy
eOQFhK+3imNC8fZu35bBcJCL2cBpEoExBuyRaFTkxCjw2M5btPC1syskWxY9ZBx6axXyKygAUerJ
58xU8wRhF9moomEMn9BZUGJkgCQVx4ISbixLsPBdTRcvQetDkz19LUA6+9w1NEgtq+v5JfbHCIie
iPU6elk1w6X84PmYrT+9A8sW3FHZBtkKAXXx7kIPDr8ypeazxpVHt422feIvrzi2T691X2qORRBM
VZlqSmSjcgbeaoVHbn4hW7iN1xwt/FEh4qpGKdJVTSdktvYJGoNMoDwQtxer+DzqqRG3NIWhhbAc
rgULLgdtzc09epDOYLjaYGF43bzKp9tWIHdEHmftoC2OU6aF7YdYt3DgF4dld0XJq+m1W7CJQ8WZ
Ppjj9HtSOgLojg0actyQfKqR0phpjSF+CTJ+d2NL9aD1JjUFpsYI/iZxdoHV4J1hq8LQrNqFp9ZS
NQrNzP4IxYQ5WLeNnOG0Mj7go73lzbjAplI+smLaQYnzIAWxwsf2PX1JZ2vsTtppGGFWejhSbexU
vQJTkr6HIjisSua6tSCDJcGtEMmTFbSX1t5ih3UWEFxG1l0zvNSt9ie6A0PmtZp6v8UZPwXAQz5A
gWUIR7Gbxe/kwzkNeU4+cdP6X736Pod8C8G27UnVQHaE82TqsOqKjiODTAJEAe9q8iGBpH7PsTKW
2SjyISjwErlbOxZ+HJ4RdPYcDLid0wBus7gFEY7VI+wnHcoGl6/fezECCPKkP6hl8ze7RfySDyUt
I8DGnyokILamh76efXni++ti2Na9pSCfOQnC/L5C34ziaqwFO5MvuYtP1xplOvXrsJn/JYclwdBH
1abthtSgcxb/9kfAJYrRx/BUC2/NZywxvUD6d75LWeA5kz0kswqzVy0ArvXJ480zOr4LNY8UX6Tk
2ED3QRoK9olQ4SXgxxwuZBmjYrpqy4PlS0ZQl/XqWiyzFMmSKXrxsF8YCT7pKCbehMGZNG1YVcEW
6KWezt4luPhtObG/yRZZxWZCe/F/QQ93wMviLs5dQ6l/ffPH7JSXhhDH3wifLIWEvXvNNd2kmsc9
we+sl6rbQPIDFznmiAwwWG13O9AnCpQWEJonTEsI7RGOcB7fSUVr/3UIdOphf0jEcNy0QBcDeGrA
Qx+LGPbtiPXZ5xCBaFKJL3pramT5jE1GBidLEHW2WKuUqZf7uchXmdr3Sn9KDr6Ike4ZehUSGaXY
nbM1aSdpejb0/A//8PcfcZF+gAEfQwLHt9tTWFSRvRzSeIUiOs+UBcWKGQWnRp7PXz4zYZi5u3LO
sQoSMD/yGehEMH1+BD4fyONIapcUsVINEBSVo/qIUThtzoAHceQpQcjgIqz6MmRRK6R6cSaXgjL+
/dj+AhwWHDWlV58+7hMixTWVtrNfFTGJvyHN2ETHMB7N0oOgJh67LnjYEdxTbkZzSdo9+lg3eRyA
EYPfVUKoi2fMVMRQr8A/WPPg+1A9yXuJVKUv7YA4ASKt0B6Byxw056cxfUvfKOeS3vdqgLCfAL6g
hFWl98kZs/ebL6NBgyIuCKy4GgzUXQqnvR4XX/MWkk6l0BAlTo4pVdgaNmq6r4upEfnVhjoOfU2b
+4vJVgWwyDZz/c3yCrLUsteQU8VmMyrFTK+rYVj3KEjUPLq3akwTu5iTnlIfWSlqYd2MNtDqgnLt
FwAL05/qf+2RCrQosia08b/z7C7GERhiYFcMKSLGRC9f18c5rraensa0YJhOM0ycSz9cl49xJSR0
4909qUuLT9815TdDzQD2c/VatG7R1NRqCZcQ0LbnaTDJI9pJaueE6rtMp6FMmc4+FKdtcvALBCKU
A66dOFTj3CZE784oW2y89Iszrx3uUhTzaYW9xexhZkEbNblTtRzumz/+QUENTsnbGxG3r2+k65w4
uKSaOlBHl2tourIoOwZPreSesS4Li+fEjIw1Jekdb8LwM0TPQiwzkVmZtMmSU34z7277S2ElsjT4
IkO1X7D0UeunmDczw6q5V/PrxNz6ZkTVfpN7Jyjf2h2HnkArNTaHBrKTN8bcSeKO25wT384NaT5f
80BJvmUBl4yjQochyI1k+qnDQ+s/M0FhF0wNz9XcBQu+ADLOaNSLFo0btZM9WqVetzYCMXpL7/th
p961jiSdAKGVo7HrLGwgzVVhs783t8syiHgbm6i1nff3VBsQWMmkAmkFuRFFX3MOaeadLzyffko2
LdI7Erg8bdhIkAwvCpY5TKX8tuWbBW3bnoCSjOHgKaOO0jBHdqNWANb9+wFsxqWft7VIZvDOKIRU
97lpHCU7LLTUda297mleZjzGZXAgqJxQY7r2UAIGbAqSowyLDCqErbg8+q+HL+9GdOULsJYDUjdg
td/8O12HGDy4XunPHQpYHywn8Sl4DEPrhxXssDUQPjh17TnAWFaM2RguhUVKHfifBUeDrIf8/E/b
FTDzlSSlDO2Fm0Mp13uPFsVmJnUUwY09zAicqQmnXr89fDBX6Cle4yTF6q388M+NfSwfM3FHMqy6
n235AjN2nEZw3PqJTtYKW6AveKzBz3CamqTP+IlaEKthFuh5aRLmW1StoSd6Lg8K+D3f1Pk644QC
YZJJnpGa9DNn/IR2mp32up1vNwNwcNhY3hZEh99rto96gHPLCpi3P//ful4kFQlAgAwmdEIWveNA
YH8uB0O7sI4drr5QQrPb5dFCBZvzAOoPaNmlhzSnh7NofJMMEpfypetxYiYI7uWMLpUgTWEJ7Cgh
2ZJHyhFa4IQRB3rSqVVKRm8jUZYzM/DsCXDHduI6IcmKUfArKlZDA7tj/WP6uoyZqYQB9KjznkEl
xIJcEL+EKFWq0atUI6uZb5DLN7waoMbs6aw7dHZc8/j5798sC6fkC16RhqEdAfDEOVDEFXwQTOS+
JXXlC41K/ILa2JOXHKfdfUqE6OCubblBpFOE8S22th7bXS06EIyD8NPZgGwp3skveYSrOOg9Sv5N
C/vnjURaHqRcrBV4sdylVgQqRg9z62F3sXiQD91ZnVwlArza1P7QeW/InNVqPitaRiBUyk4yp1P0
h/t9Kx40MCrWExNaykLzYiVedjGkerdjN5VHqdpbQcYUYbgBmyVRrRmW9/xGkZ41DsXNWHLrRosf
sc9gEkibYw81lYpQaP7er/XihH+34dCvzr943T0Ud8lBvQpGYGfLNZMjI3BnHlRiWUmgeBv+Jltw
KNFvOHoooP1DoGdzV/Dd064JhF2IyYL4AeclSQVAoTRHW50wurNblMlHvnyk34TNwzloMvoyqf0S
ZJT+Hiw+WdrpTPNJkuf4qeifBfsINYOSAKrgTjGjk/HBXsxxBIEcJdYUNE9VitY8FaapF4EIpU7M
OpyVmw7NriSseZ1pHhNAcqmvSQXUZO9EV/L1izxBVQAxUaln/0zABlams/XF7EhDjmvzhN0msh8Q
MbRj8JMEwaiZl7zDpbCZxD/RIhpzez8dYSIqex+fRuXtZ6QcfaSRLtSp/LOoWyKuJAzk0JBd1fiM
JsEoRVynpq4h01k7EBqCfcBzoums0aR+qU6gRKwIXNRX6W1IuGHH6/gUnglruGeXFcIG90H4CMa8
oFZkQbH4gzEUuw6d16QkTAlGiYQ2cYOHLt8Cu/SJtgCneiI3lXLR93o9qHMIbyZpF8BQ1bil5K8d
jkJD0+BWDuLHsrCBqthvOFDOPLvUw7wAKAPbcVq6ry0WZACGiSaGJKg1XOMxUL/0IM3JILT02RpM
2rxM7VOg8TSSrDUy+CCorGlW6H7IcfvT+XH5pqqKyLuKq8TuAA10Hl4X7+CvX03GAP+TY1K6nudM
3kHVyLwLmEAqfg1V5rzDrvd9x/g1r/H6gq8Z0zpMrwHp1/zvCmEmEgSZ+AIbZIkJw2Iugk+datdc
Nu5sS1ikefUEZo0fkXFtqdJVluvBr5sfKFFbwLIkxMObSQ1nAiCJ8XKNiB1zsXgo8StQi/staslo
fGeOl3nXqzfkjP+VPT0ZX/st6RRxFWY46NN9zQva1uHyFThW9YvknLkLnpJPrsnovbsu1MuBTn7n
gDdhN8rqQwQskCLw28qk5fp578stik/e0CZI5g8+hI6gKks6YBM8HSi3oFz+OsUcf4/ZoKdpEY3A
1flkoDsHHsBRSVnWOdWuDdEZv3RFWS9DiwVLPsorH9i6h4Je3w0BY4/Gy8FNJFH9TE1g4ItLGNla
68ZXXVJgGWckEEEduMTj/5Aj+XrZzguAPCNp6b+uGcR2VOKQT9bd6QikncMYXzoYCmyd2gpjFDXm
4FWiQyegwU86NpHpRCxu3b6idhvuRN1vI7g0ZGQkKL9xSdgoADNn8hdTj6ciYvEuSsEK43adLEf7
zgVTB+fbeiqa0nPjxsmJSGs3MMAx0lNix4A20807lZedMjKlJV4UV2LpKuCconIeW2MlqMILTE9e
ZWvonjGzH88qS3qOg0vg8ODfx0jU13m8Yxz9hXDXuFkXYYUWmLDh+K0DD5SMHZwnD54t/q260jGR
526KYEmtAxpKOzIm0yOQ99vfJkk+AaKZnFbY30h1ixM8tQH2VQ0YN2yF47xFApuucNnNQo/Hdrat
ilBKbh8BpPmY62En4gGZkjp7x4GY3ut66U1oVV4qUyPKusKTdAck9RQ+feopTAPpMZ+jS5APg9p3
Qg/jKf8k6hn2epD+t5a9qVcred51vUQ9dyGXQIMI0HIQmzl3OGNA6RckCPn4zQNvzFipCc2Jep6e
vkwNsQQXPihaz6yNH/s8gsJHlXdEWwkHutV+0vfA5HDxV6m96iwIfKVfLm5qfxl70SsCLyLxVo72
Yy5vRnKTnLq33jGRYY58PNd1Pd9/owRalYPa8sx+vOOHWZ7eeaYlCYrHSPjDxtARoBw2zpMIJglS
vyHS6TuwmLqEVd3jmdk++azJxyfu2yhB98n1O0xE4KhjsWkEF5ary5E1AbEma665/A+7m7vIoL2T
5qY1Y0YKwfcbcDWds8iFik1oLMBH0jW3KfRF0JwL7D1vArr2pGU1Yw/TJ/XxPz3caT2C4vh4tuab
gkDufCA0M8HHc4wYoq8gWVHJ6R+l1MpJ9p3C5rL4k8W9wGSqf3tR/6iBQiJMt3rr73pOiqICtXku
TmsBxO13ObuP0Fd444tJm13rSU8dfcez6Z0U15TCPOrj59/8aMBEz/Wjgdlyfsph4wrWiWqiXzQr
lt2kTPq4HUnE+kR3oSidLKym3iLVuxEHwj5Spr52kTcRrxe8cq6ibv2op0D0dLXPQxhjyp329fKu
o/IQ/lr1ZfCMu/ceTnBD0hAceT4LpnaUCPJy3V3DRRd/7ciEwOycd4A+9rAYdp5pC0h9Ur4WscoX
m0RdbJFaIfstERUPnmJMH+gY+rulEfHj0ysX1lZrLNXdSse5qyd4TDdmsGb4REk2tC2se4QFAVbx
L66ju7Z4MFtbuvVeDHwucvQc/bGaM0aPlW3JbWInoE60r0KgHL4cW3rXQatmkye37sxQ6q2NGda/
jnx01rYKzK3N/rdsp3BvXaSivfnKQy1QCzilhjTm8GmM5YgS42I06sMM1TtczYt4rTfuVfqqembT
cT8T0nf7QHp2U/HqE0je46onw9Yt9bkVwbcR+7E/dhMw7bBNQl4V9MNsNk+CMiqMg7J7qvTcsYnv
y+ymrn3cyWGe3sfrxMgQMNB4cquOsZ0x66kdrfdAMv6dU0A+PMjRxrpRiHSk3RNrwwVz6gcuv9MP
T+8OK3TaaVXo5thnKWglBPKIi8NqLpRtmnVp0WRUcRYHDVJ2JfgGf6A954RtLMK3Vd8vMemkIUUx
/Z8Ilowt658jkWFLYgrTC7wUolm8O8EiZstIL9uf5zIahWAUgOe7f+Azkf1UH0MKwI4URa/uTwlu
WYQ3mf52aJkurUI+O5m1qN/wuGE/ryNK1tUx9jWomXAE9Zn/g8vW/wNFS25oG2G4GXEXZPlMiPBA
vEoP5QqwAEfxS0Ii0YaIbkGsVfKVJDUih1iz07xx7JQxq/H+0u+ekYWX5Yhweeg98NSf8cKG3ISo
aHwAp9SaKT0qTJ179eMsEZftbwn97Z/lTItBDPTCWjNGXPRsGpnJeNkKh3fcWg0epl80bKaHis8O
zr1+0eFEjkoflcbZc0sM++C5EY6mFPMylY5q6kcrIAc0T9E1eJWlf9gX0ERhkC8IZv4IWexRC0cH
v2IGgXMH9iU99i01vX+mbrOCNVMOoorPKVzL4rEd64nHDODOcqD2WMYBDBOdTqJZtTqrn6OpARRC
zXgeaoumoZ3mBIHrmNUYTafOPmstemYy9DK55kSdHrnGq2eheBgCOwi87X8RInluR/6FxoIdQB29
MnEKgojMPsoWG5gnXXaYf1e03DNNKRcaZ39KAi2bqhbsOqZmvLm1Sg5P5YM6k/kHGe5sCyE4UN7M
AW3Ao1Ru0mgIKDPmecfy1KVFfFYeyvKPhvpP4KSgqcW52q2t3zmwjgFXjbnFKHUTXOMmNGSKZ4zB
MzZrm7dvyIT52BAQdzjpe0Ys0bgVusjTTHXPmSWzmKTva6JYpOyGE2stqP0J+Jxwdld5yNTRTl7k
1u4T60QkLUiUZWkMWinWQWvKWJkDmuL3Qldpr1AFHr5tje3hM9axlxK2F71rtViZPm0XlltkAJrH
0U0IWMU14cwFsx07Jxa4Hy9l38p0x2AViEJ7Y2aOtcANSkr2jAra/C3Ih01NUr3/cQUmOQUN32QJ
/o6+eB2Kp/qSGeAOvP5t2u2Ts5EUkxk0k4ZJHgrLzMYgAbPU9ShZbhnsW2YLAkWe0q052+EgxJ69
EkgBJyaElskiRobEUKm4jhs4xLD21pcodI749l2IKgiThe65VLEq8FMqL9QFw7s5TAEA+h52DOx3
7H0KZDl6Yh4rX4BvgcM0LMffM4ZhvOwttWBNTUC6K+T4FySGJMwFh/GNNnEqDlICqDEDFKIoMI1l
3l7p/pY/sfUigIv2cC6+aXAnu1yDLOkWnDKls/oA/7FAxvCXkRcyZYAepz7aawiUf7NuDzTqslKq
MIaDrJ+NNn2D3qkeEYeGD+jCGJFAP4kKxZCJJdFH+kxt81mRYbJNmn09IGweAI6ztIPLuCC1KGdW
iBUOHsWBD1DN8OR1xPucVSWT6PLILSbNNjgDGpStIwlBIFgI4jTKve9L7AMN5T16mkQr/8m/4fKG
w+XVChNILIZaOiVcZ72HgR5G6n5HhOG+Q/hOT+5jxiNhXYIaGoFyQ2H6ZeSD5PYtJCvG6A8VtqiP
6I8tszRrMRl+Ba6KVY0KTIyJ7P3rVBK2VVCd3aNun6AQVz7tY8Ad2qCrmmlvbw8+ZSjEVUH4leUR
HT3UyWTKibaPaUWsfjX4nHMsrj5V0KvalJKMEnHHrqQx03q1Th9FXp6FTdkvoKfpCJK2Sb/cZUE5
vbel6kc63/TiXTNxuZwVjZY1Y+MYcL0YcYgmuWVl8tVQTAKMxV+MGNwy97/5oi+ikMlwO/0qWEJ5
EKf4cjEo0TN9kn8uIcxx3betQK2S6GgZLAERHXJ4UsoLNnvXkC0BBoIDTsDKBZFBtc/ceTGe6+c2
zu9fqSpGPu8swYn5rRWrQ2Y+5VmPOIun445bObmlz/kRHfhpd8OCrhoHhEZh30/y/ewcSdVuKWR+
mZANJzjEn3FB5eIiw/1xWO6FsuDCGMygiuhWarLsArhxM68VKIBf7KAXw/hWzhnNouhvu1vXIUwM
POUZH75G+vCuARCfWFlYmf1Xg4568AigOYotmPoJ95b0N31muLka5nIsB0S4Lbn+He2ExQDVxKh/
37hAxvxSusID+K5mMu3e45rN/0siO8pTRt4CfPIRPssYoaKNJ5HxYUT5K/N44oTlGJ68kNsO6IFp
ETUa4JwfkrqlK/M/83h9VQ/1o7LXI8Gsvm7xPfS/nYPc5JmFAiivn2MdsGAfel8/YOacwC0ldnka
9Ry0qvB+js3JGP7CzXK4JeFKwr3Mo2SqV5m8yRB1GDd3HV1ErEbyLXxvh8DYAAWVmZRmg+OOKxkv
kRtRsvIN0IaI42zCqYbtbDr8uocsukbZeCbnOtuRb3i6vkG8dDcrqsd6G3hcbyxGXq63NDdxkY9g
uTedICXkUE2T4pF/FWXjCYNyXJY/6PCDqYcWuK8PNSfj3UdiCgYJ3E5HJiRbpE7SW9KtmykjiZ1/
rSeKGvwv93qG7TdPQDkl1+35a2JWQSVCHorRPSy3g8+PUHSVa8+W4cvcbbRFzwyMadA/oFtP3kf3
JefEPM/9zwBRUKUpZNDkI/Pb/3tjqQxXyIEs4GN+qNF4jyj3ww09lTu8orswDq5i7lG0QUC1tyo1
TaNYuFVVSq29shJ0wNNQw8rFJ317lkmiTUKHGaKpRZC/QW55je42vxPE7ixa+GXwMUQF6ybR0Tf1
LBwPKNy8i+nGPTcUp/hzMSr5zH1YstoT0vxqCMxkys8PRVian3pAthhE8g7YBy/uyYiujuTioetl
Xe0UrNltRVpxkIWVifIIp3YvoWsxeNe6fnfRZGDWPmw9QTkJHEbiwu4bYr7DMNSjYr6bq58nYqMK
JsgWZI5fgbfnwo4HtTDXBT+vtsGGyl+u6iHLBD1nh3cVzBBbkdFlMS54BTwwzM0VTf+pEbdhlU9I
heftyIFmmsbU35mp7sM9KPBEgbIQWOJZGYjQHf1MQvkhVNqWnh1qHN+bKER6O94yKEUJH/oDINv2
23W82UaGKzZ2AW6qKHLf4/GrHB6xx+swwhssw68uTqRSgN2U8NBAcUmk0v3twqT6DZaZOh3Sr8Uj
Tr6EaeSVOEOeADVwQ9yR/DbSihDt9mIIHegVEbzp5USxdp4bNZy/PEZlZCJqOB4gmPQkBnIadOgU
3fmi0FcvCQrD9RiK3axnu+clBo3ZoAkJUJ0AjBf5JXSUOOh4kAfeHYlhgKZENqkZo0Foym6h1Ynp
pSRGpZefEFSWTnkJgqK/JPM9CZ9oP7DBKJvuJofYnXwOwtTVq2uYwLvZRbY2r9ZPjZZSavC6b+aF
sTz4Y6O+uBajuQ4lZF+QV7rQyDFATp9AXFj/+bgaenZtPcfro6KYDW9DJ5HUrkzr3e/62lGBu3ME
XnImv67rFMLT0gRzW6/yCk68zjHhzCrktJL6BJsp62NP1ToyqjEjAY1thZw9QlJZTaYoHzpCd330
+roMebZhM2UUq/1Uem61YZMYoglUdhw4694u/EieF9liYWBjJnobolaQ8dv3iDgEAYMr1GaUgqSA
OP8fY9ztCT1cam6FoGXpQfQ/P/B1guR1akDGjurnh5sREaKyOqpkvAebb0l7MS1F15Cyf3Gie0Z4
A9FidjURdqlykVC550mz1JcjjhcH3y9NlojKVh1suFusxQO9CFwZ4Umz0roVACAslM02YNDAu6LT
HE7B6OLXD+2tU+dYHq+U5cnuOBz57Lcv0FDJdKu9NzYIdUsgGVE9UYBBcy4ODhRUUKksNA7/NcpD
wLjI5CRzwqAOTmg/KeIjVTth8c1kh138O7QtIpQ7ZA9voMs73HG/UGcMRc4OjcTdrL5DkCAz8PRx
gBJMfP3frTzPE9IQXN2vPOgKkk+ghpuEPJMoDloopt5gwFOnOzFtpYX+YfO+3jPZ+MGy6uhkLeuc
+qiAKXEKwH/qd1s8TlqfnDpyjREY8M1fAuLwWvNJzeAJyzkJw38NwOdV4qZ7EcqvrASH5DVfHi/I
3DOyL4Mgu1S93FXSjMlp3+WzZtWVdl+vmp08ByG+IVRPZXoig34Uhn7m2ehdwf7FX6RppneojMxc
I3+UbCoH4c/HPH+uDTWrchzQrAaJuGXBtdlcSW/E/EYdDnDtgOJhNgymiG8lOciyrKNsfcqkJKwT
TcM8nkEbrM9XLJGpNqGW/f3fwDV9/+sfn7w8uEA6GgXaFJL2Jb8ODdyY1FTW+5/mCzcNMUtGM9Di
QCveb+UX9fz+bkNPdYc069R4K1HM1cEx3Ftq4j8KXHG+8K/ZEKhRib5YDV97Pc1L/3gJIomBFCt2
FrdU35t32brjjtxclxo9yGZmW5mXUTnTGdAYeUF4DSzpOgga07sRJ1RlS7Z5czAX697jFCYfpimV
NXbFWGoTu3oqIMFcfsR69Twy32PstN21Y9ZvcDMy8JyMB5lz4muvO3YJp05nGGeTE/mdcZ6qPShf
fB3tV/TWmL3pJ748TViJS297dhNbaF1n5zvMEinrlL2t0WbeXsA/fKaykt7CmV2C1OxcnWd6Odwf
idwAG0kjNki/EJ3k30ivkK25Zh5KWX7cSwTaPO8ME/yR6v9t2D/AkfOzeh6ZiEbetiiIfmQ0rl7K
wD/qZ5ev7BImzBLUWm/8hiA8+tqFKr+Jw123NrdpTpckzOt1Qhiov3KPA5bY9o3I2Tj4zrWivSVE
ue6MxSuruZPP49z1Yb/swnGx+bqGXhXaLgdLX5yndWAQP6JRtHeIKUrw2WVMhzsZ8M1JvoX9Tcov
q77dxGSzTMu8J3pJFTLQhtZrRwLfaXXKcOrZTRyyWyowsrBEm2dtQ7mkN8w5//0Ma6tcy4pQhSkh
VPzr2OtTieVU2xNBmXOO3dqFFbHZevm0U93ugkzMQ+XDnuOISKQ45+ihGI+Rb7A2YoFY4UzKSY9W
qZv73uuObmpYLdAxfigOLY45cwzjDcD3XCaAcKiUuZZmLTmB9accA8RyBdC/B0J+EpuNE6UJd/tF
7nsbR4phbkK62Z8uZxjeYJAUzpso+o5PiTBwt7y+bDHVxIokVDLElZW3mX7tNl6LWgK4FmoS8OSl
2EFINhrKkdTNv9PcTZhodiaI6/eytiE9YVW+LBpF7UxpndbPH6MdS1yeaZAyab1qYwlC1ToGqaen
RTCMBDv0GeMuwyF13HtKtwHwLQ2Ldm5g+3egulwInxScp7uS5KyD2ani5Eo9mV3DJPzjYOMTJoMC
agVhpLHkkhBpKEfQ9RTCFyyhgCVAK+UA62yXzOIrv6S9j/BQ2rilGT616SiV0no7cRk/dG9ZX61E
MiclTEIXnYdDlO79mvUMmqd6JrEoUKik6sbT/5J3G0ulgL22I/oqgfMdc8jYs2ko1YVcL9pfl/eU
lwPA1JmBfFmGd8sgox3WBaovgstRRWplzs20qfIt0pkd//Cnm6/S9yUdnyR9x1HZLeatQ3/b+SGu
hIWCbmHVL1AeQHXmsRBNr7ZpsZgVhaehmfqHZbYOyYazCDcNFpIg4O4/p170oqmMD+uvYGKTdJyz
X5Bgw0o8Gabfy83uOhLUpcWZosjfoEdLzcEWeyGDRiB3LTBjCfrQ8vT9FvsBAKS+bbxvauFsHfhs
mTUDfXFvDjBOW9Up1eM6KgL+c+q7y0JKGlj5SQkUSf7r+GdFSTmQNjJbLPiFfdF3/wOXdKmsq+T2
LjibPdPuBgThgvI0+nM+ir/aRHdimubcalJB+EAYwCKx1SSt9lg75kIgp4ckMaCGlnR5wI6CdMO/
uhqq+Om6ru8SmoZDMic9u/iDlLc4Fmnuz8euLonH9RCfCTAMzK65Pzr5a2zrwALw5iMHNeZq5kn5
9NZI8F7IfTNMxFh+MNRp7rt7chbJZucR/51Zd0RTXPg5tPYlK2kIvIThn6cydp13JLM0aMxTst2U
XYhQKxNEKr810HTae0MG78iyF7hFmD4lKDR4UD8JfaMGY+i9WBZwMznPtnNArPd6lYhHzpYsDnvU
MIZmTwgEVnEPxgZtRwLarqS8EHPhZvOtW7MhgqHnbCVgQ0YI0dwMa9r08uEgR9pBXFd20UMGAeCq
9i0FuJe8wA4CXTIO7V3IIG0zI8P16wBL7+fusdNcy38v/WmpZGEgZc6rouYgwGs9ljZEhVSC4F3Z
lEDlPw0jrgTGS+TlpweCOX+wN1bvmeqetcl0KyzraTXTG4Ojw8yJrWvr4SvZZDkpD1RdSn/TAeP4
gZpPTIQdKvdc0VwrEqjFxaCGpaF6KATCp1VOcnwHDx6KafqTCrPupwOQtJH95IiUWafK7mEDiIoh
0rZl3jF5PDBh6t2C3ZL1kSMp7w0Hv8jWffbfq7KChkp8svDZwLpPrlRVzz2YAb4sxzkfsx4ri3Bq
0hL5YVG82gYK2Cty46RxFuNncDPOKzJXtuZZ/GiDWM9fexj6A2WtmpF4wkiv1e4ix5Q9b4WJtvtM
ch+upfXTLCjxUACGKmrkNyJK59mhaVNuA7B1RQnd3oIl+YEdOF2iS7GTlk9m60EImMSZ9VJ+tw+H
Z7u+3xtDc0GyHBLrFmRBnULXZyqzj1ggrGa0ptca6TEBpAr8nQcXKBfd36EbzkAvDhsZy5bHh2tt
INGr2WRDOYmVFIhraIa/NYHj84/dVQ0K1EAKF6lVYHx4/C0feWbkSxzD7L/23hDsJgOJ1xHc+q6W
2K7dyAdX98D1Q3+NQgSMqPhaSsasUp9oosVoy1LEqqdVWSzvEhnUj3Zv06n4n2D6icyoYBszATwt
cZVeoWf0Bj2hiSBQY7lruOOJgEV4UGOqoet+0i5S+6ZZQ1sBtV40T65bjPLEoEeNJae2uxUO/K+U
lwiG4fhqrlPxlnrltcOqZnNrzGrovFfdV3h0pGU2Kd5kUJLiSGmgtyPhXyw33IN1bhkJPdf1CfrM
R5OcXNyvrx78Ca+5FL8NIchd0b5s7Y/qhE2pFMXVUTJ7YETClsg/XSNhrxnMTnQll33Z7c9zIltC
PIsTzC7rJc19Lz+DnPqRqaO/ayndG/7fhYGSIeiAIeA97GR9iQcTh0sGGAyrvY0kCpW45ZSpasPF
r9tMggPF3rK5cJcj21hueH7FxZ1TwCdqqyFBGsB+2qqVYsyBap8f+wcoLfxp+6mS47SOt5itvb8c
alTYO7cqf2fmq07Xy0UgkU8XQdUM4Mg9MhD616Zmrmt/eLFyQ+durREBy0tMKBzsh/6cz/43efq2
2ARH+KfE46z2WSFjF1mkyOsQ9cIBtr6yyWB8zGDwgZU8Slz3jLQdu5tV+KcIRODCs4edjwhcfzLC
+ELQYIZXWQPU1qCbHxLk8vQNKDFa6HxuSPELHdyZehS244t+SxcYcblBsS8RiluuDKR5yB2eM13l
0BornwwMReiiJO1s6R39BYDwPHgoXNbEsrez62M0KaCBmIaGTk8AGIXlUQHwLiHPxn0MSV/3CLE7
afS8Y4YWR3T26zebfSBn+Q805CbDv1WRd6C0sWXaL82V/htPbFQcqd1Zg4oxIghsIFPeuk6hJp/S
Ud1qFoAaGr24e0uf4uZPOFsWv6JvQ4li8bBtWjzM6DmJ1ZUCsVyY+E47Ys3uYyycpra4XoSblB47
y60R1s1AVNXGxzSZKT40ezGPvZRbLVPHY1GMbS4KREJUtsxGXF94LiN6vdAU7muNBHej7RHc3OH6
L8KD5Wr5CbXiotTEQ/TOy78yCkg/ASt1LFWgfaLrPT3heTWzoPeZF6sYmrqSD1ujDWCs+CJYB5/G
9D/rIZcN9G44UTMnkJXDqF/7nSJfK7TGfu7Ti89oXdqQwMrh/5wI/n0moBLeYYwuB6X60oSVvtWn
ePx/sQbQkNLp0zHLxfQXUW7Qvbf2qWmo0QWCDpcHjYGrpxfI+Sb2Ws5VH8Iaxwpc1lZxjzAF6a1L
w6a+C+Xsyggmuwf6ZpNUx0MOscwyuBc6SBlaUnqcywdigVcmWc3mXqljbyEuzOjUhbF564RQweYj
4hVRmaREBAPDufA60hGqfBh2Lk0lhfRqoPjlNWKDn2qTXFJptWb50BbF8vcIHx6qMgnWM4d0Al+i
XSW3S1ef8hpkpes5KAkPIQklI3qGH9mhG9MHMYp0QcAVD2OdeWJiMYMfwIJaMuqQeGuVJIokyDUm
Yg0VwGm0P9af2wPYdifulEPXV4steTjduo37CJ0S1c88hd0KEpyyqOOXs6GVesnxEKiSbmr2UWRt
MGSmM/NoAHIAbkbLM3TBdYy2gHh5/TNeT/CjQGC56K00LpwkmsceZx15Sv3dg4/YAwT4szQj9/9S
TrZ8kMI9mJEMLJVuALRVxrgfCc09AGtoFXQFXIHM+9BuNmkUyQFhLRUo0JCOkw0DRNOJuFBHoSq+
fN9dC7pyIbv8lQH3dn1uq++e8KgYzzHOROBA4OXfa6nPx5B1/Vpw9oGQxy2PltKiYLqmJrPKOmMR
imySPgXngQmcSeP3KpC/zT8rKP/bKUNUCdmJv60yDK4yWVD1REfreApYWEcbz8+hmpaPJ2Ra8+rh
d3JmM9DP8i0Z0Q1BeB+WxUvuPyX+VTi5FyxaMNOrgWC+NlUnXMI/z+s27myTvu/wsg2LNbQ2hZQg
vOytmZIRq2D0Losp6KqGFL0JTVCAbFFI5+XLT/j0n4AU26qz72lr+sfS906UvB8Ow5kFXGiJ/oTY
KHgkLVVdGqLjNaktT4ylEETiL8rfH1/qvxtiwCfSBpCbegoPCRK/Q9gS5G4Fm7Ps6dW5PBPG0h27
cG8NSKWje2opVYqgU3zITf3nF+bHGyvkfNtpEDWBS5DKN5N1jTKrTnnskgUapU6vnhShvoB3fKMS
5w2LhzXUqxRd0/W6T0wZgxoipBMPx52Cb7VD3NdTnA+J7esfpFEuW3v8eY/sjqTgsF9B9KSx0aU/
8Aus8TJ/pdlXhSp3tkij0KwNGAKR419yZyR521QeD00jWXdAqQ5aHZY3QG5ordFJSg+mjtc3upV2
cf1gvdsmpD5yNR4jZz7a+6K9Zp5HJgDhrZSRZiewgB4pMYlNlVOLcffoRJ0gsAUUPxkBMuCKM9Kj
XysNhTe1vFVzHRqDXgbGlkCLywJU5BQ2E24dK9QKR8tA0Mvh6wgaig4bINvWxD+fVR6fo01QNoiY
vgUKtzChXohAY6eS1vRQ6I1PVQsMRTk2PBa9q3wEZNFGVxN6FD4DQxG91gbtCITkMnw15rJULN9o
kP/lm+LNctdjpmYYlCa74817KL9uEuOomDfrRYGuhyHtzpKA7qih/7OoDRNUycftT8qtVXeTAJyv
xNlT0LTziRErEWNxm/6NR2knX2X1gvRpeK4FhlBQU0/qw1WYfXArew7uC6y5COUExhCm4xx2kCsr
l++tqcuMg07sYCZiVZovNlC9HIunUksfdXg1phRloXqn4NF5664tomR/6j20ZVkZUh4tIE8BC1jW
qgsJt/G0FQIlNkyzNi2St5PU5spkbmSRBSMr4LsbQDoMhzDAbLueec7UR6FGPfv/dDhDNIvWbT/1
TpxfkElN7A2i3PTdqMhHcTfqt8VAO7KNKj2LtPionaFib5cSUVld6JqmGpfU00DKNcEFdYQ2DKK0
M9P+H0LA0fBsXXBG6XB0bvSFYYL6iOXWCPtdVFeJFJEjuAaEsCZ+uKk5DDZWugakdAABmfDvTz2M
s01iAW5Mmh8qSUHEb3DDWRrZkJnNVWUwNeJ6e5F8y5lKbtm4TgPJreBPeB/0NdrJs9fSLhx7ijFW
gjqL94HafVf/FEAx8IsmorVNHwUwN5CmlO3d6SDgyFfvcd+esDV4ZwzJPq/s6xZeK+xl2OWdxkne
gwBHg+1TEphTtSnq/f5Ni/VaT5p1ql+zg45hZ+p61xOPCnZKlyla6mYX5WYhm1Dsp/OvK99xWsfK
X81IJ33X2nkZjvg8pxDzRrK8WsWCpypUUXO0kocj4jhWgsPIqA35mrvoEKPZ00JF7GOgzIllWrOx
AATflJFvOBd28S2PckgKFR0bSpiTWHMsbt6ctjntHyYPoJxHVSsRbduIV2jGSFP9rrxvxbd++1Gy
RmUhn9WflqpAwWzwmfbLTw43XnnEIOIDLIThgDxrtFhmh3eXazSsSuarjP6X5x1D+4Pt55YYJuIA
w331AUcTmNzI2aTj6wpkW3KgK2Dr8wTv0rQ2dXyypCILPxZl3fLhyYiKacKLeBhz+N5vaxHS9ypC
O3xPIdctIupukLhqQfYmUwaryxxtAVSBNsg9xpdDYoYVKXIBAWAaTV1OjlLjFMAccTH3h8lctsC1
nYSpklMPxgYvHm18evt4UebXXkR0jBd2tfs+/dq1kdBPRfQZy8R9mzd7lZ+4VghYSvG63qEsOZGx
zeBSB5OWsvamBGKpagwl8HGSWmNWRgU2bg/JbtFRX9BCg8pzdISMILRIm0AkUkRWap/JBZDuPNEV
KTZWXBenOUUgkmqcGouj1brVYIqPZbcXVyVAKG6BIoejAtOSqLtnLgoIQP9Iigl6GYYmb/O+RtDB
hnEXhrxbnJyDXNdXFefko1ggNciO3D7T9J1lQaQO+4eVws/vs+cpjKWj+lzm5U6rz1t26JqK7mdP
Spnen12+Du0/mSg/BgCCtYJK1abmMEHkRHOozPo+pSTs+ZsUvVi+K0UM+hURv9iE1wERMz0GP8vE
mPysZAXmflcBcBdyrIRVa7fmuWDa2YJbeJv/E+BFpLfMYcuJEupPyD3WQDPp2wVWWRHZWtH15GKU
sBsLbFeakvcTu7PCdwjqnucvdGeNI4IFIL0lsM0eJ/P0xJHGqYwK294vGMuw1i0yk1AP0kzta5bE
kAHRTxqvj7BgqzX3bqpv7PB9GqaelKlMcB2B+Y2Ntove7fwhu6y6DXfIC+eRwJ2NJjANOG9n5iHU
4lY8ZawWWY/xMBRsSFwoPwr/3pe4lrgZSVfil/yhR/cCGqDXPczxAc/1DXtxhbQ599ujt3a03xve
Ch+R0I9IXj/N1/VvpBFiFIq3HLFobvQeCO5yEpWF1Agie3frq/ivLDDac/eFWqx/EJ8rCN2Jka/9
TxjqLRP3IhUldM122YQ5+R6o8jrxWSblrFyUDurIQdfq3wTZCLet0KIb7WYpMlgbm/ov7y3FlZPt
z+9RsqBGgRtts7noouOp2Eh4Y5+7cfysRXUHiskqNoyzKWKjrbyQ21hR2Hgup0+Lm6tODiOtr+Dl
7f1X5d+B96TyfZ2pZ2fZF5/A/efkq6g7pGCoqv2xZmNk5P4IQCwsDGKdMGpUmOUR/QoG+b5wtqec
SgcTmzy7uHeb9L283TYi23/nrzsui3lxLNqypMLHbRwEWfLRDXhwPGgjg3noQKoKG2fBIaM1PjPU
qnfxTafJ/A7LmjIqLZu6nvd42kexOaJ6L3QSDtOwZ2ZqqNN0NdMOIzkA1vCVrhnLox1RydWXBf0u
Kv5Zh4SXjNvtzTQjPSt26xMGBajXSbpPjU/wmTJskaNM0gvwiY2rUJOZaOPWJPu3jxLfTYbKmJP2
wgPpRlWZa1NCDqcxcsmJuoF240/br66tEDcf54B+KS+VZ8wKgbnevgkkRToibE7OcezFqADfNn6k
XBPCTIEOsJCbOvbiLDVtKi0n9vlKMADYQLWxS1unYP5XrsGS7p7LKkztb8JRXozUuWOWGvURDkif
uIBJqZMXdrjOjyzAYHqxwkKytqur+ty9eKQjefoNwjdrbAc+NIjBlhl9AqaPmCM/ZXM4+/kGfuC4
y1+JSc6naQ2bpRk8OvNkLmrsCdoDMYFbDkHRjV+2PjM69gtPZzUk1M8MudGvMQ0wBYmKBVbl9BLL
6UwXuXnp+FGjLFX7+n3uYjNXMZH0LJMBupFL7SbEal96cbN9uz1WUCPfzGYuRq7QI4AaIpmcqkq5
qxdG9LlNKQZiP2O/JpJ999xW4NUGDmtCn4cvDvFwbUC/tFynacT+izg/PMFItC+rm/oJMfFBwB05
8rZGqZg0SG908+1NnowdbK2D6aTJ8B+86IUOE36/uAriGSJYBHoepZ5QVi8Fl1btnBIPT5Cciy/R
EVAt0+b9MoaoCgwb4Iaj2vF90EMDCepTwtjSkAqpDwn5XmjuGcKI5ISvA3dEaHbaXeloU3FOnqPY
eH+BD3627echAvNKMFA3bH3lG+mwmcytsNRuidbNIMcZmUT/9IUzPBLeYgrRtB9U6QM0sgxr0WRW
oEqE2yTcU6auCGZp41dDMhm0NJcTjAfEsKbsC4tb7v3jNXl+Fgl1pO8yKwG2+bSXxe2XL93ZpAUL
AvGwp4jfFa9F+efpvD7S7Esa0D5gEsUxkbhY3HfsyPOYufj632rgtKlOA0hkCSLxsJGxgk21fP5i
FciNXO9rKwXU2Cdxylp+k+T8vSVY9NkZ0jO8Yo0gCayxeDft5UKNSDs1Ge2jAKhCx6U4MO5vqdgQ
spHmT0GsM+921qgRJtAyK2rc2kECCDhAEY2KWBDjZzwzYJAXm1C00JCHMBSB9eWOQJpNT71a/GXe
4y4R3YNcb2bgzzROZmCTzb48M2HMC8k3F5vhwe7boBNIIRYFHAgU0omznXsfHKsYBwq/QOs0Lhvl
+A274U6Hg1/OoCG/DPpjMZglixUc790hArtXpfP0/4iCqW1goI/ZGg92/Fw4m6xiCKBsHD5PIObn
gP+zwUw48AbDjnrhcok7dbNzh2Ile+kD4OiqVuzj2xuyzZRldwysbA2nREZZi++IxPxrwPJCHEcV
HMFGhHjMO5b8eEYlkNnWDWQLDx6qOXmAJHbIbl0jJFgg3cjKejlb/RRdVNKsvC8jIxSrUvRRy/jZ
bWsARuJFOn1boajEGgp9vjOghllpJ9NayItb2S3gHrTgFnFBk9x1xnOcuzCXuZK+N/gy7oiGLsOA
8bxyf7A/ACZ+yD6hYO8vm/wJUjN7uBZitVkMX6o4a5tzOSIsI06jRwXWhxwz3GT+28w7fyVIE+Yp
NXaof7iSH00wDVzFeY8wtdO4VMj5Fe5c1fdBir8+gPtlufacDS9Z3IAz3trt5cyh2rf6VD/Kqryg
UgroD4UCfUzEH8ctd2j2ZFd6AwRMXwMcksxy1NW0EqA2weHWuIHlcyatoc5CLTSq91bKYaTjLvxB
2g+HValRMYl98JEPkGnbuw1VWBcxYf4E09QcRdWLgfHvl0tAURNdJm+eO9iIjQTZAP+ZjnWEcGXa
5lhrc4GThjy6YCfLK1iVoH2nx06/Y+fyDgKTDOBPk38URlUgGYls3gM/MJQ/9ex2sPrpyjfK179y
8DYTRWCXENTITOrLgxFmFtfsPs1efSYT3QeX/2k57XZA7a+0VcaEZL/eltuAxqwCaAdc+/6Rj2/d
leMVHdzWircqxZx41zhzwpr284bKFe5jm8RA339hTA6SO7p/+YK++EesWXn7Ap/ypiHq6UBlVCiM
EP3rkTUELWKD2ryEsZKBzk1SjDT10XXULnTiVzPH/jR8WI42cmmyLipcsFXGPO3Z1e+QXaUhgz/x
8FVR326kaN43scdpoLzx9tLQlz8RQmznjH+Z7Jy4m15M2YTsW3SrjDWggZimEbg65TowapcpSzjG
iS/xubgyNYR2I0O7dVSneWvH3lFCaoaXr8t+XfIfY9CtKllwiRP+ba+h74vE4pmfplRl1xhA8Y5A
oQlaO/mdoRkh0F74emrfDMw5V3D/BiCNHuRQi+UJPHx8UFrJkZ6ve61iDOajpvWFTPU1w+jkQkVq
gDk2Bngbhqa4LOw8pQayHn5TmHIslDVLpfnGGXyhPXynrDuvEqs/BYt4HCeldg5XcGx0fE8Zi2/p
m1vkoaEM3C9vlONlAfotPfPekcXRAE0IAIZeM2wHbtvVEfJpqEatFH1Enty9d8XE7aP0fpXzAOBT
rsB1SFt+Qz1FcjJqvBOD2B1iq/GUzPAZ5eFEyBN9Io1JsGdJUx4Qko0FqjhzwfBSJbwTauLQMXTk
AVtCNKZ6fwGSIzQJoyQJQ4Z/6/h2lp2aQOdi6BmL0B9yZnsoNUaXBTQWogOd3ESYBgEgupEd6lOE
0tHrohOsj7Y8DIzvMnVVdEhkXEuoyq0qKNC8EKPYcYreTm2amicZ1OTrrp3hUFmHbaHeI2cIhinH
XUvH1/5UmdC9oh4zpC8JiYE5fwYb53QDrqfBPQTNgTsNl+gXY9jC+FKQQ81CPZC2LrsUXRcQXelS
yQtV5YK3Y9tBLgdyflZkfKgOGIk75/NP8szFIHOB3KlK5Wr128LiQoO53f8eh1zKr9gb45v58UuB
JcSq2FvFH74e+W7k9VdM5gXzm8zbzQrbly0xsZnVXx+UCNmoe9pi5f8PBnEJo1fE0SxGNT2Wtw5N
shYKAG0qpvpqYQUadLzL0ZpKhu+Rqvrnor0DctqvgzqDm1Uq0yZKM9YFKm8k1BQQWoJhYVxEykbD
N3oTX5qOPug9owkJEpmdK15gz809ky4emV4oFqUJrkq7OmBg+Z2m8xivZI+HJq/Pm6KQIVkgP3bY
1EOnGTtL2h5qT0oLZYuuz2FOeWfL4UeLDjkbD0nA/ZCYNyqnwY7XozscqHvLnanOjPFY6qiycIyU
D8NYaN0ZlMTKNildHEfwdxHyHQijgjtXNcK14Rd99WyfioQswTtmxvdWmkXseUPfZLsA3bmZIbag
Gzo/pOP9toVnmz1eTOdGdGKlCtyoufaBAUlvNDAaq1gndufvO7u3F6RwGf2TuNokB7773VgXNSsy
qDRvt7tDtBI1z7+XQPkDfMvCe12JkxUyXzBMQeYfx88WeBulW4VUk+kBYZk7bgyV+4igaLBoF31+
1ca22MpR9msHjXtsLwcPzQrcPqDpLC4jxUIDnL2jp1SjJsQOoqlErnmTknsbjORu7B+gb9MW1Dkz
zShZQEE9pF3vjfDgB2Qjmj8V9FB6Bda2GljyD2+ZXWmke9jnsk1Aqd+LPUQ2r6WK+X8KxcrK3TXd
pqKSsHMmOw==
`protect end_protected
