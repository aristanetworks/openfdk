--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
V41Ltr8/F+FjIX06ueBU4gJUrsILZy1xdiVqx/xWYdaLVXEU4yjRnomWlHGY29whR+b2FrtlNmb0
kXcAGA3ID9IoF2OyTWs+5lYBpLI0OEGrmjOAseMMnEbdqfBOcWeJ2FDvGWO0HHBE1kvw6ybAeBJK
2U0R/nohtzD2QLhal6shHvY6HzcTwUIC/mUyFIMnEglPEhSF0YL2i2rrqPPhRXbMFkQfmbDSso44
Ummic5JOalpB9F3XtnjQoTLTgeGHeZuR3IZc7fPWjfkpzu5VAg81TMWBiGxm6n9raaHUUR1Q9hky
VPRoWoajbhlJnBrw+tg5L4min7aJQsg3r2aM2w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="H6IFpkxUM6+VYnQLJJai0eaWU1IdyEjrWR1/Fr5OzgI="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
NIZed3k7P9JBWQxiY8ZdxbUUt4Z5p3Cjs7B5raGxZmCV2zTZnEaBugCajZQer+dsGe4+OGhqfBrq
6SV88OwQFrI8hmQTfvjmTqUAsBHnKxeUeKrjhQGcCwVlpBUWSc1YhFDNLFiB67BXVzb9XaQd7xoR
uEEiYz3WL9FxYFT2vMM9gNAQtyD1AQ5pE3jtrHHoYBwLk4Yur8x4FzZm2CMR6TLsqeiq6+fhBMJF
q+muCv65hbWtZtckzv9RXgvcbzkCpjgm4Ns5rCzpUDCc5VvjynGXyF4S3n3jWOemxg18hsRgT6lh
y9WVmGnxLs5orAn2rb8wQidnrEV52PUriF53/A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="uEMzMySr2+lL3RUalWgkKQxZ4uniHoHrSu5MmmLvRlE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17552)
`protect data_block
ohwMzN9hqskaxH3ICEg74+KwySAROgUyD825XaVfzVf1UBDBxY/wGOCabB2YrGvIWbN4C0pO9ZCC
sZ/lfkuY+ouVxpp5k/0h/1lS7k7M/1XKhVFWBEqX0f7l+EFdm/kvQevPmAxMnzh9b1gPGJXeMw3I
lihIa0sooU9SuUml8COup5aoe93DIEoN1FeMnLXzCr7+aLmbDoCZvuuDKa6VdfxiYthxj/v1emaj
gaxpGchUfonZdjc9WGSbzbeExDDW4fAoEt1an/4MagmXGwId1q1iJG9pzUzUYDKlKAejGQVXZ1eL
6BCmypyR5JJV0c8cVkdfDtGAasRtbW3wnGJGISaiwrIT55WoOc5EsWna1HBhHnDE2gPi5FssgvJU
mh4+/8M30HQ0FW7A8X4WdPqyLEVdXb4rJfhhDYT21rBAMk6/dlXReDRBmmEaop4SEL3Wvv4CUD7f
eHfXW8ceNavw7MPjthqCBrj3OkZtYj6n6LeFTiwKqjzmo6/jgTmPhGR4kTJvQ4kNM7RdKmCMnMei
4R26i+z+PWmMqE6O4g2D9/hvbsriZfABedZ+oOKSsFmtkV/4Qc/ASRCZqy81Pr9xl6GWVdXjtoFP
jjeSzQYP5Gy3CM11GkcEwGl4SYJsNVwv4Krp/tWdOWGMG6DnLRt2gqwa8zM4vfc/VYVTGRpXxfIF
vtzzdiN2bP8dHFsT8IYoFl9FQEROFuvK9XkVb4cmTmmau7m1ObduvCYroRvmtVNT5S+Y69SAEz7v
0IfzGE4sdQEZrceEXjEYW9vBb7jZiyJUyOXH1sB5bduFf0bCFDcPAgAEja8ydEAcqhjTcmT2eTXG
i7vk5+q9SYfmUM9wlkGpF2dDtIZwA3WiPs98Y0aDhMCcxNLzArffOo63N7sKSTUr0FuCdWOvcOAA
3ABx/4LyvF7P6mnuj20SwEjvPMyvuOHYMcqzkf17ldDDEy69QqvvUkItJZpWUlJcyjS5oVLDcrq8
Hbhnc0VeE8/hcK+UIIEM4wGVrqNQMl6yVAAX9uZd0LukgPxXR0Hpiya2EnXOya8YI85tquc94B7t
07JnkjTrkssGLxql6KKF6hkFvhwerKB8wrZa8OWWid47sWr4OkM3aJF/I6rBBbqLBzgQ1X908KTm
vPYx6TE93ItZK9sxF32IkxrB6EXG1aVCMrt1bHdwZH40obut0g190CZ6cVwsd4gHDRNtj6MX9XXn
8uU46qXgb8RYGikyaDgcVXVnBMibJuzv+3g9tGR4sB37WVRVp02rGoi6NOkEEyi2YvRvhJSSZqB3
5OATKDqcTSUtQJPKN0PY5IWlWJZpAVRDBRbc09inWkOBprgx83ibDAD5XCnTi0wbQ79ssNcwrPoR
gT7ulsforeVyXGCzw7XSs9BrsQm7Odz+0CsA4cQeAZ9p4IlMXYX3ovHFNnoRDuADNcXBrhFzMUcj
7qZlLG1rERtYMSortOhi0bIWqaJX9KGCFeCSNnRY+xX6N4WUG5THcAkh4dWCqMPwL0x1E5V0LKxc
J86tLVvZ53gdFy+zMs1okivU9VmIwZ14izJZ0TcYo8e8sc4019iQqhtZEFKYc7uoyF443bg2ttiX
m37JuoxJGN60EkNBkWQ0N09T4uyldihES5aPXoK4dQnQdiDHwBLY7rSZp4gj8RcisF/6SSi4VcXd
cmdA5uPdEbE+ODSKzyVS7UJq6O3TSqkLEhZdT0i1AD+2YLwn98SRqzCG7GERkVxKOFyqu46owSup
EXfe2XJMRFMlOyo+M2DoplowUc2wyIkrLoZig1W8xUCFaGdEY/RPTWnxRVPQ7pF7BNIdlzydDMcU
BSipAPM/3l1xg9sTDYjISVSnNK6cQIV/ByzEM8tzAesBuXrA5IAB5Fi6l4F7Hy71hSSOURpJmb1X
jpgKHSugbpeiejSwDrCeb+0itKiSxu6otX9V7N4CLK24VvfBZg8/ftdMx1WeZR1/TI8bW3c231Ba
/eV+iqn8sPwNKEkeLvnpW4tPkPi7zCwN7YruetZxtx4nW1y9EYa2pXcqhAqSM76mT16T7196lGyU
M9vUkVfn+u2lReOdVBYi6lGXvt28YExM8JHJbXgsFZfeCRSGuOIBmEI1dX0CF1r2qv/EzOo2ipfx
MJaNum5W1I9wv6zKdmZw98yFvmUJJ6Pj5cHpH+i/8qL/qymNwY62XHXxmRxe2C4XRc9v0mb96JEJ
f7s7i2WYVlE/ufarR9XjnCQ5frQ07+SBt1+BL80uIYIFVW6dG3cTP/NSEkoVVyz+ilCLDH4K2lf2
xvUWKrmQWEGCGCL/IATTMaPEvoYGBCrGyQEMxYF0TuB4LfWlVBFX/ofqRcoroIpVjOTIj5qGdmp9
RUCIAoYovvQ1aw+0U3yIBLddRR01SOKXGrxtA/yHxRsP7I6z/ei5+xh/yYbf9l7CShOWYc36z+7y
Qn8WguUzWHc991pCNmMhY6Mbwj0GWHx7SuzyVbL15cGHEQ+21WID5tn7rHo01svtWGZ2BtS6B0Dt
FqRzjfEDSGj1NItUKjRwot8iE04jsSAC7B5LSHfj31zizCAdVZCgSEYpOBDeWDRvbv4FcV9HC9sr
Ng5QcgiTEpmPu/Wb6nqEK3cUsHCY9QuoCvSlHoH7UzG6cZhWzVcDe7XMVwaezgfQPVIrnM0V/fgb
Up/3hD9YAXIUuu9RmudHYBV48/7WeUnDWuDDd+3HCPupHnRzxrDObGfonwI8OSeID4x6/XvUQ0JW
iDE9JdYcfwSUeD0djLl2RiwYJdrDFnj8wVZ5+p74pEv9BL9vDJlHvmBUt9ACjKp5rVzCnzDVQxjU
2AbRak9A7qfF9Oyx2BfDHLRRAS2LtsBoEDn5v9J+fScWj5CPXYclHRCbUb3B3Amc6ymCM7b7Q5Vj
Qg8OddE/RprQcOU1sWktNySAnZosde6Bsd1BjFRYX92K7h48C105FRus1/tSSx6UrlJ/cnthhq3H
7cB24ZYUzDIziFaEO3O9Rme9OT0E8GuTNaNvKTDvfiQ2YvDUNV6KR7bOv8H/eWSHYHkHm2ziFqcr
lrZDMkTABu/rweILzFaU4Muf8PSkazM+EiqXqWcRbH+xHQqB2KKS0CehTVf6GgaM+c84S429nuiV
xgquRCynjX50TZLuw3iW6RFapdM3QVTmqcFMJKyACyEPou2mOIkRhwi9yger7yf13Kac04cdgdov
c3lDOYtkvAcatllpFSRvrFCytZC52d2libwrcnYvfRmL8dfAyUU9ABn4ZNUXX/Md4sHWTBKhfIHW
1HUwppJJO/U9ohE4XzlnMrsSbxD9sVmByJMHt9w9mrJNz/c7OZOjf9jANo8FOjqHYdLUzoCY2NAb
UsHbX7Fpz5uwme/mIO0A6ZLquTC6DHV5yqxL4HXQ3i/+hlisVU1HZf9+HqPNrcaB9+hnyn3CsoKM
n0fPXnmJDniCWKi2OlIfWwJ0lVXtWJIWpxndeyaX46cLHs4OCtJI/k/2kDoIy/wf/X927x52ZzyA
uZFL6Kzs+8RVIA+D1yqtrCBpXZPfGMXRURGJ8lOm5MXH9Cv1CIWANP7t0jVsRzgmjCy250rI91SH
aHvMhngdTnYyZg+TJs+hoM2ScJxozXcjVh6/FWH975HxlwNw/hlcul+oAYdKPP7wd+m/F0ywdy7Q
OLtTof5sfThCBIDmzYaHbsPnzZdY6HCK+3UlUeprxPpvCnjwXgl2r+4PINf6X7lZJQ/D3y3Lq/MM
HTzXg3Onk08kl8WsbiQidGfHNssItRQA3s9YfvZ+eDKgppcs0CDRNnZINWE1SfMbdFZlTT8o8EyB
ZeStBM2ZihcDXIirp8kXBsEo93SkXp1kPp/MzDlQovsg4x9/OkOlxuHR8iISclNmt6aZ6+UvEA65
hpY32B8H5i3H4rDbQx1oADJRL7AQyMV8m7+0HvPfRbCYuwJSEkz2xDfk2g7X5oW9WJI9u8FYpHJc
mKcDPLA+NjuMjbCP1hDmcOgqZU2DnSRjLYAR3X5IlGb9xrtvhOZQMt25ka9NZ+u6hq+uT8bBi84F
0MyZXvW5jBn7I+H1zWkRKAfA6YDyUAGX9vMKDgXQMsWiBTwOe8sYF/GqMeVG+aUX6mQLXqloAFiq
3ZFmnFr3uwgJKsgPF/98fYC+dDjK9JdRHbb88k+K4Wxn63z5eqlqS7QknOxb0smNgURCO3ukc5aS
xWovvdnmO99XcQemVhj7qIRTERGWjEW4vtxWVbA2mKxWloZqzlTTzs5gwkMC4MdblXxcjUjyuJAN
0YK+taNIZtb89KRtF1MOC82XCfU9W5O6eFeP8x1Ci/e1rXP3+/BcMgHMBwjMdhzzLnKCeJbenVFa
btBJ/8j4FD5Pvqm3IiSi5g0wdXsz3l0f6Okp/LXYlFdkCF375t9sYGww5BxaUsy8FxMdeYMtJh1L
1k+M/bjnRSZrxh+GbW3DzsWTW/ussasUyf2m8vrjWRbSrJs2hdleZrid8JPrybU3AiK/CABSR90G
Kd8gxmwT+0W2h7bWyqNoaBn/hdyulB/QDVZ1J+j1H6Akr69QX9pgz97TZlY4wAjZmquCCR/2g4A/
3sECrgE8aFAQyKnDoasDflO9Qn04Pi2N4HSd2UOqnvTEmRLuIxvjEQrtrUGvPY6JskcCIYtVEEJs
xJvlamcEnMmC/YfLuRFbS+ANGxW/VsPEDGUaoWsDbAFA3cvMF+i0V6DS/sdEMIWC3BCgCo0t2dMt
lD18oZlBBqIsxvYWtvW1rnVRAJY+gzKqFLYm47jlDqikPz2nK706/50n3XHS4XgnlX3U5P2nXHwd
6t3/DvV7NYf/5z36jRldmVwSDIg2rCTK+gxZKM+SVx+qW7UiSjnFkHnme49lWVyg9FItOskjmQ5o
voggAw9Ptvf11fIYtkxWYKXwE+YGAyBDtjfio9ABHnxGSnNOFnA7ECQHXxnFlH+xwGfRO+CFZzM8
YUxvge0PxBsCg7I3K7hL44unBkxZC5UkhmBvAtLolcNqI5FaeFiAU6kwLVqA7iK1Akg7Kq+c5ZBO
VbiYKDiUhcpxDno+gdHjC0DRwmuaKMDeP5DQugpZhiWHsUYRfZe+iCfKNA7VybufybhhO9D8ZJNo
fOBK4LtSIFEhv6mXNdmb7QSTd5HmHV8dmHXnhc01+TzazhA8sMDvz6GWpQgnstDlkzQtTBlNCuc0
zGCtpkmfN+q7xuO3vGoZbZevinaFaTc2gRmL9jZaSPwPnju8+DFlk2Sx0QCGIwAx798w+c/sVc03
LEkWL/qLTuQhLqHdj0jHwxSUB0Drq1Km7mH85L5GatEhodsZJRnrflr01n+XGbzJVmodgtR8oXjT
cOvl/sNSdhF6o+UAT8q1N2VL9ca26fa6mPVQu5A5ZHHXoCmBdAJh0ZFP8pVEKT/7rxiykRqrC//x
Sf8CAJbwbOEWjvq3SIglPRktzj/sIQqQJ5Z0oIRfTGAxidZtAdEXSp+pVyFgmaracq4DEORa+gQ9
IOCr5A5rseMwGEafP4mbD1EZ9VrUDHDGh19wxjOV6TqK25TaVwL0Ek55A2j7ABP/4ubkndA2Iuc4
Uc56d/Ike9NybkDaLGsP4C2O931Os5XI2OUzSyjR/hCtIcb3VP10BANR3PyZv8njLWpeX7WJciS8
LX/6CBCmFbRSnlYYx7H/kWiNmxXfJaZPAdPzHCLqqD7ZggBrp027h43tlePvs+CAqgLVYDf4Ni/S
9TkB4/rE32THWl5bEsPXNK3OdxrGhb+M7/ZPute0yLLkvB/Mx2svFTGssAXaC6ybJpwHZxuW+vEB
qSEmsJ8ZlcSwkdWxEp+D1TSOH3/dUxqsVh6aixSA6ZkEPzFLMJxQQXrAT/WXLM2DEvD7cEfsTnzy
Ibk0shCWf7P1qnTK6r2sSv5lLKctcSn/x+42ig58itaVK5MAYRM+Ye9HWJp4fQz4LUPuWOy2xR87
vS9mRK5qMifmR5ZCVgdEk0wWsj3Pn88rYUooKSSvOfgdcGrMIdiiUORD7ZBac33WrDsG2I2B5B5c
NDqJlylPtSgtycJ/kbE/KDqsZlGHT7e0jixVVNYpESijDnFVp6PFEPU/MdXD5xBHnD6MqAK5uFLI
Z0/A/V9ydFO5YsaqqfTAWgWrYvgeWOU5QsgtUP7s+mZUdOgMtqMH/opss2gvPlY1LMD6EKmlBm8q
gFk8oy0+gMDTBxgyF76wHhmFzYuCut2yGmAHqKkxnw95c+zd3XatOLt0iOzYw8/olQfVfl3s18wP
T5gNpCLMtIOp5zn7gXmtYeLQ66k833+4gXEuKzxpgIezkFvhAeIGUe16oGonVt51QjFJUggCktxo
SD7qyManH+ox4cNH2qFpXu0M6SdK9P7aDJjDP9GNaq1dlcejo8lx+n7Od5lhLCwsIKkUbT1CEjIU
29bqGg/bHg8hiHx/Ux6gNBq7hV48L0MxS5PbiPYhaeah3vKq4qjOoCCIepz6N3+h4Pf74gG3hyoa
QafzOHMHAuQuoJn4tseXaD4yTcvk2j7jlV8m1osUIaPAPfedIDfkYAXq0NFhOpcoTI4e33dYR5Yn
6Bi0cvGCCyaP1sqOtcx+rLg8g3VhD0TRiD23yduPJ68zTeGPFPHmODrp/PGQF0R7JyS0V0u0+bBO
uFFPC9vYoHGQDawoYxnDJR5mZpgMW9qb9T2oquZgK8oPsn2RJIZw2O8XiofGdtFVz8tW8R6o6QSv
Xfp5DakSHBaizknseLCwPRdiTPLdUgm18AOX8aO4h8tXk6ModhYaUEI9CGfdxSwY2Ew06Lfs9Slx
RoSe8XEsPV/Uglf5WUPsJMIdgHrGna4dr5Q1Y+9vMyGtSmJhN8NdfEvXwjO3IgoabDkp8FY27yJY
whZ4XL9Qu+btxmWv3hox3mLowaKKiig2ntB0vWGY9gkwaxtwlTMInhumj2hck/bvEE8kVpLee7pm
i6DuSco43OwdcS4irNib3KPGX57aBkPnwNYdcRcki7vjd+iC78RYk597Jyn/D1/DCdgTHJommA6H
2IHQgSOgVl2CtWS6rOmJWemHx60GBzNnRjbGLu3QbYXg5UJECUZ0W7hD0hEHIdTvT9x3EEJ+nMn8
oAl4YzDUsLf/r+Ktn9iFICPVHouHL3UBMBXXDkQlWsrGm0B+18BgjNngxzTUIo5AtuHwzBGSldii
f78PD+LC+DCzTWpXSZLeJ2k7b7sf9qKzERzN9gDi14d1XGpsegRb2Dmwnxj66Qw1aLKdVdH1GWXs
60BBtViTthXvIucu6LxMwbkWaEXy/GFNvHyQ9RbrRyazU4kcvJI2e7o7anZ+tJ/84O4H4Ad7ZI7V
mhNWgMZ3b2qVGuUAoMcKRyicE89B8D3Wb1VfH2U1VPmu3ArtlM461TB6mWL4Zpnq32A54rOjOKzG
D6M9gv5+PRPN4YM7KLXLV3Ajc9dufXTrjrIwMNGuF62ldXZG16LAiRqMfIfriAwYqrscA5GMebKl
yxu9GkhCX7ezehzYvHYexCzSNMjKPTmhGwroxj64t62WlWINHrp7wUFXgaWh7+DJh3sjT8aSgfm7
Ebk3bfIzKMUYnJIUJlXjael+OOIR1gAjt+DgVBmCjx/BvDVFsA+oywn3PbUw1NsHLs9cGFWBVOOq
ITxGWOXDVnLdSRU48+v3N6usaoLjkZa00kb7b7xUJi/rmlHPn9rOLhrccuIAd5CYoJjSYZ4Vvb2g
xVuQipXPKoU97Fv/IW6+Lu/3sqMjrI+OKhf1zCjFpW5pG+FmxCm/3FeCYSwnQnh1ay/1SS2/Pyoh
U1syoUVDoYoTNjgEqNg/1i7RkpTzCOLHEDzz8HwcS0Ti9Ubr1jfUhIxQVyHE0X12863/9vLAXPY9
LmeXTbaPOQW7R5+AmXVaHlqkJaZyDGcwf04wxY7et68jGMxM4i/J5G/0n9HianjV1KIdYPpYWuXA
BRtsadzCDaQ7PuJu5StFCi83gp9q3bmvy8rz+ow4RqoDEVuggLpjeVGkGxolTw0OBNkgZn1c/+GC
6zt8PNKFHc1s+CVhps6JMX8L2jTq0IiCIKTxhcvonWWms4RfA+IG6Y9lPMQ5s6e0c2WZ+XTNcPmT
ZQXLA1yPC30hgEQ5tDHhBTKzDQvQWR4qtaMWdGL9ci822s1yIm+1Y3dkyyaATQI5Njt0r50FGb8p
6jI1/ZEH60PZOWhe5LuKfQBFQcu+iw5IordKuPcwkGh3p9IKhDqk8x0LoiqLyl/Pz0edncEIL/a2
kgjHLFTlBvuOlxs0inVx/MOcXlaBCCCiIaNsCZ/ZUFCdUTGRasiQGOEUp8Xeby1zuB18Mbt2q49m
ekTrH4/DVydpDLymzWbCeSRUPvwRr8Xz1pV9XmgFqMVsGDoNkshX0Mrr8HoRe5vRs8rzihkl9ZbN
uKV5iUqeaYpWdPumZiHT91SYzaxEObwERgrFScAIM5GpEQuyqweg924XqjSpYj72K15e28Tyxoqg
QI7WamPyiV+ntwb9xKLfSpaALhnYZ3it8A3GNfgNSIbGKVVlC94IGzwvDLqELOGrRIofwpm+4yOu
ce+lJAEneUyhQ+ZCuhddpjeXtnowuCNXrvUN4HvxKN3QgzRzOhNByMqX2lPf9Jrm8yt87ioJMa6e
Y3c2hO5ix7khPSHRwNyU2hQ8pF2OJl0RYnCB4jUaLHrRJxUbJqz15ZLkDkToreqosb+z+tpyiTVl
Z01gfW3tn5o8fuhdW10WTDzBEs4iJE+I85dbzHEYc2Gk0+jYj7F/9X2LuiiLmH5IxKcB1FrmfQ6Y
2JJHplHMefOrNjjov27FdKL17PWOQh7sWpFo8vEibgGXgW3FHtkGr4zAF4XnJbDNC8bsdOqOW4az
OZ3ZugZlHV0QI0wQ9wWhvZ8aNmJwsXHyVpPHmzhj/9Rjs8AMWI9n1cx/HoD/2kjk4nBjYNS+o/Pk
fMFj5AVooiX9pLL+xj4V2O8JbAXrYuHH4YJDy2qNV9JSITMSl2eGxkLGwHwWIwVTTlj9bsauFWw7
6/ynIm9n1l648ikVFYHo/poFZgHhHuIJ5A42EguMXQHug6F8WsyuFCe1+/3KrX/xpii7K1M08jKn
bCHS1/OXxyRO77RleHzDR2GyQpBXP1cAHQ5POZaxi+6aFJPLW+5Wof6zl5JFpobcj588a7LhqI7D
C5LLbu7OEi5hNg7jDrHqz93M11zue2cN3cQSoa2S9TQ1x/+kr8Z0ivv/ddt9N91+xrJFiV4EJTnA
e2Us5+66eX99bAkuEpFc/vha2ynA6m4GlNEcJ1Da674+F3c+UtRDxQ+lg0tbsQ4v4lfCiwhJLPJz
8ySbCZDO1+YMbdIk2bNAb7ddtvWZz87ArZdZn5mwDugWmr6I6aN4K83zx/GLnRDdDPi6mQBqnsqJ
Ikw7HT/h/6LwDnaAeEfQa07rlCyC1v4icyo1pLn6W9kkdimps6DJQUdYGlzxF0nd0yIatKsuWhfC
q7AITcQI2WwQWL0FshMtsmKzty5l75sFdxUzR4lscNK0QEJKrPxwYh15/UDHwxsZRqgLDZ0aKQNm
Ab4K6pPNjkLyToX4JX54eYiV9B8+5iqT8VvRj5hk+bAZcvBIXonoiPK0wFs7kXVGWof47npAeTCh
xfEpo/6d78ui5iLrBnLwapsos6F4NV0hITeKdxCJ9h17vWLtUyqa5G8ap9JZKJ4DZP8UZexLlUGM
UK6JRFBvapPWtVs5zVZyZJ3pu6ofU6GdyTLuKhl3KVzK3P9XSUCRmVsrvMEZyXDQBiJN3/jadHl6
G2TmNdkniTKVJgbUsvYJmFih0S+tDyGgl1JF19h5ESXXvOwU9CFb6eTFnmN0SmXpvtrGvMdgn7hF
0TB6LE7vVxgElXbAPR7lFw4RlKViuq9JiElC4Gck4nRqhCdSyfxi2qjvokHSXzN3WjAcg2vYO8bM
Ud/G9fqdMVuegxMZNiQqbGSd0NvxVGEl2hbOeHTmcdZ6PTUiLE2uHs1IronWvatnVNLwqmYlF20Q
ZYBryYtlACesSR8Gp06ubgFUGBfyLvpO2615lsTV4grs8a6tM58NVmVmc6gjytQhID9y7olZbAcU
BRzcXsgUNLe8Kz2U8eocn2/muczqRO5fKMK0P97clpy2SNKBS3iTTw8uuYEGgNZ7pcw0Gldmlu5w
BMecGoj+0zrXZPZpSnOvTygw2Jz9PWexJWjU2vyGsV2tDc+CfcL5Ti+ig9iZ0ArCko5zTqasIZZE
WIIlvvSXO9oqgAJOuq5aCSI3A/TnkkL+mTpQi4+hBt5eUx8+x8jN2V8cKe5N24ZaWvEHV/P8NWuG
uQA1Uhab1vKE9rMDZKQSTdNpn3mymHVIw3caEF8QNIHq/2xHe8xuXAQp6F+4DP89rNXfknRYbW2o
WN0U7soFrWu6WXXmAaovKhu2h3rmWbURWoApUb6u87GDoLRXUSo7pzjD19FEBy70UkeNp2MK0jsI
zh5ucPFOp7ibaT9RzjDY1Z2QVxKfwnrw+852sdnP8xw3Z6oPyC7Kz7cJ07K41Ld49yf5Lnq5abm4
3BQ167SHKQ39+p0KdfVeGBhAJeVwEVckyLNngHniz+RudiV2ZXXk6AUfE9EA6OHDkXxpTQvIr/1M
ci3HJkb4UgTQOcAxCX9aaqJqpH0b8h774cRt7qSqtQ6YKnsWtVST5OlzbSrqf8DNXBxeudQ9UxtK
wRmW6zSv2EJq6v6xEiuCn9EVKuPkLLuUsc9JPnJLlc+1qehGQvN68eXmlexdwJeQNitgXz5t6uEG
tYRFxxfi07uzsQr2sffIYIw+w2ve6k1mKgo4BFB8Nc0fpp5VF4OMNldokBypvvVMqyCgj+0ydNrw
Rx72VtT7O4ZhPj+kfiNILeIeVdsptNNa95UlV6ani5jvcYwBiuHjDjWv1U0hjdphlYYPC7leE8Vy
hNPXBSnu8COoAnlawKtwFv/pl+hm/Ci3DbEQsfhqASGls3g+/tfVpS01Uk0kc+1wMxh7pyrOIhme
poAgPnDv8svajs9GHVoYIqa4PAm5tt87E4dPRHHgvQz9Gk26EI5N4nf0hKFkS3oIvXl7nJzBbnhr
7XuAZMINxN1S+AQVnf5DBSd+eXmCR5pyd/6DEGXrAgxJDN1oC1XMAtboMXGhSNCm70EVCFLCYUdD
+BrFk910EB2qnytoYFmO0hOHKdQSRVO83vkHjLI+LuX6cDsu1E5ACxhK8U9fa7NOdFLkmt/AqJ0u
/8YgYMYBJWAtM6bz2L/x2VUx826BMeYKTBo9my0spSn70UsckP9gSbuAT/1C5RbeQyEV8GgIitC5
K4b9N03U13uNRZrxihM8qI20SPCZk5l9X7FHswQc6vMNDFoii59Ym97iL56q88+v9grq5ZyJZyc4
ueFAjGUjkgBwK/J8xMB8vTR4ve8j6nBcc8LYLiCDMH7pN6T5pr3FmLEoU9frgsMkM4xoD2j1bzVs
4KQwO/AvQOzqu4+RFWUjrffPI4mHWYfZR2CgIRJvL6ocsz7+w9TLMKbjbr8LAZaWvTloPB7yuR6T
TcFvB60GcFTralwK1iRBBhtYfI2zhf04h4bwlCiY5CJh34caHYOE8rXvN6eICyRGnPBpsrqBm714
6R4QvIq6D1BG4NeIC6850s96ZUSyGQ54mjBGoWdFeGQ/fWBrRpNP99xR5oGJDekBqkfz1OJf5k3I
qnQbWDBlHJjFgYvXNiNcnak1qRrl0rLf0v5mkQpBA/UWwDLvYLHXUS0cprUuDpycloPvyXC1220W
MY/hSACNOXFWRM0i9hyisy9/F9pgR+3kRGF+kPMW1CVtuWCv9dtEibNV0brXSUNvDK96hv3z5zKR
QhmDCRBRMRKvWAsY+9Wm9HQFlqh1LSn+CEAwsllJ/RwVaS9qNf8uugS/o49cYiJp6M/MdP86l81f
Z+Bd2DnVW6Waugw1OZI8DIVbNlESjESTaJPMChfSiGeZy//KphAzjX/FGocU1N+5swsWTsvck2/k
eBOIS9Qpznu2AxUEFq17zdsOlnOoeeEiXLBL6Xp7ijW8Z6e82YrrOASSHv8xX3LLjbalfqRsJrJM
lQr15JAr5hjMAWItQof+BSXFTCsL4Y/cCVEYJ5YWLfZpIrYQf/4fPNhduIa4WxSyN3LZAmVAiMC0
Xg+KQqmgeANEhzyS+V1dHg3cT0QlLpH3LP9C69o4Pq8sJxg3zEcJTzdSvMMNaBPC3VybNDxCLHRu
gKMKoi5FSP21w6iM4y7Y2hOM1jcAEYYyxcSx+qCxRWXAJM9iBRXOGA08ZCGULQVpW6sKFzpGvS7k
O91VR9GVbCHEfsEhL40UAywbEPXlvBwSNSBRLeFjpEvAUHsBHPNVq/Dr+qsZdxK9igyHmXel3Jfl
LWFsJ55GHji48YqOxwmvFTZ2hZhE+wVNW43oxABYMvBNHUBvXRsxVNL6SwgwHWDToR8nlRQ96pCl
H/AfXvubYW1t1TwqcD/ZKldNAiu8wuxR3vNR2UJCiq2Hn1AgFmsOFalcGXGVoS0j8zho8bMG5OVR
SQL4UkZBHGd9XN8H1eoAceWcsGBrwhJbTNM/ZRcBbDxZfSxAwUZUAme3j907p2qc6lzh0nEKPo1u
bdJId2Cq3Vhwl1gjdeVPL72I1a/fPq4QZr80VtiuIxac/Kvb4bWSJ5ZNTcbBPGBPrX6aTUU/rkHs
TX8PrL87Pfv2gkapJlUhnmkNalHQNA4HFoBh+LJrBmpCkmmmMqvYOnmzx8xjroKd7lWK9mbBYLoN
YeXhgAbkFu3avpJ8hlSPyOPqMMPSqC9exsRiQjpWzhwhMJ0zJn2I30I9N/wG8amfdgM0qzGM8syM
yY8KXxPZz7/A6pQvS+EduEyzw7WA0Odogf3yPEK7q7zyfWbCNFpdPurI5PrWKdL4Sp5+QkkcRC0c
35PmKwTTU1327XpLRAb2+6obMNJqQRm72J4W+BnGZ1PR1Uu+hDh1e6K/Kulmyw+AXmYmBrnet7oj
6t0My9ghp8FRcQ+BIlUDqg/4FS27WUd0Nbwcxe1+EwcXhoGwl4M1a+fgWBC9x4lQVjTmNjjORGSC
zaKHZoaGe3kE7ujfxDeJYMgpd0lG1oeAsRAjK069Drp9RQRJkA+qQAJtIxqmV2CSwdQurZUX1y3R
NXi1Ed0sRpQlDh/es8ROyrK+uAy56t9mX8AQxYR595Xjh6MSS6bleqvJBqkrd65tfDMmYwPO/R6Q
FqWFb63XVcfGS1SvJ0yVPRjE7amrPU7v+w1vdo5HYJ5U6T9opk7DhbL4QqUpIZFcSBlFTLCnxQ/x
X85zk51k+cmu7Zm+iZ/xuN8YxYAnvfppElC3BR+UrbT4yOTq5g8TjDqKwBF7FbmGPBq0n1FjY94x
tfUmYXVgNjjqQiAdaloILwSeKUT2CkULPHO26cZ7uRPQoVPb3d9Dsi91FwlNbix5iFnPNQ24GTgF
lngHUpaBbxJaBrYuHY5PJxzLTyDn1228K8nMKtVFFAodXgQV5qBfu+g7lPiGP89PPCHoQXdHLfYr
ZgeLvZzBACkr/oYy9xneBc9rZGnzhO5q+Dorz3iOkLKCkHZf1S27HIcgKrVDlfxe2BuBhM+YZDcw
8/TE4U9uHQRzsSQa63ufdSzBqga86JH0+8b4oy1vI3nyP3K5pyKny6e41S+XuEYc0CHXR0qdi9OY
Ap3dupl5LhAwWagy8KSDpuMT2yD0YxQrTKdy0SyIKHcgPLUELwcYaHDd5Ag0blbU9YTMehGfia09
ahRLZuWn9JNReOdVJ14BOoxGoTqforjIwbWO0A8OZFgGK5C8pPVnU+QgestPsdNs2gd1h3ndk93N
OPAuuVoiA5w058IgRTeBwNabAFLHojBwfI5bpnEKEoj81UhajRERjMdgFbM58StNW23gbPHZeSx1
bejZzX2/GhdvTTIXShEq2Lp4TT52dYFCbqEhU0jZVapEb2DvoFya6Y1QAceCiaX01MQfv9ZXacz8
5B3NHhw6TE5d//8HMKLGErSNWoJ+3mgMYK8QlOlb2zT5538hgobsFS8hEX60L0yQRrH9fr5PFzjB
8+Wsad5lEgG1vJRQeBA2L57R63Hgg4NdKmPYCPXkTGDSBvlA9SbGb3VLxPvJXpbb9mlwor6S7xS4
fwhASEHjeLjN6t88iT6Jt8iznMnG67Jw1L+vlLNxQK1tEiuqB+To4JByv9Sfw0MKk0F/zEMuvVxi
Fy2GEXclnfVWPQaGuUptnEmRgnXZOdNrayfuhu7JpViTGkPTrtUyEWuzhBcjupu/+Zfsw/ElW9Il
3EfnSxmd4eLeeoMEenvTPjrjeagpBxhJtCC4HzLDkcTZILCtcfnIstpCnyXh6r6fMmuRS0s7a4lz
wG2DT0JUDlF80DmUZEX2dmJQnfCNC/NpVAYXoM+B6uayxbXyjVNATL7RUKrCn65ab7w/VtUFYdLE
8mPbPESQw5OI9noZt4EmHCvQH02VDY3JyM2UxV14HQYkk0iwfhIHwCH/r9rsBAfu94LDD7zsQ4Pz
fP97EXFYAWp9hKY2NnG3DJTgxqJpv2MkfUqm7olE+SEm6UNWOpS/fNKAj+9Jx45l3SsBee/ltA4q
w1VWjf8HIgTgZlPH9qIrH6cjyhfSXwrEcoi92wuJ6J0ab0hLEDxkNy/mAdjBg5Njlj9DnnS1iGFP
u+n5QXO3LJI6uUiITnsMdIW8Ax65hzWOWqk95E8BcQNXzpwcox/9PvJJPIU4EbjEv6aGnuBzq9q5
SUNBys+m0pDv4un04tpsAbWqVREyL6rHuTWrDI8AMukJlS47KdjaOnjeaCO3qCQEb4NAfdXnjcY+
5qWPbVF9zBxhM7NypoFKmhN12Vc0Xs2mmofxusiNo8Ddfzh8wQguAzvpdyskfjZzDYnV9hAUrRn6
1Te3eODtly+xjJYH6OFVCEE1R1fRLQ/bcaV2in+gitw33caDQ5IjBzwCpjMq1I3giwocLHWVhamS
3J7DhqXsvp7wd1XLGDWgN3wQhHPEmJr4X9t7s0Xd9gyLNPx5/IbetuVCQM8hcaqwP7AswabpKW4k
4Ve5xBiydZTTQjFoxQXbl3OxgNU07ppJt1tTXpr6o/t5k1tL1DMF4Irs2SCxzzb8FwhkDhviUTIg
WmtPwRxioqsQ86mK4J6OQ3IvnKljTJyATuiIXdRHrKx4TOkk1itMlrUvNGg5nsIOCwRVhmwGbdzQ
9o32rkaxPcYbiv4auP3R8VKBG10U0LPRotyQnNfqhbdexm33o5ud9bmUJWaELXLOq4d65SjP62cq
whndbU1iEeo4kjGmre0/CpxD5kkxpXyNc1lkOcPb5ybvUoJ0zlbaFRPAAITKwlC0BUf1Fwfvs/a8
lg3FZvuMRafeQlC8fL+iLJSxFTDpxD75OKCgEgvViheun5F2t3oCBj/xPq4efBPCYn8bj0ODVH4a
g1SsoZJs360oiH3+bv79L6YtHIjzZMY+IGtRDa/Pe9IrJ7Nhxvv5F0yhMgjdOHnddwOYzr1R9F71
T5UvQhi0B4w9YStYJlrxdJ5aD4eWml5VqREZUO0uqvw9muDBjl/1e7tOiBS3sqTyGESUW03ry5ZK
CNugROcyewZz2ftVVkyojfFG616F4mxXBnXD/za1V3ZYo+z3TnP+iDVKdCl9/QL/qKXzfKsLe6Jn
q1B6ndd2qK64p7gS65twr+CwoUqY63CCNp7xDxjOJdFUWVDReHT5BJh0E6mX57qrckRpayPf8UQe
517L1R0T/12EdTR2UzMDUEoLXbPAoW5ZiOi95DkxiORvqMiIbLGnddgMr90mErFT0sbX9oNIQcst
lcoEJkkYc1fqAZyk759E8mFHfkDpKjy5XmALY7ABhuVG6gklX/Rl3v281NGmg38V/sS8f0zoTPph
leWH40jgu5tgFjhhgIn7PCnTu4bZNufVOdsoA4z8rOjgPmmcPA736Zjv9bDngek14wReb8mcpTVa
UOObo6zKjkc39BIDqXvmjkxgeKG675WyfeaCAIatrwZTe4L+fc+1Hc6wQvO0kIjNqpvuYw+uLn/T
VooVxr6SEUlmQNbD9njc0s8IrmUVaCepNhQ0JHTS/kQczE7P+ixIKCh8eqKl0OgtXO/OGYrVsSwD
iGto13oj7/Iamalk2ZQTTu8Uz00aCPPLVhiZcj4vy3FrmhZBI6oicLhfqBK9qnLdjaTk3L2yh6+R
gI7D0cW8PLMH70KFji/SjTzIMbAogvhnwbXlTUSoeIIiqxxN7iVDV7YfJfzX6Egz327VzxP40wUg
XEJ2pHIhhuzJ9lHZ+8HJreV/lRuGiIMZdQpgnBYsvJR98IUXVbWwDkjyXRj6W+WirPvOyvovPRrg
Hg48hRr0gbn4xrWoqaeGQUW77B4V8ZVE2vE+l7sQS/iB88ATeB2HVBhJeiikpJLXG3Kh30hDbpSG
3UEMVJ8luzoJ3CrKN4gCq+sZEf3JMSDBorUxWD973HzA46efd2yz4zRC98bI5nL1nsUGzIJKK4dC
XgYUu4uBN0d7dDwUPdIFk2Rz/ne291HMHHjdIJ+x0R5FqnNd+ljj0uoBnmWiWPed0f7sPO1/19xS
esVs+VPXldYnwpDwRpssdvT03bBAh3rDzfSne2/UVlOIHf2vkoXprCgJO2SbyZQyU7GaYhUUW1ql
ze/lf7+t6UEMccUjkv7LL6QAkli8IzC4XgD5KZA3Ycth2ElRM0tNTAVDL6zbUOfFTwrAyQ580YVs
k9QmLLzX1cF4ips8t1kGRQhbLODgLY/WkabslPXo0Xg6VzMJDOA1njQEqb2qXdmF0RcduDWY5yz7
EcvgD5zfrXVSfx2zewzkVwt1+K8HsQsiBluXtVW3T69XlRwK/DJm7uSet6aJPUqJG0GW5hoeJZEE
G5qtpvay76imhVc5chgcQyOvSNt2bl9R2ShxE8y+P7I9ZLzvjCa7xq6LrowLqgSd0DxSwoXHAmiZ
O16JZn73eqElRbLhH72w9cADxEpVbW+8J7rz/1zQrAC4UBWCTNvnunUHJYD/U4iQr0FvTYFdX/YO
kaoJzj/MbqwBblQUtcdz8pUaRk5re1QP2C5bWSGprotUyyR3tYkBL8MQ4LD4BekAm/zPVUoWB9qt
K0gRAlB7wlJoEhHeUaxnWe7dgiQxjAFUFTRXoL7NZgu31HCpH5p4UlcMP9oIY2YQrdZCf98yiwxg
sITPsResWkiQu55dk2khkKrgyDOlT+Z6IMl4hdvjWsMISuSlFadJ/em2hayRt/MUz6ozrIElw0hX
L085BxkuLXuEMA8BzdH1mmHSxSCWofugx1f51ybHXsB0Xd/9pYj0kpEF12WRi7cVIcoA23NOjHx8
SWkPnDXPwDkAc/v1hXFPPi3UVgj4ZxRNqUMoYTqgDDf2i5jgyfKxesGep09FoeRDlc0F+bNwDVr5
UA1OWNuUIMbguAtkGQrDEUtXOcnLL3r/QPeO50YuhgoimFVBRXAgcwzMwqcNoTHjyVaGxxgBm+g7
guQACZdXuwVMA2UglcyydFxpsi50/VmUTf/sy/xhLIRgrFta8B++YrtM/jGDrGUf4plB/JMuGQi7
UcHaOjThX2TFxj8c2odlO5KGlqBIX/YuwjcCYFkk7DVirW3gr0y+JfJ1qc9P1w5ZwxkPf9lec2lX
3XqXFk6TyYHpLsT3YJBJtRVG/NH72RvIrOR9+ah65KNeBq/JIxH3p85Dd8AD2dC3UlWvtW56eZ91
L5/146klcbp+JK6ZPJuMHQOm8Bgk6VRLd4+39PIVC3r0K1Mb4KcH1RbJh+cn3XqpwjPeUdbGbzBa
DZjELhAOxrR2ZQAEPCEH7f1ty2ISq5BQaWGn8RqV22MuBeLCZ/jMuA/StFSn42phlmFxWkZ226cU
7BuzwyYu8q23WxFjNY5OutPGSB1tQkh8ghmQYC7Ldbt8zJSn1HKulSVCv2aVc5r9FjzWu7zKtfNc
aTU90Bn33y+9GZDIQ9ctUB8EofXrNG1b6+F975y20vGT4mgGBmY/AI/ORz0dzCjoP186qiHdNfgI
ESrL5S/evmqt3DIaDYiC/sRICamWbB7c5T+cZXCES8XnMUuRci8rqY2gt0af2ueF8hKaHiXZKLFM
Iz6SbLLrrTmXzHHMsCQlX16cDFX/reytb1WkTeUBDx88NPG+sSKxZ1ytobHzbOHh6wQVexGls0Lv
R4zRzWz0y2U2IwpUGfEn0W1vq8LiICMVRjhdcDKqnFJ4o3qyp8Cam0gSMnA9f+kIsuKgdbFdRi8K
QnosSVvv4FWR+nGbgJaFyd4svdO9IHhTzKjTZyiQBU3azToei8Z539mjxrhPmDlTB6aywhW1On1U
bZKMxGdM9oH0p6lRUqAAP0CSC2kBxKsy7a7SyVJZSIqKdFyP+YhE6mpV6pRQ0xIb1ZUwWK0jjdhB
Ut/PHUb+/g3d6X/uoemm5Q0oimpqhVgHz58yTGtCAG6Pv5rL3sMvaJ96kKpo8E3Q4tro4GbFsT8K
N0JvqXh73ve9Uapp9lD3IDzIAmcElc2T2aKJw8wg3qemKf9G97Ee3dr7gi3qpyy52S7ahiWduuaH
8obMNV5q7ffUXm6Efr0kIcXT+omPFllNXdzNKO1zQL5A+OOKmO08Wyfu0wjd8N4H0NBq4xAB/uG2
S3ecEaKlTYCCkfstfi8cg7cvqlQhYerubDVaXiqqukLBzELwgi3pWUC38/TgIbN90t9fVSLpeM6y
U3LIf5soWlqyD8oychNJJ4oBuIfHA7Yvcw5dYi8byOIBPtcwvjOvfdVzsVMOR7iyRCgB1XEWXa0U
BlwppbuLA6n1Tsp2paeBPeDITN2TP/pYPZXGKeVsUY8g55rIacTsH7PHHlCzQcVknk2rEXCf+2mc
zSSkHgZzn7TktYOJCPJaaLXe0iaj29YHdOaqdHwBrGV7xa8a8acYla4iU0BxVWWxvycTrXs4d2Ij
3xA+PW7pc5v5pOqTS1rALUV4bdJAUxpl+3/9bTT3NJ/Iyl4MFZoA8mANA81cVW8veT2DkAcjTJOY
XJcRLLri84EuugH6iuLxV6d0WAspKDe6zBmcUSuVC/Abbj4Zt2NmsAccwfUi6sAktfWjaCLBI3ed
66RRfkztvQgikpVI/Epe13IcsK/C9PxDKRsXdb6ce3HXk182a6Xnu4BToTYP/aa58al9ohiXqXuQ
nf8TxyCAVjptJQh4gmkNglqzjwIJ22V4g86ryTywNEdMVmkwtpoxhEQKGRZpArl65eL0Pd/56BtS
Bs8NMA01vKiHJfssWCuVnMDeohi73saxKfAt1pt0120cukkWwu2xHu1k0ZW5dStrns0/01yUZCen
FHRZLshf/D0LgRoQSO6Vq0/Q5QSFlsSHR+KZ0+AgBbtPSiS0GiWz0nL1C67pejgJfD38WExKo+1B
eQLSeRcxQA7dau6Bn3QE7EhNy2+k4QhpLYS1gIAZ3CRLB3R6Fh7iHnV/0U84+BQu3vDADyZoB3LS
ImTeRkwRU/n9na/BYcdFfhjVqQqfXAB6ttj/2XvHxOVWs/JORyuewbgFXgdXjWgy1BDUblMujyP2
TVqISdtYHMC+hT2Dujy7jSNxAMyGqcrx6A3AdvRk+zt0q0lRBjsFY08R3QqIdmEQ+YMI7TijpQfk
HyzcAAxCOt2CHqiJwdhrOj0tEhekvy55/7Lb7eGttipZw6PhLGwfkUYZUZve24KXONUs7Av6K8RZ
72ifl/KdNL0WKJqSsdt/rYXVWOUQvRftKAZbuKNAzehYsEDoD5s1M3ZICg+qaOd4c32A3P/p+HXH
nlPaOnE/ROzT9GBI3OS6UlMbA7WhZHSpExQovMGQ2F5IZSpErppTy6ErzCffk1uWfeNAnCPY0eUs
ZMVL3P4TH11tz0luwatH0NxeK/wz8mnaouyADCgVB4Du4XvXdDcy4lhvLTyV+vHfCihQwZmvY5HX
MLtpsuwrG5GI5393QVP7pUYt4VlDMDbBLVBzS9gYsDoj3KjKsBQGLDiT3fGUxO1HwkMQ9f6ufqmk
e720Hp4UVv4wgYSBkIrJRIo1mUVTXoDgU8I+xjxn/Dumyhrt/WpoM+B+rg9b+G2O7ZX3WTVbgTJ/
4UmcjUty6P32GmScf9QEHAJRfaMyLMfMsOo69sbQ7bOAsJm92YCSEkajEfJApufw+JgHY4YVE7ry
IhguR3MTAEb0XWaW3Hb+NlUF1FbXp+0KfcDaDz8cKzg8oIUXtTEw3lZ+KgmQ5KZ31BD3YfrSxrzy
a3xruBssG5wuRbVmSd5Dx0S4lJBFwAPHb7W5wtWBHxqoPXwwHcAl0JG1wvMWh5MKFdqkTNVsGBjk
mWZ4+Bxw+BIJRni/VLHtVHopOlviZkMWwy0aRrbEqNr/QbCfvycpRpAxXhT7j0eUG0h/7lwySDHL
J0cAvTg8I1VbN2Bo1ouoy5nE6SuA53KCmNtrRAdNUmzhmSI5QiDNf4npUJOKKcy/WfvYDQqbkJVw
P91+F453xyjSgaVA2ig3WmYMVaAnojG6++EshtVXJePDaBH4z3tA4NjieOJd3u3ltTWM98g8t/wl
Kja6o33X88bURztPu3cqbG6/fLA6epG6tzrf2neH/i3bznIf4ns8fXnCAxHb551An9sLaWqWt0NM
Buex/nb2DW18Fu0eVDIx4OdotDHJyxQMLCrtxPkxv+B8adJKJWRG00etK+7uNdXSTimZUMigctdZ
snOOX49X3d6lQWLJBCwzX2Xj8lwV/Lag57LC/GAyzcPfxOVL9b6DxGbKFrvc5BzWAm0Hmywf3CRI
7lpW2m6k0xR3tIR60XasK9L54QOW7ddToaGKJ2tvc+59xMHJ6FDytYPWohLnFIjG9BUU89r7RF8T
wK1WNg6SY3yD3ZE4DScm6ZJEQPtTHRKdghM+RibgKVSz9jb2rvYbFfUpxw3F16Hc/RUBzNzF+SwK
VTrtqy16Uqzfvb39ravNAGQIV/oD9CQdxu6AtJNZu14VTfGdzDsNs3RknQ17gVGP5Yq8r9H9PJT4
u1s8lwANlo2NDxZ0pFwJsY2gFg5Umih0MBwtbQulRU1Jqy1LKghTfwTn+dxRzhkbq2oTwRmxDyOm
68tK4YVt58sJcTQQm8SIB4cArty0ngzmSjHiriBF0E+PeDyqsxED9xbZL9bvKsUq2NIED2sxJNXq
IFggKfsTmciCVm0SVIwEu5iER5Xv/BaAFMtc2mVGFI0X8+nV9yxJblzp38wyO7PRIsgkRhBdxfBE
/srfLBJ1cRyM3Vzl/mkajApRyud0NyOZa0HBeVpuyDu5RDOTuErxNgtCMAUMSxvN1f5enxyv7xoQ
RNWV4/nqRKk1eb2p9nwqC+VSWiS3X39MOr0aAewczCkms/lotPzV3lQfA3jnQzea/9CniHqOgF6S
NW90dcj+uEtaiDKeQZMzch76AKjcTCJCi6B1WI/NG9dUg9Kr7RgoqYhOaxrT6FC6VO7j2NwdDUEg
nnLjAerpvP2PiGpNrh+gsApxZUOuYoPUeWf5F9jhvgn7SSJNK2RDNuVOjcpxFDrxAU0akNrZfWDN
4qQwyEFyl4Up4wYTexnXrBcVFVt+U2+jeloc5KP7iEvLlc1HGjJ0HOvNlbdnC/iL/uv8Jnzm7a8j
mbdXQEbEwdrjgxCN9Umc3CcNGmyz3pFKnCt1BTTf4id4+AW5K0MBHYZNgE03WqAy15412fV60B2U
LOpdgH1aVB+2o0Z1ROD2topzNRzuOADjfW0xdBA6IJw0PHqF2kf5xEcA/VrQ19d/G2Phw73eE4dW
rc2rfP4+gzuEBmXlA24aNXMs9+LFGcnraId36CVn/zdruGIur67XZcdXOq3LvslfhRNx5VATnhn8
9A8rytBTkt3AG1riggWOO6xvOlIZH0L4FQcKgCZMzf4OwHonS7jbKzLkbOsacqnRFLL4rasOu4AA
RE7Ddak6NG0N7NTuAsN/MUvx3/FjuZwSI+4jVk1AMrR7sV5UWwXbIY7ZepbkXuj/vgLtE9rGcHNH
ZEKX7rVptX9vnDLci1A7daJWL40PA8SiTZwDjNq9qLLAEte+ZdaG0w/HYR5hMOeoHim/siqyFPQM
YRh8EMBjxZSTAGN80/UW9KKt5+TYv5az82BJf2NIIADzAhTluCCsX3XKFjS9IiBZgB6g4KiTlXqR
AUFGZUM98JiRKAMCGD3xOZc2J+Tnh1Nwg9oHnXp8ECX3hr2bS0ode/d/ByrV2trvRny10UPeTMvM
RipjlDOV5MNM5wTXzCsaBaazQobxG5g3nWKFo7yPcqC4jJihDeJc520Xjw8fZMGCJqtiXvr3ATZP
32mO117WJLp/zmy53ysR+uYt/MhTXuXqiVcE/16bZnbLSCCUuhbdJ5E5TSgKCAzq21shM+MI4Zl8
Gv6cLPQoFQ40k99RnKzty8lqLTofuc6uO2qwV6KSCLIL4jzCLvQGCrCI04RFXrLakyf7iFI0Qb1y
fOglkLPUvcP2lfX0QOQnF7EasBoSECwMrKF77U4YGsv86/ZtCfWXlqaLFxkzVNsYPZMBBjqtEFcD
agUoXwlxYY7Ifbx2Ju5ONvurz3kUgOnPjXomLGAZC+Z+oxae57uRe8Wc/g17EWWMh8TSb9E5s/o/
Sq2fEhvz+Y8PGBMZze6eSghLgpdM9WZXk/IRSNHnCvDUCfZhDL/ZRV9JG48+QCEtrePOdzVRDEYB
m1WnX9H6KDFKeKHGco3QVWZcZbT9dVZLUAHL+Iw8wn+Xo0MIJsF6GlBfgUDJCQ9rOzzX0ICnY/6b
KLPMlaEJkcBE6c/zxLhbFwLcy5v+76c/6C/IJKBhcyG9hqcvlTYprqfJZffu2sO9zfShKDb2DeGV
PDnDtdKTEK3lrH1cictImOw9EIo0fOPPJObHFGqUEfQuSqx5Y/suBOy4eDj8IrmAsHGAGnOxC2FU
6wfmB+RyFbGSnTwJVg+2d3TdQk2rMd391XUPqcR64SqB4fhp6UaQdtVuZ4q+nU57uTNGXqPXO3Dn
6zPqJgpLG0lyBqYJmuahmxBNYOeQ7vXbFnZS0Un64HCYnBTENtBX6lHD3Kjd2ZNtDezKGMEwqAnN
JZTOAWytrudMZZ9cGV7lLnhWa5/dHqv6HK1krjHj85y4/YnizFe4g7r6BlU3q/ADr7ADk4vG/T83
O0jSErAptQsjxaaS7w9OC45oQSMclqqSc2rKF04nlaJrHjHcjHnG+WTvJuDkpzByAXpGpSRYLC5+
t18P8T2PSNq8VIKRqa7OuF5P6joRYCaXhZosyYlcQkeOjFNpqRpng1QU48Xpou/frKoHUCXG/6J+
wV6sCf7OxjAr/nn1RIpQ03xMQVZtzXpMAY+HEbDc7s9Zi6sKmsIRsGj3O6bVneBiuQktfF4lw/jV
9PY5ibreTFLSxLIoYRfWuKLnLHUNadeAGbYQl0GAJ6uFMNWLduVs7CjZfLPXgy1mm2WvPJwAiz0N
bAYfHegDhx0YwxtNt5K2kcQ0jmzE/neB2MzL8UAusAnJ3QmtfrrmFENif7FBzykBMduWpT0=
`protect end_protected
