--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
fFJUpN7JdIEfmg/gqbdxCa4okEoPvdLXXJFl39BuIuAVXdWE8OfRNt1UscIqaB7wX+r5QhD6lf4N
x0su6Am0vlBGdzdgbtno7JHU8+EKBTtXDMVhzSy+rHwPYFpPMMv03reb4rWO81QOROPPNFraDpQZ
FfTn+Tw74eAwyc2b6bNZTZM0CB18X4bvdF9Qs18VNHE5cCNe1O0aHHlXtH0DA6zJEsSV5STZJbJq
ef2HVflh0jQn3gOp03ZC28kddM0XvLNWD4XvxkyRSIsFGt+giQCq1FBVp4QMxjbgyODgtbnpsOoD
jq2MFQ71Z9sxSkNx4EseDk3O6F7s24mp5FOkmQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="5bbUGwnRFy9M/xUuF4lsl4fKGi8SwWJRLo86gsITdeU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
OOJM8eSnZ+g+ojCWdhI+RLaAMaMk0EldOmvxxTNLpQdYxpsVeyjR3TJt3Y/iZEcUYxIwd2c64/Wl
Ycv/E9ie8Bu0GPhI5lkaV4cOSxE2qfEXFp6L4W12aDp+VvN4OgKPqQckRMaeVv8fbKE8jDAB6E7q
lYPptJS9uNRbpNCYl1+XAuxhJBVaIy8wQI6VBYvb/SiBm+xvQWGdBjwdJvHKToo8VQHRMXWAR5qr
WqYJoKlQow8yXpkx+QJZKg7B5LqrSCmstANry34ZKhLGt3nitbARyd3nQbTM60a21cHXbxuCz/4k
3f5bL2xDPpfgcpA7vdQdCLL6oGMiKPVTLkO1vw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="aIQyFSyXEcTg+gAacrNpR8Srn0rVLjPTBsravvTgYh8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 93168)
`protect data_block
OroVme/tiV/rr6jUPUuCNy9Q98BWG0hgDvf+mky72csgdbeLy+zGRyhyZkxtLtl/s1Ikj4raB51g
ci+tR+sLRApJrgvRZyjyVtDlilVQKEGKRMvSVNiSR1tX8aCKlceEL/KxEv51sqtLbyFbWShPOTwK
N3gpAFvOlIMEOb5tE2fIyqlOVihbF1V5ng7c4cwMGO/PqBv+D4fOa0khFF02uqVU+feLusqIUQK3
ejCpcF0Kt7Z95f7mEXkAfDGDtuepoFdpxgCdzMToIKrdZWurg3hc7UNI+3ojoi+roQrxAKdD9lxg
+qjR7MH8uvadnPn/k+ikqaB0BKLHFDdHJqlVoxHn0mzOKy0sKbW+Nh1wvrxwmXah553IbtM1VZJQ
SFZVwnNQmokkq9oIGmT14l7Yfm5+62guruOJT2RSoHkf96kgjmnkarhGHyQNWc4qdQMNswTRKaMq
7SJaKMVpbi8YJv21gx3PJYqEMVxr4cDIuxSIOC8jsQ+jtkGAo61emrZCqvRG6eEUNaTIdhhR/0F+
584CTfzw84MliizJy1q2xhQ/jxmRRbNcBKBEor1xtz6iF9jE70tKY4+UwI++BSHR4feYRXtwUvK3
KJwcNyE20GXmotsGbc2d7Mv/mNcR8mE+Wh6lFEnEvaflg7T5FyXGJNNKbRgByv9n7tafW9m4T1fY
4If+1yef6YTV4cFSDtDP6H7o+gfJmLSi8wgCHgBVGMRU7M+IwGgXc/d0nqJSnvSOLEJILmXAtpo1
jHxKfuZp2ODjHRsPc6N53OlVqK5iYr/32XZNxNXr4YFZzy45fg3IOaWMX3tzvfd52aEmRlRZ2rF0
+AHowXX5A4aCwUlKjeVjdRLBsmthr38HFEucHU6DbjO/z/3YYhTbTksse0cERpl0bAfXATv9o5Xh
dpVcdanAk70fVbKu2CzaMG8zfnyUMBVo8pWcCSidAy7KeYHskVawrvEl3/XggFAULwT54dlr1c58
sySzXFX+/i/vUZiRETsxsGxdnoryT4V6yMZbIDgy7TzmHoZ4mwGbVQbbTeAdaxUdxRx1KcK2k9PF
ZE4rYl9kaCpKsGGtOU0ZvBuIhTMvLTq4J6XIFTXjpRkYAyzF24JDvP9YmMX4algreIAEcKnGNqih
wa8piQp55E1UqGCzCTExmttswpskpeM1jBYWLNIrp80KLAr7O1x+Qz85AUb6pijyVedZ+1PkdmY0
9Dl/VGsSfuHKLQ89PJA4/g4lQtsO3IZLi3ylwBxraxw5eZB0l0vAyOGfBJ+6kDX0lD2rKFxbeIIK
pwzcVUfOEnP/qp1tb2BiLlrAjOyXWSoQrGqdKWWeFLS/szT93TOm0BML9rMqgq2pHWwBUg/hNKEF
YYrFdsI/LZNSvdvPdhbxZIgNHHLZSDy1xuqmCvVShh1k40eqnUtukPke7oglpFZTDnNMcRbeR2tl
Y3k5sOSx0UX4guyptG3oBuMhQb+ruNo4fl2LMq+K7YNe1HP9nWyX+mXkLdDZ8Lm7FOuYiMtWENvn
DCU7Nl19aw86Qur6tvfGE889v4tSbRBSx95ZWHhaU/HCGl/5o3i9bGRRhc2347l5PGJ/3eh+sMQ3
JJV1cXdQyWMXmIwlrxHt2mTdbLG6Pqfsl61mTaoeCHL55UIAoz63WDEvzFCy4cGjZbhR0bBLMUi/
FwNCZMQOy/dqWr5myi1jqYfenUbZSYMQ3lXmaKUqes+e02lq4vfCsUr8h0FQtSo6gc64vzW+JaYw
DiIXBgSCjh0TemtfZ7CfkCXRuDyGNYBYGlcmAbyq7KHv68iF5eryY0HEsuSZ9xUrkcnVSE4Fa1pn
O5UZJEGn5L08R1/RZTpoO+bhlrv5GT2mkeIW1ChlJYeBNLUV9Ypdr2JRWePE3Ghbmmsb7g0hGzrb
9N8cQwCXc50ZKw5crvV6noRRQ7/JOj9L+mq0akuZhyEuJb/br9rYrngR7UxF/F0AFP02xEJPvfFB
5hBj7x1HlDmKE7tzbhnIROjLdaHmPmbrTR/EoPCytwqpJE5goEkon2x3AGlPkGWLkPOLvbrpJWU0
T4xPmfh/wCG1XZ3NQfwuQKhbsKcW85q0QFvnn98kRQh5WhhTFv5ha2yHpGLLtkLxlssKQ/7V8W3b
8YXi9klcVg9FXCp5uNjvz3qS5P96C9kH7hDQUxhxm8O+QkntnGnx/7IR1v6X8R1OaBY1mKwzXm/W
jMddXsc0kM+VoVpkuqBNgUr+5T6nodeC4NRp08kzgw5qF8rxjwNCVxKPvVryB92zH9WGRtokbPVb
/hG7AVIKar1VyVqUsaaxYt8dfPezf9cqX1pEaslDuXqVS0GFaG/9tH97JZ+LEdf5MVd3LqxR5oiS
G1rSUAC4UtPjjy16D3N1cOxgckqGd1l5dFb8q0EmTjJKSqDeCOcwL0A4qBP8iDeoUWQU9QaBO00u
54DA8Hl9h+b2Q6yvKh7CSOfHD36QqhBX9NjtN3L2avPskrpa0Awpkau27ZsshqYR4jYB8Ddqpr6f
R1GJgrrhgYcDhQwkN4jfwXzHfRw7pF0StNvtcjla4KiCGpeK4MWkv/fLH887Mu5jqYj6WMncd+qR
ptpg3XbcYxv/RrfnP61fvpp+QRrMg2GWuJxvUoJjgRmKgmya2SPTTgV7qt6Z3j2ybyYLEmFgK+Pb
e0Mmkfd20i7ofz3pzBz8SWCQgdmy7SCAYYk0t4JKB0TwxmEu4FkJ4T/zR8gwHe/XkV/vqt24Rb7d
nA77wJ4XpX0/tE0cSBLwzgV7OHQjw7yR3+AV5YO2uxeKd0PAVZUu93XhGbZqrru+Pj6d2+/1VKeU
L0JPZ+4XWFjVtlJuP6GYS1QSzPNOW5QUb6uY1wTdmEuDQ2iK4OdMlGyp3iBD9cSiG7ERQC9CFirm
vJKEJkuiwx5RDRNz4tOMPTJeKlvMzMD24oH2lpjOZKOoM4gwNcbcg+pkaq+aPvVUc3T5DpE2Y+EF
FtV3WgdASh5Dd+C1T5vAA5rwgEoTOJzF1deLIyRzACLNo/iWo2GM/2w5sUtzGim/erlVF/CG4eex
c2n0jdsCIBbAhwPhaMOk152ltbjz9F9UsmmhsTz5EeInxfQn8gLEV4SGu9+GDLCYV5926ucMLYpi
5poUTQFJ6+SP4fvsWWy+zahKG/1hyNTUQcvcZZcTF97+mCEzlnECe/xOdeL/4S/DGLYj6XsOPJVs
tRjN8HFKvL2ttYmjYdZIekdFoNqcKA+CcepmBmwGDOjkBu9oFuywIx70Isv0SzSdIAGEJxvRJ1pO
0K9k7vNs5AiykSVqoECeAjvjAGLaFT9CFnpjbx60RpjmyBGEZXxZ+/GKfOQLlLWv+xBPpyIAN5W9
Pmn0Drou+pdv8BHqwzY2nD11cZ30LewNagaxS8bDgbUc3Bp4Tg/Vfmv1A3RUz0hRQxmaEXPMHxHD
e1PCUfFUoAF0LOE19GPP/3epOv6wySvJtkOSzd4w5tGv+EjNeDPjdwAc+zJs3lEv5n6RzXc+l0gM
Th692dU1fFD5CKtHwXrMVUMTvr0tcjhowYtrDVlUqjxHVVrR/ktIou6M3SCKS9HxOzqJss1dYPxl
iAJ04j00aym7v96+he4eDJuJkVIOc2Jkqt4HHyMvWJLVVv4YWpD+RfaCF8soXdp9n1UcCsm7mbJF
R9ket+TNbZEAITIb0DGObALTzPLppOWk4IiJIKIURfzobmFJVm/40zQmWdBgg9n/bBvqZL6Qtdd2
jfuXpEUAmYgvyRwUV5ef1DqRRASN9fjnNVcoLmIcHbdGPnceIxuvfprsVmbJCEZc0NTkikOqLo/7
izSKCwqt6fpTqOVxvEN4U1S8fikmMMhyNk3UgVlx5kFHTvS+YnWSRPo/bC/RttokVLLdrmYprVEU
b4jW3uqzBQVQk43vw13VjDNhGlf4DQ7tp+ugnFiLJ+5TQIcuOa/Jw+dW6rNUM7g54hDVMRHJ4HYX
GopiZ0HedhX49ATpLFK8Wq/boIIHA1Vfa61s/eWVy0/ZUSn3IxcSV2RL0tm58zr2lAd+iclXyTp/
7KpEApNnRClRsjhTijz8yh/+KtT6d9jzgBdHaxZXM7sSzU5/DYh4L4OPM8rNDzP6y/XisKQtGsFW
pB0+21ImYwpcNFwzo6de0APa/JR9jsm/7XEwy2c7n/EbM/xIXWcGZUDDyGxL5n34J3Lqo3+d/Anq
pAKp7s+xCCZaSqx0OZ2u98+RmAQnHTjECbDJgfhlRo6ucFWBe28cuo3t7DJtE5pGW13osJfmBHU6
WTouf/r8xh7Y0IrePdoTcYSmIRUxugzBDUxAbgIfOzz4b615nhINc5t1tnUoYfaunJCXkmF7BypG
Vi/woE/7ZBNyRPSNovY/gn9gKPR8peHSUo/40C4s28a41d1nABzKhCNRQzXmcyVX8Qa+ZN2F6Pf9
pkvtqXiSEusGWLeDZg8rOUsEZAN+xfr3JBAtfPGiRKGwD6Cl9MeVg4LD2350wAg+3UZF4kzrU0Q+
6cbYocZALy9KpSL19CzHiCjpLx4+Qi36chVx0lIbMLCQ4xDyVkJj304vTu2t90EHLMEam4MzzZHA
prMPZs1OIE4iiDdZWgga0fmXW/GxW94PHmm7nldcsIrd6xkldC1R/xnL4SGmi+Cg+lLy1y79jxhk
oMlf9s5uEJ8M7Hoh6XKIGp1lMwNI9McjnQaGKeviJJg5u1AuDA6+WMwgVm/nZnA+eNaC2rtUGEtC
H2moip7leRWIZb46a/lrjq5NAXgNum5ei488gZHicNMtrxsgwx3FW2QLI16t9UJzoKtQlvqKAnj1
q/a0TB8xJ/7lNpHIU/V3UFs0q/W+3jsiC4Dh3rSWle7CewfYL6rJaCT8lB0UNBd3f9vnZwl/ISfv
/C4i2qkEqC1/9r40lshUcrKA1ONgxzcWeudsFk+eBRENfYnDIRi360nKEsIC8UaX4/2p4fDUi/Bi
tj4iXC3vDylxNSiGZRMbKLxqrtBXrN8kByJybTaSI8X0INf6heQk8Mjxef/8plZkKTeznz1yjp3k
0EkE4HDlB2ORQDzjORrjKvK/nMhucYQP992XaUW537aP//XGtOjlPK3DC+JNpneg0OfBkJ6/nPaa
QE/1JJpn08cOa/gKlW/7lK4C7Chs4XoRepmhQsrFGUsArQRXhdQ/OG9+o2HifPFAlMfy+P1+PPCz
zS+P9L2meCdLRIZaDfrW/ZaTUuotLVDtYhexB44ObSmOtoPLYDox2b/6MvvMjwfj26GJzG8cIPEC
YaHVhwYmn+iU1bEaZEaUsuyIaVy0EqHDfYlkvdqFdk0OzhaB9bK0aYCQhK2xw8vux0gzXgoa4W8X
jGXdxd5k8exMBtT704KS0s2AXSLYIBzbMir/ZCqSuv492kTuS8RykyBrDvCKeajrbwH19yj7QEul
VVKwgbmD3WL+24uq5chkqgUWPa+w3WElGwF1nosR9ClauYyQT1gv40kwMgr+YOQZDALJH0b8z5Th
la3LcBGITlKGX+GmPbzorD0OvHsOAEpckN1wIMmhhXEJp21jYrAl+zaJGTneGYtnSREILWBKBuR0
dlLNPp3560rCo0zVpt8ocickwbOqe7lhKLNjYAK+UBWHqKW2IBzFDI27FI2zle7/X5GsmmCZTpLT
JeN3l1ZWXI+ZWHdiuUl1KJdpo6zNhGS/hwnNk8tZCVdgl266cRQnEQvCwS9XOzPhCETt7PPiTkMU
Spq6AKPJmLA2kUfy+LTGibij2ppidR+uQVAuIWCRz0eWQ7ulqwrtkO1/G4vV0Hn/U1q+gPe/1NqG
0HQab57rFg35zEkzZPRD0Ayj6fEJjEqKW43GSMkcS1d8+4hyYtQbwwR6LaJJ8tucNStrZ683BKUX
Bb4L78RlIKytekc7ZalMijNiNrtp4RvP9BMeLw9ruiHe3WOrXsSOAojREjgiTToVtdd4DPauQQqo
OFo68hQTeKgT26RVzdRhAxOxzlYM4NzDiiRZENfybtPeFlbFp+qxeTr/FcoknUlRtZ5ShkF4aA/r
hlLSyT4XBninG9nFQg2WqzTMYI+kKb1Ll2iXc0ZN9OAn6c0x+I7L3hRY/vuAkYpb5dhSiQcgAp9U
G7lOslSJv9h+++EGSGZrkBKI1jft8Ueplr8U4UNLVtqZKyIjhEpto0tI+9PodoTw76P+DfozucXm
79Af9rxn3ZHMHTuZ2w2suvdYfOjF5cQWqeaI55ynv7UA9YsWpwlNbmiGEc3RAZbIQlSWbX2jAKP+
XxMD1/TWSrZPR3GZncrRpZOVgsmXfrX7IM+RE1fYE8nbnMFCPhRxL0t8wWuLOizdua5uo7BH6a2q
OJWCEw6spzmvmWqPZB2YLSnQvKfF8FFN5x7SRjL7PFoPL+QhiiCi2X2QC7j8n/YF6T4qdzSBTKKS
jMgvrEpBRepeu1QmPrIklguwLds6Xh4ts0aXP+g8ovh8cMpUzGhAnlS5Hled9NHt+RU3BQB+uc/v
tIFo0KjqWBuFs9ypkdQPcmlo/nQ7MZlXvTTbs7CXHKDqNQ0qt/lfMOqsWz7EKJtEWMN4RZV8YvD3
Yz1iPM9JgN8acKR9ShR+iT2g0MbvUtZT4W9V8B5BS3InmRlfahiymuK9okzw/ZyZSbTngNS+3j1U
Uo2ZGMwv8g2dx42UOBuK16hPFmFrr9GpViBNzhRONikhneRqu2yCX8dXwXyySu6FgKQBglFfH2SY
kARa0UBSxEJP7R/dwoobppiRBRorLxyNth/2aUD8a27YPRoCRggFPIz5OAIE7rMjtEJb62J0wTkS
dw8vW7kR/5P8BAvzPXi609chege0eJC4aYPCTRSeOmhqxZIBnUmKDaT1snjpiFrlIdu7GO4ROViC
j9xwbwbEi3qOS7T8GMZZMxpH1ZYwZxevjOdgwpsS7aDd1UEv+8kDKUJ1e0NxRII9YziG+rTJYOge
9BsDdS6D440GxWE4lx8bKBZjK6K+ZnxnRLDhfkC3Kn4jCfJWbKDDx6FWi2fjlRgy851gK46My75m
vWg7Jrla051Vvucx1aBMlKB0bLIxFYsd2+iUMtnP0w7SdhLdVMnx2/L6wKr62cUHrzDxlnKmAZC8
8L2X7XMdRRI3G1VZqRUKri6ly72HAu6ynHt22V0Y7yG9bL+QLKKvW/Li4xiCblOy8PforQu2CVAh
OTKKX2paTryFhqguAqSlxKXtmDEoV2LTqzZ3PEmrii7ZruXmdKrCOjQeqhJ9ie747jORnJI/TP5E
Jk3uRUlXF/AHLRGXJm+oWo9Vbrz4OMWEyHGnzGyBqh+6XY/3w/MhK/KEzG+vBWQ9dMbN9ISf+akb
respkp6jeY7mktUD3TkLIVK4sbl4wPlvX/fGRuxRJn6aEf8zU0/lRbKQHgbn1PYYccRjVyxWOfO5
TcZZmmB68ohM/7euzCexTWXm3xgiQLwgeDC9Zk7e1T0d63+xGp0VnNQhwXXiiYyLA6BGW4NO9uXy
ed+bhChwxEJO75HW7H0s0hx3OjnlAFUzXYn9mFtBvSJtxoEfb7AQTPGel0QfGodGdPAiv04V+f+/
rFe5cd7e/0tFONKetUDyKFo+yLJc4+QmRuDEkYSuMrYU1C7xrb220K4IwPi48PzzWDJU2cGMdVD3
a1/GzG5O+sFQKLIFyeYpTplCtWt4QHnlEWC3gaSBCrJzSWrLR+4kuwjWsbN+sV9ByE4Sp20qNKP+
8fxDCnDZDhbuktnUZmcetcxmg/jN60ktz8tinFveiTB/bfRSTw7+4S3c7+6d5DnQbUgNBzlSgYkn
SSq+PpZHZz5/umBVyUZKlPQ0440xYRdhDDISn9hstm21Vh9xsOjkPWObdErRYQJFrXgv4yzS7VzC
hBxhkIGebr9XOXa8TFo42m4ry9nhg8MbW4W+P7uYs02yIzJDz75HvlPUhjOLE67PH0eYh4gRrqH9
rEXtvw5/egpdncRFGmyhbfN1KUEOyBcZ2hxN9ad+DzfKJZFjFndmgMStBecyxe71MvK+ReEmnZwq
NPfVlzsAuafR5WJuS1fm+kkRrjRj96rrd5kK0Kfwb3mb4p94hxYY0KhaJpKsSalr4CpYBrs1/qVZ
hwA2tz9JS7HD1UvPLI4tT+rmL6hXoM1XRg3CnjzmBko7QZxYjdNiV8CZmkSA2t2qSOBIHDsY/nNN
fIDIrCoVYm6G9mUjOY8QL35GeqTlDrzEQA2yahAhTpKAOrJENrD+3l4xK3WZsX2KbbIjBgvtCrRW
2trFb9hkJZ/WT1M2Xi3BzncrMLZcVWUMieSz+0KKt4+74IDEbx+5TvX91KOpTsY+bkc0hwq99oOy
4nRH9vCGKAPKtOPto/rjYAoq69Y4Ut7nq+5N3KLL/zMEyt8J6FHdwboP4l2OyVhgCjwPYjqPx5Wc
PmN+0ZN2q0ux07sS7jHzK5xiMKepM9KHpwozWrQ4Vxq8u8JRPINDPQdQUBJxO9kGyqVPhSharzPv
r4rfTg+IkQPni4SZremPNaeCdF5fhqd/SLJQGp8KNWIak/PgpMCeJ/erQhkaehTvsIBTMEvTp1ll
3+LNm0W91LtFBi5s9zpSUsAML9yTyQ8Z1ulA7fVR6zicHG3YHUpNpZAF3B5RDDIvCPDuWOOgsopx
RpgJvx1TGoH4VP0TBQPDhX3VxKVu8k6TBkrBlWjJ0gL8AGcLN3DFr5fpLI4SgfiGUxCobrvYmVXi
2C7EOhaawelhW89aqCbQow/Ty9evKDygmdebUIskX7rq8aYXJr6G+CPcOm4605WP+Awygs6f0t6D
RYiXT/bvuqV+e+egk60N8vct5koRnZDiPjXuHCgOYqqD1CAGq+KocvbYbQY4680eZ1qOs291cN5Z
4jUF/+vl+BD1rp6zhH64K2OIjeqcH7DFjN/NgGmLh1PhZsgc09XXxh0RlV/x+UUtC30NlIh+hvdS
nCLpeKPXfqM8XVteo6vZKwP2TD6jRL+sHuw/8K5mg0PuwQKkt5tJpI7cFbgzoq0GER85a99ZaXpu
WH32QPEYn55HybA4+mFV91ZE+hbHhXtJIxUcOoC63H5u7s0maRDKfyCNIQy3fbjqu1qGRKztslm8
jTBjU78czdmjRVo3kH12NykTIW+2lZqmrtyGDpBwuFOTV5KNL7AbsfO/lEe0hhq8Ajv3tIpX7dJk
WC1LBr3mmZ/kCQ3fKYTTAnZh4cSzQHtaLdWWrx2ephS7zJEW61aSzNRtHkHvTdSWJBDum3cpgNeH
KKIFRIlYlYF8xRbN6uc/7AbRYzT9OXRrnLaB8+ZnR3hTjY75UzScG2L3DhYKQJdFzQkBH9h21WR3
0yaBUDgHOeKFQumZyuOnL5mZ/SrOgohX1WEtR0YBwsKrABTaugZyZC6toyAbDAsMYTt0WvoW+4O2
yXEPK+qPve1kcvZyOSjlzA22vx+AsCkhskV0VWylagPDhJ5O+/2wQltwtDT+XeySIW7d/n/ZgemT
wAb3rItkHC6qfZ4xKz0qXVVGmq1ckWXAh7rAkem80kuoMRhoBHXco7d4Fmpki+g7bU/4/7PTfZPB
hToPKpZXD870eCXVk9VKUC3KQvXYeGlphTu1Tt6X8moeaO9ld4XLF2PflzvBZP1xb2+ta25d4DJf
kIr5VPdYSkTJl746FNnKP/mJMdgOD3yfpxhmbl/CJ3iG+7iy/x/hl1AUKkpMgM0lf3SVFoCVZdeY
fdQViFS4r7FEHUAZvwOl0qdjj1MykDXtqFFRTKX1HwUhWbM0J51rQwOKEs1sMpaKp7NW8cSPRqMR
xSDlkYCRt6Kk5ndHeL75C0+E1akk4Nskk5QTmjT0y1oIRZb8Jc1Xu6itktbmft61Bgq9n1YVxQyx
Z8xMW8LnCJTqvhOGhOhpOc1g5dTT5lzYIQ3lxiXcygo1Afj0Dwei0kAx3Dw1Tt/+LrfGWYdnG1tK
GWWLHAu0hBqncdc3ycCGg2BibQnoo6dpQvjMegKNEf8VRihmo9g5s5dH661wRzPnqFf4RXajD8Lg
yUHib++3tsPs2y19mkPDI3fB5HKZhqzAT5R5R7+fUXGx3F2HufykvjJRsDi5E4pXRar3ygy4u4dK
tXKJYiG2+LWPMVYlfe3nKLhrD/v2exAx5lmrl9eqFQd7Lf4jrJCGwBhR5zLdqgtZAMJCK49oHpnO
KzY+tcJWNpHB23iAUoRPxYfBRS4+6xKCIkMYB1oZ8aCpINJvqMPh4YVQ45usITbw8WfsO4QPf0TP
la/Dutthoa5v72D0P492TwRdMJukOUgXhz653cFIK5OXPzOR5AOTKfgw/FKNu7oZKvSjHsZ3kygv
8oC4n728ZE9c3oCXlz5c7hYtPDwMRdVM+pWLEXksnmyMlh1LhVbdyQ2kyQzequtGAwBEyB1+as9U
LiL1BeGxB2eVJrwoiZR3UEFLosFNhEN6LHKQQKkw/pkAbQvUHJR6UmAy+ioxrxMwfLJgp+c299nB
x5gwtDZqI8iUSCzsT25rNW/Tywg9nnxLlMDkxEviUlulZfyZN+cv1rlSSf3zyhQn0MhtIlXRwXtp
hAb0X1wDlyzmCuYG4Y60fo1GELsxAGWgKMNI5Dz7tbrpKGmRkI7vQCkAyvylBLLpGS2woB56M/6q
h1pfM6dQox+UfigWVWyYp5Tw+kpQ+qezBZFoy6UWYxh7FdxJb1kbTO8AlAup5phLDExQcfB9vq1o
7dRCt4pVdb/tSvjDna1q2pxUTSWRvmMA8lWXYZNDCNKQaBOpTxl0vsz3upVJ196kDyrYwni2sj2A
ZLVCfFMhWnj8xvlnVzxz4c5/QsuaoU4FRdP7UtY6vAjvcvfoJD4/Q+YYrmP9BVTmFSTIheS4G0IO
NUULZ79qATDEF0W7/kpMze2V2O83Gnr5NQ4j7VGtKznQppnUR0ZsO4FLin3+Axx+tS9miNE7C8ff
vE5aacRIhOYbT66smhoOgdaoUm6XBbcH2LuAfla7ouljUhqNgZfgUm6ucoLEwM9Nf4DV1MmPpS3F
kVIdMxKISVGkY5OQsH1i9OSAQpwG50Ly6SQ7zhgx4FVws0Db10q9a9WukMiTkUltXaZRUBIubrNK
F/SPmCWkBTByg8D8CIYdaYFwZnMFSP0fNpSY2lU6pUzOpoS57H5EO8LZjS7baCwoZXa5rLy5L91w
je/wKpG5VcfsuFrUtcVUx6RW3ovayTvWvRaAI7fzbMoGvKmA4TExs+bZrbnjhLzketFVamev6/2Y
TUfu7QLaVr314UOXNmyfTFUSA07afeD6dd7MFMjjVDfT7TH2QGBnAneP+tgSgHurk9j5ti/zx9av
4/tbGRGWV8CJd92ihZ2nV+bKtitNTPpSTi1us1m2wgYi4RFmPyhijNVLVy1TRO+7Ggn3SyNg8vM/
tqEussbL6omB0jiuZiFn7B8UCdXnJhsLNMvwJDqThU95SLLaSu49tToty/m7VumMyIMK3ZU+U27p
X1cuoUGV8pR+Hlf+BjUml+IHmCyaArRA2CCSmnv70sMJubGeYrl0e1fY3jc4zJISy6zrzwqPWQRR
TJFFbp6NrGlvhV+t+jVpM0BEmzmQviyDEMw/Vc6KtC/75t9RwTmoMEgMjp+7dir62lzorwPdArTN
wPNxqoDNypk4KUd++dWkHwySprsu8NyXAl7ubvgw7NTgJ3zDOk9QvWJbrD3ZD6BQ5JW6i+kZqHuL
KWKKhUQf8Z+GvSlb8qa6ce35MmrU9V8qxj90yrsdzFUmrQrCJUUm2AaCAw+8jINvh+1MY8rf1J1y
ROp28erYKOADhljWF94lX/pxI1v7mK3KjO+M3/72KYy13C/5GaKbJ/FsTEJYo+qJ7C68bm68z1EY
j4/DgKqcu2DbhZi1EJMnW6T3lDy9bfGI9yRa/IyEC7sUgBjJX+hLyGh+mnV56p8bZg+ZZ935AeyW
SSDzHBP4HF3hUcRrk3LIbvfywHKjWP9k40ndvP4u56At2s42M1D2UltQvRXr4PxTyHIJ9DwtQplY
orsv65EwkPjsNYM1x0SsQ+W1nFuTriE4ToF3ly+zLNmL8XaASfHQqq3kCwTw0YpBWed6IHiGGn4G
shY5ekcU+YfnuERn2PdriVfeG9TmIxl116Luewd7+epVGswqhXrXt/RkV7cWL8nFPPQPdwKZh+YX
3T3f43vmTSzTMWCQLWNmdOGiW76YWxgKwFUlc0uDW4NiQ6havt7dSMwy+nVuHr9WD0D+zCR+ctoN
+u/1vZGms1qJ5Z+Gv8xu3oIPes3m5Jc3qm1kneYVj7jqH18pZj2qHui3g3r1twfORaRkjyGjjIU/
XXcH3fZvjAWFNHRfvbYvENJ2Kr2FAbCnU/fMP/i5GR2LAir7IgIF4GDEPLL7NsJbAjEgCoodFIRy
CMMBbpjlB87OETrMzACq7HOmfFjS/1/MNRQvZVDgdTLej7Y/xxI4uGDHvh5lrF2O/IDKKEzzdzEF
XN134BZjy8mXYXE5LUVfbFKqqqWLWvBzsNDsJB2wOluA0glt3LJEvx1VnVqQl/nJVbblVh0NUpPx
Qq/wLpnpYPO3rpqqTZu265IGcI80xsPxcZHrgAt0x+Z73eqGsErhrt4UEgP+Ay9FLWsxCelvHhgC
gahFy3upihCQEnYuX3UMquCI/NvIid7fqQQIuBTRc5FzoEaExkVSS8Abw6wSxpMRlCmtoA3b+cu2
F6n+UPjquJlBzVFHYaP06Wsz8h/+vuGVoovGwI60xbxHf3gS5/a4GxXvXE8+VgZC8BGwRxdZMDlJ
ldThJXNvW3GnXD5yttXsbcphAwWDvfhXXv99lH22UFOC7Lc+rVdsZwH1do2s72yjPAzL45vNlCdx
t+wciZLaFhNuCk0qV4+VkF4z5Dly0pGCa09rHMlcwncLLi837n4WiTPQ/hEkcVzFTfNIo9KFH4Ih
rLkrby7nXsSe103HvGslZlDocaOmY7qi68EQNvSWpp5UY7vhH12u6cLKXgQ540IbhZ/zZ6NYQ6PQ
ZwsN4SPjQ+8vJ7CZdPTpuJl30F0CKgqUuI80/1FbYeZKwd3Tq+lcqJxmFnoedCKdav4hiohIfM/s
GRXMdgB84idpvMECsI0HwRguqrQqMlZTWYOaQ7sJdUozH9y16BqXvQIyXoH2y9apaaILjpb2A3vo
pRIDpjdgjueBUaTzATsTFesMfB79B2TxavFyJozHFJJB8xNUYnfayuQilQwFTVqa0nbN6L4ULlMG
WzVegb1Bmf8xgPTxZCC9FEpWlgi/R+S7NnKSlgyusjTJ0fW+w32SNpkPzWHxo0Z5ifk1E+JOKA4G
Cxps18SOMxAWnXmlgMchbC4zhPQKl3pRIjLDnpdV19hWl7aq9unX4zV1hynew7rIuZ7bszknyJu6
ZKce7nzQpfG9+pvmXIlsEx8B9/cjxXx77pqik6u2oRgjApw2MWE8B7LhV//fsdUysNhDes54evZc
em44a/SG+mcETDNZ5+hLXnmX5Jbz0F58qYPqSq8ryAV5w3RLWnFERWcShexWukzg7rJa/hbiewv9
2ElD/7qrSdHsPUT2PYR46QEwLA25BrH8ihoRp/UfsLydWvB75ywdQ3TDPCMoEkV10I/Ptz+4Ut0/
u+v8raiqbSBXI9yvbc3FTUKATjjzwzpxxjZvL+SQ5FW6vtNyRNqcCLo+mSDv5j6Al+V3XczFYt3Y
ELTxn5Q5uVzODBm9yFVGLpBgGVRtV22OwK0j3yF+hvL0VQiI4VKCMOylPb/tNLqiD+J/yM0F3TaM
xyD0Qt3WBjvxPO4D/2kAPzhVE1WdywOF80sHffaTt6PTlyU/nP+t4qDyXZmSKNzqk5sZjyXt6LCS
Y5g8P3wHoU6tl+aRUcUZ4LOiKYbgJjZ1BovllOn5LOP8q7e0aOwer3zvZJ4pT5Hi26UHDF4uPmPi
+VNT10cAz4jz/fgFo39PTiAOfm5qgENfoIcV9Q60RKrxSw2vGsREozRjk9s906RmLMWc91C0RI6Y
r0d77B5k17bSbDreLwnUVCSrgG+9Xvf/iaVTdgOOK6ES0Mi5ed0We+/c9O2np7sef80198pvKV+D
ReLRnWzXFQ6DJg/9RVrUpIOaVvgPfvDLi3stCIxyTvU6iDeNsYk0yp/IrNFP/csz8PaYI/GGzkia
JgAgoss5D2CBOK0Z4z8yKxBhtOaKRJXSJn1pJCijZp4zOtmFw4ovED/qkCMxNVsnTKeRgs3PTSjC
Xk+3Jk70Z9uvVVuuv8kpyGG/uA1yaNgkrEKE6dQE6CNWShJMepuYupSAhL1cnMr8yI9PULPgszTO
SiLC7+EwE79nVGYmOPJyYggrpGLwOXQB8oxBE6pchrN1U/4nilPQKlAZcn9Uv/tOfIb2UyvZpI8h
zhYy36aQmtX4Fg7rLkjzDDhHn1RHW6V5GPfct5aapNX2bYJezq3f99G8Ux0HUEXpye1/OqFC7QRV
9cUT2cjaU3t2Pz0ZZyfOY8EEZ7ORREFc/t7sl2K8TTi98G0WJa/kgNqdDrqcW/MUNT3DTmd6gl5p
G6esk5JcJpa3HNBLEhbqHARjqN+G6vdHszz8bWcrX6MvqrHdgbCsWrLXiyfiBjTaEOpezzTyrNKx
cOVqE/9KZlJ4nSLJPz93oH7KrKn3M2E3TqYnJFwTsLqJPfEJsaP2PivPujQpiLTPWYIdr/nWvHfb
l3CXKf2JobMu7OdyJg2h9LlLq5DXxHjAtr9W0tIyOAHlK70LsxxYCn234Xu9Xah24zJb87hj/nme
NK6BoWqaNvk0E0FxnNfwY29eqtYytMxFdU6XKOT70ynv2ynk7lWA18jn/XVPoGvN9EY4PC54mVRb
kGP6/+pVGDWn+NUCIxJryv1g75QsjQa/juS3lHU91HgoNQn41b6/FhD6PQJrkRD0EGP17SUcj1a2
HiNDWYW41fT/F2WSdsMB7ZHauf8Itxh++g07nXpQWbzuCXuuS6sG1GW13Tkc+bJylfVlUJ+KdRMm
CUa2Yg/LccS8v3cK4oFLbV8FZ6iPY2ixcBsWQ6Igvm4mQYhp5rNB+woR4iqYOjswU7GwhokhWP8O
6u4Qv4MnduFppdjM4GRtQsN2g7CnubFmHa2xrtCqib/GnaoBJCnazcISGMTuOy3d8q87O8/fWEJJ
uekdAZW6a2GOw45mXuY3lTt0LP+xlWXsbM12nFlTIzqtVQ0gQBuato+REY2HukU36UkVT/K2hg8g
eVWnTX7c6D33aJrtVMfHqTYWpzVJlfNtVBB415ilPNYb81qzApNI/suoyLbihCHD6GxzNNABX/VN
RFHZIoz5NVQ13MpHYTeNw0J/hgHMATkKIyxs/UXBtSR7wRr0t4TxlBf22vsKQyagfjNTwo/4FO0B
0PgBK3asBhtXvWNrO6Ywb/nxmUsMgG0gUO/SN0IMvVuJ1l+wlgeapJZDlAgglPUPF5MX4OnR7qio
VkKmdO12TzrihLkCILrNa9jbq4NtSVmZDsOMAhOfK7jZN5VwPwP+8vf/RSsgU1/XfLBBrqUEfD5b
dkDiqK95ycS6vYeh0DQalpqPWFI6t2XdMidz4fYf3cfryN5nw4o+ILW8It457ubV2dUMXeM3fKuZ
1lPgzthDhQyl8/Qus0tbvEBo0aaW0b41/WW4i63hGA2CoIFb3Qc2yr1ltpZbW0gE0IjTMfv1UWq3
BaXZ8VdNNMScuQLYBLOk+Jk32bUnYug0m3g6tjj23rbMGQDRA8ItRvvkhXHdJhzbvis1BhrFHICd
pA21R4jxjEYIoeB6tJGfnkGfU6o7hPn5LxVIqNwoMvs4fb5yoPBa3paVIoG5TxXBKhJllUSkV9tz
gcoDDKrl7nF1jNdGAYbL090N6GJd7BRS4z8pY2WxKIcd6yLFCLrHmB9ol22YwVo1YO+7skuY1rkl
3iWWP4S3/cWF3/SKIndZDQ4tHqLukV7anbdc1Ntx33nNyucDtddiJcZB2lCUTLMHqLg/jdq4zEvR
BqJatsbujAPK1rmLOs0nfvAgD35XgbAL6YLN9YigX28QED4qn27cPh6tvXlwvNBHI4UiOAM4HjDA
dxjbDSJafG3mc2TptGBqNdBTpXBrsV+jkDvg3HeEgDibZ6uUNtLbWCfeH4YoY2nXFQ8+/iNNaumS
QsO/ORRFz6xDOsB+mHnAJj/g9e/p3sro+84wf3C/9E1zSv3Jd6AhmdExUXlZ85mdipfB6QW9S9F1
e/YMZxJ4bdzn/pu7GuuqGXx3H41tEKNOXvUbVr3bxLKLZxp4lJG10PaJa0jf8dEJHGR2ZSMpZ2h/
+lfE9Q4wNVQNUygCyyXRDSnYFDfm1xk/uy5JlZvfW6Xi4uattnUWngfL2p+JCZtrPWQGdV69ZKHv
JkYfyyl5QxuJfm6FhaR6/WqHsvWkpihZSHry936GnfR1AWkj05g1JRBdQz+xsqIjp22bdvjAtuA8
h8YdCjqbyIzpzvvYGwWaBpY9g3qIMVboEOx4QPwBlWjLmwwwQsEBJ6tO2qpeTNnkOlaYdA+f6141
oTDAkN2p/uRNlvHhLQaDaPddPbtOLuPk0zhj0Ejc+LUX6pvJMMQDyuMxcBFpbpOAASgeFdhJBIAh
9l+86CWdIpK/SbKuyo/8KXYH8TfFGBFO/CIIl9R2+P310G52SAkCQTJNoeBSyOeFcpd3/3oyq9RQ
RTv5bVOEjsFJ/ZzhPbajXzu2jvmxS0YUolGTIq/PlAiq4mFiYrFFfI+4H4gHmN663raz0f397a+s
YbJaGGJUI6ft+Q4CvkF0RFNVc3ZGMscTstRVmp7plV2A9mjlHYX+DjdwVvxP68tDE3s1o+7TsWdI
kx6zblBmgWAfuP61euK0fcHk5IEUrZCXtzxuuiC9UOJ8RGbllHu8+KtpJJ/FqHEGb9uTrSv3TDTw
/ERggnP274Yv8qeeq6MUBG9aRuweqBSrxuQrhvmQpsNh9Yz6BeZ67Ncw3SFTo7Be0B7m4Dui+ZAs
Djjgn/1jfm+qTmwN8WQt6ZrNDd9H2QTVZ2dzrMk2zXWJITp7j42uAF9pn0jRE4PsNfri3HUdhHgB
0j8Nip6SwOFwelhaAtEgfosfLL0Tik/+2vnYrL8DP7XmdlAA3lWv+8qJDVXsR0hJstDXku6htTb3
5j1XSDyBUyEHCgLiskkFTFnhy0/LzN9FzFIH5KJiejGcQ/PA2KTGtPPcaA5dXi4fXqz3+G7/s5nK
Vt9WXoTFcknqTxG0oSbsQc77Xq86eTKS00CBw3Ip+jzTJs/Tl7LoUvFgxHJLD+GQBXpUvczuXo1i
UGAEAkVjv8H4xtebX59jOsAN2wFv0TNKhukJS3d18u8DfGs1MzXCYgVlYq3JXcfERZzF5M3nIQ2h
4GflgRWRJZIzwtZCFJ4+wYg4gwX6IyfrMHJ//+tXFA+nUmsfDkGodEicefUuFGP9wL9D6rNYHehS
J8lLp1ZhE5COLodpTcywulWp8Q9o8+80vJUdAVb+7q/Z/09Fff1w7i7+HHKkwb7XG2DU5RXScG9/
c/dAd22uiaTfTm7qg5lBldVS2j4L68nzt4ctJq4f5ZTIuoGrhezL0UJfMc6Omcu18G1HwMeDB+Zg
HHjiO7vbGKa09t2v5UjtT54RC6e0cZEKmRGkeQJri2pjMTqA8w636XOcxTFRmcLWw/XhHTjrn8Jr
W2t/F2pmyp5g6LMb26rI1KAnV9PtuzW8KK5LytO/3CKiO9hhr0VvMWzVSNGugeEdkAHvd5pkxuJ+
7NpewrVmU6mr9Zl+1S8TYk6ikrwvLAwig4l4wTzvgyPlIcveTGHV8ZKh4Wvt1PH8B7s0yI8r31Cg
YZCP2bJBLIgl8w+sn/Iu4ieOuHLfe0aTjtRv2QhsvDBiMuAh50rBabGl75y3UdNatRXvjYFivdQR
hcOv1QTh4UimxV2ELiROxzmRVDomowqj6dFOPekCs44YivjfqMKmjqIzY3BasskCEtF1E3qrwG+E
b/krC5PFsrN1tmm0rCaycloXZXa/2kK4mQA0GZ57ZruLYPoF3tZ3cssGyM8oDLGPfklhtASC8YIc
znO8N36QO3KYZ8hXj/NW6pimoSlqZf/N2dT3eNht8ERnIUUnZs3G9qXIiOZgFueMeX9Vv155S7Iy
jxONZK0cmo02bYXpzuTRdFexmln4Wo0659mT7dbtOmuqR25qpxVM8CloFROQjBDWg/1xdP8GM+Q6
CIb8oytvh5hmNMnySvLC/EZYkS0G9Arb/kJKBFHLb6FakKnzPMpEb6dcTz3Vhq+JbzZ6Hl8I686s
PdZfzYGWpJjetqjHgizTE7flb9hbvB7L47c974Gfisxy0JSAKAFAYTaXx0A6r/Q4aOInXZX8iViI
vZj3L4MFL9PChyXglcPBtFpxdDLe5NEjS/Wrzg6dlDyW9A8ufrDiIhgGj0jERJUpcyYAAkuEehHd
tJYtvV8dshzijelSd46HB/7apGk8Ck+cZn06EkQoB+WAUDZoVM/sTZmfUMIO38SC9wlZ5wGgz0Yc
mhZDg+beJud/Lvg2B436QdIbFA5dRFIbF1hrVo2OIXAIwfs1xSEkPikdmz98LOwV7SFMKwlD/IdL
NlFGh7BiOeuxoxvenXTzRUSIOcVmE2UsHttvs1FDBGMscTR/U+QsdH2BXGfJ6sUyTOGz+gR2HPOI
QKNcvaLOOISIhJ/Cyd3jVJcgqtOldpOvH9mr6dbj4db6LdjUjWserQg1kEIX/rS5uR/fkdcsteg7
LtlNr8IIvP+bkgajR5DxgfM7yHI2G5aDjs6qvvfjp+9baaU04ZNnEgM/PCNKZCL1WzPZ1H+77sNU
razk8SoRJ5b4HVgVTJPXJ1xtpkmLgPy0aU8PA4NJ0LuSAiDKotkdKVpVLVEPysQWz8G7AQ99kKs9
JXpdKM4hoNIRaoiMg9BJfy2GlyFvoDsFJBbFBLzJVA2HpGIv7R+mGz3sbhqpA6kGAEoMqI5Pe8r1
kvWAvE12bAD6vnLNsVy744uE+NEqteYJfInpYVPLx31W8ktXbV0gD5fpaDisaY510d4aLO8L5K39
h9QojZ8A2W52WVrNTzV9AkLRKNfoIYeuYpBMpeGqrGMZpaQ+UYzr81szwMx2939J8fVXC1AkXuJ/
KpMiBNO28huiOKld48/Pt/U8k2H2I9jt6sTIohAyoVhhdY8zyeH8uiUqfEkVgmsoOzjKRxZFOT2f
Nm05q079J53j/KanciiWHEQKBeIpwoTfmXayFeaU+Oh8fJ7cQi4IPW1m4nEo7dOeEe0b21+UDMaf
3r/Ljusdq6QTm63khV004/yS8BBFsXkg3KwpOtgaxlKZPxz9/uVyC4BgYgkiIOcH/dF9l/xJKlX2
4J5OR2a0zHPngpvcC8hzUBUsQvM8/SmARec/RnDKZY8g2sGZS+EBbyG9KM28pt03WFYQKKbHdBbv
7dXJNFCjLs9y/T1N/vIwAGzbLUhsOQXqVhAlXgKMifNty+9Yi8EOv9qrrdi7UMbh+sn0YnzNhP4i
wJIURFQO/jh9QAiDlG67NL3zpzgsKW4bV28Rhq8El0YisvS/BDij/52/bt8n0myPoaEMqraKx2ZE
IH3UCyfKFHO6M0EcJJRllxB7nufJVIbkTK1tkXffLOvdQc9rEYfGBFmfTqDZLCNJ1y6onK/CyJH3
DFHmsbPyq4/q86hFmrwlGnKlDQSF8MBl83eov1CbtivZgP6ulJYT3Vq6WT4FrJQrIk2YRbXozj0B
S5p1GdLhnWy9Zm1I1MbhAVVfHQeKMUdG1o16x1nhf+PQjxWJycZIm57RWB5+4ulsdCcBnO1dhazp
DKr9U0bb4q8Bwl+JFobnaolEjiQnomAlid1/XIuRa6mdlStFUwUN5XMpv+b6uWFmbwhLJbViLBKf
5Mk6lyMZng86r4GcdlfYN6sCZa239898eapt/Gc6MxDcJul+6OYUgGB1plkuWnuuRDuLnMdgOdUh
XSmdSm8tQDizu48xZVAyJTiCdFSxb//dP/0MKseUO9FzvT6ImLBxYDmxHfa9M2XbGDHkJcgyTnpp
1ungePBVqi4qTlQer4Wp6vL4Uv2zPSl2XvOZsZ5n0Ri5xBqd4X3VqoUW8lVIVNF80vdXpWl/RmYO
1toBWvRrUkL/kTloE3VbRJuKVKCuw8uWiJiF6TblBUVFlsx/YkYN4Dej5waeQmLfLH4nV8hv4BsU
5x7RMJXyrT1fdMKdNeDuecWA/yt/yEQwfE/6TjPObEw+kGbDiTEta5IiB//CDQFkmYzr/vMGKon7
AN6DFPUnUFDyLqy5uIv3Jl4zf+ovGAo4B0GczixbxkrQ8ey9lSnF2lyHoD0v/tv66bidpF3ln4oZ
UY3U7C506qZ8jcYVMd6iQQZUZu3vaHxfPz9Di1yoKGiTKthW7C84yfIEg53dsMSWav4BQT+jbOgO
Da2FttF5Dpc+KEa8USk7gkszgZVsxaeAQ+rG94/2Aktl3v89g9Z05/gycBp8DNec0PCgsuwUBMzb
kb57C5o1S29Hs7y4cFPp+CogSyW/2uCmVLUN818r+h/F1ZyWVuL1f3/AALjC2Lpnz0F4MGE7rgji
kH0VfjN8OgUzOwG8QGRrbWTifqIP6v9+riRwbK9eWA+JVVJm9+1QihEh2naBRbuypVYBpwQ9tDM6
4ZnDQwAGqEBdar6DIe7Tz5hMGGXMFE+eLtNlMPHf6jq9c3b0oevzpVpT416en9gJ0QXxXYXsP2z/
ZU6Ns3dPRm1qkGOzY7Bn3z7ccoJQ0JAXJ8e4mw7rZUQq7mUGCZ1bortl1ujzH6/rd6YZlXsXh0kj
dxQWWC/IFSc7SEUE/+7REzmCoUlhtPy1SOXwK2W10bmK3uvbZ2XyRckkGwqnOcIufHJljid4VlEq
jXCJMG5/mZAyeW7AVVIp9Xtj2KwKBADy8KQtXjYbj6+4cfjzv9KXefSstznukE7bDUhedNlrG0BC
FHB8HmLcfc0Nh6+bbI1USg/hV0e4xWknx3CCUSwak60xPaPwN5cw8mKMWeF964GG9GpOxqcrHje+
mhMZArg646l3TnWAf4CygI9QFGq9s7rUhFpg6q9yREBmWQr8LOqDsf2mSkr4XsDRd3fNyBTrgbyg
BsjCSPlziIPjWKBdatCpddw6tqU8w/uQoGzZHvCBsx4YQnMAUizO3x8/Yf0WEo/IU/ZlFOkWo+Qf
aejbIeBImLMowYAlp3DICGSmhsfghQ3b5IIv4wf26palxjHRCfkv/fWtP7T6cul7VP70/q26zNuk
GX6OQAQt8thXTm35mikjLH0u5CYrSSBhEcvbiv2dBWX/gL0nrM3Kc+uDwjnqRqadvid3J/uYnzWy
S+Y4zbi9UWqEyTGbcoiqqB0a0J5WW1uZx0FhEO+0jTaT2Z8k+glrJXHehI6U4n/zYrv2IY5mfCsk
OvscLWchUUHHDGCeY94HMlXPdtHMxdndE9ibn9VkGAOATdGrFOpPf7RXyYWe+vycAqyUjatonMqg
4NrdUZjOMGxmwDV4+WcLuG76GNhg/yvSrS10zBI21YPB2pcycjbJwwuRSBUHmAwQGLUpSST4g0Aa
ZlUapzqA0RNS3clE0o9Y60zvsU5+kg7nAzXp8M8WJLC9qhzfnl22Aznt1B/vHSSCZYmx+CcIiIp5
yBHM8IgFZzNikU2vdwnjPz7NSmWV83KY5nizKLEPv3WfazL+PbKq0Wx6n/nYVuEW5P5spts8Qx5e
O5yvDMtQrhAhjOA/2rvesytfKO6xqa8rabAg4Nbmkmo+0YHVI4ZFsXhO8kXgGG5ADBWC+jlOOo8J
nei/atlVI+9iHrWGYnZRAPQ5ouJ2/plKmyzJLjeKqiXKevwlA3ZdVR/2/Rqv70Isv/Hgu7EM/Z69
/be8J6azIu9TaJRWz425lF7sCuDr0QqRRqntfpnPsHclRDsCBNV/ZXn+15I8CppugNxrxcLSTMaq
B5wWs4/5KYTIwtTMngPV2UICRGxWmX9ZXpU9pQRuzs39BrDbr3NkHGw7FTEAWsaSh8Ewavt2rVsU
t4MYrWAcYZSYJIXXiyneysmTCVhT2Jx1BkFYPjVD6Rb4K/oV01oEHoNrAQBvWAgAR7IaiSk/WqFZ
zDA/p0CFwCIpAjQvR/pzZBCONBgVL9/Bm2uy0gzNWR+gjHVDwmMgN+UyKuwJptHFChcloTN9Dzv/
sIa4dUF5QhbbB1akoaL6WPWDuWwYA3ZKWMyXRnCf6wqVPZOlvDJtzLSKWINr8HE8yQ1HP1IWl/QF
3sksZ4ACSVNemRK6eQ844fc0Rvpuf1QN9+WJPLE4s4Ek6yP2PobUEZHSAWYV1KQzJHWbZJldofHD
UVmoGxu7IZ8XD+1ZGAnr3tSq0k8EIlz1eQRuykuOsmDXUYThbzodg7/ao2sre93ihufVVs/pcSyl
El9eFk6sls/6oBcsGONSqpXuazDTwJPRcaN9ekZmm0yKtb81wyd5YN+uMqiDdVt+8EhnUU4Rbz46
UD7Lffdey/boQiCsYLki1Y4sN/+iz7Xewa86usccaYbGSZvPtQOOmJYJh2TwQI3Y3+Yhm1geezfO
28GhGVg7dD5Mr1xlbkRz4RrioxbbxjOfxwLEAGMUt+buK/gyo/YzqBvbIZW/7OiPpkQP8bWZjJsg
XyYjn2by4FErGpjvdMe+HOLccVLIuP2++aBXcY4TEXkMRx91vEaMeYnc/7Q7/TRwG2YojZ7U+53M
YyyO9sQg6zPJEASNhr4cs7HLS9lQ9DwkrQDnVaaXhQRfzGYZI3JA+PpbwvF2EfuMtetBA8TRnUgF
YZrqO+0bBDfHkhFrmdfg7Er/ueHw5AwMZ6OHUHFo2CJPjBxKeO9HBWY4ri5932W6bHRvNsFUYRHK
D0F8vn8XCcs9/Y0gZ5dAafxr6eSJ19OkHFasMxbC8zecL1FhkH9irvadGl1tQi85TYCfi8/uqwnX
nOPQ4JNtcijrGZPoKmGf6Awik6p6tKwrQiCH97nYCHFBJrN9EJOgWKqTHvnNJ4YRonNH7h4Rnrfh
sP3zmo5LHeijaIrxE7niP3lsXT2La8K8Xqv2mVxjIqLxa7HW2PCTvtsIoqCs9QBDtk7X7AAUnWOJ
7spL80eKUjAkVqh+SONIKctcCjF1pNTgyNXeMBOyokd5vMZQsXvEb2h/6SwjPzYdfNuDu6hnEqCC
MOzQL8aMEWgRLXohnhKHw8siA2JdgnX6WlpGuMvP1cszL+HUsdD2f+HXYa5riv0GK5HkNMwNcHf3
8PjteuvnDqC5zefBFZ/gfyZXx6iyIg3af/aFJrar9yVCu61ZoPBIc6tHIWiMcvJun0fNE2rqpmc0
qoBBmQMtzJoVbHuSiuN4wpGq940iCtt1QVleUMNNnN+HCBlIcD63oNAhAuYfUmqB70KpfMJwvfKZ
Gva/BuforSt2z8PlyDkdoIREWQjcTq+I7qAYZdOuToao1OizNM6iIYFqC0Ce0i14lD/s82t/ij/h
hSlfUo6WOLbLsv7y+BD9332wIuZWRg/zKblU1MhizlYENBpg5mfs3/Y7YnsxL6NKHk79BNvD6LzV
gtUzuRjXf0scbMoxIa/Qkpl46Pxv4d/5TplQVZuzevE1KD14/Z26VRaoMRqRkE0pCu0+pivdT5mC
KgklRDuQ7LUy87B9G2sJ6VbtN7UKcWffF69u8S7tD9e1ZGprkXujroWfXdtpCIugwO3EtqdSYdPJ
jqJ0iQz3wtiAwWyBhq3a3PZfyfOzsdN+3fWcMd6ySVSH+JuekMREx+u42mgUpF/uzduWD32HYYps
aESyg7dxOUd5yxFhCMaFW3xq1pe/UlLShfthhSgcewQ5KeSFZ3OHMrqcmja+DunesJpZwNFfrJxE
qeMUQ/B3ekAxmuRBHiXJg4oZ6KF2cmQZu/rlpC7Gr8K9a/nlUn3qShl+LKG+XNMY8CN2kTzMPY5H
2BSV7l6t4WTinSlDd0ZQODj4w36ZCXTLjHFUlzWSeoorwGeilq2bxkui6QrnD6dI/ptutqdUOEr0
imbWy8YfFYT49CfvrBDG6NtqZhOoXC/5Zmk9WAX4OdQKQZecsvdKjHHeOupLHIyvkSfZtEygDxH3
aI7CKY79p8mgaSvOJ97NtuSjrILi7KHv/qKbVV0R5orVhq3pF4HcGIilGs7sqclbC9pRZaOZpAC2
Sg15YgTHCQ2nH4q7dSNAwFzHmQx8lFNlNvuzpOFW/qTW0maartp81dVmxpYWBkHvUCZ7td+HKzAG
15l/gv4qQjrRg+cXvFqvMbTSCugHstA6uTzthOtleRb1GsX0UPNHBSLuD+mE3ZeQzMxiq01XzBJO
D4Sk7pRxoG3TEBS23MC4dggW1DJVm7pL9ARTZNTJRcjyRtFzSgQZtA4vMIAxUUHtIw1t1xSfptRk
fuhdUx5sN+J6mG0LMHT27k2hhoicB0uhgiFi36Mr0GQWay0rNEdPGSTmE68d+TWtj45/uIxekbPx
hh4TxK6Ajp/u3II9WbF85de3fSzlyAYOc6Fc87fLpnK/BSz2/cZbPs0fDJ6Fuw3Ku5YHSKZi9D1R
AuVoXUEJHrw7AwwwREOY964i2oAt7IXYSd3WTPIg+NOFjO/RHlVQZk3d54dN4c+yh5IOq6/wZ1P2
9eUIJ+DFDvwzYK+09CYvUOT4jP/SCtY+OOIKo/A6RQZcxea64WT6uzRIYHmI6xPP6RxS8473qJqo
7MBtkNMq/B6yLbPEDPmVuQNxEryc7/Kxi+njrBApnbONLXv/addO9onk8DdeDcxIi+deqO/Ttizj
15BvLTIEhAe4Mw4Upxh/acZtM5j79SF//5AdG/wjgGeHYnvdBQrsT/j8nT8ToOdU1wmraoYCTAXv
nkQ2gloOnfdItmAl/PeptmofW7PUjjt9E8XxZQL6yurg5mOLWnaR5l0PyD04uK6SPpEZVsgUcL3m
bA729bnOYNv0AAjt675qdVXj5i00TYU0Qjr7ys4Zbto8qNzdJ+LIORHO+vfFE4kpz1+b1r4q4h2H
AjYPvh3rkfGxPbHMookrEqjICJ9vuFqWnjspRqjLpeSPSCbogCC8ixWbP9HGaZja1D5+Zhk+ztu2
VjInf3G+y4qHAPUcXuO3tk2OIVMDfjvC1ltZtwTAOy18K1yK1i6umxOmYjcYvaLuSXvYMqkilYKk
lidVFYB+g8iZbEgxQqxiojhkUyX2kj5A4/tBkI41B/ey/i1QBjCqPnNHkS0maq1FgqklixVzCfpP
zqFj4aZYoS8xi0IjyAGJ4fym8mVq+xOU9qnNy67DC31S5QaH0uymQ9BgrdRxvnKEBp7O3u/tNYck
v8njvTQIXIhvbMrm7H9rfNeIUOSNhx6AiV0v/IgrqOt2cR3DNMCTRv2Pv+1rGAZCo/3miUjkTOje
Q6kAzOa7fex/KZzNBggmCQViMr0BEM0D3aew6LHgtoVwZm7tFaBxUtliFm5vUyc8vFFXUDoIifZA
eJA+/jg3pMdzM5BD/4xf01KQdbnQTBEITGxUA3f/f/Wdbf2Qo33iMIE3Eupf/lmHAYhyK7oW5bZP
GjXcPTQ4Af8TnE2sEEVQA5PnrYX0JjWgyonBQjods2RrDIXVh4nwzzgPf6us5cr+IyshEFCrewkq
JOFZOBOsvTUS6DJ7VN/MVhZ0kLVp3bOWZd5z+pHsu5udaSQzUK/AFReI1j39sPQGej4sg4FxNuO+
J/+g8lTubvXvKPMEGcCGfrMV7Z9GfH1txMzmUeOVrMi5vvInCYZb5DuwWPy8u4Qt2tyH1ZytmFZk
ncp66YxayQg3qLdbarS+A9wFWyrYF/fBmk06jA7mp28BL/qV98pDuuF9WVwBCYUzK7bjM5oUFESd
8bjG5Wr44Br5meyX4jO6SI5nuDwDLz2hw/pTqhAD01hMxdqLNwkJSfWfxosShsP/2CMgPG7ebnCR
PYaCAfR1XVY6mF58H4su/fXLIBO4WlkCWGWfnG1yt1fhVPf2dlEcuIirZMvz2U5HaMC0lFlXRinu
dneNV23op3Ix/mcH+/S4sAfYpZ8gnqxig0IQVViWHYBJBFC6ZlU+ptJqO0919SHzKNwEF1Qw2fPQ
tMXiTMZiA7mX0GaV3LbM4Sx1N91pn1amcGbs6wc4VR2fQbYpaFa5zztxMkGGXLhb0XTYezkMwkhI
zVb7ANV+swWcJF5M4fO36CPR7GwakOjva30tZOuSF6Q7sEEwjZGoQi3CsHxPK1uKpd+bYNopJDOL
RWg+ngkTZ+jPMFsL8Nf2WBwhq5XCkM5INBrzhYIWeuhW1vgGC0nzQPANEVX6X3w/I9MQgAGZ3e0v
rrKDCOipU7NQqoCGhcn5el17WjYnCB7aYTWFtompO7cMPaCxMymsFdUv3HyfwfH6pjFvuwO05F4b
YAFTc8SBdbFd6Pd4WRj3bBRTBTk4IgiwMJsiWNGEVK8PrjJgdoGYkRnMxlctHqwX4Wr8BSj0FVHZ
/UBmjfXzrwT+Qc369ZwnsRd4lE8v6iW3hSry/QZi4tiE8AVdXJ7ueSJYJiEVzZsM91y5FQKd0nWO
2Bb5+3pJO+VLnyEPTgbujcALGp1GG+uV3rK/Ispr1UO78U2Dgs2mwwaq+cHSwr5ig+hVjLPv1agG
7hCd3m0/Ga9zeAtW98HJl3ZJhoV0BQewqiCj+TL0wUZnAmSWg4sZm3V67AfyefgFn9A124mXTM+F
R3XTOcrz9Hyahk2ookUtTojMQ20YY9eAYD7KLgSmb3493q1xS2pa76d+hPfujP4t/5y3vAUF7CwY
PwSgGburgjFEk1P6jIHmivQsKzhElDJtC07bOz8hpg13DCwpm7kpW1Bcj+HYw8QPEpP1ovHViORB
JEpN/xFe+kSm8F0pEsb5LeV4vDeiBhNJRVcag+KiYtmv0gXu9C6xPK/HTWDIszZFISRD3WAwKz/Q
bBWSPHfVB1C+S7RP2dnaHIqBwMAIZm5+5MVHa4eAfnY1lZn1DyaSjlFspbo31DoQFDzIRSkgtfUA
wwTIgV0cwDnvUG/qjo5lmP7g5fF+hbK7v92rGkMc4kKszvEBGXyT8WteNLzDLB4bV5PRsrP2nibF
BQHpdcyxEwhKEakiCHboKK28IGHqDPk18LV8d1jOPTZ7rUn9TAI2OSFRIt9o83qcmDhvlORlejiW
30wIdRmF5WAwQaw2oQ1QiZP2yvEzmqQAwdX4SL72wC8jt6lPNG+oFNv5WfYCd4d5dxVGwbKGYyL0
lkKz/UMpOdsqYDYrN9zMi+93xZCV8330MljWQxglJvfnP7x8J616IgVamFVj6SiSnGLjAhducgor
wjFtWt17cuD5WpZBGs6ifVBS+Iq5IyeZ2PqlDNMw3y4OBPiyVYHEbu7rNUgi87ZCNDj1VoOjorrJ
B/cNwXyjuK/nPUGA6WqEiFWkJt6+npOAmiCIpxpyWZ+ad5TiWlmd12YRMcZeqjnC+cwx2gCxJpws
HOLhm3+LavMekBaz3Qymq7eFmDadV89zJWSlUx/lrShWpt5w3bfb8jv6loymZdwt4QtCjETLVZUJ
5l4S96evr9WtW+KFktEZQESwBqmIyklK00L/Kc5urq/d+tAk3uqcBGcCG+83uynZ9xZHUDiqN9Tr
id57h4iurOAN41t/kolBq3Gt+QCBSvp2drnlwYeLuDpagRL7qrRAPe2zE8dNCB+a7J9NAWhFxWi0
V6Mbqi1n0KsW39F+7Snnb2WcchnBCG9L3HkhlcD2fziMuyfLshOZUGtjyfYa1XCCrP2hVmUEh6fK
glcvXMwzBs9QgEE+yRDz4UaVA/7jhqU6LY1EXz1dM2EvkFc4JdjaQm0Fi2ICMYeYBXv2zJzr7b9T
a4F5g0ZZ9zVuej8z9ShIRI8IpyfYztCxxBqji4w0+tLSutde+khT7SF7hnc5n9h4Ca8bbeM3RWGX
LxBKMoEvO4pIevPmbtoiIYDz4EcojbSjaHAYnKo55Dz1DFr2AqWospILT7dXioJp0J9NvuIH7ylh
PYLD9Qd7CQ6YXmNtJBwJBbl31hmOgkY7J4jiaNbcw+CeDnuX2hfTQaANAjRNv1MSx+oUH3S4/SOB
cg0GIIBY7TpXhdBIfU7vF6T1MvjEm3afGuCrcxGqUn6mr0zHuO1KxLEosRCm1x8vQvsjTbhM9hH3
A+iDTYPRdOvFelZ5qccmMG11ciJD0ujzuoQ78I9TL92FO3s1HAq09xMSVFtDimwP6ZCPXI446UNu
orRtiAeM1A2NQ71D2CJt/K9vM7V4la2lyPnT9paxfxze53FqqkSAEWCyqxCwvHe+SvQFDmBN41KR
ZqrZOWiBg7GTK6Ybohr3gwBDOliz70VaINR+t2eHNknrrTvGl1S/fhGBSWm7QeEuXE0wFlfVzFFa
/fVLazJ2ors/BNcrifs/wpgH1fYEJ5cGOUhDvjl66Pe0Bkd0CLiPjv5o71SLqwmsTVfB4QinR2na
ZG1Rsai5l9gCeX3tMFi/8t7x7z+6op2cJ5m0H3bkGUpYBVghBwh4JpHpYBAcdEVVKf2q8rPchP4P
VCSEsTnnFacUgz55DT7OUU/49Xc+EE2Ev3LMFtepDkF7r3KIln6Efl5YBpSjHjwQ0cUHoWs/XfJ1
ap5YAWEgRGcujSNmu9A6mrrL22VLgipqDlrQH1HqDOBn7m6Cyp7VQrLAZI13p7yO+geVLDeh6/Is
XlvMsSYHPSwjPaMcyrLWHez5yP74y+dP0K/f28Yt+lIZXVuIc4TGRoB+CuatAGmXFgRy//QD+15g
GSEueYHhm/h5NM8OAwCIAPy9MPN9dNlvg8GHfvvtkqxvJ+FaPCbyibFXBTFIyAO/TYpOsDqXTaO/
nRTyXw6eRMrwGuaHR4biC0d2XsnkPuYqWdzKTDrp4o+m7fyUk6YAMpF6AdElt4ACSYvWr6Zx/vDw
+rCj4K2rG/tVBRS6xF3Qs2/sCDxPGKryv0ZkLb6pMIB6eVCDvY0uBIK3oepCuF82zMrplMM+3P67
iN+qiYmAkZ6Zc4iMfztxkSm86k+b7raeXIvEruCgNHidJePs4SMsHxUlge5BIUXdQS1TK9aGntkV
/41KK8dGLlLbiDlamesfoMUVwSTfFsJtFHZNzdv2VsEo7DqminMRD6AgVoWbmGccL2juYNEgqHRv
TCN7JSG9u79hrk9Qg20QnW2VsZiP+NxQ7z8JXJ6EnZFCIMw08ePWUF9KHeGq3b8Nnoi8D0s+UxC8
i7S2GLGudfW/zExwXNdDTgrajzS0jZX0Y+uKLro2UG81Q82UHWfSoeWwcB6SPQM7YBgU46Hx1rAo
8vprU2RvEiRnOdtfCftIXlQOr8ztMSEVhSJg8JLK+K81gzXVwc+hzrZovS7oThrZD3USOgKJ5uxx
DkTyFsPQHCEbUw/WItAJoUn5H246SvzqRiv+CLZYbOGmILYDfDSFfqr9hwn3XJp9NaZFj2uYf3Ir
Mcx/h2Y1bhKZv8Yyxj17v9pt+Jf6hZU+4I6wFboNJz07GAmwCWCyMReICd8exZEmFOaNW3lSAqop
MBw781npoglfXT/gCQEifWr5k4cKDgNEESP1XcwcCvcnRwmp7JJ/c/DUn52s1wBQa0c+tfIKcM3Q
90eBA4BBoLcXvPCk38JsX/RnrdlzZ9QbcXiQeyA2Tcp1TZu/O6wA3s3XtoqnWZIJqLYasBwZzrGq
sPFsl/mI1vAdJAfufG4i4w8JVm6UavM971pNjyG7xu1KwPagtcKRApqDwvodPmG478Sw08koAYvo
sJinlXKybsgU5VlR8sKJbVz83Txb+OWLfqCnYLX8dlY0mpoomqyEpEZ0OrWKevqjkc3WnzAJDbsA
rfBHBFFVIsOZPa/95jleLSe2KqUS3kX29SEiuOMbjiIwVbkhn4zRi3l//NW8sPstHljsigRmyuRY
41Sgarmbb35R37upMrbP/ytfCbU0aC/JSol+MBRU9r1n+dXCyRrcgD9FgPrvupfmMNXzrqaRGlOm
kNfci/SCEMyb0HAwYCGXbGyFmJb4Su/DydM0SbR8CDS7zk+KexlnyUVSyW3Hy/07f3dtjulsFFH+
BctFa/j8yC5jB/5jGicAvVHD/aN7kePU/H3jye7OYzTDKBqY8N+LZF/7Y0TMJcvr8eLwDvnuxsEl
4Q4jb1VzFbxK2S4XNtSlOMHmiw39/Wc4vl/ysQrm7CYA2ov/mOZ6ikb14dqLFWrTWjyty6tnBkpT
3MEDQIdPnKGWcHCaJ3VHCZEDzwu+vQDV15KinZ9KqAGDW6KOHCKvsA4BgxBhhu0kw1OSmO6N/zsQ
U+UCyf9EviXOkqL5tSEV8sb7+qiy5jw8xr+4XM4fbOeBN/dbHraX/OoYH0Vt7ETvJGBMWldNJpfn
rEsn03z0HcasnQQRCdArGNCkQ0ew1pKGNur/y/WUzfbBHh6PMSyWQtx8BCEnFbxV1A1qos/w1R3O
72UqvUi7sLA+uEFtvOejdSgeXYrN008brAQTyS38tXW2yoBcfieCKrakxejwkg0I8192LVAjeTyA
D+xir7ZmXyUk2h4RXzfBbkjfn2FT8+kAyx/ktYg/sBYX2irqTh6zFHNWUuQDvZzB2i3LE7WeWPiw
34fioPJEtzoyRniHm+3Hnvs4lpPzq14vcqhk8P0M0DMeZKNAdU2fn0idWXUr6kwwd9VU5p2MuiK1
6JeiXKwf7nc3xZ/fBaYYN12VkuEtOgDjfw1gDPvZo3WLseS+ElY7OD6eHr+JhRunTQvLyH0IWa9w
t+rurv3JXT/pSTApyLlOF8KHL7ac/nhu3v2R+iAbPyS6Zt9HD2/sSs8nO57yeDmEvxRlMPKKMkvA
DiGC1QbzdMsrqGMJSY7DixGHnEQNRE856AyGexh9CSN2KMKV4F6y93uHgFRP/oDV8s85IEz+NF8s
TO7BH/TZZACu3mV6x3FCV19Va+c8ISYlVNr6vMX00E/TD3G7E80PgpIlPwS9sFEVLw1fzOQ2qYSp
GKzlADfr9apdZymFeSiFLZbNj2MaWQTfXtXUlCHBf//euTv3kUeOKd7XRpyCxECLFdrwdChknq3x
y1jOyhQj/R7jF1QxAWJ3KN0kN734oSEYmDkL6OuZjCv0BchSpHG5PSvzHWKqqeaBRMp8GhKNbtWW
NbA7KNYUt7yd9wYRsFKqn8q1IMd0TicZYVDfSlyjghGvPfXwHaTBRFFF+IlDcr7jUApf6Qre6+/U
YutbKNaWxyQ+y/Xedoo1v06aT1yYj6UiiGnUQcR9mc9Ymz2yBxxyuqK4f0Ol8d451KP+BaL8Y6BH
d1CZ1+N3adnhSkCD45yrU4PfH3jXciaiX3SkvA2U9dlRhwmpKceF965FqwuNBCErA+I1ZVH3RmXq
IcQ68cRFcNLQ67Y+qdUwYLwSd+VGuQrBV/l2Mjm6GC15Zo854eQ/kBwJ/83eho+1vRI/Iv1wnrMw
7dMLVAMJ837OFjKXfp9j/CxaO5VVJYef7PAYThB2cyY3g+ro1592ff5+IMa8LV7xjzzHXa3SxsMJ
TsULExSBbUbBc6buqFKoP0U5kWaQhfZq981+2U/T2SeYKC/Qipz2npzCEmrsiDv6TqC+dDl0fDIZ
aLOKFLlKpd/ZxXny0HchaGGNgD1Sc3ngyBZgCw+rhLUUX3mNtvhisOQfV/uNy0gO9eJtAR5pjIQZ
78afiV684rxBfsqhQEY5Mq9VJC1s/mxc+iilmOxNTgdvP8VJ1Pdmu3rNpEajeHUdWjgat28xLMkj
CwKUuyA0d4VFzZfdE32zYpJT842R6oXLCqtfgUCUh+bwXAq7DFbBTbFOhdPeCPkOXI+ZJy+UBOYt
rLIqVg4q0+ZsGlIo0zKjL9cxcq4fIw6NwVLEqc8FZwhmX6A/JA7sZBvU15Q9MjlSN2EryPl5BuEv
TyzM9Uy6hxpDqWYTZcHoAAJI3AjAo14l2JA2/kpR7s+mvv/5cR9wFDSyTY3CiAqtFgMqyrp1oJLa
jLraclPLQcAM2hmwxblg1bXMejdpHp4e2fHzJLNkJfgWXHOWH6iXYwIrXqnqonIYlMoQo1qsx3/x
VJXbMus5ZmYCkcLn76smJfsc1k57lyVNgfcYK4QncppweMrYQCqpJVB7xdVpukF/14hiqKUxIbJD
7EwvA1mrol5JWrJVaU3WJI2ojmXFOd8PamTRQewgpitDSVmBqXjv844QvBTfMgi0LKZHJaaZxxXD
IStHMOSCdH1AyvWBtQIFhJzoVh/5BSO62Gv6wGnhJZJqeo05yDg3AT0ghXcqDU5Wcy6gCiRECznk
cV8ru2fi2Wl57pbS7Yz7zf79lohRqr3ulseUm9BxdvzpVNr2eKQ+aONNzu9zr6kyB/sMZnFJkVHX
OVur6cDoNPtX8WlL2xTgnWW1TCA4TxAvgY1A7fBgvPwByH1bhPxIHtAyg1XGBBa/93nQm4nTL9LR
HitZSbIqui8wkQjNUypKbFBtCWRLDtMvTkaUMPJnXLfF8D/Au0pX8CeLyetKN16bdy1NocrG2tf2
JeyfVj/i72YCOs44Uu6P2Eshphnmtq2JnyEL1zqX1bmjVUAbHs9D7pc0sJEig6kMELyXtr17cqv1
19Ck4OHZd3gvtHB8NZs2nasfe+FjJk7Pmg19N6k66ZhbC6YrqQOlNmLnFPhhO0/gN9LhQYfYVgkr
DmegFQpjYBhrj9KB9AmmugIdrvsBbxTQ5Tx75H/Wt7QgG4esgg7xXCXNhLticYvBr5xXgjZs6p0I
rpXE+xm6pvLwXE5593DtibDiCILUDv0DPJ9trTnWcOmxZmmwtcU26Vhf0LnaeIySO/04Hh7NM/Bb
a6xMUF9XXiN3FAFQP8i3ITXDo/3w8g+OqWafYeRmj6HCjV8okA5yXrDKQ1/flCDeC7HYjAziqkvn
bxMjHd/gIA7GghazjB3MEVjeJ496r8d6n+6Lx4l8q4oZBBMPeXg54Xs+W9jwz4Mk/Hw56/nT5gAZ
U49REP5E2fsPb36hhEXcvGqka8DFMwfwfCVNmCQMRNB6kyP3sfDvm3Gf2FdnUQFRBlnUkKT6F4sZ
8c7oNMTk2x39fCsTlwxfHvpknbXftY7LfWegCevp4SCMW9o0hDZ4HRtaFKKECBatJdwBaC/e34d6
YXgOgttP/FUo85pRJn/7gGmNgaGqPgsgz/3vmzBRSILIjrfJqiExwH3fpeUKsJ/2HAxJniV6rJGY
FKy+z93xcHaLPXplfPvufqf0GGtE8NLQ7D/r/INg0GF0GcUJBQ9l/BC/8q+H5WWpiITVhvkQYveV
rZEl+LytOTn+AjsvkNiHbectwR+bUv+E3a9mqGaY0AMBaJOpe6J9i/T1fgCLNEAM6JFICh+GyhEk
419i0dJruxQ0HsxzI/J7YEFPI6wByxv/A7nTcXANbzhNav6rYxGdD1QdfR9p2JrnoISa7QKx5Xey
CVJzNScgWFEduc66J3YZ1IrmADM2I0CKqIpDuPVo5QvFBEcPNDDs9cphw3ZS5hWyBrEISHGptMru
8eGV6qbBOSD704odGoHp4WFHYr62k7FDr0rWCpi32sQt6cCHOBRSJO0kCpQXFwjlPQe/tp/91x1E
tYFp9zZd5h5XwG0c36ULVSKIFK886gLjhJEf7GE8kJgH2/F+nrt6RgPRgjVE/keN/x5ZM6lP+TK4
gEBzVt1sEqmw5OOEfAz+oBKyA3qMuqZPsmnfFxqOF1CaVqPwnaeEwRdwX8q3bpak6gZBZ28rpn+i
IoK/EbxKIaKVgSKK45PaiXdK1+mF6kljNmIhbHs8nJrKgCPprqQIe9ME2R+pfNAPQcA/pV1qLYjb
N14Xs3TmjG3X+6mjKy4okfwPFs370LeX6P+1IYY6KGBwSm++W1/0uC0WvF/LiPa7cJZoXrHjO5/o
UkXF2cHiOpVWCtH12jLFZSzpgG6yiX4+WKYE4nL8ZzlEMQJNHs+J3AeWaVt2ozsKJDn3MhaasrSf
Iy+eDhFNW9jR/RR2KP9YcE4Lt0WB5EOWfAZ19QEbyyO1vAG0iDUa+StjhruozuFWdrpLGIC5w9Dh
QlCG06j0PzO6VaD/ph+ZIHmxbUgM6bk2erBJU27pKvekDVymGx8OPBeGQpf95G72GY+fgk8He+Fi
K1Jc2fLBiOqC1JhFjYQsgotMJE9W/ZnxGbl3rUFz1Drtfq5UvMZADexSRByFjWsDu5coPt99yZGQ
cD9cPwS1WrXryv6XKKnrlKCqzxlXjfsbSSc+u/EWPw3kJXhZ5gi1LeTXLKEGqGNnRwbLLrC3K277
aeW6x/vUHKzSsQJiSg1+g1T1hxYoh9uQLZ0ddLnaQ/kINCRanQ1se2IjkyZKQtpyzTOuClDFn+t5
7ABilx6ljONhguJsOlKXsptZvcWfmmJ3h9/FwwCq5zmOXe7l/f33Yw3Q/t+zy8cJJ2J5Bx6clRH7
hpCVA6K2hzfkKxYsZYb0uI0yw9wTnP9odKHJ3neWbfa7QZ8vsZfiDclGhvjlug+iP1+mafEIE7FG
6/ppwx3HosLnyOhrdMdiGMn30iiPXbPadch37+LVf5V+rwLFsGPovEM8cow0omXzqTFzXMXW6cAJ
Db586H/95KDAR+pE7/LzGER+XkaL6dFev2HtTEj15XO7spLY2csRw7pYYODY4Rsvxoi50rgp2vhI
cyFTN5SKe1UF+FJmVx+0Mg5qBQ7RqDhZR6L/WENjc/23P1pz+q0LOLusw8g/j5GnVVaVrkbTULmy
poM09JmydJigGDxh+NOhHpheI2m0N/1ZKh3pi9G+3Y63tEhN5Xn0hyT8TPtGh/V+lYQWps9oohLz
Pb1fjW/qsTGHZP8ipUbJE/hQ1US1jlcen8DU3wckwJTdzYE35ho5o5Xx8Hm23m8YlVqFguNRrIKZ
X+a2qfwg34HVzRF3HlhFOwhYfuhMJzy/2AwvUypjXtD3SVaWmhq/C2XFDPZ2PprBodHilFRhQaPJ
8YmPQtH9diZT85Xdbh6lnagVmYkc2eUHOOMZ2YjALA6A1IBOfchjD9AyYYA207mQ/VZGoC/VWW4G
jTybNhbrKITk7+A4HlCnGnIy8/kqk0StYCKlz/K8i3UfcwA09KG3NcmjfQQlIBgFWE+JxHLuC9Nu
IGlFSAqkaJAt8Yyr34a1ygeCSnXolASwCnFVgLHgFn0BsrxzygZ1P6/pwwL6eZxhzyhbwXT6gunD
qIb38WJnmbbhUMZIAH7imww2zFQMWd7r2WAVjR6AnKrdtP222eMRLVLulRexo3c3pHmaSZMv2x4K
d4Z13EeA0PxsscipQV2L2m+o2c91BIbwZ+UhjWLQI/hFYXlDBAVNGxcNWvwjptdiL36h5Fv/0zVY
xsfoCn9WosUOQV5GMT5ilRhnkFtaxuHkNw24pKAYSdc8FQvIy1fhAu1IS0jvgKaL8xM4ngIsLUHv
HXz4VazulbP0L+V3siKNNBeBE4HC2m3b1Px9Ij397gfutpCR+N/nRyLe79R2oM4go+0xHZgkCUx8
kLMpwThnAfBFC3c6ubIQiuHyymTajv5M7K2G+Ykn3EKMeyEPFEkTEPzz5YYY7z0w58XTgJCET6DH
We/aO/QE27XAWhB/az76ryEiWj0OwcxiMEY23QKlrYtawLMyZ6xFUta1kOB4qQ31Y08rD7Ff5KQF
X+IJTV2F4dHm19cn2vJq4dxObn8+Xtw9F6sUweOyZHUsLTT83c4pgsW5CFHhVtG6+Z9iHtYBu62G
h3TG7bQVqY/TB7w4vO3I23KLUV6jr3ooYscAO/GofGryuaddgYh9CaNRZnFukevm1JmF6DNXz9B6
0bSxaVPCXAHvqiPJn7sZZnWTMHE6SQl28jt3dwNg0tzvZnjRlFDUqgze7zDXRbqMaV9NY16XfxVJ
qTt3+ykFIpiyFdg+kZA18fhYIGfNa4M1JtDFeYmDLMzgkhXbwx/+vdecMZUviGlGLOaBJKOkjMp9
VJJUcKb50GSthYJVQyYIPiOxAx4TXphybX6xu6L2wN1Gz2zjF8mgnhrtAeuOKjgIjP4TX4bDX2Am
DovBMkH0SIjk6KBK94V9Upfoq3B3Tzas1XdqxqQEeXbHBFOiGfy6Qy/eMC0jkwRfFc7icCKS90YC
HJ59hq/iCJULmWvZazcEpX2wf3k9X+VPNb9pwstOPVhG1Ja37L3765RtFr5j7hJUEP0N3tb3po5F
jrqJ0Pa94RjPlYWdBGoCtM4PFIe+vXtOH0JN0cB1e+vvsvg6+Oz1uNPgQ0+RAb0InEDNabGpBYv3
vaQbySGTwio+nu1EEx3+rhGpdaojpemgov7/sVQIebu3cKXlJ1L/mePaNS/ncZQ3OEZf2HafoFj/
mfWRt61NnXuRIbN62ECLAZxOKI7DRu3jfSFcGXknBa3BIBhRvsbaNajaIBkgi66HLuBuFceJRauB
2VgaYECijTDzaapzmbLYQbcmhlayBUCeJVChufydPuZTP/AtZrElZ4034jrekxxn54brqJ5Z4tdV
QVKcy5vqm5zUwfmrBC1jmrw/Ujn3y37ArlL7oh9WGqblwNUsmRsPideYQwt5TfEh2pDVsEvSDn8u
lPDn5oLrQ/maDZ6ndzHNbdrYavR7AJBmGAzy9e7LHBrCeQKnE3HpS4JIJ/LC3jY/I0e5t2Wkd4tm
STvpWg2GnXiEc4w4EGzXDDJ5aqoSC1775UVsF/+2Q9O42gt86ukgautJXTqnq2JASLHKTGJ+yi8k
Pmd1ODMtvEkQMpTqvX0/vMZdFg1yug6GjUIlYGYZINGlS6581b6OzZavFJfLxMSuMny3cTZoSvuI
3s8zpRqJeN2/l4Ru/HvWsBAIkXztRu1Khd2UyYhcn+E8gh6txgu8uHRLFN0GnLhhlD1vJgNihRaW
lFL+V3qrifLUNmivsbTMGAgsxgi3zpPD63wtzEwbpFD4jQohHJRCLgymg074Z3AN4tHKt5RQuucw
xLvOR3q90mrgvSCIaaPKO/ksDkESs3GyrRBocMfSmuDke6CNM4+bjrhf9uxCTLmY2MXzA2x6lqHx
n0uvG30H07lyC8GNWO3GQrB6KTa1Errls+IF8DSIJz5fVSQj4gbkdRXIoFpV08NPUpRXO8Sqjzve
2KlPD75jmLb1xRHyYVKrwUdem2swH3qntPA4b0RnQS8OdK71AUqEwugJVB7nuhhT6wfKMfKblPaL
ciAvoRjA5VKpQ/59a8o0Ks56dPeAqs+N3Hc+d7U/ars8bF8TXFllS5ai8DyD35Qo9qjuMN3AqJ1D
ezHhC2utWKnOZaVpX4c6j8ySVpaybR9MwppTDoZwYxz8iVScUJ4xVNUba5j3d90m+WDhkB3293pQ
EtG+RmwgXTwEb0i0zylkqiaCqg3zY80UIciXvTwaJHO4Jrg2BmGdokbELL5DcA/pCidrKbjPpaSP
1p0dpH3L71E3zo69vEaTi8iX54bBgKGZee+5mhaDQoskIt9xYNGuKmKkjZc1d3KGIvs6YaSVifx5
rRFizPSCNKn/zvW95qpKGsd88aJ1GT3kCoWKrXG1Bs45wf/visr/jxnBXFE0bNs4sbionK3jfFIG
v3ZEFz5pMtbxMc9QwpygTF0gVs6C6qbnxdNpXo3lFj+kgHoEAr2z09A9XS4i104RJgkXdV3DoPIL
wIppYcUfrH1Xg+h5kC+wwDlRBKWiQTI5HgGARLk1naMnGctdrUZygCoIRB1oioyIROulQnOReYRH
Mx2Ch1sKpDH39pzPJwOW4ZFMc+JKFwhoA1V4UhH57Bd7PT8FEr6shgKaIYYXdOFywD63BVfmAYTt
7syLwGb5NKzIpAOVFcCCg1q+Ila4ndPJdgonoeNHt74GY1NCaV1Md60oWbuZEzvvZR2kNJ0Ce+1M
v96DbOcGw8J0shuJLju69089ziWkbzdBwHZtLO/5DN38QkCDtqisslvj60KYwflsZLj45zo/J0cF
SYxIs3E4nx7zLDSDhiwnCVbrWehSNfgwFWd9BO2mG38wNIJUZI1VQHzU2cVO/jqy+W/DYrUUSl+W
6zE2XIEIIhYJkRNgCnodkp1PnF7TRcTIMBtbLj+DaKNveYfboX3bbsis5rwq4NSYV+KAgilSd4V+
lA9QgAnD48FrSWOSYGaQxO4rbdK9NI9zsJBfsAUTs+D4afmHtZroBIsRoc8i/mqDwByrwtwtmgIF
ochlibMB01taA5em1vLmG2871g+NfwDqAWMz7JI/ZcXlIdsQvfU4hHNR/Mq+iixlrQgddtp/pYoI
KHZFEfFkknExg8KUXzlTV9jMrZBYmTPRBBhFw1Pgo8ZI5Ox1LebQ8urZ5hzrcI/aXMGxnw/xZwUq
JaD9HSoZbioIKQQMRy8pz2Wv7qJqzbOAa+/8uN4JY6ipWGr22UmnrEsQ+P6esXgL90rsG3dfWouj
G6fue0uZu4iCzPATkbf8jKj4sqpCTWvEYwqg89ctGp/L35N4Cxu+ROoNqfSxpWB4Y5CagB29v6vB
2jv44AWl/u2HYzf+nogB+NsXPx8lni2Zmtv8k1YDIOhhOvYcuYIirgpn35iWLtaBfEN508znPeEo
kuLLr9UEAjxEODcrZoxUQXAdsqb6CGN+qP8MZfAdwKMZw2XeI4OSA9yWiTl+aUGs9kLPBpNie9+h
skQsZgsW7hdgoAA/euO18zKpaDV6gzWyi65eZ2PYknawT5Y/Qr69sziX5ThftQ59vEtCYMq4GjbM
fxOsPI6Fug7zUJNTRMvNInmfawLXuRjvZlUEvsgSuX1TvyOu5YlGl2zj/WRV+/Qy9S7CsgIhvMwC
yjLSqClCj47OUufQWNSLyr/WZChVcWzYMuUScN4wpAd9h4J0VSEi/7A4io8mlkf9/DmsKOpjQZAH
UF4IcQRwY3WqThZFMhWsu12zdhiQVIrOzijkhK+CKLqBX1X+LcxkBl9mlE76rsL7MgaNcoJyFq4c
Snuen5hhSI7GKSTP7BJCakyGkYRh5J45lFGbpeK4LUFbCJN3MfooH3Nkzz3nPiB5zjCaRUKRfWY1
hCBBlLqKBHJLbbiG61NCsWu+f5psjXr/4GdDab+8yNI49xCwyPLkkC2HyNtBM/XPuEYfpF2wGLCq
A1YupvS1RCPmOTmgApAtHchXrzuOHYTLJnCms0GyOXL4/9WSkRLtqz9QTFwJv0YveWXO6l7FLxwJ
O5Hu5gjZwgUVfwWaptTZPxQh26YCbxwWFymrl6cU9efanfk9prRIN+VgeALDMNiEQDekCmVPawbF
IZZlmc2MAKV9JMjJfVd+X5qOsTpBIDWDVauSVusE2Co/nJevCTHsL2X/NvbdmU1itp3WPyBMU+0i
DdjIDh8h6K5yAd1xTcIwCwfMg+rWQ1fKblVm6MCi5EHAxJdjAO228t7zEp4f8CEz5t0GmkR1Dmke
1jLmUKGd99RY+gIymhU8Lt+oOckMkn/Te/e99kSuiXbFyY02nYPfZTu/ij2/0qRhCdzzd65kXB/W
str96RfssBQ6odpld0zuQ/lvdKMhvBEb4/KsLqEYaZNjK30E5wgPPcKF4ucqQ2Rv/0FSHrefVMQb
EWHvlaIImrpPJ324EaDi2AHqEYjUyOa3YCmOTNxJMiNZ4RouuRSUIH8rdYo1/LjW2f6K4JpIxOBD
Odxrp2c2HcwXTSxHs91/LEyj+ZpZtkLvpgySp7PninEToRuPDBDN08N9pO9/24fOdVOSuDnKkxOc
NzzRdcJsTI+T7fpmWahVD0dn1KL55dxFeC7OszFb+TT7OOr9wvAb/dmpIb7OgU1/eJhMGXUPJAXU
V8wdI7f4rm9EpsGw6LqlhFL0vBkzyLwpj03oAkKyLMSh6iYtFUpcKvwbO3q2ZDJag2gGByuBT3Hw
dZanswd1hLjGuBymwBw9WBms918IZvCyWzk0idyu97gCNDi9DsfD4kKNKN8djFPFamaZVazcqzuF
ISyNGC3RQ7FecFREXm5YzIChq4v9LUcbdZPAOtAccJkNJ28onjo0AlR1XfBoUoXArjPTYXSYCk0x
K9sHoW/ON79NNPx7StdMNczWVSm+VIm2wzTHdXniA3l53Lp66EXzQ7EwPEjZZKLeZ+JtDLnuHRh5
anR7TbKjPE2htnOte/x0RrnW7tIA/OwqUOKfZTjojqYEypV9YlpJYqunSw4p8Y1p3nhagesBv/nI
GshJhlmzawdh0+jAHVphzntipEy8+OxmC+YH2WoJRoLPWjLqAX7Gtek9CgxWIgZ4mFjJvKvMVEXS
EyQ2EVzFqItfEYG2eKF6XPVYXjzJ5I3fFYv5H3EN/fyKHXf+doXVyNPyluGLY+ToriGAu7LFqE2w
V4Ma5L2X5VLcI0Y7WgrL6gGZODbqNKS9xHSR3ihD5NT/kYcjtwb/XuJSkyvWlFmC/809lrO5d8OM
3UUUNR/A9rroCLWCUY2PLLQzE89sRZGhIKJpQD/UPlKXAqzYqfsKpUrh8M1zNUzRdAEW8fwCYkD5
drxS4FXc7w/e2gMRkzKz4+lJFxZalSmXowQUpfGqiiz2XOW4ViytpsCsAuN4vZDa2qlNJSgngt6L
+f58YfZWs2/mlRWn7zlxvyhzomlVM5BveAoMg1KQ72TOEMqTr1TR3ZwBCvEuQA1HdzGiEXEKE1Ew
rFTkRHm6rzQqR+K5nfSjxLbEOblUNnVM3J+dgLu86QEkjo9foJBLycIXRIAWqSSAwfZrbzq1G6EM
b39Eb4EmWOKP5dVgmL0QgyefwSqfXC1ZAkZJi43KqAZv/CzolHvyAh8ATM3M33nFJB8V1cyxJoiX
hIKoa8f2/nnM6rtchew4M09PyQg4Brq1Xcf6YeudCJ1j0wyslGf3ReQFGT65tTB/ulPF+lqz+O/T
ULdT7pSnBfAUisDo+JUnILsHzmrdXCYq+KIJumxhcDySormGuodQM1VE1H/sAJjgZYlgecx+J2vN
4NEU1+SNijPd14Zg7CZGRPZ7j1SRZck063BM+JL5tDJj75Z6Hwjh3ZNY6I1cz+zAgB+pc4U5va7o
iTlWIQrSIk/alALcUZKNX/yjjDNWH+x/zUTO9MYo8QGMgmrnm1QzAp5IRTq3rZLfRwooeLbhiMC4
sz3hd+QLRfxmmj3gWtad49NitceI6PSmyIjo7Zi4VSQl6DWRdG/GAyWiv0Yw8VtGO5moN40Mb044
G7HVSPHfQJWCfBVSvumYs1UfFiKS9jqv7fxyeSsTP/rXFjNXAhXO3leUi2QBYUqUQAVuHNsUEqKX
MSEquSigXXkCnKfggwvzT4NnONYEehWrGbrbawa+ctapRUNspd92h8jfY0xea7PY2PRCTd96U59T
qkfXSKy2NJzk03FYumXn/8W/bC88IZcEZhyVPQShUJH7NS2INs1wtksKZLpVU+ZavCgj2DY3CmIS
uedNQGkgT8xFV/tmHB99QjTV6CN1SgHq4vkvhR4rtaCqOfZjwZaTz6MkGCzPmMicqKlkeDla8BS0
Msczs5GzDzGxXsCJp56vuAjcuL5zlgCH/cT+VhieZKr9+aqdmlZ+mmrdyMXmk6DEYGqTevo19CTb
4dKp1WQ6EKQwPcmS+inC0EAXi2BpWNIrfH/x0YGUn9H19Sm9Mjycen/aIYbwdRFnqmFwkKrBKZJi
A1QiGhyhwkGet8KgWFdjf5phboGYw7KBPxFh7hA0fITw9lYtTba2QvRBocRpP8mzPRheja3Xw4bt
zxGgFBlmvRW32yJih2b59hU/sXDUR1VZBudj3F599qdgY/+IZTKDa1LZ6OroPpkxqmmX2C9udj5D
N0mQqu4hcoBmAPl5ueUmWKWswplB3OJQUB+BKFVUXQUC1Pe81j7rriCYrYD0jsUZP2z1IAnlPi83
VVmJL/oPkOyswnT8yfIkto+4is5z90EnpcrRqvMfreGc3hwxsE8i+hgeUOOXSWet//0nYo7jDsw5
+ZrGV1EeUq7WwskydclkrajRBBm4SYe9srLoM9BPyS2zFYU9nPkyJbCiVe5Wb7owGxiogru8GPSC
HBY/1d8LP4ahQYZ/KTCbuM/e4MKxqCUCqRxmHPrEdFvFTtcZ17hMt67fdghX6wRT3iCjZMq7bAm+
/nc2eXuTerQkoKGJHFaO99y6H0ieP7X9ypOJgTcMGwZKH1iQ+33Q+aGqwb35cS453y9eCCEuiu93
b9UCg48Z3dOAx6owCK71H/YCU4pEP2YMT/EcDToju9BCxTtKfH1pTHAAtfVgGPAXVXDHDEWRxvNP
MQ+0nQFAi7cr1zhZ7KgANTPzngL0XOJ1rnod371usHB9W/WW07JOworhJ6eEchSP6WqQXpM8M3xz
OoshBvifbCPPSCaX/RJ83THl+tjyFn8bhRqSfjbAh4Rr7mMgFiBTYmSK+VAbfCoMS6LW6qgMh8ZJ
6Phzj4xX4cxfNLF28YUlvhaJxC5dJ/Mw6ELPKQ9FzaqxMsT6/INpKGE4RHyTgU0gM69jJHVRmfpE
MbW0J7kz4KMZ9X6wCo1/U9SJw1hPsG6L7YeL+UNt7SHnl09U07QT3Q8Oj4uUa9SZxrbThXOvM+rx
/7G+gCShPjHxenG17QshAU9NX7VBu7CSUQ3H4TT9KEdoSAUcZ1bxKpciDZ1HA2Cx2v03fCzB7Dow
Qc1j3r+gb9lfxXX3Lf8vry649m8JiuOZh5TJdnO59K972SylCHe3pzQu5xuoMMveO/dGwr4IJfsi
72qroTVgZZCYqRdZa+INMupqD9KhhQ911WFT07XkZBnrRYa66Br+WX1fEbazudoZXPkcLB0fSetT
PJv8OuBsDGMI3nC/MVOl47XEh1N+adsSmhpuF+LPpMXJxuHGWaU3KnIeOfuU1/RPDJ++yxykZkmI
IczU3GSCNbRegJfAYBi+4p7rt9gxZFa34vPjddYJeN3hFREtVPLEiNG8Ob3pynD6nDF+ydQL0HJX
4hBHpPJXsFktGgeRT/wi7byG7OuwAb7TUPXA0J25ig/qs/fel6VBuFqbt5Z4fYNWvII+AaP6hKir
2RJ0rnUUvr7Eekc8fKvLA8WUn0pTP5juib42OkyTwgF4qlmQazgQU9fSi+tycJkWUrhzT/etJ70c
pYbI4yJ0191vC4NGGil9Fs7NCXbsgwb/7+4j5tR9k+CRV0xsojBJkRb9YAFY6RCQ4PA1EiDBpPGE
jwNgEAmod/sZ0NO4l/tAoyUSmCQV5AnIl9UjDxZH10TkrRDF6FXaKPRTR0pOcwd/VE1TjqoFU7R1
VqxxPweV2q36ZRVTn0UzouejGNmEzLlNuPL7TN6XMAfrd8P0sNytJqvfW0o268434iWbxB7VTmBR
cLghoOzZ82bkkRINQt/BBUmIJHi9FGvbj1w5e4qStNNM1XgJNMLezddvRN2zpydMVnos3pOr3eWn
Si2v+DOQAqjYnQC9oaLBvAXrdMx4rbve0TARfE9ubxXXUU9pFoteDnjIXMsPfg5zSlup8YJ1iHcM
fWSrppwJBRz62CjzWa147H7+gSH18/hGRzQXlmsOnoDcWELDgvRYN8yKA0vB+NkEtRR1s3/XydVN
JZv8R8Xgk/pvVNYcj//itz3qYzcy481Sllmt/2rPd1FHsjE7ENs5Mh0R0HsbzArIsFLmsBQIplHc
+dauoRoUVDXC2Vmje3GiTLR2DB6wEOFlZ/YjFSOQSRlLPl/ybDLp4WWSmyjJMYtCVFs09nhFxYHh
TjHZn4pWvwFRwmptD3mmPriKov5hDau8I5IaHP7zHbIMeMkjcAL8oZctfDQXnwMDMPNP7Yvqx2HS
TeyFJ+PgzQk0XqSbzlftFafpKRpRilVt2DAhKzXcvoCLQQ+MQH8U3CRmfW2N3UQqiiv8bw4zotVo
sdp2U7HygkB+2/52i+SXv8Vz+eIqGwFS3ejasBZvivgdOQrowIK2LTRf3FDhyU0n+eboWacRXkzz
4j5k6XMHbS9uInRi7BinsxYlPmXyEE+s9mMai5I02l8HdSKrpxhKu/VNH7QHIWBa/cxNDgrWoMsi
4NlhdS7e1uz6Vfzbm8eZLUQQGXOEEJsqHI8AvJnndrCQnuM5+vGktm7x+8VyNSPOoIHg3/DgBq+j
/8jcOQBZ/5Ew2/zSqZGADCqj8ylrzYKV8JiPIqrSWuiCxvHUsq06UqNP+dp8Z4DRtAL47+Jrw+fj
LmG1UKxOcjOZYYUYiBw5R1M+f1DQdTc5R8NEh3g+JfMhL8IZL/EuBe4aiVjjcFbMTShBOX8YDbK2
PqMyKnPELFxu7+ijmbH1NY2qvrgZu/8EvwAOv65ot3syKe0KRPVy5n8hiu/PxDEsJGsIlF6ku3bd
CKOM3Zaj95Z673+qCvjqonyXsBISrTcjgu/rmmPLFcBXh/REcN/mhS36/BLtFoO8AtsqiQsJnHDf
1NA5qbIkhRGxr8YUwbhRe9fwIMwjNDCcSAtl0a2mwYFDxIbBNCXGoNGVO3YZSESafNd0lnqT8nYj
idzkWSNFRJDlSztBzqiwAxvOAdmVCiZneTBeFJVGl1n6XRQr52uvSb1D2KhNI/uD/Zkvpr5jQsgs
V3WepTuFEH0q8VXM0XhX8Y9Xc5RT66nzVex3rUxTvK0ltu53bTtZggplyZPgZWyNYlqAVKKfxc+P
7MegkwKdTIIKGAQdMQ4fX/ypaJwtttJVlDUmw1rKxpb3hlGSOicMZwiqcwkRAiEJ/36tNrTOusXQ
jKDUgsOPqGG7s3yxFJ4CR5aSD2r/igHFMsKAGGDXjeAAHJ/HqbXwYxY58SnZtOkzJLTCl5mX9UQB
03WiNbzg1qjDHBdRea3pXSfkGhVSlMVPByWwa5GJ8iGfy0kmmCzJj1o+rh9rpd7W9wH0O2r5Aa7X
GoDPugyi1vdOdCmTAaIJjihIdToP3LMresmmFxzqIvYzobXUo0Z+bASpwGju2kvS3NZb4D48q/pR
xRlAxNN7oM8Hfzf0iil7KLLboSFiIMekI5pcoyreUqQY2rUlIn6+K2Q/ZzaP3VThLJy38LG7a0pG
tcESba5A73EO+8BkFUw7HBUlyfiiKod/1vTp+ps0IuSImmfbCeBsXBsMoFZOvevSZ7CA/8Cgb/bO
XvydQbjt8b+3W2vdEHOBbbkcaUP0OpwnxCvuVdoP6let3TQpyz7/j312uOg/sUFERpKTevcIj4K/
XpvEzyywTvAr1PTDAiRA4ObSgI0/+iHN4vF2N4fuQqoW8csRrULR2nxZs3jcPNi3RmZHuq/2Z/AP
JuaZAC9lQNHLhGYm1jc+vbG1pyDMKcLeIJbLNWI0K58bbxOLVqIsmkKHcKr+YfgjM754UF7S6ABO
G5+qjGH05S+hYhtXoo7fez13jB4sd9YYiFjbVg0VFQqRCkDxIqfONmBFxZySj3GDV76Ncimc+YVe
DmfCkPF6u1FRzuznw4T2CML4+diAkDaezYhGedTn1L9vyQyKgJ98dP0mOtuj/omWLFEAMaAKm2s9
gqTDk03fR3IRPpl4M995Nc8ykyW3gxhRZTW5QgvYXgBme7sbwGtGMhN8CvHtw4i2okIE8ql59afX
kiGL+el3psUW+UmuNQoUY8qMIUJoP7S9s8nRCDfN9bMlZCKc0ilQwVxgD1rPGqcPUEbF1KAKkULc
NTAkFISoYd4F9qrZ4u/JT8r4TKWY4UO0Fhq+WT7oUMo0HIlI2cpDMgiVojHhF1HgWrM5HfI8FIZ8
Q8egWU2O5Lj5WiKAEWCtIKdRpoz1S/MUZhs4bQrjLD0yGHMP8OeU/ax9JkV3i8ZYvh3cGHDoJOHI
/O9evdACaecv/zKw7Tc+bCoKFq9CYpk+9lE8QyERneTREJgMhAGY+erFEEIDOv6uMMT1Bd7UAct/
AdqjKc/4tRlHZRTPe1xIw6yrNyg9DM+oe2l9VIUYRczLDl3fI0chBz8aoQW9Wq6NpLd9tqVOPw0W
VFuBytCEweE6i6Pzoa+9E6kM4yBPLmQRKcIicwD3FHHbSQeOu/C3PWhOvu92d00rzTev/IYyD7b6
fCg1JJcGf/lvPWQiFWf/DXzqHqzDVOpd3WopqxlsjfepWX7O8vTbf91FigZDbJk6Al/2Xd7lL4He
bx4355CRz0USZ5YVUF46y24YtSDvR1b+duEAcQVa+cj4lGv3brqMJiFovTr7nOHUgx8zYPy5rW4l
IjqWfy1LAQ6Yp2h+ChEJdvM/IwpI+BElGhee4+z4ZSASEVKiOb8CpG8H2rh42e7ICVjmd2DQKE++
aTFigJi4EGtOfcU8lNS1Nuw2ruVhsgs4jpe2JMjOnVC/lHgEtOUsGeSO4bVT0KgSIK1nAddqusMv
w6K6/0N34Rab0l+4XzJZRu1YbKYYzHLbVesWdk52PkzcGX5ezoqLH0jie/Stpe46hJLEoOWVk01D
ztO1EXXW2B+/1G3MkdBNgyZ86CAr0FMlvWhLa7GfALQdaXw0bo+JOBrcSe1EJLNSCco94aquDTT3
9VfttMJyhYDxG3cG6FeavaSIRy0fgL9h+o5n32pRD/TqIpIpmEWnmhRW5TpZjnsy2sdAZ1RqhH+X
WTYM9bbcOmfkNx+iNAHg1G6CSYg3LF9uTCbzTCZaI1jnI2oDegr4Md3s8SKcOj+xSB+UwMl9oRbP
KzZ0iIo1Eg7P/8QQAZ5+0eGAWLgJq2WsyIeH2KCmhLl/9fDaslePG1fWDCa2gTOW2GS9ZSgOXDNO
UtLrNMra3eFU1MQGbPFuY4kfmKFwJeUDmylomEzjGfvnxhCB7jU0Aalj4kMO9foBRe+IDowBBw1c
VZRLJVIWWeQzopDVHBY+yeNCZ0cGqyS2GrdBuO4J+zJnLIsyYAtmbshw3QAJ8203E3TdM0mMpJwC
HLvhk+ihFuuK1ixZkau2rpk1BKStGbeZkPhGjxZMwHHPjMVvo6r+y+iXUdevHVYFQJrhmywN8kyQ
eukq503oOkpZCR84EezDcMoe9G5yj8656T07ag4pBvIh+U+e9vls+8O+zZtpx9PuWPGpYz5HDYp6
Sn4SxJ4Q1bkVJTaiIBYhjWRE0nyP1ZBs7HwKFWnFcSoKGHeXyh86ffLJO3tC3PKBio1aGjFktwP9
70KsQKpWCm6dohFfVRI3lIsbcUjnVlFbpRee2NA0P7nDiHz3YV+PnDNTk411ermURoAvpny93Fpf
IozSQF32lDUxIwyUD7j1tGneICGVPruvglNTBT8qFtCbtDV5DR5H8+dBAMeqkiLpZXaBz6z3pOKL
HI9z+tSMzI5RAj0A4RohAbk+/AmL8U08dfvkRUz/41Dk4WkWk6BJATk1S1PlclYzL9MaqM5jOuw0
F1jea2m36mWXmTKMJxMXUeE0bQIg4/pWv6BFw73eBvHkqwuo9An5aHUcy2wHGUM8tLT0O86n8d2d
MmL3AEV2UpTSLUDTbbkoXeu09Q57CvNK/rjPe02BHlMxcAliOBxVlNm0rlil63UcFyLzcGvpQKFj
TY04QDhKQe2C3jWlzsC2Zp0TK0BbiSwXEcpHRS5TXkgBugh9V0C+db+n0u4IK2DkCmS7SyREvkxp
UnmlB/TyiobC+D8ez7iYu8qIuwux54QRrgbDiIBxzivzQi4j3x1S81DaYJLROhtImjhN57m2qQTp
UCDsbXTYaM/gIh71EaVbfGkXecwt11T/9jMDfTkjtITaoldDfGVeKj5lzDRi2W9/k3+skU2k+vxy
ndwiZMm4zusEDuhmyRhcMpONGcqI6CVIIUjhYbkAOXmwa02FCKfMmUGPYgnxPOOCo6xpRdITZ+kH
tQS51RpQ1VtHONUJjG4iORZRjJ/T0Aa+FhX6WJR73cpkzt4QpzCHqBHZdATLQlilTu60qxqNTnC6
TlgAut455iY/hfHqUnt0/ba2K+PUEpWF4I/zsnTAHZA7k4YHDn1bIQvwuK06UES6tJSw/LPA6Il4
QPJBufS9JqgUOENGHRK8okbY4CxmJ8LOA7I/9ziMTllAhP33zjiRktvjcBaGeBlMvjZsfYMx1u9u
ZBW491CYIYNB7SxYAzNoUIt8sJHglezb3JBIP3MyNqcSnCMgkpzDt1wYW6I6h1+dJlSr4037qR5n
lRIWpye/0f10NQtodZa0xwjombnud65r/FMMyoz7QdiMS6+cjbtKq3yr2OLot94cocKpBp1sZj3e
7aR5O5sr4t0ejvF5SHK3ec8Wm7jv9gUUkq001wMWlhgWRtiC/Sgy5Yspcflq+h4TxzawFhBWFh+R
6l2ufG8FFgQvbcukaqGkSZTw5IgerULxgYqmLwFSeooddPPfi97IBrX3I6bgI75vDRzfhEM2iYGm
n23PqTnMa/tjQ2w6BSQamvc5x2PZYFZq1cHuY/JhUfEcVDqiRuTsog/N+8sXpirQ/CL6Xm5y6aCE
2Q1g6fsZrjYN9f3IEjKIO+sg2Rx/c/W5O1DbPiAYbzrUKs5/fgmdNJv8jwxZw5SnmYYuyQGDlJGC
gvoFkvi9LnfRn1jW3HdFARVrf/hPgrJBng50i7DcQZkKyvtHgWGNmM/CwH7vJm5zsNiEn4JqwHP1
b4sDB842+xdkqXAl37Z+jYUAtjm2K7NMPhRDTMD5USbjffeeV9cmPuDYV90r81AA5mGc5an//Jxq
vx3D0wEQp0S5pBe/ZvcTILa0H0MpIm+BE3s9SMHFbErDn0hYhsaC718TFAMZxr14GrlW6UnQNXYs
ufPe4k0lpTH33ef/2o8adEes4ECKwTAQy4c5bQSZLkH7ndFLMGiI+NZiB5lmBNMolFSi2IpPkntd
7XB2IcWGgPuAqOuJboTVjvzBIdnO9ndkom3VtHtl1C3UCZk40Qqcu5Q0vA/1T0mWJh/hGvL2UB7F
A0isD5eEHFFTsj3ax7etuSGqMn0qJYEb0nK4PN00UY3Ke6FlNYixJZQibsWZbVBeO8LhsmEesi5V
lbjIyk+wpNsQGRLQP2vZYRkeX+wiU0OggaR2UbGoxeU6p+wIZJc2MD/Fmw2y7SkoziSIGHCS2y0d
Xww5RVWunzCYvSDpZXnO332zZoUuvg/EEYY+gbUf/F2aBZMSI0dnEBjHj//U31JiDCO3uoZ1aR92
oIbaAcDAdweBpN7DR/AsOTy9FBt2Nwne+fP73DxpG+hhM7jRY7Vx1CBxugFwdOadHe8Vf6AdlYKL
JBNEELLBXit8hMo1B9Q0UAxTiYlsMMxDl9sV5QKUNE1TiMLRGfX54+Im5dSGptZrNX1BEHgY7/Lv
cas9kTsYxvXOIVM2+DZFeDNNcttsh8p1EnnwSMirkm4e7dkHYW1ExmRaCmXfEIGHG5RBJNVjCt9u
Mb+dG/g9a9FKhfo903BCkW9urooTzUpaxpcn7pWw2tvDdh3aWlHt/uJysdYtDzeKBqY/3ViF8t8s
uAH0snkJGSoSfZMHb6gLX38LgXHIZb3XMOp70vHSzk08lYclwZPnplbYShnDkar9XEkCl45ikXAb
gYh+o5QScBtH/BM8GaPw3RH8qN0wktUq4HHTFjv8ch6AmF5DhMlHLXZnOAx7WgDUuDh47zc5ODcw
I/uIS0bkOX1JUD3PKDeHU9AtFL2JB7TBKsTk4wx/q2aDyBESgUPI3Pn74uLZpsdp3DsMQgDLqWz3
Cz5ncgYXWHowr5ZC7LeOSm3lrYzS+bfNYR9ZOTURbT7fVjU6J1oyaIuzskg9Zm+wwlUDz+Hu7I82
S79ZJKj0/TNEn4jbLwreqqPeMnnK4FJWea2gpP/ZHE7ODV/h/Zba+EYZ5XlIOKyf+QZJNrLq5Cvn
L18GU/uBaaXDblQ35Nq/rjokGo6Emrb1TB8/AVftwuXXPHf75n/L9RycNWGEBv+3sieeEesSXW8l
SH4uxJbmwvp1H2flOczXGdDdN4P+QSLLObYzSFIkYG048tdvo4mYoyVwz52ED3Ha3DOIhrh/aswp
UaTSIFWW0k1w3nKfiuraD7G0H+jonilolNScQ3NLErPywULFsCuSGmcI5NWG+FqO7Y3EXHxRsR21
02x8Macv20gQF9IDUUgaNNV0F8aIhQ13OtRTrXR4JVnjDQpX0gDqp6FORW0vxTnvOhe5Rx0y/YYp
4T8HqJw1hFkuDFYRoqULASUnEYD3x6YSwlTP8ulASidVKZhiuXL75XTumtZoltljaeUVRZEHTKKg
fkN4PRFTQzEQLLHBRrQrYoVwkdXia1ebXkRebbzCBrlXoQ31BcqNQvcD3vJPyfK3l9yIFy6hJnQG
uzlBJfnOtOf2NpPSzXA9VQXqKzlMZ1ehKUih6Cb4taLLkyVE1eiP3iLnrHOHmaytIfndrSax+Qvk
a+BB2Itx/OUsrggQa3yzE42wxrUfJLShiLMWcoJjbvzMhsOH5pOdJYAB7IX+1AIb5YYJ2+d4/BBD
qwOuLXS13pUvpOuAPt/0hAmii85xshNqN5Gmm+wGnaxgFzbFQevcmUR+3e+GTrzSWJqTIw1pQ7i4
uCJ7BnnwiRCcbjDtifBpTeU05DcA+hGT2VfSKZgewJC3EE7y2Hhh25AfmTwIL9Kgny9C7pRnhCL0
XrzMqSdYX33Mq+7eA/xtMK01Sc4iAq0cDfjc/q6Mle2AUdDgXisOsMTRQHsKfC/OBCzzWsJH+ZUi
lLC2+XCpb4thXasgLWzMzFfxl3+F9deDFgykHz5gMAANWOxE22BuiJY3pLE21re99QqsxIzHmMsH
q+J5TDIW0wgii5sbfHGUEfqUDFqQo+j1Tn1aJN3q04zP3mKefp/D+8rm4v5a/nmTWdMsO4I3IU8A
SVy3KK+STkM/gjt8ytO9YF8jpNBwa2+KHpjVHnQAX2qZtRCwE1r/3KCpi3EDmvQddpSGVHCWozqy
43FjOv2N8S3JIeH3nR+SCQK69jusoRMV94km9kvEQI8xOYnZJtAJZQDdf2boftO+Pmq0th4or5/1
KTC9abH/f2AzR3bO+H4rrVElnCoAYE9XUWW5QdOPaeQCFSQ6pltndluhGsPGYXqCdHv1Y+dhsTIN
ervnPx/o7g2DKxYjBdOFxhXUg4YWN3rx9HyY/Ct6+arqM+h08Bum+XTXhUIbWbm9afkzlBxT0uKB
K/o61/w5wGFG345jxcnVhCswfeUESpADndXdTvPD0QEVMWgJKT7fUy9BmPY7bEQD6FKdJPZm4+aj
wmZy7lwzJ9Ykvu5BT6aIliz2em45D6QmDUHxyw6RUpmoP52uudRhy2f595MRyuXcQKX2IXykXg9f
Wh7TKGJw37TBGH7beoRGLbaYZdSMMVCLzfFL107UOaajg3sPr2aUg4RxN4fq4sw7M9XdHgjBSU1X
lq+iOVhTZC+y3tPG8mUao7IEk5Xyvnhe9n0PfL1s5/F9onR7EqfyFCE0CeUetF4/wZGEtgUK0+Fu
achnxMELdEsIeJ82YgAIk/pQP8bPTcirhu6+611YTKRwPKu5uplLRScu4pNfVMjj7XmOXwvg67WW
zda3N9gMI37wbMnlJ0IjWlhy6WpnrbGmLrGY0qhq+SbAobIYLYE60Z+0bhiMqCtqnBRkE2/DTwGF
Qr/HuERAXgcYSM3hs/9iS8HpKBxyLUaQ0KEXubdLWuboign/NTgK1yaxzl46KuQhF4zvUlaPSrMs
cKszjVKj9cBa7X3s5H3rwbX89F72Qqrf90ppAJeTW1La5sKGNCCozApk0fwXUfMvsnZHMM1VPl/A
gc0zrOQ17wj5hToeOw0FWeQ0vR/w6S2m6NgogkrRLkPcY3SniXsHseNdjL7QnFroMbqqhuCX/CsN
8TYf+fHDSqGxslcqJCnf+jx4NJuNmRwDHh0tuko1gv4MEOh/TY8/e+Sfwbt9Nkwkyen54poxnhY5
zNQ3QCMJ7mhBqiYKCZo5aIn/TgCisDJdVxl3G4ww1LC91Y9sZCllJT3kQvbhgf+rPqMyafqUat0D
ahippaAjKk1wjDA5eJvqIzWdlsMsdPna8mPZwFqDiiIBBVFIdnPV06xFWebpZuqEetXGIH+v6ary
YV+D5TcIdAbzv8wjLP+xrci03/fAr506bOooR3qyx6Iua7tGt30Ypoml5Nwymp98Oa/MHW57+Ix4
owQQFtbeSy4gS8JoYWPcXiDmi+ctqMuiYu6hJgrl8Q+QKm89AKJXvOuKfbDWui5xPAyHjIN4Sze9
3L7CDU6r1Vx9kEMCgdxObmywxnERTWrj40hdHUmCjO9sJg7xT6IlwVsx0y5P/V5likVSfOIXapTR
24NwjEkq9JMYUmp64uyxnLS4cOu2goXCigI9Y7muLCzu/x6ix/WwhGNZbjKe5aYx/bcqmDCmijJp
Ch3PMfyMqCbWQOqDbRowWSYBfZDqqqtCbhtPqBnT0su3O6InmZfGaEXFRj1o8fC1YEfjfgZoOKpW
uQvSl3UApOwEo3RbQLI0+cC4VTjbwIW0baODco1DW6nxr7YnT7ueJO8n0TzBn9A6eqKZRmr7FsGl
QipAEE43wEhtlVEfRmqD+O67LmAmKJVSxIaOkuIBTHzoVEDljAZxGucXh6iyScuSxgYSKVPWCAC3
8MDbJUZDS6ikHRDyGDzrjM0+4uHf4EgAFBqfAw/Qy7A01H8H0JqmKG9DSaeneEwlAQTc8NHSAqJS
VTcU0MzH6Yop/KSMuus1nXmlAdfkx1Et37PzpUuMq2HyBu6RRzTmV84p8JpAtH3r2JWXEUgUKIPb
TF60HeymUtUgRJA3LqXB0pTuxewCMQFBsyT8sP1wNMPVGoCruMH4V2RgjZp7CjTdJvIF3muNHZda
3DYn8h0pzWdzGnX/4wN+oHM8OkUpS3JZrztSt1O4maH8zg6H4n/UOxEIloLzNtOcEpUo8XKRPEVF
cTvwAUdvGkUEEGlZFTBHsJrGQSM2jBEmmZnd2NHiITJwOkMa43ey8F9ttf7txjYRlD1nxBYh6siE
NE2mBugfH9MS17jd1dnqbL+Kpivc29U+GGP7GnZCVusuVzjsvWzAqUlLheGvszLut8d0YiKj1VQz
Md8XxvB5tBJJ0qzmZM2Nw1ujSOA/ATq8VOg2zieQl3TQYZT8BKsKS4VKWD1vYub1TtxWuwI+kzA3
hIkom4IvVHZYaQfM1tg/VUjWDgxtmaQwxQNNw6f8nW5S/irgqTvc0PnnskCO3YL7P2QgQy5BnE0T
ED1Gw3Q7cxyfQR8o7yCZyzCMaTlgmzqGI/rPHgdJLDGX8CJpxr3fRqMkZ0Ufp6ak7FDCN2EuoBGT
pqlef/77gMO0ILJ6GE372Q6zih4k2bFAVfaNNjGvoF1kKE997pvCsmv6vBecCRyuu3KkmfpKSOPK
t+DcqvIyY8YknvIC5DZ72xLH0ltQtf9srKdRet3xse3O3ZIrWIV/xaaaosByVcNqKT3A0brHDH+Y
3g2hCQRJMMDcyMSFRl9l3RXxZvEvlW2PbnpoYU3tqsu/2iiGwSnp6FSpseBKSbaMf8gQKmdq3D8d
OtnEG8GkARNhSC/CNtIgW9uALb9RaKgAl9kuUwPiNopbPGEpmWFymfZsI0Vhb5roXFIoVnUMHKZR
PVlSNoeWaCCGoOSjPVQUfe6oxV1lSTxyRSy1nLkFAPiBvWCB0MWo5jh+xC7v/gpFrnAbVMliu12R
blDNulhUdPhmMyjljZRNvBy7Rhl2beNhFcN1JJfYcOmYd5jsMVec7pjYGVkxEv9iUFKpmIYs/iAq
2z44EWQPCK6kmqTVAyw65oM7gngZ3ANl+PGBNM2LTm/r5B3XEaM0utKHajgpk/DLMpcIdl0A9KRF
3L0F8TGf567SsgyBOpmbtsfs4M9q4Sz7g0k2rNBB7/zJ9YR6Gx7D3mR4sLUGZWdVOLzb56OAjf9B
Bm3gDMddtMpKGGSsitVmXQbo+XffH3i/IgiE8STEtEhDGlFFYu+GmXWTPAByg7em2IPzA96XjRdf
APWI4nf+5wGDutVtWUmPVyXQR1gEbryTr9RjC1jby0fikwxB3Bw15Vmb4YHkIF9CTlULmH7eHXZH
OEdwEJINZMd3kvEnxhFPypTCMnZQqpaTrQIAUWkm+JIvrMd1/hCiSpSSjfeCKljyPGQbrO2Mx5Vo
QJzr2KPnEurSBrSHhjhWW8GNz6nQ3PmrKS75AseOKQzOYP5d2vRyyZLRFQbFRcJm+IhmfUt0puyL
xCZci8zyFPZjGGhH7tRsaLwIkZdFkFtwT3FJT+MN6XhnbgokmrVcyERiAsxpxauGNTLXkOVwU8o2
jNrJbO2X0OiGELNIRwpkTQqP560iqfZlM7RJqfz5X0cr0ZC+baSNJdT5td2I0B10kyS+BO+F6S7N
X/JDMj6WsBzEgJAq8xcblV9z2cbwmCbe/mMH4sTrs13X+aiRtAtXOYF7Qef125XkMJ5CzERHeTCQ
YuYz+BRGKMrgMKz5POncr/tsivmzeXyHU2S9v8y3PndmFEe07/Eiwxj5bLXeAXKkgJ2geAxUYVqW
+nLljOvDniVcWQK6ZTG0QtV+gbsAQ9H16QbnKfXJ8yME0AWKKM58jyKx6FJ8euxhyMqBQ+PQD4WL
6HvkLOyCUryMfVKxI6aba0q9pJ8EohrB+1nCxVC3vpppHpdYw3rLGG9XiEfbxTGg0FMWDYvlKvkV
h7598AKDJitz2L69Z8KtFOqDNiA6daNft/igjbJNCV/H30f+lrTGEbLyiHQ/bpMcLENpuBjSxUJ1
b1rjAz41Kc0rza2QiGC2G4E8+s1H2bBonDctJp5WaPSi/9VJ0TfSIA1mkRORbNeeETvFj4WH97wX
mQb+TaaA3hKa3VwcrPxzXKr+CB6bM3+lPZeRPFfI1VNOnfjiF1HUWGq14jozSE0bB1jDEVV0XeXt
ZYcvRQIotSEKRltOqEtulaYHZAFz53afo2wNFTtl4x7gkONq6P/RJ2ed8yOZQXIO7BDGnJ+tVgqT
Q40Pw6E7VS7bKa6l/FdGSzKhFF4kVNEGlkmaTfN0gf8aid1KwsBm1PTg8Vj8HJpFdZVEN9mJ35jm
cCy76aCAkFQG7KZGgh7Iocsj6wWL49/iNQQKJL+KwgpAJxwthEJpLdqRIiGD5aDfnWZFg9mLh3lg
vZm9FXPJRxfJImpyVVliSft18zSCmOLnt0QR1cRXMErZIRVNwAYofT5nyaHtwPCl8LDS/NcNw1iW
2nwgb1Uk7n6WmgjV+HvfENeXaoPjVA4ORMAHBn5VcChXt5zUF7lOQRKzDPowh32lPpmJ5RKeQYDp
eJbkkk0be61WMAXFU3h2pgy2VYNUUqCwACe8iB2ppBjw/MgndXX/N2E00DVG2T7fzzvhnwYpnrX+
E6BkF/aCeDTERqsrydOshApPCPDzAr/Pg4drR7Isosl7BCyt7DJWLB+srmQwXzVZXBv3f0nEEJ/S
fdMUbaIUsGiDy8krFJaqacR3NxPncKJcxkB0hNeMzMxhn5KdcIClD92GPUrxvgmfywI2LB+hP6/p
7Js+GEShY6O97b2staMpe9Be0JQTwD4eueYqNDPS5idMg+jQ+2i3e10RtBRt8qNrHsng8W4TTHkx
uOU0PVI+ZjKOfYlux41q+wdRkUUMGprx7AsyS8zrCb7YnxerXU94j8AFfLB7io+SxVk1rZQqYSBU
QIj6IgfFGFvsN7tDr36XavWrgmFdmUDgud3C+rgQe3GWzl1xGrSRQFnZtnlCoZYjoKe+IDJaOrAT
CPZJMqGZqMaE8nlPR3aMgxTugb1Sqde919jM4psYn3CVRZWhhaKIP2C84c47D21PaVMT7fdM1xoF
nGkK8wEnZGXiNEkTS7Q31JfhgFv2EJsTxtduyZ5urS5noe/L8ty12ybClB6dL+AE3wxxsU576qGr
6v3RkDBtwSbDE/3KdX4/+IG9bNGraA8XAxqPYTeo4TeJ5Iq+sJ0O+/VLcrHD6FK1eaJgkEbCHfR9
Yv0EjgV9qobrZwVkU+GFO54pSNgjcIJqLpm3nf4E9yDSL8AJbl8zbhazx9kOWMx0ee+tYFHB7Hg6
7v8VlYb/Q1Zgd2GmUg/tYvw4bOktpAYAG24PFmqCUDAPwm6FANJk2hPp63q28TqUtk1MFwz5+z3Y
R6Mye71su9plwa8p1jM97A98sr0q1ttZ8SDbjPJncHOF9XeP2AdCw9EIz8Uk0WSC3dygt2w7+oAM
DelGBJpiORssfriV4E7YV8t/RwhAm48GCZs3LFC2e0SUpuAdXswUmB0kr7G8FqQUoK1dB1zp2XtK
jq8WIOZFYzx6ZnFoctGVVkH2bNRJo0oKChe9njWtLan4lCa+29UMwT64lDGn2OZLVTlpJVGYUN3w
aZMVip/6InQ/8kiH8yrLRIdBaa0yqix4O9I0UNRnaW4UZ+gAXUbtCtBfL/CCQvFQpMsiAuPfZnJ4
VNf0+42I2npD/wjSVFBycHRGKPxLSwXA7wO8x9TizLzIUZ72VMAA2SVaYeUwLIZIpWQYoz+2Ao7r
1GNQk+rogau0b4foOMHQMrSolqG0jEsIDzvJqK6+OMHMvQhgVYI9Yu81kyN3cQaD7/NR95wm54Im
afjZi0wAU+K48dILi/elXTNqsGEFDPUedEq6NNtiyEnYCmt+cyknPhmo/wgyfCyuuDeRll9qhe74
cWhbuB1WLgE/P5bbD/qsz0W8u2aTTYGUi5OEqRzHfql23M3u3+hOufY3YT9k/5nJwmQH5jC6sFGg
fm6GXa1JF8AoY9aK1aDO5PJsjJ3ekwdTetcaFatUQgftEyhz5z1Dtf6Fz1QtcX9kQQjY8DWxVEBv
L2C32Fbq6rH38pW3cFj1t5kWL86dN2Hd+AmHCuZwBrHwt60W/IJQTM78tk7HjZ6mhTDZImqCnb1G
MgxeCI6rH4XZ82u9Ora8+8PQ7ZTw1zNGWKnyexpMlXCvaHJPr4K7wx1KLLVTXjpZ8Dpr864+Y4k1
zYbZMOoRmjwMtN6hOCJ7dXC7Oavy/o7T2gYIgDmYCxhSdh7VBbj1Lr/pIZT/8cUGbCgCql/y3n1U
53ZzMZPvbeTuORxw1qzNT1obdsfhC3EdpyetaZalanEYVjQ50HhYYxUdnz0/S32PwR1yRAA5av7E
yoKW7+zhipkW/erokEwrVVXYPjwN3zCRMC092HEign1l1Ble1qTRZaMLPFVdoAgDbWKYrIuDsFQD
BkppvTvHuhZLCuV3mANPQSI2fPQHHKvc4aK7yyhjR3VIR/8y8YJRgJbZ9yujn8C7huBI6hKM+97Y
V3VWGmqonyDrpyucdxnBQV43tKRtx9FHhp1kC+IOPVANk+EiYR7QSqZwGB6BfQHSolvh3v6zeKEc
6eTN2yKc5WjKZRIXjlBptUAZjuFJrouOmm5FAfMcHjGtu2471Gl6zRuqvgUsiTb2A0iGGHJm5yPa
ddWE6sxovo9b6CWTHPGhyS0/y+MEy85DtsVO1vz1FSevOvzfOUGeVx4jq1QafwfqBXml/HTgUpYn
xOr5stP1pXK4nE9/WeFGqmXcwmcRcFKM5ziJksJh5tT7RQMWzxTvDdHVELJ8JygpvA+QrHfs4q7b
INQyjRuNj3u8cYnJM84MXmS2CkBSsYT3KIpzmywIQhnhJts34JzJRY3iBXxFyJV/Ee3YYz9tCGfo
9cOjPTlQuCG9fQefextK/ryzN+H/sc5dFqFi9yYRxi/+5q0sKoujx8pCDRaP42e92qb2mialUQGH
ir/Zlx/Y4CSX1WSn13a/4rZkmm9ZZKeXVO3MW3I1XWvkCdvXaxNhKe2hqyP3Guf2WpeaMB4enb/4
Rgc7GyBMp8CCBw23QMqvyD4RZGOf4JNK0xM/b7XBLo01CtEUXsnHeXmqhItq6Xvp6+TakBsp19x7
/0PT6voTHlXV4Cb1SJfWxdiXDEhk9c3Ik/uC+ST0T9+b7sInOb/BK+GQpm439RQOw3+I57Y0L6Mc
dU9nsrwaUZ9wdQ+MnJUynRXRiG/weoSCBLinS7+yv3LVF6kkJEojQoZUZDDkCyGZNfipVTnEGoZi
6eeat6TnYf86RGbQyksAcisjb9/3NA+gX+oz0J89dKgjdH4knWyEGiYgCWNKp/zfrmI0sR5Nmgsa
sq6FsOUis+r3mf3y0jzUAPpEX205jADM8+poe4xmk/e2AqzbLrDs3wR7o1sDyYX9eV8IHQbUSZzK
Nyet6bDyYCps8mZ4V8T+DGL6KjUE/hfppbuvxkeSP7P3ngYFvurkx4/bb62QocHih7haj2DSe2iM
OLJ+QYNt92zqavAjqjPsCat4Pb2bMxCGraxhoRMK2Nwf/e3G0qFW6mnikErlK9bOuiF84EL/1X7U
0sZ0NBHF//c5BhUQDWu2iU4eve1eWHsTP7WyP82aAboK3WL+VwOaalmFVuodOmllwUemOvxsFOe/
eYRMeRHsUFnLDnpjigwVoI0sNPKlrFk4JDqhb96SdcrC91TQI4WG+vYaCIzpiBZIj8jMJWBADRy6
Jk7S/6+SlOqNO+xV2rxKrrcr0Avw+8/vXXlsBcC0WFCTjn6zDF92X2ByzW7ZylI8cc7tE4FWwMJx
ncQBGj3IOts54+Gc2aj+9mrI8xLlBlHrX+79XmImVfVGj0mYIxGa4XcvXSJx4MBiLc7yc5rf07Rn
nVeYajAsUfjKDoT489aQwM3Z710A5bn4FNeV/H26ipPov4EHQlDH7JlFPdS2/WtLA2SnxdKItlmR
PJNKprzgpjVTF+/vVWs3wQ1W6/Uv3VNyh15+BQuZ7dUNfLpXy58WE2GYwW5K9CjdflRI6at4P+Yp
ukYf3fLTOLu2BZ0e0KKNbVm4iJaVP4SwMbPy2VHm0g0qrvYSpOTV0LVm0wtDcsXsVU+At5hk85ia
+G3gDxiTI9C5gp75LMEecbac/8wORI20MbbmaCZoRKOG5MLbNtCNEHekA3KgPgtxFOKpk5Iq9/Z4
23Gkp/Pgd/DoJW+sCF+A/OzdppDJ4/UuuSZTmAJfy3IY8vpqMCWOXSoFJ4ozWPd7DRo3+8ns1HoV
dnydCLHFe3HHZp/DCUUb1FlpJnuXPXlWAsDglFsL/gvOpqQGD87Iq0WWMAlU1QFxokukLAfJcu0g
9TxXWrUu+9C2Epogr8rTmTSzq4+FkhDzEmQH0wk7rzPpT1S4JF9LHRhzSX7YnXx6sCHWbFrSUUWv
XJMl4csHe5p1+G6k4Cmagfv4OZw49oBYC1dJrs5t98X6OZsIpfQo2bZHus8JbGNFC/MDkrjgDcfF
+LTi4Z3mv1UpXproIVEoVXHB4Uo/Mrc7TOsZqThAwuxwMCCOuyOC3ROKtUPBvEXEOYNqihkdAONw
9N+hcBDxMqtuS0Fx6WtVRWq6zLkzL8Nn4QT9Utf3Edcge6SQILmFhjXR6YY04vFARG+auLvyoHpV
VFQ4qRwYelej12UtK0df9qLCeL0D3xZAllaTx/gE/6e/S/H3d68C312FzC5AMLZx/NXoVzB/51rx
gpKtgjfpdtTHbVOP+rzAWtHVovEoz+4o1e0d61f3I/ZbSrTMa4BHHazkYvj0+2es9sHmJI7DTYHm
lR7wmux3R+4XQ5DUxSZ/1NwaBi0AnieqSzAoOx7RU1PY6v7aQx1mZXZZN2yJ/K7k5dg8otpIk25v
KQPshqP3u7K6dAHL+eLxnch3miqMWsmGMMvX+y+b4n0NCqSGUXtkUEzifF6Og41gBw87NOLtm6Ea
XGXwKeVvTiPAKKFkd/BJEtg7fj0Y+OhACjjwfZSYMCo52tu7J5HA+8gnSc+9Gh/bS2JfLFFXYNhg
v2NTBVRWQKbLSUTrHmN9EeVj06StKrOy7YMU+kAls5FbGuhUNwWD3MmAQ7seqLu9bDq2VBX36tmq
GnOldi6pf2WiBEMgot8GNOSLgfWexMPe4kO+MXNrvnUKvsGcNTnKtZy15LzUlAvMSuGxxmtQoaEt
7RjzYX2V68ICV9+ZqKWZRj+RcNPVd9hdohSKKEkCp4O7E+UknZoQ+eBQWyMGSnIj6WvMHN3nOg+V
MzASUuK22XlSXl263B+tdlwGv4lHl3DMkd/oBNL8LkSHyGu8A3uene5RP5ettmoAWGaOHe0gSzKl
z7MEff3VeZQu6pk4dT2L2kLlIpagjRuWEyMASCTxDux9E3w4U7Z4t0iVtyF3P7b4KxKxpMJBqL8l
zzLvFzs4GVkYlby+TWF3snEOfIyDgzjPTJa6QphpbTDPfy64kv4JkgqhODLMhbgHjXJ5li67ec5F
bE8sGUSu8Mn3BlvJ8tHcsHQ7bzlBUtfB8G9rKfliTgSLB+FBA2IfOjnLy5a/vTrRkzR5i2WLFAn+
UdWcmZIk2ecRMiqyKOlJ9LwBaEiqxIm+uCnrX4DoiBG9sJJzbKlBlgSgyp47dptyAL4KgIQM1WSD
oN6squw2GOrMwYRhSc4b8zMwhJ2+40PwH7mHQVuItRs7FKYvTlKYXD2QzwJyT/qXUcCgbYUEO8Dq
H50dCN0ODH3fZ8+cC44cLs9KC6J8NjXgLVcjKrENcYm/hrLz4Pd3fl4gU+ppbx4al1BFA/X6JNqC
8+snWHZPV1BQeLa3A/9TkUPI1hBTXE45xKetDgBNSJuEJJbsSbqjW6Yx7iXpuJq7tMamKjeUamDC
O1jDl9j6KyqT8hAPsdqRyjXzhhRmU6ttRebbxP/0hmS6QzsLSqNX4zZTwcSJnRxpM30jMOcVjN36
EVk45ZHMvaV12yU57XhpcnU+VxJ8m78/HzcMijt1HT0HXZ6RgjfD1qvJUKuatKYmbepwulMsg4Ma
jjP2ZAOPGOW/bspHbOylqbN4TTlx/IY2OCl9iXWeYM3TelwGg97garTRfwLNs2sQVn5RUXsl0S3Q
RsAZkUFCUNQ9Et1DC3PS41M32HKszRdFEC9yGi64t8fy8OgMi2tG3RE2lavXPz92VxtUwF7m8grT
6QVhs3qPEYPyY4YtLs/atKeJjudZs5IxIkd74nctb+hAzf7oI/d24ms5xXmqjHqTIy6N4wytEJO2
MRb3hQ8YSqfAp8EGRQBZNqOg8Ob1zeC8TB1pNxWi6Osv8G5C7+vh2JaGc85LtYQ+0EZukFk4up8X
V8dBGbZlEHeI0wVM92RfrFwb4BxEfTpBIK/F53OVjLndyJWKYxC3am3dfukflkPeI+ZZioUO8WaJ
IvDE+c+OAsW4b//xCgfJ/bSP1/dlM5Xyv2CwKUblt9vzaj7zJ9EkRyHZQt4YC05FMM6kcbQqRQ37
QP35ZG+fBEXumq5vMWxwjHCQa5s4P0DtxizxsgvxsNjyBWvddSDHq0Bp4P25uQE2UiEgt4d6nA5U
Xrp9c4R0Mq8dZwoJSGw9TLmOZWSI+NtfCeWPkrhxVy1iEaBL2GSSQKS9mP5caip6+9+ku2K/6U5N
0wD7B3Ezb2xVbDdhlbOPz9ptIaItX4+7TeScJd01yhHYpuQHNzlk2p+9ZhDWYRp7g10ct52UDJ70
oPf7pkg0wdXfnOsaPmOkbCvx3divn4zmJiQydtSemIKmo2fnnhYSXhPtDImuJJSkF4/2BoLY2+tD
DFhHGX4xnvaz0p2t8cWaTxEDGWgvSwDqhNGKcsmGLWULr29L++8nR044WJqra8lPEARjXluTpdDA
n87xZLjHWjvfKWFcG7e4djL60u6+FLqnIC8K8jdQB1f5u9W9sIZ2rezwrwf2VdY5RIpxj3f06e7H
xXeXO1xKioZYCwn+3cZ3I0DcNYJYkzOsbnEO1Oam3siz9lsvPZbGKWFUId6pFeFw0bd3z94TwhX0
S8+SlhzuUNLEgjbiZV4AK6ZSnrnMwKNrOY+k2LoNTgm4EohdWy4MeIJkzEHczGMPRCTPhIUEw/rG
ln1CKgUYLIjxyDoFVBgwXpA4eyuedhpsherWQmR0h3n/6VW3CONBVmZuurwN8DgUuJJ7+6zFGJ1T
vA5BKweHxsloyURkPX5Tz1jsQxti+jEiUY0xNskDpG8/P44ZbHpqYCb3HOnJ5fnEk9WQ2oCHeekf
uFcqNVHoOPFB3cSXsG1AIR2JGc2vua9nKgpS/JGiuKyitPP5YRqNVw5xtDO6rdp5MdQItFLs3OnX
Qh/3zv4S9iH7sVg8GZDZcy/HKOqb7ta8Aa0ZfNV/3wbLcf/ujSMoytE+tE4YJvWQqv+pCtkEmEWL
MsKlhgCaPn9K/+aUnS3f+JNZlB5/4N6AvD9h5jUXfn0MOVO++SIu0KTq8eY6eSISmOVx+bkO1QTJ
gqs+vo8DUUpGuszZ0kJ+7Y8xTDbvaJ7wBHMU4o5sNgbKyaIT8RwMaQOSrVkgLYrinv21BAH3WEof
U907wx8FZLKtl3ObK00ombhuS+zhSYIpHgBmS7wzp/3Q6Q9242hX0NY/J22gAzpjGjm2tXmYEmzy
weOvgxijylhgX6vYcQjHx9AHy2hzFHdmLCjznR+8a1yyBeGwNEadoZypcX5fm4milyvxG97yAOSx
lMK7rJyEBJnIINwxMT4s+ftHMaRGbhqLJCJTVE0bb6cQehASOR100dqNf8upD/6vLC4Z1qwUax0z
I+UQwAmvVU8098ht+1d0Uhfe6dSFX3XXCFtoLZ6DERKAP/x6RW8TD7h7VT3IP3uoNpPjvnglMfFn
g/Vj8Tn3PDgKdGdVvzg26KiaQcUHYbEPA+lRSdbcDoq76t7HR3rjvxbzZcLS5kYDESLcv0oQY5N5
URjvhsMmnPLp99inMn5++CUXhmd2AUVmF2A2Kc4RIA5A5WytXVcDuBdZT40/sm8uM12shQWobDeG
BhcBFljl8y8eWPjYbOxdjrpidr+eKEB+R0OFkbjG/DgTi1PGE5BcT9Hyh1v/pcotFfG/ZbJhZJnV
XcG6cQ2yXboFngncyInWW77yae0b68yy6HOX8V5sLk4n3ksPpO86J2bN/7FzTS96ajZRRouRNTK9
XTzutQEAQTAv1djIVwOhgL4lgcSNn8AtCucBXHDuMggKpe162eO1qrm3VWK0F+AKG7jluwIdhaNr
A77aVTvXrTE9x6xsWUu8q1KHmNm7GvnwYMRm2KqY1UoxpvTceLXozDSLJP3EaRrChr5rBa28aXZC
s+wfWFB2fhdONjPbVR8Ja6N49IXpLq7x9UuYcycPQRUmT5aCliRhmZlAcsBB361qg25Wv3K/dCwF
yQk56skkQSgHm6azSw5KJNXRa9N+jp41nSSTFxtthdmSOST4WZrpT5Za9l1fT07yKvDJjIshLpns
K+6NSCUcxoBUbmqWE1ZDEuhQdnJF0C7yBfwty7hKpTUi537HLoS7tbtLvUq6wdtI+ihJI060Rnuo
CV5TZIO+teXZQe8q4hvUtJMqtcEJYdjodxJbMYv0W4hRM0KldloZ23FKzJkMmelFLyAXv/kh+bws
LJnUp7esV/cZPgqsklhC1mkStTdM90xIR/MP5edJ4bq3uOSgKzltyjU9IsseE/6TEECWf6yIIHcv
LHMHAzrCfGL4XHnIkq8CdzvhwuO+B3x8Oq8xk3b0miJtdUJkmUSzS1eY8q1q4B/SD90o/FduO6Xh
zDxoN6PXIOKCl9yZA8pXDiwbOOmce2u9POppVOB5tW15/OE9mSty/KALW2lidGOFHzpUZJ7VYbbw
5XxwXa8kiVVWmi1fEp+KRwJXa+Gbw7sHAF6IZBrh6zuXlceI8MvvCCEqwWq9reOuW2nS2NGlEORq
+RbJTnL1UjyjnkhCx0CpB+7T8WjTvEuMAHo7MlR1RAI5CuGgSlETXii90lCAEyE3ISiUV2p5z0wQ
Y0PDBqs0uSwoutZNkzqrHgpSZBM/DpCyU182tQLU6GRy8s0XUveEYlLyKfRy3/+8x98y6F0CFdvz
GysfXSprYXbFmzXypCiVVRII39vzAjYs6VDk5X0yu2OhxulMyQHP9Dw1wnXBWrGB8DAd8ce36MQb
UkuHPDFGR2kwZvnpKQPx54+GVVZ8q454KELqL5NJJ8ISAMwHeIUE1VFRCfQ+p11SoSHdd++rSsGF
QJ0DTIDixRtbov5sT9jZ+j09YhC1Dx928Ywc47S4vAlBZ/a6b8J2jNd74Vl1Nk4pKD1yoBHTFUPO
9Qp0RjlL0Uje6df2rUQ6H9m7hSnN2lllblX7KudQHx7sWQzqPz8bFjC2Gl+UI9aIIreMPV5Besj4
AGT/xN7d2emKWz8zi7TnvqSW4QpQftBkapuwmq4sHtUQWTOmjEx1niMX/t97Yqw4NcKfu+C49QQM
S8vl3e4bgbmxWIyzgUX37OKdBOo7xLc0/Wp177RIBja/KSA1Ri+2Jqh594ZUYv64ZNQRow1WWnPo
dJdp9hZ2L3i+5zG5opXbYK8cTqP3+vjodWSLreABRQLNrmXORf5o9z02ji/mHazI8L3HPfyrsRdy
+csgmyfRgLOlN2swP2MeyKXe27A5uLn6Zo6XjEKeV6cNuSj610m/8+ooCyfuy6076UU5oopVFQE8
wBOo7sIRFFYCBY8UYUxsiAdOgJ+H3OQoC6fcmbuAh/SWDI+fM4HpgvuqcRiiI+XeoFazP2+0EBS0
M5RgF/lDBe3sgKyRXP1fC8KBqHZ/3q+BgHSPPU7Ng6iR7zqHtlZsvrldP+ivRX6LNIVzbOPfMrk1
4veCeWgPb3DsIojrdC16myBdnvqRwwbbIDfKHVJ8n4sz3QT1isL1of9CJN5cY3UY9oHUa/ecBvGV
PL3yqCrlnNSaDNmbOygH3M/R65Fdwxn0Im0vcU9VSQLO6FNmzAT1mtcva37UdBessPwFP6y+dtfC
SJdW+w1IMnrIFFhugqetnXL86W0Vme6wSx0apFY809pg2ms+t87ZdhZXvV/4yMlE/RMozqPOyOua
d0Z5WUOyAvuFBghmpJkIsmWkuZMXOrklJ57wfKcl6TXjEv58czlaI4IUuChFH4y4l/xjo2KqakAZ
T5jUSuJtHU/CvFnIZ0d3Rz17XRzyina3n/tB2SSeo4AtX2SXicGdWz8YqTa37S3c/9m6BXz2mPk3
JTyWoDnN6bjg5Vwc6ny2xhHhcbODgfKLRfUc4nw7ORB3+Z6gL6kqfHsKGCklqWm8VUWQqqDG/58z
A2p7Op0iaMEwkBHrsueeW6sC3ZYmIuZdTXvVGpi8vucjcUQ3cEw85QTQQJ6+dKQd91mdxz+A5wwE
Iu5ec/d7BVvxuSHpfBgfLPNFYWS69GGo+vS83GhySwIRT7AqiJq0JCA4+Wa+M1uOwBPEW0jPAtFP
+oGfDgGiT4WCJao4iexhv6xc4hjlSbCXoe7LAdb+M6dBouUa+6/Nxw7SJ30OU1Psv8B7Nw4PP841
MgAgrm7x41h+JnuxYfx79XceE2fD0eYu/euRrGggumGdTmgKXwYM/2wM51mqbyBDSpJEApy9SKa/
QdA2grFO+wp70Rp7lv6IzFn2T1T2DXk9HDfE65fmlMYCWdqy4h1sq5t8+MMHTjicPJRRCd6x/T6l
QPKotUrzQheCpC5wNGCjZEWb4sMWyV7ZDba7OcVbt600v/E6Xk2gUxyz6uQeSh3rIFZNa9o5dmaB
1qDAm9Klo16zkJakzfGa2CkC2M5SyJTMQ4lE6m3JT2NXuz8Ykr7uJmLAzCc6Y8g4nS1N2WrLnnUg
+2SyzXYkJowDUzGC1eVug1clsHTZgdewkf1wStczVxwMk2/AWnv3BPnDqLdPJDOC65gP8qdTkLRC
bRx6ruTXqMzSuPWjIpCl+omX+0Cci9uhP/Q2Lq9wcAf2gm6HkK36VG4jYB8DHIq/cMhmfSeH92Pa
zJF1SjNucF4o2SfV4F2LaWNGruubo8vbj1Hj9ZdGUb/AH0CloCsWVKdA/wBC6XqZJ2rEmewmmaAI
N4bl/gWYPtWiGonszuAOTNkZ0e4DvLSPk+AgHMNqcPMViQ5xp/BQM+GshVzLPetXwO5Fq38PNUql
2CIyIyZgmRNN/yfKPKZIvYAMWQnYu1EL4irw4b3k6PTSNDCTV2SpceQIyoU8CkYVD2PSwLna8o6V
njRLOa56OFDoMnWIe+hxEbKp1D0bW1uDOD8DqS+9XkpM+J0CTsXisIMYTSoHWxoIZAVEXaIZ8V0o
+YxEnlNC4IdGarv8yC+KpBsoQpbQtPHIrlkb/aiFTxF1mspmTWdmgIk3tCLmrYPNV+2uhbl9FXoC
OzOCLYpyA1r5GaDomOy3YahKBigJqLNrE5+VIfEZ8GkOsOE/+9/u8zvy2xRAw+a0fJDHa2jJQsO/
lYtgV+sfH67sAcyA+K5MlFINuD8wPsOIEvUDG2CKxYVA+UkofZAtzdvU+pyhkao7AKharwJFa+Eq
YefpPBPMlQEd2qGcnzahsjTppjqjsDtkpPUB93FhEpZYoohrxS1x+r/DLyYWq/wCSD8fgJPyBHT8
YLY6Dtp0hKmulv39exAGMQ9batErcBGeEPuyz68QSnv+tvn0RBhtrTIovbjsPmBIefnQ3JIy9eyg
49ASNCAcPggYevcGDpiuMjNnRZaeRMSvfz39tNv8CJqg6nHPg85/8Ib7Rl66KhTDkCho8Gt7b62k
FxVLR+y0FtDOtdLzU//T7tGiH5bwfdWGtgB25Z+6wyb+qM1WZ/dszJ5ki2/w6siatRR0aKM13nYR
3E42eJcgt+3TBTKhAOZDRwCu6Bqr/Ap2e6cTob+TUy9t85mmY+4hEB1cz/zHu1iib6rXf2JsA6n2
60WRz4GTsF7dQGa2ragglR5ZSk1SNkCu/3Z95ac898RMKcc0Z+jKgPojIRAwAV44LRXUhHDUH0aT
RKUUBDhowAoiAjfdWpL/Ya1PReV4pThE9zSF7HxtksUUgvLbUaHDn1EN0k7CqYDLO/+UqCoT+u/i
O2g+hr+iYviKHrD6SxILBJbd5YH49dcaqr76ubx3LG8RfL6d6YAQ7lJ1QbHTVHz66sbfisvdZXt/
b/fjDVMIzQhT3eaYJViIOWvThS9Iiga70ZG5sOiv5dP0aLoIMy20Hogt0bDpyryKWIaakZxACfL2
lfr6VRZ7pGOzYOQYfYqw7faRDYTyMhiSiaIsZR5oOJd81FmGq1zgWuaath5ljNJiB+gu8uF8DHZc
nLTW8URKqd7NN35CuP07cFONEci1ArG96BdM2hRYT4iuquenGfTuzGqQzHjIAJiuzAnjWeVIyM7C
xSt06kGL0tJRsnwy5k4pCwMDmt8D5jhsk3PDjdKO5tSQ4PftObR+s5vGmSpkVsB6CJH3/7D0lC0x
mLIkicqF23577xEM84pkfHvSk94YRnAlAZXKF5XCmJIeLHcCuj1P/4Pgoyj0jThqnwx6Ni2wqe8l
75qahTleglEYndovM8aN1OUr6lNxpOQkrWUGgSXtZmrZf3H4TYnwzGJLXuwwjlnHfPJkHYC7nkMF
GE/D2kAF2plPuWW3grgKlMDiDC3mYAA/tYTIO7RXncSTBCzKLDH5bGvchZyDh083txYf8W8v9o6n
wGs2koRevyg8/lkZW8WiyfWZzlB1t6y1g+Ay/yYjh7YYa6l6igBDkcFnHlDt9AU25mYGkiEJzkmg
uhA5U1MrZH0u4TZv81w60AKkQP2QYBJL5dlbV9envCanc38396y+YSby1QmZb9QTpqpOOGL4E0+V
AuBSv8f3cPjOyBpd4bxcttzHsyOBS17bYEYqFqUuXJ2UiJssH/0O2S5NMGFEiuSUOL8+rr5JuClS
Jfoqfqy2PLcFDRKRdGMfSFo8NWP2Oq3k5VxLoVfSXT1g2br0gz5+ZeGulQ743uV4h+Otk4cyH5GO
CUko/aUKaUE/U1gvfei5YQ8BihVHZZAGS4YqlcPyHiW1jHE5P7dhNYsjoBuGQUWwq55dh+tn7MQl
uMO6AXV2fSMcQa/R5AiGbWT5dzniWlQNrs2e3lZPbWxivhtWGbpApsOHV4is35L7L5vr17cYxNTy
HxyJMjeA4P9Bu0J9PyHSmdFgjIGz01naVStWNzo8hT9kSRFcUMt1QPa+XOJ1OhSaaUzulpPpoznM
CLJMqcblCRnbaeEEq8biZE8DsQKfpDse2ggzm0D6zoVENafQQH8+/OtAF3SPl18E3HJ9vODoV8J2
XShKsNKC3GQBKNMLtcH62KbIeyXVdnRMsc3VdMvi/zWVpnPikHB29yv/brX8CD1znxLQqTDKR4eK
xs1S6fvoatDtZNpFxQv6Ma7y6Bo+Zs0GZNqLslBhqSp1w9XcuBJPO5BD1UC997r7zBHEKzIoHKLC
gBZXGDOai9g8Wj/O7GJTcKuEP3cGWQB648BTBXBiBLcoEtapPeFRk42NETp0oEZJ5P/wmc67qrpp
xaUbrXM3ZFkVkIq9tmo6ByAT3vQX1EHMKesuIofpZML2xnNPHmHvxWalEBIzYbksgUroK0KtRIre
MR2j5ExHs5R+/5ilCxW+we2LBcBo3gYhlV46dNsiFc9DOJr6bwGeQiEg1UfYHTUmlZ6ax2uFUHaz
qoxTgQvSE+EUhiVqvrpuuuPiS5Y0TNHbukBDWiKX8pWWXOiRR9Nh+LFo6lP/NqDhpscYyrYjzwzN
Q9BwkTXrf1vvwDwLfmJxb4J34fj+At6BxrhGtRTMypOMATNKMA4QcKCijqWbBfgkd2zLMa88EYk1
rnZ9LafUdns+KJyDDgXJyFijSWIoiEqK28QYPFqtYhLJDou4C70Cy0fasc/i98IZhxiuqEN7N6Ku
OB0d1gBDSLWYKWZQWzEjdqTKaAITK9dglYC2yMFy2zC2nFd/TgD0St3w9DvGGwFXcaGgKsB57GrU
cMagSvbu1y6cRC9bhFQ/d+4RiqJGvtRK7erYNflP/8uqHrnVeKXoPC75sajANawAFn8nrHpSM2GK
H04PYOQGx73RhXZhvOsMGoeAXOyazMcoLpWUUc/OkM6kQhG6i7hmnztcKMMydTTJdSB9e7Y2VzPo
lMtNg6rvruYVNfsddv3Gg2zfZshSIQdrKKPT8zdo9hgsdEPbaUkFQUOzXhF+RBYHsd3kgrRAoDTv
0qtQYE0GyyvDVnkPmbtL2vx9y88XkgA9kNw7ZWXN4wl9ru5ioxaTg+iwJxg7/l26gGBUyZPN6iF2
/G3vMbN9tgOpNx25bo8bkCvVzcqWTL8YgFbjVTPfmropXzZRdtmVYeMDkArxky0Uk0dKP2BHou3f
vBfB3vKI+z62xga8j3UHkHrLk1BlnYURWSrFqdhC3b5T2co1E4MeqB4uqx7ZPAFIMNPlEmsZAkA+
2DP7oKTp6P0A4Ue7b3dxCb+6rPn+PEhqcr0O/2oK5RvAZe66NbUbV8vRStNTl6yUmMMxhJ2M4QPk
p/kXJ9kef17JEHpknZy2QOXwdd3BOtXd7J8CwjOEM2+S3GTNv8tOlNjvx9WZzjTnKJi65KyTONt1
iWuIrkZ7UB3+IaKy9y1+lv2/W6gyb8mge/cAe8HvSj3cpe5+Ni8AsSBztOOi1jjXtAgHbsGtJF51
Lsyic4QaSZC24eyyJEydtV40eP1cGvbf9BW7eulrnX4k7QtQnorzhMZWwgJh4UkmxgUAcuiI9Ork
BYqF3UpHwl2OEO+IhbkwbWJQbpoN8MrGXgoUdaHCOXIupIPgsgtRPDItA3PmJjaTUQqHPjp9IWNR
Oz6Rlw9su2rJgrgVXz8xYQ9NnhTOs64pYxTFv9aZcU4UbeNnRlhArptJrQbFQaU/8K646jYxI3mS
oX5v25WRI2r8aQgSuhum/3lNERf7uY3uh2KpGYed/m/6T3dghorCiOgqySgOs7DgxrSPgIX8DAik
+eKcAqxd2nvpAeiwG0ghkYXDgv/6zu2qOZaY7+gmaOCsGk9OpwchMInVD9hJUCP3jQkYQynREJIH
UX7YsqtOZ94zflu03c/B91tFIT5cTuWX4qcGeAFAAtaXQfpNXF/vuuyzOOlkz+GXmAp0iYLkH6eR
EJlYBnrnJxSbuozNrlds3VCY25Hg1+1rOWB7iMqwkwGu8JiS/+cYJ6JKhvc2uCy1Hf88MYHvROu4
v/G3HdM5Cel0ikckSOUUgIM41aqXXOY3PR4bS3vVaZeDpQvibGdDYo4MIarvxpP4MxjdxS7/xLSM
/ZVZVemJlCMA/xsriORuyrTfQrhIVRhIVJNf0HfAcON93NlGgmBGLdZkQ87QogJ28RaqIigChaey
HLGFvB4WfCnyLbDgdokd28IY7kDrbg+9BrA0O+bDnRh4Kcq65k4vDKU66DPEb/ix5WqyyuEJJ2NI
6O6zfenmreLUitBEUtwM3J0Dz4MFMKnBWNftwrW/oBfIhZF6HGIJnw1dZsVkP9Oq543dtpmXhAvE
Ubah66iINlbWzLswx8L93vlS5rftEyyTCkLkxmcz/6ULUuX23xI/GRrxdioprESZqe9av3wWH2LH
QiCnO4OozCQD/5tKvye6j/7qraHQLjAQnbBmPJgZzSRqlpt3M8/zVqxI1tQ7TWY7+lPc0wRFkVL5
ovrkcva+MAvLfunCLz75XMY0l4VKAOeYJsYafZjwY1zZr33j/I+wYgXwVPTKH9g+XqVeXK1tUAfm
F4cBTyH81gF29equNndX9Y4BY7M037JJss663moxxxgqEjsDYWCNRe2t8bxexDqGHggBNB/2qi+p
lavhcUcqKZPBWA/9W8PRHXqHpQPUy9+/pZvbiqkopDLyQjyLcE+1qRW0hLhPpGedrrTus3S5Z0MT
dUVEUw2zXDv8oySAcG3IzqIB+HxYFgJkFQ98y+muv3JUtXM4xSTAiZnOP/hTWdFzeZB24UMyDwRL
Vtxn5H2+723ErM3Ew7DeUqp9fnmk1NqveOPwnZ6sX805sQGnNY9YP75YL/XF9lIpKGTmjHA7Pt75
kgY3Wa8GR2CPkgYiHSy+4ygkmpFSPXRpMEgOkl0xL3RrbEm92B1diEv83QryyO+wxmqfF1izIMML
yTi4Wcf1n6MeLxb4n5r+zpO7w6g6TCMhoITnq2NeRK6gpylF1vlGAov/ihqXXdTPCjqpEWGRPqgS
EY20K0J4AgMHpGxgvH0VoMf0mqY4nSGaOgE88hdLdUjZWmonfQcu4u/m6O2ytG+DTv01r0Qj0NfZ
CyqrAPKiNOTlciQcQJWk0z1sswn+HoHPaSpPNs72Oc4dGv6UBHpMJaBpKo7qKS1t9YiRw5nWh3Jw
hBctKE2te/WErlj4Q2gakJeWD8skN4JGRE2kt2mN9V0LDNqG/u9MqhnUA7iUj2iHS/82N4oMGCw+
s489y1Emk3uorm79pI2OAzkdfu/6qqydpCKnPro3rXHb114ztLAQaQpi0Zgqnub9tL1iyV/O5ClI
mI+cOp+ynsYKO/O3BWV0Ca4grJ7SeWOZuczlQeXuXVirDCyBL+eiq4UE97IHQoctdyAHCIOae073
vsXf26ZXddghRP45rbUZK8dqd8rHzouyPnXnQTWP0PCet8CR7r4W0FNxbheF4xg34yVuhBD9T5L6
obLy4wX05YlET/13j36vYw13/t5lMNLM7B8URbNYXVAS/YPMOJpd16bv7SXFgg5raor3pavlDevP
P40Ve99QazInUK4oYlEE/sTVM85uoiHUBZHIkhJhjkm/FrU4evbjsHBFBZw+wqFPBQnzLYbhvEcq
h+DWv/1ndeJ6XBjF4sK4S5qWCSL5IQ694ByD0Vz2/oSwPdGM/q1p82fLif+U/LfoRo/x6mpvzPaz
SqjEK8WVC6Vd1Z+TxOMwSZ4THAdinzj074+/LHDllWt+XeUItDVBXAYL1lXeu6cUzBY4KJAzS+mo
gJ/tMJXiuX2FgOJn5HL9botSc9OobL1ZzEfQ6GJ6YM6CoepJG5DhYmaqOQbJQerqGRKF87oFzUwb
DVR+jEJv+Owgn6BjcKGp0iQrsNX7XTxIR2odVBGqtI/uMSQiUtKyAOlaN9UIEtlTktkQoVyEbRtI
KY7kx77Fr4h7QUuuS6Vmf7+JH8zUbcF4M96BM+ViZal9cMTa/qiRjpN97REqQVY6dMOzzatE1iPL
uJx8qNpFKHZB2LQ1WG2Q6aKa2X3TNnlvzLpRFuOAPrl6x/Dq4pW8tIMYxTm4ejWkoPTmca/xpeZy
SUIN6x+wxvdV+51Yvh1iiawEkdriO3XfdkorTH62aZOCNZXtTX67qu3P25lwypoxGJs8YUXFRrlL
NbJuaBnXxr6MiYBs8Qcfc6wCJIPEamQl+yCTo+Ac+TIsA8h+0+VsrzzpABb8te4PtKdAyGZ7oy3h
ktRk5CH/WB/El+qI83d9oofkvUmb3SfOjSgnvNLSwCewPdtkqnGqoGnNBnQPA5PrwgsyM23/5OcZ
Z9fLFi3YTk0FuM7xi0+C4O9jnShX4jivGmo/JB8oru7mWQdECkvlOjTNnpOff6lxj4jeUo+GPNnR
OxS93F59dxyMnX6K/MxIQ6n+T+JA7RaCHbKYhbHEd0jG9AHg4rXJupldMlyO/4pmWberkwy4s4Lu
nD1yfLxHHQfW5qAV7NK4Yc1e503S5bhwrly4Tp9awAzB0dPFsn2EZjVqHnUHe2rNigN4F62vuCaR
vEUzIkQpEIH7T7weFq5z1Z3bTJFSbxN5mWAAXBCjZT6J9fqHKZHsrYRATXqibJLuIuENq4arYQl9
sknluxlOLhCahqtcQcY/GqH8SSI2V7fVpie+Cmnal8edGOuToUKL/pTqjLDkPQRwP4Jozilkobrj
KaN4NYG5Ky6z8EeNLiePr1yuKtr0c81/T8jMIZ3S0S75DJUUIK57fm4pBvuzsnPTrdg4kh3V0DHS
Cy/f5L/gSFMS18eenXUbiAF29jXGteLffH2kyBs2ISjz80INy4JGVh72ebN2hbZXUi1n5qjxuVwV
C3pmig6dKfG8FdJxiaQTOqI87/W+IvIY9+p1iM3OgPAWAsdC4C/4Ign4rBP+y95w+kRB0DOYbuSz
egIFzHpe8xxVByUBHvJwG2KikXDIv7IA2KXr6qiITNYqEZVxG+mSOkPHzbzRLUpbWQ/D+J2GWu7U
3D55rgiw9FkKRVt19RPovp+i2Z3OpoGuhQVXN94sfhbv0c27gbk8OrqexJZJrA7I7VnhB0vTpR4n
ifWgNWBLXBZxnEaz3fwArzy0wdwHQKNp8hZ4R83sBGaz7BPMbxgyKqzL5XbubmBuNVTcn4Dk4AWG
cT09Vp5gqO/BuB+V0QIpK0H770jBKCDIJw4sK+fa1DLWNX+brATzqBTnAoIJtn/clf3v9N8icoQt
Jfix6wEhsgODv+6QmJtfjyZOcsTPDgd99koxPpVZUA/s4f9JKfQp+4DP2lbsurrufedQxOnr/g2g
dfboQ3X6d+/WoRqnT7WfrDODfkrdEgOZ2Hap1qLGNzzt7eA37HO7M/0SwXmyGu5syr8ObFPMJDaB
D01ztqfXkhbc6GAEVzusS2YMc/lcpVj+ezdxZtoiPZ3pl4DzY9CDL3x7JnbB57cN9h4wb4KAbotb
jGLEWmp2LmoIIodCltKSwkJ4E3okTo6BvzWpjei56Tr5e0SNPIC2LtuNVKO9vEahFwygsfBAWRAS
xNC5gquvarcCIcBcME0mGtvR/GM/+cHxhIPWKVOrtiuhyghBeynv2l4MeClJt+XZ31+UWEY+gkGf
WOcmTA27ndWvrtHKnNid0ZdUVbfn+x3eY5jh4MxuddqertKG2P9TDBUcaUyV+I8H/Y++zI3zFBRY
Ns9TnwAII3SeCn+836jXm5CBBERuQ4chYPw70C9nF7dN4ynbYnhVrIOLZB9nWEIZKKVLOJCCAP8x
vseM8lQAb0gexxpkdPOt4rMCrcclqjBHn6tGe8wZ6gpenJh3KmrjwHdO1JJj5FhCeJGidAILI8Jd
gVrLguCB7nlG+gm5sZ0vheILhrVuT7YIGbbPw4gJLSMWFglyVt2/FzzQ3zcSeMe4g63ifSPhCT/j
VCjrI1tZCNXBOf8wARkkFsGTk0GW2X2RsAL+06BzJfK7i5VzEXwMSsAzZfc5IAqoZsFUeg0dcQ/K
u3xcX8DCmn0TAJc7/qMqvKu25QNqpNLqTGi5NahY7wezz9RHcms03nyoqYhIDG1AADAT0gkftyEE
VzIZfm1BpxhfqvdEAV1WDXKpEAMFB4ni5+OX0VvZV/J9ttNEocj069cyBPBi5l+G5M6L2FqCxuAQ
4oPL274V5hXXy8AIB1N6cr5UUjN0mvqlLDtUa4D+uFsL0Pv1aFHPHc2g2dsq8MLZCJWL4sktLMj7
cSPVY3BWP5Dg4Z3Xtr4LXh4jw4EZw/99UCVWpoxloWAiYbfMpVMZ6t5CGMoVknmxqYG+tN9/Z+3H
sDTese1Fn3dVIicAxToiULt+h0WJRaZUSvy5EfZJ9llWndkjO57hbm4hIyArVgZ6izj8xFim0Y+m
1u4L3tbCMy1ZsIxOWPLi+qYx8n82BA0pzViJZgYHVYk5tlErYGHjwwjOH+hL7AkVyMdlLiXDibg5
OJsuQew16t1/646WnLyN0h3g0G7SqxWz/DtmO6WRlFS6eVIh/LC9xO2wuj4OP8Xger5SWyYyNgLN
vwuayOd1jaknXihed4XR7CXmGGHNS4GMXVFep4/TCQfjhXHAUqsfgABbkFrjWRGTp4taQ0emKYsB
9PI7pOcxt5JQtv534GgZnCVY2pkuh0RxruJ1UvASHv+0XYF5XXfwMbSpF77gD/sytHYDFc5n0pWu
fdFfY5594DKYtmzSg7yBWaWSLAYIioPjMqiA6XzqEiqxj1W06RlbQJ/INGqj3ZeNKfsNGsygQoNa
HRRQt867M/YmHFZeG4MZQFVWQKFMyl19OC/iWD4VybVfpksffRM/fVL5ADrHgQfv6I0Zp9Os09tu
AGeh6e4d0aCFTdwDA2zp+9EGdXwmjPimSOzFjIX5crxQNff2LJKuI2+/oacDe+yrGy3lvPv2Nfu1
jUn881knbopi8eh7kP1h/+MrMK3FxmDnejSra1WecE+T9pjL2nod0Cdl3k+nwnr1cluD2rsS1pW4
YjRrbSGTcMrGFsl2v+Keub/8Db8I6E2/EsEnLcpQJEkbTNO/4BfZa5HMVz+Ew+CsL7c7zhO8nwTe
V2FEPvGhEeQlxxWeCRYG1sTy9gJE5kcihvrzc+IwNPMeWBiLQrokv4/FpKN7ze0cSXu+efdez12y
eWdoVPcv7OMzOx7ZB+cf0jDgPzmuuYuY4qB9Nv7wzT1Vx1bCDsoG9V2YL3Emk+ATC+YKWhiQzzlO
CKUo3iqVK4nx0md8ONnxxOEXnPARp2aMsBR94kCNPkxxcLe/ta9/lI5cpoIoflKM6tM2CdHW98Sg
iTPi+/EdlzNGdji5vGqzzTo06snwWCJrqAmPwQZyPHxkWvsMxjyJuIt5HGa8j4V7bWs10G9iMOZD
stjS8Seyaf+QhJMLrd+M4YDF3erENbfUQmxxHPTYKUySXD8nKLocCR9IE/MRe2YDd99LocCod1n0
zsBRqu7Cj0+WXKBoFArCF58mGklKqq0wVYu74EVCa+ZaI8pcv9Amf4FfG81NE7eR9/sZ1cP8tjxP
ShcZ6EfNKLzsg0eHQQQW7qK4Z0ABSzGSUft3e4yTjgQy4xfAk4dLWA5CIoZitYQArUH62vka2PAG
iXVSkgLUMaAHYKRlbaVrByXFMPcKzR2ZakDBqH/uNUoGTA2V4KQSeDxifMuuFqL0DqAW5j0oWrKG
rMNs3OVPoztLEthy3j4dxXVscoo3SlMzXzJPg4/lYjBcDGF8QGle06e68wIMqp9GZAOLPMizvChZ
XrrIDcDX545QZcz76zEBR7o7cIqimAzuryiYydT5XuwaxJRcXWlGCVImSZ0nMy8miUNFyjzPtiLP
rTVMobqqj318PnpDCvuNzka04QTDV7w0V/JvqvZTvksXyKTzICsXLO9O9qWi2PGxlY1L/If38+Rz
frRhnr/oT4I5iFRbWt7Tda286oPcjnICVNul6ENA3lhmuOQTBWqIfMS1d9yX706QpJp8gBritlfG
64gBBpbtKXTzUbuVeagB6+R1vm7dDIvzQZ+jmUcdKZlTKBrCyN9l8jTtkp4agmyg8ZvLUQtO2EAv
Bgl2RdJbvYENE5SK0b0ZpeIEfZpF/nNIsuJqKdpZaYCl0Dz3K52i7Q76zENOl72oBqNOVaP+ZKZO
GJk0rSR4J70qGiXrHw/RCPtZBpTu/ocH+Hcf9IGoudDde2tG+9+0/z2ZutkFWuWHC9IPpPzd0DSa
Epm6S7N6wrznBC9WRnTPC2TfL6f1Yp8q156UcgdupmSGeo6lFmGTo/O8iTfvbyXHILqo53GyR5GO
ROcUD5JOim4Fp8PF0NJqBGK9k+hF1Uhmvz4ksHVQqNEj6GJ6gtHFO2aB8RsHWRU5Ig5fx7ivD0ft
DV3a0befI6k4FQYxeiiqvYlSn9yZKwYEW89++xd16xrRR4zGQvDdK9gfrcbrRVCXYUPOaAK38k7Q
zNrgBQ2r2/kIXY2W6BIOVKoJYa7K+ND1Va5LPHzpwM1JTpOzL8SXamoS8iepgrBni3S0U45/IAOP
rqMgYvJTAmoAY9OJKU5Excx2UVAA94DAz+J+qSyoDaeC/qwO0yau88X9lcx1zufL8nCxBFh1i6fH
ddXlEdrS1qHhQ3QAMVzNixoOQx/uUA1qVY8Rf7mh1Iif+QSGxb2qxXeIWuKndOiroVJC7FJLux00
NJ5mu1iZqsrqOqLz6d90bjm2KrvD4aIUJ+71wkpi/5pnxT2W9pREbj8tP3zLgd3k5N3kuKo3OuNb
KvNPf/zjQ3iRGiryhTbsbA9RGRjUvZ5qUR35CCdsbWXDRYa7baCZfl2YkDk2KCHB4kXQLX+K7Y54
az/UlCe3//Li1rCR6RIV4cP8OmbD2MZMt2wd2U7XYnfazJN4ucg3gJqR1DWT8JuwEhe7Iry03eNJ
+FBUVVJ+ynfrFWT43y/geU1rP3KwtO2JTjS5IIr/MWziUck1H8D6dFR80ozKXYQiFAfh/7YP++4h
e9AgBpEImVdckZag6CLFlJ4Al0uL374GSoVyaykXGHTFtPAZCexV7TdcO2MPabhyeULepC3KXTHO
Kp9/FAbQaTcLb8MAr73DDz7jUW/rb3/5PyQo6q827hNxECDsWxDp/w1qnxLR9Y9ah6AE0PBzOOm0
K/rFQsg5VO4aYiFYPiD4XkNVCsq6XJk48ZsvDAtFoJSiSL2bfVP9Z8baZwT5nSJb2/X1HOFssuDP
U+l2kM9mIoIbdLsrinVyN4+ARVo5vOUpH5hWYgeKJ0AoDHuBPUU3myxjtDQha1KQXP0rktbmq21d
u5OL2vpGNEHRLhj8vjhTsV2dfwgwHoVodAdzYaiJtSPb+QTLz2D73QgavJHI8OOBLDIryJ8JD6lT
44DZR8sKpiGZBGPb3ay/tywTZc3GMsNOnUc8gViq9Z86zZRb9jW5F61hMJvZSrmRtnPnjT4DU8iz
wgNtRlTLJOY6Lh8fpUGm6T01GNnQB4iE+RhJU65JpsV1hagpooeXOnLXZCcelEEQxnpkLX8eDrV7
HfV5F6jIq4/oxPYWbz/cBrmvGoduzzXwY606xZNLUVaj8LlOVnW0Ln1eTqDJFvGd26UXZEtteinG
zUuzdJHOuNB8PuCNo70h8TXJCdPkeL21d0+0kNfj1yc/W0xc2dqHA+4DWoemtFX0EbcqsX0s9G4M
Q1nucUpIVq9MoGNb9HW/Ds5geZaBMK2CktSXBqDoh1M/vsBCYMfoZjPQQFLm/qcaaq2y0kZaQeOm
hMBN5tvx544wTsHCDjIEUKgV9XxIQmkBv9et0KdYK8gBdTN7u/Ib/gGJls2gQGS+p7J5ouBwT/hE
Ftf6tso8WBWCSj6pXhPSI7Kcp78Ig6MVIcBEon4jqbJb7zY513BDqf92Pmq9Qc1yeel02W85/jRY
rAb0hvuOq1fzecYRZ3X1r3Me7SXzgiZR2zuqLqKPyhpcjYjTfU20LdTOsXgrjzm3BgA+CCR4CJxn
sWW5sikc1teCdICWf8GC7Q5+stCC4nx0GHH8DUzFTuip9SLhkJXHm32W0oZZqNyELk9zgAqQP+sw
WACczIcZI2hd9AEiBq/rX8D9HBWCjsYB618sDOUeF490R4AD1gcddm85nVxmSVD0F7vmJ76MpZHN
CpBXACBH3rsMFHnTQXj509C/KH+FoA9b+0vwBfEVosGRphqqgtHmZ5GFwia6MDKyiUl9ON6KBzCV
Z712MxNpKvJ9S5Co1SQ6d2mom2Gm4o89OzNgu9UrWsPWPTGHwf5BcijZG4C0RFpcmxk4No3gtaHc
Foa6Ex7n5Q9MrLlXA5LcpsodW5pBupy6JnGAZOxu43xBPVH6S+rMIbPGQ9yGJoe0zejPpfAkx9dQ
EZKitsLMHE0b1gSlQ98r6t9dmwm96esVF8meVvwNsRVK5pe7Fl7Xyv1J3xy/EeMRB1LAl6rqmCPk
xOvxWt9ysmAMXLAVKEOk9FaSYwJnMX1L89BuDCSjBKcUtMtyJiUvEYlTwhYsawcDPnEu58qz0wJ0
PDlvMFsuL1Uc57f5BDXTCa5Ir97xLF7Y4+2A6mT0EXWpBrvyt4ny5/TOe8qqNGasmKjehseDy7qh
MHcbkMZ0E3RJFCVSH9UtYOYm3YCcd2Vs3zQ1fa9Ai4V7qCQAK5cuWcO3Tbx8kkSIkAdPn+c7MbLD
1LXMBzrccReffcuMq5bMXg+U3Nf0/TDeKGLIrX4oVOZihPQEG0psxylkYJdk43S+1TRkIEmnICHW
Pd+N2OLSw7KqISyDAIZr1KERbKVXfEkJ+Jf16Tec7hX6Cy4WIj8sOKrXa4eZBL1wuEEv6TEa2yiX
eMN/F9SN+tfmoxZyjwideWkcIaR5Mmr5Yz0k5dtIQx1G/8Z61HbYxC6nl/qnsHkU4scWcbHAD69r
tKAr72zV1zwdaVqarETfpna7XUfE8TppLuJJQeVrXqeNK2zQz+Wtvvmp8ZFMtgVwz05EGHbjrcDZ
ML2TeGiaRpCwV8YlHA2VTFZw4b5tGxocxgKBfctnZaDWs8menRd0X3l4elBGNCpZAmr9RTjJ1kaQ
tMGKStNLhuNv4gSJiRwHXmxaC7w1tOSDSaRe9Y22neM+d1jQMkiQyPiHCp4g+iY+Z+XqefFQjWav
hu41205++Iq3f0BveqH522rNZp7fuwkWys/oIqGUtXAqTr5u0CVQHmRiNnSdyw2VgXWCqQQtzWxo
0Z3v/xLoFt5JJ5IFq2aNp+EDleD10Nd3FJroAtFJYJw20WtlV+SeZzIamW/TTnO6p08PspDjVUIv
3D1nNMt8eSlKGYbVodFa0MuH+qoUevt5izdSPd6hV4jr9rjUjhm0PAfiIvKFyBby5OLMnaVyOuE4
b2T8tCLwmDTr+zi/UtRK/0Z6Eb1AuOOtbizDwL03DD8upXa00qzNwtDiD6gj4SZVlGHqXu7JN19L
wIFjgTfmS1QdxFEpZ1UYVXBQeicqSgZCPEWZ0Bly8cLk3ouzzEUAAtDmlOIh1daYNCJPAANTMNhi
ZUmRkjltDfeJ5w/kgC1UG7nhv3EYrxO2eZbUrU0faPUYxdmVRbPpDblGpyrcodS7zZK5S7XwPOWI
zzWBBega8U4HZyggrTh+zXfjbrFWFVnQpvV3BYiXzjVnyfOTLcBlnbENspXZ3DVLEJo2aSpHVN8j
2RqiaLOSbFuLP8dzlidAJuyaXEejAOzygLLLwzypGTlgwHN2tS63UsPAD3hf7ModH502pR+INpJB
WRH6u5nDR0m8dneivFQ1zDf5ua9Kj4fLNJjf4QYrEGONDyQgLpsEydfbIMj/pEpto0XhY+2Bdv0P
gmCmJYJG1NnsGvNOyGQ6zBTkIWzgoUfxQ92NETCLDFhJM7KWm4YbI5laTJjcW3bXev4ABKWWTt/L
HGLXobQJJDxvXthxJ0JAGfh8O5A3BWalUGl+sot02Pyd/gREjMVBJtiJ093KJF7nlP8nS7FdPP55
oF0kW5hOTKCt6YsO+JGkTEC4AsCQaPAI33v/t+a4Pq1KPlPgAJODMTgyYWB+2g2K+DodxPtQZ1rd
3qLe61b/KKXSUNZMC818IXl0FOfDxYSxcx1g5UeEAHQRI2PQ+YwydqedPkaUBp2zqVDBHKNbxAgW
dDCuW5/aD8oxbG4GFGtc7gDKUEAZn/Ij2lqQ2XFw1mKcAv72JSnuaKpJtqWEMkciCPLjQ5K/JXRy
MRNNlaiF2W7f+dpmK52pV6CnJCHdjZgjnQwLVJfJ2GCOneBrtqwKpoI9f824IGIIHz73M7G23Mt6
lT2XMMn/m9kW6OlWfOCuu5bRP02FnO8foPvJrRygQO1g9z5F5q8BSM4KFcydEdjSeIcEqOkW93Ej
k+zxE2Blut/MMNN7HXG9P9VKEZ6XXlGrNMSVBBkT0dHToZoPQcz1F1lzw8m4dNKW53OpDm/lieXh
6dl5j7XtAAXvoYqo9IT0jpt8VgG9mgKbhrjjebDsLfa0clJo1+eZ42JUG5b0aSaNiu6ssjflP5tL
KZIL/W9UfAgzRe35ABcw8QNfGYoOULBoeqFRpQ/fLz5nHrhZLMZ3QOch2kcjqPDttUGL0CX8MMlt
ij6qVvhQXhA68FKhpyhzB0MBaU2VE+O9veR5jTSnV8p5FCXyvUF59jFGG4X6q2CCtcvf93CdiOPD
vOpg+6IqDWWn9Opn2KCWEyWVUoY5nlhkX9IRQrO11CCqCTtuAm7NijQUyfpfStZ1qUCmgNxx+UIM
JY0b1VZDBB7bgAkNvGASMQjqpiCSK5wgVvYdOZDsOoOgXXler0gCvHFVz/1TTWpLHPk4l1i+QOEt
H+H8Rx2Q5+KqO8W6IFAwXAHSMG5dRRtqQM4fVr/di3mKl04HjRMARdiTpcyL0mkJ24tsQCEqvsZa
jHj+Yrv0ZllGhZ01PsX5UNy3HNn2Ye4mZu3Bs+Amw2y+p4/CDT5NZwbbpdYfm8fECBquYkgeeaQl
aKN/GDxrt7ynMyJdxhuNpDz2povhk9MxLF4Y8D/MSlRrdXDuJevymzTYsbhbkz6iA6wPsBafjVcg
dwlEEQRiBWNshT2HqGiDYxOcdhxUwPgZ3yhL+LgIOhqftm2hBh2q/BNJr5cx8H6hluzNtj8+svAU
xnTwvj6Fjkm+QmTBXjivXumG+peHOY26/Sl1UNaIlhN9ERqwu6biNgG+SnCK8PIfrrpw84OUCLeK
j0KZUSgTBMXFO2+Y/1sniA1YX8wGVVmzlHuPZLEfzGRHW+OiKWrhZFdvfo0xAmvDdod5i5OCydZu
/dqLkGLDdOmdxrdS2ZBGa9xFTz2OixOw7q7hHq4QPTPSbKyedtNwi6JwblBK/yRduXJJToLnf/uS
jsLzphlIOceRwB3vr2uuuKLPlfrbO0pVe450RNmnnCGAlS89vogp9a0Rb1pAty59D8crlftb22tQ
bi7c8O4YbhNkyRMJC0CJxRGMZ1WD485ku72nTAEI/vSNgsj203O207t3jz1zQ8bfy8SNuujxogAZ
4L3wbnM20ASXqDShZPeWTYDYwaZYV7qRlojOFg9rd3Pq9OxmKk/DHeAS/DnM7I/dsDHo6+p2E87A
nMz8gy4tNgCmNu3161IC31BE2GihxucEJyajrOUyhgq1haDXTmqlLveOsGON1alohz4kc+sw8aiS
Fdl1et4Djt4MMdd7oa9ASei7zj5UWzy2+A3Xtq090pNwj01uaAuz6YfAw7JkRUgIhcDRv2HLAaIW
flymp0kOMWwtECY3lRjtkIkHFBpcOR2pQaMgl89KmZ1Pedq/WY2pQJaxNid/qBMUxRg8bP03xd10
Axx3/joquz/sBxaO3JocP6gDGposYgRXfO5kwVBB/nQWUIzhjdCSyWnM2RjMZEtQ7tZHLih5C05X
JReBi6C3igDZDNUNBgLHiN0KwLW+i759NTKpDskB6gwKhMP555lQZWUahXmcD6AfPaBcYi8m3TkR
5B+WMNsxWQ1NUy2Fq/RSRf215d0Fw2xDZU5+0IsOvF2QgJ2srCTlsURPdjxz351NELYFX6DGyLah
Cds41Gwbm12z+WEal9IPxzLbyOujmja8jcgVmafrdOUW06nIxrsYzslw8BgyXLuw9wLtZbCvuo0R
H5DQQUsjo/B5OTei/b/hcmYs6ZV08xM1NuWcGPejtS6esr3btZDCoW35TnObuRgHumifGrCfRr0z
/MItzpDUMUbNQxZArNROaCZ68yfzTeAtrb/RT4FwKJoVHNCYOQypcS0YqxnUi8I2Z1kDZABYsmJ3
3ine4bMF/R2qhQvkPIClM389C6ymf6Ovt0+tXQ17WFlRfyhVSpcLb3CHAtG5pQzRHpto1J/N8vIO
1uFpEeRH5BiSgsTyyosZQEjuCgOP3QRgFY43wKQXnHWduliWxtGl1sdMAkDur1sLy4co9T+P7Zxz
rPGAdiNzvdmUZs1Pcu+dcFpOWmaS+SjAO1pGcmNFfVwyDV3NkojG8e3SiSmjYoJIrzapmBHdJn/p
uKHMEBRRU7HvscRuzSyP16FLVp1VGrktIlYX03HqoBRThdvIexs0n39rF5xpg2wnAKXfe8zPSb8a
pw9G5EtNrVmtwdzwqHpPY5coZ6HjHexY/WfecRlZtAS6quhV9a/eJ3+LUlCLjg82m9yhSU9e2EDz
H6zUGqG+BiblXouRiAz5372YH2by6Vl1VcNrsBPNAxIEFb0raJjCRyB2+eRGlTBdl7jvgFzEcMAh
ph0zCIg7X3piG06oSYcln/MB6XnYGbZFvTsJRzXQcWFdBh1C5c/gIVCav3PwneMhml/mmLONiAdH
s176g9DVFSw5qLFPprXgnUq57KjBkskRB96iWTM/UP7KTDk0PvExQcYqXjQ8PJlt5HZYrrYzaXp/
VZM3k0qVz05Z3YZz1oaUWcA4N1oBrxJcTw9UiB0eHfiGXoTe3HXms5iWiPGo4OnQ7LlLWKuy+qmh
Xis6P0CGSbBlaraDWrP/ouI+R1XLRAPYnyQgc2gkJvZdcOPZ/MDqsG9YCBRyaf+5LhgeiOXejR5S
lNtrE1YwZ0RgNubYsik7Yl3NZBFcIlc8Df1d6bZT6mqZCyDRTnyBHMh1HwAg4AnCbuM2/RX9NWvM
bCB7ngZQktUQAXJwCahN9rvuBoX/N7Cl0R5RIjFQgHYhuY7OzI0C3/ry7OUxPo8+vhosoIaZ+EEQ
2FyZ+hKUqKxndV1usz5eZ6kZrT7Tw4Dnqy/wnUjgJiHf8o8UWP5JPOtkw8fTunYKtEav0XitDgqB
QDoehWXrVq8AKfsvjtTzh2Ah+R8gAQ/iZM+Xg60SR++9Y1MqshGl/+SvvAkf40it0PR2Rv3pM+fN
OQ3Bx+wfpNM8SGmPHNI14WlSXRS93UTq5pnqy1JXed3A3ZmvCxM92yADV2Im/v7MbhUJd2qEeG0g
67HVyDKLj52ntkqx/YLWVk/YAoVRy8w+lovDi+cwQcA+fAQGvxRNr87RYaKjN9YEsWzyBoPa+uUA
ut6YS/1RmIH4BhWeC/BZHCKmvhooZfWbfXNseGar4y3nCpTzSGiJvZd/50mqCBDoisBMk3VVim/Q
OY3yoWmzkO7oy3nazyCGo3HKyJ0cn0N3OVJQmXx+PDsPkLB9t4M6KX1230nZes+q1ptEtFgLtLsp
GuBoml16bQdVhm9Qu6axC75q1vgLXc4tAo4IZIIETZoJEWp/QrbiO//Qu3koYoRAPfEBm2VqE7Js
6GeZKENIJVmHGSqBriSXS/CkNGO3ZV9EP0YfkINno72kbiizZXlmZsVZy12e3wdt4rf2NSNXdCTA
yAItasgi0Kziq9/5FfuGg+4XlgiylrkYFEuCNfAZu/Vnfj1CrAq8lrmWfaWNxwlWoLjxWP2aMneD
NovxUjgM2QK4HkazoFQrTgsjLai/x/+n4KNpLBBHe6lvlSPoG/AFI7a7mD/NA0sMIcDgp4j7Fa6b
N6MthtLHOlr/fRRQQg8HR2U81NPpH9mir45WjRc9SmFAE2hJx0AJq5dR50D9z0hvNAvp10jiPccW
IoxZ7sW1HkVJBPlamAfFJ4VTNaQoackj5nkERGfGi5LqzT/1adtXHIO+LDrCCIZixHrJGTH5EAFn
16n9w+uIMzMz/n5WxQyeATxe4m8uMd+wCNLdBSFK5PMNM55APT15ncQ82Ajzny8RCVbjA8/8bJ59
aoxOfQ40J0Ee5YYf6JBBQ19XabwGligWgbPTh+muxMlZ3L37tHOBcfYjnH+mRcJbvb23x5LxDOJH
sJtH13tXxMiv3FlP7M0WRjkUXuJZZ82QHtyzcaNKOHln4D4QRTEMYgYmFTQ1v7qssv6HQGG0Llla
jnJWlrR3c4PcQGg7hxDAQvo3aOhsN97Pf3FP2frAFEZ3bkhv2YO9X+cChHstCYQlugcpm4rEA0tz
f+jQ5GV+c8o0p2kWYrg6XhREPY2uFbAZGo1BdVY56MYgsmjUV/a8oQA/eRO/yLJ4OhXbkzxAVELE
HlLswz5K1UVN9jq0zGHL9tlTJPOJxzZrpVyyJ05bfE2nUQGMLKlma143NXh5cke+reZWpl4a0Rt/
DICqOMvTVhBOnR9QFzApW0kkhbNoEtfbcFRT1URv26Mc1uPEffC1eAZWuBCnFYih3DUCaKP2EmWq
HHzIA++GtTcUCzUuYt3j200Nfp+XQz4z0xjMb5pDiTNyWPKGGcl4X66C5l5OpWGkeHLPfi54oZPQ
O2IUesNA6SH+8rm9xHkbzAuRoYf8YnF2V7OW2SkBVRnm1tOzJO5XH0cNQ91uY7tx14CGEBeVdYlp
qdx3Uj4OBfnrodqKkESP6ZDRfRN7+aommXzXJvakLW434K8FS+nb3s/1KB3Pw3hL+7F7dVJOcUFN
q+o8u39b91SuX2Ru3yiy28JJB8+SGrAehre45KeqYft6bYWGjAV10hWU/NLM43TkBc8Y6SRNz+PU
6MTQWU0Rk1VUWrdcppl9O7TuLLw+4cs+JzK5p7oX+uysFxWQvBqVAnFOfeOrElU0vEMSbH/VKNDT
zj2YfDTcuSUV9ZpbW5plI/47DVjaB2ReUYXYizbi5aUokEhn+3tMlSv3N80B6MBPStct8RUUWNXA
y/VVKqH9JGdpln1YPl8x6RmhB0lcCjo/uc3arycbk+LGSVU7Jki1QMuICAfWP8M3GfOgIfBPYOFU
o8wtCk/mTpRAITxKANKNSKT2QLVCuiq2dX4Lf7yrO4WseG4HCHXlWP/EuGuvXnr7H0wjYvaG5cli
GYlHTAUW/UFb2WgCIzuFtrA/1fLC5/ZFVL+xqJvzRRXKEp6UlCojZLaxbCz68hUPbN8feCWCJeEF
uz/W1CTQH9Pws+SxiUMpGisO4MQyG9Oo8TnZeAUC4kZVtvBqPXKvypfRTE8jPcR7/pMxd5BATHHp
AX+MgXlDY+T2lc0FLA4NyfMPw+XvIo0ilsrRkolXJa4Tk6IWBWLKLZXCj0aALroVL++fLGTjQDMH
ZKav0pb4IBtGocT3FXMYxXZc8wH/qzFfrRBQafZuZyLxEBPRI8+Qg88jw2ysaavGeJAwtkUYAsZ4
NhvKjFoosJzOofWQ/njm0BIBYd0im42tZ0Rk0Gw+SGOMR/uUR38TjGrGa8snBz6mufbqXFHjZ5e8
2omOtLqdtbTIUpjOjpOyJ46nLM20NX5efYjKkv1Q6vG4BSfLD3Yg5BYhdJAj1QXCFwtsP/okl6qV
F0N6eQnH7yOwQVscSchkMD/xbuzSv4wz1CC6gpV0rBkmDgXSh2XcCHWGf19I5FCesEvgrvCNSCGn
nOFJ35+Z6mFxU7QXhvJd3DTjSEcmghMgxNDLIsOijiBRi5og6frRVdtHA/j7HoZ5Wnd/EJ9KpmLK
lNScvzNOm/5SKaJ0K9i0sqCBQM4ViR0wz34CvqiHB8ka9ulIsXTChMO08Munc9erDUCvw+FsVUN4
jTnbkrlBDDQBHjtRt8S/1J429DxedEsj+HXylyRcAM6OAOH3KPUQBf9/FNZVTsfDHpUdMsVb1b4t
rlH7ujecQw7AhDU0KY6lvqB9Y1Ei7AVu/VnbpirVMuCgGCkICpFhr62OvykRHcPpXtGWWDZLDmh5
QNPM7reVwvu4HtPtaHmKYLuReCdMHtTjo/R1DFDWZhu7Ool3tIB/p6Dr2vWuw/ychFe3/4itPOFR
5QnakqIIe8UwTSscGa7nr12oZQdk04u95oV9eKayw2HDP0kHKkGdFP2Y9888BoDloHpl8tWEn4NR
EboUmX/y6YZ+m00Oymo/VzBsKJ8shRbOlx5X50sMlFooWZgkWDcxLgI1N2wTCWI1MLvQHZuPtSTf
3a7ovTidcAd4MMOGRMO0NU6F8X3J4ptofGFOJy9d+jfGrjq3GgD8TxiMJJaryRPV7DUNEwRTwqEf
B5sYV/YOCN9OO3LzsB2bSiNfww/jwv99grgYFzFpbMhpajql0Ngr1tjQPH/HIZnNaXp5t/AfiuNY
ZRapDHWk+rWN0IB58+ZJftbzJRqsEKVHfXGoV+y4QT92yQSAtGm2LOR0W12TCOXpzlf6z5SpL/BD
16LlUIglopoO48iK4g63KvqPUXMr0cb1h6jR3jg3EjQbZo15nRaLkxrZ/DZLuIh5L3oT/l6Vh+U/
WkDiwmVaLgRBLBBKGMLzbP8lIkg/XfDhOxzqEJSzyeMhHGSUlwKkGPi1nUJm6rOXiJJDBilXWpnC
RVxfi4zsdB1XI/7Vopz+/7CiKxzaBIQzPOBw7AYm0YprnCQxBe3EJ8YS8H+MZnZFWkq8Fi/tsn19
i0AMOGHx1kwJyacD10OwYOfVjMlenkA/cha/kmDzmsZqux3hjrMoKKe1G0xtd1kj+ZDwWL+4B3PS
+hUL8mQA64O2GUu2Y+DOHVdVCUnPsk3n++IpGUlS6EGiKlwP1xQGLO6UUVyScUu16TFZgEo/krPW
VjR3qApUy9yL3JgZfCpBGt/0hBBUpgt9/S1f0D4jololqRpNY853j9mcTki8M/w7Z60tP8WaOQQL
5zQQaPPB8DetIeiWlioQWveGXkITs4inMZYbleFyjjQXAFrG+y827xPBwtuLoQdZg/ZYdKMlrnfz
dBtoF+77M6p4EIXzLq6q8mRXkk4f+P53XtdPe6yni95vLX8/uuzlt/NuSp6zeK1TyozHJejSVGGO
Bwz9mkXuiLZ6uIpxHVdAfJymQXCqhkbTxi4Kff0UFGggiwLjaY7DT94hKlCPCJ503ardPtHImELj
p6ALcS+VNawqVOkge+4N9vBtGlrCvTcL1UrxihjH9L/1BgMSd1f0lRNO54FhHj8nQR8I29bBwW+I
bWez6icJz+5V6pkUj2pprlWjl+D6LBFT9oIuyixE4qf7j3ATQpoqgq1KFhXYrfXR2ng4W6GO7TbQ
u0L7WWXmViIRJmt5Skg8A/WallI2pZVeodhvV5TCgBXWUvTBmxtimiqe5AHhoRifo6uBaafDe51p
OsvvusCzrNutl2uKcCO67LRHO7+ReNPpVUVNL4zeTrzKb6VF5+fK5kYLulsd4I9BOGqd0D2VgkbE
c8IS61AisOO8+RkTt7RD7VFQQgWL45j+6t11wn9ct+d80SjIQ8QHaEnEvp80+A2jWaJTTPjF237x
AztHiXTMyFr50bQEy1KUf7Q1xOUSP0JwiMY1gO6aZwVEyHFxMaoKWqyJVdP9vvclvfU7NJwukOqN
YPJv6RcNKjeflAGmD2JjUKsdQllgQEUgSbrBVuCedumODhY5SuXzX4EAlo/7D34Je0behYyuLYgD
rTfrO7knlvldGG4syV5euwlGdKsD4O9/5OSWTdFahJ8r3dc+EyMdARmB7gs3J/Pr1RcYDjsbsE76
6SrLKN+/fZT3PkLyUrSuj8glIHu2tyR/27Df8VE7/Aec7dhJk+jaLE7pelWq67gWKJ/ibck69bss
PQykMBwa+5SvVUU40hb22SlpBZahloetITZ58ejVf+t5Zrd0a9BUVfX1G2QGMG9BROCYBRYoNdyj
mUWmrjI41OgDxeUuM+GiYUd6bVhhL1akOm8+660e7YfhcbxKbnz+GlLWUOjB/F0ahw7YjXIFwRyt
HX8vb8spTlF/si0aHjlQoKWXYQDIHFAwzLhb+tEmkX1OB92esEKSjvE6HEtQk98Fk/4yvqARrOGY
urzskrPoLbMAoDmvyo5kuKcpQ1EvcvYXYKNHlBp8w9LjYDT72Mu2riXfZFIJBLi1AgMzpP7HMOfA
JGrORNRMAVWdQnjTz4YeXqbOnk092tBFRD2LKD0EB8vcLEno2CUVUNUZAzLglI+P2NjIpjCQ26IB
n4BZgAkjf6bMT0yIdoN/vPje9lP6fJWfz8kmUP42fZ677t+rhcNJvXRpMiEJpaKXa7DsqA1k/fou
qo0gQQNgQT5xsBmDZXQCSsPH9LFtl8RjGKwHsmfV1KBecQ8ufY06yuB30OpL0E2/ePheiBTqQGtp
8mBXehsxk+m9kk1xzZa8eUiF/Tp1+EZHeJqf5ZRxTnvs0rQ5AxAWAocZ+b7hUjbjP0FY7CeVNLkP
CzwmxLfHIU1zoMuh8u3tuq1006V5clQMPPuyGzgrVwE+WUkpr8pwC34hXw6bQpWg3jNtVlVkdrAc
KWRe3WGirwYrLNfbUAN+jw4EXWydD0CdPjsoMtrT36fefQHqg5c8eQ2bVmReiEtfNT4K0KWYwYdM
yE2CZa/qDK6DRTmJZCIIAXohWYJx3wW0o7wQ4fxEqf9ZcH8xQMHtdH/rwTdhCTo9q+ikGPTcP8Gu
189wuCjLSM8jTBnrRTCxRRDsW4UpCO0Fr7qTWI4z0fGQFV5G+yhT4Oz1jlQd67t5ribXRrAFQOON
qKuQ9BFqoDY72172mgxbbxXSYETmg6mR9KIxJQy5KGKqsF4dX5xc4jjkOVm6mu/4H71uicdOCULO
fHSpAeNeKr2pu8CeX26W/HZYCYKmc29uG/cP/Zd6raEmgK9dlyLflJh3Iyna6c7wReULOJRQ9XkE
hAuJOsUA/oWVJXE/pweOUzgwhWIRTYYi6WPFXErIyP4Q8xd//4A0yrleLKReUSn7109QGs+LW1WR
Ls7RTwxOlHyTZo+StP8+sBbpxHvmmdQEFAj0jPxHXeLlkUSieI99h1Ua8P7EKWL2vV3H9v1M1cXZ
Rd3j7bI4mfBrLm/FITk3nGJ1/MA5K96BBESMiezyicglwFAh0DO85Dad6F7H9aEauwYsRT63IwET
klnT5xPoCntJuT1Zqgq2pBdR2mJ38aeVlGK414Q01T9a371DGEm/EeOAGDBWV9J3jpJYxvFdyxaF
stpSLhA2ha59sCkx5d8a+xY1S2kZNd3M0Wo/8XvoRKTNy5WbC/20YJvbvpJ/1YkSE++3B4hZKvCx
HWoP0fqzGUGPq1uo2xrAMF3tToaPw/vAdt8uW47ikl+qwEpuKd2BeVt7Amfl5+u0jNIvRyKItTZu
I2+zgjS8ODxyo6egvBxIUvK8ehmV+XFrECnFM0PUT2bwLhVKLgmb8BJeFoZOnB1DwxP/LvIhsKxj
8pPxb0c8N3vkwwchhbSyrUDeTGGrQaoLINls3tezhoYUhhMu0T0zXCW4UUC2zYJWnaGqIGFKesnc
vRL2S82vT/a+PwmRXMs776+dVOf/tVkxIOrJuycTpJ0xgtvAACUsfvUf5CVY1OINgUuEhfePdkqN
BzlpX+sbIknD/aApids9wCu9gPy3m0tYfNapyItBiPXjfysZQHw56TDzEH2nnqVNLJdwL1a2ZD2r
klVgXXuP1K2PkeEXaeRfJ8EO1MTxi47AGVQNteHrM84o9ILUL3qHKcelo+mYM8g7wyVz5hzUIaXN
jl1roELb7TlYJNUXJpnFMD3KZhdqIXEpkR8Ib2gVUVWXT36nGUfsPX3jsLftGFg/+AeJMU5t66gC
9ctrtkkJstrYmlHRKwUXP+RFoT+DYWva95DcSIMtIM16bfxMcmPkzOL+MmZo//k3jyS+u1AT+wrD
3HDMgaXYWWanOjeSpOI9ut3OS34/l2cvMp5aD7FbcsNtUT/+8EoQ9i0zfr94JttyH1gQOtPYe5Zc
JWvGbjHjraUpGUsBmRR+Ii6DyNJ7v9/x5Ap5oyxP7njiBl7Ce1Dn4vOEap/rxN4Garn7aU2HoEz5
aYnXXR1qqS6D9fSgwd+fK2ZlbeYuFln+NK9vf1hNataKxRn3twal3wo+zlkrCjhC4WunRDDZWB7k
QODjN/6Y2zEpJCSjIGAy01grV3vjqq2EV8mmKD3xKUrFChf8iFJLJ2PVprpT4m6q0a2zUbl6KdT9
5QF1zEO3dU+68RUpafr1ra3qeV2bBP7ciljd9IMC3ZrZWx2f8eLoR8Ne0aonq/SFbbGY+srYj72N
ZiAJVJm4/yXvJhtd3EEooqbnyGKKay1FNoPsFR3SjN/ySCyIkGAXMeM2BWj4pW0wArdLsIw+s8iC
Q/wSFv1aChCormAH5upp77AqGppj4tK0GAphaqNx+6e4X7Shb4sWT/UYvnXhxVjlWy5c5Iv+/rs7
XEbo6Lf1VpnQMDyO/eGpD6UwtIf1xCG0ZBV1QAJQ3qwubQWtDsJ6qkPKKWDhw1gPFpqmoeEftBST
i8NUY3P4SuA0x5PBIu+iVszDfcVGg7RGGpEseReEnni//+Y4DVGvK+vCoVaXoAuvz4mZ9s2sJU+d
jWzVbllC33LAcSf6ztbNCzMueK1BHzxOZX0HPFaMvOWphiT8PdZJ+hJ7H9IcCuA4TlhN2yYUGOPL
f/tsuqPFQdjFKTJswKEiA5s/zpDXqgEO1LcyZbGvmQwrdt6JrJg2YYUh4IKlGWm8CpJP2lOpiui/
NyccyVU75KQ33OTGRyouJJM0/gbczYHneYXwavLxqT/1ssa/x7CBdEbxQQIQhhEwU13MceCQpz7S
EP9LNn3cwT63apb/Dp5Gb5NI5GKSIfpr/DoK5+GAuL63T52cj0WoOpb9EUvCgU0UqQZ2rs8L54BV
hnFYRAZM0bz2Delymg3MWwSk7NYIBgR55VYZJHDUZilAi7Gynj5u4mi2Q2CcE3bwg3FKF608KIVB
O+YsaurqQ4PyZfOpRejZpt2Hr4a4TSr6wl5IzG0uWCFitYk6Rg54EVMlY1CRyDOl7k6pUnUD2tH/
ji6QEvHZVP5u1qPzXaQ2RlZaP6b2zJf3thUul9oG61kgQUn1F6vhaU50dhVoUMbYeJTfufOrtElc
MgleaWAdk+lySoWOAqxk8KYN31vBwxR7UcWQEKdldl2Mgq05J0O5sKEBRdbkHynElu1LNkMQ2NaR
Zc09QQJnNMjxoQjlxBNWxclBvhiNFOAajvSqLI6q2SSpQTt6aed0VfwquKJuKC/OjkZ9SxoPNm9M
1aRB/E4SIHVdy/N4mHd7NwWPGIxrO6I7+LVbByMadn+OySOPoE/ZdZfnwJrgrtUG9+pGXu26Nf0U
eb/04fne/03BBZcLAfHlXOerHH8FAHKFYO3phNJ0X05jyWjou3jr1g7G6nt2C3pPcIIDt9FaLKL/
YUgSl1K7RyFqePtl5Z9tj6sCgQDJletDl/ijd/km8pawn4oLvqK2jXKUKqgN5+7L4YtiuysVHyjK
fw/hCqrwbvyGlgmTa5C5q0KZ0HsrpQEUgU4mw8wDIBDRdIxY3ThDEZrSA+vZpoeAlC+mCprFQuja
YQj/i3mQv8BFC9ohfTACo2dMFp+k8aXJDxHhfD83/9e7tXaEcRCSn1JQoNmOJBVeqxkvMapZEVDv
Ca7SbUjZu+qlRqr2sUaAIy//hRe0OCq256eYRaO06/C1KJ176oqujuBiycrgfwmbrMU6nyG9ePq+
oOf0TC7ImtD2B0E51rrT/YArqBEK0k4Y7Q2PceVzc5pw0sNQ4jN4Y4MAj+t+tAaRPizEUg1cXc5e
/Re/mc9fZe/wQMVS5GXXG9zczcOeXqZWBC7E8AV9uizwQthKC+R0QccceY622vk6HlGjo+A62b3k
BEHTiCfbBNtXxWJHMgG7zXFtI8OPWOpSAOBzQ9ZqlsYMQzQ7Jt8MSv6Cb57tNB+YH7+UYsbSDoPq
GBQACw1EuzOePn+UtTJYD00MQCj2Tv92ad75RhYdMF3OW14vRimthsn2IDpqFgRAsO+jB2lnpb+f
2wfl5cqUMzgrp4Q7iU83SRn5f9OQtHD6VZCCA9SWfaHNbzklMF6ouHiDKdrueaod82AeBcwjSzDv
ILTGDYsfXIwto0VZd/5qtoYdGWtde45BHtpxuFzYE3e2xntPOQVZITBQmm/kzceuYP3oYNeozKei
PyZfQ7Hj9nTskjuKDAwFarXML5gA4dLALSUwY4rvHmjBayQTBT5wgjpTci8D2txrls2j267vt8g9
paHr4z3IQUkNIqpT3t2XgfW3UYHYW8u5YwrCmM+dB9Fn5T6jNKLfWbDQlA8wsrD7dCaaN80ukyIW
exDBN39wIoTaJdeUL8rJSPfPqPHiE22moGENx0/zQBGVvcRZuWKI4csHVpqPEo8GZFSZ+nJoEs9F
yAfiE93UOrZpBOK878kLBwv3IlrxVuO9AfpiMChLLsMIHYV7ZizLGTVbepRej+3+56aH7/s/1xaX
vEHdgMyAzrTnq4V1/qSxOJccECPDtK2GBHkgIg6v5n3D3rpGtz8tNUct8gv1owD02IIjS2PARs/K
H9dg8FPtjp4MVn1NN4jK4l29bf+kYp5v+SHvygblw4xArLTjQElsPCyfxrqDg1Npm1Wyxt4wrDeA
5dqEMyRayDTmtwI6MnVWooh5ywUPmKrM8Pkc3CWhoM75Wz90nuisOBpR/LhoUhvH2oMNqx5KibiJ
jNf42HqPIkg9FHf4iEwbd/kB6Gy7cMxo9Uu7llfGAI+n6pSL5J07GRBkxpchPQ3lgB+/2EXlOApY
twjzTwN/IWr3CplvyTmFBq73TFUoStcSo67Dvc2sKTsjJinj7nDMhQ3ofiuUaIxFNFg5KFaxte3x
a4UjcYxs9MOYbWWo6dhEDgCFUBstgRQS8sMu524oJV/p+gbgNVUbXhYTDarsYc/e5xOqQNvlFntU
epWJNwPf2qaEKKCcU5D+gwkXiFy42vxr1h9q392NP6JQar8f+HctdH1AaylgUWs3ZcS61Shlm5Km
I88goYPY1kTSNU15b06K9224niuiNtKaylwwpBzgWUGds3EfjUieViJIF5ChR36l/N0ktkzcIoBA
zy224T+qpy/sMmfl3YY08iBeDms/ilcpMSMLUnOO/mMDHYE5E5In8WO1oeb5Df7Hvn1Efu2pd8BG
VGH+IYtzUBpfmRTQ78wkG5bXE7Z8GLPsjl3tTTSThpZDm/HvyhLeim1PNqmYNgHctjl18hoeR7vp
SLIArDG6RY+MiIxyfhUS6LUlNl3UVAjqJynASZfZkMNK2t9HavOUl0Ttik/4LZW6d//EZPkgH03c
J1Gp2ViA+fW0i5EUVzEH0bq33SrE2DWDOFyhbLxKXjLCJ8KnScv1E/QRr/a/YavAJUetBCFF4wtd
aiHyJ6hoLOYI3F9kEUD4glTKGDh0MxcpaRaHpS8nrKBLSOQtsxKwsVNwaFNEBPKnlK/0LwHgtkON
yZEgVzm4UoJqjWYUcgBXinOTJfwvF8udxcktcbHptYLtvCGCsDEYHwdk+IFTpeRE3PEj5wTIJbuT
yyRJmU5Pe3zisXEoJBbwGA8tI185hMq3bOwpIxOSvbiUtpCyPxn4ZOCJi5wMW7GEO71Ge2cO0w0l
apKnJQWY0lNe/REBSk8OF3Fkr2U4mDVO6rt4c2IzdfVQdVsHl5b8SdHt41J+JC0zBuN9iGkCRMxy
JLFqoIoGtekO61Ijb+x0RJL46KSstJR9Lb+VX0fBLK8xO7kBM9jCMfzwjOmc4U9TwCv95D5jy4Bb
11W6BU40/dj2Z2/328VAkxWitFeaOnp4SlLDx7ZpX1iG4yXZHwYlxKYTxbLQZCZvyWyvvH2eWOsm
pZV40e9n4GeJEfPXAEiba0gj/XxGEBnji6YlyEhVxMoG+uTBx+sYr5ZtdgVtq27kXec4tpVLHeoW
2DhmjeRBt0kEyxyVwLsZRN8wIfniZcFd4cXUEwPYEqAg8Gpt35tHyUBRtoS9sZDeB7E2AsjJaprB
AkZq9r4jqDGMraDFywVWwArwtdp7ZKBBjXtrKjvFe9SeLOMGcJ5mmVNueUkpfTTbU0PR1kQorpGw
KE3zyi2hFrJqcWFeW3cxDjWsYzCQm1suqrNzat1Bs5QoHVYF5WbEqknR+xSxa788Q7jrPgStvrTX
JbQbx6pyy1Br7b+NK/8fI4sBGzK8+R4hGa83F5iuFhvarbnYu+K9M1rXbIJncRVs1tj6XMcjsI/C
h6vMu8a4kmbS4uv7bGEnayyCi8hq0C83UwmWaqIobAiN+9ujbNds7PI3UBkKfcJch9m3SUB6VAK0
kEWahBqLBcTaWBNQElja01bDnhAYF7q7x4W5ix1L2xdCk/wjoHTum1IJcXOnmctLYPdNrFhhXv7D
9fjqki6Loyl4X4rDG2zR/JywQyiA+j6G8sBAyubwJkM2wWI9LYML4nV496hZkJqDsT/Ed/gYUdMq
THGci49RGb6wUTwJEr+NxA28kNDkMgddravTN0Xjfv8HWsp57le9R2NPzSpdH5kGey6mVxzaq6PC
UfsHKiLIGFQdTwEuR4T0lndx+NTulg0rLoN5sR3Vk2vdq1dA9BieRqvKq4VDhDwx6rqvBx437sho
Dka3OarHQr+oOvZ8GtVYEAHFkr9GKqwNhZ5HlskUP/w+eGl9XWlq4VBa3kOg28SALP3LjHSDOqiM
MijFfKr4g827D0BfCvKKtOuuuPsUELpScML4O81jR0U0Yg8Gf4JYLKM4Fk1yoXHyj/hiLjl8fFB3
1wz37HZSSXhwuzVbnT+ZoRgMtwPPJLnkNP1t9L85FBFexNgxnWn0BE7Dj2jPvrPFHH/Z0GdXb10e
ggsE5Yea1zM9s3Q5D34xAIZZmLPrF+5goeDIbS8NuGo/8Plxr+Dic/VLXj73S+bEgHUYaBAAUgF7
Gpc6Z4caIw3FoqfhlaPbzrt5bIx9SeW3XEtTBJz/856nROAD7cGyrcRgNfN9QQwyD6DcRehAJ/rv
rsiJYGEzuaAPasry/sts4+OJdGBtnaYBzXhWidlwxTV5eEecLGRlFu9UZXv7X50u7BY1E7+8uZzY
xjsCUC3jDt/r7l/On8Nbg+XRYF/qZ8N+Hki7VC/t04BLVt3lB4pSz0r1+R/IMuRqn+7DBRqINhLK
nnbUbDGvCLfCIbvrhDI7sLh6ycF8MC2oCPxAmk9MCF0yVVE45epw57vj7QueYToe4gIUbNkV4ZOP
a8hC/XbZGV/N/mq/gJStdKaZdH6NUqLLVDYLlppAlk962jh0DjVTbNk7Sb2EBESeH7Dhi4WGIO1q
Rim/X5ijWaOSW7wddo+i3D7yEXuIaC8kEk2Bsex2SfIuuy2lptJNjtQac2vxd6RtDs9kS8FwWNZw
AlkEN9SOF/KF+LH25HxzlpSrpM7jqTzkWTxn8bZular32/GPxdVpmIv4Jt5/uINaL1kYkc9/vIGP
8l9QPZJWAPq10Sg6HT/FEeHb/+GnsV/oI94nUuRXpoL2FGjAXYeGD7uxlCIJVPGmo20JdqH+U8ju
i9MfeprNfgvOLb2mQOd0fBfjH6AcWV5oBXcNDPK0hZZwK6nWK0GWLEkKfidO9hTTVsJLVo7LmUNB
GZUSfXUe2sgMNsZhbSEo6toX3Oa7VXX1fpOXFow5WskMCMXa+uUT1CQ8uaOn0EkLq6LwES9zyiSY
kV6OeEOUyf8cfgbYtqIjGrXY/UW0fqJHwULgGn7ZmozWP38QhMzL9d7lLRNERF3Esz+07PM3CQQm
87YVEwN14ziD+tMrDL4gIGS6qMdo3tBsxn9lTr5ANS8qqBdZYkolDpypgxWwiZa8/RdOJxcate3W
76w6RPYsDy5kPBr/cvKyJdxhGC5QCNbiBsAtgW0L/jWX9XtdI3WvK3fE6/4eCVPlUBtlJ+toHkYZ
qmVmeZSiiF2uJZE+HdhGVoIvsmWRTSghDojo6YzxNJ7wprqtwv2TRC7sycshSpr7kYAkfuIDfYVg
1Rs0bJA3xzwIt2oCdLk8n7jbfkft1GX5oWagg8V/LJo5BMWNKPB9+fKB9Q6tGDz064oK3Zy1Gx7T
49hgJAuxQa/8XVhB6MNe41u5qOM/OqMCzbk5AcQUj8Xb5A7hsi+13wvg4b5hRi4SNbPqqohfeSeD
3S0tcU0xxlw1JZVywYK8I0/E7tzPLN4TLU3AxG75IfBExEY0fWbNJ6FQi9AfzssIodAyG0O5cgqP
AgeCbX0fXhG2zy7pYy+XaGav526f0Xly3NT2upr/hgto782fASP3fRg8cQ763d8xty1F5KOoBXJk
cBxHjlyni8QGjmx55Q/Ngojv0PaHMfoAu1iU/KzFTPA2ax79GTYwbxbCynAkS64IUxtnr8jGXu+3
9fC9bSzwM9Bhmh2q/CabCNs9VHkGPsP9PAPUOjeBuLiUlwnsT4/Knf6bNdl+KXeMlhYDo1HRj3yo
3Wfr6Y+2bAn1yPklk7hIfCY8hqiY91Gq6GtoTTJOvZqVVmAueUbR4oEzIKZh41iOvTuszHhAvXI8
QOSJsVK8IQvV/vzOKXka+zsVIjepDd/hXoESZPQAcEEjpkCl6ST82+k4ewFfPBV309a2kLKSsHob
QEFM/CpkPUSPpo+jjMkn9a23xIArseRUCvqB+KUnMXXWFCtZgZWt8eU0vIX3CAyfIt00Jga3lA+V
qI0EFxrij2EgzerAI0rOZhrIBrikmCdizp96kyWnrkQiXGROYRxkkb+L/XlyY96gNvBLD9bS3YyH
r5SMab4uKRjtjGLrE/c1ZfXa/KbTEBQSjMsWJ+FRMpTLDpkClbTQHOMYYRtwRbpRHd6GzzNmWAh6
DUCg5jykF5ui8oL2QATXTz9RA10Q45V+Vz0FAFFEctW3Tt4F/kZUxH106SOcn27xNx/NJbKiX227
D4nBoqoROXthrIPPy/wtfjtlOLGX2N8UmStYBnuhZjfOsMA9ma5mmlt2apTIH8Lu68MqMXKE8bSp
euSqwhjyTRjdIaj2k9+i2UuSuG+j0JOW23e8d/XSxlL8E4L9PWXHP3rccbnVeThaE1+xi3ntxhxk
vq2LsaoqQQaq9MjzR/zYbatx+aGgU5vguGVkYdOFg+VuhChD80X2ef1A+bK8IPYdu0YrshE9sM8i
g8r7WhHdMfhRGxblhmDXh0bNMFYt7OwND8PzQYZrhleupinKfUv6IspMxyScWtUehF1AND56T6jg
7+kx7fNnza4wZIDfq3v18Mwd5h3qzFm7KDDQexF2jVK+31jUwHkksNLybHSV9XA7atifKkAeHtnj
h8jbCQdJVVkWho6+KPfV/h1+L/Es8LhDoPa+ZKwinyle2d4RnobBp4V5WT39yBBMN2OJTaHWAu7d
/PtFIx4FmG6BKOLSRDcjgnur1sc9jRUICzxowBgn9Y+hcpeItW4f8VgsnVXSQ7jyRn/bSZSmWOXe
ij2I9zoaDeREF9gIYZ2l27Hg9/5bO8tnjVLjj7mudmlEvd/KwI95esQWQVB6tf8QioL7VPYpCnyf
UX0VX4eqxf4kxJKoSaycIfWB7c2Ph4UzAZI1PZU/14QIxVfciRVCqKWU65wtuUSqCJlzR4Djgp6d
OYjDzYcGXqxhDibhb64PH6Q1Srufenwq37ypYHQKzBENmX0xdDCNKHj+41xTd8Atcd4QFvQbQCdy
9mYnkJRzoXfKfQWZFVppM54Gi0wPzG9J/wlaiZXDxLvi/T/TfeUqPdhUSu580kEyRre3Sho9Mnys
xg+djFd3fkhvtUNRXAZDkgEPYOPaOU6KduoRX2nqLXOtV/J97NJMikMhxds+LFIxbOoZCrgf9b5C
7zF9Qh/2xN5LRKuIv22TfTsQst6TOzKk5qN4EGRCcus0RdcoyAbbGV9ZJtoADW9U62ppnR8K56aw
5Al1kB4AfBhbLYmvLO0X7yD3w26HbgMVwj2D3NL2aZwiunKrszfIH4Lcr1opAHTHuWH9B9EdINdl
DB4r9tdDIq9rjT5Xl4ZQRV0rLA+Cc3lTBo1xO3YbySr9DY/Y2XI+8GmhFiKSq/Jdj0+BbvQjYH5T
KOx2DjKvjoREZZMJxf3eyBtHAn8+wS2c3fSacSQjOQ/k9gHD9wdlLAJuplMnTd0W50MlczcIOrGt
/oaSVNFfB9PglGprXSKtyi7HeeCqu/vXESPXcwA6jO7+ESrnneF54E0eIv3vFME/A67dTqSmDbrw
RjPiJCgscQ2F08fU5qpQrUp3TkAp274mr0Pf1JLKKos2Z3KdDhCZSyHJtgFIh+AJcak1XN8hmxTk
GWkOGqoLAoLSbSab485NUE+QdIZ5AcIfPIYEUuBoMIYKPTxifP9xHaJ1WoX7UsPDN2Q1sQ7QgXg4
hK2UuBsF1t6oAS3IA8+aElBtc3NnyA5NmzG4NwGIeyViJrrLlmGqA/eW2QsM2sRcjWWF0CxNloZ6
eCq7rltwj92ROT8rAm8tSHqu1zqwzd7c/0IHNFcvghL00O2AOTByiXvci+ZAmRO9pM8gC4NodGej
5C0/vSXcs7ghpSPZCFAUr0mCVHYtbqxAzEUszTd61qdW1S7rZjdMnFmXgyAVUFahJEwVppsabOwB
SSIoDbhonbIQzILvgLF46Wp1zFNHRXdbbgNzo+r30c0PVRwlMrg2GspfNx6untLDQCarawWpIuXK
fNS6wK3Xy2VsLp/q3JBtrtN9S8wzgAso13JurZ+8UjgksQ/1Yhf0dqKSxNYdMafWxWdVyAnRICiv
KZfS6mLFKP0Y/dzR3ToUzFnNGB+lk4wrt7chySRONLZj7gq4nea05EXGFRF72miHItNLIKUoUg2R
zn7hEPKyCCFbOmAphFrh1BOOcREib8Qg3RqN/tNISjmKPnQvpROJAN+6HX0D2Mwa0OCYwlKPn9ot
hElc00IGWv6NypMVm1X+5BnqaWV//OwE7XMHcPxD23AVYSL6yfLIO8mLugAJv4lCgZ/Cik/LF9jS
SMaVDhV4znG440lMxUnnk2X/kpXU7pey4pVRNF63wXYcsXk4Qe7kM1HMwJYNC84wNukSsaDsU4RM
qFTYfYWVThoMHouz1d4n9OoamBQCsBxlfewS5olT64xsL1KiEq3qJkpd7Hjx9FvTLnEVuirB1zp5
kc+1F6eiH8SkB65MECft3tbx2GbWHHZDvfa6And1QicyFOjXhtd2xqciisDh2p/bVF/xE70rYWII
JR3la8LBCKWUpAsbmXnRWqtIAFskrUyWC38F1aOeKtS35aKMmyI83T6oalnWvYt1HmzN7Sii/qCj
LX3Z2h70BLpA2GhBRcSfa147YJT+NxyMzDipsFMbgOAwU9EA6xF2KTaMf74pl9nr9AGD5DC0T34W
LlLIg3NZKMNqqk2vJORiKq0Mh7Pjz436/UhGX6ahoaP1kBSdRPyuO4zLjFEm9WP4wmsWLlqR94ZE
nzNsjaupEBGSgQfEO4qzhIv4sVdbIbDMjFPt/Vy9oxr44RQ8OWqjMpAU7zCKc6AV58c5Cdc36NWO
dScbZ+UtN3XlDygKAOEhO+yizb+0kMc99DRMI+wnbElweOm4kmVJn8dkdbtF4sckK4lTjiR+eFGX
5bOUaNOwfVLN2S2DdoxKxgtB9t34yHe8m9ikfOHkdfDvK/9WLWzR0mBL3mvw3vgW3CnbhKB2k94P
8HM0gzO77p7RdO2oaiUVDZSUmK6F4gedyV5Lr0LilgR4WCBpg2vlxQz8fkKO3UeBn1SDis10IT8f
YwC785BvY0e3yyUl/C6lZusdPAfCzuhaxpucC121eWD7kZyrp8M1hEWcvxEyOPocrN3IlseoTkun
Fkrta5Ywi/UyIYNNIVvEIxlGW4Pjk1yOvE/03DoMKstpCAA0cX5DUzk1zGcwiAHRRBhj2LjbPtcV
RJMMs5u2YtwkekHp+sGRfhAE2xFAPHr4t6jiNqY2NvE7tq6BADLa0PbUwIpEVKMLZPkKRzA3yxOE
MyUdAxfwA3oxcRZdHO4Q05DvB63J0lOKs6Hzb0O1u7rH/udk+p6OqrlGV29AAGW/3lVVfXhcqd8w
9A6yJ6xcCWj+28YcL2MxiJv4E59y+5ueqV1RqGIlIJG1HEd+5L26OiNSRfniyvqLYpjE/tEAaRgf
P6XqXgWN9qzCxuyjiyPpsga5iSpkpmR3nw/lDi7nN6bdFVYGtV8tfmhqR3bIk6szIlYCsE2rVCiO
LgIAiV73tfCgyHA5SdrFd+CZeJEhprQH7BkfCmyUifPJoIIS+P6AYJlRHK0U50s4shFqYb8TeWDn
HFimwb5ZEuc3HH5a+3/djIsdbtAMD13wFkvgX6IFvqC+oKE1xBBwWnzfAcETlLf4crjpzsM0vvpY
N3RF62JWYarP2yn+2s9Yst7VdnLGmQFbHzsDN5TaTwGlQju4fuZglFRNGT3lYCn98WZRRhEaQ+ji
+JrwOxk22XT0XKkGNTLBx4bJFXEPPkyjnkVzOzGPZfkHX/2XN7lqLDt+hjaJ96DYcy1use7oJIho
2AZFpwPESsmL9Jj0OSj2GF7ZA3a/mepXokf+gYrQPE9+GgQWXGYxx+U/FgLpj1cXGgsEn3VyPKwe
ozdU7/DUnaw7D2Yd7zd1mKgrmufQsnBVvql5Mdbp2Mi4dUGosmRp/EHWXq2acianHeuldlnccZOB
re9To7t2yGxBVCvSOVCLFXFOut+LvlFTCZzH/qsJc5KKtPCVmXdPkhlB23Vy7Jh4zyktZWwB+4g1
11ZcUY8Lru9/+r/V674AJMihbJCy5D4bEjQWaW/V/vRJZ+5imCikryiPZsNDtCoag91sKtCilpOy
wsJEjmvHv890cSkBoXgbHj/bl58i2zfOVGWCLY7ct1m1RWMiOUDgCbYqghTLe77ZaN/QxpUdXuos
79AyL9SmXa1Wnsl1tkPfgEGmudDoN/S7ihS17wioWBsqGmpLe0NWyMv+3bcbcjCsu+prvBPPybNd
yZtjvFFL5yZsR/n8WLWzT34WfH1hk+NYWIiieKpr0ovXor5iFnt7fg0C/c0TmKi3uWXWOZr5g3E1
qOcgeBWpLwf2r3FYWdIHs/o9g3tJCdpo+iSOfrSVZNgw0HG+6AHIXaTf84f6S1iAkgpiSmwZT44v
STI0BnecRAVFvjkQeFrfgnNC5ke8cwe6f9Bpxkm4MOKTKU+zHCa09Br5L8Ck9X+mfK6Axaeuta9v
790eI2GD8LSTFHgH9jC+bG9zIEvu2sBzmFhYj5VjqrzgnK5SzGeqwFI7qhMoXhTosA5YU/m53JDH
ZjG98tdyinFahMe6cgzStwdLbhrhAdCi+62ELCii2uCFnWkHgOV8K1UfsbAAQdCYX7o1IFEYm2ZR
T/ZZUMBNz0F/gva2AamWblYUwU95E2jSi57a7G3y0INYorvLE0H9vZQqtf4DWiyMRJRnGepHar3m
QltDDHaR9xSApUE+bB56P+ylZ0bxkv1uH4rSh46PMEXrUy1Vn+CBThu/Kl4+5Gk/MRHrHSMbGtYz
BXSHt16eQZcds9HrIjzaDDDGSeEgJVfaPhi/y6swDKzPRiXUwA8MwANEVvHnw0sg0tcF+KWGJUy5
+BYxcoQVuiZHYbNi8d+uh5NloPoxCzfJjim2EUhouxgo7bJLt7JgfxNGCMgShiD4/PDwwgQjaHDP
GAnVgKw9a9oMmia7Hhq4IyoX9MBwWX96BXvVpumjMvzSIpQdXUz6PBWToGDE366qumEhsZ4VVftM
xVslrlSFag5kBhzo+vhbzainnHPNtdP2Br+IrXc7qxcAuajDE+gMtDEojvAqtjf8BJ0tNroxZvBK
icOJ5lJ1IUd1YOdKrNPG8lEBc7J/4Pkudwa1O9vIAHTg0zH8RJo1+E2mFVLkZzz0Sv0yNRvwT7sY
o2G8cV30pjYYsC5Tf9zPC8SH8OWPI4q1vHplI9ov6mCl7dx6AxZlar8CePF5wFjoxVdavdkNjlKH
FK7knh67dpymWFu9FcIzWrbjuNfQj72Pq2BZOOGRZiF8yJ8k0phOdjpyCl7E41P7whMggYnhnVRX
Uh74JAUeo9N8n5SEygy/LfDPj2+FGO2wPi5XpUbR80GWhSb94+RCvwyNp37ypiv9I/7riWzdDPco
HHV+o9mNVjBJ+q6qLW96JM3lpAcuLx60BTtulGh6tgjOy73MaP4zZssL+C2QTCmV49CEpB3WGh+Z
4k6pAwVveQ6CfYM4b4ythB6xGBfdHZniQEbwOFaLGRoakNevFizDXsFiug5Nn4iMgyTLueFauest
2140/SLd1LjmbcJ2XsZfCcXFlmdNmIGm4vNWXAzM2CgiWLQbPPdujab82moV16Uut248o7mUb9c+
ZsrWgUE+YA6Qf64ic3v6Nvb1jXkH10UP0mhVh88Jx3wQ5UW7qGRuZZdVwNN2NK4rB/SSOUYucXB6
sJjEkRMySGyrqXLjiurnOY50NFVugPa1+RulRiRVeIBhy9eDYVs4Bf+saghdIINiKQ0v+g7ulITs
p3+OqOqimYe8nlQzeWUAryky8i19NmiKp5PgzIDHtkWlh/fUtvlo3T33JHtRzq6Aklh0MzQmOcPF
6PfAxWSR08cAPO7/hrarWYM7abF74bge2scY14L4gh5pK53BdhnB7ToatsHexRojK1fHHqcCGDdw
fTWb6SCPBVajYGP/Dyy1s1EUTeCQ/jgUMgZlR9xeUimRJCWdJd5TaC4YpSX3EH9ved/bk84W6Y+/
y2QoCiefCp15KOjWvC2aTkaiNTM4fLiI8MSz6yAEUOZMKc4VdtuwCR5j7Ts8sZCmDLiZyrOFhaw7
8or1GyWyGavZLxHVthE4Rxjs3ouZjVLlVQOtdCJUSb1P4fFWVF+RmeXpYxljkQUHkhV6DWlTtS2J
0OX8TvyUGs7voacd7WlTM2qs22YLsIWj6URee1INppdAesIO5EOWDPQjzUK2VYZYOK0sKLOQGGck
CfdQ5hybOAMeXAp3lk5WvTOw7mztvpo7Jpikr3PmFyZrxS5iaoCYQg8c7D+G6QrhXCf0BQmbScWM
YT3SQvlK3xTU/Z9sv33KFAGQ95nKU8PjmvHah8u/NgkT4E/zzhXnB/c7Ndwzglgu+4rigXVF2/jP
yRGjjBtra5T0qiW0vYwoO9//8apDGsahRo2RArz2YngvFPNNCT7nF1HjUR9WeCcwtEbXNOrpuoyO
Ya1hcmy/J5t1CC1O+E5zyp/s4tRjvB8608QtO1SyH50g8jhFhUIs+WZG4AU8BQOtIghycVWaeF1q
CDh0tgv8hEtOYgTjOMQTntMEvi5LV7/eLwpmqgpxFVdb8dSnRu8KzDxt1QDqO6Lzc9OEuGeinSGG
I3jH/KLISfsyj0rFIooKTGpfdyYI5xH0YMdYQC/1XI0EL8vRbaFgh0a4r775W3h9A1iv3MArzhto
BzK6ceoLaDrVATO56OuHIV3atwIe9zsFmDVKUZX9YDEadIh3iN4RzNvADNfNbjJ3xdtQGJVBeAI7
s/L7zM+MbrC/R31Z1Ml8allwHi3q22naB1i2wEE7NiYZfKej3dN/2lAUk9LJtxZbqcSTvJa9PZIo
uge68+ekM9WRqtDJK8ECRq+cMjfqKC7S2LLsArcHTyVsaLJWiztbQXc+eN4JVFZ7anGDzu18tp70
TSBh9u5QPRpDERYF1ZrKW5ILTd7lGUxi5B2CUYow0nWwrPxHys/tWWB1myVRW0OuRcO+4H2WUFvQ
1viEzLZ5lZkyOk/DTHZMuCpLn0osJaN3T2njwYdnKwXev/XFlzVAg9eG8oU2hLI3yjOzKE6LjbmZ
3vb8zaUuT8MaRs0axJPPFVx/Nnx+/8XNp96yHc1yOLlTLSDp/ltN7zZBvUy11d8DzO2F8IC6AHGO
fA/AeqZjZPrQaNRJYmxbgupfIp4I4hOMfuMHR5urmeImIRYM30kXcfR9jwlrY4szTLsjdY7Lutjd
yoJDrTiyEqxFSFVZsNZ2ATihVYuO+VwmvvDyaY7sRU8YBqWZtQ6NWLuaGWMP80iA48HxzAEiXWcz
JuqPbIuLrLnbq+X4aaQoKP7vNJz6Rj7yitB+vz6iWE2wKWA6xUcJ3G3b+RZeCItDaT9nqDoh2c31
pQw7kg84pIwjPyawFPBarIoWbE6zhjl9Nc3aNIi870TrfM+flW87hsw1MDMo4MiOdESxggC6+0wF
QYUng43DbAAj3RqORapA5P3MG16iLK6bR04v4PKoJSxIrjLAelKa+US/pUZ9TGyMlWdJ3/eLgjDT
kCP/A9lB0YfZbXhAWWOnxSk667eUkU7J+33ieirKhToOht6+BNeUvG6eee9cs2aafMs7ScaRqexc
hHfK3q3CaEfhIYw2k56+byIQ8/fGjO7Rs+8YZ/WlGVAaLbDTgeRClNrQyCGCKIxfCYfUY4nZtnu6
1RZh7K8vrN9iGYVI34Fl/SRZZfTl1ytdzXCqjXjzmwz0VV8VauqMn1VwxnkapLWI5hxymDOZonZj
xNTeuwIqVRC9rOFDjq7PL2HRTkaWMiQPpQC7YJxq4MxI/ko1SprLM1JiVePG4sv5SuR4ADu5jXGy
38QtvNMAvd8v+Lk7qMfMJW665AwuQmSbQP64CV3RJ3Mef98rX2LXcHnJ5BadhPqfT8ywr1VoXm/q
J1QXUOGtsOsuSs9QvnhYmD+C+TgLw4HdOlzhSkfdnVMV9WAJmmEHpooCUp7V+/Hc0QzpAcpaWKe5
5HXHz1RfM/03yNowYJa9dHziTCnprCse1C3IRJj4jhw4R6tLQeTIKZoXyyNwPCfp1EmEr9BWmD5R
4jV4aIMtgOHL6zUwZEz3/wCAj8Ne1jBC+lds9hEyfAxJjjb5Md36sp27U+gAWG0MrncxR0L+17ae
V9JBlOgRz3bEnbcFvmAYvDvvR2kEPG8gBccDQfPKVo5NrLc5ZRomBupI7fw2BTJ/Kw1GVuZkI9uz
VpXlarqBTlN++OhvIcyt61Tvsd4wPSX82uG4vk1P8+eBjNXkf7iaSgmNVq4Pob5cGDDJ2P/rPpfV
1TAjlW7RpYp1/udWQtVf1EC4g08VLWeWtwgBewHUbdrKWgDNkgbeg5HQYnDHEG8tbAj5Zd5UwTfP
H3nooT1QsmgaDANQlS2/IKKej03E7vH/2JMbVbqGzb0VVGGuQg2MeF46NSb7Fn55xZg7D9AYbiK1
1ep+hZxC896on7FUX9BQm9cU0M1Qir46Y1dh6wNDKGUvsfmPoLRxigUesDyewIHD8gZv8IaDj4uC
B+KeVTQz7DlwTpsgxYN05AjiZ57yOmyvamvQIwYexyumR0Ul4qnPedmjgzjXId5HAMLvX2aIk2xU
vdN2s01douoD0td1z+tHvd69VusYaOyqMIlPvKIgpq8ByvzaIRi6E6TrcEy1SWl4wUjbVwVjX272
XjdRYHD+Wdfbuv4mUsLBESi47h0fhwTLOZcOpvVb7j8n725lAGJ9cJ9ez1eJmXPHGQ8BlySmFRIk
pXaR3M5UkdTzwzB9XtkAitIQiXhk9kFNfDJd311g2KzCFYvctiCrnrkPg3EJ4Ehstt/Cxm82NMY3
XmRG5sZLJaDwXigOklnhJDSZ7U3Fvf3Yd0egicmom3X/dnGm3f3j7I5+Aea4A2EqoGynmf0IXqpO
/36Y/fEmgNBOibJq93h+0Fl3SVYzqUzUFWRkphrnGrDiVT7uGR7L38EVGDhUcGUMzUGrY2YBXo4w
uD+FDqoRpmV50t/oZdORM11LZ+8kYEqKMUD4O7DuPnpoLwPSemPHHe+sOVqFUs+pr3ciXVnOKRQI
knQ1szEPXmiLgmlM+hlZv1Gzallg7CZemhmUZhUi7OXvRFFhgKno31VYdQrlTPn8haN8wpv5d5aH
oT4p8KKl944+9MiacDMnP1gccAdTIaJrzUm/LGw8NyLcUy6XIy3TPrtOVBhryHrf2juqmc5yB0kK
tzF6EVkyFttofTx1sjp1YHB61p/hgrRz+IR9BfoD8YNChoZg+HaWQ5wOedn2dEGWj6cJdd/vz7Q1
UqTNmnbmfrZOZZx3pAyIJx9i/3RRzWDhlV8aN9xVPMZBoeYJq5+8e3ezKZZFZoX0RfgGB3fC0KxT
Q4mcjHlgnB09s56Jw/PFg4BouBUIyjMKCdidcUQeZ70lzI9yUe7i4iEoCthYGI6kGSqWjBA5hMAI
wVLXnDFSc0OJ3lq6vDaqIempwG8Fc1mOFQCkX+8giwoFqmCvaooaJ4DlYYUKqjiZc+2uwuDD8E0z
k9CGhKA5WFUJgmcgWOTMpATHvAwpbO9znziDW3a04e8q0OARsTG/sVvmHZJe2ObHng2gCdN/g1PE
fBrThMaZE+9hXL3IrDDg7Vg/J2C3sPcPb0gZCBr8jCABH2OH5FFUntPKEmR4Sf9KBuQqwVLP+XM8
oHwHzjmbWaWZmy8crDhGbGZ4jNFF/DGEzc8Nko00H3VXHNbskrFftk+FRuM50UD6VYwh3nSrT8xm
sjyYdmWwbPv4acNiZ9KEl9X+ccXSvJNlAuGBRL3k26bgURviujGd+PSVY0k2tLKoem7XqL6f7sK4
2zdqUiqBFPf8Y5pQ+Jcedsnf4MK0w5bK5OiCtksmm3DftZwyYUB8C51zOU/IOVic2NH9P8o6ANdj
XMAed4IU/tUefZP1e1fVEx/jRuVvU9P4OtxKhN3JIJmrO/eEWnrsTIzhoRWSKxMz6OXXymhg3fZX
+2Jvq8SDhxk4DzHBNADtFWQLHv+/bkHoGP5Sh2VAd7aDxUhrFdM6xecFWpxPQn+0M61dPAz4aNtd
hlSUCg3G66KGEWOmzphTjmpEL9XBZ5XZQTUmvXMOaR1OVZgpZa04k415Gsk8qqtxMLx8pO6kBB1k
CTuXLpw1p2GbswnETw7FD1ndafE+iTFYsSNhBquvfJCiC+Vh/Z/qCnvxdzhOohZjJp5HtdNPlf+N
LlZAp1TxF+SeGbHeWld5k/u/J8US/pO+JoReI3kv5CYGWMl9vOiw+VqDAZ8IiKmJyw3NUco0PTjF
PM2oxIT8zJczcr2MBGKhy7uaelCJaU7ZzEh1w4ujs7XZvZaUJ2x1fInsxag8a2kAh5KcFenRc1v+
H8IyEtOMeVnLylMhfGYfhN/qFikfp875XGUL7bgplnfodTa1Qn06Xx+Lu8HgIMyeo02uedzkD4g1
xmE78IdBLeYzrneam5nV2+HdOEXrbxyo+Wo3cYyIajZwlN1WQOyCV6KgNSoGuzkus5QhLOJ36Mjw
2Se7EKk6W1mHPInL7gOK30HNetcIIaiJdGdPdyrTEUzzS2IgICywlVXmxW6soHxRj/+eW/1dLKqv
0uQeEb6eeB0xRVtNtVt6t/4VL/bDvWvcxQYtfiz9hGPoqC8HkRu/LUGTialTYN0UKS9FdIhTSc8v
0oorDXQmTHerufhkStGyZ3rHmEkOngu7jZTj4aYX3XB2uJDkpfIYSWNRAc1FuJJXCKG7GSbrBcBX
TieifC4j+sfgN+8deqSPt8AnwiXEJmKG/gn5gvrcbVKXOeL47qN1wGY3mpfL7V1dzNgd4Flkb7AI
TwMzC51hHhG30vCMuyJNXEQc5Rz1owrG9bmbYpgtRI0qH2cXe0Yjz29PtDzPy4n6DI/NrDaY9QBW
KClA8GEZ85S26JRsi1sFGbbI++Z4QXzszVc3IXMxQl89oHM8IZIgGXPeR6r7JNhamwZpnwWK2KtI
KB5GvoFU1lfB5xDyjlIJ1FGp84/y+xGFJE/Bu70Oced/1i4S5TNnKNoS9IH3u/Mc3DxgAHaFyNey
Di3j2RuHkcN6EGRAv+UGOIwYf80wR68+1yjyzXpk7Bs6/5rPv3vIVuPo6EGKBr4Qia7Y1zF0HZ0R
Pu5u8VQR287AUSsspR6lH4+TYmH1TZvhVe7gMeDY+3nPa5TLxCJC9YsrcH71NQ/IL3M+ThnlSt9G
4VxOHDOz11uY1ywBJj4eOVM/xv/lHtHVRjNmmKYV3L3tjh4GNRMYuxdTFWXfen+g4Z9Pw+U5GGAj
6JHnsxCHMCPPzqUBVC6qse7B2c00DaD/rw7j3dqOglAY9k0eJuC7DyVZ72qRSj2sBJVxUXFv7g1n
WLyIKvd0K19tkB/ioHLpRMUWy1DyEkLsKDDiIKFE+MsIpGtLdRaEnlwcwSkZhs+DIeHTIbfS+g4X
mhCsXG0NRJU9wwb9obMuINNQhFpgtiDifbkE4Vl/c512wJbqYuCVvezK7/zK+UCeS+IT6Ao27CUh
xPQ4tGPhP/cClS7GyJMyh8l3SbjKwQXygYPjSp/uHxesufR+EmD1S1JHdznIhjPvkJU0XMsXX9bz
HW/w5mqQ7IPnPicUQrO2lZeQaFTvds4YDzb/oU2EkPFrCzpycXjXRpuofbwjUJio5D1l8JAvL1LM
g3cPZdow+D2OucplBhJQhPhs2LGKbUK0WQMy5WYZYX4LNmfmwYeKRKUbaWlWXzyl6HxA5xG4Fspc
Kpd+xem1DACgz47mDaWnMgdLS27ROIahcf13oUOmT73jmP09GAUDq24h5l5Pg9uj9clduO1aYo8q
kQHdbC4UfXcepLDlG+XKb/lYycC9Gt/53c5zsV9hs3yPN78R4xW7mQYWm8neEbsbpAzOjNi4jIbN
SFQprICvIj95j0pjpFFBU9GaeNXTV0cbhCDPQSf33zanX0GMeS4S2BzB2bZ2WxBkYCFLGPuNR75e
21Cg6dCaOacxdZC85B+5d8aQpC1NHBcJicEjtPlDpBFBUXZMcQ/B9hVT0J7+709A5XBtIoH+wcDE
WQwGCjoMm+9LiRqEY25ekQgVwBabSyPbvpFXgdy/PLc2n++RtmpYqcE/7CgPjN3JOwu8nfMwSZWw
+SE5qTspdjmahYYmIJ5dvGo0wBTALnqbx84TmY+kFbJvIWtsQZ3JtZ6ix18fgTeWIN8btf9f9K0Z
/g13sr03kzA/Npt54te7hnmm5dWpFmIo61LXecYg6devmtJ7JmvIk1kfsTq7t2SlyXEfg3tS2y6N
6C59hutpXCl/oJHN9XhpxKieGzmd3kinqijKmNT1/UeIOrlOterqr1ld0KgVYzftGOVcfDnzbC+v
B7rO2EkgElekvBZzCHZpcWM/doFs5bl8ihys5CxNXzNqBneCLG1mjPH2bTD7l8GENrw7VXJWx8Mh
IOOiiJ4OoMjGIKAOo02Im0zcSSo4m17hrR84J6oHAZMRvTU54fPEiWeJOT3prW98wX3sp96rfrOs
R/VrU7FMQpPlgI/+O5ZB9KwhqeXO4/EjQz2mQcWMoD+7u1LvIV95itBVMt8Dcejs7nTkq4UxExRY
0iPFqBTsKSZwW9u1nQ87NOBTHcSIWPYGE/5iihTbdD90WIXyxKw6jIwg0965rDeqMAgJGYo5UaNv
9lCoaTKWSuO998Sit1UEt5Fpn4t4MB5n0CLkd5XGAIvdVI+s2dC3LqPHsOBLzNgMLhu3G8JPzQTx
M3g95TTzPp4DKEM3vDl3zGqwqO0iTRxTMeHQmz/Sf77nmRO5m+x/mdqLIb4otr5DpaAp73lYGWxR
24bmKbOMY491Hl3hCNMnMbdFF74iGAYmk337fraphQOw2jz21EVlRDB0Jf6zeV37MD5uRFhePUYx
pbmB8QLVoyg/qmzHxYxb0vR3guVBcxKrxVUIAlp58qs2C4deSbEgWuQsHyNcyeNp03ZiLS13JgF8
ElKUOfNvhKNGLGzBkgSGfeY+TozOnibvl07idqQhQ2M781FcDilqv5pmiSBEkCAyp3J+0s+waDah
WcL7VzRazvG7hQgEjMyE5hjygrOnuTSXhXLXTa+RVQw3cDzR18OAIxrodmbtEJa51WsG6nzXDk6/
4um79JQbOqqAhMeAey7JDCTcWJAxuq04XxsejHzXWesgWTLCCcKBOp9IUe+ZxZ+CvI0E4kMT1jyA
EdCryGwxO9Bq3xvVKEwWq7L93kx4d4FZKhq1PzrN80nBslu66zvR/T/CccTBWgs1izykKBtIoEIF
ZLhiOzSpRehVn33/kJrqiKPZE+c4cm5KFrraSi0f7V5Z6QQckbAc0dD7LJ6nuGaWGx6Ob1Z7IIQO
4sgds+gV2kefM65P2fgEwzh5lL4LD3UvpX89lUbJLUBqiQ0rf955gov80tjZujdsGBRbNPOiXuAh
vS3okfgArT8RLRK3lbZ6DIqFXqAiJdNMTrGcDwOA6WwP/Yj/xCMOeVk667rNMvvhPVGCyEk1i2DS
dI+AEwqiLhIrpDSPEf16bbodj7P+w6DqyhfiDn0XZ9HsTMMV2YlFqm8zvQfujzV1/+l7ehsT00Dl
FeKNuH5tVE6zL2zD3oJuKBxZZs8nMI2pQzfyMvPj4v5exXa9r9dqp5RRkKKehyT0b1jcUiSTOjhB
tN6QWb0UJ5D618UhVNcngARW4lSKXwCsQT7OaUi6RmQgbJsLm5StPIeVpmoep30krfTka2pmZr1Y
eyn92ozVrFI3L+vY9Jv3S1k+TkAR/LiUNGWySWZVThVFf9Ljk3gXa8NNBZ8ji9rZp1Ga0zl0PwZK
w5nOgaE8LDlcTlSERTMgXKGdhFvzD6OfewNR1o3IhPWC0gF76QtxVGD9gTdc8MRfmyNB8kGycvUO
mAPPaX6p158KCPYX/bUlElVETtm8Zsb/7uxWhujfLQOvMejOve/NzF1U96MS1PycZVAF1LLG0Xyv
eoi3J32iOBI+YV2yow2lVoQrRwQ06+XQJUucQhU3Tm7GiA61kEdltViljtXUjPXHLMvs1Oktr10s
j0jLsyNVlRpquL8pN/q8lsR+s9tEN7RYdpTLHZh5TSzioZFBsCKQF+UzqcUJ/oy8oiQSPlXLWXsI
UvEZlqfi6rJv6tRs21G4d8wQgUpQohNp3XUth9evLSzlX/01Yhm6TuXuM1/l2vaOQrh+rPt/VMle
bUQSenMUEXeBmbVk3Zi5CNBCuSSx5F3I8jZE++0/IGEHXLCO7aQiQym04M9PHrSns/05WvPY5qt8
dHpUnE5nlZtMLKaATtbTu2dcR4IqtHo49juV5DNmbG3q3LbtaXzCoMrrALmEr0sRIVRy3cc4vulO
vzk6w4ZRa2g1ORs71ALVFdeV4ijM5QW7xYDsedO1N/yQi5x628hvqBLm6sk8ZkpC04BD0xkJ+Pin
8RnmZ2Z4UztXB36G4Tu65hrt0o3JTr3CfQuKLj7MI9eM+E/KKhlq2Zekck3UTH/RFGN3/mQD3At3
RLC7tyT/IPn2clQ/pdao+LrI36Rj/r4blSk3nmeOQykVh1x+fF4NXBA/Vq/DF+2msTy3ZMPgpTns
ScJZjP6SgQCyaR9ZfAVjjTmxcoV52mbPP2bGTsEznbd01lV1xv9f8pRbrlCrlg55JlubG2lOGc4d
arzXCgoWzaispMbvQhKZcjyvjnB+eEZUfzxmVczmxVg6AUbLctcHIYQCNTObs9bQc1ElvtoYk3wL
u1D2Fd1ddi+ugNwDgDs4loUmDZJy/fXe/1aZLs5oa+btp2Xx32XFuYGOjzzVuDsJD5yosd8izkns
7/UsnznVzLuflvEHdaXVftvvSwZp4s/IG3DA0ndRuC4r78Y0zG7cYTmn9P0HJv0t7edZm5njZLyF
JG/t6BLIBcSWwL9pNKfnX5o0DN+uzWw20F1FnG+ssEoJKgd2C35lrHUr82qDW8dCFQt3pbuvQHv4
o2zkmj6/B/wx8/na10GtEOkNIWHqsM+Swunxxde/3mpN+idHQYFpHR0Yx64gWIThHPDliwk07RD1
6GX04SbtC9LDiGDLN5L3BfDc6jazXktSDQMQ48Md82JRc8F4VA259BUf5VLwK5LZ9NClQ//hQJpM
MWWkxDrU2auRCGJqyzYU+g90jl6NFI9gS+GRIMx/4fO3ougM+dgxQsRbnzLvIgFbA6KPF4xlE/kc
LHb/HjDcfCDmGSgRALiijrq4ZZq7TxnWD8kv8d/C570A1VZ4tT6bNnjA/NjO9LHoufArjSw1bnqd
wqPrIUQoH9JluwcAjyw4GGHYI7O7W9MiKEFZivZA68jXtGgR7v+9Nf0lnmbUhg29WAIvP9v4dq5I
U9CBCYWQ6PfIovaiHJDpqtOIsB+9+m0cT5uce4/5z5pffkGRF/KRSuJ28hGsj0NQJrM0EvS7pgDi
TCA/c35neroYjJFL3EFgEgSMzWzedyaADCEbepAkJ5aZX7ZKLZtaa1opp7jnJGMtCSRRUUnGitXk
5y5oM3dc5MyLb2OoVGD1WqekfL90bbRoMIyFK0Tl9D3OL1Qy/i0Om+2YHvpO65ajtfw2ov0XXEDz
zIFPXS3UxmjtJidpa0Qv6NZakiJWAwqrYCJen9oAAHng1BdhWTWGGYtq9TGW3drGODQUqvMnYs8S
oeEYsHJU0JPED/GayWl0vz8/u+43OfBeF7HtquT1B9ImTg8ESjTSFHMhNsGsy3JwduAUkcYp2HMR
KqEh/WEwsSADQBgxaEZlw2zi3Xg1zzRuxbdy50GhQ1xhf1XSuHTCU9BH7/AcRDNPvEw9Dn7n4f4H
1wYaPzFCno4rYKNukd85zuGXppHMcToyxJTP81hha3n3orNXY6I+NrUzTP09wvS8rOI5abDjUPEF
ghzSW15zpUzaW2iA9zONae78jrNt9Cp7L5b/tVF1s59tpjeIOoR7iQVLi85PCH9Ishs+N0hFhI2T
a6y0hngaCmWGwvQAT8CYTz4zf/q5plsYYbeKdlD8IAYjXEiQTITowPeC1rRNoQC5NCoVQjyHOwud
58RYBke0jLwVr/pM+BkiGBBalLIBninQk5R+XkSqBikvMnvR8ygkP9cV8Rr/+Uv6gv59cK3TEurm
xaS4UqSOaANB8XVJ+7qQ52YZikF6c3Hw5epx5nRkpQxDui/1wJspMGLg0zGQNiJLEQWq9Ai08qUk
V8UUT6ThqYh8yogFv1qzqzrxH/61VnOmmNl/8ajNwI6+nK1S5S4Llv9raiOJc79HkPmO34lOEnML
GDLUlWEK2yrnaQo1d8X4NzZw2OQyFro5HXfmWZVXUsy2Y4IUNnUEwttLEZC2DKoTXz+AD0c0kjlG
yNmge3Fc4i9kjXS509p+NXigJS5KaT+JJpo8aG+ZDmNpzfcMj/q9Y9M4xxqU+rH/++Ny/fqumVri
+Y7PDW1NXPy2dg+5vyhjtrM8kw8a6HlCtv7kcycei9d1sQ1OaGjTzglHLnsbYje1aJw7dymzO184
sRK6UCsAavsdgbQGAk77QHir2DQVB/N6cBHP3IKtTWlwAJqS/37zFnkkjzu/mWyLPmThO4qsYW37
WltqrGfm9BULEIrpYPmgMcCPVGGMTKFVmStk7o/xpcjM5SY+Qxq8O7Gg1Ws3e9ghH9nL+h5LSe/X
LWmYA3WiJ+YvJez7RlO0lsqhYVoKSTB7TRr06WQZ0gC/JdaFlTZShskpCVLCswnVDMszIV0GhH8L
kcQqs2LvjkXEauYILeO9DOPomlXrbDwV3Y6dkyTKqNz02VNDesoFkyGNwiAwoXSruM4PAf140Jop
SwlUkTQ99rFjZfEe1475pKCiTqcsNAYnQhj2j4HBUYfpCa2PR4vAQjNtnXJMvtRVXzAKpF0TnJw8
D4r6ZbSks3+RA3sboXpWOusW2o4bY9iLzBUWQOR2rn5b83bHYHF8fJUPvg8oIcL9SWR2To5/MjLr
sgai13oRTz70UR7mSAPmVXGHRxFzQO9FMmjHhnv4ez02fxdeKYdlojvT4AmH/NPipoAmcZcdJExj
sirtpiR8f7h0ei8bGpljbBavGTrNtWykSKUB3ZqwYMnVeRvwh80fv6lN5LPI0DXSn3srWL5DcPdj
PKgUmBvGDN8lHidE+JP10OnNTjKt55GfYiNeR7Lg2sOrtzREW8DJ50uN8wo91wEpR69H5++hmpg+
5gITT5EOQJjPhrHmIboWMBirvmnrIOGF28R0ocoEd4Q8qw3tShIeoDltydtDWiRnr8gu75tvB90b
/gRpFxa1KtLyAlAohLHOcjSHFMA/kn/bfURLnZARwmTzZp4DNhBbj9xM8LRqRX8VBICNiyMPVS4W
yH3+qdyssN/wUFk/BUjSWsICevRPVYmPzIbsbmYIi/Jb3H3jQAidJ/b6yRL7U3axm9MvLjvB4DiZ
td8zKBAhrDYFBhtiWNJnEzipjRSxy/Vob7Np9WCbQIuouKQJ2xxP8KJO00gvxF/NH9Bd+zpHUZ3m
O4fbTlSWUOhu6p4t3511UqDZEv8LP0RhZdiG1l+RcfyDnAgtT2LSAGp9FQ6GMu567WvsKzBcEkKB
ZhSZkAAnVmqbW3j/PpHtU/hbW/NE496E8CEwxTgar5X3KNm+ggxGWN3BXqQwEKKVuvXAR0/d860J
KdqazABaxlhaYNFDVsDYLzT1d/MPCxSjxJLHeGpLvf73NcWNdPFiDAMJpWBD4tfw49dJ6B0gH4FK
IvEiMmj57L5FRJ+iFJ3kKuWPKDFz8Gu6QY/XJnCWu6rpfTaPImXlrc+oFkZNHqjdfkF7Q8Gtxjga
QE5PfD6ng0TZ49yQVp74FI6sMBixksmpZNw4iJgmG+BqnrIm1dnPSqHEsFLjLkE4h3T5IAp7Fk77
R/+dEneV2WjUdRHKYAGTKofUPyg0BGp0QCTithZCfg5fMFd+V+x0kQCTeFKyU67c8bRU2RnmTB6j
3/+08o195EVauis1piL89KliXFFFB7VaAWPPHCaCxXIBSHXt7GbD1kZfeTG0vzbM3Dlev66rx35Q
0sIH6/MgzX/0ipv39ESIEoGx8ePuqGaIjNCGITql0QYcNui7vYDFTpZFKuLy7/VKleznmlguFtVE
XtUD8qoxgsfJCQSsDFVhKlS/1fcKYDWGXKD93F2onRo2DQa4JVDpCBJLKWxe3bF6etpu1pbZsOxJ
mYWfkeleE7g3XpF3MbQIke4oBmyY5n2Hr0s3tI0AvygOBWBREGcwks4avBt3hUAiQyB45f3k9ho9
vVoImLysw5xscxncqhM+hsFEPoMRA0xRMecDcIPwZOW2BTD7emLdVTNpeHmOxsfsERpv3FATAtqU
GQe436KAGBdk8SpncJuqig9ACUbBmu1pY/jVrB9GaZFfGxche+7Kn78IY/odzy9ZznTC3ggvBdn6
OPhf81BH8t2AyMiUNfNUYeV1mIUy3axSXGEuYqsBXEbGLfdI5M5gCnz3UXccEBopAX4p7Xe7Tqoz
UStMvKokPXfs1izqYMNvFs+8G8hQd1LSDH+HigY7kO41bL/e6TG7344EnROe211NJQP+dF6yhJUC
bDy3lD+1kIZgttYUUpL8tzRtqeOOXjUUWybfvMv9dYWVbqAySnRzSQyhQjsq0lRmQDUgQj8rh0Bc
RqlWY4QSkQL8v9qVzgH4756r1phiaj4TqSSmhVI9TYnSBQY/V3gfi/M2Y23jjQ69eegs8z2TATyd
+bTeqPFJFkO7YUlMxs7XIfdSb65bp1myjVr2p0plOhjBO7O7iADCxgAlmInJs6Lhi0S4nI6/Omft
R8Iuwao72eK89Mn+DamG+l7oOPTtF4rDlubGDt3zOCCWxWN5gacH7hhBFRnCReCQMRqQSdofBI3m
rvB4RI/1u7YJq7kryRTAy/MjQG1YIQoSHCNlrSjLyrD+mM77RZMY8A3Y3sQxnf9asET8m37MPl+a
S9RHkZCiPsuLECTRccp45OME9QhAoa9Q9Iw+6kbfh8/AkgZOhmnjGO1VF+u/Oh/RbgOdYdZIAg6P
g3iymK1Eogwyg6O9KQ0Ho0Q9Zbw63MKxdipnxOtQrPxY8+6AOvXGd1g0mXtczWSywXOqwfJwYDSv
bIkFJUwJXcrcco+3bqOKZdgYNUE59sMN66Fbq82ysa5pHUsT7jKYFk0CBNsfwOQdNR09sZ7DmtBC
Meh/dyaVZoKStFG2jpYeNXK2ICwOpoIpiFioH9c2ZcjyI9RBBg3ZOJPBJqrE9BT+IcizyYWseFZH
nNs1hDeou2zS7zt927vKuTEE/dHdvbstQgrz6lqYzPP7ve6J7fqd5LkxM/73bL7mGnb0f0Tru20x
yyHI96Q7FYMI8W0DD850+ylaV+JNIcKmVaBqjTQwhEovPc3mmWdFtSsf1spAtRvXYoU1q7vQXxa4
QbNTCPb6RTSL2mF6RQLgCZKabMmR1Nk12CdNoltWtAxwi1uxerzsOufdqSO0RI9N/BiAqnPB+xo7
x1ayKH+8qo1MmH0USE4EKJj+UX/m61qXHP/PaPCMr+uNjakLgY43aPc8bHy5GpW9pdZg1W3zNFkM
JZwRL+Cwy4vNsEwrMarSV/kDplHRBhgLzBWWvWCwSj4ad6DBB8SNfMxEMkaGGRap2n6avAAG6bUg
4Jt66FWGd8efPMnX0bfPtNWL1EoyPPVUEY8Uju33obO69ZmWSGaepbnekPH2N90MkPyORdA9pwZ7
6zzlKs8zfxXtySbxrpKBl+NOqnP9cjGEND9JHhWM4y20u3SnFi+VhXL1gOnjmQd7nxBDNbCATF5N
lTGokyEYNHlHPb8pj4a/bDqw4Iqb6cKpW0+2w9zaeP7w9lYpbEk2DIUH08aYV5XAb17IhI5QuzRE
vWbbuMqMOMTGilqklYJeBg/M9xoHRpg/Xtzs0jK9Zp0E8zmhmvg962uVF2qk7kCmq2DQ0XCI06Yk
mdaqcHX0Ei4wXbVjpt0V8ZA6wvLUzCAHJSbphjbICELTY7QQlHBfw32c/BJAu1eHjCd78LhD5v76
hYPzzLjmuZCeiR4srbHiE5+gTs0WzYam/J8w/lkfVzsggLc8eNAChOdtgsWhFLqjueymy0mO5jdp
HlUiKsjVX+/PToHz9Y+N2E8h8JT+RLP3EOpjKZUnTK4XzYBZPOsTRYv2PuPk/ByemEoEebe/gw13
56Baje9AkHSok0/rBU5IXs+3ILu4A5dfjIxYYOjA2sZaKQ0zO2IfmnMerKJyDRZRZbdcr7AsNlD7
iO1YftClF2h78BR+iqCfdwgdEYVSEXaWKn2WztwRBsexW2/cTHZQDkSB54Ai3JNo2kBqMnrK6ndi
qRO+Gj1uglp1MPFQOg5i8c70Qqj4g3/E/ZQh3Vu8uYVWPe0QsBrjtwBsDCi+nIytqObW9PEVd/Xt
spgIFoTkCtqNQRgBxW4JohSznY6cPAG3ZZkSBBHyonsNDoMoYFGzBCjNOIBKM/GcxYCDvDSrdQJV
33nGwTs3KTXrl6MLNX5UaMo40ZdzOp+U9IHUmzFGtaok0+OKScr1ehnifLBeSQH8hmTYxmLxjzag
QIMdFWztJLuxz05Fr4NplPItINjQ/FsVAmrV3nJ6irhnXJ24vgGhnEx6N8Joxki+WaFsF1fdAram
UycUw5qAUwlvEa8X7poB5Vkb8JJZv+dG5mBBTqVyHAQMjdvc8gu+DqMXiQswmI2TeEMpvjccZ0Wr
ufzStwNvC5AlDeqnRdUh9E4keysMDKMW7Cvyt0uX8FL5gEH3lfXtfk/mVVvDD4JFy7GX4TCPZVhO
jjmHXsNQJZkCs+QKeJJWk9Xz6CLYmmxbe9JhlTkBcUgNXe347yMfDq5x3DqpXI+SCIbdRFz3TArG
O/elg/xTXYbjdEOczc8bu7F9cK++XfGEPaHLZukRjTLzNowPpET9W448g8G7Mn+edha62smBpz52
9DPWE3XMNc39ftIMkINlx/iKyJjbqKL2sXopBxWfX7LWCGFH/kIWEkGknbxOHYmga6avRy/fXWXE
70zTJM8nxHf0KHiEgxOJHFZlhKMcQb8BXmCR0+gpmZfL6cHd5v5/VT6cs1kjvVDEAIdYoa5NzAiz
2ReUelf35lQ+B73jXYJz4YWCuqqP0qUuuS0AbnlXjfRzJ/k8BK1vs6lbYaOWs5PTl6J3VKa1kj2M
4arOPEGbE5dISyBximg5yBtbriR2/vWEkWax9LDa+pZE8gqHW8vRYWWQdJ5ULCPf4LG0Cuw+2qIV
bjAlZKy1TEYu06LqP5YE+oK+w38Bilc/m4A6BpdDDM5/6bLLUhllBeQr1OG8KLApRYCoTSXypvlR
x4cN6E+3CoFi2ZtHEOupPILOywdGRk13ybIsVuCMK5QT9DOMdCzOc3hI+6BKK/oizyCJGWl/x03j
sYnbdAaDFfhJNrwA1mBRurcSt8c/b8auVBxahKMZHoXMkTVRhc4fMxMAlcWDB9H1m0VLxevvi1N+
yfhS0klAsYUp6XWHHNSdFzmwGNJWimM447SzwF1+kU1RO4VPxOLGo7s9fDMv42UYmy3u9eRMen4W
FTGBV70o2D3DLJLPLuvKfRMXfv2EWAM8TM4J1dezy8Wk1ONJG9pm9vDscODAqm/TqR0zRfaGxT/R
uOc/TpC+GEoFMW88oorirzeTQVkUYMxvJBz1EqWo3qPY7i4B9cf2zYCwgb4GYvAyWAifE/IeDQvP
vUr6T5cVhpf9sevLy0rT08gPeIR0Zb+auPE9M8TyJBGNsxYQHtwcm54l0fylS9kaITBDvL8WcGIw
iIXB/v0oIkwGzx4SbkSquwIaQuuQCjtyYFE1o8AhyuXWqFWRiDIgb03ojbC/CPZzqucFcSyqZaR6
KvX+KutKw/y5UR2Z2rZzHgLLg+wxRnJpaDw7Vg2wFRmPHmdE7COGsPUnr3Gqxurvy4ivW38HnqQU
8Bd17ajMqKC/2l0LJ/VG6TnBakOU5I/l6AH7Plfy+Mzo/QxLvUPQAXWuAAfM/9zhz8/thJN2lY5h
/xbpFIRfaBkzt0wXxz3BPzxLKny5boCsSIrmp9JqSSIcaeDgrpA1CIL4bHOAzapCd2HMmluARipg
SrjMXi6Bh4Eo90iovYhgFAJuJgQ9FqVSGsBao3L/f70vQbXCrBiKjlJDGVE8uI3+UqzxtzD0UTi+
Y+AO1w79IxMlg37dePrGvuo8xA+PW8yizQZSqfPij+MViU96nYVgsUXVmuN7kBlKdcH2GODsQGhj
/Fwz1ZPyPi4onedFMY3u9OSgtMj31KKN492XcFgo17mLshHXKb67P/ojnfKlJ/PZamB+j+O0JrdG
HARWJXXrMKEHNwrjLdll/plUc5yqRwShjCW+zXfnHRaN6HHQcB7ZB22hW3/Z9MaeFYAOAwFOvD/v
n3hEW1prF3rtGfapCdJ6SOu8NkrZ+28S3CAjVu+2LqwvEHfcBy302vuyao1vzhEvbDk0Sky7tPkI
otcvM0n420K1Ane4FON84f6CK+nyP/AP8/J7dDAGvCjCGo85jrZ7nVIbjc3O59Dm76e7VMsxX9lu
+46PyATzzLcZBFZpYhdtcfDTIKrWfe0SfpkeQK3OnwqlCD7t4trs3DeyxC936bN7JIY3y1/7OeHI
h+3LoJ4LAOiXchvBYj/llj5aJBsGxtPu8OPfz9Ck4R03n5YHJwfAEpTiWrVokhvjLAxumOdOrgDz
a5TtXt3Rzcch/e2jELnlCqr6GqTKY6YnBLwOtJLne68011QHI2mnqkTfXBV5Cdqx70VoQAJ7b89M
FQm/iqpmm9nIto6Hi3hcCs9oJwOHrtYHqEspqjz2l7sAaHJKs3aobMUaPHfnYI8kASBTreGBVk81
ONbBWpMOnwLutbuAwLltAR029y5usVuzGFCgRj7uwyeKUlbp5gt+QRxr+qDt7chGcZ4JvGnOyPOV
smIa38d2MarsJS6dKzuDe+yERBcdFz+pT8XJ+/8h9mmFJLzg5uX42aM4EmMP4etKVa6nkpXsWDy7
atOqZE+/3KeeAWEvp86snX1E5i6kXhlmoHqAnvyowVHOLm6HuNiPjRaWevfPngM+z/2RYFpW8hh8
BcHfY5JHPsCkRZuhubcfaUa0+a/TtTKBAA2y9U35FGZjMp6h0fxe6YziuZoJa7Fo++0nwHM/UxIt
TGXToicpRpgoVd6L0EPXGOIKzO4E4nZOFFm+Uk5vz848yW6ARapPHPCe61Hp7yRTKPBsVHelGsF8
w8dlt961ESHVJTLmi6opa5Pg6X3kt5shJ1Sb0w4ET4IyQXNCSqZnBgFvwGijKOqnMqqv63Y4WoHt
+FK+EkJplKUxOC7G/EezoUTaF1JEer5wBpmEjVw0228lUXj18kw7erysyNbZ6sY7GKnwyZpezwCJ
5PL52IzA11HFUGAuRwD3n1HXhLUYL1Nvkn70k9D1chGlCoWHZcPsp1I5+mRlp73riG+hxJiERsCW
wWL196RaNnwXWSMDqvqIt2YbGmcbH3ayJfjj2e/P7n4bQcNTbvyCgnl4yvPsT+9cJzch3y2hY3GL
LxHnkEwNh++wUrWoNZ/mE2Ra/erciSz2nobgibOwE2OQX+NsEDk/Id9hvZ9HtohsqWwDkSG+CNTZ
IqhLORc3DyibGimhS/0zr0n8k9jV9IpFF+0V+an2wjtli6BJX56pzwc1S/rxNGAwaGipLyR4BVW7
2uYIHiz9aPqty5WRIEARheh+IcaZq30/QXU2TJ2Fs2ltiRwVyaFveNZc2TdQ2cUEjUNErlBPLy69
b0G5rdJ85GNxQb3e65fVNcLemQJ855yJ+pNtxzid1Fnix8yXrHdtXPuI1fY+54j/K8jhzcwuQNEV
qYenyNk/Kw4ZNvZrzGyjLibfMzXFIdl/ZIDeNa3xFncppuJR8ay8hhIL91pvpbemVq/CQXeRUw2O
zi/hXkhCzF6k+3oJtSC3YVqNq8lKOwp9SGlFxz4A+jyugAiSquSPUGWmvIUN4UeF0veQEfj4TG5K
SwJEC4P11vjUx9GYPbSryVBxoR18ysgSa+1RZUMy87zp0hgkTJBrv6QW3Zipyp91DS2Bfdwwra3X
w2o01s9R9lHv7uOEyvsp3QbEvL2bntxq5A6KKBZUx7JgqZpuGdMKz6s2iX5brnZypysWFb2GKQwO
ADIm1721UNWNMBHo+r+F0haEmAnpcG4Jp6nlwWS8zmHsJ1dnYB8H4Mp2m4FhiCoStY5Alg43266E
GmW0HTS56H0HimHCf9FlAW01LEBWaHHDlFm/XuHEj/VerL9FCRUB+5EjnRGCdRY+MAxF1RE9mz9I
rwh9j+JBUzhgImcO/ol6/Uc5dYsoo3FA/E9+vWgAmn1095JZDr+Fo1wdo0UtWrf2bnF+oDPG2dkw
G24QLwo3OfjOv+NyGDuq5SYEH+7Aiog7F8/KDSEbIkPOdvS7PJp0ZP4gRh5lZHQxmSOUPzqJaxcJ
2+868YgLQ+6HxQzHQf42qet2dgFxcXIiHLZlux72cSkPCcO/In6CLoznKxO3KFwxUB85XEEnzjML
LfwLZaYa24kFjDmboiKv7IXMj4MtgkxP7Brhh+qDjJz0s2xL6JsCnYPNpoSTGpIs+toi0ZIG1/DN
SgKQbz3RBUwtl8HpSKWhLJDNHlkQuUmhQpx87KaN9BdcdCvtb2CdTbxPwaVBHq/E6n0knLrL4t4r
wVz50j9aUgWGoJEzhFwHnuicy5skPha7cbdKMxq5G4Ku3ziV5MM0HYzTWzvXSh2KUXMXCwxqpd+k
ZfHkejrPn4+zcNwcvleOaw68M0AgvaEpi+zfjRzKilhi7oXHi/af0vR8HZ8JmPzJlME53b9SGtS9
rneTp2thVLIdeQWQG7gtJ8tdU1KZCnuFZ2LQmjC2dqbk8ujphcIMJI7ouhzjuaBRgDOLpGQfUFiF
2yYKGr2X+0qlp8ckFba0sXYq3hHwJ1g8lPcRUFmJIL1UlAzYNdSSu5Q4eIhIDrcYKgHZ8pxqOj70
H+cy4v/CxoHs0lhA4R8aP1kK5JAMfCd+plPcFeenaKRRIsM6bpakDNi5dsbbxJ/9g9RHfLsJtz5n
l3OyCgvo3mDFv4VQ0xxcHJEDUAnud8q2XBHLsVJmwoV7Mun7Tn2M0n4JdeGTAlwHGh2/mCSimeLS
tC2l6hGP+b/lM7dimqv4AcK3uZwKv0jKjm2EzI7wEsIp9G0+Vvxk6JhGEkMnovopMlYqH5cemKjr
32oYaRgAiPA8WjhQYcUoUayQti6zUUxEmqY3vmIUGoEyH1trM9V19zJNuABqC2tVJlLGBv9+gWOL
hmVlBAALbUxormQhAVk6DzurCsi/VmxA0KxyngRJ7L57DhToFq7nBXvK/3dLw/8j4Rm/Ni3wTgcq
O5656eBEhoZp+WTCLCmBDux/qZiTaJ0joGJ2wjd6VugNvMM5UFLl+LjP3ChZXdXdRXO5xh+1Bkdi
i1Ipz3N8tIT7OTClbMsjRAK3AS8EaV4bt+dKZgTRbyzq9RfSADE7Xy0i2h2vUa4r+nSFLeUuQjeS
1iZcbjzzdEH1vTrrnKuTvLaq7t0C/AK85C3YjAkhgV0dITG85fhKuOqFYAgkIZ9/1yod3tgDXFcD
uHJwNAn1OHtgAfwqVjDjuuFI44WrJEEHStj3tgpMt3XK5Of0CZqUle42KqSuYbHxDQ4Z3frgbbQE
csDCvZR0jhvujfYvPq+jtRoWK3XKOqyoZBa3UTJyN3qXJHW3kbqOXiYxW7XCNv9eQwJqykf+ePMd
D+26Jv3KJAAzQWRBYS5o5E6yHMzIme6d1wPkjJsmdDETkRu+Bubx0oHjan4TZtNpVti28kd0P3fk
E+1ViGuqY6r6qePY2QYyvfk7ZC7tB33YRl7QJhXMMK7iuY/Yl6/vyfOUF2Fzx1Ta2HkyuDnTVP6+
K/39raTnmpRI7o4UD+ke9cDw5AKwNADwIHMMEM+mBWztLjOT1YnwvBERgfpGkx93Vr+wcCwntH2i
mrWK9NkkMhEgw4O794Vp8msVYGDHVQ3REP+j042pPPO61rHz0iQtvzUyO5H+Tjh10uweFlvMRf2u
fjUJ3ZpiNfCstm8DTIQrUlM2IjHbNJI/8a7MwHlhZRQUuFwaFW3/Jqzuf/3yZNt3Rciy0e4pmuS2
g4La5oDYNwSZL+hCaYRC53lMWz1tZXxEI0JJnbKqyGwqU3S1JsmnE6p8M4eAuU2ZbMIWHVRZhOqZ
LZuZ6+Yv+ZaLF65TLSUvXKwok/3JvBR8QJH0NKvxucEKq+n6q/eBUmI6Lz7L0mEWhVencUjwSwS4
0WCnDRm6o8AJHLhiDUxvF66zHU1fU8Nw+3L1qVaXEThLEYz5q/CHXif8v/KbMkr5ZG237CoG4BtU
Oto6v7QjTuLH7iL4sEoz3DKg2GAwECWqIZcdBZDu/1vsnZtgOBpxRW8Wp1XEMFrbA6Tyf8VcE/nx
HYBN69kSOM9qgVac2KMP+7KxlryTjjSzX4qCOn8IqbVGRyns/hoxZIKjD8tuVQI78whE8ombrhje
aLWWpRF8exsFawCRXNotY0MA04eB1hTizCIpWVZq/OfWjAT0UHL3OHJwiFAfqYlztZ1nLa7yDjiP
Ug2RyQnswI4trbWSW95UV7ESUKge529P5dzecPm7j7rsyBVh3J4BJaMqyHi6KkKndtbQdXotHpNT
EK5X9yVY+s15jDhNYXiO0/08lbISbAkcaicDPNfRh+SGU+e0GVR1Hx0oKPLp7LUZIYa9ODa61cPi
STbvzlvmVw4QEKOw2agRjEtdMl5xSMrcjEkVQwsdzeZgvQK1Y66J92pkLPqJmcZYbXV1Rnm3xeQD
vZ1WM4P88V7/8ngW8WPFbyr0JS++IOTobjCFexGp5Yrs3S32RQR+Ru/IyxvqNmz7g4nmBpAb8uxE
xOLKfkZ4C+YAA+rK5/c+0+yok9Xl3hpkQHNR/m0VqIcpzDGJlpmRX2iAiVRbhbkBzyYC85jC8vWS
KGca851K4auGRvlCumC1a5Kk9KGc+Lc3i3vlZJfmiMBHHeU1M4DFPWa8sLQ/L+nGAEyp7UH461X4
OSiKvbaCQX1UEwkiMnbFhC39bJNPUoWz56IasjfxEZBrgEDl6JNPLo8oEAQca/ZtJbAXy6ojcTms
WktlD2y5n7/8QLO7AoZOPNdSGZ93ljKHO+Bi76r6f5mj4Spas2QoKHDsovREufWIJP2ufg4bELYV
A0tJ8BCH652KTAGEpDjes6jPOpv3VgwlbwZ7usyrdLmdEy/xgRlpkuAnpxdLOeUSocIxRCYwhiyM
Snq2LIDM1WPM5F5aL1h8Chpfs0sQKztRXbsERgsz0q71OBTM7mDptWOMkzF5Dnv9CjoT6eO/OBFu
cjyT26w3l6hI2i+ZjyOTTShuDV8CmkYcl25QAz3qSkSq9dSmCw8yYb5CGPTfTUvJ7VHQj2vAb85P
wy05oaG/8Ztx7Q5KsccoAKq1WXgJiaUA6hba7Dz1Unwj/9K1ekxSjyOciV1ACMa25fD1O5K0bIau
/+XFwdP56l+9exzm6heeRaNXaQlnr/gkmXOnFU5hZ+Z0xN6pBxBAmH6GRq0NdeRHpvo99u6GmPS9
BS8K1D7TePLFL4PasLqS887IERLWJ7/STGNcTCHZXIMeAbHqjgjOcU2bY3wLklMTM4PQ4kQnsi0R
zTxU405XuRbyLNLpD9KQAg4n/W5EFpWzuOQmmDNQjLCnPyRxPPnMtsjbEFSDfB4H4UgZuPMkFlUD
MkvDbNwkMhjOz/8YQMFt/Z/acNG6YauTenfdm0dIIr+JwtGaUwUci9DgdqvkchMGbC8MduZ89D+m
kdtKG/SJYSSp39yumenJd98TjLNMr2oZCdqR6utYkeSHhxrRcAB0j/BPGe7I4TQveIWeP3f84idh
TjkQPH0Ez41VbK6qhiUhdIWHwf8BwO86gnZN+Mc94AgcvrDljFib62H1w/WSYPzcVISWy3ns2I0G
z8WqULysnAFvu6ryse1cp3NXyY0FUFjPMfHpJ5FGz7NI5Nj/EYEKV6kfKZaerEbAAzGSbaLxd00f
Fk68dx+W4uziaj4y9MnYOCmaFHckmx66wF7bgTFm9ceIC6AZd4R6O4l2Ux+cP2aic9AZDLdXuVgo
tGhtD6sE0Rl4WAk75/WXxqkws/TxuZXzTLj9J0QAwTepaWxo4e29CyUfJASKRps5fXd4ULwmWR8w
5tYweeiIkmtvKJfIpU97TqHksaOLbFuGYEEK3Buw9tTnyMsBiNrTsQMAVad53/92U6AGXVrWFhel
e6WzqW+WRvkFtiYsXod0zu4bpY2pI924pcwNYlk02crHJS03pbYKqJwKcUV7pxxuMYfvNA64cvDH
w+m1Lw/TtQ1OogVW4sAJaEtyUXz1F9Fq4DuV///o
`protect end_protected
