--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
RjMqNXNWOPdknRQG7nOqLyx/H9kWXJ153R63oDHR7naPBnPEnA6HKAUBWBUtWuMBsmxwsJUJvrx2
zdhf70mHNLRzpsIfFkuk9Nz/fOYcrkH7Dpi4hKm8LeEyy+t4i5BQNMIgQ59f0ojWkErd8zNp2g7+
SPi9+1ljJ6JM4GKovdWPHBdpEOlOEwbjTPvwtJIvI/kMyr2u05pmZO9Bz+1rTrWZVJ6pKORv3dMU
BVscqGraAiUQsQWFfidEJ/7wJjJl2SVrNegZeLS8xA75VayrBotDVrqCcUiRfoeYL5d7BfUPB6T4
iTSZzS+S4rww4EyWJeBtYSxt+Gxp63DyfA0ofw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="a0PQeXfD5w71cIAizRZ8JTVD5ZdZBgp2B4GaBaTxlwA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
hDXqxogRtsVc4ucK8P9GO2J9X+P7cuG+1/Gdd8/zY4Ud1euroZxOpUhHQZvEymkmHP6yLUuY95Ka
UsZPL2BTDDU2BH7g0AgHXNUj+jp60txHntY25ObRCGNuXtn2ow3hVo/9g4KQviS7+wZU4sX1nbFf
molmMQMBpexAY2ADjNnZL9/ksE8feuq9YmSPzqJiE8VNOE2DlriHNgk3gGaq4t77b/FXipnaDUTa
dkYH9mvcHZ8wCp5xZIhEfDlfEas0SOIlMLQ0NvLy1KCrJXZwruwkHekftR3EUz6x/EsJNRsxzwKB
94r25YAgTl2jjwTWcOn6emZ9xP/9EfmuOvN8VA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="cw6d5qQb0Zu1/kq1nEzhBmOEpV2rL3YjcGkHc/K3Mrc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12336)
`protect data_block
MPN5krcM1X6Ff/4b3QnUQ6CRnJLwJFfFSswE+Ix8blBWkDT0LypLs1tMG6B+r5XZ2fSA+9SSMOv9
6tKePFUQZTCSS6WIaPo93pMDD8Os77ZfYQKQAJkCzGSxWjlhEPb0pytGRe2gwFsjpcVthuma0+SB
w3mby5551uBtuveDS4EaqE4q5EEFzrhtssnzVTOpNbQWQ3GzfvvOrggsHSdLh/v3MvEGLRYx041+
cile4e7sPtycK964MUVSS3YlirgFYBc0hdWck5DEZPxjfoJAaEH59GMIFV1xRu1vYZlXj2efM/yN
DSpIFO0FdDjRrHGJGj/5Q2+D7rKUkjzG3JuCu/BsycmY5jLVG06oj5mEJN6wMqFylT4aVFyWZ6ZB
OpJF0+hStiqlCCn7Kcne6IRylzQqnVeJPC6Fy0Y0KhgzPOOvl4dEIRymAyzGV1OnUhOeMwMg05sJ
mQ9DSUg9pLN8/DzUJNDyI77PB4DeV0IqPqBKTAJPX9ThDVcIxG4Ddiik5zQqjZCYM6vkTVTJG+8b
HY05T5VyhQTi2CemfkMDrBaCxJIUvg7UyZfRzg/T2oaxd1+usKaqoNEUJjpXUWEAeXZa9aGECtda
+cXtygcdaSHhjDBx5n7CgR8GTfpfRhQDAwtdqX7y5Aug/YOSuMlQMiKBobbIrz8fixBF3QtJf+6V
5d2yKv3zinYnHEtm1Gyvi6xvRb4Yfnnvb6oP5CZamSNjEfCI2vmo4OCZE9M6CWVopYUSfmNgBEZj
6B98C799m7bZGLlz1vfT3MGQ0MPijpq/YABsrxtZNHLB6vro5o9DWJ8ljqoUWvsCFJMSd/1yvfaw
5SYHNcxldwxR9vUiHLbqyXYifMEYUfy7j3sdb6DrlMrIElwI3HmdKCkxGvKc2B6fCpX6e6muysqR
jwj+TlrAUHnbs7POgsRSFZ2VfMbCgztTOwjKlesRpuMtTqFNPp6ah1bb+G6YW7dcUV/oVA9i22aN
G+0YdnAdHx9LOXewIGvPQwrcG+gmSaLEdfmAachigMpHz5LF7nAd1BGe8Nywi3HvCA1PKJlr25vZ
n7j+yrDT5szvdbnU4iISgrQPU+pnHGFC9blhDy8Cclp08HF2ErHFNz4upeyt+f26o4ycVFaS2i7I
nSpFZdDhihhU+By9oBdLOtmw5yS36grZs8rZQsp8X33uDaVJYRRS7jXiirHIznbEatyUfn0LWDYN
n6yzjjcnzBt/njoE9NTaIY/FTmwDmkR086Qo8+H3YAk8vmdw+CrU991hjF/4VhPmVjNQiHpeOVuz
MPPhY3zy3xT7yMgAaFqLB/R/YyUPmMCgCgiRn1N7MS2BauC6CL7nCI5NK3AVswiYJsrymm+Zxf1F
Oz0j+RU8EwkNlTa4Akp4QBOonQcsR2Q3L7l3sSU8mSo0iGqkJAlIU1s64t8Ado7PcBifGD40FI8i
crMGN6Tj4k32QDU23O231aUjosmaMrqDhdhuESvLSDEl8vKETtvlUbKSXQujP1NSuqnZ3aq4aHw+
JqNn2YYzU8y++kYIwakFisKxU+DJrWfD6VzTFDUa99Pn1MplBIDbO58rbiwcehH3KGULLpg/CJ+h
DzBWHY36a1NFX86K5SgYePxdZQ9gUQXOmkZhs5v+OpakYsFRNIx+FWMB38oQ3XlUNiyXdi2V7sdK
beV+r+9jIQZJJb38Q5MVXzlupFpiZqS6fe6A+TB0JrIhO3xnqsWerr4IxtVUXiN9ZXYJ209gE5Iu
wLHBTgeVRYfYcQ5/qdklR9/MyZd4Vg/itD+dyaLDdED5PwE7MhaZO3+MwKvqmMgdbomwkeGJNPD6
pWMKPgN25TZGy5PguZlQb66TSsatuOmBQXqqu9XjP5DBaP88qo+eaRg3mAwUGYsaMEg8YdsL70Kw
xp2BcVbX3zXMoG8fuvaYlxHgHbzXRCUZic+xH8xxrBoOYF6498/pcCG/eFuhHrq9DnvejSgpGHSp
O86EEUlYSZuMEZnD72DQhufPRgYTSJSBus6OwpM+dKc/i4iXBnJ9gSy875fDEbqcUCmaiFCwk0/A
V4g74Lp/69bIom5ozvfdETCQdH5E8w1/orYTKcoxMwKl5eyD+pSrY3Ru2JsfFwfibrTZVMDWNwvb
E17V5b5+BUaWnplIGijOIWxBWzobQiAVNDa/BVrP2x43n6ioVrtpN1noHDTuDrCiixSZ19occgCT
4TI60sBty0vhQwT4/3wn36jrB+Z0p1z4VvOv8Qx8VaOKvL0A4ZjiEUrbbePEOzVnzWB65Mts5BeJ
HU7AQeEAHiJLADMs1/7XyNrK7TL76sCh+1xGbrUSB8+E/vmWRAI+bLoDfuFFMmpHhcpZdukjz2Fb
KtaVru9nOw2VvDNK26IY4P650qvx2qxMk8WspLkl+Lyte32BiLFe7+yd8c7h+afGCznWj17MUAJb
ruaIyfi1c7b6ZNL2IkEEvhk4iogJxzHR3eVjzCapfRRJq8MCV9qgA4cAmnJldfJRSjzoZWzRnFy7
TquqmwsllF2sEQL3YmS29A3wjqBXRxOcV8i9hqbrrXGMw7Uj1yEdXlU8BUrI6YZPtJMb6wMhmaIO
G82gYO8chSlWaJZvDfWkPPhuUdkdXG5g5h8JMGSmIi4IrsbeJa5x2QlZq4smkxgnmrCjZLNskGhX
HMFOrYWTlpbeSOpngNvd7u8aq0dxSEl65o9jtV7v981lnmhnlknYFeF4HZJuNlAesfY8zv+EjEss
oGPQnjc9dA8HqkmqvMNWfTJbL0D9ejbWp+I3shXNRUCQtVSyTiSXC/+KKB2uI4QoRwDaOgcLLwca
SOfZyKlJg1DdySyqaMp1sZ1puE7TMqK81IR2Hbp6PWe1NtXA5/XnZ3cFg8m+ePVr2Jaamuftp5Cr
4Ws4Gup/uNBNE/ch0gvC1LLPQdDHb66Eq4OkPxUiGX0NyBHF1Kx7VVWa9AvuI9TRX3PVcz/7m4H1
o3SxIFAqqa5SO1iWF0qh6CILslnH9FZAAvq77HfETQjCcVla3aKpqJnqPTb3c8x5icyRPlmDfrKC
mBEOZyFbKIyWz+QDUsp5zh8prTm4KQim71eBajGBKGZF3+9yIlIlZH/Nlnxyj8uowXW8Yv3MKshG
4tbZri0JS2z51EQC+Fcgfbk52OLMJC/yFiH+8YJqDMVOVom4wn2WWiYrGpd7yPhFRX27irwNGW4z
bV/rpl2+alsti0miHyb8CiCB81s39I4TBAhtelLKIKZ0fPrP0xinYcRkZH71RVc6VKMiSCFG+zFw
YyWl3cEbwq70ZiZwDU/9C93OND3GqnhgJEukF3iWtkIB0tinfRDwKIEiWS5GCM2FZAiTd01PwWnt
GsEKt9/rWYsY9QZFD3i/A8vFLyn0Po3YZceRjNyYTZugPpYHfhAnYJykjSmQU7/3w0/BKvxsjo6P
D63ExDdv4DV0IQZkowKBgII4hnz2blq+pZYsd9QJrVDucWCAKZIF0lSAq7NHCkMOigq2DghVkjZ6
wNOUsimpu2Q5/PjOfbyu49eUl/f0NrFOuk8vDxsPAZjRuUJ4mZYExOWWRJu+IVogaLOcVibqsFvd
s5ovRkIBIgVWLFHZ/TCOR3f69CsFBY7MvKt9SjGJPTC+DRpV9lxpUb8NHnamJQXDuFQ3sin9TLPK
F+mE7+xfEDkD3sbQfp32Tz63Y6NpQi4yiIZf5ShON48v79UHXtVy5T8PfGnnViKhz0BJdyzdsSAJ
e8MsgZFem0OpPJhS1KI9C+XmJBSRhW053+2hxdst4+LMU2/DisuJhDmOSR0JoMlc7mqu2//CZOVV
ljUPuCR5xO43du/Aj2TICLVm5HtApvmALKHVim2bXdVvkKGVvC6tJTVJhuQ5bnb8TX167XXYKuRH
5DE00mY76Lo/MRB/0M+kUao18OWm5e0Pt7sFsdZLt7PHmWv+IwpuibIdJbaLgINzVZmxJLK/ay8G
HiQFmwABTjxECmd/DvlOpF93OPhkrh9ub9WaE++Bj0rEqBNnJEnO599ftYQ35GyWOC/Y9awL7EGV
2fp+uU1IO5JFPFuiUr/qrUuIMyUvRdpmcAsnT/Ieme48ErPeviaNMtPAFOZitg5eT2UiOgPWhvSO
1a9eE/6gCjlJFYoCf94/6m19IE97MVVeuZEWUJXZkeHJM1Mtek79z9almwdJ8rk01hipWwsLlLeP
WQkbdhaN9xK+/GHSSv4wbrGFnkxN91e3/GyCnoGrSBE9eERLRT3JjWymzKrSuygiMuKDX71nqD+X
Z14j/45FiGUIFPmKJ8nD3amQEFXMUNq+iySg+jnh/46dholHEa7T/Wv5HsQi49jRvxhofMU9kiSE
K0wNbepsC4eeOSd2g9Lnp7ua6ObD0uexzGM/KZkDsPi5bYvPo3JwOOILFg4JKg/huxmKkErvEpiY
FNSl6crY48rqHhJQZFDwudM5SKcT1Zxm4bcODGYGjlYR6c8RWxEc7d3e433gcYZ+/pagmcFeCRHF
RxzDfZYvufRsTYgagGi8Rhd6HXxHTi7o7thfJjzYtg9a47nbKgDkx6w3aBVrrHAMrlIXNXbEc0KP
3YEEQYA6I4zMty8i1eomQCkqaX1cmMFUYLi3BPHJSbO8MG6JDAiv/BBvLAeaYfY4Cgd8VeqaDyR0
VnPBInsEt+bZKDf+drM78osk8qYUXRVi6uf0MvUMocFWteulSAMVjmXQzBG1S9abNRP7jLT+yyi/
8KOxHhetgSJSXYJxOyld0uGsW9ZHwOnrKK03y45tmx7opAHV6ZwGXFHfyp8f8quL1Csi+rI75PDX
FSkNb7BMmj6JLw4vrG/xaOJGccKkd3mUPBIUVKlrfJBUiS334e6nKtFGAy2eskxIYrjWZxBNAu/d
348rfq2XbK8rkdOT3w+WDaaZ+5lVMbJu+bOwmK2ejry6u+P8izupXGvSqrf2uYKbJdrY8cLdOag7
qLsL4C5y/aZrKgOdo1WdVLo9dvvvxV2thYtKD2Ene5v655VrdrBa+6qLfPYZYsP3typSXnWpjzKk
d9u/hEbix4fRIpeUEE/LLA/wHK50TKmfwTTiy1zwfiUfcmh07OyxepBGSEagYGLj5AoOd/kYTAnz
x14Ts/qkzLUsUXWxpGeKudcbum8xSDnev+8mgbnkNHuE/SUiBdaMU+/Fy0QM5oxOJWA3+jOiILsx
vjKRFewgS1G4JdQF6c4TZw0zUmB2NqvazMdP1s6hEBj4g4Z3uD4LVwDvMqFrdFbj2h6mMR9r3MS1
kqh+Vz9LfkPrP0vJB3kVpbbkr9R1Dqpwa/MJpxls6xe5Kr0Q6nFuZPv4H5pD3Rr1ojsc2NCqEbLx
myRoWCMnxdnO0exwRlXFtiwvevxMEAclUt41iAfx5Azy7/cP3FAHkrCJeZLs9xPsTP8wt4j70pLP
Fnmbhj854MMT39u0Td/aQ7//VCx1FC+HVyq8Oc+75h/Xl2lOR7FyLPpMjGJvUpseexsX6EKVa1L+
CAxC24agX06tbSesQSLUNDN/4/gdZtmrEY9oVEjH3FjwQsR9Ed2eqIHRpTTs9S7XXBRMA/9qtoKZ
QVjgpWEpkvzCxEqmQ7tGk1r9xqdw5z1NtUb8UnEN6+10xfADBzqckDHtjLWTs4S7z3/NIgiqOu9t
/lBGqcHx71jWjvNZatXgmIW0On+M3HOhtfkQOt9rL2wUKWQFm60Ae1q67oFYPjSSd0wngU3tyvp/
qeiQEYQ8AVKjyBVeGSo8fEZzqQ0hIh5b/Ptk119e5udhgGxB/dCL1O1x7tK0jYTRts8TKMqtjXNW
AShC8MObYi4vVTaHNFriFxcPjNwXoCsB+uVTeqquUkZv5OuwV9hVD3PNeHxLwoVZX7CjTCSI3+uI
5bZPHa6MJcsocgXgWUy6USF2NUH0VhIntBgWU/9JbLJA+sISYgCoCdvAN1prtiWmZMm8tTa5WONK
GK+XQg23Hk13XjkTNFDtZulxOv6KcBVvTLaszhsOXslrtTVPusFsQbxgy0bTA2ijRoTmdE97Nc+W
3o+PNt73PyOYPFyV4ADe9sJHwH7dkzmxqm6O2W3XhaXZn1jTwmUh5cRRBjfmS+DUGaUgQzf5200J
dhHfs5wqoEgHro/I+wkuGbzP5X8WdqoxbmFtRjM/WPfodShBH1af1IzlnECd4McKYouobxifzy51
TDjhVRNup3n15kY5wDl6exM8+KMMz8G8/3r5r0XzJP8ciPnrjkVoc1TNNVF9L3dCRxecyKwP4D4c
MVogszDVC1AkwH961yU0O7wTzLJQq7iOXbE2sOFa3W5D+B1iGXoEmpfIrMIvazeomno7i5s8ghqS
0IEhJenAgwUrP88wIsIKGp03b9Wc7zHjbpN6Xp5V9YaAPpIcehNYb7EiZHYqX2hwblZDg6+tN49r
JXW7ayUh/6cP10MPFfM4HaIi/1lhTJOVb75RNUI2P93gilkYFqq9ccolneFmj/9eSp1lRaOjWEBD
qEoN9YKJ/BZFEaOKHlr8P+NEfB1zWLynlXN+ZpsuCSB8bNdX0qez2md/n9i8/Pux1bswzGV1Wc/1
f20U4ihkNsf0ibYw0gIhvIIbWHWhbFVF7ZlfVHEVrkd1UKf1kT5pUxcZUKOn0Ajj0WzHLeD0vwd0
4YXG6qbfeUC7oP2slCRHgLK2yKJQRJ392NTJVvA4VXixy43zd/gJwMwPFUTOYUQk7gmLzm9coTmm
oLwaiH+J9we/2mAIPHiBt5gZIg4mh91HpZxCZHlcY0JRp0cxlBwlK2UzDW2b76HYMFeeuN1L6k8N
ZQ3SjwCKsBQLK/oMI6O3h+NcPWLli2uWO5V+KgShfe/MMGL0GqnxKcPSQBMZvx2jmM4nT99Uy/Nc
z+putVXIeSv4U7YAlH+61Yho0X/BaWp/CLTuLJ67vg6MrOfFZ6KCt0lwj8mNZeUmbhDtFyHK4bpS
VOQMXDmDrAH7qCMketMPrPqu95+SqASNWAOakpFg+seX0CcSjE6I02oQZYErmT5Y9ut9Kwvkb12j
POj3d9OhCSnc0ZdGz2Q6LXwhi3n7fAIYgk3bmbValwY2P307ZmxvmRIokzai7QEcMnTS104TrtUV
j7e+LBxcuMEwkkiLHp2+LpgxuFnvmWCDuQ+KcaAz9VHOCLbXFeaJIAXHZ3MA6AaTLVGY/WB9NZBY
+GyzP61tpJRP2Zs5+cm72w4Q69tWjPoqXtPcjRFJiW4GKyyqDGZ7AGbzfalahFu/s5F3/cc18xHW
8R8ZZPV1ZJg16ynqHPAaSHk9EpKFJWfbuy9T7Tvxbs22dA26+ixTncQAfyi11J1GZzp4756kxVYf
r+pqJrEz/UuUWNXL976TFJb66xZuxJXC10zTeQkEagKbSBzuONNQ+onank1swmx9gX7SGDQwulZo
fFMVEEja5YDHusTn0f9A2ro+P8gNsZrVP1vQ6cVlq2pGZFGXjKZ7b3DZSJMn90zpir2RhQaqzL1e
tFZrKd8yo5rsS5Ul/9kXSOYXsS3KsfBaVyfszBVMhBxGVqvV7Lo/WbDs9u4vwhgXillM/I1sbI/6
E+UTbrSNmnxbRZdV+QPfJdiVR8elb/z02QBbIslmklAxR4VMaxtUPl0JONpiXI9fBLxjDjwQ6Ajp
+s1esSFZoohJGhporl8+IPIhkxvgGqlNFfNKEPnWEL3Ea5ljo6dE++q0gcrjfp98jfdzXjfOgNrB
K9uF89qDPXsOIg6RaZwH5i38ot850OUMQaCTxPytdwpxxBPc97ug0y3gJkhEaDP80MPY+gjvsbQd
6vunQDKjz/3ipDeL8vtipaqGtyFLP4vxaQ45xPWDByKN7IDCWC4POOnhqBQ6TN6z6/iE1+gW2XaS
DKwmO2bSjSqlXuqr/MvEuJCwbtRfaO/luBLeuxjKLy17T4V+QX6awAAWFtz9Wic2P3Qet0vnrVYc
8uNB0bRA71+Uz5Ff629zg3ZPYpVc5bf6Yil1boW5LL9S58Mn4diDKSfbwE+ZPtIYu8Qs5P/gyQlq
a/cE6tn0zt3p3+ua2YjfKG+4i/AWlmeO3hlXpALNMYjXSApU1bncfnkd3YHRux1UyTSOaX1VjFkV
9G/rkMK5cVeCKV6lDyO0CAZ0Dg6jbyUoSjUMr86X3SJLamseYL5qaq4IUWiaNTaDOWlQ0kLhwaYS
uq74S+d/7tTJNf+aRowWcYabi7Hl40Gtxh9mjY4xwI3sfsRu4cyfQ09pabXpxvCPTWU1QPAp26wx
vnnHU6LW+p+GuYtnZc99ceKxxoEKyWheeDRopc1Hw6TvQDuXkOVZ8hgSP7symWHS9N6qIa2Ol9t7
BDA81zJieGBYxRBCv2+USKCWz7tZVMjwuKfv5UThJ9uph/wuNbHgqzeDkBRdLRVN6nkmS40ivQ6N
nOoOlHqqyOHb9d6prLhdxhPx/4lB6kTMmC4srKvIHAI+gR38Ca5jxbxXNxI+/kgHYF9dF7ec+o/2
OstU0c69kZuNlWBoBzSYBBA7K2kg8DMjZQVV8exFPfq4PNsLg3N7h9bKksa1nXkclTvAclSsp1zI
bIlHoz4pmaTyuEzYviBi9KhKaDZnpMu6WXuG7n/68NC7sTeRWbXQpVDGmP3iwSwn8kdAbD2ERM7r
aWZk5VW0OVkqpIRTKOmdYIXZBXqupQg7XxriKH5wK9pbVZU8eDdGJXg0dD0o9rCpbfb/TQswpdHC
l/7vIjjYrzW3HhBAxaS8+D/uRyv6TBMbfH1MZez4ABExmHuQCrDHcd5N7j0c5PkiPdEQoIgevb6K
4crBwGKX0i6s+7/nXjzjr6zcLvaekz4Jsd1LriOrSOyAtFVFdfR2mFjtGjdj2icsxJ17Y+rSbbpV
wL199WkY1lG72sH4Xr7SybmNCHAANqp/iwcTRq411MFRnTk8nn7dTOqcei5oPRr2+qSsBXwnUwmp
wSzU+w4jsYHhEMpfTtUT2sHWExsVR6W6d34Wnx2uK99t3/sS/0d0Oycwi2LCYi2Lbg8eokHpBMR6
/JmgD7FzTS6AHinUEjK35beD5sxxc8fk1sFbnjYlmRm7Fi/uRVM6qDAm5BzJOCLqDU1Fnv6zmnQi
0QO8uTOA0N5Ua3ttsIZ6KXlh28lcZEhF8wIRIr/ULihzaWx+QT6W6oyTumJxdjk/NMVl/5mTocYW
0ygsiHvNpQ+kEF0P1hmyTt3toP0XPdaZ+JGg/rvR/xgNhNodIpm3Kn4wms7tqk+fwdYAgZrn4wO6
XXPykgpRFMaU+68vF6t91U8YEX5yHu8SyRXjVfTA40ubhVUY5k9uz5cBI/96AIIVMHHupFDg5PQV
KxQ+9ExEL3h5tLncvw3MabX6SLClBlzJCB1chOpa6nZt4ITPL0EyjZXxUtc6eunAG64Awi6WABkK
ZOYtNLbJX/SDGa1QZj8DrKF6PMm2MSbpt0VTyF+U5T27E760d+DCrx/GugJuU6s2ucZ2GJJnJ5ZO
2oJnayvmRo7FfHA1VuhAtdqHIxpb52mZ3YEvfevCH9Wfeg5oZJlRxyl0jz2zbg1SHa6cIDbwT7BK
oEhGmkIUwUB4gz6K/d6qmzEnIimJZQT3Pz4YxGdwNS0EwmPhKS51hi0BVgDIf/jixPXfF3tJIKBX
gk4kp5XUMkwgmV7LLHubhIiTe8h+Cq+BM74pMuo8iX0C8vBQEMfRRMvHj036pT41ALW6r0s5lZJa
J5ObZUMsvghY+vT4BhXEPcS6D55IQh0obfDS7sU99dP3sh9VRNM8MciNCR5t/YVEuepEfING+/yO
m/bqTof0lR/nsscynsaEV3ZLsyCfMHS0UnP6Zp/XEp3zHeo0AbAIPgKZAT08awnBF0kQ//Zm273Z
OI4vxxwa1ZWRpM1E47aZlN66YM9v4XjJKsRON+I5DTXGQXeUdCSNdZg0VaY95h5SHdaQ0YAJpR4M
Y98xBv2GY1mD+sLqxF8bhVAy3d7YYEFCACjZPVmuQwOP+k12uqAfYJLm85vVwmOVMq06Xw/kAgH6
cv9LuieMH7ISqvu2inuyhME5eC91IU0FVPG4NVnBL2rlrUgV6zF8MDalSaA7NdvVPBnBuGriBDgC
YIMftx6tsuf4nnqn4PHmWjEEtjtosfmUG14qK5UCtBKYJVYQfBNLJ8EzSmpIW1iObUqowR/kyBb2
t0ctuhhh14k4NYfDJauvELsESv1+0D7rx9WJ1fTrqTFV+DiWqYOLOd5TPEGSigBCG2HaW/XS1nHS
6A/w21M8UHCcnIq7qQ8tWhooNymxYRbhlKPuL+PN1MYNZD7A9Vf1Kbn54V3y7UT8+Dd07Xk4hdND
gE5MsTQ6ENUcJPy529FwUpb5A2YASlys74Ae8zSj/XkW4t0PKKDWV3VX32KFSIA1dXDc4HhmsdOd
/DTKuhtEhfdHwawdKlnUfjFhgfGAZKldS0JAFj3HsP0dajXgMLwdNrpvFaWDBHv8UhH4ld6ie/GU
gtGTKtp930ERSY16CoMWKg1YsoFro++90RIaiu2GRRNffs6HuF+n+1G1FNWAeg98aaPLPnquYgcD
icP+hrbFugcFt14jiNFSugoZaxIbxS9W5DU3yYLyfpprlJOvc4pLuY9dLQWNDMVbtBcgjulf4SSK
wt0DQugn9kT0MCO3NCigpvhG7RSYOjbgb9VOppqCdoP6BP3/vCy6IfmNjhKYz98MaoSKtuYMpLPS
vKXlBsQFd4fW1vkI+/OMPEfLMzzU2GPrL709IzPhEmxUhqSBQNc0PvokDnjkCd0uy4OTotIPRya8
BdYwnCQrfclBUBKuu5r8NUBGZlz0+d5gB/EOY0Pqu8qo44B5Op9+viSEGB4kETJKzszNYOSdzbPF
RhRREVkA555BpFagA7epOotrDVrmu0nGBMMrELBppsVKsWm5y5RdCjfIm1mRg2izPuoYyfCPlkfJ
Uibfu5Lqi/CETUnfeaMjGUzCcrtQUiITzk7J1qpZpiZl54vwMq4hLb0UY5w3x0F7ho9i8e5y/3Rf
vvK53PUx8cQk55P8zN5o/HtoD2WVRODGDKMeoMQ3RNiREr9YhbdXzoQi4urOKouez6DOYtwtpjF+
0Kay027dMcC3S5qDGoasBC6CXNd34H4LleizFQXTqFNzSON7gZXH724FdmtxIKGCwBcmRqPnDgHO
zsw5f4Rm4v41fDc2ew9ATUvMPYvn7zC5UcTEHZUhDiwgPHluB++D12ncUXYk/ysw22iECFBheWK1
ZsF+VJ8WIYQCBKmNLUHfj/ntJ7cU1Ht7o0GLnx2vQWImWgfRNVHwJ7hQ+KP9JmrbWjtwbrUD2l0g
4CbD7X3vUU/UjBleNy6uRjOVvulKrdjfaB4Lu1dT/3p1hK76NPCeE7WrvN6ScXll+c2SqPt0AB9G
G8K5KIDCWsQyhORHdk0TDot1+MdY+gQsr8E8EvVM8xLT5s43IwBC6U5uZb/J6B0A1yQLTYZdMcZp
ugu/ASOE7PsiEeLqpi46EWfSwYb7j1dk2enXmlnLSJFER+FwKuYXYaHoe07Jr1xIB94Vh0HGm1Yv
8QlDhJGPJ+zWTsnliOY0lh3WL8v+B9DeaTWWEQSSG48IjtnWbIKxfAx07yvWH8wN374N5mMcfsx0
YAZFHZgTtm935pyPKrijHgW+SLAI46XX8DcSx9NLy1TTIatRyMd4ieuVZul+pmaAv7BFbSNVjIv2
fTC4GLx6SKiuWmAa8AmOKUf65JG82iZncDcgY+3v5Wv2+07XlcFSHsuc0yxako0YA1wA0imRh3LX
34oqt+mMr/v1FUk1mtJrbWveXz04GFlRK8VD1rd039CutXtJPbNkQf4kwMHhQ2Z824nPDSDOvcMf
Ju8Dj0Am3eO6vK4O/mwGGxKWqhWCzocRcAmBSthJmZhCHnHiKx9l9Dpc4mMZh8O0RD4bC6jazP78
ssqbGBX4/DBqUz6yVmTkIl4aVJ0Oy+WOLmr5rPM6iM4RrxVBJMOYD/f6HzPTBB18EoEWz9IqgCuG
R7c7AlU4V0eqr5Savo9WIJfcdPDqyM1Uib4o0ZEep4STSizfLfHWZScmvDgXOIlD/uaRU7lOpjeJ
nWuxh72k+GhXYYue19W5U46OmXIaw/CVYCiAe1Kh6QdhtwVkvpdHoubKrtXUF2Onr7IMxqj1uKnG
BS+VWdRyKsuA1JJpZiYELuH9JbBFGqdpWm4OTVWTs6nNEbb+cQU9yAYAxhSAFbgiVgRd6VvKMxbF
6Ssdsyq/wqIjHBQAuRTklSKSifr8/iYfstb3fN3h2oaeo4ddEmXWuA8ri/rjJEeuSU2TyjGoCx9+
afBZbBl0Mb0yYqZnF2ofQ0bFdVJZbgSGfq0/uSnKKkLTN9MMD54CavravZzYNdo39S78KtY8MZN6
AcvNnX4ef2GRUWh+pKKoecLLIfp+c3tZlWVFy28lizQRNYFepnmjiTJokGPDz2QEmYaXC33hRfiK
JH5EF7f0RlfrZUEqkqnfSwRT78Zypcp48gOHJywDUOQYKOsmVMW0Vk8CjAlLyEjp25g1titArkfu
Dt8ybwwP8HSyfOpxXc0Rnc0HzqqOddLvcpHP0/ZKA5VPt/XvK4bKub4Qld7FA2nMWBIL1PBB2Qsn
WI8KytYL4YHw1bhaXMEjabOTp08yBlUK4T2ntzPFjhRzIfd5b7DilytoCCMbEjfXm4q6WnKoeTkr
2mdidCYw8B4Is1MU1aAesbxvuRGJVIUoOg4CWZKkwUhQKAeuVg2xhoYDa5RXktWeEmHgmaxI66vI
xchPpolv/WQWy8qiauM76GBsvHasRe39iQVK1Q+S9/tJ1UQuTBhpFiHswIZQiCsd27l/QujSow3h
wOPPmyeN/+UOVEF9s/KCggjhFlzqaKwKJD8f/+u45lFK+v7gA7Po/8L1Izrkmnq20U2WgRcWyxSf
5hBfHzdMPp2d7jk2qZL6nSd6ynX/cuXYUUB3EqckPp91tG9mBQDAwWwkiStAoWdlJTQVyFFc35Vf
I7o3zUVWTf30viPqW9qYdfz5qDB/DEsgaY0DG7ShlePzE4i9R6IRQx1kloaZQn73lD0lTwe+e+GL
txLGHpuyCJGvs5VoOUzdAyWqolnwZC6Lbx0pb68WGFq4LmancOQj7CbKoEiyvLtkd5ZcrhzZ4ULk
u1ZsqBmIGF9URe2vq0HoYOeeD9dPQBianabtF1rfwbez4ym3yrFQBUnLNfca0ucI5QaILq88+HZb
GKdSvvsIRZOT8CnvQhyJSbXEqaZjUDQHbJEC3YivvLMCbKEg5DuEVvr4MnQPoHECjQx2dO8zC6Ji
x4V8ov59GV25g/LkHc3Tlj74rbqd1T0+T0RsRi4+YuLB97LGdwcKO46Pm6j7UNyfqCWX4x05G8Ih
08mkKNQq0+hHCwKYG9LnvTo1hZ978PVB5TI2BDGbrpusA2g5ynYiXNluk7IhZFtENhJlhTD5tdr4
f8BgXy8QCpSw5R84841aiWpa9vNG5+UsMZTA0K/ZI0mEFAklIWWbSquTdJGwJa3O0w4xshtc48a+
0dLv3gaBYya07q96IY8huoewhH0sMXHzxFfOcnAsQJzifxMH0osjDHU1EX9sdJlbnr8WymsZ+zAL
NkHq4iLhFDXyoob6Rtx/hONLPsLiI3EmQ2c1EFEJHA5WDfs+hTiu9xXzDFm+rHvhGK7e9MwB3GPv
JSCNux9bifKUlZNj6zV1zdqp3IuR9H2Hgkxqgs0IJQv4qpfnbbV8dQ2hq8gy1yUpZSTlqWbh6M0p
WC3QQdA2TT0QaA+sQTaXSZXyQx9tnqd+vjqLQ4Mmf5DDBFNmUqyV3fH6rrgfLK/lC3L0+zSrw9cs
TRQb5w3Vm/IUUK9VutbocuE4u+1fs0L2i1HelfCMyAdsu1cqn3PzSa38AEievFpK9Mg95LQvZyYJ
jzZkq2M/W1xQ9/34MYRtcmgbJShGhu/Z23kiXBVvPFpUeHbSGodVpJBMzQtp4E5FgIw53srgV0NZ
Nn7uQxxK88UqrfhXnIk6G7NIXEOOrKFF/MVQJxDsQZkZZ0rP2VV2A5LxYpX3VJtEC5NmlGkIg94N
Y1nk/hpWj58+rkiXJHVRg/ttWB7Mh+0Cwh0HnJ+xAk1l8OhJSgS0CXvFJ9dyK4FCILkVRDN1E4I+
Gp0VsHXeU8aP7R7F9LGNgC9/8fKHJ0qz8VYFPanUUScN9oeQ8AIOgrITfm8Son/hvj57pPqRdIjy
hb0ROQfremYehrOy9LK1GfoR7cRuoAuilnWPNSSNRvZp/EM9Gx+tZy1oW1NLSOiHKqxf4GLl4Uml
1/+RVBADTXb0A5op8ASYEr3E0IwrTtYfokF8KH3LhjgSH3tzHOOK/kH+D8x34AOARx6mIT8h4wNq
BseYuZ8jeQ5f0nueFCxuOnLrXe/FRG2yRATs9gpfbfu/hu/HkPSomrvoOfS8g0fFhczvH93IypJk
R7AoCuXBPTFF9YkacbdmdzLf8C4CGp4yRSWTy/PUTK6E9rLXZ73VcyTaDXxmq+ti6hwGkToZSVv1
lQBO44ixBWiTPYRs29sDSYxfxD9rWZ8xkLHeCZwefEpD7GAWoLo5vBGs5zvxp08G2kHkx2ladKd9
hZ0c0MLApFmsk9c9A3zQzHkL8f9cxWZsRDZH2+QMonbMtHEabMWRvMrO9Jl1F2vOMeC7kCgqs688
tGnn5WlDw1UxDAPLS7kW7ZDmzv8e9Xav3LvDN+tSZRh4glh12dNaEMVcZgEOKdJ+z5Jz58svNxJA
/sRTfYYR6ULjfn+ugP3rYYan/6HmCSigRdRaL8TKqEixM6kZX8H30MASM88M2dBKeN1xzhDOfpjH
VCP+NtOIL0hu6j41KLzofdMdmHUb9b6bQD49bx/MoYMPpoiXfthZWlFM8g2IXQdgHhIdTJsOs5d+
JC+6mpUYNBXywVLQmxWHBsmYiIuPKOm0nD52mUtSa3GJwj7ldGgxx5bdg2TPIlJmtSIF6+b+7xz1
p2KM46k98CYu+iQjuIDF4CO99N+WaoC6WMurUVyP3oIq6756R2uh1sVnkzKr7Fu2Edi0fkrp4rQh
ZiZaKPqW6W9pkomYsW9m6FvwXB+XlfwvsqRTgYCr/1ySdr3c6zINv3mngw9RFEMa+81cycwLF5sO
h7d8IG4lbVriwKNQGUlSo+/y+B0Wqj7+iBmlm7HqAwhgUnKv0BEJJtNcqu+c/DVgbJ3Y1wzXX3m7
0Zz+pMlESEga/D692zkr6W3+fKcTXcyYw4AzdCmETxJYXjDiogFDBAcpX882/hqhev67T43+thMe
z1H9Dcm/TcUcWNRmdUu9Koeb1IB8WAD4UpCIxYBw3AJ/EB8UfVMKktMTKiKS78QmrfGQbZnvx6BU
sRjXDZ5sIoXu30V5URrzUTtmBFVAahT6BV8TvNsVucEB/6wTaslvYk7/8uP9QRu4y9Bp8rmGd8KT
T2XWfSy1/RilxyE1mexUe3/H//XlJrie3oWRy9ge44oKtzP6EuwwTiApuqiNdxtlX/KfEQ4tg6e0
jLIlOGOYcEepAKgednGOQMU49bepd+w9z3BQHZwXP8VFOA2O4tg1YURGFlxRdC4+dubWvqXkSvfQ
KEzOonRdF85oYQUH7p/aXZt1E87olOIQjwvecLd2rGYBhQmdJGURJ3LCw++QEBzj9t/iHkGUYKiL
6L/WdbQ5JPs9nT8zjXDXaOADHURHn7my+T5XKeCqiTkjBEEjYLqkqp2J0ovu2E/10V1rxErDwfEa
1MDIXdJLEEManV8i6ddynL05+7dkb97Vt4q8SplznMdQVsLkuoeM1bwvcsSrzIAlGagDT5LktPAa
QnQhJFyGY7jSEgxKySReiP5AH/7wtXzX52XZBr0ornuDcE1RbIVcDubSyGuczDMiU7o8qsdThLEu
qss4Re0t1NJUWf6e1kN1jnVdh2kQS6bJFg6yc+AnB3wBPnc5cFZcV6zDsJFKQGiqA5RDqJkdle4P
gxTG9E/CdDt5PaKaLId9NlbVfYK9Q/ncJ27ZSOVN/4Ae0lg4Q4fuLGLUQe3Mud88zMLR5u+WV6Q8
gjoH6DrTQqh+8m3LJvqMCQ/okGSy993AarO9HEhEw3VTpdEzp3YGw/R9GV+CY33UqCzwBtQ1OGdI
4FTRDB3A4072s1oXwvdVRUHOcYVfs9BGn7Gaf9Jfz7Ko4qP/y4afKdHzQPBNKPMFvrsH3I+FQPJl
cei0eh1eCHtmaKMde0xPlv3MCB2sLojnkStr/AxFpkbiwgtkw2FRFo7ZCr5vCIRrHjtytK8PseNR
8LHQ0eGMfYN0YdJVw50NUu3TwUWKhb9k0gbICqmxevz/1nE7xnLQL4KuqPidjenBsWJBaqkB14mn
N7zmAeSOIfY3JRSCVCdtMuHHjhs99vTbcHfsietDrRmzlk40bRXjfARyWbzinv1zQhTQLQRJmWX4
oImw1SWK1x81eL++qNgh5PND+MaN5OdQWGufA+VitI1nynkEEaCUQRnthd0pwJV0hPr7xu3O0S3Q
Cxmdg2NprigkhNBt8RbRt6xqTB+Mk1Q2
`protect end_protected
