--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
TMO1TfB1ifGTFDDk12BecCTttwVGy6DR9+vRbG8VrbbmaCnglrKjPpOgmkeYq7r4J1C2QRn9YAKg
3bwVGT2p5t2EoBTC5TgpCUu70ZRqoujN8sYoF6ECij9ELqVaiAixDEKI8NYzOAuXxJ/ZPuXRcy6G
zCEwWjYSC/XNCUXB1c7IqYJrD01y6rOpNxGsxLGsWHVdNfgZuwWS36izAL5h3KqqRDheLxbj1XE4
GyK7tMnz+8z+XiIsipmOp3Qb43lgaCaIP7QW0OSlii3ODxfJgOlXNkR+KO1s8lQ2R2mqwqIG8xdG
luasG03iY5wmaZZP0q6cQ8yHT1XOvVX87kYPfA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="30ywEcArj7UNoWwCl52TgtRVvPHthfLADKSaiM4x6jw="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
T9j5Jiqd4twohMgxa0sKpMh75AbREDNuAgnSsRfqsh1d963ZIPRY5IXmZBqWnCOm/FbT4493wo8N
h77X65vFjXJWIdfvI/tfwVcyWk8OeUnFShC1ndhLl1m3WiBUV8oWfO+6r7jkmuaU0uKznaTTjqQq
CHw4z6rEgGKmDS+1EQJlD87kHArQiVsQvVvdnJKd87kcoWsEfCpMbT3F4cD5gTDEChL31xsYCXqG
E1vCc1xTrA2ILs6Ri4DL3cIXi+x9xLaGe7yT1g3O7iiy8MfAbtSuM4hlBHJHjpbBDnNTCLQ2V13i
qdk9akqi/F/IeBKW/9wJXBzgYMXYT+p/n6K/Ag==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="jT+sbu8smT4l6WrpGfwcjY815z1tdJttJGphR1Zkxpw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 68896)
`protect data_block
VAFPMc4iVGfk987rO4Y2pumIIUOfnKexmOXek1W/MBBuk5FbLZ/peG0j+Yj5eYA47kZuOmbYWVoM
R/fUKZ5yKNV+9QhtkonS6R5M320DOrbDhDd26VieHsYKHr4cDGbiIL5fouj5AEwbr95ZMBDtFxDv
4nz9wFT4/6BTDKyzjf+h3X+2E72EY3FQ0riKapgqqwyvCA3U1mgWWZRVUKYl31dIYhYSscHsLTTU
jIZC2+oZ9d52qGqAFjVSyjPvw9hVMZ83zwOpsH9+WjzBE8pa+6eG7JwiNm0qXHtt1BCybLDoCbtw
bqwRkLQAKqMR1j86pENSzFG3KoG9xCVjS6/Y8iB6aeTJjlpPq1UML/WOWWgCC6f4yCPuM8NaXg+s
q7RkPc/owashR92DIsl1Afasif7YDKH327+us90Dogi5PuaRWMnJ3jwxmXiwVDaCQQuATEln8D7y
nCFHwEjLpgGgC2V7NPTfNbsIgYYhjD12gEB/VLMutWkW6Srgf3JO7Qgxqrh8Pa+7lHaKLj3PXeX5
+VNW8kYXf/ZsDa3Vn5MdgqJV3MpXE6nmrjCA04FVngvRuVszqKoqmNhdzLVl/hJD/nDI/NFxupY3
ryaZCQ041MOMAcNEL0Yi2XIFnQMyqvfh9KxjT5B/SWQ0MYclUilx3rOHIn8Rm+wHQDq+tODFCAZg
NdJokORWseP0rG7F9FJm8x/z6jqGscLBmt2viUdjSRxwccAJrwKgTVfuUKc1JdJfkO+MSdpl1F3Y
8QGGSINwpSUDPvdZ/t5QboTy7RQ8ySWh2b/Z3VHTlJhaqQlXuWn9aS7W2lafmPyQ0C30D8j+EOJ5
wEXF3HlmWltTOt7HWFH039PjBB656bK59TObVyT9mXLrXYaaB/yZOgXMkyHQkGjELzfRO0OE46ne
u14sZ0uxAMGatBArsnD5dx9+xjRZJMwuMqNmF2tfKZXSj7FvkDlfkQHKK6b4i3fD+Pn4GN5mR7aL
gGN0QUNz1z4uMmrHynYY72B0A6bZfKAB19RjEhIRPzmGMcNLSZu5NIDO1BD0OigKJxRlWiOmj/lq
2Z6Evz8Yo4ikNsDh06fxmEAicAOCe3/qEhFVga07VOTTPkratwsyEsM2fkMWanE2cbQR8GiP5lqY
mpIm5Cnsi3gQ9NNFIh31xclzdMq5K2qJ8pnZmavm8vdEeuje7iejEwOUM6nJVlr4hwNO32GO68Zw
aAtfikjH5zqs4cHkOJ84BbjfBYYmt9c1TyUP77kRQauPLpaAjvHnaTeMVPAM4T1ANZSdEUULw00W
yguV+W2XhR0jSpDfBjHwFh8KCp3INKDRCmdIauv3/vG3Plgo39O+oDH9qkBslR7fO2eX84aJjKXt
Xq0UbjLdgB6+VGtNdSrQiLJy8wEiwdD6s+gQFQIIhSw8fgf9zW89IENYx9ISF8ax863LnOj5lD1R
L6rClozhdowBjf+3OGKNHjO4M8eu61Req4NT+865tq2cyTulguzMYlrPzlKVxwcdG/yw93l+Mkjl
glHaaGlvLWPTCREjpYAG2xp7woCV7T9c6HSogOTXv/B3jXDki3WNyhlVLFonAzvmGmJHLeeDyJ86
2bnRqTmh7euEKOOP70kcwSV4KeFGNJaOmWtX5wG0nFwwsFxzoo4A4ksyWLDg/JlWwaEyIAb7jZvF
EAK2yaw7aw48qa4KPmqj2YT5HFFwHtza8im5JE+m2L/AU/jAkAaykWtn2cmo7L/008AFCAqRUipO
/2ZJ4c8jvCBHg0dJr9D+qtnOH9CBu/PaQtdDzsaWW50c6VV+9kq0uQrU+syHL1Olw4jjz5UEmHmY
nlSaN8Xi2bQDt+NbOwgeO/W3Crft9/Hi9a8ALT2M+1afYQYBTJ2nVzsqig4bp7YryndM6/kOpa12
jFLaJlEzuvEslIbwfq61wv/fRDQPoTNlVP8AoLp+PHnQcAqw+gKyhMAbzFraWEQItCsuUNy4d1Xd
JZUe5XJESSTLMiwCO0kHuQ8RSwEkrMMeUNj9K3dnW/kLkJNQZAnNCcQu6KVoQyGbQloD+dbYDBbd
yGvLbACDQTmHOJAQJ1Jfeb+M2tZhkiqR71i/wFANXOJUoBhSjOS99KBvgnBHTGJZMup1e7jl4+fH
6ezmEuLvOrFnMxfFLNdoy2K5HIh2ikKew5Q0SGUonE/g9EdNS+Kbo9LLWuUJ5ZacYgMXSpLuCCZm
/ZYaf6BnP1ksdLKaVJkl0C+G/c/qBB5+QJHDxrVUWws6bBSZeP6y5Jo0cPS3M3YWuCVNzJuJ28ma
1s4nPf6Y2BV1lKh9S7TK+hJ0PfONfJkNlHZJE3aOuiOu+5QRHcUDWC0sPvXoRsDAyQPqBP0tDFD8
YWsKDXtY67omgY6zZqyrj9+rhSQLcU1JXI0P8cGHd0dDpZz2/9H4BmghgO3pjECObybMzampBHix
ylJGZMsiZMhn7rx7ZgSldFUh0/e5c2KWoQahDIA48XW9KiEbNVIxR8iIrJkSBQnEGfXpI9H3nfiq
sZKMGDF52sNLu389MV9VpQJuXYPTzeJBCBdDpL8JtXJCYfNqwX6muBfTbpuEvUGTUIjgXSiAWyPS
WSrMM1mbKBYEe6LbAhIC0BnlLb04PIwBak8nwMlts5ZBlj/Ihgf+LLusHYZW61L9eNKu+/epbPJV
8YVrLJfs+FW7baoVIrZpSs9l4ppKx7vxM/3CjFVS2CmgkYOUYjFySOpDnz0HB1boHL+PaijXf/Po
nMbY0zlhqFAsOFxuntsNKEy94v1fTxJNhBLe0RWkX6512Q1ykL4oRJto4bmoX3nGz6tIDw2Mw+i8
210FbkOh3b6nehsAkfX6LtZW7sp+l+y96RprLj0pXh0X1VYRd4f0TfNxF52Zp0TvX6s7J7GHuXBE
mtpIvBGjDubtlGOInDpTH0e1LAxtKvpLDJwpS8tKBfLS6Qr1b2nSyrCXTuS9oY0O16MIMU6s8K7a
2OGRi+tS5mYM3/ohRN6L1YEU6NDQ0EIxJe8UW1ID+QU3+SbosRbui8UUb9+oRuI6JZPKOEEXXThq
FmdXjaRyC/XN4bV/4F5hHV02H+xBS6/jxndWTSr4NJ+2DF7XLs7rwzihPzKfIozsVU7+TPPBGY3q
2jeJP5liBCPbfuCfSwmCkk740XFn7HdZa5DXuVufFqA5W1dkLRl71J7q8ZAE0Ajc7KOhC4yNqNBP
+Qzbzr5sl82htiznq69uYh9tqeqEaqXaKGyViZxKWpd5ZSWYCLzDD3JCnInPWO9UkMmqOsHEiw5W
vuIWNwWq5UL3iraP2uB5drw2kL8MlNtWh6iNA08h1stAWCGI8rZaYmp1h60lrxZ7rJM0OeY8o0P8
FKg/vCvZb8tY1MOBMcE72CVqWySH+42KuwFjn+0jErfiiOqZKEJ4AlQ3ovb91SOgREH5vlizw8YB
/S8yfM+m0dnCcypFjKcfrBF/0VFL9NKMv9CJMxWrGidsB8otY3U8mHK+0fpiqxgY9ZtMep1EMWiv
R1IJz8uinl00TbEUKdX7oVlUBBTWtoVXyytz0fLRXa4JDguKi1Z1OSAbKgvrXHrVCvsyAkK6hVJi
wqjo4TTMLaqAU3PazrzQtjuPn3l3tjlZyz4Y3sRmpe5xIz3ILQIcD4SLysQnb9ggs5yN32VDU1BT
RTv7VBZWupxBRI2hLl6yQTFbGuiGN/9v3Uq8EB3O3/fk5XrZOlzXcUXMNX4VYA2thNYGIZ6ft7Lu
mxo3tsvr2DVMKcWHhDWZkWIS7m1FDNZUtaj9LCNB37iEEPAhBcYbuN7kQ2o61JJsrw2gCkeiBjkW
uIQBThm+nN8B2QA3LmPBnf3JD6Ju7EYtF+e3L5jM5BVKJRCNv9Pr3fDONLN4H9ltWbw3uTZU0TpS
NgNFgk96ki+3kK4TL3eIlJCQdndzaQHryqg4oVFh7pHi6E+yLwaexVUSgipRTxYysXmpvoF1cUdg
lkbeyESD1GgqeXuZR0KX3Jclj6BrkdRoavPLHAO6zFYatNt2ROnkAw6MRcllwXUsuc3e/RaiR/HL
M5sB8oqfoEf1q7mdWVWLr1gI+JAdvZmFJtSe7NyGvXjfMhZBMnrOdOjX6rMvKTOP2iKdWxB1Hsmc
8jiHSpPhIWglkiYuC9CpMWzC6vzdtsKUZhIkT8dm2U79WfoIONa3X+oUshTi/FeEjzNEdHGrn9Bn
T/yIQ+ZZimEltcvtUWBQRHNz5nJVXTlKICPwZLTWu3s0wEgHiazgX17FJsLcWXVMm8SVX8f8Rr+e
B7Vaqb0jxIX99icqgGPoHvPeNXk5cyArSnlOnA823Sdiepnv9EO1exdMZFdYVg6jdpgWQA5dhXdR
aHcW//ltj5ZID8rTqZ8P/qvqLiBa6kKDVPacTNXf212h/djUNIzapsRv5Ke3od0DRA5G7XfOChLy
oqy9Gof0hgl/E/v760vIEPdXQBZaZXkW80mEsPPPd4MGVEtWxryFQERtmd79qtK/4Dgjry5MlHvO
hXYxbafVJy9oyWCRO9nm/ga895drZJd1olULWo0nc6OyHphM5/5Uhc9xLHYPOV635tcjlmPmeLi2
HW3bn5u7z59I5luBWcwnYlVu60ZGX2M4SXfpQ6rodg2PjWFoiYgMbgq98g7M6A9leiURWeoYTpM9
I+RMr1pOJtQrDKEX2rjvMvKvk1iwHziLtwEPEYQo513xVgb8ad5pyvvz7VvBWGf6w9QR9GJpnZgU
5m19a15hhehvXd2JQCMJeTcNkvan1FYL/OkSAQFPE2+rZpwNH2/Kn2nfdNn55xNNFXBQa0C7PWtT
JAM772MLPVeLCulqG0AmVPW9TwM4fkNljYQ8U5fTpeCbK4QKPwm72fbCWpgGyqQV6+Xlcpsc/n+y
cA+m3vDxUFMLyIfL6xQk2a+Cs3SQG8EbR6g0Z82iCroLji1eCQh3qKCLhucKYAnow9vF14whWbUp
/SjTy5WwQwDMV6kCSHsQ4sRMWnY1zwwf6zkuTIayzt/c/8FomWBr6MvYTwZ2skhMgF+uuGWG8qTb
z4yyhgly+vO9qAF9ToHoGPViA3YAb2jKetcqysCkVoMIogx2UcN423EEE1sKRwYu9DGQRWPAairi
rLNF1H7ay4M3jUIwTpasmqyDlIaMgHJT2Dxse9WYYG0XdWQdk922RnD/b5CeKPrBfdtvtBkQDHCf
pXJdZ39h0732FHy0EkYK2SxQyttCzr6YdnNEX3WuHiabojrLujbmFRSaEgj4g5WoUuM7Q16jJYGN
FFo0EANN1x/V6JNeRhZ8rKHWegVIfIKn5UarH5sG6GSMbM8BSCRz+bEJLUT2kS0t3TjsUXe9JjLN
AGFyFZc+J3LaR/5TJ7RBvdneTJmvt1kpRob2g8GZX1ESUgSWhyzOyMUVPRZps2zSJkGv7Pgo/eK5
FVGe6a/SPX+J3JcGE4GmyH9fX7gxMLzY7drANbrYsgW6egHald7MNFSi/w24mTmcc3vL26tjlB/I
gMGBKtJJT93ufM0glOuxVBWOI5iKgEbdDqaD8xMu2M91hO0L4RS0azh4Zqeq3rTGEASceZ7RW6Rg
Mvohgzm4qSmQtMR08ihbx3wNTmH5diHil6nVtewykj2lH2JmxO46jjye6a+NoYMC+twdV7zeMM37
+dFa/t4QU0vdeRRgdQ9eMwA7zXjqNZYyQVM/Pe6eIw7aIZYJsiexEbFAkkd10CkOOlRBgTeTveCY
guJvMwVp/bfxDwG3P1v6Qn4EhkS5FajJpW6UZfLSTYOz8suxLbAtasSR+fXlQFwl/ZLHRqLXVDqp
mzb6Br/Bl6zYj3qeyzch8xMrcMZhLhuBPMLqhkXAGgQYXqk4WuzAB2HjrDpo7cftiaCJlmLwYeOm
iw80rP6JUTwp3bJW5Q6m6pJuGg7BUxR1VxfJDj+EWXVEOXAtAIm6EtL1Tjx99NOaB6hVZRKNILtN
/Nz9N0WuXhUL5N3npNAGpW10mN/voYoPpoQTT7lWFfnspRlqkDoYlM81Ebt2XFDCm8Ue+MGNpV4n
kPwO3XPLpPYGLRqVpgobf28nn4F1fuPnriE89eyBNGplBS8iKId23QqQClUaQYPkLr3ezY5oM+F1
7AQwNxvRvnJgDDr9AqsBsC5U7VaUgrlEpgGC/GK7NT0SMbb5n86Xi1zJAork8lL0F8LwtEwtct4Y
ohAGq6wNcU2JKW9gvRimZSx+55h+JEVzJQ1d7XNBP7svy637P0hnurcSOqA7Ks9hXSjZBcF0bEqJ
fjHWZTBFKxNM9eWdaYjJYlNhft0D0VbBYIkHCRU7ZuVgmL3r7YYgVYctlZ7teJnXYpy3IT3aR16z
bKl8a9IXZVBMf/Cuf85f6WIqEnheN1qS+aEDtrCxOPJj3T8G8o+120KIeA7EGhJcqOjSJb4E10zI
k129cF9cCVihwQlxoVOjd1WGTK+ibo/eYUADwbk7OLoX7/gVYAlG6FIgCKKjf3BITAcwFBvn1UjJ
FDaLYWk2I7y9Q70lwr46ptiYSOcLG5tKNingoEMlWr9nGFDFv1/1RAiLlMf/Dq0mzX8tkSNL2RVd
bmI4fYXvWgTpvZOz206CUueL4oRttahQPmvj4gZRlcdqUpz+Gv3lCNbzFUpjb+lc/Nbgg3NX8NqI
nhGTLgmn+WFmOwVgCpef0bbFsu0iZs7ooP735rL9mvIaQtizdNP6pmO/KpmtlYjYexgSXyN0KGIB
k0W9dZZ/6lMRhMBrvRo0Hcz5j1+VZKXgR5QAbSEGRJW7bkqKjbsruorBcnEZ5aWZ5ERnTJbN6Uj7
7F2++Pm4CHW2nEcyMw1cuoS2L7d1BFoPKIuUxfZv0FFKMKpdQHIzwCFKoPb7gBcwWXCRgKn9FaKN
Sl3mhJhc1HS1ESYGED8XIKnBXK9Lq8FDVy62TKeQRZz+7UeXSK4dnro90xrDWKxdhJhOLMAOvW75
JK/wdl7NiRebCcwlPJEWsRodwcM5MCCjKEQd53hKZSuHnQc7yoVVlw6usKIOE2k7xOsw6JutSCDz
b4frAFH+Rv7ie6C5VMNQSDsT20IdzXZnFG5aeTkJS1CWjlbwhqTV2lPglaQhHOGfU4WL+HiUZ3rV
X5BMR0E+1vgzuuwIiG8DJz8uTGULtz/6xHzAJgReG58eDnKngYCNQbWjahkYhPXEQZ02nxCRd+W1
Wclfr4b0c0k3f/mMWCdsTaOzCUxmFZqVS2y30bzoCX0mNvfDmpeDNPGqH0iugXbGBwQyVgPIAdmK
3pB+tKXXD+JzejbCjduBRBsW/eT+bcKK4HLYf39BhSQN9xD1drVxQM2gwqcTCDP8eHbVyJ5X2tc5
hsvLpmUjw+MKanoqqCHD8HGlQpk3PZ3JSc/cUAxo7ybsusWQJq3F4hg/8lObsKehKhKiLlpIAtBT
VcEY8F78oxdUvYxb5HM0KVaBycoOdXJffZ3qJp8rkNE6P/i63qg/owDyaFJE/fVz26Ok4QNOq5qE
fZoiwQ92I8efCeZ9l5xBaroLsf4crvpLvqPpM3T26d54XGfjd7rHWKLie2yj5tf5G9otKywSj8+q
Wz1RgD4ZFHNbaOpPMubJCgS5fRJdwnN1A+PtzBqqN3bSsgYGv7g3qF4mg0O4qJipSMIlpvMEMROa
gSoI0mumua4eegw97q7bExLJMTKxdMRH/a7kSzN4sxDvYZwisHM5YNc4EsPMEIrn2jaYYRnzUhxR
zrXUw4Gu292nGlHA8BRkJLJPcNuJnSArSlaOY3pNHuWe9wqp28TsZJ9baooCDBeVWfklkc5aER1S
qTi0bUp+d638+LqNQIgfvF6RyLd46sGLAm5zgRmEtKvnGQJGOURtT5ricthlcW/ky9IN8gdglO3N
I8OL+5L9xQJxVmiYM7XIHanibdBqJHcXQmq792WrF0vyOE2qH55wDJtaL2hcK2MxEQ4fUba1rBFu
7cA3Oo+0OkEMqSPsrmx3HNHOafQUcoa+ln6UkJCL8GMkHbz07hlfaUaqGOAkXlcRbo/zH9S/C3jb
D5GpUt6nkBvPngaHfAbIBPQ/fnOkPEW3sJGOkz0dgyiZD/+7EZ6hrtKg8Mt+LNvhg+swwg5RP3rm
8ta+TRGTtNcP7I9ybfaERPuvjCb/Z9uwYMEyyTZGroRwtNTJ0eXm6md2ZQYklXUD2yQx0511V/Se
cLpj3ptRBpJeRJzyVmHu8uiKK3NGkAiwwR8bcAjA8OtecXFnSAyFmu/dgMfhPNyb/g+xvKEFJ3xd
QSWnl+r1/7wSqFirgD+pH6xGUd9hcMkdhrVHeFGXu0B8L5HLwmcL23H2op08hOIaZyGKUcc4NQMI
cxpCuMyZDba0vm6qnqIAzWBW4zx7Qm24fBBS8WE6OxNnznxf098X7w2mI8JmsMmmNRe8Q1EW95Rp
slfy7fG9DptMhH3V04QJO1tYs3p/E9uKXWSyAjFt8JQP4IPexyCBw5Y994jpH/Juz4Njk5156fQW
eds520qlm60hzPLF7404PuBXpujugEDBwWi8l0EcoRu5DnwajjNTIs4l/p9usKwZtmBTt7KBQgbG
U0547PnngmE6sqLzGCQ7L9BFErAqh3Sflvqi0GYgufwgaYhuCKXXZWKWofOMCzmDEeNeOPK37a6b
Ag3RPoT+X+j9K77v8+/i11/meGQ5O3GhYb1MGkJSeT0iWFNpP22lUxFqumU3EkfKWJVpq/fDv44t
SJQpRvgQi+iiiuajtxX9CYOPww9IXAXXQMHb5WDI0za3EYXtxlj5kWPcGP5fBwhHVApxHmoW9ui8
jNnhoEbg/ZIJazqvkHKDa4v8PfjnO7kbiTdUJULUh8sSARLO+wUCOh+bLMApaeRI4JI/0HfojM8s
ayNiAzjWGxpYtfmxs4kNi7T53VhyhJ9TDM09XjABTw0odBm5JYcAoIRZXGiJHR74048QiD0ZcGzj
xLNH5ipqLB+cMB+yNt8FfgzvVwEN+qlf5X3/x0psGxRgca6PkmkYt25th2OpnboJjObstwm8/3Bh
rcPTCIkqYpsHpIoSsTzi/KBZ5hLiwypMq9MfK31vcBmi/giJDO5NzecG9MzPOlyKA59hTECypLvU
uYyqbRVgT9gtHy9qtLYO+GfgAvwR5MFBoL1icl54AhCntocsMCrFC1JNAhx15US2l4GEamO5LB2p
aGjxAfmQD031M7wHMVL3SyIfUqBYHECi2LLS2fpkUfw/xU59Uuj/rfY5ROb8mDYLCVHNEJgpaecY
6j7b05atMOLCZW0U8x+cBClX6ieXvUDhXCT4f7wHY8IHHviCjy02hIESlGbk1qqdjDX4K0jDWUgP
hjzpIIBStjwupyJQqbvbojanlMCmKhGA+jMiIYAVpGHIcRwfSR9UxVXmwFNV+p+EBvJMSm+F4JLI
K0SzrO6rxkB2i8G45kheqgHRSVAC4BDcFqfHsWq0BPm6vYrxPe1CSPqgdcw8zaN8kyS1FRDEEvxV
KXq4ItNQ8x/Cm2nSe33El0cNDGbbeKrZe/ppfgPJggv+c/PmXv4P4lsWFn7dH0IekuaGKwluhaWz
qDD1O9/7uTuC3RyNl7HhDKFk3hPzpLIOadeI2emudCBuIULk18hqTUiemU29adWUBbxM/QDgJmQF
An8+vYOY/xvzIfUAKiS9SB81/kruxe3evHwaZaSrIyiJCz5g4NTdh+eitHzmWpM7RfeFEIavJPUN
t1gdid1g2u+5r+UObBPvCmSs28nQ+Cm4kURZPhYaZoiQAw2f5dKzwHmNSwUMlJBWNrhdLWnH/XRt
+5wUZ5nOcLA2btYDUNzJ3oFTs45sqWmmxW8Jdle/+G/wG2Tg/Zbyt01kbf4WTItAR5mL5GQ5S3AB
8twQaP2IVwUqzO1L3SAVcnc2P4/uY4i+y20IV/VWJLS6TL/4gxDMtIfGsmok6PVxauWYNFU82yp3
aDhVFjAdeBPQiF+hRbLd5kkx81t/SazL4z3lvyDFYLhZ/059OXzR7PsSgpHFNwxcdgELZQUz9a0V
jRc1enRZLMYLiOI/obxa+sEh3vbieU9qHeW4FTWTlap1Fb026gpbGKtoeo1ScgiErL7/q9kS1rbU
B8iR6O0hfu0r4vwscgzmZbeVvyPtOYf4GfUmllFQICyLQaNRrk42Qy6fh9NCLw0VHODSNtikZB+W
c87ZxWusiP0jk88OdwfeT+82naunXEaIj+kij4W7Vq8viZtH1jUVVtK/Mvm12RolvRXkrg41sct6
Lb57hOXle7uBcIB7ZdSLtEDpO7LJr8vxH26icw0xLf5dbbI12PcsNwoaRvC+CoPsHGn+nhY80r5L
bjDNHaUr62oqoQqz5tJKlPbjGWNLJK+75TmGveYouF+TzoSncBWxXlOjNQaTB/dOV2FneFPOTlwM
T7jGDFCi6Fzx3qzKpR/9n0e1YqXKCAyC0NbwTqJyvXoTCFFeDNpvhLKYH4OovWmZunt0kX/1maSc
RingpFQ/b3RqdtkhBuBzmB8rDzCj6s6XaDRln/XTeeUXiJ3ToQLYtbzo3i1poSK5qGKg/7F5BsAr
sA2XjAi1ni72ZZ3aJIO8aaD2X9uP6imjDNID2zlGlSvWWep6QbIKQwR4wgxjkXJBHye1Yv65rSrK
jjQu9JzQauwwXbKI8Fzm4SiTuyfGMHK+/kn7rNi6uXZUmUoAjiZbZj47hPaNCoMGlLWbynJCyfb6
JT72MscqAUZwsBg4SPAOKDJh2M1UaruyxvnWIGiyHino2okoyaY4pjpFEYi6EwJHubAm3OCu7vm3
KlqwoLM108cE0AeN+HSX9VzFLZRaSDLplWOcOqd3JwEejV9SlQeFFlR6xS5i78sbnbHxj22S2NsN
z0HSGMys/ORu8IpS+nKOEVWi8ycl5UAseNrEilcSdAX+ohM3CobbGphazdGLofDvTXidL/LrvDVM
1lutqlcno8MsCoGv+jk6wg0SHe0QsK3h3ZYteMBTsMN3GsJQH5669r7YJXGcBuJoDPdq5EIFeUUz
tgEu6ZijTjLNYeZzFw3cDZzCX3FSMxPtewEvCmszPQ5T9zakkA0+4iZxCZp3ttzBJxwKe1yhpmNY
7ciCJ/EF7SBwAiCLw2/RH/QuFIiMx62v1MXwVIJ+stjv9lMJ3mgfvG34Rhwxzuw/kEtigFjQb3f1
xeyWWxIBlu0YjpfwBzG8h9SgwGFnFuaeVMTNt261oX0Vhd4h9noSJPgjQiGF2vjFQ7cSnO3aWead
JS9/QLGcBVHT6OrPBjiKbZITic/eDAUg5g/czJ48TfUVJHAkEs5tFtCd3ujI+kSZBTUrz2/Dqof0
jwHbKxyXPdcSCtR6DRHdtBhjSwJMf/t5p2QCuRsIZbPr9iFvkEH5413m5vB63pmo8yFA2EnJ2Lxy
nmy3p4yeihO99SUjnfQZWcJOzmiHsXoy3RuUlezVd6Q0dxEpdK9Wmqj9bSVGuaC7I4Aj6I4rJghs
hbzXllm2AEjngfVzgq+8+7ZzynpbVBoZe1cAtkvf8EMhxQ6tTXMxBeY5ncupXUoLoC9sHf9q99cP
rkisu8ikgia3eythBpY/bUlbFkYIO3aDP3Val1nN9E40jE2hEqf5n5LoPsnvHojxo1rBbnOpCDcT
ieEeXiUAehDsMy7AWjZTEWHd3ND13vowT8J/w5uzJNncZ5zKVQaQdb8XwaHEYpbVh/QCj6ug8D3X
8smkO8OlH/+7BTF/MDdXrMC+VhZesbsgrSS0rP+dQR0Pg8/zycBNnl1xi4P5FxWlGa9MV2sTc67A
JQdFgTVVlyHyUc98Pk78fiRMZ7oraY0AQLcmwblS8Bgt6l+dglfE1lz8+IVcZ9H/VwFxF94lHvqE
6Ow6tvjFa/OlQA/Y8KutDhb+QRJfvPn8aEUJXsvpVW3bt7dPf8GVvuFsVINHW7h/1R1H2vdBD1bu
dxMhHYnp5O+b2mMKwak+sHYS6F2B1jUKh0Ic5MQZ0qF1mS1qk50HB7xnKiuVmpIdA7BCu2jfBLsg
6ZQ+jY90Z+GKLpnyRQFXHpLJzjtZnF277fRCGBk2/j+FKQirfJZoVMFPA88rSyswqQdGeQwQ+SAN
aZG/MR0Iae8drKFt16zCDFTbMiUH+cnLUZHsczEX2HJi0/E2B7paj5IE8lKp33rhcxP690JUFMK3
CK/MgEf8WPrvoq+96esMV1B+8nX8b+S5a4kHv67iHjp0uM9RoW5CVRkTDvT16LIP6DWdKt6fmhec
nBWMCYhcCEj2CEEc+yf74C0v+a6dsjilsrH/fBEb+UQoBJZU3YIs+uX8YceNIOa3GBqkodJOpqya
xH+ZGZlWGP6S4kHOB19fvXqKsk6ZzIKuOwGzlBBjD26YMNoCpWgB16nAj2nGLq6bgiNARn4eD152
2wdHCXC1QOP4eAtyQMKfAaTWZsK861btsCOCczhCkgJhAKfZdNmAY6bdIsEgGW64xwwWlksUosvo
Gl5M4Lb4yxa+zwDMpzjEBhK1CyveNx/Iwwh/iZTK6ZGq9/rk+yUdsa4XiebUEjsf/wyqeq/XU1FN
UYQfKPe4SRhuxbRn3I4Bwe47Jjh3aL1y4h/LR2XtPiP1dE0hMOqePZfgzZcKHDYiUK4FsizYhcty
S53Apr4IlsAnKCuTxJ1d+IdE/AHCDlEaAnCJ4MH+MNDinp+N3KQP6vPz6iOQwp6XBWlh+k3p8f+z
kgIxLbMYP+iHyKIuLFp2NBQ2qQMzNVWImWniYb4YYzQQ3xMhvY8qfroqG8rxGZnoguIdBFo8H9b3
cFI0S/eFqzskkGBZGczyC7zhu54nOU2vEifpqg0jcECsJQdiLwYbUrnoxYRAIeu0HK+Nj5EIDznY
F1vHwvbKNrKkAffAivFOvUJWNXid5sqVZgcLXO5mUSYmS3jS8jh68NEsz+fUQa9INiulUYpxyWLZ
PtGAQg7qVfRJTbnJ3GHP857wdbvsUpYrp5rUWUhdv1/aXe+31FSDSccZfK+0jj5IwqCIVC4nWTT0
COQ+HiQ8jKdS4GeZCv59/FT66+LkYTtd+eGL9sJqefKIxvrXuYG4nvcSmjs2sb5qU4hiaJSiGUGf
9mremkrHkVL9JhXcpw/PiizT0ZDgJPS3CZkri8erTDdymWGdl0pLYw8zTK+mzdiJmzKt0XwG7vrf
gCFja+KpZ3E9v20MqcXds/H8eYrsz5f+OqHBfo1cDotBEhzuUMoZDzPkk3V/LQS91ltSN+jGi2oq
r4QYlq2JCRMYS64P0TaPJy/QZ4O2/x0VyAeNdMdQWxLhEO7JnUk5PDtlgRJcC1DyEGjIltzH+mcF
6es6LDgaNUhekM/yVu8jWdOrdke8UQ9QeTyVSYCs6LZ7FKdT6C7fmaJjHbcgA+KRb2Nm+GnCuhRG
6CjalYz3tN40CpEQ/XGY0O0OtYe9AkYoQ9KvCvfmNTp6wHjLSG/b+TE6eKZbbnRm8NnrJ98nVunU
wHY3l2vDGQ7KHLMt9vhyLlVho64ZLqMl9UT8gSUTTauzuzz1kaakr39ROHLFVUB/LOo09zE4F8Bo
1ojepqpeNvg+Jxhgb7wLK+9dU5n5wGu3PFEoaqhZhTk5k1mWLQvt7s+JjRqhvNrCOvQAYoXMHeD5
hEigUQjTZEF+0iol8wMsiApaDYXdZKgg9tj5VJhCrvQccRloEYkgDy5k8u9u9xlXy+A0p8nx5vSy
ICiFeq9MClfoegxhEA3GY0sTZJGrsKioAmrH21qznizc2fgbOIEvQ+TYImRm8JZe89aLAf0GM6ZQ
iWYGomZVuA2evCRoEf+vDK+Ivb25jdNPt5MDCknnCt+KCfTQFtjcZ2HDSOAQtKxs+N8A1uVgxpCT
3xoJjLVQSz0bi+1NrzijTB7MDPPm9dk6UKxQJaeHtBj+XyluWYFv81K90Lzy/XHzo5Pjp1Hc+Ymz
zodzdkTFnOnhpjMLv592i4cByR1b2ah9tCMTZ7UwVEGqzHivB8tpOPT5YzXj+YDajLZ6e9pzsZnh
4LBZ+j4DVvKzgv2QG6PYZYSnOQwFEfUyRs3au8X5DfaZL8DwyPzXgaJLkZFb8YLaqNxWO0o9qzGA
o023Aqll4mIhJNYBkBBNpK/pGGP6Q8tgq3r0jrkOEYl9PK8um/MELBxQkBmfmilAhiKS/QdSafr8
ilRTEiYiF96gckS4N8PAKUXlgi3weY+9FkxMN5Uz8TQLPJj0NnUGZhHnK2lpkyAktIebFJoqurgB
2IUM/bX50HiDti5i8gOKam9cPdcsUoy/ktQySV6tPYq8PXWzvkWIQFBlRVK1oZhofYti+bEhs8os
6PzQbuzJttSzHXjREtNS3YeARXapTv/LGGh0NknfRYo4GIkmQHcxrxt0sDSzs0NqiMGclnz/lg0j
yBmUONbuajicrSPCYY6V6KpEHw5JnDPW1Pbmemgt74OZMP+sWlWPNbYg0LWBawlmQhCcXmZnp8xR
TZdQW1VE95GsaL3GfgCPbVS5ppY47XEoFtp8PxeTrnH63N2rwUVwFcoAUGkCDYO+zRlxjzKMtS8a
0pZuZJn+eSi4Nq/EopnD3rdtLe5RKy8xTNQIn0tptFeSrV6kNwHLfHw8PFGd03B54yFX3kSLKMdd
D/84TXEgS/nBO/7YbjLYfY+jStHzS4L61R24nRfLyB7bwuV7A9OQ4CPWkYOafmlIVuTAOTQmpdRL
+UDwgge3IscwoYQfipugy5eKvjq56vdY0ofBHdhQdeIC6ui/+IvA23JmjektFxhZL5tT3WMtTNM9
xvZqcUTwX4YFvKR0GeZ8o0RAhWWT5ineeVCcbwb50CtuhFslbNrtzib3/rdswS8/YfuS+ePW4Q8V
O/xeS/1lkozgBwbp94D1g84f1xSQXqnilpQGbJtxS66i5CyzBHBahSF5WbVb9YNwn4RVh0f0QMxL
3rWP3X24/7U+cMxDptEf/NNud0HhIw8QPjeF+eje8SELmzi4oytvTEU5a6ZGLU3+mewm+FDjaRtM
v+bwiLSgQWGzRbA6lAROXLC9ZX7d8fpeyOfJKnhCVzmutNAmhP3XFYF3HHL4rIRFT4EcOSRlzew0
ocGw4z6V+0UmTFMMz2Ru5ERxY9u4pj3QuGElqB6YgyFBfMuEOurdWCimWZInJiympcQnMbA5Ul5J
ATMhP4zGgdsVxm0+0vyK3CZpAZg74Jvt6qjW6zTGkPl7rJ0TBoff8VdzRTovBWxZ0sWso670xW6L
ca+r4CF4WlwStqSqm+1E9kKDgTrb03xM3MqqjbNXcEOBE4cR6X8y6vNyAAiPa9cZ09ORccWK8rdO
PHRwPrpWl5jloC1ALjQOAHdTpG23MEOs3bNDDZfFXwP35DPiWN/zpDE768N7VKFPwqppjF91rGZH
87i/Vu9zpaSemo7YS/dNL3WBi1d3CJTv+d5e+B21a0paQWkvLRAkGbTSHWODCzBEc9Uk+wVP2evQ
fAkd29wOTFvlVhRm0ceZyzjYgkn75hv8H1nzHHjs7rF6FONOj1AJwSXhBsZARadTAWHcQKUHAhIy
pF37b2G0EyMXd+E1iD54ejezYuPe+LVCMf6/EQ4Rv2d9Ntbnbxi5E14e/1HIhO1OjDIYlU+EMjGg
RhrM7nmCIMqqokgblBzlq8oHa4+Rf2WuHBo3g2qUh8BdsoATSupIHZOA3BEZGD5fFaoFbDOTybj1
D7Y+lD7h3mqe9O8uj5mEpryDkHBQ0wCcVmUs1QMvcnGX8fU0eNmhqC3VCEZuduw/YRaiSqVXedrW
cvw1gt2VsTNnwUsY26XS4e1KF20NUMAkAqx+ZH/1xwgs0N5bjFtlQryGAjRNcjykZxXvN5LwytXh
QaXOMBAfFuPXRI5X3GfTplG91zblZdpJC3fcV1Zt5CmLhmycoV77DS369ZNH1tFCF6L6JKqulxty
ThivCGRjwa39ZzdtDDaaTv1ChzQW/N+1L6Y8dN3LVNcgHbjbP6vDkjES48tKIDCdVC4xIbQGB6uR
5iNOvlvueVczYg+MfhLmH5vNTg0Jzqz9NBNbSUZe/yBqHoEG3awybVBW66cF/VOLZmQ3zj6nCwMY
dBabS/fZhE/R4nKaYf0nfQc4fNi0bgN/zuoeYv5YGzSfigxqX/r1XEbCjuqlq7szWQ2mqfzrZaTF
Z5LEGE5oHeKsufDtEY4aJEDlvK1QeMQpORpijxFVB0SUxRykvyrjJNEepHSXYQB5jksqdaiFzUv9
ELZW+PAdDDR6+J3Jqend0Be8C/0jYQ96VSWyjG91gv2R1co/8jNfa54gNHjbKWpKIB1n7x1KXmOC
74s2Zi70hv+pXxjsFzFwkh9gOOriHFMgTOkNBFgXmqcfpuJGcR3+24u48ZC+GTejbAfT0VyYfXyR
rC4i20rjhFXvOngPz8leIG+Fd3GMHBeofxlOvoQ7DpMt9VCebMwi20/CoOzVvhc8kQ1WmZANW+rX
qLw07XpsIwU+B0iqIV2QaPJxTAs9rUtQc216FmsTV7gA1t2KfIcckaSG58c3Nh387TyxKlDMcuhE
YwG6vGQY9Id6fZaFecWpF8qr5AS0IlQJKkJswgQ8eG7+wFyWN/ktbOtxBKwKsA5vDqna37RgNZJr
cGAOLZudYjcyi7Nnlp3QKo5JVd8JTw1Mhn44vJjpZnc0rne8vxeENB2KPHlXUAFqoe89Wj6Td1Ti
9ZTRT5srn+xkh2lZNOVhjZwIyU1ToVkoL4tuHcv7iaMTzbM0UB2TjPwgdbUmNbu0dWg89e5XeMZz
nejiOXIcvT3CnzM6NxlXMsMDDzLI/jF268IXNxai27ji5VBNHiUwwR2wH2b5AjFjA1x/TBiHfS/8
6AWrwd9G8AgFP+K+3bp1zO3fGwvf5HPus6Y55hooDOCUvUQLMcH+tO/zLmvIqFc06c4273eybd3j
gNKgGg5ZV0HJUwwQMVi8MvhxXIG7aKY/LSiMUeBkr7QLzwO7xG5PK1IlWCHV6FaPlgfGrrAY7Th6
pF2sJ59ANUwvVFLc/2r7poG8XeLuosAU1AfspaZ7O+M5oTEjpLuP24UqaKoBS+3G+40c09ppNrS/
FF+ayKVJ9WwoaQjo59AFZDByzcQgcEZnT6jMlcVflW2WQQl95UA0aMCdeSFgNSfA/EHDQFNj7NIE
bbUK3EqRJbXzwp4hKbb0tKThmSKtbDSogqSm9vPt/jRrmnjaporQH4PwPGbDlDyBJlCf1hJYHjSO
yhNsh77DZz8AnfCJFDshDjVRYxxt8SRk7EeBgHEsxGEjakQj3Oa3Y+yMFcZ146pBBHJzJuQVNMij
/Q1up9pJwT1jwyVwg3D1kM0m+LMwFeGH9eCslOKjQbhJUeubR3iED9+gK+IfbQ71h5ACJRPgKqaZ
6TiUmprL+HSYnlCG0QKwaeopYiIYAcNgoejeyA+oca5/Yhsa3Zw9ecoMZD+kc6uHbsksbtpmlPtA
mjGnExfrDQ956zC7/10ri4MuEf/FlU80CfqUXtpPhseNTj4yfxZHqGpQYrCdwIJjuYIB0vZDJHix
XynsPDvPOIZSUfe/hibSF1kgzwt/tCfhiKUo0YtjD9Gy9yfYz/AmPS0hUzWAEtHY8b1Lawm4Ds4a
mOqsa5yj1+Fmr6elRh0HidHAIAGMXngy5DsGZyZPhQDEsUyxyhcXzQu5CxLzioib+ZGTvkmFhnFH
DJLUl6+31nyxhAEyXW491JhHpV5dreWbyc748pxHhjbAt8maFcLCI9YxzVv8cAw2YfV+inyGcTrr
zUOfzjV7TQ7hKZ/0BLDxX9uTTnypTdeT7cgCpOg2OmPMqCd5TdA8kLW3cbaqljf6URvXYwfxYMdR
UspHfGud+vZBHzlBdZW5sRS1iGt/tvsF4aLDDf+VQXr5flrIb2bwH/RPPGUebBvSx1xopjT7YXXM
iZWkcV+UUc5iUzyxe/LU8Epc4NdTlYjdy2CdGS9uYoaT+lHynN5ucQO02Iz6mWi8oPEanWKCmbOq
pw2qCDyrM/W8/225ym7KpN5GL5GuVsyD5yA+wz6mM9s80k2A15HdDvqK4Y9gHOV7LRqEnSx9WWjh
1mQjMU/ynPa6fmoW2lCH11CfNfGPZNBb78R/Ll9FJrCHmu2mAOs2lR4NPvWZ/WYz2wOtDo4Ro17e
fP9QJ9Ec3qdR6Gg/Uxh58tcKyAJ7by2DqUTzauI0PkaJlTdIYp6+1CjokiOBVmT7OqVVZAi3k0yt
vqyn3XpbI2CZEdgjQZi9LEHtphKBh/dXEYTyJCllrtJrl2Zw+osrMmKJyBiUNXpUd1Rz17LcD166
5pph5NJuHy5KNEQNvcE99pUTVPPgnmbU2pKtkPDhjBbOmTj1cJBj9dfik7V8EZ+epZnuFQHt1kll
jBnE4nv4HngIW2dbfUql2+LsK74axShxu89kNo+X/HBYtNZVHKwD4dDTqmgHYLKEHMYEV/iSiJpW
eT4hIOMLqLHi1ognlw7KiDrXldhBoh8rcy2xgfCqfYh3x8uAuH1ff/QBSv9oCyUIh2teypEvY5ie
YimVM3i+BHz2C2ZmJcGqmarQpCFJICWAtx83803MWsG25Wd8k5lm38mG4xGg5NJssG6l3SK4BuN+
Df67TO9dWyg9eom1GUlMfaLblK4TtRXwEK9LOmuNCFOKXs7DZC9nidvz7yIV9G1Axlg5OBO95ww4
aToHnRzeMdzQphDaQRgRjaiSnnvY3ZVVV2qAYZTm0p7PZO3VLmuXAlGjfeILBR2kB27NtB9IYHWO
M6j/ZM1MsvzhuJmzlxbqo7a3MdH2qgdviL2GjqMBOr/F83TKOHeg/9YKe9idsw3YBC3p0znNZtAC
UGSSAAyNSKgz3hu67gwhBBtk/DkJqesI36E3b5oO34oHxqpwWjDGhDR9TNIdThSFGILRC+H6DirG
f+4kh521hPtpDMjPTJF/ftIMPPhm9ghf6SR0YJ2+WjVs39FjDrQpwptgl0hKiOJWUYNIJCCfsiOx
j222EHW/5LDfyO7O1CJXUVaqQ8ceiTxjcOd0lDVYlr07cEu7dh65MMFab0WvRO3KdY9Gfk1IXzmK
hMpcS/FbDoVd8GClIFaNvIxb/t+DE5mSU++QyS+BTvdCkqKnzTADomPtcJvWz4LtyFb3LirdGzeN
5EQKchywuTah0ey+UE3fZV1S0gSO9uVfe2hTv94/ld6QtpdgQ9V9PvhbdmC5jSryG1YH27nVyMuD
ZlatQGS8oNCFjPdAuids04SwCaOzWM+GxkY2PpvJ9bQeeSUBzKjB/LuxdnY9dkQYndqh8GbB2zC7
VH2f4jnu22ezDzEMpLFdd20jpOPwKRWahAawOytOARpRyj8qlXQkTX4Cj9xbRoJJYxNkKyFuAx2W
PRQkp7MAz4Do7HJpj8TxTK3gHk1DTKm0NJDQm+oLO8MQ/LPN/qSwEQ5lFGwfAuFNLqNIM3VtU9il
xL7s7vWF/aKPVNA7dmTtkiaF4SbUC878ZiKLROrRuJikP3bSmbZ4/W2RHQcn0GY7guDTb01p1ZF9
8Jiq0ZwCX6o50YXQLrdjh/un5XgX+I5s8iF49EL+STqhOjhsFloV3EGe0xyfwVoqr6v1CDO6pq3z
ynRF7ovT3/4ideE3Tgrsfvv+s2Lj3+OoUfWvDOI2zdaz6VOB56zbAsGXxtURXoC7a/eOVRBwKddn
OXSD55qeXg0eUdHq1es5umm2r2xOAxeZu1SgPCGYHqfzedO9H0G8BLM5vUQFWPAkutu8EAMuPg3N
b2YclXNuAdop7f+eRvjmyf/fZ5XBNMx92Vsy9QPTQQMsqa7w8YBu5/uhuHU71NS3kiEzI7jb8fkM
Q+hmnc1KRiVlGkNWmqF6uzRaOKR0xm+wX9QZhBav8lyfStmduTr0ch7iDSNlztsbxiQXzM8gfT2n
Lyy6wfFigYBh95mmH9k5F7VVGGTTdWwCe55K5yju7PAuB/sVz7+Xx63G6IYzNMZ2y8OGQ076fjHl
6KMci8mcSnhuJlO8+muVvTUUUe7FrWwKgGhAk/3NbyKMEsCrYKmiP6DIWjBEeLmb4Rk82WWJSLFv
tfnLzRx27rylK8DI9Eljd4e970SJodVlfy2pkQhQZEfW0LLjGEjMQkDPhWlAyQ5lKy8ToplW/5Ze
Y4b0s+pew7WqymIgXf2ieWAy55vcgtfTJRlOtNtBFeCMT/DKzskIAYvHMj+Y9DDYDlTGRK1+F08k
qbzL014+R/FZbw8ZtwaforJNimDflzDfTPhP8VXnMgXU6aEQRwFd9Wglva/p3VjCInpUlRLzhS3t
H2Ekacy16W2F6bDXBLRBAZ7Ojnuae1pQL7kgCk4y9wMnEDhrsML+auOX3ihQmwD2wwmOGnDQ1MgM
1IFYrOiGySnh+nFyrU7U1oP0vXem1Rgc6VhkutbXcxTvSAExqOlJK2po6VT+JGy+iuyMoOnB0ryN
/AHklcS4iFgONxwBITPaUDs3f4qGqO6YdtZVJ3v2Um9AYTNmTpfiTc6A5R8LWbISl5eWQ42QPcHw
vPiIhSvb1Vc7ylcTyC/qeaBlgxgM1tDgZUCgu4S2T/B6wejTZCfCHnbAz99hAbCP5vshIAU6zI//
tN/Sx9KiLG8I1UgmN65Of8p0l+ggJcyUnahNMqZA7BVB3kjR168C8foSMYygefEb4DxNhbsd7NAP
yYceY2WfkH8LXQ8pqoDL0oRmd6mG8wOQ6cKTwm9cu2H8J0nKXLXht01OMjRv2711y8uf9PDSbn3z
zrr4KYNuocNBVrZPuye7cmsBIhAIutu9EIIp/NETVOwXRx8wSxoVMArZ3twUybK77J/mLqhay84x
mVsbF2G7ruTzeaOi7EB1+PDXge3mrlQSPjWQe5h8GdJqT5LPEJwzNIgYRM68o3y7VInkZRV2iwNA
mMl0srpWpMb1RgqnLOV4E6NmznXHWOfbqmFygrOEq9LAQlRCvvN7wE5kptUoDCGGLpqluhn9bY9S
HnuXppcMQqk6X9NydWRYriNsEBcFW8DibxL2GR1kxdcEYtM1n/rW6rHJMmNcvT1DsCtasDFpXTsV
Y6OoGVKTWNysDDGvmwsfWAFifo+psbJ0I8bndU/jUM47bX9QOyfEpm7XeCCA3AQwtjOsU+NarKps
V+P4LUHM83XZUXUjZ4UtQRglbJnPlfVoBFg6FOF+fZX1BMXV4KpHKmRfjKnX95PayrpA56DbHjSp
n5XsfCMQfeymzWZMR5cEGcPg7AjUKAqfFYAfoPZNYOS2ZHvV6A5KJKbhRusT/EcXKtp7XPo48nIM
LWgJ030OgyFCQ0JGwq4K2USx7iF+HIyeNrh30rPPFxFEN4XXaME9S1XwEDsNTH8nbjHEGKF2CLQe
7ltuzO4AckkQbhxO0U2aRolO8pqz4ljFH+lz+zDAhatYA7PwKpQp3lncG25+/72abxfQmYEbcERX
+e5vBDKb6jzYz53kGrINett5D3u7uW9inxZzCtJ1gjb0473YJ40oGT8+PLFDlc0JVKLKNG/Wb6Uy
NjOnWvqKdpz7X7pLJUBkPil5dWpRQz4+bwwvMiXvvVh0U/LVmdV522WwZFeBN7eib+zu1m1evbu9
LJ8zS/SVicrr3x9rJBj30/dse63tTlDzmUdn0IhEiZ/3Yuf4LT4P7M+vWJrla/kMA/W1gKTiY+Lm
4yEmIg2EDVpio6Go/EwlffqnNVbnLFA4KXxVAFQ8ytxt/WgKbwPMa4+V2fo+ViUOLtVPSEoIW/rN
L+b64WxeKLtabGiqmFIsUqJ8TrAYyVI00+UuGUO8BQNBLbUhzXHTO6CdxHa/WubAQOoulVZWdQeO
qXAhI/DgocuHioRN0eTq8H8SMSrrxUSmRrQostZ8GCbEbEUJVjk3iiW0SHXQpyHSW9OG9ulvHSig
/LyKKihfGCM0Jsc0LHEOaX+tFch46G/b98aaM6l1YSednXFIiH00Ob4qPPJk6VlfWP3jsNqgSrwr
pods/1b8wH3/A7bwpz3BsZkRNeAuRBgpXnLAhv16HWUO39AYxOut2rhMOpKqGBH+++/P4SpVRl9C
Gi8tEaSiKFJ9tBhtn3aRgJ1ZaFfVAvgYn7PQo53c7eNXQjqFPKj4u4qMR6t45nZO54FBdraNAxRa
PLhe+kfVmwn9/ibtfs6zNqSSoyY1rD2GaB/uznSXu7YoydbyrsTOsUI1F4yQjGvcRgZsYN9ZQqNn
QKiD9GTjv3GBnXdXvwAX7TI1sFVRXPrURa4kLdin+apINzy7MMUgT7kkmto4NfSB9evGur3f5+Ai
u2ocXIOWfPer6eBtYtMW4ml1Fs0d69ArluM1zAX324n1pId7ciDcnB2WoyWUhuME8/jNFiEHjoOJ
Ry3RL7Fj1cJ1iTS94d7YC2beT9NSRNosqR0zxxa05dMozsUqJ8RFTHYAB/hIKlzMf2nDBkFSt3yZ
YZM3RSG2lc1O94PHrBzqysmupya/eH/m5uEAGlva2Hz+Ptn4LI+ngx2n5EKNOIY52vu7sAEwWjqd
Yl+CPDnAJ9RFOUfcanmWS/EmK1SbjR30ynpnhdAWFj/3IyZmlSGHsd85rQjFrDEwsjJ1bG4xpfDb
i9q2FNDRJVmd9HWzTXuIVN5LCgG4YxanOc8GJuPClmH6/DdkUhbRXBXtMDtP9gbyRre8XuTp0fgm
NgPLJwGgVrmN7VIuc7ZeACAlc5RseSgnZOCKNJu/WeXO4h4XzFrfPmu6CwuDcFTitHJmcLTVjlH9
Z3OXlGfEXQ8EeyfHQsgLOPpZLsZddRt6VLsZve7b+7GVzwzxWI8UB28wLTtVmBoQwyS6PVVWrxOt
XiLMDrI63RVWfUO25Bb95iGeNW6qgRLF1yD8WVpCaIJhVRbB4GZGM1H2f9omBHmxUx0GThMECKP8
y5Xuk+gIeGnH5ZlZG7yczYztTayjbTv7spGN5s04L5GmAhCgXT9Cb62IWpDaugQPLH+SCwGe3+5d
hvo2zW7LCXv3UhBR/TnVj9HGOghVAFjkvYJ/Xl0q830Ap4U4T8/WtWlzESFMpNNiRNokNoAcKmeg
Brp2ahteH/EauJh9K8ra98RKy7Od5jXCZk/hT88TxZlBUGkQBaDvBnXqrSIV+kiknb5oYYTJ2a2v
HPQ7OB3tgX+JaFa6ztpeUYpHM7WGGbM1fguv3NJtOh/zUF95f+IPrbkMabQK+bymbajETB7VAOyl
f30XcRckkrftBZ83XWyngXi7xV2v1vKQcUglDFwyQ/k1JaPFVHnuRhDtDPejFEfL4Rw04il8Cuv+
Llw5hvZQsEW8j6GJ/gtSfqQ5HRZn5KNWCnfIO1g1K6c3Jmf62H6oNAK0zu33kShuxd8WbCIh//eQ
AlBZYY7z/RciFREPumnZS+NFKEDi6HElS3HZm9NC0T20r5OMSuDJmh2JC2sgU2Tx3bwt0qZM0A6j
qTMldd1KIAveUKrMiy3Wa0crDuIgMF0EPDyvbx6RNttTRT4vMmsUGd2dgWhWk+PLLYOZOLdyFm4C
KI8MOnPx9xNH1Kkz/hcgFCnY9UeS7iOeT8arQdL1y4y7mZXtra/CsKpFPmMvzJgvbFTgJUlkAwv7
+83JcmAEk+nY9975LL6wcvOglnrZDUbICmYL10Lnk9wR3nlJwc6rZj7i90weV215Rwn1dzVTRVZB
qexUEkpAIUD9jJtfUOqS+Cwbcfu/6Thn6XtCfLL3JILqHs2jHptCPDKchXzLsb7ZSvcwgc3Gskcf
71BbtmZjhubYDRhYj5pENbEiy4j2UbxIIgkaTV3/F0E6ESGOhpT4oj+cWjDx2j+TJI+erpowT0J5
lzyK9l2i7vkTLxyMkTAjuxLtVWTGMAnuaVw6iF2St4OKR+oJclLKKFzCZoOB/pc4JoPWTWFBsgEq
dknWcVurFrL0SyjzzEbJeThXYRDfAA5e6mk1IEcK17zszLTFrsr9Px7SkJv79m/lXMwZUFoq94P/
/ENGvljPP/BnymGunuhd6YBE+J+TZVqLH8PYWetvNIu4dQ77nXCLkheyyh2c82CD5vXWKChTvaxj
zVXHgy7J479aAOOMx484eFDdanPopv0U/NUc0qPfzfolKHQ4MavCGP8SAuzTNCiV2o+2zikyL8Dt
FTz5A8enWJ06/G5DS3lOWj6TFuYGbXYkTZkNlSsp9k0Cp4a6dOQ4ZQ18tOi0PHKjzuXK3xhgTsFw
d0Y5hbcbEr5f0z/rPBnNjX9QNEHtzf+DVaHwGUEOSeFKxgKuUEpg2qHof8uBJbi/E1QlMwkre9z/
Ft+BgD6q9gDUBnRPAEEPKmk2i3mNg3a+vx/hISV/kSxDAQgS/rsgZQTdmTjcwnbNZmgu0LVZOknB
8jPlim9+01CQ+PQrM3Xby1CCUCY6zIIF+hky5HoluDSJIPcfQkjxy1lI1ZcFry/hUNwmjXWKn93A
2enLJ321DHGmphGhJ5ojlBaMbuJ/hu0UQRzloXZDq6fWiKHjLyF/BZ8C2/riNB+lD4fhqO+i8eN8
aoIJH1GBoD6Waeu8ai9Cf7vo1FAbap8H9LfFJUv7ki9BgezItPxh2NYq/c+g9cluZ9UdukrDNusZ
eTheDO/1yRYZlOHGCSYtgsq+OkJHXFLxBExnpk/aw+y1eR+TsGhUwAIlPZUxiRr6iYDKUesolFtO
AAvLVNX9p4BJmVKKNWOzECCrsHSRosuFaDgNt1H7P2Rpm6pWJ8dsibjmnciT9qCnvyJvQpGuGIYx
zsD+UK7Z9nC0zdSFosLe7IFDPDA7aucPFy0oV5rwaTOeukUlADtLAF5tjVluMqVOJt3oVgEn+pRH
7bVMrjn9B3BS877VvI+kSEfzifV3P3C8KBG/WUgRw7m4nMPvq1drhHV8TBQpXXZPvdNsiWIMdUJo
pd93ksPGXu1q+N6SSRS8xPBB7AL/so3O3MPaw5YspkLJrwURgrWaHDOmIT8EwXXRSG9mD7FFjebM
HipRjHK2fQDW2ugk90WjfOCR2TgsGLsuYJ65WgzIqUwsHh6bYVp1s9Ogu36JGcY+YUDQ8nZvsu3e
5h7EJ73irKY9VqOUBa2xvnyuz5wKnOw5XC58RotpXmkapTvk7cSmwAxkkPgoQcjk6beyGpDU8BDn
2GbVfHkbBZzCCjpbGQt/hRM7Q+MFa8hfSPZfASS8Xf2eQkKrP0BYg6jts9YdlfUqNwkYxLweOC3I
+O3tul2DibkTKz0unJHmFy663ethPOcn8TXAkjubXvgAyNs4ndPJWdSi/5nkyI4fECoJVgTHXA1a
VXLNbQ+W3zBJejpMpz+obb9R4ue2IlnnPIw3ABCcE9feh1LaCImQ1Xr42lrBKsAaSis3CMpe8ber
jQrbDrstczg9OcF5Z5L+wZgSF088VxPExMHv07CupGVYl62n4Dq93T17KVOf4Dee8MRzMClbdEA0
CxF8BbdgZzqpB+YpAFgwjpQYPKrmWe2ZLLzZ6tqSVycADpbnV3L2nWNg9tF39jLPFoEVDLDlifNi
WOToYJ3nh/GzYWtt/M8soXlAMj/PFraEzLpiFVl5uBNuL2lFwa6fHEo6CsCN+GNSUgkfLHEpKXJq
tQRiXKDgw5RLi/8E4YODfjIc9bcn4gjBOogssKGsckgPdgNb4wvJ/7EWK2MM5nz00iU7XOT6kXow
qttHy03afk6SiCPJFyFTo0ADneJdXgyv34YG9W1062wRyeUk5kp2ebWrJVDVtefm7cM3bAs8ehnW
8KyFKG4aOVUTHN+2vuvl8vfVXY4JlA0C1hO6kHr26ys9oAJHys/rn3Mbd7D3u031Qkb42ZkgbaYW
fAZcWuaAxm06Aa9GLXoTsw47arxcBQLDSCYJQvZey/R9shvWMnp3yANa/lT3pRvQPGAeLRLXuNAU
SMxqbrusvQ793R/U3DkGua3KSb3p4RilLD9M7edKcZXgWaWdeAWlGrvctCS61i0shazxbQFMDU4a
0UFr38U59i4tUTvY4eV/Teh7zIG6Q00lYDV+i5LJa1hLD4//CQ1AZMJdJTOUvUOBa+Yh8gU2s2DY
HN/ZW4Cb+NoDIVtHPE32nZWtKfr3CnICGw9l+b05vcABfkH4GSisdFJxvH+H12CLz1wr/g4nBA1U
gWGIqeQwOO2OP9Ai4qUJ6YtMburSMKOEzsW24pbciBtSykwrbFjPLsl6dt79kcAAwOr1nUeM8f6G
2vBnkmn2UMcH44XQBbwS+zW32hd9EUUiOBIBBCXUFHDUAWCmmAW6PkCN4w37QkQ/ERTUzpfc4xrp
xnRWNZghtWs6HLAUNUEZM7irG9oO2eYY9fObSwR5sBJsLrnQMnTh55F0Nygwn0LtSNMDG17e6EKS
kJ+7YL9z3KUwqF9LZWp8JPynvJjgEy9HzzOOO7aH7Bofp7ra6YcjwaAdEV6TVf94rX5CbNuYwvpY
aIXoRJmu4T3U/SNuIER0yiDQU++MPSiqu83sxHl6KJddzSN9yZG9xdcZJA3f+hH/UmeBGlmFlUqj
UqteBWkwXfwbaYpW8hbLpnNJLM0H9iGmfm+rUyZIh5+8RnnsfbhWsHz/oHIX5N9+13AaxRq1EqmK
RPiy9bfs35+D7bmB++eJTLc7jEUcdovcnMaWTW4+cAv3fH5T15b5KJehbnm7Mejd82zqc4GNHMzI
X3ZEiAJReQbI7EVIvRJBMsQnkbugF7Uf5b0qagAKH0DzlMH/uxs5u4iRrBqdV+dIdGppOAvFdZLa
CYEI8zCprUHTtguDwllKR91EDVnXcfReU1O6KClsS2yNmCCP9ZUv7pELlJnc8iFD8709XFRs5HXu
M9ZNjKG7+4FAEduhBPkZF3LqWTkz971vHUkDiJV1gt/nKyOY39YFneJOAFHviSpkvybIT87Vl0XW
FXktOFulVIzicijF/7GsOdgd5XsdgYnK19q42ylDMAPt0bhpEPEM+Tyl0GfqEPm0UOm52Vyr7Kns
cka2Py3xdSzLK0upQIEFd8/2p5+nfEqgQAhH54gQ1+/5SqLUleJkhjYh0Q9BCSNTtMMN4UjsM761
ZsEXbu02783VgnwDGKmlqiZTo9nPO1GkyS+gjlwbFzVj8JYV7Dbs5IOIMx/MvkJmQzeZdEDEr88M
GZdeCH2xQOhrkuwqaidzsZkPNmAhJWhlx8mwhy1JP45QTophpKY07K8YaN7L39rfJzrKMyY1p/pV
Z0oB47SpSDO1wENziELG9/SKUx21MNtySNSaRQ9SvV6C7pTV9v2qVkekv3fLMwIqvgYHne2qy0Bq
nK7gibU+KP3I3MbajpMmr/d4HPkiCVPSvKnix2P5MqU+rPsj9fVEGHU6xURzTB9bNdekx+TXAz8x
yoGp48gTl+g1Q5Kc5YEG5ZjAzTeYJ9fBXmtJ5sv4JsYhhCXcEAQwXfnneY7WBEUcrFkLltzu9nXv
dyj1ymZMS2Al5/HqPrCCGKZb8UceyAsVLcZnbOezjFktis6dd3Mb6hl1ZTHreHXwlwuk1loC9x6E
Aamz/w0ERH569VAVH/BpaJpiTAywpJvSWtXH+PGTkVmM6fwbQI6GSljPQLK3HMU1R5s1U1DuVOK1
eqkYGnrhbJDprHhsTLWha/vo+nq+sHTaJb9zh6F9BaLRiy0WxmXJICmgPXOtrXeDKZX4NBDmIoCC
ZzZcKKKCeBkrWWc2QHZ55/8mN60l/mBBE2G1BSjMjFHn3I3P40l9A/4bMgDFIyo68cdUOjBdIUqG
AGTGj58Uu5YoX2YPHgiCHZvI1SmwSuUsoWnBwSm13NVF/U6GcQLVbYo++iL+exlq7Ijpkw+NGk5/
IsskRp/rKRoF7d/cLfTsq69S8vvLFqUqq2lznnbDtUyGni4GuOQ1eagpFffov75BtxUfxy4/Ksll
mDcQa7d/FQ1JX2lfd+0f5vZGcWJTSG6RTkPZm2vX1ngiSYw193TpWvWR3mOmJzE6UWf2Uxoa1KUo
yxpBxIby2RKjgqEOjxWybDrXsJ5aEByS9jWMSEuqtdDgYTbBFKj+VX9juQU0ZnH5LeJFHAzICffI
8eUhuOk+8QaIk185NSWLkMEkSpbotIMVFGRiZ9YKMeMBykOwRxcMO6FEoIujmMraS+VjyYwVlxHN
BHolFNH3563ATUFMslmlFneLFdYJ38l3eiX6U/mRASUMnwN2TDZN956ZkrNTSK6oltXD9UxbpB0I
GQw3RLJhWYRX94FOHoFlvPgYPi/+W39R3yBqVSNjf8ZKai3D1X13nH2m2EqUbp/qqcbZtkAZLvIV
Kz1GQrK/VMvrzdeyB7b8CrzbAtUemt/Yfv0+8k9KFZIUxuHjFL8T5P4a/Vz+Kq8GLxkTeqTEa6eG
4HJ6tsMz/OZomZ+oLYGF6cJQKeZ8GDTTmgjSI87ekSpNQA0C8mUmH9YH7Cap/k0SSZq31WEwlCIg
0w5jMLpJpWHFZgL6VRrTrTdYKc49wP6jkZwi52Q45Qd20DhU3QawdYfSzMrKfG92NmgIGs861uP1
rSe7yRNcyPz+FNbsrg6XmGoGYpBphyiDc8O2dwX4tOY9cnY7TebGfJVCxR2OVccpHVLdh30MnM5s
xVoUEJfmgj29e74zQxB0Cw/h10uOuF2AJsvCCXzZxcZ083TOn+rcIJ4YjXt4Y4il0nbfoZbTHzJe
Mnwn+u75z/yPwf2HrRwJR6Y9W6h4di5HKAHHdrqzh9uy3WBWTBTZsQeIX2eL0cdbdCiTIYCYHJ9r
ezc/28byr2GHHnazXH6js1BXwly06VHtTsjDkhCNTkdZxq0LO9LE1WFFdfOZhrBQHprBnfaIhRmx
AOfN7NlIaUP10pjVEIUQZ7UTbz9ABSotHARUPyxgT05j1Bu6zFGfj4YvMpXjHHYoj+6CiLdjiMWd
hbDvTFnbWzhhoD+/2r2VBaEVT24uuFaZZKzZVzhbo1he102YXHQckLTnMH/DJoMNUOLOLU36Fs4u
x1E3eg9zd3OpiryUAqyvvGEEdsMhEn0WtDk3gxYXOnhuM/5fy58SNvY73XGL52kSyExRLh7DjNd3
FwG69WZprEYwcWKfiLqYx45s884rNoNuxyrRZG8Gf/Z4NJLnsQKZvQqcOrut2aGULQrGKJZycs/+
XvmS4ehYve43NHbThhQPz+66I00r/k8z42lr0O6KljuA5Lp6CY2BDrUUV8GDTyeh6H1bIfD8xmg/
wu8voeS7d/+ZVU1lVEX14AEVBjCnNhyvGF1sCp+Lu0UFcm1msNEuL96itiVpKg2hG73cgBIPgj2K
CvEr2SzeBx0tCNQ4iBXpkKJuyIcPW+yg1KWIxxLBFgMmFzdGrB2cYmRZeQPV82f1SHbHYkgPRIQR
fl2DfK0CT+UctqxrdouqOFiocRPCCyfu1JnIOHUOmshDOHgXIT2lcl6up1vFG9Q6PsC35TNQPq3X
D7tNPYtGMKV4yAsv+Fd6wHvI56sNyH1EqgXy9xg1cmOPTB62vbIPqflMypEUij1PTIi9eJo3kdWw
IsCyDiQifnYDYrm7sjVIwp0PvFbeb5fhdlx7fQTGP4SuxNMudccDrM9vljJwoT8ZFDqmpX7k33dt
RC6dTFKYRXZDP2HeWUQowhel1i1UgZTmNiS1AGdhmgkvTEG7hWGPLOpSUgnkAOmCumKOuFb4/tZG
cjBSOIqn22gMu8gMDMXiVxJROUuxpalRefvq8UHBxhoK5na/S8oMj+L1DmsXr9oGqmRRNq+hslUs
UxiSSaUGlHKcHsMG1wavW/rAQC4iSeb/eKFw1oWkegnunyo5BR0QKOCqtYGThHhxGaQNuS2S3iNe
pmnP798UsPPMU2xGuV/pCpcurDFkMSNKVVq96CSzkWscPp8+CG+7ckos50UhkOWY4kIiODfRrxFv
36gcpcqYryUCNPzUQwDdJxiXbnzY0Op5rwOs3fBJjO+wqFKEQoXGwnbI68u78CBqGMpAk7ju3gbu
qc9GYa7sr1w4UIXfFk7DwsgaTWSp7UmIAs2wcCAR5V3b5cBiBWMgXh+lyFox7wiOwKNQVV1tBkL5
PGHLRn0ncY0jfu4PQXd+PJn+95Tg2SKtcIiYj030UXvcpkyct4lb3pcq8tFG2S5XQSL47CLogwAu
PAA+NpInQkrUux3QI8ujSgfbnnxIvyIw+j4wql/QyXoRrXU1oUbpeXiVBVrXvV2ifrwhcteixRGL
svOM6kWWIRJJ+VJqyFqRgdQaGsNSu/0Alr2J/FzgFoMdc4OoshnhBgJpC/1y4SukXFkut12E+JKw
suRIspMzKUNCFRRBG8Q29BB2UMfU/sqeijuib4PMEzSoO19q5o+hTTaa+8nxxqluqchVsmrFKTmf
1Erjd7ThUkU8vVrRMgYeC9wOxKkE2/u97fMrXD5uG8AnJrW621YPWqlhwFS4TWuZ9vpb31SjR/To
96OfAGHhdfu4zksXtq4P5Va+lSE5o8MZEFfJewjiKFM018F+vamOn8iHPA2WVPsKpn4fJyxDYrPl
t47b1gb/fv0FLGN5yhjwSBsThnyg079TjM2ANBMTGNx1kERu7nWJ9pw7ECdGWGBFvpsucufTehHa
uRFfE3uqS2IySAfxCJsw4ifImOwpM7FQiWBvU1nq0YPeGCewcqE8tpy0e9BfCN6Rwc1nLkE/jerW
UFwHNKXP3864EWNkpN920uAcBmetOZJ3PemY+G3w3v4JW2EQ+zvgMugNZEB4CiaPkcc1AD6Fq1K/
wUP0nnqARqrVJolfpSjynrVW1CUH0hXMBTtAkTxMto+FihqCiFJnhtgRz2BQd7vH+EX1aw65dQyB
XWp95/vxWMvIMFayFurQH5TcrbyPXnmnd5a4IFwhINEbedgOVInMHAQ99A/xJNiDo88YhPk0E2hM
g7nCZghmBerD9UvZlRvwjSuWoPg1mlIjKqg2/CmX/QFXdb1DyJhVcrY9GN84jRtzckIyl/Os8FNj
T8OAhgLdphS5GMKoTCw0CaIfJksRAVbaA9sphvYclG/b4dPZC435wJARGuoVd1mS7apzi5LEl4EI
rxr4g12akJ84D37wL7jGDBUCZJ5ey9nLCcknu8h2hXsIQzeAxQrpAta+t6Fek4qB1CyatcB26Yv0
J1/nukgxnEG/NcL2UzKG1mUlPMJiuRW1mrqgiRTQay+axsX/Ppe1jlo//E1arSJ+ffvJheT5cEDK
OHzluYHhmMHve0BZrcqWL4w89QJCvks61VYpeN6U/yXCk3nQykWnnnnzWdFpn03Cnkd3RZsFFuNP
4ShpjSRdiKf28Xo057GKd7FIpflcvb0Nrh+0vSayXfNOJ5kgHKu3MgiF/hYcEbs4nIdx7te0vPlT
PAMumxKyH8E97cDB/nwFVvA9mN2nQ0b135HiccqVlgc4C9ZmbkwO7mPd0zXt8tHa/ukDB4MUALfM
7+gXhE/6GBe1YbOYGYrWpzZtWIlp+g+LU0eNrgzvVQTIDTWRJn2V/hANeFd2jbkLCQEe3k+gPedC
wrmMuPxywZ4brck6eZhqv1ybU7CSe2xMC4ay864RZs41MJsDpg82kb4ztkfXjFUhnClg9WUFobMV
G5RPd4Q27DP8DMqcLItMGBlch4rFDgPlsU5+iKvavZGz/uuJijQen4PpgPQRRwGUyxaxsNyQ0nbB
6WtfSl7mCnlwnG5ALx+TCm0nOVAFk1n9LPUfe2MjD+O9IlZvhLasly70nQglD/6R4s2UBLTJ+0b8
BS7CBpIa/wCURmgb52LWAmjutbwM4t1fnZ+lYKYi7qSapZtFSmHxhS848edszIXxb3L/CcD8n8BL
wTFCQVyUR+c+3PC+Vo5SXjYxaZavUSEdcHcj/aXVFgli0K948nK2jjhHr4oz0Egdih1NeHFg94Q6
cGfLuRpyeaIpGq+hVNeazA+tfBs4HbG2DfiaSI4HllCqQWsFq+KbqqeuXey/7uO0eCPhfdGlR4eb
eZTYChyrGZcmtfpjCmIiumMdZ/imyS0wmlBlph9zTpN0wjOz26ve5hl9wA8hNrn2XhJ5RkgOnE30
kgvDbOKGK0bpR4iFBY8w4Zc4zCUZtdGulPv8W++eKcke9lC1lv6D4QxdCG1FkBjtmbF6fmYNqAh6
RuYsS6vKuB0bHwOXzjrgG7Px9B0szVkSxZb1+R2KRnhyDSRigPJ8eK3bq4BnwNZ6S8Wud1AX630Z
esCqg8913ChMpfaAxFym4HUlDtMfv9fsSp00cJ04fzXuFPw6/3WvtTU/R9+TUAv3l64kHHsh85iY
Quhnrl0V6KQs1mOqhv839V/1egFKR8/8CuWnVwSe/tQbWcYbtFLvbxFZAnDQdp9AjGUe4iJkieHm
VBv4gtbjK1UYzWCxdWENjdjMmLzQR+eZXaDRpnFLz5guwyH887TAC7HGD1sgteNS7yElOOdE+bKJ
1G6MowhuiaJvI5qUr/WYW94eKf98CGkj+fKBw5WNuQDdCVhKpakVQSttQ8EpgfDkuYsQZ6kwwmQo
Yl6yhiezZ22McvB1KTL2dw8Z45DtBQlNB2gbUjNVUjEWizgqd3zYlYlQKZmFLdzb4SXgfiy1W/ln
AemlgCmjljivGeHqHa2UuwuJcIf8TkIEEPYMiP9tC1PKUw7Q7ltURTQuJggkWXah0TRxtXWCsLQ/
VbCeFgdWGxbA5v2sdYfz/nZBcm3wecJVDp89/5Y7kqryHgNRf3ICyWNokaeGoGDYGpTxhXosSFZT
cUeCi4KijVeyBMpncsvTP53k5ti66Y4E2qg2xPU4hYabxKtsJ8fruQ8cX7ZSE0S4Z8XB1gtqlQyZ
O0UluQOp1BloME6ZODHuQyYojMi+M44hh04xQVm9QOSzCoquHfttB21TZX2eL6zTrabMjIs0IJ4G
CMmtsvMZxC73vt0FZcId/4lfKbpweMBN8hACfcpPvygGwyiMo+D4XDPNt6N+IwU6kuswCt4R+WUT
mTbhXNr8MD8ufvrYFx6V63AgY+DHxqCtpwupUyeCxzAQmBAsMb0SA9wTzutF9Ie1OonwWEgVHYq6
Sq/0pxswqYuNuKOzJ4OsXx143426SL/336P+2IAkOat3I5uTfSqj4gf0IvkyQrvHU29wLV6vKdhZ
0VpUkxWTPo/jEgkTwxjYudph+9BBKUMDNp64dI+UcFHhlKZpyqINEfTmq/0t9TupYfxv/0Z5Yrv+
FZNuPUJhUyHxZZ/0GazF277JExKGT0ofumUx1IoTqX7eQSJkwVkqIwBu5HBb5h5CoXgy/m/RROU0
qGNZD0S8cATHFmLkhvQsJH1BYY9YD0F0fB1KR5Lk3o3TDMtCeeX2f71LFP9mbuVZ2nq9WtxOQ4/y
3Yh3ngYdtHO7u7OmBAPZZEHKj1tip+vwE9u5T7DXbv0MYKUCLbPnfCV/at3eEbmDctDSN7geAV3a
28mTQiWA/EO86zFQMAYqaPtH+jD+uahigAxbIwFCAgySYPhmxSzk2gzIM4ZR/K2nlYmJMbJgA+Tm
SdbW25OGZcJcUpK+HZBtomcstsgE6gH06oQsaafGZsEkRzAPyd/PCk81eIP/oEz3+EkvPvd5gKCH
EZ3Tah/xuR0XMV81VIlMJGfP87hUpeaKSBO0Ts6Pr3anbhJEcppIfW1T7c98eVQcjST7o0rJ6XTe
s6waSSk2My7QV1KMMuv4D7zOP11SzJQqSpzGT+5DcVdq8RdIO7ll9tdUWBKIvSus4MenFAQzmDiL
V8hpLfrnDV0D8+O9mg1oK8ss0Eg6neHzCic40xNj6ZZN/OMdw0zrBOeR7sXDrHrFRPlRQnjXV44h
eBRhXsIUtyYB7NV578BbLSgpW8onwwH0yM+23429AMG6Om6vEXuzC5HTuwPnfR1u8AhNwJtG5nki
zQeoPgPqtoBrz7giwZxgAdw/bh02VpmaaBzKQ4aowrrLFehvQmleQtGA6zz1OvuzW/bWZ33zPQaH
bfoMeErCCi+wWXhVGruL3vEOIdoP+AT4Q295QEiQl0M8qGNu1UBiHz/PUKnH2CGUxSMi8Az+1GjK
0smbwacS1+AMXBsUyvPcmCACrs8ezvBtKftGb5Je/VbpPz+OMLffo8KW2ki1ajlEId20Sa0bdlxR
uHz/f1S82Km2tiughLfXe669yz5Z6w3+onAX733taDVu6MdMgNVQmolS0cVe9llbdvAAIpYJycpQ
mS0SB2OaE6LXxRqNxC9Ow09z9NVG5roiqGwKPHpdPetHx3GTWgMtjfShPCwIZww8jDD198q0Qy3H
KD+LWdbIUtR/jHzK/W5QYADbpW6UvYBDa3Zr3pjaZUmbAWDNWtUXWqN2qdgHrHYhgC/nCPegXg/l
L7/hnQuFd86P1y/jJqNIrqjZFazwYzzlNYQTiUwOQhZgdGfFkFl9YB7fCjXFJuQREL4j6KPmuavJ
prdvE+yd3htNZ3i7qlDB3UdTtHav0noiOhdYEbJp/dhKrMbO5HabTxo7KQ9Bozz2ARCUhnbM+rWt
WkeHV11/9PDxMWyL6C9spGxs2RXzY8rAVKpITAQWfwg5LRvGmvajMwVxIrNSCfoB5T3/AjbX6Ncp
kln7c9yBnE0rc5hMmcOS/jRVv5Pw4ftQg723y8qMmfSdnGoqZrUwH8jhpwKdV/xz/TWi6VGUgfYx
JqtOREsKwLPk5iXXqbnUPy2Ukv/TDjM9OrUgbm0w2EjL+F7f4W09BJW160I70Tjy5tKPSD+z5hvd
SDdoMLNKWGRneoKwb/PXkPn85qmvsVEogfiP7AinKtzJc85LUNaPG43oTcC1woIY/2YzHV6kPIDt
h2ywGpIo+IEGFIrrFktxuGcUtWvNKgwSp4lSDTl7Kwehmcty5CDHHZzGwxc4uSDLOO+9LM8IP6M5
zBnZiEel9ijq68IHCafS6j3lneP2o/ZkiDIKi8IBTdVHg7jXsP6ZpU4sim9PtXW6D2Wv+hwyr+Dp
HdGJuqzmc6e7nag7Nr2dxnQucvXj/QCdif95OLuUz/o1wgmj8EnMCBKwJQOj/H0/3Ak93wzeauBf
k3rBfEX/jSK8BFcnwGHhtTL/S2GhJlJFmJvS3yoox37fKmDDq+SDvUbaI2535gMCGAiplpQN9wec
FLCRlVxZMAtquCP2Fq2YNYDqhx6IqbtlhC2dEVg098XrE+o+LSGBOTFxq5NH2/DurQ5/FrFYvcJn
73fFDIdeiZRGHrPkozy+IhBMn9GU70jL3JsTLj1dJykQIa3Pk1t+eeqN8X/XZi10aMEQggqpgn18
IA1zA6Cj5kt60/eOreP7SfEv4Wrd6uolrnZtr8QN7Al0tbQqaP1IhBvxfBobYciGyZFVKZZLJdc1
7NWl8eg+zwJ6cSOe6k/ZMZ/cEkx1OU3J1ZqR2QlkIZ3tPo+ZQIvooBOtcIlfGo+D+5zpZzhKFHtw
wOXmSEQrLP44aRtBd2PpEPq42pYHX953mZbMCFSz4NNuW8Jc2ADYyK0ECz2/OnG1X1uRCSWQzbwe
ZdXwfIrw5OORRIabucxtRfO8W9a6KInzGd0ml0HaDOI9FHWwwLteVLhwv42muaMnKouWea+lKsB4
yAZSGNuaiCHGCW+3UFz8Fv2DxXeLe21pNqqHkcjnOcmxN2wMb4ZiKvBwNhC1HESlvzktEFdNY3U/
lefswcS8SZVqYdw8GXIeaGj9bmTBiTq/7VcHSFpnqrSQS8KJGMim0PPHNyRKLiBmzZlRN9sV5D7k
qFpQzrZs9OtrLOIYGdbW4gliv3AlUR+Yld83Dn7MnV5SFKCJsMRiUA1aXivZraNdCmv3P686F4Sy
cUSzUfjjG7X/SieNuXGTLtN4899QxlkCq9s0JKYDF17Y7eZJgxv/tLlJ7LQHoNdwprGZP4Y0lTzO
jcoJTjbOdVb1QQ21UhGis73YDQqNB09P9fAX/KsrivVV9GR/vbfiRx9lo+ptFpTTunOpYIY4mDBg
gi+YkLFdn4h6Z/UGBtc+t40zE1ytwNj91nPuPk8400rAeDQQJCDStOy5DmeEcjga7bvTKy6r44hR
y1k3dzOjiC47+JyGpParGWnVulorE0eCgBBZTCGMrfoIzjCIA2IPj7LG+ncwXg6jI+pEuaXXzW/I
GsNU9xXFad4UOn4r6FvkbX+dJFKZBWpoiSRub27GXqetPmOuxxenwUW/IWLrvnvN+y2+mD9HW87q
ISe2VfF3daNWJ8Hl7tqvRDBwtfhkSbogbK7LtUTZouNsazfs8HbUg4QfFseK/5ylZF0EdXnwySKA
8661QxPuwnFDQUpZkBhyfIToHhOlcn4Cyx7pAG7T0lcqnMuNnTVWndxr/xCKOeXZlUir1v5YQfLw
/+mhayfvYQUTEJciyA7wSDQwR9fXfoiMlBSBsWD30amlVnlWWGpSVQb7ASPSr0JgCYHW4qBJW+ph
zlPh1Gw0iuSdbcuzc7Ds8m7/6HdZVJcTGkpyqN1xfOCyXaNvlWpe9DFKCyAKUhuxTv+SiXalXF6a
npL4zQuZPz9/Gy1661owMWCxo157Bi4G/kxLvmXIcuF9AlUW1LkpNmKylLQ2c6i1X0Ds7hlG+uTg
VvAZRNt0bFzuKE3fPzv0DwTBwvaNlcDWnV9DbzS9/SdlYA8k9dv2GdAx0pgdnvuthVghLyni5wQE
C8zn0biqMzFykX79EvFkuLVY6T9e8PS7Si/Ha0g+gqu24rdHABbEzOv96gCA3GLOq0NrhoNSzWiu
bp/QKQbKmqV4iENxCVGTsvOHDbe51Ebas4LIUmoC4j8/AvLvXRMgGBarsDMXsCxJbAq5R+0Spgb8
d+5voURh+XCOvlQKBhyNTuHo2nipihT5+mVTySnQuBcZhrLGsp+p2qfOoKRXUwAVFPDN1SjRZRge
T7BZY094m5GpRwHta4iLUj5wbWciJUrbbQ18R6uJ4Q1NBjp1Pv4IHaScf7/Kz8auuQ4N1G5AnZ05
81AJ4VlFFLtZqkbIJhV+3NCl89EzX1nawwVKcG8GfqDnboJMFTydlj9jjMvlCGy+X7yHogiI+T8Y
clt8liPCLxbOscQAfhtvZuQps9fYv0Y7t3YievKRo37itufnF5L4zg0sO/dTZroxtBX7a9nohMCV
7ywbs5NTF28+iz5TKaSQKe7l4AHeuOPycEdfm1VZU+vBtlERygSz3WwxMhE1ubMABPC985n4kqWs
065+YAnW+vJkQYdywEnC+PvQRwDUsG9Cu0R/9brCiANN2dq3yRozDOwZ5OGd6l4tCDZvX2KEoEve
V448yVNxNovKsQJ/+g2lZmT9ay1TwcqBgqIDoa0bP0mlvRmUzZ7E2pp8+/AEpsqJ37rWJWQ1SnSF
xHGL78K3sYJcUDCzLFKXfnAMRAzb15RNM0GFfdhpa/g87Q0t0bLMmbLAGg/cqMcPQDotBp0XVTjT
mXe6Xu7KiaJGNDCZkmnaGMfgpvx9apCqbg8g0uWytQghgi+JvDUJ1NqavzsZgYP75wjFplvZXAcm
BThaVQ4hppk8I0P/km2UGBEJkrkxIH/BGbN/TPYc3cJ4sf4796aaHTaS7hEvzQOlGM5CsLkb3zPF
KjlbTnHQEQ4xIHAHVWuYF1XYPhA19cPG7sizEJE1CQeAZ03YVLozG5ngCt0LIqqlkmdBjYlmFWeW
RlQ9Mh/kX7WXPS3KsGioHHAKdwHvSexNsItKCgCoflD2KPyNhX44Ue7a40z1Vi+2I5eTZMrJxAmP
9aF+8ka3Sn0hj61azxD7QhTol9Q9E0H70DZcgcGzuoXWtY4iCh8m/15sMx5XazRh7T8u252/V5uw
LQ5lCcF44D0g4eaY1njv3cTDEhsqaXP3wV7TqFVsW9Fo15zx16h7RtXsmrXIlGe7SDPw+pTAdsF0
j5t+WMRj3GGDaiiTZtIbcegav5ZgG3qRysXg1eDV223WOw0Cqy9y9ItFw+xWZuJHKffas+u5QKl7
MeC4R5AkWbHcVQXXfM+iEfqHR2oOlTxtaJiUKacNf0iWx72iyStlunSuk569/pEU+MRfGQMA6o2f
YAd4mWR2fKmF+YYT0palI5Wngxl7Pt67AbxBWmfzJ7AnDPU+Y5WbuyQ2FxJQv/8LjIZj2OscdQxh
pYDNEbiYceAfcyA7wcyoDUdlQjuqAss4k4W0i/Qfrfy3iE0ED9RNVCsksMtGHx/EIQFDJIJM/NeG
K5Mxu4J5ABO0c/NtM57cIxZxy4Rl0WbNysgGrwimpNf8SaULeiKUYD2W4hvUEgy8UewMzZoF32V/
2nagpS8/4JOcsrOKqgrtwnuvquhu4KmZR6G/RDexjBEbF1UoZScfhkSqBjYSkVfvPLJUhSYOuWFf
OtbzpNEVfFnaeE1MecYDKamT3Kq4hhWeXe1wU83jC95vc6VAzRLRU/+Q1acLXHPT3Q9sbpYX+R8Z
tFI+tUxfX7uzcuguLUTmAY4G0dvsPJ3V+fnLEMBr56uWL5/XEnyPusXGhncUAJWLhq2otdIOwWa+
L9cxHf7xgTu/fsKroMufa/Et9TB22y7JYraT/BKAk/+6fWOerBVSm9p0svxMgEdvFyjSRa0hZn39
rubFhRuJh2kWPetrhJBl1q2VkrzWR1Xj5o2gsgsBIvIow6wNuBicHS4xl2vC6dbhC3e+WZgDvFq1
WCn+3bcJ9hNJQWrcDFg3GyS56JBDuPnVJeen+GiKwiTfNZ0Aonaza3WqZEgYYRSZavmHygskS3bW
XMGHAT4KDf8MvjOFMKh/gJ9GrR5D6YX7IrDNYGrjVHLZxQUGHg6+YT8a0ApWMe9XGpTEISuQ8NbR
k80SzPWYPzaPUFwpb8AkpJcp94FIWhTGh7hywfaV4NBCh327yiofTdbPrkSMawy+DI6M+0OB6VVQ
FFgm+8doGYiyvBeMXtqiqoQhsZT8+aRA/nb0Cov02Fis0+ZTOeJozTTv2PM/5pHdajgCx5Ycnugh
0l659KABYenc3L1uHDQvGd1AC9Pe7sZOOSC50x7GWNEuk/e+1aT40ogxWFPkSLDRx+MmZbcoRotX
+OdQIKW1bmosDceksjn8CskfImLH0tEkkIdCvVg1m/jGV46fO+XO7buLbWM1weveEalXxqlB6W11
ofJc007TYXCMLDaLqPwBluzrmQNo8mr3cjELlR+xxR/n6RYfxWX/2mNwI+Slul4qZlOsugchK7Kv
WedTwyVHJ3ONC4E/P+obu85C9qyOSWdm+PlXGJ9+9BqgkvLyIpfPCpME5eGQXNQ1ZUQr9YN7KxrX
5ZeAV5gBvwdp9jc7UqGalOi04lea1JXP+GC+OnlL3e/lGDbLRv8AYi9unzH+EcWnfOh3udu+izE3
RvbL7LY5wGYYSjvLatMg+8lcGGyIotKTteTVkXfMORux5WYPUV3ryNvqob/V2mkwE7dXB9n3NEkO
augincstQ4ob3RHkGLkRObJWi6IUwjZG2GkgSLHNUZekNYHk5tD73sRgJSKBSLSWs8/RSdqDQufH
Vw3eoZ9XSgg8KKZOm0xh1p1MJOIZkA9Uo+ztCFUnsLp1IGpiD5oO7ldtMfxxUuWgnx5RNvYx/waA
up6RCFMIPITXaVMa5xpflt6jp7oQMXjos7gB84Y46KHdQZaYTrnTn9EACvsF0S/MAFheiVLVkmGB
IwCDxoDpb1FyczetdjUUVcy3e9MJs/a0S4LujcvOyAVg7wTj6MBLD2FFPcNuQviDcUbhHdnYFZpx
7lxbEjodF/WCVi2ZN8+s9tgI1eKvWLOsL7CcCUJSWDGdUdKgdqH1CGEWnUf8paPVRSi0oltnc8B/
QkUAMAytdVrJo9n6n2EZvBIrJ49AiNz87MfT60gtT7iFHGu5gUcLPBrMLrBHY3LBMc53H+FX+Ta2
UxeH0hT3KguJF8UwTAlboRiwqqFbNel4b3jFI2FTJieIXHzPRmyZabzvjDXCN8yjoOW3X6zBcY1C
VifNvnIEa0bfN0ZWVfZpFWRxYm7D8iYe8FBMkdYa0sJ4mJ3p35JlwwymCJ8TiStGiVgrrtdnT2Lz
R6y79HfP54zJd+Z0QFMPtxsOkXZeHOwzw9VKhTGJ84Er3i46866+liZFqgJbR4HUnyErm+tx/HWu
BPF34TIkfHRjUuXA1YNokvEPSpbZFQ6ybOP+QCTXv/zI3Nji9uSe3TitlCHwdNugFR2edqMNKGMC
jvAI9J9gUe+x+wIXNMcVtvYsKLfjFuV0TdUBt55ydgTV3Jpe9Tj4Tmz2e9O8f6R12mGXTGCN9l2a
lvsouCY0mAPkJ4RjCS1VcNiIN2+6YOKvAMiLDjIvEm1FcrVUp6TuG28A3z/MV4lgQM47TF8qU9lk
9IxqS2oFBBFll8qi5RFTGNgic+CEpsV2GqrqDAsieXdqGMIwZIK/UHTqDrvGfC+gvDEaceu+s7Wc
56xvNk54FBo9RKPtWrTiOufD2ZLkgwfdvWj7XQMyUOi5Z8SBq+0q/IwoZl5SxScTHJmGPVz8izM+
rPngTAq0s65wOAuwMoVHXXTm0qBBw3AQ2tHnN2FKc+llfkvnZi16W3MgHrUcqee5G9xqHdeqyk91
9mV+m1fbDUmtRX7Y0zL4mLnw8QArnC3/o+090geeYVDSgHHKbtxexDNP4aUVdHtR+bod1m/870OJ
2Bc/Oasofgm8pL4dIlshzQE9NZX/JD1YGMgpgW2yxsKcMuPm9hIVxByt+w3yGqoQXjbB2aTE7aGV
0vpoO6n8uUPvxN/Lda96yLTVRuyLDsBNgE+L3dp8NLzzqE0Pa9id5tNSSV9kVNpy2/aKBC7Kfu1u
J9V0cRFiypBCrpc0SMSLeDiU8K2FB83Kf4juDolcAHwSz8g8OlQ8d42zBWqrTTr4ffKvjhvDYZmr
vlohb6Fc23wK0VwV5p5fpSM3gfNLaM6rseaX6+1m2HkKDNiQKuC4DvU+sfALl2hseM2wNEtMLb0e
4AOIh7GGx9lF+T4pFZ4TWlGt/3wYOTDwxniDCkkJdbbAVdO1VdwJDbR9TnbNGOzi33QeDMOL+XHd
T4TUBVYey3wbsLG6SGNpd5LGcWRsgZox52HxVUd5JVgM16SzXJ/63CPZHtqlZCoUH67spZhdTYYA
d75qTHEh/bJazuBmfnoqFDktcJjlaCzLNcdUrNoHIRD7MwwgY6PWhye3iNPxeYeyOOufqgY91EQl
sA90gkQ8LnkuhuvqXiiOJ/BysVu0D7AtD8tkO02t1rKR08SFYIozw3U0VTjwcckSb5eCSawLvyYG
/lsqCFvr/eNVeKIXrMuPBd0H9rnrGa8Nxa7eL5wn2KyiZOKsaQ7rR9sCzKZ1Nf5YepMt2J4gPmVW
a7nNCSb6Sj4urmtaVBD/dwqe7wFd9iyWFMdhWBd+PeQmu+pu0wRkn2UegedhqE+lCy1q9W+wDKG6
bbM6J5Cz5MXBrcdWgRdpDq5301CzGn4m9FNXRIWX9EK+alTmlfNN5Iuk0kzYMZ8SEhmbLdyWQBUI
ikJxr45kCMMHAhsxDcy7gsEzi7ed+hHpR9XYiBxmUwzNqPR916fxkuXVb2mqcrW1ylYXvEZt65ED
CNQXkESLb2SkXWgRZN0Creq4ANC7FRnXWoX+J8qelH3SERLBVA8xQ/Z4wg1VC12UdeRCGCTmQVbN
ioFZ4DHijkUu6Czxlba0DRwrFlcOgabLYj++rSfZx4equFh3yLGQqgEKzOIlGxCx84ZTKktbCWcP
E20eZu8FbhqFaUDTUc1sZHbGzPL6cxBJHnlWiVdPwTDKnkDggZzv3QRrE9gQqxKZ9VFAbyfQJ1Us
/hIQUqLtuc/xWddq8Di/yT9xtuREceM66WEx/ISCg5kgrWAB8Eq2WTPhLhBmwFYCYpyi2po603H6
gb5hnpjKz18wtoHDeWs00X9VYC4DZ/stzSeuCEzLEN6OZP79G5QLzUZXu98rtRo0stR2WNI1mm8A
IUmVLIrqh3+1NYaJ/gqGIdslItEwPxuMZ0waWaIKBGdgEO+N+PBHHLizwXwYPLrG9uSx7foDF5o9
N5+hlqwf5XGGiDEaB9HLYrgpXmKF5GvRCt0osVU0TtZp18Tijv4tJlp3v1uI5iM6jp4etPfPSvyj
69pRQOQwmqktzRJq+9KGcU3R6+Flb0R20doOfR+1ATW6huLWnQUfexGKED/Dd0AkBkwYMsBOYIWr
sEtEEZlz2Ft6ofRiuCWjgPgtGib9TPEP/yW8Zs7I4KnNy6ZYDsYQPugEiLdr8R/8VUvm9PRg7y/z
4v58kfZ2sMZohcwmBY+Ou2FBz0Mv4fO9fTU4HwLnzDzuM8eqdI7EH4Id1Wfp8PzZ96UNRPIaXu50
fban8ilFHKtfYZ/0ARteR7dWgq8f6lv3ycKGp1rdtrMPfSMjyHwNY32PviPsSKcp39ouWAdWhLE4
CAqOXRufXz1hfx2QqigS200w/bA1AJtYdfDfAEDlNsDXo4QDksCHrUiEXSjlg4oNt9GSAr+/W4Y0
shG0YL4p4o5hZausXXyXsTO0qb58FtsT7ScGLfNL+ifYEMvIsBv37YLj/5po5TySVYG6rx/jcJI3
D4Uzy+vs4cKvGz6MGC59JEVbbB0EW6wA+toAOKXVRMPwAjgYEGt3qixQat94Nw5Tka1jQSgmNBrl
j7maBzSdFpN0oNh19HsWjIXJ1FWsANOnHetDnefLBBh4EFB7RzZp0QtNj7FCDEFTgWaeet8pRcvq
eUuwsu79wSGj0fw7mtU3lLonmSa/iSIBy5R52oKXdQdwXWCFL54RfGpdT+FhXBWJlqUA9oh+xrQ9
PWSt+LQN+upoKbr9fyP5TgQTNKmmi+1gL41ZOSknwnojVn6ts65mai2gtWcxTcb3YncJFRqJHuUI
afNl+GAKnph6k3xLzcBKER4pRZ0/w1Qv7kGCOt3X/EScrTXns4rtWVKvBdyAnAC6138JV6n597SJ
jSwx44wPnsTOlpshrOikIRiEWgnZQnJpHTYf90S2Uwi6ZVX2psW3s6Xu1ahE5Vu/iaMp/0/z9KUi
zQ/XP3Q4Pm7tj8afzvlx36SY788mrcYelE8xpgp2CF+eCfwz6pnkktEStrKhFdvmreVwWvY52PF6
93WEpIMB+LGAICfhrUZlixCudDjeWk6+W6wcZjZaH6cHStHSlBGavncTiGGNRcELrPhScdxeiLhQ
DFIfRl3NsDHGUNLsKxTTnxx1gmAml2642xUEFlEy4nkBhjwtfvy9jq5VSahIvnQT3EegLDgSHeLW
HurbXVU0Sp6sNAy3YK2TmoyuqiqrfrB8Tz2mfZyTrG+8QrjP5Uexb8UIVk9Lyn7cLhf0amIVLrM8
0AE7Mn2e1GuOuJAVmyFiFacZuqhmTyJWNS1cnV2XyCYvpJPVwOqrlou+p0FO0J1xkLhU/rssKmX5
FOeS4Ge4p+KtvDF3C7xus1x5GTrPJ+lvEKyCAGOJJlNHK3XPzOPgkxpOTVZaQug9KMgDTnYkUiVH
YmBR1ktHmRl+exPeTQCUD6whWCBucHdCkLjRbdpGCQ2X93iFbqaD/OHHD/zxKS77C/RW/4fOLEj3
ZfajW7gQkg5BUhJWtnMi+oHcQbm9rzsjLAPj5tWc/i3jJOwrMKNzppjn3JbqWnvzICHyQMhlmrIb
Eb66RttpNXetWRaeEDoH1zv3FXSsva7vIALckTUs7kFGAu7ipinqq8eaOtwk8BuXHa4zXwl47pxw
kIQrB853TZ72IpvzvNgXJa+NLpNilyJXgGrJmkeQOOtw2g3LTsCNBZc2TaoYJV4CH1B4QX1VWrKD
5QxHQqUle1sLv5G1ngFoC4JRRZBjVmJE8r+NukxiJ2z1ACOIxA7WcJiovlPdiMrjAZnLZ3VzMGtG
bCBSI+OaaEFsD29jVaFX2SNx8GCjoYyHz4q+heb2RvcjvuXpNxYBsY50sEpfvYZXj80UG8zGnF36
jCbSqqeJTWQCcnB6ne4it5gvM78Q6iLT15gKKoe/+wxLA9cTnLjbknVz/Z2yv/S2qKUaNVT3jNSW
WknwAs0kLFtA3Kq/d0S3Sg7a3yLPYvO7NzCsvsX+t0nKYc0enRXcLp3Ug6g+gI6PrzdtVP6BZ0aI
GstG81nwMILqKzwe999MPRDe3RGD3XfExqlxCdX4FK32DAQZOGvtiy+Kollmkjl+lXZzr5l07B7T
9qlsWbkjq18ZV/JefFkLj+2LtN0W7OYyhH3WLdpZCqLShoaZPePihBE1DwHhUw5CAjc/Np/vZElz
KxyZMZmkYFs+5Jvh2ru+InD3Gdc46Mdd0zZ17UCwdnOxZ0ZwRNOXUXf+2i5wiaRdbLhgrPdjNYsL
kz0s62b3j01ca/t+vK2adOFw3RXdn9KRlFcRZFGevkthl2U0tcp35AuWd6NApOxE6fsGODF/k/rQ
pNZIf95+JayL/aJeGGetcJvyeTHBZG+RlVnB93QBIPp74hg1+k+5H2sMu+orvozjZKOCpATXA1HJ
jb7MZw6qm56gNA5QTW6PndXHS6cx5uq0D4/u59lhnGd3lWmg2wOnoSANr3aH0YuB6v72H0pxRWGr
SJYOYuCr+wYx3fTcaPYr7N6P8Gk5MmkUe3oK9AvN9TlJrNIJPxkqgX74rlDbkdBj/7N9/UIQB6AF
/hghtKZ94mLVTpDhffVLXLTjLb/54VXWTnHjjJvKJjuEy9fhqieJMERJxHH8dbLhPleZ1pPEgwKb
KjELrxaWEkQDi5zzwmjAPRtNAKJvFeJoFDLpfto5R27pIE1z8CMwD4I8mDdhhPppZsd78wPjjPjW
s9K6FTSlmDMdAZxyGJJx3HW6O7LFWBGB50cNtn5NWH8eB9PIfSMpCMrSuE84FQkUIhy8h4oQGgC7
7N9s1O9LDURHYrXRhxFgsE9SfewYWB5oyLbP/+1JY484OpGxcX+xiQ75kt62u0J7bsUzOnkYQ2eV
F2TvJ3D6uTJQpFqCbylKMrHmP7LP4nMFgbDxJ3BaYku28dabhdO6GTC/hmaTwuvDsmYlDOZ88D+p
8AaZkzpAu7mxZxItShrsbaJ/2XvNYmxkynHWYGh6WvDPOresrUeR2JrLkzjpOZtNVA888yzXJvwN
34Bh7+Hgt+5eVyNNnnTLXiJTJnf82eWuQDZx0jDY3N+ystCEYChEhGR4bjxvqR2S/P31uoZlXrxe
y8uq+GC2KPi/QnOvGzChbnJKywwnpOOwGGfzk1DyYX+cBUVSRocTzxdlCDVTw9W5G0+WSp7WDBXx
xjggmVS3Za4G7o5LKXo0GlaZUZUsgovvu4hwprnsm1EW9dNRJH8OJh7/5OGWeNdHWoV8AwdTjsxf
7ET/JoaZwQ9Unn/FusFETGWlrFO7ReNfUxUuYq6is5LPCPKCnkw4tqx2LTwnwEWbCqbAIuDPK6Vu
xsv9yHAmoDjgk5AVgpl4dI1F8/Tw2hcFMyOgV8Nhhj7tv+PH2HXGczH3p+dm71es2VTs5DsZCr30
OG8PmVOeGsn3lEKizOMqcsAC57URlMR1oPixGHncB5ygD2eHJfD/o+8Zj1L9GiD09PsGV3CsS5Xi
yvuZFPbbLffhTViB2yJANEzyYuGO4TRviQchd4VVefzl4Okq2udXWmeLjthqUV6oDEACqUifkUpF
jK/NO9s0ZSUC+Ju5Q3Yma+4Yne1h7worU+4Q6/5qbRR/fNtUBliyrreF8ZoqRRa0sHatQJClTbZy
eo+f1kSfkl3Z7bddG9Wcpt//Jul9df5bsLf3EV8i1NIOVEcX2Ex30GtkVek0mT11AjG5TqRxq6FP
6gdcQNm6YFUhzRjyIYmvORKMGEOGYzlpNBk9fgTlXJkOavnjfHdq7aXNWuEp+qcd6KaJ0PoIWI0e
gfMVS8vYvsE3kIO1fcBIEdNqAjN0XjWv5B0t4ROBHrpk9Jo17QIi4/jX7XgyxggM0Qlh+M/Ca240
olXUHX7ndNnMVzeNUlhQZsJFBAIGqn4iJbwxci6SR8SZIhfPhSiiKUJ2qZGF1vfUevmqql8sSCxR
AzJS7M5eF0YISOpnsbBlFe9t1M97eeuZ0KVeHZVi50cKM3m7x2HryYWJ5NznJkfzSTgG0dXmI7uX
fP951IJsS+QQ80Zad4sBS5wiSoXoqvmyxA6sx18pHDJQnCYFdV6T7/pDJxGj2P5p+Ljv+3tM9oTg
jG+l28uNXso4Zl/nLgM7NXbknli5lD2pFDWvMS5Sxrdn1B3h/2ZnSEpAAltWz8lJ1uUsf8UFwlxE
nyE+GNHAx7wFDWq9z/mus7wlay6aayZwEk/MfiaUfobLPKEXOBdenr3ECgcBiKkX426FQKLHlleo
rgjiCtcy2FOXJdWGvtnhhITg5AdJ9SaLryKP6uFKPcmpWTxQC22ZsjaC4lCNddZqDCZ8ePbzlct9
0dBCLy8b1kyczjjwkCv1wRGJHLPXyioRwMo2xMBZkCUlum8m2GmaDm4+tUbcf3W5+ARvIkOR3rBQ
8z0mrU92fAJ5UqoHqzfbU2pPkfbAT0XZrGvCbWe+wk/du945MMouZhFJ+KzcXIMGajgajzKzZgFG
0mxIo9UR/2g1Em3UGYBKqtpSKIf0YPUwjbkYs/RXW9Pg1S47HdYPF/uKpm0BgjLmERi3DefUt1Yq
GtAzlGzVaBPAedKg+XdidKgMfPlOB/V4fAMXTTzBxUQOvqNfUeAsYJObOwyfafmqekugmtoV+OnM
zgdPWgn7f4KViE4rUUXw+RBGIhSmGEk9kYAt1aMNBrA4OOdkjhfy9BCitYd/hNTEp5PwNdAwk4Ys
ss+dfVKfI7DWph7mb4qLhKMFFuceyx9CKemnAI35oPtAzfJtdRYa0yYB3BdvcLXzZMhlQbvWvK+l
xmJ1MX+TYbAqyN7SvznqGnHViBGoNOX2ve9Z/wAcl0kVEUzBwN/9OMF04PXIbypcCNRotHJTA63j
rWnYVjJFFFp1eExFzKpoN0iR9dmJRzfkyTi4h4dnhI9xVwzUNxqSf2VRMPc2PPYF5gib/YJCLLip
BrApNm7aBaJ1nAmESTUSfERt89kBVz2FVueNtggAzDLk0QEOk0hqBcD06BH52bZ2n4B3vqOXLDRs
E7b62xdmpWL4rcGbQGY/dPJc24HZaAN7otDPD+XzpoVWDSQ+WnxWwcutUowaAftWhZtKMeH4dk1H
gTbmsY4t0WkxF4OQxiKgi1r/rpMGn0Hjou3Zou3YWBwEtWMDctWal/9Fa1qgKKUM42F6MSB6Hk2u
wpfw65XB0+3SBlfODYTWBGmJO7PaszpIgsd2w+9bWVd3c5lWN9nKWSmhMowL/xr2FRD2IZsK4+Zq
lDKtBqWqisAFFfF3Ay9cpMWZcy+LbfO3XK+RgOBH61cCH9f13lRbJE/rjXZp7dGDjwgQzplCTC6M
J0devp3RsJmdpKr/UbuIfqFoRYt+ZrIrxg+XnES8XuB2zW/V9EqEZEBNuejh0/G5YL8BFyatQZby
wGo/YodJ0DXimfCEE9ldyqtKQ/5qUmTug6SzVBEd3YIGPsu4Kkcz2+oZxto4Nz9XktpnMYifRR37
quarjWtLveHZfi6/2aYGujUXE2IL4CxhDlTM01bkSndanXhwtr68kuI6Y9Szbj0uNHbJtlAQglD8
3unPHVh7stSQv/Ip861/AN5ZLzAThrTAL5Dw4MmoTG4uq2viOHz9mt6/CUPQmyYkcZkSlKfYCQRe
HEE2turtUTpPgsJAeTGyCcD37MMZjUBzwaW86Vbot4yHKzH2q5Yxk0tZjOvnLP1lbXxLmsVcfWh1
foGwLt7/R2Y0GCKtEEpdoTR6aObtX7z0RBIkAGROoPBCm7dscTLfv+PMxTsBzFKHWB2FKw9lavmr
sTfBruXgmtHlZ2/TtOpNCpETct/RM3THYRU2PE6PV54Iv2ADNWstwylfo5sA2skrpT72h0HkKU73
a33/0S0i+iCqD5AkpyhNSyu1sHPkW8jopVfOtf5D1aBajW/wTvU/3hEEPNFQxduNPfIJiG3r7HFi
287nWEs/ggw82czU9l2dRtpq1XpSGUJuZvLUl1VkRMU2mAEAV9udwdc1sCgp/uY4jRSpFxZYNETH
CE3b2XexQOBbDfDOQ4Lk3sA+KXmp2iGtYPEoZgolUQyUfM+0BO8NL1xl0sTrd9jQMccVY6bvM5FF
s2gZMaymINK902tw5zjliCGA0h3VHHv+ZKja/jqDSHO8F7kRW5me+bksm0iXUwnoldyOdGgw0Fiy
LQDFxi95YMVTgSTbENqv8ZnHeU3E7BO9pktZT2N/AZHfZGfgedLaVW31YbvgcT2Ec8MrFGcHGoTj
9ISSn1PrDjYmUB0FSX/YXPo88tvfxN56ezi8pEev6Z/9oLcyur9+tF4fk5n4JT4GLG+0zZuCUWX1
IL2Sa8TU7NInwos+E1ikaXZhWMeZ0C4S9LKJqwBmytXUuhlb1E0c0SqtDmcmv8HJZrFdaILUXDHf
NC2jP+WPWLHdpPRD/TncAvaJD5Zuj0Maa+UZrAJLRh0CcSG6cBd7MZ34rdz/x8GAFvUKyqzMwB/9
nGW9FSECj7wbApQn0GsA7EwsKAuCGBl+Z8SZIowqBSzlHzKLfqKkIqZPhbkQ1IUxHttL0RHx6nAH
uJuLZYV6Y8xJQDHhTsIkeCpVLqtfZj1HQFYGwTELUyXGDQ2EpG7511MGqKkXNO/w5+NQ5cvGYx1z
LVEed1Yv43kqq9mostVQjUuMqgi9jQrqngvBc0G02B9bfQQMJTImVo5zLnwK0+dQuxO4m2EtN5Aa
uDys4DVIgd0Nvui/zmy8nl7p/YC6YJe7lDFsoW7jU8Y8TbHMbQ1z+CpyhY62rEiT82pE2YpIUtEX
DP+7Rzoi7Fj4iZYKQZWH1rfRIsB6HEF1B/jcPGiO53D0O8cU5eMPNjLDmYYmEHesbHQSoaWoTihs
HFGWXkUQffr5yn5nZ2f+BivtXYrY8tkG1LFkmuDoF0LCbCMx0UkJdJS+L7hemvreSrpLsm6MjjGb
juq+0UdirAXTTMZYyBN/VKbMbmauX6jiqc2UDd3NSreJEnZRWhVhlsVOizRUHVWX7Vdb9SWQvcW2
KPNihKamT5gp9f3PcdlEssR1vIhC530Bu5KLeNs5KoPY3uruMi5Zu7f/Kxu/fntdEUsVvsL3jp3n
eJUgMyjFENWca+BighuAGihEIummJ8QvnYnegDyQdQyCVH9E76FL8O2OmtoykiSpYFOm2d9+MasG
ssqe6AlTxOSPgj5GoxeH6alrKEvfQYkIxLK1Ak6UadOocUKw11KrUE8Ek0nWsLhnmjZ5N2hfL/X8
KEdCceNcG8btA5Q51cjPstKd/QVOG5NGRFqYez3v8b5QrYu3PptAtYbIuEwC9AXWn8PsiY5U9Kmj
sGNqIgEet/I8fhC7LX/hiVw2De2NURa72fIBU4WJIOemphFV/LIfAZCZIWeJUlIsd0yrurCn3TOX
nhBorVQ/Ze3vOrciUIVKHKipIqtzvKx8nICNP9TCAefSo0g688BFtWbuE3BMD4gP/qHOVWskcnhT
ckWn1z54NmhbR4dtD86yA+0v8rKYBLz4XANyfpj/I9Oz9Y+umvkRDAMSpJkuZ53hStDsFidmbu3D
hUxfnu6mJDY9YvF9JPXr5iiAC47cZZc6sfavMloaNfGPikHgfvIX9WOOIY954mHE0CH1SS8jzcnI
Nnt1PEbqYOeQvtrIAhLzBA3cLKnNgAngM1QlPmbk1nCGtmt+2zKCNfj2DkE1RiUccPHwL1Js5t+Q
/mnXgVM3JUaDdqIzbuXYdVyuWI7SZPUf4cywKR47QSIsfkuGgbFThavjXTTphAnxj0/QXRM45xab
PKshLDoVeq6dSfEO74K8eFoUKN2uwOgmndg7aYJ/ZilfqPglr6R3BjEFmgw9ZmjsIWmBNfTrhexR
OBxzzgRzklZ+/LyenrxvD7ZKz+N8V2BD2dRf+Ufe9ViY/C4Iv3b8KiGoIvBhCXe69baeic47AwMs
RaahYy2ruKgZLd/IUh8s8pFUioLYqOkevW8t0MxlqnMZpaqjOGVFKEmSqfFEYdfjuWp0v9RkUgyD
70MAAaR+v0pub7vVqwEUSAjUnbls+K29VJOX8cMIiW5rArazs7qUAtStVWnwOlcbQPgpIZ5LF+3o
vgTbYyYB2jPPl/kT/3SvIUxmnQX+BMMvIu0jqWARoEBLkmJtVUiN13CnO+3juxc+xhQ/dbQAGRql
1ZVinuvmDJUglGS3OnBbso8axBIEsBvh+2xabBxujKulN3IKEJkOWJOdKrTtYvW+NPFjHpiCfS69
e08vol+a9mUmO1G56pDrYC5NY/VfBX/QFx0VXvPHH7f7Nuw7DcAoElbJfSeZpCQI4rK7trfMKY/6
MrJEu/wJ8PbzumOOyDpQKxoxp5iRYVQJlNFoAsV1SRXY/Hyi3ZFQ/wHy9ZamL01znMqoFRws/2TK
PUmbLuWcA+fZmJsXtldvr8LwSxGBCRpMBcVEnk0wdN7FUdbR06OBnWvdwbKAmXGDMGgacNsh5jEz
geYeOXtTUCCg1gS+16VD/GXX9o0dk1W7evvDS/Qp7am0UhpzCJhqDvroB6nFqTmi/7Wi8LeMpEa7
bLFswKs/E1dyQj6n86iv7QYmKEddGm9EmZxxNFfRCUwEyDpC0KSbF+5wNWZX1+8VScco6rK/T79x
pomnR75Eg7x6CK/kQMJtD4yDd5e7JdzG8HjVIsG2iSnklcnAlnU4ey3zvlcBeo90RtwL29Yqq/5Z
PyMDQ+iSEu6ZdzLs/dmSlMwVB/ZRbStqBcCAlpKZeHCXLX2bREBI6qg4NdoXeEGd4UfTFnK/wAGf
xl/CPlAJYgUvAiCLWPA/Rz3GAkl+A2QOmgw6OadzuPvK4ijsoQeRt4TDQBuiHrXHP7RyP1jieFSm
ftSvzdVScN97w5einIpfVbn6tWQps2AiNkKNV4U+t2Yyt15ze2ZOdrcIPdDrsEh4jTig+7Oec/Dh
ocTkfFwkYJkeIrSnfgt2bOXnM7/Z5Bz1Qq/kIokV0XbPhsqyPKnPb2acIWoteRUzcG6E+KcLjvZN
tkuYXEecYv8jrtp5h4pKNaiCa69t6XWoJhAiqQgrchYgVQ3UFzENGom65bBZ858A40/aqf+fhOBs
M0D6dETHRSq92Zwluuhf9b8WEMBTG7wW4M/zjr0YSPXvPk1H6L3IRfeN3FhLbAMTKmHBUbQTPq28
LCnrFCT9er+lXWRdBkEfrm1CbENOpZfIpBDYzjgO4TA1JTyiur1bMwaclpmEY6+lX5SoqxceQtkM
T/8G3+cALUeNMU8zf1zWMQbcFS/TCNZyMcrJCFodw6IAhwOR3OsQlfsZRWAHVZDznH/lz5C8m7d4
51OfOcQ1P8J2ceofnbdLoJbX+Bf/+pnh9p8E74t4GGH3zXPp8VuBmCE6IgVFhxokgReFgq/3ydC/
MAHEMQwqqUyMnu45xM9rRiNHWHKU6sM0qvQuc8Bcpu9pbmFQ6ZwIs5Xs6lq9kpci0PIsL8UDnfMe
azwtutyOiJ8CMKrNlrRyOzd9e+knrAWreW/svkGvPj5LyHU4YXWViWh5++UE5NGzOAre756ktRZz
D4Qs4AyBJeYP9mza1DXphuZ1ooXKAdCRpFnj1zFg0jC/adn8ReCWNV5JTMaI5Y3W+/SbTUoVJFb7
Xek4LfI/niGaeJLy008IT8pivxEv3eKsdmrqaCD18RhnlIDLBpgzKPjfPrTs1Bcc0fYWlLiMAK43
epECOlqPHa8rd3JIzLdwcWwBMQK5rC5Ejuc55UTrdZVSVPfKwKjcjq7CIjBRzRzczRQXdGOqYETA
LLOd1U24fJThFfI5ZtyKM0RbkKm3nK4s116WwlY8uil2zDu9aILjirS2UBG0QSToCqNgeKcObKGU
rwrL9UQDA4xVZ7RoVBDKZ0eQSfry1hSqXSSNeU1SZmfflgOtKX/f307Clc2v2jlyz7sV/+GmmhEX
ymucg8lqamgfnBPrYCmf1fHeP/5U0LBTOcKYclqCxzJzJPUxdKvi9Upi9Cb54t0tdkaF7P/ibrY0
agz6T9iULT2honov53ekxQdKXGy18JZFqy7KnB6FhI9Mcp1CbbUQgYqPMqtvjBzIGvBWpuNsRXAt
cRcH0IZMBI81AVzuIpPT5AQl2K3PO4j1BzBsn3UFy35Nv4b4rJS/ENsB6MXkOU2xwiuvm/cfDWww
W71MjqzPx+G3hFv+aVESfiX9l/Qm2QspK23W4TKqtYuOfaQy/VmzWzKpI/y4F1cuHq4ZCMk75RAY
Add7gG5Fl32Sn6q/Ryzj4HTuCW6gGT9e2AS1sUFWnSpol81su+OmA6ZmiBJNkyZiR7Xw+teG9tF/
/OHNT28dCPMvi8A8siU1iXuId8s7RtLb3wYiTHKsi1g04bJzDaw+hZbYKzCSfNAY15Dp5gyeNn64
1zw1taCJFwWzluyqINZeWv1+2BGFSRXtNbf91FdYbmHEyy/Kg6430pmUU7cxt3rlptbCY6m1TQUZ
4lagrUzni6KTt2FB1PQLfTh5dqfxzJ1840P0ERMvxgHHMdYSi9pHXQ2OcCXOYMBlKA4WskdDnubR
o0AP0WVvlTXu/KJFYASstFz2KZfEetGOzgEKTsIw6Hm4qvqRRmcimyB1w5XKbM+V/w2kgW4mTxbf
jjtYQp8r+Lf92iv+5XthN8nJ/Ze1XNxXGDZxsjiF3lfuc7fVfGfTba9Fa1/riVRrlXLDIIary23H
fgya8TwkQ+xAd2mOiCkheulE9hbFB7b5hLJlZbkESaciWaRY1wJ2VXKSNj/OuBJ8uJUQJ8KAsSrW
3cwNSzRxzOTIm56RcEBaTf3xBbjY6exmgrYdIhKpK2QWyKNAT/O/C1XAg3wAeJV5EGygwOm8Pu14
iCvfGZRZbvs1NNS6f5TwFuFlSOMvlqiOTs/lkV9WXpCecJdGovp4syTYCgcX8CCzltduNgmqIu6i
55G9sMdRGvTiHOfKRNgmQa+Zu8AK96hBKqEhYdFoh0PdSvAT1mWzfhQNB2nf9Egl6uWwjDKR9Emq
9hq/5J3owh0NmD9cmnGCJh9/cECONVa4xWezy1LYgXh7Hie6ra+QrfEpmwsGDQIuCKtIfYOYnabR
ZCq4CsAY0M0a/Z4nCNKrgftPYLqqaFk7y2sQSj5Lz7W68+GzqB0YyZKFyDXQjrRrzUp97wtxuXkf
/iYy/4nOwJqKaIPBocCGgjlXZ+ZR5ebCBCPlac6zHAFTVGYXawZ3JmTdyJtFMZmLPTXQXV3VvPL0
eTmrdsTmbQGijuVgG5aWZUoQHfgRGninBxQu0a8WLF8hEtUHQkPsEtkHnh8+pXkZTg/G2AJIDKr8
9HULVi+hia1/c/H3S+E1dP+hgZ5aObnp8O3CqaarqDINjwlJY2EBZSBOuPSmoZazna8FoUy0AdAD
UF6I0cnBphk32KnKwnWavAG3Aj+rI3+D3y0CE3y+jR6rDVGtdKAMnoFSfJvknE5rXEaHWWTVcdfD
UWfkbvbpDcJJzobddH/wY1FLWYP8efxIID0+fMP7z52Xclkb1YmIjdjtX9SHkR2qVqA1Xpa8v6xA
4zXImimVxvyMRmItZoMtbko/7mTazhr+HWzyxLGhP/fkmYDBdwh8X4/oxXrS1kWyAHE/NhcVLiYE
TT03SeBGx8af67JWjh4jfnuX96JazWtzrJIuzGprAsyVbH+5/Sp5IWY0NHc8qQBzmK0QWOhyk6tZ
kNLzrJgH51UJvjyhKKM1Ne4RrCoSjnuWysd2EPhr6tKFY6u2zNEXgBSbToY6bTMwDjksPFoXp5Yn
VG77z7PkpZP4Ut3VASqGThrry9xyyqhEtTkDRA1mSSn38cXwi+mlLnnkrTTDP2JqwAk4WRqxipnQ
14VqYbG4PjWoLYsqSC2LIQ0Gre3qJAfrZvPz5c6ZoGdUns78qi3f/MvkZM6HKVrUnTeuEGxAqhlC
qQRw376wyei+gNCJIdcIS+y8K64g8u6SbzQU34VOQ0uk9ajiV8cydHg9CmjKUBlqY1ZnZqZYwzLD
Je/XcO/yUUFy/Mu1t47zdjiwwCI5AN3VKvDyLQBmNRA+jNFywl6KGqGUgsfZmWHthQOs4T8OyFhm
Amugl5cuIlQqCbVE6uYUeKkUKWPM7X4CftydsyVUtW3c4tY9zkrI0TQnPb4hT7q0fTcjicgxhko9
KtTQdkDIoLxn1ovGSozTwXMT5kmiiT18ZYBEP3qRaaZeTiMygTiD5oHtS8DHNMVVnBU2fggmOXiw
ABVLBW+LGImVmIaQsy/2lXMmQTcilELmRR0TKTLHrfBoZf83LoTwqukYCkHIY+mW51YwVeIr5T1Y
WdtKzIanTRvux0OHF4QDb2LOvH84Urtx9uKjBu637mM7TRTTjCofGLzkVQl5vrCY8hRnu3mdQS9j
9EDFDX0vNeU4RY8QSzNH8NGwoRmqrHKaYAjWufe81PTwepQLcTPVjTUjtOwHeqv85PwXT+tsn+hu
p4h200scQzndZg98V9WKbliczHr4VOdJgsKisO+VFwYMS5YoWjo2SZHHuG43hkhnYmS8QsqBadpJ
x+O+OOTvRilC5iFhQCfkQuETJihTFIYGTlHR33ZtkTXu7stt2oESkKTs49zjhZdnpoiG1tOvE6Pt
7weFvifdxdgOsJNN2kMnl9JfmHiAX7VFPAj1yq/Z5ERbWjkVXKunSj15fbBIpAe/1/TlqcnPzAxr
aTCeIGh2IXuyoWXSOscAyf8+g1U8+VmvT12cdmt6T+Nj526kL808TcXE/cWp4Sa2qDZlkl8TocHJ
Edrrnmphw6v+JyWWXZhxUQevhT5klCh0s42h40p4lsydKlwJceGDkMkPUXqbq9Kf5nJicyCF6axM
8IUIH/9EPSwfagCHRoQDZU6hdX+Fj8axr/uEG4u/Z2Cd4i9qCq5uXWVs9Y9bDOkxgQQngn6Stw8U
opaDdsPtAozEoAAck6eFkGpXodCt0JGE7Mr/Iq8fU0xtYLuNUcQxCuVzFJl4u9iywBhq+AZL4dcu
OJn6pOnCId7NGbwAzqB7tvHDhzsegUBokrknDOioffpV5cGIMpwOketd3BMrH2dkxm8u4FEEWVN2
EDp+HMkdebOzTcMZqsQrajMuGEmrTSTvpMQCIRGqUnPwLk7YcebSaRCOjHIr950k/9tnsrWk4oU+
oPb5U/pXvrNUMB+/wNCue338OlzcnM1o6wLQlNC3OtbplweQLHHnKGIfRns5wgDvNXjr4EpUBoyD
rI11CGH1w3Y9W6SaD105380ZhMj5eBFEEHvDGS6a3QYIrMOREz/+ey7k2kn3zVqhOBeb9lHxAhSP
XtvR2Iytkb3jErQ9iYlY5izfNvBbXzH/GppwI4ttyEHuPdIEqSN7W5SRg3R7aexvTqmM04SmQ3Oj
nbdIvzC+f1IBj+DJ1Bp0jzz2Ybd7WCRvAy9tbVDIZufs3zV8wuiNo8j7OfE/V+O02ejN8ZXvQ6g6
uxDj9mNxzGQBZB376/E3zPfUId1q29joVDmYun4z4V12mMa8A06nuLWJsFPw5rhswNcvchJyf+TY
DA5gRpf95Ym5sqfKSMIRWdBd8Ry//+KWTEOiNblfsJA/l1P0pK8no6mCSVGJxDm+ZI2R1O4RECfs
CwUDDFohNbhs4hfPItkfgL7PW3cMZb6WSMSSNsgwaCbahhO9PEHKAjWUWQfGGAo1/TiIH/0nGSPs
RfRdeTIwKKpe1l1cLyKAfIeRxyWF5vvSpg5e4cIgPK1xoywLTRq47jwy923o2y4682PpQusEL9mz
2GP0y6l8tRnDRAVLcoTG9NqWm9OOCDpMMppPdn7pcn6oaaCDJTGVEuaEWps9wDG3kUqM8xXQKODn
yFv0QY0ySIyx1WvXUleJrhxg3rGAno21TUVwzEW7rptK2OzBxmL7MDddA5RJBEmDn/c+XBPdbI0g
M2+kw8Z/NqvaroHzZquhmkTd9rHtLyN3oto33fCF0egAptGkRSbWV4cKQmnO8GrqOo2wgadBmzrj
94Gf98yJw0QxESl85Kncvy7IFT9x5un2nBjT2SK/dDgKwW/0yD820/zqCy6DK+ic5IyZgxcOhhUC
nYBYB4Kv0zubvZ9u5NpcFmc+cxPxQfsQI9cWivIZzNz7NMllrFFSFTMDXys6v+xGoGqLgLBTIPvT
o7JmixH61m2Z773+NsEAok1y1CuTjyVOvUq9JOr5bZsfo4rLgiVBMx6PM3+ShLo88zKVJ7tz+8O5
ZS13ge9sKdzlTni5hEt81LN7FmXZXVkxf09QkVhsCrYutibpY0ectbrNaRMFs8qqBAo5BO+sWRBF
0MhUg338D8Ogk23xF583BDI0N2nmIHlEhNfk2PqqmveenQlQ/8F2c/xit2eaAeQbGXNnmQJ7/tys
lLmYxLwTQyaZu/jwmBuWjNpqWpw1SFkSIdlfWwjVmJnzwgS05P5wn77D1wb8tAau79QB62QR43qe
e+IcPEsBgnVCEQ6+/mUU9M2pg6D6p047S+ilZpfc69Y6ojLWoXTd6hB4HUL1mXP2AIDuorfnBceP
6iPnFL944gl7XidRNzF3F/VOYcQSoOvQKwAv0awSXdpHbEDbf7wZBI2Vl9uy6Or1KmXw0o66jRzg
f7bHyFQ4drpwDDk4n2O9KJKxdJYwXuhA1ggPH1Qt3otRjtTOK1cBsCi4BwpdsD3XP7un2YuyTzkl
DyCIpgb15EylLws+Jrr36xLi+EUYyz47Y5GxMo0j60WFn2BqV4hqFYM+rYBuQ8PlVWFy6p8K2W+c
IXwvsa/e5xb/VoXu19/AyesCBNzGwqCJjCUwRTQaNxFYKkiK0rWdtPw8PzOLG4hbLCs/Z6dPbgg2
01LPAM7BInJMKpzDs2pXgfrcjyANyPHWKhG93yiY4mb7FKNKmjTEy7yMUogZcMFq8p+c0C3VX7PP
uxMqLsHWxANzPAXNj22sLs1MBFEd9uPt4G137L7gdDdV/2K70ujwT+Pfwqx1kPDBkQPJaR25ynfM
FBQmm5LQqanmXmF1RjKJOLzJOxaKx1kFqdqhKqqFv73nv0nnRFlTsxoVSR5aOVj0PmuzDScVvudb
lgnpmInLpYgPZLz8ntcjIo1wDhCWESmZCE4uzV/zi0vaWL8GNL3qAV9Y4wfKSupVjeRgXZlbdGuR
sP5KXsaxyZ/RFk/hWb6u+7utY0hTgOiHkZlnp1v2LYnMAA4PFqsobWf51W2HiLaUIFPi7VsvoPQM
3ZkcZ5C1BxWiLM1zcSY9sDSjqEeqzUfNAABfKRqNPB8I54VeeRR+JC3FiWruHHqPxsY4sHnPhaz1
Zqf4goXSSKY0dAfa4gZq+epWCcRvxn1v5kIZepw7m2k8Dgid5tE+QRcuJwjIiv3JRoit18HkhgXN
Y5zY4j4w8xEnwBYJdxwPLvIpGYTPoFrNGHQUCHo9zTZEDQlTM5eCaKV3jDm2ndnKpixBeccJLqok
Mb9BV/IH4H74WoIEXnyuSjkcBeVBpUmQNoiEK3Y9LT/PzRQ1vMfYr3YQUg2rk9OqZ3jrQv9hDSs8
VtWh8YfrgNhROElnZFOeWEltt4x4Bx1UXEs+KJ8Cpt6hLC2eq1ew0YMF3zKePdb82UndZldvh3bu
o4fmPGo9MmYSKl4ECAmilOl4++YLsR4ufdAsZYZGnQIcXAvj480ixvjM8fh89j5qfSHKRIus/NT9
jknxyLgO8suMme76Irfjd2Scy7Cb7fEESwc5Hu9X1WV6W3Sv2fcQTtkr6INm34VNtNI7TozqPtA6
O25ETQSflADjjIbvONmpsTLH+OgFF4ffogj28XftjSz2oE7J00I2h/aG9UAL5MjN0lxkxs+lulza
ooIEOXajZ0S3ivsfrvkaXsDEM+C/RGuwJt1a60/vy23nPpVVmd4M6EIQf0MjfawKrMTo7xoYc2Tp
Jh2ydarGe/Om3Rbg5XQDjzhoIgetY8MrQdavvsRy9BSdb4xpQIFjo1SpGQ0UovOE+Oa/DnZwXAHQ
OChJ1D77Txx0lDEgyMEV9PhLzcwjeFqxUbRp5ZI2pB9rkuNlzYeS+RcJs9W1VUJ/8cJhlBxoAANb
FEk+gg4AqCDEu7RNpwI3C/SY7z4s5GAzw36ktCx5DBaivuWmP4VqEwxf4GwESmnBdfif1Ny0ZfPQ
AzltD1RFLceq5IxQ1bxSrfYvzXANEjC3EZ0CAXIxtj0NXOTOcpYtTYKWBbGtWR1t6erpAvi4tgQy
+KmUcnaVrY/MHRWazqXnulX6aRPB8yELWZkmco0q0WlVDHUWpEjSnG1cbK82bBL17qOYIJqHLTsh
Nv9Bf6b76nRSIznwT8lMW9e/IIwLRRmPNC6NC1ck5eu5Bjj5a0Ng05+R93puV1N2/eGQLueo6FCu
c31heNlhYsG0eoNZKD7QvdNc8ad9xCA6TfHcmc14J4g36o9kOAnAfSHUSuPS/Kf6kQw5CU7YGtBA
Ah3Rw9TeV3BZHOU54ubxoc4fBcfaNNnIIhnbI6QOU7cZ+lVfI55l+B0boopkYJSR4i500uf7l/Wk
Lf2qYM6IgexrF9Vwds/R44heiBcmiGHi/QKxFQw2adbecaGOqL7Ff53h0ZqDAE/7xng3mI0nFzRm
nHFPN0x53CNNuE/OSPPKtxpJ5m4hOR2ZyxI8/tmIquD7E+v/8YuFusmjbgbhyNwN1MeQf5hEFYOt
c838Ae5rL+MTeIjqDp5tSFDklIaCn57cRo2w3t+BOM3/wQOfB2JUq5nkRWfSj3ucwWIoHMphOIeu
DetvwY25yMkzZcnX/jceXwPoTWxDqHvuV2ErU5Sm7zzEIWZpOk7Chf6Tp7vHnK3JMECpJEPPFbl1
pZ5VBmqIbT4LWW8TphjHQr8hdUEq+O7C3q55trGpwpr5pDf5vCtpcEytVtQFtrN3OTD+hkp7bW8v
QY3XqtNztJoAPAFWFRym55U+NA8iX4dvRxWj+rVkdYOWC+Wl25Omg6igub5XqFp7oyp2cV3BZZTK
nUT2qMCbScH7yCB6yV/lRcPAuck8CK4U6uZ7mZEaXIW6juSJi+f8+HB3YbniWBF0AhFKzARXDMDI
GffeAsyuLxSEzi6TGF0Pi1s+qSIya7SKLcHD449kXjIGCwvvMWFCESP0sOUqnKKj592YePS2+uQA
1N/EJBVcXS3Q521u9reWkwcpCbJrV8lDy6BWopbxmy8oT4Kei1LpKQ7t0i2qAx55Lf1ub449GbKa
W4v75HSpsfoVPY8ovGWGI1tuX6rfrZxDYusfc+qsLqvvEEg9W2EDoF3gygodkZRnETpSmRScVxTZ
ClxN6e3PcvlBY2c65optfrL/qUyCRhgZMJUEHd+sGVIWlYgcvcDLxMUAZJi3P8oPWXCoqqMG8RSh
n9Z5LQD7vXq86aNqUifsj6X6o2Z2Uw/AK14Ol4JX0ZhvEJsdPCngL7tbYmeE09+fpxxCtXwWkcxJ
GEglefyM6X/gpnBDtLCnj+jWIairlIt+AXLbj1o/5NTxyr/+E+cs0NNaLhjhigvw9sU9ljrbeft0
7pYDq/GeUiepgR638F6KwkCx0Z3cV4hZtjPK+Grz+rME7Wxe06/3agkumyecvA3Kfmjv9qfS6IGF
ekckh2rhYIsRJ1LPa+31BiOo09ke9hCKOazabmR9ibmSZNPHkFZo5zt3nC8G6U5gByAtM6iBiqKn
x1oAshzt6/VHD4vmjcY890adkKYPVJuRNqePZJKz5U/GrC1eoX9KVaLRcovQJM98ma66UIG49av0
kUtmTNi0iq8iAI3cKw1sVJMZ6KFNZmCLHexH9effbsYE2SrkQ3yaBX/vzhp8nafQLIYz/HgDrYT5
AwoQkcaOzfFWg3U4XC3HjG/6hJMx8YdgNWbvM3wcb/EElOUk5edvxc+/gZrsAlVDLDzz21nCYoAA
kSofl0lX3l1STKFlrTERKHbJMsX48IaRAUk9zLp4TZTToJA7zbJjQKAtbaVEbkhj43U6lfZPrdvn
CtfpTwlJkWfW3Ll+741npBLMn3FA3uYCJdRzvzqIE+tI41uapAoSIt4lrgWYB1H4wiZzAELyATV/
/2sB0c2WTs8hE2fqkXlDodpJ7eCVEKouOLce7uyBYenQW5COjv6BOp9Ts6TpPzXan6ICUAaqdC5P
H8mklLhKyj5JULC0uprby5HhkJjZ/QNiwNBAgKb1lN26qNJc9V+Z9XLVrxq6H31Od1oHr6CQfU7Z
7ZRq5d6QiZP5s1Me7vMguPayquFrDD9Cj7wSz9aiPpFCSzXTjCMgSlfNEX3n8a0CIspoLiaXSUg+
9wOboUtORMqnPMtN/myeDc+2iO+MoBzDLmgGlFjUnEBoNp1nhATo0gm4/Hq6+j/ECweQowZ8+CFZ
0ZPN0cUpfgMj3KxNNXKh/3x5bxFqrSUZYqIRR4VZc6OOp2C3y5HE6J0pj+XTytpHKFjE2/MxW2ii
wDqo14D+VO7FsaOHKFY2vCVYUcXkvBfdouVJL4Gj3xBv21yvMk/yitM4wm+Ectf1LGjtN8U4dfvP
d7KjgRKTmVhWXr+cFtbETTAu90BCWanOOqWm95hyY0ADpxHtlljyhAT9JHwtiCvNUot3e3LMLnzQ
R0GrGB55eaDVzybW1bIEeLYY+QFnlSjR7TYuhFTFxRbuSpvif5RFFNMGFam8o/SpegeECLO2NoQq
hUgZC+zthdsNqhslCoDjH/bPkbuUys0SimVAPBeikdjAeIvaAPlry39eRXuPdwznww3Yx+Vvrqvm
y4fOqKZXGxFK10IOcKuDPE2bLjXhfCGUjEfjfHWtE82+Fpg3Ln0pAkXqtsCp4OqCYwhfY2u7EzQY
gpk985Ji23mNTpAJCLyvH/dLjVeyZehICL3QTd2lDHjAT8ezOUoPmnMUvA5lpdn6W0lk5fMq3gvZ
uGBFsJPx85MczwHWzYitDcH3uV2ngT1tY9WXkmoa1Ki19o7YoKoj0YtK5LKWlGRuK3g5fHGe6Pgc
u1Bil5k1u7+eHon9Aw+UapD3Xy7p4epBm+LIsJOGkUMIT7oSjtG8RKcxxID1HlwlK7C6r1ZWFGwx
PMMzL/GCTJP01NME5h4Vk7f2Q8SRVwUgZh9T3WcQhwoJMlwxMZhVFG2OdfpfdLO3bvB5rh3vbodC
gwkvZgg44dk/bt09Tf75JxKBsoS9I/ixaUJbQ3okgVDCfR25CASEJJDxfxAO/dHVZpWVfye/ghTA
2lPF5iKqmXVT8PW2OHmQts7ATOhJohXljj2/pHeN3S/90xPkAuPDCneE4qRspqLqA5N8JEzkLr5i
2O1BCBRr/l2AetX+H48DQWuT5rHjLmpfycTz5/5OUSFSS7+yOzHvz2It1E7bL+gt2x/2ev7LSTzB
/641dRbf8mZM9u6R5ZL1J+ux/I4Nrvg9tvyQjdYVOvFL0Xj6iGsc3AfclJ0NSqK7Hn6SmuSI0PdE
SeeoejJAdFLTvCmAYAvemhvMwVTTH9FC2z9cSXg9YV5RBciYxxhE9P5AyyOcmaNiRLOYpVvpG5mu
GC0bEvoq8aYESwgwI6RhBt+li0HnVCtHn22BpSDXNUUxWJyiQP/X/dxODU77EUBdiUGXmZRz3T0K
VT0RxBK6rJY66EEo+06Chbj0ExgkrFMshEQQwjPiGdpCOzFMToKqoRQoUU+RWKZBy8uj/kR2OUIa
QyH0/MfNgaBdLlPmHNh+fHnDmiH5e3gCQ2evVkSkTGJJisLufTOYUTF9ICrmXInMBAyPVIvZF24j
14/qYjYWYVyiyzBOtcNKGksGxIDyNts+9zxF8swO/3SOXOnGWogslHBD8PfllFBUS9wzstVx3KP0
o8tNd+eK5ewQnhLTvKULIfmioa+9Wz/dveYr/6LUdNHTMyUC8oYcbEjI9WC6FzAIor1vQVOdXDJK
3G2wbi/j1F6mkkEP81c3R83InTQgCTrFfVw4tMqSozzLhayOTmXqM46D6x/CWTlIcnNqorGAiRsN
u5opaduV3HjCRRXYt7jgNg22flsFqcBikv/sSYaPo71M4lXVM2Yy7MqrAKjHgb4N8es5ET7ovBzG
eJyeIILs8bcISwmCt/zQWK+hiWH9MvXqmaA6UttedfBy6+xnzryxai4cokbYS6uQ16q0jyPkVFF4
YnBrDX3TMmGTykAZApT/xtjnLz1jfuBgfYr0hqPqVwHZB9inZZnfQJZt58nQkNAegDkn5b9wElqg
zJ2IkO8foN9wN4WZ1AFx18yWKqiTFYXj6AmrXU+0fx00xHqoySMh7mSSDWl592olccf5r5WESJlZ
FUGbkb9/EdlMKVq2nP8hZ1UJaWAOuvPkyoEB1Wcd1pU0jmvPaA2ecT2hi76Z/cPaQclPRn8iqRv5
f/Mjhz2DTRQQEfV5FGfPTDwMQgEL1ksHPPasS7N+OSYcB7vu9MeN+US5qJtK5YSU+MaaCi0NeyGu
XA4in9Pt6mu01/WGdtpNJDkmqzdxOH41GEn282uR21M+XBFDL89HWlYkK3ewNB9HqR7c6N+qolx/
zkTlbDDJmIcJLd2rJddOH5N7tPW2wUzRJCCH8KeRAj3PEZNise1JtAjdnkiaGIK+b2vgGc8eBPT2
PZOYoFofvbKtsf0FHSIlvB9DZ65Wlp8kEpVEfbBppGQH2zGZK8qwDiomypz0+UwYR9o50f4cnuix
tCDLWjnQbDbUMH2NzOulI3WnHom6WPlsneQ5IzQ4M4j+kS9in6/hR0gLjCaaGFdm8sjvhzDiu5Qx
WsWHC3mPcnFW8QXthD/oDPkjuctxcY+P8+CDmi05TPgWesU+nqDcm1tvxrRhWHzhP2jncDuL77jW
uk4a1EPP60YhbfE9UbyZSWpV43HZQ6K+YUEAhP0CaygDg2Ir4D/HihP7dzyKQUUuoK8q3ftFV6gD
mx2ZHnzN9Zm9J9U9nmAlMkdfjFXY26/rUCGj5z0PFFNDBqgn6CpTU3e1Oo00FmdTpvSmHNq6tvya
OqjuGySmiS4k1WPxqpeYxaQVGgkGyTC22TcQ8w5xO/p3q2LK519IOXwns5bqom3IcWmJO1CziHv7
eCqN8NhQ8tTbsSv91vh/UyRUwwGUwbvenf7oHwB//HKF2/KFqYsPgsVlXasJztorAuvTFQ/XkjuP
oQZBpBCruI6DmbDVMhsisVnTFBFi9CT2opxuMFxJzrGrjPc2ofSDI/oCRtr1YMnaF5grn4rMQuRv
FJa7+tzzZNDfoLDIKFfxViWTmQ0YeSGV8+5NX45oUQnvyARZSD39G2xlopQ2CMu+rtTrFOkGc4HB
YLp+l65lnGnLq4DYn2TZdJME8M6TLrlZyA2VXavW1eTfaxI8HtgM73f+S12WB0stsZ4HxJgfGo0g
BLaXJL4b91IXj/Y7ybHlfL0h3KXWTwPmwhdakPoLRnR/uhAu8HezB1n4UK0q2/PzCFrPkvuKyyjN
9zseYHK2h0xcvEniU2zLF3Gb16klBKET8tGJTEKj8DC0ncImzkZAGK9IIltHdWSAfd135x3p5hHP
Xlo5WQLsfFsBRO1lkMp5H5Swz6KfUH8D6lNQFWRpYJ6+2C8S4S5sVT0fLOPmgOvS7GVQvOoSNuYP
TnhHl3sArQHwwtOGjgIhWiC9GOySm2nzlb1SrtaWOxW4XErQ65seJxK3fbv9OjkKS3pW+FQVWfyN
cZvgeayin97yQdnKP4S+ZwN6BCsh58c91A4QNU+oy+sTPfjHlQLrVfd0/99uXGYkjscqpqRIL7XQ
tVgdmHmR5YhHmE6W2EXFgR4g+0PfrW41SMi87NMY0a66RzqafAF4PntdJHFgHoEiBjtKn9IYUEk8
XtXlNDR7pi/ywe28lRwfmxQzJELADdjla5pUpAJko29ZApTji5v2ZefK+s6vK3Q3DrMrQcvqA2vq
F1yszp203wWiD1+W790orVvrcbSacfeHv7ejLtHoeCBd1X4e5lQlHWpqHzg3CCJGonCEpiC3301U
magYCyhaQErMeX1d3AByATszMxxBxYTtRJ5UswCTR4I2w6OFIxviz/j4pdz9PyWMRYmRxjfXCItf
wRiq10BkLqvb6kj7VS93PyTz0j3PHXGlJuONhXnQMyofBiwtaZV4mc6WMgWAcizzHjlM2x5aotel
GaacqsT4hXKQbW10d3mc8t9DtueNZfmpcNYigDGltCRKYWuufrV3PByDlUqA0RAiViG89Z8twyyJ
S4HDmQIqkEwP91VVwmI9CVNqNFPil5U2cuae3DnVsf2nT2277uFI/U648eem7GbA3Q0X78aHEEjZ
ykBoF2/9MRayo+nd37Css7ZvSRLrj95IROxyzV4Od43RpDY0vMeXcOQuh/wmkvfIj1odRejxtwLm
/lnsJA4ad00egSqys5Jp/XiQ8WZHvimR3Mj/Bc1fCBgn9Dhz970N6p5LFO8CerEBpSwgSfeV5EhI
iNgLNnutCYhXVrHsBSpSN7vGw4UB6KRlF7lGf43EHG+c8YCQDKeBDrguNGNZ0ffytNstTCkRLv48
NbmkBkZl08CI4/MBwjodNIh9Q1sBDZj+UCySgQVE+E/bBhJ4Pj0Rj4t4O+jGkKBSPyjMppOZ/fif
cUoqFnQdfp4OmsPq+8Xaan/b/H1LbKj88Lw2zenLDHgicdEoTLUfgQNtHzWVG2Sswufzf+dybkBJ
KRj2IRl0cFtOP/HAWO76Bycjg18AHT2JlvU07vXh81siXSup63mER6uN/tUPBx9w8kRtv097eV2w
kH4sBKpbIZiSe/5t/VwBYwchqJchopDuIVC7SNM8dXvJ9J3ma6cRI9Jw9D4ndkwd6a2xH+uCarhI
SW+mgWp2rZRVxXNTiqVZntVZH4NMr+qnrIrJPrg8g7wX9FKzwttTGMioygqX2qtpRNTCsV8NOxll
1xPZ3mMoLCh2+ayyeqhgs8HJ+lZ4sLeiQSZAgjvA3/FdCJzCRHeKGxRDz8vT0h9X1VwJjdu+VoV+
d9CZW5s/fH8oIU3MZZSu2toHlO43K21/AoduQRFm0xJqw/wIiH+eVWNYbkjUV5sqCH2YDye0cn3r
YFi2k4HcDmQ9ble/WMS9yKovkuhhrl0JA4cvdWGNrH8hmVWM6TUiThv5PWTYOvrDtl3DFVgxMAg7
SjwwEorohwKrdutioic/6VtcA9fBr1rWmY4S1Pr4BomG/ZqODSrQ2C5tS3qj91tIljqW9zKPUN5R
1ulfyjIthIskbPZ4LCY27iFYIum/JvQbZcK7AjwvmT+YQSku2pvLoE4BBKA+8jIMe1je9hXraSgr
UOr2SAHwoDhWxCTlM39OKj50oduPR77TyXecTiTr+zRZ/1KLiCmsclwBJyOIhiJ1afTmRevxFNlu
9bz2+TJHxSVLJg+ZbKzNFk2Yc+NhgJ8iBJeUwFbBkZQq/01H11gnUwKecCVJJjw9FLSfbGB+P9Qz
WHUIGH+TnkfvF5aqr83+0nFFZ5c7fiMcnuV5wxGgVLRxHsivkjtq2qZQaUunKCjC1oss3wsPyLPh
KfqZ9ivZ55pFkkK9k1qtIauK+wDAv09qY0cKQPjahOVSqhpImBPPM8orCvQT9AHOdwMG5LLZTcUb
ICm/gzSwrt1jaMbfHwbEWyMo13pVmrNCb5AexvAtfMKilPh2QEZMEnT5+6B+J3ExnknJIQjFFuYn
TKvdegKfa6uovEjE1MrWTcpuUg4jEittYV5hlz0NrIIbxjcc4KDJjv7ozUFIX82AozqyHQvcXazy
56gWrs7T6sA5+8zo1C7JwJwbqaaLF8XywgugKDy1VxMkyYjWnufwlIeqsW12vkuuJdevmaTS75RH
HybxxkShVhxyLg1QE+uOYAIlaPGaukPvWmYRnhkqKWrMadKgNjZEXUN2a5f9G+sfiZfiiijHgF7K
qPBxVsn6Glhf0gjAcWNmXJzLip9/OXLicyeHL7clhtPeViyCHIQAgW31gruEbMwOcybXnli/Bb/l
y/DMTePoi44D+rE4R0jdvJ3h6mUwukRY8YaI3nTj13727WxbrqREthu7qYtvQ6XuvwbIu8LpcD36
ocHwkkTgMQNVWRG5r9Ky/7hf2LHmnr5iPt7vEorY+b/IOWuPciqnwtURhEpzqfUKeWzIpPWby+ag
YyzzpFNs/0im4hdJXVKBDI2BH3WzyCPMHRxjRbARhTBJAITecfegAix/bKff2s/s7xy0xqu6eLDG
2ZGikdZyQ42c77cqNkqf3pTgYEq0tArWb+zpzWc+MPS1ZGY7JSVfbvBmLzCE0DlQz8Z3P7XLv7X2
EuXmhOBa/zH2xyQpq7JRyr0jhpgI6AE+EujUNgaIeV+e3N1ySH5WaDILIIPvtR42OW7MaUCd+8On
6PQ9UFhOeos2TjoTH2TYaQnpSALKZeH352srvGrBVZX93oDeDHXQGSd11PG1jrg1wYWH6D9/Bj17
CKliy6UkDnNR/LaHsQMWsn9IIzYdZZbpwyKEmeIis9zS7TmxW8pkdy3J28sVUisuhxwgbbKs9qaV
kolr3bXjCroLkQTkbuJTeprG7N1NJ76F1Mtt53vwjwCN46J7P5H0OniQF9mv2fMU64lwXfFjpVy3
DQhg03196s8qS+/bY/DD/QaNWMOrlA8BeKNp592w4yld9T2f5Z1j/RYRqVg2HFngzneKElaJEQyF
TU531LMYDAxxIYlzeXe9XsU8f0FzgnP+tZKQ1UBi3BQrKrz9b7Xw2yKMAK8vVaRdmhaN857rUPXZ
xLoxlUEDn8JdnVIff6uNPYV1XwRfL5IGS8liPkJyYAyoZYEHGi8x0fEYFam7VAdN1sJiUUP+U0iD
bYkCBs+20UEUZQDP+m2lpfN2Gro5zviIqcxU8fL130v/9V0/SzNtfHVfbxW/WFfpAqoEyjgBNo43
gRDy4fLPPf0ZBZq8P23/KZWMKm4n2PiIdVxAmLGw6ye97XkcSX/ZGe1RWHjxfkELRBYT1wUf3vj2
6AUDc8kIlYHF/2sxsqAW+58iC2PXu9gJD5gzFCT8I/P37u8UohzvwsMRhUi1llUMbH5YK/3wkRqn
G9DV0pOvvtUuj5zOvHoW1Ma1oi9yNueusO23VX3rqMGUfJoCiH3Nk5u/eft4OnLBrblgJXqDM9Pg
2HbH3tn6c2oBZPmrJDhGdCcGwtF2gqLxSMK+Ux+n8u2WIBWfViYB6gSQxUmx4HnC77U1ChQIi7T5
/y14VGbRNOkqGTt0rFn5IEEGtKZVky/X8UtEwqOswHhyTYneskgCniQbDxPa5Q/2uyBTkLcrctjz
9Q0hBG20/4Pu3o5tqsOyPZEJu0pCVWPPQjCmNLvAkoU27TijiqXM+cVl0KWHUCMdh3rnoBVKdjAo
wGPczkvmB2qkUyJL6W7bIGOMtRQVb66c4NJ3LqP6u1GTmugKGOJ8Gn0ENqN8UH0XJ4DQpALsQvMT
VFkdlvnzf+M12RRhkd3BcmJVN7FqS9KIZRdIB8EMBQzxU5k3okHUDezCEzeQleJerKf+klH3ryWh
Oijj5CnRepn1p5UX066eWnOaAKCfJfI9nsZJzCA+DTxFUZU+esfdyGA4YBR0iMXR6Rujt5XwvnTr
CfS0tld9vc4cwfoIDuKETWUuEih8p4D/U3n+M1RYkytyZ9d+BSepvkfl2pvnmlTRKci4Kun5gDWV
eRr2Q8qFLCH1lDinO5Sl0C9/frouEajAkwSnbr9eSjeTKqwbT/XDXLhEJQOYi6YtCIaga8yyAacO
4CTi7+uHF82Dl6mrUI6Hc+rwCPis2gmn1P7p68ejU0UbTK0k16RDJzPb0cI/CavUIjEtFDBOQNWc
x3XeNM9M7RPHyGkNKH+SNQqmF9nd2NuIMZBNiFM+Q32EgOpxwcjCvFNd+2Tmo/h4Av8JopPJ5Hox
KnbOGr4nUoD8shjf9VGPwpsMBFYSNHQO6wNyZAJkFtw5u4Oj1wQVQyqp5BolYHH1r/In+HRRmfYz
lCnn0+9sAqvYDEg/hpUq7Eph2LNm0zMwkqSE2GMIYWFLquRcLkeE+dfMfBWkeK0W6RDeL2H3iqur
odg63aCgtyo1iEXg7v4CvFpcvj5N1ZLQMsVF9Ttz+q0xe5aSwcJe2NP1E/kFKLYLB3lsh4oNRCl8
ZdaO0uVz2DfLkkshDRAm2rT80lZAIKYFpF7rp7IB8vmhrdRQ0Q9OETOP4iwz6LFoKODMnYg3anN7
sTdXn6YcBktNoPlYs9bdFFRi3sKIOf0uS79DKMWfOAGi45XG1+MksFdu1haso5h85jtmA2kLf4bK
l20Aml4bRIwQeggGMnV2tw8jHFGQR8bf+PxYGyiw4Jt33UW0/7XFUmbLWgAIkCM/zh1pBA5soKhi
bT/qUaZDLtt59ThnYmlUWto0ZciKzkoP8IfuepaFrOb8WEYdOnB5O8gWTVlEloD2r1p45H/lpCSw
FAidwuGVy/B0m8vwBxzXk/2FT/+07AMQv6Liu36Y4+pf5Vva9qtiShrNLYYTbtan2iU3FqlpxYv2
EzMFOQjbtGZbsv6CcKUto178cuPYbeAnQ1U8YFWqc7qQuCM+74MUXwMvn/kkfoxAfrpus5Vn1uI1
fsIMUAovA+Dv21wZtAmD7UanjwfoBLpOyCdoqb9GwPqxDuxvQQxEmFOznevBOaGNRq51eNVMnyco
UKv8pwKacQPeZoh/6ubBDRukyFfmcZPRVpA7GaCBbiSMHr9DRVJQ7jTKPEtBX8OT/4usdhRV2Q9v
Ro5YP+gYWT4VmsrV4+DNukYUJ3OJU3ZNwKRH+/T4Yh+xtbrW8E2esORYYYo4hGxkF6vrSPEkYhDo
dfTRKGVFRcqEgf6gKUaxMnNMpKtlX1WOc54odwgSZvnN/vxKtxywD5/s55irHHpl/ZmDtbNhtwO4
415aG9MSR4jHje7mE1H4wxw2qCOoBrRMTX8mdj1YaSEcz9Bn9wIYgxZWhekS57g0CdddyjVpP4+q
Yyk/q7JylB/7/rMccnHHFcWF5Yyc0Uy34QNzQRspfWWkYzrq95mSGcuSEaiCvkvmvTujOvBEyG9/
hdL8zAgA8+HY6hJGBH5sFoTq2KpaFClqyAV+HNSdfPUSZmEWJ/woFDXfpIMQ20v0L99OzbpVyPPi
kjh+CQ1IQ6zRih8bYMWlBvvEBS4hD6zg1udrHCDGc51uVOcCdBzXQeqaFZcn9cCGdlWLPdER6Mus
TkohGJBP4EzGVtJTSJJPiGavupKFvN6LypBAvq13i6dnM6fEtVtrxDZzUyPWW8ZWcuaqfSfUO4+6
a1Co7MVdEzSDtyr037oiSjXgJqfqESF9QGtDfXr32mjklJKuV5jqKsOVL/djTmeyS5wz7KWIP0do
H4t/bYBGH12B4kO0zZKYagKjfl6B4VMCVnT3c/GrKix0pgLFrr19LHIxKutiwO2gNQzryKXIxgYF
nz7d3od4DYHFNw5qE7DbLyBSkE90xui8iQnH+aoRDL15XDcEylNhXbOWCkufPXIhe1D2eY2eRkJp
yMPtqLrIcaKBiZ4YggwrkJcduEtfrwJdyqSkda6+YIXgXhnQZkJLOivwbkj6rsyjkZr/8VhzJSho
NxxNiyViWaa6C9DonsmSStvx+8iO7vf853mNUb4BBNjagVra1eXqNgNrvWwJAsWDCkZh23gmJUBD
I7Y+OrkgCGbK9x+jt/fD5ftCsHoYtaBrjX9OcPhzYtLOGRhMWtR/h8qeISvmbkkdfmkf4ZSNboZ2
noIuTDzI4nA/4GeEhzjyxA+24ACkMry+YH+uQ8zc6UOi5mqFMS9ggbabRB45LECfDQIzs7Y569RG
0cekfxyDHCZhYW0zAjLxl/RHmntn7xZCxeW1aY8cEig+iA09geXjqtzl9cgNDdpq3eE47jV3DzZ5
lCoH+PFzG7Z/Fewip5RwTPbLzmXac6dPU2ugfrWoEwt3VVQkRJ13slXFItn3mIEBnx3QHwVaIDzU
W1yvds6fthhlvfD/tXYSIHQ9Zmnn9mzrzV3QI04iYhxP8owiXORQUYCPzDRnH7tSUYaZH7XaCWPL
Meg0bIyBwzbV5bGcZ6Bgz+1vtYUNA6hUYmNYPox4lEZ1gVCSHQzMpcHTuC7Q1SyVtKTNWlay6dYU
fX8eZlUvmWpuG8l6BzORJI/UnbIdb93rH1STW4QMXRuOAeizpCQg6ifktCwKVXhK1dUOv03bMzTo
AfzEwf96rLaIG92BgfjsvgwK8+73Y2bu6Vl30+socDbmf7JLdPw9nZzQ4xN3Ch2+EXc0SdLGVf9J
ehD7FKpPMf4RPzdG1JEI/ZVVK40B1gaMcy09GAORZmrbmDyqCdjgX3B15oVAEoAXUL4mKxU4X9p6
QMvDhbWsEWy9ya7Sa2WbwoiouBLcHONK4OYQpyzR4/teregShMCCXsvbe6XrLdJ8xR/BqivUazI0
wDwBMpHR+2ImU+wDLWG1hVkJ8uw5a40tDe2q8+E6Md2Obna/c1jOVNlVtvxjpeuirduCYQinhCmS
LA58P+lXhUg/QK/daGWHhXAYSl3vq3ouh9za0WfHXX8xO2zzPLrJwJwgH1o34FaKjmmx0jvVa/Qs
MlRcXnqO3HHnAnLTboJwnpvycnnmCe+kwDsBgunND2ikcrKWlCm69OqaMcSxgYRksndavfwIq7F8
uIKCkDHjXAzCFIAnGrMWUrJme0nyE7+WCe8XCMN0ef+cCaghzM+cmf6Ndyr0wfMbEUqcCgXkwdpa
a+2vPNUOYFszOf4xP97ZLu6c0cc2XbpRi+tn0GoSEObQrvj3jvvx86T0TTICzfY4zGCtCswFk5LH
cMh7bVleI43aDnkJ07G27xLeeG3mQq4GZDTpkqb01TkClY2gDnztu12EY/KdApfZS5C+gE6MEUls
eoTuo5Dob+H+LC3xWgUGVOvd6BbKy7qvv8PYo2K3wOu6Ni5JIjvvxn45no5+iPPrnfbG8PYjgkL7
TKH3SQa+fooYUcLRkLXz99T/wHe0aps1ONdNhnjHVaOi0tS17zoVx6Z77vW8kSHD5gYAsvHU6g2A
2LUBz7lF2FnZaQ+NRAQQPQhk9RAQA4OhxQRXNCdg8q8eLkIcYqIYQ3q/HhkrUvy3JP5CwIw+ovTl
GWjE1FYXPXMMbqR/R8hKBDYhMRwE7xKwx8ipajZ2kus+7fafBa1JWdiJ8V9jSOjSnDHyg6kaFTs+
GlHuTmIgWz5rArBNExg1aHxPw/hLVG3U0jcc5NLcYyuCq/RAwUsZEnYFIdCd9W/cHOr7cQKhPmp1
JS5kV74hMKAZxKHy1tnnJGfavo9lK0K1qrtnE/YS5vWI06YLUqvMRjhaHefh+xTRE6SXr76F6Etv
JOBu2N1fHI3JbfEeKPhPCS1UwjUZLI0+qqUmMoszG2nY9WhkCYqIgJhvAtXa4Rf5sJHhdV7D3F/9
778iF0x/KpxFApMusdn94tZ4KbUGLKMjSO5Fg/ip8obozTSmMhEiaI95zaXSAdHTZ9XPuwoni2Gw
5PakuD8MJVcL5jDyXxkd6YjnCVQjR0cizMceqbjDc8XLuhzT+3ChdSpEizWygRJVnpwhzeqKhl0i
15+k2Jl47gy+nLtzRVZRrsBObIXZzgCUkqGzglnpDF3v92i8U/3Lk4boQT8oayb8scOboaQ1fgkL
daMgr9EttqxaWRy880hKTekQyQ4XWQFY9IOzhwvdJvhFUgMx1NsWVV6AVFKFYzhnCtHgShPQzjOF
bjzcvC+21nCv5nsZRbNZqAI4zQNSlrw38Vgld+Tg57LsSt7gW2M7ZPnwSuiDNw7TQ6OZVIMYhGGs
JjkZgqlsFHpz0XqyMaoUmNCZro/RSdurV88o1bGrhgndgR6bfVDG3kPUYgje68BVUXxHUBgoAdAC
Yvcp7gPl05X2VJHFjfMy4PtKRYr/h22xDnoxa89tyqx3FB6jJ73XzC0XtwPSWnGm12q8qt4//m2h
sFn0qpGkIR+a0E4+DHjrtFH/Dj/p62Z9x9t5W0wRSh+8U/VhcUV3ta8R5VEdYOeDtIytvlVW8TUo
zUcu8xli1vZFJWAyaXavu9FsR6nAa6+Exz1th5bYllgIKelbT67dvBHIoCj5eEONozfWTmjF9obr
DogxM+ABsZOeutyLZOaNHNjuJFcih7cNclCJGLz+xBHDtx6qCUStXQk+ebmZgO+iXlWvYGi7r3pW
aHc/rF/4Z2yDdxNwFSZ2XuWQvhPPqYPLM9+wb0KbZq2PFUy3cR83XPN4m2kU4ZtffGFwxZVtEqLK
kUwIUgSAalIifEdNmBLY2p7A74BEGGFbnpImCecrCG6GmxiM1BMDZoyfVmCIO7fxLFMus9TIOKHQ
GE6v+jREK3DNH1Jq1ik15HHU44nvMWinMzeKhasSsOe2P6BP6RXzgPpEoAWExkjF1O1VdejDX8x6
73LqV3D8SsxJjb078CujuaixMOYtFgHQh0fxOexEvZ9MN4EhIecV4sQ+P2wN9fBD9eDENIoAs3qF
yLv2vSzhavLdwjVEMgZY3YkFe5WtGAkZ50lOIBHGX596Z8FnL2hxTFsImr2cBBGBPgYXKB71AgYb
9LGldmniG9xBoD/cCHapbHedFQibSnnxFw5q79FKDdo038wvFCpdUxxykVDG10pSj1+V8hwt+A9y
+dLqyorvv3kHTa7WSpz+XTgAN6/UYId/iwCx6SsQzOb24pAYvBHfsxW7qBk+6xiGLBqRm90tercY
UTOQJtRuBEk/MZAwwi9i0AKfu/5NgksnomnUyrxGdFDimuuyn2for4VcdSPW861jCyVoAe2Qznl9
Kxnq7v17o7tNBWHxPwLBHae/jZjOJcG4dGnoxVwjdz/z6bLaD98E7D1B4+ojyJ6eVMxcaqHgsIqT
iQ8zwgs6ArHv42FbRjCOjaeuTUoYin3W2dwKobwILh4GvPZS/dSfBtAyLvZRavpDpJp6GBDENdEB
lMvfdchMowrCCOpdR9/IFJbKPO8/CmNaQC7T9er3r8Be6hUEc+jGYmYYOqjoONz7Tjo8/5pnVr9g
6RMNf4y/5NVskywAwToeqCLG60WBqjXyNIwnkiDooYUCjDSJcdmtRVm9jqquTBgHPeaoNwVdyrT1
oKT9kM+1rrilPQtBGfBQ1El6+qTTcoMDGP/FcBzbrW1NRTMvZEZMcMnJgUXsLW+l8pS4VXq2rqlQ
GwKd8SU7ELDEoJ/QHf6/sP7Gdk8qIaoUUK/Eg1Gp/1hsF/eAA3dt40QXMwFuXJcK9bDLWnufa3zq
uznaWRWn/8dj0YDSstn99L2uJfeJ2IgxhFw1ZMV8wsG/sNSHCazrKv51H8BSLwfE/GEuHYQaV6b1
0/WmnJ+Dv72eSA3Y2bC20npc0N/VfRyM524QEhDrNtCsX14xhQjv8o4Rssvf4uo20Z+7cF1yi0HS
RIJf6/KIi/C8YZmhRO7acGpBLnUzqkmObmzidPujYj1dcBfAkX71h0F9B2iLSOHsyoUuss3BdCB5
AHg2DH8TTqarQmUgield1EiX8mrBILZZubpr2GLhlE7doOfNcvDDXXM1a5hsLf3Ia6S1gVvV/p9e
yWrXLq7sGc3Y8io8UNvOHw7RHcY6JzCQi+shAIBXe7hdqg0bDSpmyGCMAGZ4cDJuvELvqHmsOn9k
eLJSh3wSG3EBYRFoitjTIHrf2ms6NzDhunMWohxbGyKF9zbeVXcivjiYie9mcfzrfCqzY85ytc8Q
OmHZ/fPr++9Zaw8AtpsWBoWd1eyqPAMxerukH4y1WZFEfuKxx0IikLh+tjmrbinnHCqa3k7Ekt5A
qZ3PVvuxdhX7eWnLwqzoKovKq3ds6c4JMeZGCiQunLqJbZgX5GuNkNr6DEUW4vDpFOg8NaixJhmu
gY37lqoRGjV7+LzAt5QUXNiXotXBsIVVyX+xgB38aFHqeFxnQ67PqkBZSn7tA6h/sqZZA2zOxxQM
5thK1cb3+CiUjQL9Q2hWfAnKuFynet7OsQSS3zCVeXJi2/ToIrR070IZmywTbXgfeFNh7hgUfW95
TG/u35UOnbP4udCv+SxtmaW8RS5CZhxhBsModn/CzDPxt0SlQdrsvXynWbL3ZpDX6WDxqEnj/TQa
fN8h9ALiTnN+MI0u8K2ygZmwU0zaORcSqfMHrL9vHIbXc6aXyeYFKyUr2ldmqfY+QFhWhT3iJe1W
xRboo1ZRjpBciSBJBaneQTlITHL5NRbKz65htRzXvycGUhC+c1+d/bhkB96wGx+kMw/+EiF6ZIXr
3hyPGFnuxBZLLhhJzWRY0i7PN04uNMh3SU7zummslX1QiOxg9NOHxI+J9FZUqSWHor/VAyUxkMtD
nvn6CyPh7BrO1Uw+6kGFqiyjLCuWnlaUQitbcZidFswsat8LnJ6YkglVyYLf9SDvDEWgRsSXRFRq
7FOz0RGqnzUOcKrB81zjj77UrkLx6GaAXsE/qiM6ipa53XqRlzpXm62eXf8d573X1c56WaRo1B+4
TpUmRg/3ZGyEwZKHnnTlUsk/40cajxDCqnqRABbFhaPHFsliJXVVWEXOPS4egJHyntZYRoLOdCFN
HdOq8mII7M1loeUflWa/QPeMYBakjszDjYxullOO2hq+FYxdgK8oWgv1VsRzDsy+nrBxr8XyUXth
hGcRJDv/BOBwMwIABbS8Cm0ez4INQLzB+RxVlG84jxUtTdEwv4X9VZDbiacUh1oUrvUhVvzcy6dJ
KHAPrmj6eGpKBQk1ymy1xVJYcPqpxIGHCYC1hA/CI79DZNYjcCNEuaiZC0U7m0NyQIFdVCe0j6C8
rtpHeE+0lkZUqHxXTW9fOKlSwFwxoufK703kSODG24flaADSDWqC6AswoxV9/b6NcOzWhFWMhPrW
wGiWVpEa0q8zTOzo+CNUfkKJJ/NZltgHVuenZbFsaYs5vLau45VfBm4d6PYhmceMWUjE0TeRZibY
MYPPsdr1J1H58NrdQpZLmeey+/m1av9leh2+l8pHIQH/GNk0J+5iniqokQXAc8kwhrBWpKoORrlY
9SV4GwQuzEoZGsvK1loavtNMW20+sqT75PAWilGgXKQkXTeOhaPzTApBzkNwTiLB0nAtIC+wgRTE
O0QGvoyIGw9qzUK/m6NWM+Cu4ztJ3PFyKs8b6jZ6drs2PKsPste2upj5t8eyzpROZw92LNzW3xKU
XvAWgniodXEVdLBBLZnfUJnYeu3cnYnCUGfMvHBv3NVPY6nBpRgbx0qpixrphCSei4Bkx/g60PQS
5pBGKU9OY/r6NOFFJApqobSF5t24+/K4fSPD2HJtFGmJlw9748B+RIf8xYe2LgTyRxnCRELbItzP
IIhSjcJmH2mSnrg2Jmv9ZljG6Vx2mCr5tcVfFK0ic4bKEe1f2V/Vw/afhI9vWue0nUpVZTDCgVOi
tI9mTRIrs4GjavQ9iy7tdOIWGKhTfn04suSjQhfvQFvjB3heo4HOQ5jBTDsrjBoTJB/RKEWA2DEX
3aaIBI77T4IIxm2zmmFOV+GEaHKkeR/b1cUZqRhlS9BChV2u5D8j7xbn7BDLI2yTTHcfbiWLhN4O
r6bc3BZlS6c8JnsVOeJWdVrzYeN58psA62qrwmAi6PAFDXJWjKX/3I+QUHaGUzy5ZE8vFYZOWe99
fCGJAVOAqFzyhnBvTgGNzQmN7MagG+dqzo1sWOzSHK6oKsDhy2i2tgiCTnCGEg8RkzH7tHJbuk3/
edOwpDYaXSfP003hQZ9iU182+RxuCBmYD9sgM/56d/yxDQXb8UGXE267lyeGulyz0BD2lo4wYSCM
gTyiRrfF5sMsDU30z87zMW4mu1SlA0QmQJdMpLxn+qgQ2kHOaEKRudicKJ30wAEd5fToyw/VxGgn
vlCAtb9OuQewVKBrn8SbKO1Gw5Je4NrZy5/V26L6LIV+np5TR4qG8l4xPWNDU1HfRL3iOn3Ykla2
MXr0PYT9n5hIbfpLjbqOkUQN/4XE5z/wgsOgTK1oKMAAxIcedttWsxMeB1ttpnceTwxxt/ou+qwn
j54BQaWShsVFILUPsTLKcofvXqON767dL5CqB2tB5BilZOlB1o8J0LckwLjip+3BrkEJ/Woxs5KG
8eCdLLf08aGFiGgOXbGBH5rY+8ixclt4/EUgZx5L6ggVe7lEbhW4VgI1wvmuheVSQUlypGbG4XSz
JFbnKnK+ZO923YpgDT+kezZxnpghChBbcmzNaP0/MxvGwxHO/4+QEi0isaYuj+WtZ1lNXiRiXHXJ
XpXYhqst+vHdWH5DbGgOPGYsi33YczxUGcMta6y+fu85WyC40wRoIEqPis+5sx0xAY535hcaRWy1
iQShb4Sn+DBTujais6EQm0pnq/cI9iqW1emYJCaT8glOJZt3tAD/aLI5nHmsLPDAM96WsTiZsbPN
VunA/1JGvVqHRilz82gVPgg1XlvGsKm7Nt5OGS50tSPIsIl4RUG6eNtubiMgREj7EufuXMu9FdXG
l0RPsrbExaIYwHpa1ApZJUC5TUDcwR90fQaTUPXKDlVNnX46fFFGAmYmTzcav11v/oXO6+RZmI+l
zD2jtNOJ5T4dbVbS7qFunjJdPCbqBxWchfNzfvz3a9fsf9aja1cwJA/sKbgBOfBfWxJuJZpKv5sC
pKANHc0vbPe8KxLetjotyzYcb4JhoQk0/c2k4L78OzSbZdG+7IWW1VUcG/uim1r0VWGrAPvVe05m
m9qkZif/Kqq++tdqEp7WFUzz+mAkDYB3x9Hjapz12l6EPmCfWg18menvtQnjeZJz8sVaHQpHXENR
4womHr8m4O5o3Zb9mhNIkCbJYFnl7tl++3YGB6vyQK5XPCViAXBjMfpxnCDY8+rjH+QMtb3h8K9n
3C0YVo2XuEBdbI8A7Tb/PRUlWtnBJoWaEKL/KUXI9xFYMmG4rR7CB1AfyirBn0JqkEQrHH4Dz1fc
0FU2k4v/qKnCZoxSKwC+I5pV5wLQvu3lOKYI2vuaRz+yWtEE4i5ioKOhnHLqmZ/q6hyAoaLFfKJ3
6y75Jfae1khx+6bT1cJtc9DuHGTym+MPWWBNWaMLs8f2BEeRrE9HrrT4g+WUUpbVBusIUen4qswI
1OFMAbYpAqCn6JtGK9VbXt3mvNMift/akgKVIsJ2Fh7dxrIwyHgxb1Co9sJy2xTW085J/bgmLClm
cEAF0+JCgUx0y5argq21fUNDSf8HomhVIL30zPjatX0OoxwwLJCwVhfjBm2kn3YALLioiRIm/4mn
q6ek7vZdmFznxAtGbOIp2gmkTVx/Exmo1N68ZSvoLvH4Rt6kPea37dUp2cfNWcHHyVnL9HwB1wVz
q4WxZ4Z8fNi0KquXjvnurMJmg3Sl+PGye1JMX8keKwJOzw786rE5pZc3EZZMAU6GaJGbryM5fL37
Vwl+kQHji1wCfz8b8Iq70iGzeDp4RJXvDdel9pA/VDum5H4izG9mfw/F3WMGdYiu0HAXl9++MIRd
YPSrG6UCb2G2bMzQ3oBL8cHciGdF3d9uDFmBqNStQKDnoSWeatO2Sma0TGfcdITso0qeU7tXSCQD
0pO0Nu/W5e7/euh6noSYalvD43UO68+9qicfATw6WwM1igMLTY5gynFagehY2thSLiWgLTg9yQUz
mQ53dG+O4AKFPZJqE3s2lCqdOdlcs6DMkg0hof60zaRWVmNDO3N/sDlvznW6sZ954gT3/uLV2lKM
6ss3qjWKKvpGenXLzypTy0WfwMhvEGy6ZyfygfE6rC2vPzA5aUvKzilEemO7wnGZhL9KW0dfxnoI
FGdG1/u8JofWaaY0Xp8hgDTX1jEa6HJRm37LFktNnFxOPVfeBtek+LiMsYf7nytPmKKx/RBl+9bq
PJlrDdi11fG2tfhS9wh+LSbQU9V7TXRPuwzqnQGDIwdnykl+NAIiNlh67/94HViqDjxj+cl99uxN
Rfuj+wzjAgtpgtWOqUR8Pan/YgzoziYilw3WzNWHAmh4KR0b9WZ/DWpUYJ84nJexdK0cjSByn2Sx
lf/R7d+/npCjpFaHTipX6wZOH2qTH729V3iRKhAfughnAKjSdLiNJwA4qhXT2IeJuvdS8HQzz3cP
kfi+LjUFfAxKL3wMCBUjpZ/Ud/VMY8Ij0AP9Rdkd6RXltp70HZ7DrYsNXDm1Z7DaxMNVIcxnbZ/n
t4RKELA5Pvs4vlPWbotEJFdx8jFO6FkJOEKnG6wnLPtRWEVj5ZgEQScd2XZYWl3UdS+coAwAVYxK
JM1N/25Xbv4olKHscDD634WpDkvqQIlrztsVzNeBPJjoioELgrbX0YhZ/1Vftqaww20hOMOCCvMr
y4uO6cI1K6TDLeOLG1xXAPJjFT8rnC8MZ7gNeFiBDJ9ooaXeWZ7D0e8o0ecWIO9Hyz4r2Kv6Iduc
X2OO2H3BMG9nCOR06n/BK8ar21HuoT7qDeyEOEuYAs60+muOdAAUA0YPyZRRm2AxwtyRv/AAhuUo
nVrFfmy/zy15tQtNhF+U7n6mgIgtm46IHemWn4HJQloyQ3XuIVOL+9CcsJIbcr31slocUlAXVgGa
NpbU6HoirGL+d64hHXvtCSGowxCzUi0NUeJJbL0e1vcLrWqhQulvyACLu7K3SSlh5XCB7nRGm1N2
N+g2aNUDp0zWCW4gMrTlxX2fylyGyMPrND87klzNU0gb/pwa8x1ktM95ZD1pnMWzUFwCdkhBsyiD
M0nfmt0vTgPe7NPi1nf112fa10+KeAMU+q+VAwmWkLBv0i+J4GSoWuCIuKnD8ZZwmLz7FcUo8ydL
yXDRdwy7Ygsd6lYLrmqz7QXjDY7mvOdA2Qhkw3uldm1oza+L2Ip92WnUuRPhg2+SiIyq3hV0qLUp
iGtIa245TXEWWNqw8QZY4HLsMsDAlUvqDD78Eu4tgFfeqT1i8pE2hR333fueGFp5+ts0LGB6gywn
EU9D9DFJV/FGOXmwlW6rApimq7lUknMMBjhMw5AR5eJfHtc26zTNCyiQBGIVAcIXZnMPd5C4SZQa
sxaFOwgDn8vDjUcjnErHULunwNPc3k390IDwxujK9QXcOATbkBKG7U4YLc5YWcZtH2HzviCIBgQQ
nG/mA8y3haeYEch4rX04zIMfEy4xZDTPBx+jSpUFtFMzoJQkr9yHjtVvuEe+tQKI9rin5SwCFEGw
fOw/Yr//tumshYMImLO2Ih4fBo0CsghDgmuHAAWsn+TeDHFbNhTY8bhvQdzCh/MxW4jC1NDEn+QF
xCQhXV3921y7Rrezt0hHCvauNAjPO3SNF3llLoCjWv3ZLvLXbDIdccOgPL1DakUTjkWzn3QtYrCM
FToVCT0+Sh+C2otzOv+7TnzcnhNtjTwfCmRIwFwvTb19Q4jTpuRuJ32jefbNNaA0QCBLpYqYi2v1
mlrvenFnlNlpE9tM9rD7smWEw2bPboYuQn2gz9a3liB0c6rBa0WkZNJ9SF6M7dpgP1ZHhxgdZ1H3
z/4ubUjWnZVonsVwoek3t1ywBSkHqTOvyHg3hCgopmELutfxY+5qIp0kSwWm7NWYL2tCeME+EPaO
quYBH5hrRJT0fzINjxKwxG76wcszKg3QKLMrJhta3NQ/4yu/0iqS/pRfIWoAcQwLKF/CcdElchhg
0FGkpgVTGvN+K6blF8uqkcCDbrDFcIbhWaeV79WbUOVYI6I0zrGTQIvren/OfO/NpziheNQkHhhU
bDu84S1pd0z7en5XeWohxppZgm6LCTNXCDg5zAOtl4Lx4jJOhAXS0orJqRzZKsTM/d7PLvF4G3MV
5g5ovqdSRqQUvPbYs834y9JjfwG1fGWgzyUYS8j2KKPy4k6CIKngJM+9WkK1OY+KhQfn1X1Q7tRZ
YUtrIaSrC4M+kNh+uOpLSCJVVkbhMjqaOqZ8Z+fhYyYU6t46cjnU5MpGjy5FTWrMsTV+9QVCXXew
mkvKEIykRG5fk+P9/vVILNm1jNHbYW/G2UdWKFYHMdUse4SXeiyEZnnrA0De0a+vAbDMHSAccNTT
gianx1Ku5gh3ZjY01/ch1SHTuwrKZJ8wku1mu6Azapz765XMGecxIMPakrADdVSObNteChmpmLUT
U46sIisokEC7rRndROUaOu10lDao6ODjrKavc+kiFni6l4Z4GpY3OfTI0j577CRgmoDVjTMYktKD
jUoNVZg758EDBXx4iwTAPlU+SVumwQBJk9TQa4fzzK7w/We+9m9gqi07qJD2GMdJcyaO+tcYI0W+
OSfQtNLGnEch7YQCFI4aByADWaMZBiNP1+ZR23V791MDN7acawSVLQWkLEp6gp3s6y2vF/81nKOg
vuJDLoWcpJRmtdN9dG66mHOFnZTX4hXTDHtVHbS6EaGj2Nwwt/UTJhKAXd5XM+FxG0DDZpCGRSEY
xRxENIPXjtg1Ag875HihV7RbrPlnngqWKwMDaqB7+1h+AtuNY0gwphiXmpIYR5x4CynIsebL6Txv
9W+upSjuvjrb6uWerzCC8mgGlXSlVkylPKDkgWzrJnNS84HcsTq8ssNXbYNIzxTP4SFApOzK33tp
VzODDoRts4t/WnFJ/f5/VJQwXksuLk+OE/vzhbstP3WTjTqbP9URhjM8+ix2OfcuvuDPX06LL01a
L0rHunbGUerJm4bEq6y6miW/aF0vm2+vyTWNmAEDEZU0moFP+ElQiEd2CLQBQpIFxGMlJr+EA40F
V93fiGgOLL/bnQwu2Ps8tb0O8KGbO8HrtavpxIsBFEcKmrB4XO+KbGaM1wF02emciKOBP8gkUbFb
oR0txGIPZXiGT8Rci8jLfTf+oymysBd48iObwOGeaTnRPMs9AwyYVxJpEZ1efOh652j/ll5/+nsy
j+f0xazwX/DFtHjaMahPEtJQV8t/nYnY9HfzErIbWFDNnylboe427tEBKTLahLEk0tWXAI/bUHs/
L649bbitdmDSWIkNCX59/839K7znx7b6atqbMN1s2BiPzVg0OyFrP0vFjskPGl/9e5UrPd1wLvOR
bJGcoBXn+cKcW0sxcN42MHnkyUqguYVkB1CjSDiWzsVx2vjE98vopn212+HtUIvruluc5Bfr/ewq
7io21+ILrqodYsU/ouU/pX21EMCwU8M8rAQm2TE1IngyVNBhFU4N8dO2IRUzN3Qe9I/sE9Onwegx
zT+gRayu2XI3cw/M0ek9OrvLcNslqB6PCAAHVeUZe+HqhGeBQ7taSQUPf5LFO9gbINmwyaPAHDSZ
ODJBS2UVyBUJ/hE7pRwVqiXxziNwLOJb6ZQpfZyEOaZFfh89VXvZRHG0v3VrIvAGzuQUzE4/GdHa
brbGl9JDjP5TjRV0Ui6qtjbK29PlcNfV522KHnn19od9xjwB40Wf/eMu/bC1m+Cac+hE/o1rXdkX
X62CKR6+RL45lBBz2NFA+vewD2UAV9VM3pZ+U38jUdNyQgAkukbjPjMbinJlN8bSnpTTpRtwKBis
bdiEF85UckU/0OsVT0KbkQBtu/vuePi8MbeHFYq0wuH5WeZLXWuvt/WUJnJenaN3zrAAgE6l2cnV
AmcvNfev44nQMuIszHYJlaptoGCiYIVm9F7VXCDl/gFWU6Us+DIJdD/FVXN25kxzbTtihv0vxlGl
JLGgzi3/F3E3pYk4MKv7Fm31DlwfHv0Yk9T6FjZ7o2Nt/39oe5S4JTYoYKiQhv8dtZGSK2482IsU
vxZNR9bXqpV7ke7kg+101vZD7l4+SzIJE86JlH/IzULiqx3cmvrUXJHql93NBbJ8A2ZWO07xoCv5
Qmlx2fVAkvMe4TAXDEUnpazfoc0NfZWG9YGTO0lhAQwNmU5s4xpA1Zxl+2GR99+0vd0mz/1nqjmM
x3ZIcAYMjxh9Xa406PZalHQz+GPxGD3J5y1/87jqJvewAK++4MQWMbHXtJDN6ohYOOJ9JPHM24sP
XXFYcX69jbFQLiwRwP3kykzTKTBSwlZ5ib5UQeO8wB5ti2LmHcJtLrin7z3WPpStKxyAs1quXoAX
Lamt+f6/tPLUdplcYpucXlrD8A2RmdrOhHaYyT9mowhGek8P7wXh4a6txFkio+s4hDHIyz5fZLwB
xDwXdC9GQRVCorJzO/DJezsBF+MD5IbPsLK32HO26IR7khVswiwKZY2zFKoC7UFYhG0TrANzAFhP
MoHyHKPJYPxXjsx9C2c67iqRWa5hskvUXvKZ9xnhNyYQjTeDcnedqt1sZm45jzpFm5G85v0kwf1d
xW63E+YCQHHyyu7j9N1pYhXa4l0ADFzL7cYL/HH903elhxBzqbh6AeFJLBZdM8RSbcDn8EF2oGnl
Zw/LjS9bmdkovUtT8FpexYczWjVLeUvapik632lZ1zY0CcSlFPWtssWJpJYkKlAP4Yh4lzWP/JJt
A+397+wzW4WhWbxtf124UJx2U3LwwbBpUJwljMbDa+N6gHnnZBFAklROg+Fy2ncA8AsyBkoF69gf
SV+QsphkYZmSSHU9z/iuqSFppHPcA1M69Eum4Gh1V4KRwnVTVXn/+mzwYO8a1I8ErVVGbR7/dRHS
V340pu/v15ep2zHzuoif9i1lg3pFkwYCUbSvxjKuEtoiIXJx2m2S1AZF17fMYDJgQMHETlvfdPZT
cPAZjrpzmudVRK7Gxq7dBwobgdNCctwnL/pVTVz1TMtRRd/Tf1lmYjUbKQ7oIbfRKKp0Q+RS+bpH
wDYOm7A2VxRWdoBRzet5EZe5ULQMh0OXLVqiRGpKErw0qB75SiLRg3qNNbBqUWgweBy3BXhKeJeI
qDdZQbD8eqOMI+Owqz0PPueySD5IyLUZEL0bR2ut9OxFDsYo1D+XY2O1mH5BwLUa0OCTdwH6sWhl
FeavKoya9so2uyFP1OgYKTHZEMdtM7f/pCYLGyLXOIX3MENC71IIAnozePj35aOpAjtzh4y8PdJO
Psjpt2n00Xs7WZLjEYyjOXu6x69gSaPp/dx39Td1kSgDcVYgZQcicDnCoX6em0U7fP5zFxxanUvt
0yK59/R1ewg3IMbJEfWKgrhHOLTugPKy52YdfErt7QWtdhEhf+X3kQwnStNB7wW+keTKTI7kpORQ
wHIaKJTgHtLOOGGcR1oRaLE75Y43665Sq0u/+PF52o9PjVVh9fGZNnH4x4oM/CSQPOvT4k8WVb22
IwrKW9jNbdfm7TBWUtO7I1LojKr+yupBs9E7J9diNHayznIv7t+1RHzB4je8Mlk6j7h1XCrIyb3X
74+h/JQ3NM0Y3ZlbarWJCjPb4QybyxHwSWtSrHyLdNfc+ijEr5jyOrUibFQZmWQbfopK9H3cv+4u
oT0aefO1YgRsqeXWsqa0lW0Fww5a5NUxN80CCUWmYTJ13S3EK/pNwkbf32qI+5/Po6/ScQPelQtL
ZQoLLolu85KbvnogMN8znbJcVmrolBcKRVHkXgWprJHK44pPjs9IxM/LgMuGkM+d9WOVQd6Kldge
VI9J2sq5gKL6Z+PciMUazldDciD8K2NjUcJGFSuBJl2Y7lnD4Rb6LFbRIM5v8lZ0HuWaHkkTyysM
sM2PA9PDThOgVcAPIuupwLgC4DGLdx1hgcvBIeu/OhDK9bMIpUPh3Dx9a0XDvuiuob8jzthkNak3
zW9hUsuLtvyhW/ZnCHEP7uPgkXmbkloygxohaG+XZI0EC/ME+AKCB7vvJg2uyaiRC4CCbDLZwIeC
q8UUq+HmTjZcaR6YWlZVGvScLd1WJ2/UvLTMvWWOzSQR2PC9+7Qh+KZY9XafxcGin3Y0YMmD1XiC
qmwn1KaO2GfxBunjnMAIzGYZ8OvW+ld28lft36SNMXje2c80r5JqWujFUwhF35bMI7F/SDL65IMy
Ufom+sPsFEHwAqsWJ0KAd+w1bnBBbr4KSfElTCmQ9jEIf3kxie8z/3UL+8omODJdRwWkPTBhBVPR
GoLOIWz0sswKg7AkZnTNtC1rNhYXOBElAkHHxV4wVVTpmy4uJSmL1GYgntsPAKATjmTS9B65foep
I68fQWiztUy0HjAwH1mVWcefeFEFqDc8/wcat9uAUeznvoB2xm41eVvDr1vnPI/HMWk0FrdZE5hf
d2x7fauFMGVID3tglJwagVjhJEB/+tT3KNZySODPt6Lt4kspw8k7ln7KUnXcu/Uj1M07POT8VMag
mOG79wF6fzxwboQDnB2Q3s7uxyrEczDophVGk7OdN3L8W3PAhLLfSBHoYTnhxJEH0J66aEcTj+aR
xht+ye+50QcYaOfI/D3/nGc3DxOsXN38c986VPnYOLLYYYeVegFCUzNJ1QHY1Ix+VcQBvqyuXRCN
Pay9mfFPUTOAhi5RCq64f1Z3pYDXa6yZk/qfnk8rVrR0GML0ighd6sJjEAoL6nYciCtkWC8Dr5jU
F9SH1jMgzWMO2xm5jJppkiPwdv1in21ZJkhTdwzby5S6oGc3z5/ZhwRBtNSK/FH6lBm5IYGgSkVd
PNEVB3+uksEuLqrslYcqUtaEFoo21nb/Kde16+wP5AC2iGqmUFHlTpWkFeyjpe3ITvTOTCBYdNXy
AUCK/NrTGOajy3zRzXeB8TFSTsNlL//kQN5Ou5zs0fsJfe9xq0FLZ3a80Nj1njhOsHpWOwcwuAZ0
ccBbuaVX2RJXJ0z3N6LFe0XU/I3b017IIi6uMvZiY9kY9lwBR2MIJUI/P8gPY43ZMX477WzvguJ3
9yFagvg4mCRUjxdixFY93Wz7ADWvwgTjnJHE/pcfJdjGsFJbfCYK3aZMq1BQUVxRqGL+2EjpxWT1
fv2HJ3+tOUPat+xvCfNop2qvwUSLaRZvyhRSNTsMXAwPCE1ZK84pNNHV9qqgDpPMq0eiwgeAEn2F
kKXVAYAfccYOdi1HDFPI22UBOCpRLkafUsWhX+Da2Jemm21fsBiATU6UlR91RXY6RSipHT8vTkSP
ajHWJaSJU0oIRq09zWmvWeLafOlkFP73r43iEkJwKhX6LIjqAXwu2KXIRv6EOke1hAser6cSjxTm
ctdVhKTI37hYAH5F+Qdj4dNxOFjaHmt2Vi2uz5guH+vT0pJ7zICaFy46jzJnbbWhqk/wjAqi9jb7
OsYFsC5MEQh5391FobioPmlYAU8mnIizkI+WDwtqx4fBx5DSI0A7gMDVhg+2X/dXAUOjwQN3+vC4
HjkDvLmqi6cZXm3lQCPBG0K843Q6uL0BVkJOeYyCDWoiY+RRDKx9PMSgv6h7WMMQLDhamsdJJ40G
/vGwSanAFzzKdNAR+7zcURqoAlyZuQER1eGZgXDQdGE3x4TpKJZx5VfzXthItEJGVl93sbqojuzh
s5UGmz2MsTAUcajDpw3c9ctC/sak+NCJ3ygprU1wZGgXBoRZ5tynOGPc8bhmbyfuKeyFk/spuY64
A/t7RSurrjENRR30jFdlG45sJfy06KdGnJlpH/ZiIajHHoR2rmmPY0bQNefdjV0IMimGn0fTXiLH
t1ii5Az4RYQ83e7DhZQ0pNqrdLvw93XCwycGjtY0Z2ilPJctbdyoDNNPNFloql94rMW3wN8vvkY7
hJe9HhSb7PBQPoRryVIFwIvqfdIsOI99VPx6QiRA2VMZ6aimx/s8Y70Mg2uqBAvt9vnslUiTHlcP
3QKm/ReK3R3sAwistOl4a+VRdxoqgj6Jzr8cKZutBcfENFI97Is73iItn2LP2zZv88C8DxbvJk0g
AynWEb7/y1GcPQvgtdj8ucICpwGrT6e2pqj2FkBDeHIy4Tj7VZMV9gSBCsX/nf4ONd7Q3e59c3rQ
PqfIEpiO7U8nIdNE6dcdsz4PmaKStLcZe6NiljsGEoD9ziINC2edpt4Cob+vHrELeddSxJFwAK30
qBBL/VlJjeN6Tz+7bDRd6KPirUmicw4/eewo0r6GwRbqzj31UeWt4RDA9pKZ6mGhLoEQu6+fMyR6
lVSFiVgxjQG1PiSdqPTlw+aIgrWb9CockmsZQYdUhXD3gqeamb8boSIzFT1DWHYndW4QunFuFa4m
F0PwthdWJSIt2qdjdydM8IVIYMjKfBJmcPPHS4Xv/RbR/+4YTTmm2A9QruhpXOFI01I5m7GuUSFo
lpvQbLDLALOCOMMgRr373A1btqQn+SyQxThC5FriLEl+a0ojXDplb/A/+rfXYCPkfINm/WX4cd7q
qwcRlT29Azw37yUDv4nzGWWzg3NAi++05oHhzQKFjk0+2+O5ez4yF8PSpqZ/HrFOFhRNa0gUe4Y8
lWDTRQGfWNvb+72VYI4GkXhsj4u3bvneSjhNL9P0n0cBaPYYaRREq7A4RrO0yfJFno3oPBOsBfI8
w9udyRKRmsp/2yeCXH5OJFlndnclONn6+uEVIyEEZWjJD8IpdN7vUkpD7CaSqXRgO2EW0HD2yIS0
sSLgi6E+pNXi/e70XQcOcvIUWTWzCDAPkFQBLZgMesEymvIHSbBURLuXHBNTF19kGS340c8FPMm8
Xal9WH2jxDbcN2IKnEv2nrt3zeWMFDO/PqVD88uQZIB+Iwd85KmvX/JFeqAEBm/5hV1098ITV2y9
kFvnR6p4FWYJj8i2qg+TU0kLbCWZqfBDgCj0V3bAOofJuei9Ic4AAct7NDQ9Bi/c7+BaicU8c5qr
weuUPAb4C1mpGwwrM/c8j9Jz4r4C3NTJy3zy4jaOskZ3G+gJQaxp8PO03NFb+uHcnti9/511DDQn
rBI0zastwVPEz+4cYoFr4fB4/7NCxiVujea3BhNot5TnvA/Z3L+H6J/c+Eqt2WT+PA/fqUiNYSx6
oxB3lsb57Y8A9U03vKz1OhfCfhM/ME6s0v4ZuyMsXz8MytefwvW0idIHT7A9xTdoEqlPpvsw/ZXI
rXTx0uQvifyjeL5QiA49/EbVR2j+ljOtjxGRIfJSh0t4kMiEytwkoQXvsyIA08mi+NzDD6s9Pb+V
j95g+JAW32BByl1QDvRbV66i4ZOTq27zhwDmiBxdeRzOR34tZqovqAngZ5NMvaBD6kuT+2nrXTn4
hz3UndSNWnFN5kltsFmgz5Z2R4lF+UjvnBxnLDQm6L2WxU6UQg2R5P8Zn9JYc/0wJvcRlCa9BwRf
lAiny7Zf65LQbpdSPxZEvD9vL8CyKgoaOaQuk+f8jIKdJ59VKdX2mNtKmDxMu1Vyea0HzD2Wn1/k
2wpc7zcZ7Fejx5jm0y7l7xEuivLjc9N4j2RsN7cXvyDLIlcZmx3jTsjZfWD2DeqV7+rBeTZ0+kTV
JQu/OIXtmVUt9xAQUci+zJ+++ZQnHGCLvXy9ZVUCRGgLvbjmarJTcXSWWLGFCjM4rBR+4zKskAC5
mgQBtADtQUqiowO50Sfu+mCYhYkrZ9JYECHDGSdcM9/CYQdB3xbBxbsZVn5JHoQJMQ247HnVQeST
/7tknVH22m18XGQZMGvUrXU2FXCz11x1BIvof9uT12n0mPQ8Ku/62sjK+NR9tBjz99UGu73NaDV6
tQHoZ4G0cSqs2G/PzoqstGvy5VN9C7X4hoHt683aTxxNPhljqqxtkEVdSiJLBJ5NqtlnVpeDASGj
FeVodijtVnEGQhkN9T+BMfCgD7w+JpF9Rx1dIlu0SnK1Oatw1M9Jxm6yNCfBnusinwqdOnaC5Vuf
C/1w9kD4Sk1gkut32Q7kAR9XkUrDQveemBS5GVxi36CY5kuOU9w7BtDtJgnFFjaTuNmE/is8YZBv
x2Dg1hfbZunjbbfwkesWw/Bjxch7pmjImhjywKSCuUc4YSioFqJP/daWrqJiPZMYnsNKyl9IFVv+
t6gETMThRmGLzoct6vGulqol8JmxDXvuNfxW6AWC3TYxhF0qec1WhQVeE19kH5ncxIhCcFgTO3jf
Ft6s7J51QahHkit8+zGmwkjuVQoU5XzK+zewE3qO5SYjxW8kVw3HTcsTPkAC2jRv9NCPLXQRSDIJ
G5WINW8Qxw0Ssyvg6BGW/hFQc+UO/TfebEDRXFy7G0BZtENnr67cYnWTUDC4xQs7WodVA7ZAMdJH
nM8QscAaezMmBzEc0l8gSrP7m4LDPPd4cFwkM1AHbB4RnyrlOP25l//sooqZvKZFq3KWKxvNVlY4
lqGHGxWlbCc9Q/awb6Mtw3Cm+08fEsb4WSOouDgLtO7TKxaPeC5KId8jCAkQo2qTFFdFvJ60RdkN
kjD438JgIkV/ls3WVqZSn9IO/LVoahjP0O99NNDv0N3Am8F7vllyOdRF567cL73A1PfHN2TEu43T
LD1gttz+yU/wK9vwDw5PgtyzMFQ/cp2smRnscGChbjlwxj0e+ExfunKWHmsZxHjCegu2MF6QFQ2W
1lV9HNyysIBaafpLXgN2Ft+BkESJCvVgXFZuCls3ihy7Qfx1xFwCpw3o4Y4/YXXuIIIfg36srgAn
6fSDVXgRost7Z+4dOn5ivpfbluOhpaN2k2cqcGH6+gBq+uYR7t0NRbHwHaFBpNJT4e2rLZnNqdxe
SYrpXoc/ZpC4rT7JGJaXhjohOS58DxgqvI7IreYrKYtPx/RKXOzP8k9N355XNc6hfFtCwgqUylPM
jPueFABZ43bnjsKgjzTqhyBXwfIj/QbhsNfaBQBKXvRge/vQwP/vkKlQo8CvnQsM1Re/jZotcd8t
y0CioA06nQoNHMZztOyYL+E5co2qhLIpUBFq3F8pDtkGnz15rWrUgTly/myLKAWUBbiTMcExm/BC
Y+u7iHrg/CLUygpEF+3xSy1ygaDIvo7PyAqnSVrjwDlWnhGBKIGjbWqv10Tug7qArPVQyLPzHFkR
2mj8Tm1O25SOSw1WobNmfeqUU597/7ZdmnRXmQjA2K/ARk1rcNt5FZ3rNuuzdbxaR4MH/hzohuvk
aa/l5SGsE6lw/0+KgmDG7M1GSdAsvN0uk9jGOX+UfvoLsckp/bx/PTzNRz6wZPkiS+Pok674ELUG
C/B+2VWPpVH8OdGNvq2BOlZhclEWzv2Qj66e+rO8mTZAyJJL5Q7NGTv++H1YPL7FeROpwucXRoe7
eMczaogdyz3U0fKo4UZnsVLhXXSfsBEqqzj+P0x19JFPHSQvf7Q5ZgDeOjZtGq0ox4AsoC1bhi/F
W6FSvoWrCEKS1jUIUc2k0ZKaABl3IifhfzG5gaPd4ILnF5KrxClK2bxVNOmC4EuuPPIyCptm79zj
U/VE5pcwhnh8xPmvUOozdHs0GowJcF8ueIAHC4aQ792rHxVh4eaR5NnYLzkamvDjASxvJJpEXSFs
uyr+Jzw4x5jzWraXuCOOgzKzCxtkuh2Paoq/ym10Cr8wv+c4S+p/QMa/zEuiqKsyKiQB8XabBFSf
bhbSqZkKYEBy3ObUO58nqVCCYkHX27fHFqBpYA6S03fwiyrwCgbVRDJqCJUWsziOPASZ6LG4YILa
uLXZiddTMPwPbXB7gF1h8aL0FbyXBNsv/7uCewiMzLKqskmscm5e083nB7pDpnvdnmb3gJrNWebD
7v2WbU1btXvthG4TzRsLlwefAp6zU+UoKnFGUCwyccLJh/GiqLIKlRL6/Y1KinpDv340SjMiGZGy
QbCtxSqx1KvvU5wBKQqts89ieRCzWhtmdkC14vEglXTf9muGVOUtCUIkN7AXA0eABKtTRsUxkLQr
yXNjlImEyoKaqjwCvekCm43ORBaMbuewc6iW/Q/5ko98OR8EZDsJeesiEbqqxWdcu7mG+HFjhYjo
9pBJbdES0wR7w70y88dXP/UzgjpHkQsfvzWYpDlUJbbp/+0ZM0heHAfyIF8UgC9KJomrHUJPRMab
chryP/k5yTrWT5rkKMGs2n32I4YTFvsli346NYnem7VdWUinL8zxdexK/PsoeOoSJw0sjUL2rlDZ
bkVWqkS6Dh6NwHIHzZF/fdjIG4wlniX/L39mp7KxhDKLuKS/UHlcc5NfLHZfyNqgU+S9myfSFk+z
TN0TITAuwxUaZC+MJG2FMpVCDuS6sU8wQqlj/8IWKOT6kU380cf85NT/OjrQiTVT5VnkLdTuFZrq
FmqNBQ57WFzQ6YNee3LJdSlTGGuGgDXTD2orTIAGI4PqL3SLw7W8n2gtrSuTJ2XoymWhAshWO4kw
Q8okFE5aoJ3T4in7/gmhQmwkp5r8Iu4jeo6ouCFSgw0tx6wgVGE7V8uWk6PMDyL1hPYI2Uutw2su
Xno16MlUHdajF6Xl8GjV9q3URQyfdxr6nCRjA3t8BzrxqkybkuFRhWq8TAaeznFK8kgd1oZ/QO6m
0HB50mifupgNZ0f3t0HiG17hM1Au8suBt8QOiD2sd7VWMCGMi4FfvwU5jxqzTdQp8JZYqJmP3EXq
/taw6gFD35ITNLiflP7xFCt2fbtFstAcqXAHNNNE0Ig9fV1b/UGhCBD8lRco9eaZMXcOVNBwwRh/
T1N782iP/S2kwB5cwUli8Pl4tx0ezClEfck8oBSMjfh4usVxWkKHpoTPU1QqviN/rMZTxYhlZgN2
eJ+Fu1nFUiJxoabqlXl6h4uIuszCyINdPjf3pIQROBNT/2/WJCeIKFw+aHn4QnAiPxmirumFyJvz
NOkfacyFKg9NLNbnmmKRLYYTNJcBwQo7Y1My/BWMfBuUrZlhE5BENSTyTjY5maq9qH7odvk7jdAI
EDya+T1RGzNu73cu2aqfHOSbdY1LUKRvL6tHMtholJp2v5u2bdBZUMOzGE/jbp8oiUOo4NGPFJkQ
Qsfyzp3gdfVNJDAmEbdAWDMEGt17qyTxce6h95SxqQ4RugJd/8gbBkGlV0FnUzI3mCIKzMAbrjt4
yMtbVwnG2+4S5fMeDgSIVttQZAazJ1YdWYnMeSYba8JZT2BvWlFjOt7Dpbf4WKMBGkB9pB/A2lcv
Ru2x8ba3YPRj/nWwbvF1+AIwuZOeVk05KH1Ll97sTcEYOG3EnpZ33mZVPIXaacOp8/hw74qjNp5M
4v5dty+kqXJPwr8g9QqkTzb2V6Pyge4NnbMcL6VM56aOrNlw3n4mTX1SfsGSR7UcspR3DYrJd64r
2KNXJzgTK0PI0MBCZiVQCb/45G5gWNpIgL1PlaPO337614GH+7ERiohqYTGRkHqjIe6PVCYtyw9x
btK0ClUmIlpQ7c0U+ID/dF68n/XXX0IvWMLiHv7GB6JQaPonfy+Ttcd8xOybSz9EPJ4w+ekxWjsK
9vU3rDEr9l3XNFrGl7H4FSNFhrEQIT9Cprg9Tp4U329XNEU3IloRyEqKfynMg9McGKy/14xUPvAl
+jU8Tb3atpc/FbZnCPve05VgoGeUMnYCQUGOutkW/1j5kfZ091bzHINxHfFObjXUCoYuFYzk2pgx
EoKbDlMJY6pNlHQ0DGRgjICMKq9MSfAEtbgiZe5tZoz8DGw0W7dGFLr5CA/n74g1jv1pTjJTdvD1
HVrchaDgOVcB8iR/rRTWWjjouSwy2KbWGmc34xN3zBOTIKATrwa1WuhkbDbE6k6CJxP7e9KVfoSA
ANqJ0AwVM1+FdiGvYI7sBdZ9g7tQia4T4GVsumlEc2Aw649E+6sM4imLfc2BJ/HUTxn7gp1rQB8I
YVXPG+ZDYy4lyzJZ5T9WiyyIpdbv4ZEmxPKKEWysjIJLUF4XmeOO9gd5SDPvfezUXMNJUQM0ZYTz
8Gr4+cFPd6N3dB1B2HuJhGBOpDLrfIwNYnlIOIW5/JmY8PAREarbViWzPhEo1zuWW71Rf0hFS2xL
e9g1O1Je6M4B12eBGhPdfOWxQ9aXyFHysZOdYvSip+8DUQK/x97cZ751oWtzs0udBQIIAVZF69ZM
2e8swxrV40AmL1OLDz705xVbwjTDjx3Hh4s6AJVXyysrm9rX5dLSGUzlJs87viYKMcqH3vsFF48n
GiaYAYJaPzHIDRoUQyX8IOkfw/qZN1qdRP/wK3nCCxhe75ggbwlr/2ehjCHBLO37gsFEYA5S4iEy
z4L0HwfmrlLFXCjY+1zQoE3PnHwWaDaxapHdiReg5SFbl3OkwiEzh2aV9a2kZ/AcksCHoRsK7pzU
xtg2b3gZYSCSrvVviXCGZpb9WUimy/l8EWCAwlHNOmff4ucb7BYFIT2AwW2mYWxLAMFS48LnhmuV
fPW72bPePcoatJImx0BKT9hnUUpXkjEyRghUz45PHuY2UycUohjsTtzL5NcBlCidgwDkqcLj11dZ
vLzMm/r99Xc22bfeVGNPufeJPq8g/did3MBaU7y7Li6LYTtINHItNgfyczF38SSSL23kDO+d6ecp
XG/08ZkdUTPxpYQF9UwZF5FZbHP66KPmZUNJ7AhaegB4T8EXiV5b/ZIE6Gh+vlR4/VsGpAxw6tKx
KDhBazFnUYXrU4lCfneECoutqEU5WXxKBVUAFw6bNriAasJesH8AEIHR99uQzPhuWzkZ5Ez60UVH
qfurkTpzRHCSVaXW7K/y0fPZWMoles7LyEfBlN3XIUt0pbn5xOiT84KOPdhUmNq2S0AIYZ0xz/a3
0S63oOQCExavA77vl3cBJfOwlfz+rn0RzpA3gOHe6sL9Na2fceFstP2XIc/v2WOXWMD8EZ3Y46Jv
IayuMOVglSlr87F9annQ2zU+EeMTP/CoDSoGu0i4dOylhpVHNrw64RquG0nzGeQwNMXj6iGf5ZuL
scCuy/tTMpWOl5yjw77MyTs0pIbhJtcpZDnV2sliDd/aMaFmRfAKTg==
`protect end_protected
