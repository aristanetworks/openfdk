--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
A0ArmZy9u3lJK3W5vDloK/bWO32msDjriiYeQbIeAO+z54eJyGKxYRJgmpDfmX45wLZ9/lXK3rXb
U8ZAT+0jQEDWmKxCJSEww0HHPKSEaViXLugaROfNRqNaVcBLWqEf2NScg6XhGw8yyqSShS7s6U94
g6JP8aE1017UdTO/pm5l3O8rIgbhqbKGWaefNS18BW8XYd92K9rC87Khnii66SEs+Vkv0P9H0onm
kJvHThxk6eA1HoYi/hRI3wei8xSJK+Ls5pMEP5Gm3V1pxzSGFXpeNCQfE4e0JbVuMjc9ZBHVkMXm
PibMqOdaWGJppfF3jOJ6KN/ZUzeBcosMmizRPw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="0oD7hWtc5VWg85uqb3toxcKfic83WdJLerQHxIw5qoo="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
OXSUts+ORE++rluiiYsgzBwDbglNP614lxcYL4R0NGkfBT7pakkEaRL2JM8dKLEQEhOr78W6iVvh
NGkDJpByG/NcsPhVMgTIiMQYnZyAjsKcVR68yKh4dY1bM13Fa00wvCd9v/moXjZdw02sUpQ5vHxU
9Ei9ZiDUPI6I/XceynW+dP2liTmwJIdbLueXR70GjReLfD0u1abjrkbZGXi7p/fUazbl4brEQhJC
MR/+9RtqBQxLNY4WX0MaAISgeN8zhc2gERnM61miLGWJ7JUvjidfCcEH8rsHe4HxDtZcUPCCOFR7
6eUtNCRgaawZKP6UqZlUY8gsbT1yImH/uLPsxA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="PkmgGbDxDT6ZXGmPvKqpYMniGy4lGC7Z18FCj6zc4VI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4208)
`protect data_block
YMjsqYN9dcWvIx/G2XK9zYiIGlNN6cnQrrD1oy7imcw2Z2j4UvWC0zsqRmBfkDymO0Wynldc5rwj
GCjM29VKWIBiX5VCC/IoakiedN0Ae3bRWCKAg/okgT4CeDMDtdZtxXEaVbewcX94WD1zGMoUwyU9
ycoUnMguoH085kyOrzlDNV/1TmLj1QaC58aB6/WADsorAs3clh/MJvDl0vuLyEhGIvZHj9Q92lcn
caV+1xHs659Bp5HsBTruemgo2i3AjFk5nv/FbOr76mbMCzE1O8oagNZyVX8IVMO84gDSJ9xfAnx0
jtbP/do/gKBpBf6IM7My8qoPDGa23Lb7JUxzKJO0/IyuRni/SInkaIA/oCiR7EF388RYCd8q+Coj
p+vx6+EgRR8rHCEvpTk01H0vG8RzCLN7jeDsLhUvF5nfFOZ0xzdy8l9vboPlhEaY0A2l5mlMXqAo
2v1q14Um+LPuNo+GnSHde5xLk7P3JJ91gS9FSidIoC6RVXMca2gbYEg38U1tcNgVWujozRlatWLq
+yaiuqUFgnUiMtfSB9VhgSvaVctrieqO48cUsic9VSFijOG/CIeqb4MdPPuXjKGk7DLl+QQSJPy7
27+MhA8MuIj9RrwbbJRXIcUU6TIaUwN6WeFUXdZHxOkKTOQPgQpFvj8wqBMNHTodsQnV8YnYBCcf
iPk7l3WC7f4pmxlh34w6LAgZahKKElg346wi43iIIRAr1elMPcDo3+iN/H9ZCKnjcxqVr3ZFk+9Q
vEKrt1P92g6m7GAOIA1gfXCg+0qLG7P6WyPI/SGcTsfap9s+AtUrH0cJkjVLhsbTuz2wNGdnEeN4
sUjNUcVLEZUo5b5t7erdmIPeziPd36LYOrcqjoI5mwiG+atdPDdnRsScizMFCmcIMTJZX6fQISWj
pMBPnXtBMsQXJ84TAb0/ukGr2XJwiQ+VzmBW/hKVdPtUjakmYFiAqbaCv4JyudlPqMgvec27d0dF
TyFKZWmUQ3dYyGunZJBMMHhsuiCHKbeHllQkKOb6uvhaO3xuEicR1XCV8YxV1eHId0gU1q6XaH2x
5WKg8mMZRjLCjYC0w4oJLO3MIOUk6AAXjTxl3uZ1wZUN2G8t3K3R/2yAdob4nMr7My7b4qHoTbNT
yLaLvbgpLqmxasxCMC3FxC1j2iPRdvE4Nut/1KmpgfNJye8C4gmkVbo41gvlvDXPt+KWyHs4oWeb
yorenjtD+WE1SCUXP4VwwlK1ZkP3yCvSnxHMlO0r6mdB6C+5rcS0pIw2635Lhaqk3rlH3IhYlovU
6lXHzBgDcGbD/G+9UdezRpcqhRDAfCiQILCNFML1NDmCMevPvMVaSHetXOia95RsowGShEJzN1tb
oqFDzXdc9t/of6AigPEKr/HiXKw966rtRCl3B6a2P4o3OM9ugKid+4/fFOTUi3YDZE0fqpnDDaqY
2w8FvVqDJL2O7vaa1Ib4oaAZDT4Ysuriu9jJjXjGHRky5lsqJnHKqVmZ3kptqpNJMOdJFq0PXvbA
f8XNvSSskui+tF7ALiRTh2ERuFQEa3V53fZ51HjEbf3/YHo+sqF1rL8gdZg0QR6OHaR6PBj/rHIM
4upvQtoWF7hcPPkxSOnoxCC5Gwh3sGHTrONPvKrPp4WEzrAn6JyFZWuwtcSN5v1Ga6KZxM2+Ide/
VxKUS5BM3GlQk1w6VVOckSOOnrPxSIZc1E3oiRJEhKbS3Qt2Ng5TOu9jw6smai5xZ35waLlfoXiJ
uJGDFMjEzhBgN7/Lxw5II17tx4JFIvEA4rCv8IDf4Z0f63dUdpHc8o8tRRx6uiE33+p7lhzfglhJ
VxR+Urqr7m2pU/ts8oVHYuru05W++1gMjwnBIGw7x5/k+baDsLIz3BjEGIO0v4dE0XPlXW+wyWy7
O4nct8sbR91pJCt20pZGY7NQcDAESq9Qx0zjV9DWKog3dHYpFdLLDoanDIVpBmyntj8MPOt337B7
9sIN9mWViwEXtt1Emh+arfImDZpI/yegcNYHkmjuWnXj6OwwiGf0YWtFqkxPixOfvKKnFxBcA3+/
Fm759fF3Q8+o2TQnyEfGK2oXpoN5om8xCuwd+TzE0dp6F7pDTcIt+7T0VvBCo52G0OmWDSTUl0Oq
xXvYybR1T3IEO8SRwabqXthHbI1tmkorEY5hb1EZ90aOBSMJHZnuKiKvnuJiie0BnrMj1s1hqwKj
oVoaollikk/ftisJ6cfCCNJamcboWfjGpy5EzG+mTO0xaEKb5JMkfHNnIa5yzBqVpSc5zrkLk2/4
gpiZsfrM2YezfVeRt4KWalWj2gab0o56UR7us7MsedaQxTNQNQFSgpminPWrbv0V+iKUjy3lkS0A
FmqVuXsoQ5dLe0Lh/DPxvLQIbY1MS+HkEHmTA9AYwNwHDH0Toyz6/QMatpltJVkcyecWD3EbHvfI
gqs+cGZTcL7MgGrW/zDtSMxLfsj7pTNoH03ds+t6pzqzx3RhRrfBd0td8azlSMdR3cgLjmDvx9Ct
6nM69KfXfwkmOT0u2irSDD9oN18vJ9/g4SoWaVh2Hl7EIPMpZXy3mwqJ6tL48poLPOtNLHmz/2YY
0sQbDH8xi+yCq1cwtzGnDK7w57UDkMsCIHez9Ne0sRu8vAnhLHY7zBIRKusSyYBKgb477oxUr6VH
Pm7NijZ+5WhVBT72qK9nEUVInMy2dRRQ3WlxxqNKkRWcj1PzuKgVmxAWPYjvOTBCWqW/rrF7cBzX
Al/o9i8AlkGDk2hOnA9+ChIYmK9ZrQuSICjTQfdpWklH1qPqqOJvdEaJI2ysGqijORlZFcKbNG31
TNg5a6l6wJM66982oqJX2RCcmjscC13QIkGzNtbsX/Wxc/audjS9GRiuW9C/I6cLxzjsmohflyCF
W+/UkDB9ETW716p2w6e5xpZIWV+wZZzR/X4pSOaieGZbK5qtgAcnv8XF3GxwPnmMPFuu8b1Ysh6K
UEP7Z+SQjw3VT/p4E8g0BHwahgMeRpJFa3CKOPjjvig1h9NE9VOksulQhJZXmeXx429RhWPk5CpA
pGOCgie3oWLtZXB8ZqouHHfMQfxQQpcvo7lwjUfQ4PVyCjzoC2RqElWhSa1Egwr59jogibMLSc8W
cK1VL/l0IM9uEth8jxz9dH+VKqkq+rCrpMUvrlewRSEnjIZtO45wWmmK5d3ta77wJoZitU2WfURX
gCgVrt739qsmctqCGSMT59MwMtpo0CE/sexaeJEr7Gd3+6wCBtrsGoglIKlxFDY3dtswe9FQZJhx
EXArsCrn4cJxTRyB79FiDle6YhkFwetx9g1Dh5EOlYkO+VWskF+qSMSz2X+eZ63tNXeGCEXeST2l
Ysd8HGVMeSKkBgln7OwiJy/QDdwwE57KTBVmGQsdbw+m48BFInHxDJlCsmW4tHgAYs7cBohNRhQB
APq0EvkKSMxWer77KQzmqND5a9FlyCBvdFRPH/Y4GK3iUtmbXWHImwAPJg2ZgUrzbZ3BmPOGZ4s5
8wrYgl/m1YcOXXkxGxtXmKiZ4LvWdnekPSRZisHDQXJvRZ2n6gN587ojPC7ZpbTjaW+twDNKA+w0
CUclkylIszoi3Vm/lPDz5gAWLoPove2CJTX/b2Tt2XFTkCkIB3nSgZLuVsHDNRL6e2h2V/vMLPy7
R+cxrdR3fm3ZwVXp2RKArW/dwK59/XAFCa7PlKQO0QtC4HsKi208ADDVqUjCrgrPbCdPZRdRXtI9
g+3jy6G04RW1n0qwhcuCjNwbUY/Ff1aoZsu124AReQOlkZvkClP/SE3xueJsNrfgscM13YiAf8oy
+jBzTjknwr6pNeKbagnlKrszHMqhhJ0fKfmfXFmYA8rwog4mreJ0ZdcA5nVP3wqfnI8hbo+ShMMg
CCDgQU75Ky/R5CW8OTkJMxqo8fAndTMyT+rI216YaLkpIOyqXeVlwxvETi5ObmUwa0h1N3bOZyjw
wj475h4hcBxxfGwF/tUbeLkFmZF+GGOyKLukjbY0y9Y3jZ/80duRWM6A9cmxINUqk98rcEvRWeOr
h9KX/pvIkRacwGUjvYOJAZENHMV3WtLZ+DG2ERr4kUNv4xuq97iwTQ2UbaPDNwXwwJObZL+9E+W9
hXkgyScaP+UqRt9IaBu4OUAirsK4g6PscXpuf06znCBrwjwSACsajTlMdsSjwQkxuo5x/7sEBn4a
Ekfz4EOKLGrgRIQVHN06IkRlQXSL8wqsee+BE1kAHBflOHVim7PrCyYP3xGtV5vOLKVfDRnVtdO6
jPexl3KPd39A2xAtTF6SEkNnWzeOK5Xeqg3kKWpd6YMvn58eun4BIczk/2EX0OVxqZLvkqAuTUj9
heyadStWlpbQt51jlmeCH6GSQoHGm+vwwaZS5lxKTUtJ8otHgsESyOzpawb1+EtG9AWT/MRp6c0q
hKvE+y2u1oVG8Gfgj9BNwZcrB+pcXO4ngUpC1Z5phyOwh9og3dOOeQwObVzkxxK96umX3KQIoiU5
iUxoP/oHe0FpPpoX1QuBO3lsJnEOiLKM1HMUzAgrc2utzGr+TMw/1tJcLA2iRtKO5Y+vK9wEItgx
eLHn/T3M768EY3tpYKh59LH02CxDwHaoAccgPAWNZ9bDNZsWBrXUQ3ylo+HbK2Vey0yA3RV+uvJN
w4qzL6G6Y8q59mQyQXh6mmbw6PERhNQHpAOSX0QGSr1ieGM6fMe/238T4w8R06X9z2IZYzOAZKyT
PPUkc4TfDOnTR+lmUfQMT7H5736uSWSQOd0BJ+g8KfbgzU+pWfBjSGaKtOzq7n9sNrf7iGPmrWNj
n9bAEzeLv9dO8MrFjesfsa/wgusbuKEnfw4U929rka1GLGdu8VuLtFuh5CR/At642Fg7PRPk6qPe
g+W+EfwrjlwAXaUtCzfSuxQnkknL1pWMXn1yAOLW/iZkhdUdf3ZjGMz1Ip/t3lCjCJELq99z6+2K
k+1On2yayXW1e5c9Y07CTzNBb5kUKzlBUtpjdrLDCJBct3XjJ+qgqGFFMcUaK5yMV1kykUpfr10G
c2x7DR4p+rYKSJApGpxzV56NH/TdEOLHgFJByMR5Y7U2cfbkIjctplQGYtjLE1kRpAm6G+knI75Z
Kk48rkkFFE9Xql6wWoNIVPe/PEhWrxyNXbie1XKxHhWlKsFOp+sIawkuoQqWKyRHabUTlLDxzLE9
GM+NPLKR3Uwh7d9smELWRYWaFRIbDOhOfXfFfvzJQUEqmTvH/T2OYmeQchyAv1kmm8NtAVCGrqjK
cQLmQfQJg0buAySY4Z8ArViOqpXPR7RncMq8C1Ks9NaeH/GU3B0sGhimi6YNokPxd4IjRipRMiDX
wRRfPpKPeyqNvm43SfAknAhlXhCM/Y9RL8vAFYj5mVND7cMGkgRoYT8R4QXsIbGeSd9hwH8jCP6w
lMsahh6kZXmWqDbfUn/jxHpAzUaWGlG4UBHtOgYDh6zf17wE+8wkRMHZ0Yr61f+fhpokLCrm7RCU
KNpHDzjksmd1VJVTG7s6Wox8oeKuKmFrVNqIyl1phxs/Zf8Cqn6KgyXsvs9HNYFu+uH0UuYrsgvi
yxzMekHmnpHeMCmgzM2mRJuPHMUs6CjtwGQVNeDIEg+LSIuUyhODsGdFFZH6TcE=
`protect end_protected
