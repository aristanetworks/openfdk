--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
QzofFtVNWRNoe7gwZekCRc6LL3ac61dINKxrIOomoguXTkFzjOl0hNF9QO0+vVB6pyGlUo3d0zqw
7yxuWmXCCxvbQnqvq9S5DtzfOmsqaYXJZrw2AT+nZyHADWEhpzvgf2cYbhK4FfpEPlbkYdUO8KuY
eqoGTTWxfLnKJuXbDahYsh4xaVJAhTtDJOOEahrbFk8DpG9UHKLu+TrdToAquaxC/TILK2K0z/2+
QhiiBVnLuinosZnUKfLCsxMgpijdTwVADE5MdToBb0Obl+YAxV3GPChfPhY3kQGO6lA0lGbHaXN8
lHnRxY7IUUQF+hEpGGc3Ot1Q5JmkqHWEsP14iQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="kEmtIaoaidwuBop7p4jQWe4v9zcopg9KTCFYk2rf3jk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
DzXbXiLsBiLI40Qa1UFvRSseyrOwXz8vtVKDhsiEc6TVE8fb9A/dZMAvYf0P7/hyFVaNi/kErvqc
7xT2ZcumpsvU5ojIesvW7l3dVWfg2XdMvbCk7j9raZI3SdhKV2M0kraQ9zoJqMmMcIn8oJ8PS5i1
m2tUNa0R4bplF3tKBUXtgeFv7WdUZIAD7A6jrVp/lGIQcdO2YdGGJtBZeKNo9OnUApWRN1vdwR+8
dC0uEJaNDSIBnhj0/njxToMKJGIXxY6ei+l8k7XeeppAYv4uer7BsX6Z8DW/Fp0gv+1jcJk3iuJA
evWvO972ZXpWfNaIvI7pNpVFISF/FUeImO1lzQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="uOmL8+6zIIef4KSWe+sGA84WMSXv9b7Z61vO8p1JRSg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22816)
`protect data_block
Yz/QrXIuYhlsC/qDfGBL8M+gN9y2niGUhiLpMLJXDAyhk9nNPAP2cPLL0TgDw+jjlYWcX+Tg+yqO
t9sGYEBql2YVP1KyRlrPsq/QMEtO534o4JkuhXOlJgmI2e8TkI2bN8f/3x3ps3ic8OuUosJ052QG
BYPpbPcX3yOOMv+mKnN138R2MPlLaYKILTqjaKTAgDfb01UDyZZTm/FUpx+M762yWKN2yaIP20BB
kc3+HZcn7GOeikGAj78eQNfOlNmQoF4DbC/ZCPoNFqNPdT+kK7BQhczu+lykGZwIS6ixGTNrR2zf
JBS2EmeDYt0Dub+YP5qLIxpRVzQCuFq3lRG+fdwQyy5/QiuBQLpAMExDd4RoaeSkS1ZGeucrZPmj
KL94EGhTwfdQ9YO0WPvhoP++aLW20Tdc1qsY1oJ5RNDsApHbUwgXIC1WlhHtqHlEly18gdyYELjj
0tSZWccmpqE6vzvIVeWpiDKOvmOAsDRiDsS73pbqHScpBilmeXsyd/h/W9dB/9GFL5rulXOL2OCC
fh1EIm6HfGEtzacGGRBZkwpETV5T+5hDBNMVEYZsGdzkgwRHKbn5cqORYXvirM0UBem+DXvzJhJx
0l+ioASDKEV2caVgBtTNpchCRLfZiV4GETSe4IM4tQBvC4tLO33o/w3dJB7DKXFOFa+xFpwHWvNN
/C2uJ2cGPUub8Weldgf7JEUD7w9sXoxBU+eNcLHaMNMpWtYUw4jxRJG8/Cb5kWKm4B7ICacbcZr2
cnrWkig1rJTPkyJw4ESlDna5FxgG3Wl15llxEo1iF7/Q1d5/gHm6W9olQ4QxdL/86Ha/PjJXoe6Y
8qa1BLedfq0UJebwJHwwtq9LChk6X2NSlMYDQI22Vt2Ka5eJqf4ySG/WT2tTA98KU8b0js9p7BMF
ghuxjJoGtBGLpO0EB/t5GA9ZGh80G305tsrHUUuS7vUp1nAFJRqvl7Yhz3AHbx18BWPVn6qXQ8dW
mDyEcni6cQCAp8TF+bRovuFmbPotzpTh25d/lt23RcdJMO8oENYDmrvNI1sgqDjpe7LZD3oQKWyW
rMwsastomC4uNnqzG275T8aiq970AWtjwYdzj0y/dn39GWf6TKlYV+kLgJKyyQ6xxzlrc/Oullbe
AbSvuGtMmIa9biUDGr58lUNi7a/qPvpvSxFxnB7XVaM2X28lGV1aQu3oqVCDcCeIasF8pnfefDKa
cdhetmVTQ6Ioutm34Kfdednaa451AEe3DciTV5w5lwdTA0sgiJ9zS3QbAGG/JTUY7wqEOk+T0R6E
nUbuk+OLQt73SeNXc5gYABzkTCBVnCp6Y9figvslW3L+7oBJm05cxmaBUcO9enQon+Wz8jrTKWIS
5QHrp2szUvGeoGJZtMOKVIc7xXZ60FWq/8wHBilIwpUSYub5ZNKLwffm7Bk9QtDIHHrPdion9cqD
ML/Ng0K8wVWeDjnyz0xMfLkaDuEFbYyYm4uFtXugRfl0dY3FvXVfNSpwVtWz1dCV1Z1F8sQduRJM
xhctRZ6yM5iDvgVn3Tz7lGo3L73G5lgxdUokdvLcq280Pn5NiTy2yzomYfDjkl/mOVSk2luwuo6E
Qd6JTTtJtAztwJZtIo6kZks39P3HeZRLZLhvA1uAvw8jcM/zFR02z+NGXQp90vFk9tv0kz8+cyLa
2cOJjKRwtVEen5QJbId0ao8dKpZ3pU2M9OEb1Cummq370bMsCWLUI9uhoYx1qfffl+dDu1/+Ae9C
ihUiWP8/lR2Iv8BErb63aoWBZ5aR6axuH1kbxhxIhSjn1nnbB6jVKrIWgRC8MKNn0Tdv4jJ3p20b
GMGB6tv6j/ibY+FYpG2zEQ6cJ18/Z8JoOAUq4VJLZRmEe3tk0Z2L8JUzXj7DquUBFnvb/aEP/1wW
jRa7/ZO1k/JFUMsi/4sc2stZcA5byggX5EYDUADaW7CjMQyDT/+651sA08hNhfRHi80QMRSJdsZt
biqQ48qFfyHEHkdCjo3xg2XDQmAEmn5qz9dMcen40OLOdI53Rs1wJf3vGnAvc83FR7EsDvuJoF05
arXIBr2wOVTw2tOShyz1tLGl0z5zlpexBMT1VJtif4pltdh3ENN4Q8kd6YcjuO1E8/5BPLR28e4o
ltCnKfmr4P//8sQXPnlkt/ccxIfHNEh00BFqy8LmI4PETa7fD2PzaNh5wnxemh2a7T1zqE1N3G1c
dGsE7FqtYQYZ/lFl2eoM8hKkHCqyVmtz2MXwI2L6lgSDoXRlGZ5DjbUxDJAopxDD2tB951Xr9eAV
GS8O1JgzCAZqKx4VCFKCHGBfbORGQY5hE3cwyxnliTf31duCJRrG6iteZvlBkKyuqKyRBJLvSlJM
StKNH4EZEUXGjWpPtbhFBwPEMA0x1/dq3kOO6wsvrnaLwuoKrAerzV8CuEBtSgOIqfxKPGYZCcKC
+jtV+WqkSbIsRDyvrhTQvyXjDVRxINgvjCEmim4nKPrfjaiLtYJUcqPNF3/8MGTlQp1HIvlgolss
KqqH6X1S4qVrzo3Ra861v3IxQLzmPK0McQCU7YvDgL3VDIpnrJL4SEC3wFYTtqYh/39rCC2FbYb+
5Yfa9XKHNnT+U5MpsMwez4gKzmW2qaxVLdj4hTQ8seVZgnUUXrjlM79aC3T5ERK4XE97+jjFXJwl
op5goO4eGGmpj4j+a9UFeLzpgHDeMmxL+9BXl4+sNBa/Lc/1nY/+rhrWp8u+XYZYU8tHYpEzSGnO
wus5/po2p4Dtx+2ZN4dcMO2kruBf8UsyhW2DExsP+dQcj9fxhRuD8MNap9SfMkrNjOvYQ5vm4WFd
E3bcwTqJ9KYg8ZEYJawx8KuX200boes5MRyokJjEoXFfIPZwBi9SX4cugTcWMpG85iEb5MroofGm
xwV4nQpYJqCprrNcBjeg1LCU4SnBdij1QXz0Lu10jbqDrWTMZFb99aG/aoKBox4LjSgF8YPBIldn
CaaRZlhODikciUTZqRJq8ivQ0TvzDYKSsqcAspTr8FXfNcTZhogvBxpbeoLsD5e8dCIdeew7b2zw
Y1+kZdTnfZCrVBvabNudG+psC5Wl1ulKkcZu8wH6KWUMsOIzF1cYmQbNa+P1Bzqyv8lZ05Zk/36/
GtF7u7lprpj1cDNNfG3O/g+kOMgS/d8QkOjDCl0gX5Mr8NygudJaI1V1hYCFOqzolJ9xm7li+/nM
5UK3PlTLzzW3gJgccR0FGT+ATmHGO3X8Yac9L/hMWX0fEdYZ4zgqYHL6ZP5sl1kCBh52ei5/oIxu
JTJeHCo6NisG7Y44OpMTxAW4v85ZLwMuLPsn7A0auJ21dUFi+cO228fPlSDl0JTSoU9SX97xNZTK
4BO0LnpfsPV/mT19fO5tFKlYCqRdu+CnZlaZNAca9bmlM10j/rhhVq+nJKCRLVQx9cz79cn5xB17
pejf5UH5fRAi5bV98pow0k60e0a/uUXYzNjX7bFa4lEzQ0qQ/MMC6N85qGUlapVlrNwjvPLUmbQQ
qeSPQIr0nsuxoe6cFjaeOZh+xRqLhEUXdze+ipEXFsHoGAgDVj5jYOZ7ejkKxIw/l9K/AsK/HgpI
yAKrrPQs3S/Hibw5H6Msgzp5bRI6iZ0KY6Jd+WYMbhEVQ8gwi8Fdvz7GiCpZeEwQghFE+J2gLK/r
mHCDHRQzF7i7ICWGOyUa4LA+q+M7LK29CantDJTEyMPznWZAUnfF/IzGPQrcm+FMfyp6Z5U28OlE
pzY3DyGdtR7WQLiA3pb4oB+CiaczqLOqsms4wlrwXafNPAmceEf28kQ2dWRsb5zO65gqnUn7L8zy
M26aCPG53Yw7Hl9V13tndOtah7EDydgySHEAGPNjos/xVCDCubnw2w85xAhh3e9kf0m86sa+Yamw
3FcdiUtXGwf2vNZzZdi0U+UT9XJK7VCRWmOsHHYbnXnvuAd7zVMI5Lw8BO+tqdMIHOHq8n7c4QH5
QNpe15o7VT5TkXNAjxz/kKtjv0iff8vmjeyuCviC3R+awBrGe/ikm47gK3rHGTTal1wfM38RAXTc
vsnFSt3kwBSK70KNzZHcDHKEi5VMBNNEt2+IypD6v/8CQBWkd+IArUgJ1utXwgzWt/oedtv/t5tJ
0xfMFVf39Hr2KjUKrTII46MHUBavRzeD2gdAGaYe7YKwVX0adTgpUfqoI/9aVS60SdVnYMdvPBJR
Eof034hFCxnH9KwK0nBOEbrY5k3RS2eYSSAv++6isHxcrBvYo70GXW7GaqIz9QgGCe2+r7YIN33p
mXvNQSkjV6d++GyYAS563k/q1oSXMdJISasYGP6KuIlYKI/OC+4axuUIkmFfgLnh5MTW3Wv/O5El
kg/1kq7Tj6tCl56vzjHuXEiHAZeUYQus5o9sujgcyglDw7wui/lG3nuG9VA3KFaJnHNSFy/Qr9TR
4xawnImpjofo93Fw6enhAL0mtfW3SVNZSy9IxyTaYmgguuvmQ55dKaUDmsbFC7rJ8uB47Vtysq1R
p3OfMrGCJtPvXnRUsPeWb3RE/Vnp8OMcCuwHCw8hn/xkX/0TBVpbNh4P/2bFY2EiG30cEcgc6AMA
d7alDfaTHpKWhGcEIaJWWmdVFOvcd2wQRSC1zEWvo+cp3X+EiYTdwj+uf08hZDRvwEqtdkv54j7S
X6Sh5bar2+0Bv1ELWwb1F6X1Ucv2dNqxYpIXjvXWZFsA0MyWvp5Oy8JnIhy3v7As2qLaRwOD0rzQ
q4aKNP98Hfn8PfqtPerk0o7MCsLpE+rN6H6r2ZO9GvnvkqzXaqiwHPUiAEwf5/uKUzJK5Ex4V3Bb
EmfuksTzJ4MJFzoLWIWtaEjPCPl+bpG7+hFO6xCa6AuRoGYRwgA5wTQGO0he0zQrrrimBBoyv3qw
NQtH8UiqWhXK0B7rbH+exFgXNP1e7ozYQYh1d8X8lRli3VVqMP/CpD4f3mW9ELmkn/v6drkeBf28
mB2moAitXrxTQxqAshuTbhdGAcK7QGcJevr0gMEw2OB5RKRPP6zkuKAGgCkVpTRVH4E4HCiXom+O
MSvVP8FdHPxy4MRBoS6JTB6qQYzpA5brGsxXPW2BZn1d56JbGwoSSxvLwhqDMe5Nj0Ve84a91TTc
W86xB7A1fAaacgMq2QTVdDfDel8lgKK2ar05qpbJ4BDuhjflGDxlFUZxkQGDJMBki1JeCM2SKIvj
K3EFtXdyoVU6urpf+OzaxALPXypKFjyMGHGB0EqRD+V7yUz/OFpH5DnmccT0atqUJ3rFxQZxLEiN
0HUDetheSm8dc6EVmjkSx3VrHWIsFQIks9eE0yNnfOF1jlSqWBkaH7d2pSYHMp/AeSpSRMAMdKca
jJR4eWUCDTuI0zBRXSAPIs6aC+eiK5Vt6YLviq5BGdNmQZ9dbO2ihVMvofsupp/33ZlWwp6wHEAg
JJo2UoPXvGTOHwyGv+1ckJcsFyUF5RjdTyZ2LX2XyJWaipDR7DZlWKWVwOYSu65NrnDeqpcrtPMA
O5SXRjMvSrXAazPdOVXM2Qx9T2qwhjIAdVKXHeEaVqnAVPNCOkrK8OLli6W093nFFRelhqbR/u/y
v99v6FQLZwR48KWfVcoqxFbujeFiHbT7crtRuhOH3BTWAUqNhmzYJhqJSbhSxHaJuCx+f2tFQar9
n3x3IQKFYfF0zRzN5QSdn2UGa7qtTbWyBcBmzsrsSMftqqI6A1CKFfZMyKiulwwyOZSPmpMFyjFJ
9tqSdK6PLKinXr417L+f77guH0ZupgyAQT73ZSPpaoLmKkMckYeDXcorEAOSfioQd2Q3TYN5YTyH
L/rYWMUlwk+oSRV8JSe+FM406wQ8x3/ls25SrGJw0qvPNb/lw4THzq+gWWW4yqV1Bh/sEF8mH7FK
+KQJovLtk3RPf/jfbhIdlOV5ZiaCdCpr696j9LrA+rILZTWNeRbKDk5WeJfPSLEggzHZR8aN/jo4
aYwzpjXVlYWcgA9iM11ZFzmCJA5N1V0zVe4ozOfyASObTbt4HCR1BzZvg6MfonaW4ja80OnzBHjP
PbjKJ7DSOVKOm8UTJmCvbR9K5A86DQ90usbmLbKvGZH3vVsROaV9fFZN20JwYyAF2OBXnufk0x1g
j5HbWFQb4AZK8foOuhABbkLuJzFPGBgHIl/HGNtlrxxJAbYvbL5vaygWE9Yu303N+FyinrRcgXvJ
5jagCkhVxDK1sn5YgBDYehs6O6Hl4f3HO2nRKyqarc4yHYYX4lngC+FOjp6npqCFlzGHGy8Ef8HJ
RKcWFoMXwrWfcdHdjnRufpgh9Np7ck6yufaEgQOkfZYjVR3CtYZ/0RzFkHW0LD4Ob4Mh5Zi1Dy0K
giL6YaZCYR5Vx2m1cd2/aFtAerMn30JZJm5CVV4SmL+jQ7wW/T71JfCCiJgOVf1ZyXiAfR77POay
bXcIS+Yr3ecs9EldXBAapKVeWcisiJf3DaapmqD+KkmJ5YPlnZD1g81qTk1WlnUMbD27NQN/11u9
cKSyI+2pSMaFgWxmylU0vLCIMpDFda90mH/3/fsjf3wjmR7SEiD3cNbwHW1n3+7IfDwRMOAOczzf
SaBNkZ1XxjAOoiKl7E0A/Ihnj5/xshY/qUSXRyHKg1H+pYxyI/UsZtpTGoPWUbHvIp+PDrIbN8r8
3M1Bdl6mdIYW56RUuYSAEn9MThURV/oR5jh+ONIUxpN4likBbn+usKunMr5k5h38S3bTMC6ple2+
n7GD00s+XR1+48ciGTUF1C7rOM7X372RZ9q0Vu6hQLtn6mtdkvhry6dYDVoSwcLNFHFOv0AqBVNL
mRkbE7aO7OwGrqAhdZgcfIEUZT93dh98LM6xaLcITp4iRBliBpvCQUi1rbH8VA1btmEGvWxUmTKj
leOsayjgQzN4q6NaVXAlTlqNz/MMorFpWOQh+jsBzHu9W5ovr0bvbOTaBfTNNLdsVdlMfTDWduJ/
l2EBBw1DUluRNMxCKiUFuKZCbFM7xL6cTBwHP/oAx/I1asKhzQl30lfSgth29DI+KUS1NtKnwsdP
RflgwTH41Ph8ynFjajXQTlg9WBLoyFjnSTKQsnUGI8VrX60CqpHD4zgPcTLsazsCzVAD3YhguIqJ
Tjt50dZVPEel5g9xh20UmhdXHvmMQ7dJunVrIbRI16aDkeRMUBXuc7B4ivUQa2Cm+srrxgyQaSr+
TvP/HAM+Dhmj0Okmg7mnSxLLZ7KB1QP4vNtTJLjZKqh5flulY9mt06xwDGhp/YScHAFNsuyrxxb1
4uoIgQHu3JaxO4mo6x+rSySH+ptAuyWThAmPBvnmygmbsri38xjxXsF2bi691dj6lYamh3M1S352
byDQE+xWEFJ+Aa3HE1iPM3t1/rKNUXA0kYe7lvsiCgm093WxfC77aHGZumEH4ULz04on+iI032im
hufUmuDwiuXAseA/x0fPWzenNFQyvtCV6r84NKgQv3pxRJyArIpB3vrxjE+k6p2mFV9Es4QVHG03
szPVYkNPR9hE+7oeQQQT3iKlNNWtRD6I8viQMeRHNubb/KqVKpfYBTtuoepce7HCeCf6Iys5jblu
VOFsmYBu5zyXeaciaN7ZHo1Ok4bZGuI31b+wWBWH0SUwcSTVedCyUHPSsdt7E/NuzshLdaD5T/ec
pvUW+18DkhGjJGVXspAUoLs5J4zhW/HJnnnu/gpMMnI/u9RFiZzMF+lqVJwXNqCNzuGEDrKz8sw8
tTPu1Q7BboJJUzUqNBXJDlaXVhiavaK+l/Z9h1AphD5OXbSjpE43sI94xPEwHGhD/kG5nkb5XzVM
HFWnuBka2dm1g2GzjZLRHTvp4K8OxXyntkZSgauxTAkSgzjqi1wFmMuv+luIsMYkv33+o+XI/CEV
uQJyl6gU7lPDzQ90Am9s/zR3LyGOQK/zlDcI2Qlz6gJ9CsgI0CohtMjZtrpLJjB3nfh9AkSOYFw/
CaA5I1Emc7Ul9KIgTy877Mj0LFpPx0tXQ4iAoDSaN2yCGvQcdgkmDbxWMYM0ndOx1RzuEQwgiV6x
zbINxutWR16/tEfZDRyNrTII+b3jJaTUGoSThtZa8AmSTpUmfQ/yTBGJyGgokK0vm0+O9IWxes3l
7VHrltkBhh6Mx178AmjaG04NLyM/CwDma1B59f/BOIMFnaTXNVQt0JdflirfXJuMLgQEAhMpB7Aj
Qrg2p3ibkZwWiXX2KmUi4uEP+8oq9oTAHyEGNjqILdmBnDOT2dLF1dE4RplGc+ibHZkiXpzPp0II
ORRXGsFa+bw9LnH9zLx3/6UOKkK7Fgv/PaWOSxaWQu9B0jU2yezmli5y/R0JdxFZqKB7zqXMq+fK
k4SqHeNN2w84lc3ztHyIW0BLwIb893kaDiNQuqzh8vFRz10tsx1/7cfOfNqqF+l3SpHZwLR4z16u
YrN5Bc3vjgbWHBoSIjNDp7TNIAbwpVMfFzaRsA5jyM/ZOTcj/3USoEGGNuStIP7r8cJLbvRh24Yi
3Qm62H71eNuY0wpOs5OPA2rfgE2e5/SzZ7Kfq7oHb/J7vC4JZ8PhTmx896ngr14GdKMWXlI+X4bP
6wv+lF06XrTWb5joJZTsTM8OFQ8fbT6Ykm7nHfL09POhQ7S+Xdr7lOWE4MIOAv+JPDtxLe8e58LV
SjxyFJVbpsFTIQTJjxHmWGFuj63us0/ualO3hmgou6LCRyHXf1FBwPEUE6UTAg4HBOd6F06LerdI
1au7cVSgTeNRb+caAl+mbMzjdLn0uLAshzAWbGpRuLvhCP2uo3OmqWHGMZUVN9lu7t2/A5T1Af5E
CYxQXaz+osMybhFOHltuml4L10ihl+cYuHcZ0+Nlf149ofQsD+IurCN8cjKXqLWRit7IXQxPw/3v
ILQg6M+5Em0qUIiv9Z9gzsnFhm+1dNbLfgY9PNPKweHZnc5t9FlIyVe/OzqBpO+Qlwjo/YmfazRg
QjIyo/Y5GaffgGvRtvy36AsD5o29H/csxf431vxjn8nujJ5kGY6HO5G6hEJ0+PuZEJcZNdOKXCOF
HVo/a1BL1beW0+oq/5eSY7ibS+YZyhrFXecP5rjvMnQdjQjR6BKbYkwLNbHgwTCavftKe22m/C5+
JAK4F+Dy4cqR5XD6XMMl41XpF6azT1GUWcKV/TgiYdqSl/h6mnpd64Lrc4H/6okJZii7jnUDbyE8
cGTfPMf4SrfnLOUAkbtSckzZZEtJ3tGYzks+FpsKowCMqzOPG+ZNmn1MnbwHDsnGf6qjpZIJAHX+
yAptLQO/9ndtm8hJ+bYfJbhSCWPbgsEzktG0DwxW8M1QmIrLuI+pdB39niL5b5GKkVTKC43KlUcm
bx6Uo+r8e5yPnol8UrDYBnSiTxVkssyIDK7hyr8fYpybV8/YBApvlLKfjPiNBbATL+Gy7YF6YHwW
r03fws6q3E9rFa+vCZ9CSm+Mi70oLff0VU0SEo3Hmod2hNtUFIGKTKhNFXn5dtgnD6tJ2ozZYGFv
/ND96hvQT10HX+h0KqDfyi/bKYj3+CMhjqqnUAemWA5BlXy/WHhGBiseKc9eNlaRLwq7FsxHrpxD
4xWg1LB2rnZLPnLLOVOQ2jPal3OaNcesDHEFugdYu3Rjbts73dYqvPy/fol+S186sr6JNkr3u+y4
gp1HhiXISavvt2uVu+7Q9JLCapYItvJ7T6T/X8YiBeVldtEMmv/fu4qcR6e5EEF4P1ScXwBqULWh
86AKgcyL292j9FLRhWb2LO+CyTrP082cvx5BnI74tZyZN7mxcrSJX9MrOKWbEPQXR8d7tqCxmBt5
cSLXdYVvcIfQ53Xa8cRIf5/jJ5vrR6ux81LuCsnlM4Db0+Z7A//xCcTDVWctNBL2X3g4j5x1keLM
TyclrsEeejfob/mydqKbXaKlhqXVvMpgJMsxPyDr3jcAWRSv/nX1Yv6kxfNSMSPcWhmviRuyZOuk
UtmYmE/2zQw3eOF/an2srMyVkGCoPrJJ0vuyMzzXK+Hqt76zNP3olht4BOv2kmgDGTpSMikZJEyf
lwuWVbrAFJxP40h48nW31Ek+Byq3LijW01PLnoR6OiXTYM/TrR/yTSmOcxkGVF2APdzHKpEqMsBP
eVefOim2kwHyS8NJN2JFOMi/9UFQ+bsjT70v9iahh3NkJ+HwtlWlDdIG0kbUS+SsFeBjDLvMmbbB
iWHL081ayTjp+vpAhC7lU/p8Orv4PU3mun9GlW61U7z3U0271w5/dPZqkGFaU2FWAsTCys87E/6L
zb5l932f+b33wXheEy3QlMud89fFNqZG5xJezih3OfjebB2omwKmsYtKTXJHgRNWc7xJv700UlKx
vh5elY39mDKZk2vSKPC6wFSL6QaP8EB9GzDXHECzaKX/HEk9tS8MtG95rvEqWuz/JVQiVIjhmQPs
ger1E5ah0lalmrcRqf3kmQ8EDod7BPqMj5am6XRqMZ5sIDkxLaHVgh8Uwhz45XCzjTPhNZ04JMER
l176nQMAfGiIl28MAzuccPp1R8DulN10FiFFnxIGzJ5CsslyKXx0lQaqE8XX2tMaCYVXggbaYAVY
nmJsABVuMrL0XQ9esUL4xJLs7KvITtkG5gAj+Tfzphi7ksjYfiucJ7oeeS/MSrnradvIP9FDSi9y
avvNAOaHy/4kHSylSQHriCauj6UEv9s5Sqzrc+XCYI1618BUyeDd4nDVjgb2v8mEmeF6G4u6lNj0
Ttpw+qOQ6SWrKhzPojiql6tpqALa1nEEefG+3kP3Ap8xW1oIHy+ruiPiCZ+MXqVDWOz+xcfAL7eV
q+YjoeAH2Y5U8jiu7PSaG5xraVzy6Rs+QWITw8LOtsw4tHfnoGbzRdkwCp/15EimTj9cxI8zMUQC
gir/BfB6Tp0aRduftdlKOgxPm8eJ9fnDVg4HXWiSosGPIi0Yayt4VOLRXFJceISqRQmzTPhY1wyJ
2rxKd90BEdwv5J4ZLUnRHtFM4M5Usiwy4kh5htr5kHvwRHg8ag5sY9GRqdrqAc5Pvv2qLNQeHbSn
wBKE2hnpnejd5X7HincgWT6099L9j2cy/pxCCch8Hks+THeOMKTuonGCpTX3hK8C2J6ndrxRXYI1
fVuogHwOK3hpkHwaMJe0RY2mHbBICgD7i0/ZLPh2NuH8yM4lWkeITigugUmxfXURFzMy7HGPCb96
C5eJzME1V10YxQZVPGRAE97R4dPMTO1xiTmuxEcndkZ5GxbTg5p6XqAkz5bA6XQqr75rbToi4wbS
cmNHAboUzL2hjBngVbW+GVQlQhONwJbfeNCsy2+TRLFhzPlZypULbiqvgYc6/cIm3lvN/Xn4ZCiA
rIcPh9jo/DrYkGnl99q4PFq49Kgw9a4xhpEDYL+BvNVUCavV8SDyrdIdeBQ8QiYBwAiNX1Hq6rcT
aVc1fDQZyRQThZmH9RRfzGhMYZnqR6ga27orPo8/aRfDZ2oxZEMicwcRRmW25t291SnU/+cOSpfL
lcv5vtmwDFZa+X+hixzK2WWVGN5AeQPRTbL51ca7QHP7NinVEnCZGcin5YAdQ6txGo9tA76M0qoe
AQCTTIUIQAS8EWh4UYQRxHa29/SFZMl3r2KIL6Wr/Fy+ZtR8fDL2MLOlV/gADHLedfC8fnpGrz62
etiUTz5dH871hifjiG0o1jLPdMQbkjKRaits96PTmOhKpvC8HdPo+jxYuTK08EHz/Qstd+koia02
AyiWecd7CO+G0TjNZkdCEOiNg64SoYwNMXQVOSWlrzF7xIG57KH/PJsRNFqTYWqvmYtx4I4b63M6
5BqbxEfNQl6Zmqao2UzEenHzGOfP6LNNFh40fCrzMYbeft7d2Z8ZyLVB6QFvfzWmi5/F7ebBxv3/
c00HzM8DbEZiO87fce64UnWyOEj6EkzyyVuPovnRg+knKaeLE4m4AjRIrQ5tRMd0Orm/OvtsSktS
Lzq9BWncfmn8uv15BIz9klMatsfDoRqF9k4rniVoCF3QuT4/b7duFnuGFKc7VnYpTxj1ZYwktcUN
YMmq8iDoyIl1LoGXcGNZUFZr1FgJqeRj7VrO/gWPVrj9V17e+YUbHSg9KnIVjdw/vbukaA29cqKY
EKQRjZoBU1DLYWM4P+4MMpJN8FSzUHaDUbhzPj4qPKJGOfpaF5ILYfy3BgAqC1GpOiRsbqIwaomq
M62AMhtL1RDrJUBt/GZ/PaTQz+D0G8mcVhdvY9X8TWb6FhKaIpxVCV86xl0A9GtMfXDeP++aKiRF
nQwkxfgjb74OT7/KOZWStrYaQoRLYqzGlecCX1MxUlobu2cq7umhuZei3l17Ii9uuNSqBu3CjgwC
bS0kQkQwkx7gmG8CcUhuP9eM6KlHJ+0EXHThmkXqeJu9cUwbEOAnxeNGFcSbht3zTJuR8gdhwWrj
nfqYhwJ+0YhsXEYhkFVtDPPW6l7UoaSiwRa1mwOJZfh0VTbqmF+cNNX7qe0L6/Dj8mWf+kD4Yw89
EfSoRq0PYXaFYwR2UFOt1kM8jDAn9f7ma2PdrlXPcebaOAchjxiZ2LiixCCBX7t5oPVmaLuLYfoo
ZuaEK4ZG5mD+mWSpHOgeM5T76cKt3/ULkTAysvJtw3lvtfaZSe2c7y5KlyIDRfUzo7ClQSBtQpHk
BKbp8ZZ0L6cq3uB0rRUuM/xe4yyBIGHKJhPwiELEA0bJI3uyF4MnCEEahl7968IXodDqZ5lmIx+M
FMw/jn91eeFrNMrZ32Y3u31dpd5OHZpe+LpDGAnEF4fWNCf+dbhUb+DFY7Ksm0udgqccLVQucp3e
ItYHmA77b+2UjTiU/LzocgyXLVssydgngExFbC2bG9z6rlO989AzSDHaVvMlQhMII458knCuFS3D
VMFLMRpBPrHnIer7600qV4Q/fFpkTSfxV5TpnyTzdPUKnTTCTq/Wh+ZitudClyeowEubYESF9KkB
H/XLBaYc5AencI0c1mXEK0x2YTMWHzaFYhYdkciKYXMhMfQJQrfWJ9YTqSmtpXtxTJ2RC7JsR8eG
Lx3PV55Y5+CRIt/bFNHQrI3Y14CwCgkh4PjF3ADeSqx9APXquvmjqpvYrVtWaolOFyACo29DWsIJ
+KLoIxLwla0CnLQDJfeZi19b1aOrlogaq7vaFSzYU04KQ33Rpc2zOo8PHsVlsPJEAP2Yde0v3aOl
e3nN+pdW7Ymbtoqtc7fpeZp7NH3MjgpC2ft0jI9Ay3WOqZMWDb5hCt7z40hVt4paNrBPGNdYr/yu
G1sKAdrI84vYBxW8AQiCCP5fFB914o1D6tfy7++3JyMw1ubFv61j6LqzyJcgY57tbdECXzmR/PRu
Lf0Ov8BFuMD1N37eCCw3Kcbxn3cVG9nM3cm1UdEvtloEj5isq1ZBzGAZXWjcfJ/dg2962dEsEZTU
loX6i21QpsDvCZo8q8i7DJiCSNEl51BZTELVuCD2xt8kh8YbMer17LhMfzN/372JyjqhGyDtQ6sa
e4q0FgFpXqudOIyMSb7O1/71y2Tl6jFDpCVJvXSfUNAUtAMVuZXanb5hVe4IJqG4Jokhd/LgiiCb
u5avdOYNc4Tzn4P1pthvhelIsbKmFDiNia3O6UvKIx/UPqO3PokGqrddxUs+jMUvLM+wly0OTY86
XSsRV0n74b6XqBh4ZxbSiimiyAxmN1hGaVACZmS9HT8ruICxqMG3WgzjT+iiB+T8JaI1V0Rahyaf
4gtUISlSeKbxarL3Jcv7Aqu4fc/+jZo4EKT/4RCTcLCqPHYq8Mvis6nBtay2E0j0stB0bh0CZoS3
cektD7yVSg1cBvHGcCbB0mzTuggRf/lLNF+WQJYTq0D3fIchmVH7gnv4gp1mbuUcNqi+T696b1bb
XDnd2xMP+1xunUbQ0vOZrXxOj2PjxWuXmvLlLhDMj+9SHZRXQeLweXp83iuwvYnlIRgnBfMLBOsf
gOoO5mYHzgXbJSkYwQ7klR1TBDc5656v2+QPazhEPIzLK5FCx3Jd05YdACqQtOxrwR51l/xPjT61
QSu7I2DR/KQYYmaoUHFrww/Ep6KgE1FG9FmGXtfN7+f39WMR/kjAddgaMOljfToSqYD/n/NqZWtA
l6EU768z/woP1tfML4/XoEeNmpneo6T8CdgD6l8vKNqFHaoc3M9DaWwEj1Ta2/UlNMHqidMIjeAE
5cbBuhtLJdYEFM/tsmxm+R4+5WkLoHtBFTmzbk4CjVEx+Z1hXU4BL3vuQZBa0czlttKmA7JyS1do
6lTKpdm/hpYUDnBm/DygVVC5GZM2xiHfZs1wXArnXFZV6C4lwGfmnTfwqEAp0NTPKL/OSjQRNwGv
ErIiH4RA2i5PcFNQPTEZapnSROIXctPZjVmA9RxwShvNMAyJ4cvBwfuIGqDYEYIAbbgGkCKJ5SQl
CeZTAr1V7DylhBa5cdZCVJTHP3IfMJITFCirMryMJSz7NP3DJ4S1zywI2xnFtrh3Mz86Q9jeQZ6Y
hSGd11DtsNkgzkto6n5pTRdPMVkwGJgV1NjJiqPtan6xoTKy+Y7QcT4yJ+IIquG40EsmRLcKGzPt
f9OWw1TSTSAq18KjbWA6HcNHO0mpw+fZBZBkpmcZZmagD8aGJdVeK5hd5UjXqQaRoa3P5psUrZTz
0Os/80YjmgpTXNSwjLmC8MV9w2Bh3z4XG+2x4HmDD2hOhHriuqdXFMjZEo8Hmt76qQZ2oo7KbXG5
yw4xRvjTUtD+8cH8KvRNtAviCP4PKaaK8kLFJkH1U9S4qOLtUsC6sCldWZ8jwxUhTqUxXcRSU9r0
1HXBIudRZL+liPpTHJ7f55lryxOC7AYqDi1G6YTkEfy0HnxvzlMj5qYZ0zmnYu6+7lVVUc5fCjSZ
0hCTjw1gdbxETud1zZNsct1qKBrQso89ig17PB/lXJZ3Scgq01p+qxoJoSgwPMO8lu1oUsa4+AQL
HoRfdfkyKfH+idhAekz5771u7JgPz01vJuMD6z8HbRiu0eaMSsc656zmM7yuvV8ba9ChWGqcyOkZ
vRYCtPH840+y4cy//HrKFVte/Hh7xRSNVqO0MHbTermzDr96WTqlyUX5TEzefEcqpu8mvwABmIun
1/ayE0yMe585gY166ggiBEnM9UKhYCmQPRaB2q22hkdPJzYhlHp85v6PY1i88D942yi1aNa01Wjx
bgs6J3FPCU8qaXwklssvl3HRvYVEPES1ZZzPbSOxUsoqWvvfUKNdZ6K1GjffzcW3juex+86kCPGN
CpgOKWVSxSpBM+dvB91+dBGDZ9BHwXrfVLsvRQQEdfCCqG5Op376ox53p7AQfgCipjnLun5y0Sb+
Rhb1fV2yZCMINjESb6oBwlHYkSns6v7onPo09I/KKeZV50Ac6yrJnVEckUhqIWA1GNMNer6uE6EM
Ns3nKwuDGc5pJ5wJC/ml4JbwiDygeBB3GvSUcKfSKscgviOb0SMBz9RMJU5FcUOIF9D784kKRsWI
DQKR8i+fsODgPzLfhrPCEJ6SGsI+leopOF4U0zNFocybegxh2eJXmgcrMf6+ifnW+vk5tgXLAh2/
cJ6HVJ6MKcKhZGHrtHNOitApDjU/4HF9vVEpR8BUNuBxgLAzwcsI7yuPZrW33IXSfBYORdM6X5OU
mqXVeEafQZpdrNyyKaX3D+AAQt1+PnYYjtkTSuYKeiaNNXBMOt6z8lpt4LnnGe8+jWS4BTW93M4c
GoiWMNlrOfD0aPrTTLyHHcR5uKWPGYYDpCLpRzjYcCPWPo2h9aig/xsMrok4kTChvaZqkZxn/VTu
E6Nk57WdPUSH73RZJK6OTaHVEWAl7goIUNMb9p2v9kLyRMoqISUCKlrF8efCd7grkbYq3mWBk6OD
pAabZ7RUC7PFpMSABDAsHxg7T/gMhd/Xgw6tdN5jKBFABon/swV/fihC6DHOJdwuzIKFUKfvNijP
6oO1KL2IXMKtfQa/NnpR/F5YaibfVYPIPvQ23OwWKo387r8ninZeSGsQWNQXvD/tIInnUfpfXS+7
C6O30Z/7KUhsd3samvmUVQ+OSIdfrkCXowSiSNwNkCU3Vpx/tYXIRzUHvEyqIOq3cesKU4+5VBMH
x9jrloaldfYcHqagmWCworInscUFGoI2XZtqD1wEtzPcd1SNkH9L831fqIdGj5uIqFblmYXgT+Vd
3NyV7te+iNJ7aFBt3JDWbrFiu+WIlaRetlY438vHy2LaF/XZwHCSqjJCcNrYXI0yGvCZmqrTE7KV
hPXA3pm5lq8JjQniWIQi4cTRBgiAH1in7noApvqXitc9kU4L8XpmFkOXOpuphrAi3WRfkf5kQiha
3S1z4M1aAxdax8rLetTkJhbdDi+OZGsYrQiTOzHNbd/jTii02pbrlESPmlMcyw5uV1DMUPX0uL43
lH6fNUxPYVTVeZhcskUrf0Orwjz6qBYtocQL6sEkx+v+e/RJ5NDGbwBOdzoDhXO4mT944J2Zvksj
X80i31bYavLsSz6qsHrmO3wwWRVGkSIBudfwpkAekN8YQrgevxvgjus7q4Gn8z1AuCP21GJ8F/zb
ETynn1CGZV9KaeWeOKiMeqXzy8ajSk1NLVPZ52VTJdJZ3CW/Rq+N5BVGGZuLuLbfCWwUVo/+BxgR
D/S5+Bg+BaQTwV49gO7NF4VNtMAmHUhq3bs1XMZAOBLFa8YAYZ4vNFtYmHKWmw7MlfGGre2ULhpk
JChyMC4d86/vrVZSM8HwpJJ/2WsO9UnNs6M8nCdFAaLWW7a93RNqUnYJ2RG8nnLdM1j3a2zA+jS6
NBtvuvqXdH4H0UEboMK9hiupwxBrCpoYJGCCwWcMNNd4VgktWAxLCGh5sV8IdzuHSmKc53U8ZjEH
a4sOvfvvVK5UT0UQ+Vh6hLS+k0V2huw7pvdEsTERrzFaJBeqXYtSm8GapVMCaaFgVzuyM4IYk6SG
Z5vK0LHdUoy/2FP7qlNl5sc1SVMf06hGNKR04fBVeq9zvB1Fv3ZD5MqTawG8OvQ1i3EQczjzuQAr
M5TABSuYplN7FfLK0ihyR3kMdThLHVvfI8oKWfEmpshRVYEtRE2KCUzWg8N+wCuEuvhmNhCuU+Cl
w38tijbNb3/XOYnVFSa/ZjQh25RgecYmlliRYM+IMEEuilR4C99p7d/ffPPD+yvqiiOPfrCp4apc
y7LP0RuIR7pKal5yUBCl3mlethcEqc/lorstJ+Yo1v9ccdMDkopkZK4m51MfkOnwc1RC0R+1hljL
oC86yV/Rtbmn6VkqjFP36ztXY6Y48hxsjkicc6z48KAKieNklX0G7ElA4mLk/NA8Bi0lsfxG5LOz
RaZzNrXij18j29JNehxLOWn53TkatKT0iSR6pKHjIm8w/NohwcPryMay9YvsbXRkuJQNTMpgcW5e
KDcj/oai7gNmLkBsAPnR1CfLpWPKIkCgXRsikzi9jlKJdN7SCoSY9kfzkK4FqQXS+d1PV4AJCkyP
FJmBNmoPHJdzlJ5eayeBTjlSArajtzuPTlP0O9u/NemCmbe8CQsldaVZI0je16f4CJCihGv5vB6r
j8TaLX/uBjMfBGEUSB0/LWi9sfDyUGcTp/93SY2SJWuMjJ4E6lXY1sil0zjtlT5nEng1BNFI6ldU
bS+8sfVhcboMkILb2BesF3NBm1IvLa6xWFn6NTh3K0DsqKJYxQuaJPov1fCSEsHSSJ/fXeF7ZCT5
0HioOvz/s5zlD3q2WY04V2AgB71wYXDDdofQ7o2txIb8M2I0skA/Ln0dslTMhLD9dumhfPthFgQP
rFFUTOgwHsygoRv2Qa9h/ZFF16SXW1SVOgP1rLbPlK84aBxEVMXb55mdoLlOhIQLcGZw7FYPoCbh
QRpJzF7lR+V1tlGvwPq8m4nF6lyJSeJwc1IDEqtT+9jevXmCRQqCrHN4K+Zm0Mi72Kb9Xo6TY3va
NTWto0GlKCaF0NBi8YDs4ywe+VvxIYVdMb/L/C9MBUTbZ8Tec2N65MvSXh+nA1s3U3LZ44baRl9Z
r4Sp74h8oxxbUqpEfbTjVPYfeflZsRyYrYObqjf0WJiWh8jFZcXYggn1Z7+p9gJYZDnCm1yckyVU
IBVkk0hrAcdjNjROZ7cCZIJJrKrvFsjHNoxenhRUVAJhQ0isEufMHiNoW/rAl7ccR7Agnm7eXG7R
bbSkQJuTGsBC9y1vJytPkoHsQMHcBVzQOmb1iKfvDSfTYoZahj/yfahz6wYOG5m8D5N2NRoD33sG
qZiYsCb8CQadVQ2wR8hCk1pURba+vX6/K+FIkwFiRKCJOh4wzgMZWVj20RVmuJ5LwX3Yfm1NmDsA
qSqWo5Nc6aOs983UL3hvUwNaudwgCXH2LHM7kdZTAAY7yQSlfZFPWN7ijJefV+ucZYGMgnMrGv6w
yHF9LPXNUTmc7H7ROqRJvYe7pXqS2DNxd7HsSOawg12WFPIvPzBPPl4kd1w08N9kNJuQhn/NP8oL
R1rUDB0c0NeEDGcP3Ze9VCYdfFiCaCL2GDbmb5a74Z/bDVJgXmfPLLmerr/dy9FhCKOjQPDnQm/B
SmRZDMncBN/KKHOieakoEAuiD1x8n71Fr76CSvxhOgHznFwVFCHWweo0Njgt3gGwladuOCCfyZLS
hCl2Icr/jqEc3BS22k3T5Zf1oP9rqLM8LCNG5aG452TddNRMYp8FoZib9MryMbAJBFV6Za5j0opS
fkVinhgFRBsnExkSSQQsnfNmMGXnY1hiR7Iv9gqAORyPAdY7Qm3Gy/w8iIDQKj0EF64K7KSMQu6B
a8r1kExKpqr59vKSYk+y0L09cvGzW+9KZ0vUDnKCLx/lG2g2ebewMVXwsKweAbSwJNkAI3FEVLeq
mT/NN7R7MsQDkQ0dYLU8dXWbgm6yU7IXhvFSA25ghOtq4tAYltxTfMsxYA9yyrFG6Z2sUOXl+xPe
XPlosgoAIqQ6ju3fc4XYQyJTNlhYsmdCSMv7OEqES5hl4E+xsLGt8YzQIsqG8xvd3lHzmDUpQPEH
32sy7+7lXn1UYODJYavUp2tIYJFVQlo+yciZs6tvz6XhjxNZVBtUp5RY5hpq+0v1uJpExxaZ6WFS
xDdSGBX96OR3Fc0TLH6m2jZlpq3JEKPIuG64j8l4URtKxSSGahXSo04gm/feTdwHfpXQPubKd6au
8YXTAeoEp1cOjCRT6FTzWD/dcUNdlXEY7yaR/dMGIRV6jwi9CGDokv7lzZoro3yzYo8KKufiTZVz
nRI7PBDgc+R7UE/ho37jpYeys0y86MmnKZm5Fj3P++rRSE4iYiFqnajeLALjlSA4j8tbQQwWqxAr
2jbxSAbifp9b8ttXR5DKExADmzILsAAG69WR32+QTYeOf2MdCL/uCa8XWrfYTHyNuZfHGIvh1hKx
UP3eG9Uwjc1ONOyu5Yqa0AURvBIpHukocKzLAdUCPuR11hn/zGkb8vUBCn/q/TB2fG13WUwh9fGA
IeuKGNWUGORTrYQ01xA3Dolrz5ztHpGpR9Yho00ovDm3uL7TaVvIUqsDRLnJdiLJ8hjH671h4eQq
voNmXvcdCDsmuflP71DsKU/yD1b9FUNo1QJSeaZS0nZ4+PUYLq3uDvGLdPtkGBZRCJ0WHB2599KV
PJMLu1DBlhTDGMxl8ZJdPcqluk1bMReoVEkyHEVzrYAOJNA/psN20rayCir29PInRYnoOioI4+fg
sj5AoWSQQQN9W+7c34rIyWV/pPwP9EbqJ3qGTD9CY3tjRaIM34Up/rKkycPK8n0B4F4vkvobDx8/
D31mRnwUGPwllS2ze/Eu+qvbDsw39dhpegADZu+QG5Y5rczbJKfow7/KdriAjKUHSV5V3EKdXi6M
e6vhHj0sCaErdpNg0Zel034c/cbSXhqZcwUazA9cbGEYOQ8ojjjrhVySnPJIM3bFSNxUjON8SQCc
03zQ+HYGmpxIuXj4vh4K9ylwaxwThnp78h+VcFKdwZvGfyftCC/Iu3YRi+H1HSglQxocDS0ugHiP
Pa3qvxrQiP6WzVjiUI1ZH9ZXl722Y7mC080/Tpsr7w5gXvh261Rxre2BVnIVdEXR5XhvmT8Uzs8Z
lkEm2xMD0WjT7vNspUg/FLRzpVBER6FhjX1+Jee5zyhsyyce08Rve4ljSS/ZDZ3qnXkftnvMYwA6
lvJdiHefXUY5wOAAgxwXX6G20nRSkvmhKChVAUZdDIU1vT9Rl8C5bNZgZDeLQpBFExj4OnyPHoXd
FGzzknp+i1vbxYu63xwO0A9P+5E51BCxseca6Zk1zTfVP6Lr8tJCcjU6rWLFujF9BGSELRC+9zEq
9wr8anOPUFlx8/06e5TWHZKgUmJ6XokLzKBX4mjWXb2y9Pg2E88Wpft4nLka4oVOJiBvPPcrGiKv
J8Su7tuvP+Ky/x5pDYZgXqEHVgNMQs0Hh++ipjD9bTeM6/vMCM4IERLB9mUnmBat0DANr1p/nweN
Bh04+mHTCcZ68sZ9Vb6PB9RviJC1qv7QISLezrYy814p3CXL1zJTK/w2qOE+C1mOEJRsz1I/GmEc
MKNXqy5vSaXKljPBstazOYuM5Uw7ahTy2xD/2Vq+QGfT2mifQVwnwe/FlqP+Rm+NDYZQavZ0skqG
OSRMK3QvCwis0Zrnr5EoYfZsJmtw8ffFyZ4w+BJ55o5R0htglWFqSXNdG2+mP2H4vLDazegPvZ78
6CNZIWHq8Z5Jzy8Ti9+b9jjAu52ItZocg4/jBF4Mh78k7vcthamHoZef2O/+FzR6Ah302KOLlnxd
OJT6t+KrbJzQyQqS6wGGh6DUNbJxR57Wsf3DBMkklf1NltP8imYiwuAbGyd6aMIfALmwdBvqrc6n
mrkB2hqVYjCVpIJXldKUuT5ocGLiDuDC6Grq1Kwaqv1LSJYmey1BYU/U1Te7up8zM9/QiEcJ5kM4
2dto8SoYUW5FxMtnAymzVtymTgWBv9MdkE40gqGtKTw+pvuRNxIs4UNPBPW13kaw8XT1JBDQykUw
AbGlMNL+izt0sUEFoBHN67kp/dwK3cb5defuSIEYUvd2OQABD0pCGcV03TQWFMh777xO7X7j/HiZ
RCIKTwyOTmx/BBUBb6G32FX0BujKtiyUk94ctt/g31YjqT/VTQg2cBHeJ+Pv5ypa0prynLmcta3z
t+c6q3IQxFXaG9fwg5NTqDgQ94Dm+Vi7D6tt9YlTw5jSmi0Qnzne3ywYuCo3smMx5FzJVZQvLjHe
heTf9TITwZKSSFqHbboKST0zQjV5O2MgBqXf+zYhslOkUoH/wGj3QEpA9uAOI59/LBsFXCgZUTeU
vW3WBEHRt09H2HZC6ZFRZF2v8xanVbnaFFOh8RbFyeNAeUSJwVs1tZzJ1ELD4XdQUeAqpZpfyy2n
OjgtCCLz0TDz7SZcSkHSt7AdQ7u5kenwA2YAra1aDKN1vHfJwK0k8whH4ZxSbJBDsDQxHJbVF5jY
QQs9TZg6qkKm3aS2i7FJ1t9eVCqjwZttRGuDufaWxoDVKzWBQDUhmBxTyzOBJIaqTE2kob1FlRvT
ZjF3+jJY1ZN0ms+iyQ43S6AEqjam38ugy93tI1Nnr1dOPzPJv/N6/fZOIrPf0RWtEnmUdmi5fgNX
T6vT8o6cbOGHZ0kUm9BdPU3HjAv+YgR5ey/ajvuycKljtVSuWub6kM3crP9wCIrgBgH5Uu30wQsj
RjQ+IZfWKvVrksN1IzeUGE5/EeXUgLOXio/REg3sz+EjGHZDKO9ga3CK0X3zVr0E5rxT5wppaobF
jPab2zn3lAbCqEkTaU0aV7rb5FniBf1a2di/S3vf/zf76o2v22/HBCEkUS7FJLAHbJAgJ+NvNnG8
xMR+hygXT9yBPnpO3IWf4E5WESVQ50k6oxHuJ3nRqiqV48zNogJ3f7dcVFzx0gZ/jftpuC8TfeXE
VbO/hCw31QaXQDgZNiJf+x5xfQD1oDu3pluDgId8lMFk/Kclr21uAvcQdlFpckmMP9CRmqXxPUQq
qLIKZa5DwxSFGKmDCel3M9dwRMrhETMjQGn7jkkaEtuVYpmQyutjb3LqLiC3Ph/EfYqEitVMOx2N
QGRaXKsvS+Ftu4R9hEvT1SDDEOrD5pkqs2sJVKPLbie/FpSLuQTOERMzEwlB/VmS8iq9/kYQYIAG
JO/LwmddIaYHPUngFipdwUWU7Ug5Waw5D/MGqgsTZp2isfuhgQBrDYlNKsWnO8+QPeX3l+k9pG86
jwTVXrARfYzet978rQavuWbdwiftHMfcUXCS0OwgiIVU+8bdTmzH7ez1JTVBKuXS/rn/cJM2LO5G
LJknfvDOU5ySaMzv/w0oHVuFzCuWS0s1Yz1IFCNmKp3r4ABPVoxUMgYHqQoPs9YTL4XO3L4RTy5Z
E5c6M8481dqXWfgddqI27YsQv7rQpY+qCtGGHzz5M8clpfrbedj53LqQI6aPdibInEq6d+IE28uO
V+zBiBqjh9xaE+M9DjuGt7IO8/vFAwF93TMcEeeylpC29gKryEIZAiSgNiCHg5jQkBc0+BvqOshZ
ySYbz5MfWzuFfq08qZJFEW60FL5CtfHTyrd83Oq2tbkIHzWAQcWHPEsyA4H4LkmfyI3sDDnWju80
NWEzsKc0n4tOFMOAlJjl5ULNUkfCpfW3xABKYUTFtPvjmM+1swfKXJCNJINrVsS/5C136yl0L7ue
xi73BD/ZJwODUCRLEhMg7QGRVoxxqheopO66sRdfO8gcekHMeJRLU+4XZ6CDrXbbih/45y/sBRxl
nojgrfVmWnSTUJjoHe3YNlqqjB19KoAwa16dPSjh273sgVSJRxxPmNIKFm25rX4twXYzTMzmSCtN
SkHIvLNDWmrD6JjNKnsRQmWTmevDVg2TjDl4vJe/UJrV+tGejMlZuvhp5WDQ31dfea8tdmTGlE19
ssUwTNiPkkGyK6F6F9ZdA3JpiRmGGDs7jBEjKCLMsYxOl/9k11FextFuA1Iy5hxx1PhkHzgz2Nwg
lRL5Qyc8V3Lp0NRgwxvFQ6PTPEWkA2eLd8WNBrPFDPn64P4fjnJJpRA5/NHZaMHn0HSI6b4iGkJL
zm0hqzxtKR6IhoCG2Lr1768677NA9sjWsK6nbFDviHQ0BvztsA9UfUITMNgTMkolJGQOFqhjimvg
LQyE8RIUzG+8How49YM7/FoIIH5IK03qPJXr7+bLNne50fDDwqMMNux/ygvpaL547mEkUrMCPVYv
LuXGq4vW299PmeZ4Y6W1zMpB5MILDaAChpkXBq1iczzJcai1go8FDrLSe4GDAeuO+q4J1tS14Izi
u02a2uPPW8h43jiqwiPkxJ+lG6Gqmt3uYlCiBo2iPnOtyIXooun4WviWlsChJFKzEEfaooX86DS+
cystVP4GHgy/MJb3u3vuG7SSpBqFJg4BmPbIuRGMEg94urFYubs3xuTUU6QdKndvIEHtysUcmn9a
4nYJJpi1RyqILXav4HttzTXdLuVP1Tid7w1dmjT0/C/G3SF0iszCAO/5I0HyiGZQcwmo2r46mU4Z
EIf+Pl5ejT0JB0Wm9QSmydcCHwFLhCBOqz6MaivchMVRo5OirbOVtWBnImN4hBLowoazXGWIkNf8
MnSkBBjzNn0sCz0Z+44eofhjJzFBHz5qYlu3mRufF4busrOgCGcNUH/0ccx3WMRR7vZeZIIa2NRY
751i2ZcPhSeMVqoFQ5r1g3OLyXY/7oh0X6NZ0onOiU1t9sr/OJa4G1iVZfGeiNnJHsmVQnlOr+WT
6uQkfOu3Pw58gxg8xj9dkSfV1hZ/gYEuIZUnIY+JkibL9MuX/8rnoMydE3hwSMlq8Cm0ip3hi+0j
V9XdcKT0ScGZ9bvccyKxdfBP2X3cjLqLsl9aH974VW2YnVFoowfsG/VlTzst+efEK+SrVza3rgri
4v7GAaWgW++CzX737S+vWi15PIMR+TGjVr4B7fjpjHqDzEmDVHx5fCbp0sDQhzxPDaVJGmy6vFon
lQJ78/newcZyTyhTgTt6jkvZzrNSMmByfVeV6c1mx4VwRudGpyZOeVtCEWcZTVS5ko1lznaFbVmw
nHYscL9GWkMmJKMXjsfKemfvcPVoRDQX9QHwyzN+5Cw//Q8sGjgkZ87sKmWTfj2SuOokniqB038U
+3HrjVMRp69cIY8MKWPOR3w5AB28g7UAzZoC1DPkWmkshJITSu88/muhqlwJlyYpRZtS0NiDpM5g
nBikaGVeMSEgEOBTUQViqQCWoNAhTchoVElCNFt6w/3knHbg/LYl/acc4HIi4UuUPXCyRbNmnr4x
FX9KH8jSfM5w45zVxqwFIpKzBAK8dFCJB3WyFHuYp86dPFpY8CB2a/4xW4598RzNwsmqHd3YpFp4
zcDEiMWTu3sDobCBQiVDsLiBKBA0/tp5iCtQvX5e96mWtuVC+ixMUF9s8IX9R7wZnOr6lgwynyEX
ykDXiCkY6eVFCRRuLKchIw9W/y4l6pJozxOW7EZsqijMq26P4SFKj5TRaIxS4VBSTyoee7ZIKqOv
Iz79ipW14PQeZrifBdRP51Pj0U6V1GgVDcSPqdoXgZgBxL8RHD7Aqd+0Vn76PGFE/Xd399qXrCWj
oBtR6C9joNicb4rfFa5x6ncQogdelbtOQfxdDKyo8i8Nq5oY5B+MvFP3PbnRzuZKCoEu6JQEKb/l
tHqcz97l0jWYJqxMXot6997PMbgMKOYpP/TgN5N2iWAW2KTIOaGtl9d8h8dtxccuRC8HAFGqXqxh
145DeOfwolQY8zx0E680j6suBKokY1NT9SMAr6XoQybyqv78XOj3fQQXsbxsM1aYCOvfI1yhB+OF
f3k/iUzO/SMiFnv8BPQwpiLJ8I7ejnUp2vXQb3T1cEVq0UaleVjcg/tRT2HQ4SaQpf7s5ZbBRGCj
wBAiMYB2XX/cbkCLSRfOyj2QhHkm2mOhZNgfcc44jaeoHBtY776qusmCwftFLVYVKETjznsm1W/6
zO/I5rwtqRnR6CintqTRg0SNF3cyT2yZzA0qYMulX3vAvU/9LSsi1et+29QIgCRkpOsnRYfD6LNj
iSgOtnoMIXiP/r6Kggt1RIpqukKiXCHQMyY9bXyIXzpRWpDL8DnKwaPDVAxd3FiIobs/g55A6o4J
I8f7hGsppiCihPgjCvvogHjWEBSG8zhVwmrlZQ+UzC2TabVW9B1k9KmWJyhI1kcp1FTnjtAQ9Pcb
dPhuUESGoR+dd4yEI+cUMvusfjB5Q8hbwJoil08xae1SqOIjUNRbqZ1b+FIsmKRM14lVdrKWir+S
YsX6GU1i3c9nfD9skw7bk1iYQXrxDFlphywfBxzLyIujSQQJUbYwLbLcyUwZOXT9uO7kQze0+Nc6
6u47FQK+8NpZXRWK0ZZISw4YZ870SlijXSoFbAGreSCm8c+scuThtDbffewyND9VQkrkNWl+sWRQ
ZsLvWtQIe3ANEByp0CXLm6WRMqHOzT6trGF9tSZrmj8GYAat5ib6jpV3VuxIINmjP4Msv+uH23sY
crDoOp/2/NilDFfBPokrJZ3qTjUVYckjQP3STeGwy90yZ5qfmFTC8JVqjJiJaWcBpoQ3+2By8D1M
Pg2aUFZSwnmRKcEiK8MtXDGJ1l7jULy/x5A0uUSu7wiXz3cog1KDN9YBBmtXQEax+a8VTKf562zb
/gmKBkRnC/nWYLq0blsiikKHRRl45CqH9YVXP+EDdv3dgJU+PUNdK3PQe0Zs67B/61YCK1LlQlLW
7TZhQPLLzs5flvGwAwuZCyXZeYvW3GcGy6cKdq57mSI0hFMu4NFCUkomVb9EpPaOhJsa8nM+BNYu
30ITTItPn52ue7rEr8n1EmM4+8vX6gTh5zM1uR4nq8IjYxYnPAkQaS2UREHtWgAfSJLbnsgxBsh4
8nswy9zFHVUgbYOtUNwULBe1CoJpnDQPuorPKtfyH60CNVxCpYBqSt0Uipt/RsbtQqPjYOYwgWKE
FwT0CZ86ygLIQtyA3OneXMDzzD+jN8x80IIKrcALONBmJ6DXJgrs5QAE8GfFUuqyDs2EPf8Suf8c
o44kNzSliH3aDuUgrhNF2GZ7PndeeScl8jZVGdJO0xwiluqLqlvSD/sab+KvCqedfDm+Ttj4Cu9+
5ER/FrXinkAWt0znOTnjruGpH5o9RLL29oB222X0At153ChJFhzBJkigRNz2vvKzy06qH5iGGbeP
tEWuOiXhNFR92KiqAy9+67FgKn7H/Y6E791oMC1SeFh4mmWSqwL9j7KtfFY35BBqNYwhuK0MP39t
BCURh6xzQgUX3oMx/J92A9/AHwJxJF3tSCEVg8Q4pY2AMxxvRTEbn2UP6GRj2mg8zlrT3r9c819Z
m2rVdTNSOEI8NrSxwe+Nii4sSD6rjgI/Xb7M1m+zrT3wzAk0xC13GpJzZZBajhGPonGKWhF3DEVf
FmxxX/ilI0VoZqviYX+LT7nCMhL+zJGSs1agW+TR4JADzmdI+wnUCek2mashKSxgmSjkgRzbrvlF
n685VwiW6cZ41FUgMuwbpFWyHJBUwpuqwSdmFsWTykNNjg/G6ACDxwBYbNslFzXcNw4yIWfD/GVI
l9JbL/Ob8xJ/Nh5P7hn9BK9liyj175PDL9yRYLl97MK6VAl7GBlllh2PpeZMORZ2dqiApMznB3bj
eu2uux9DGjIHYwkKAZSyMb2YM8ycm/NeZQSvRjHllutz7br5DmQxTPgNADfkpUWQGID0LKAc2XR0
ydhSRQWmldHS0RrJwm+/RoSBtjApJ3A/ljiH0bCrNAXc+ua361fqxXbJ+NA4kPsiOaX2iGhf2/u/
syGUCf4u7Iyu9t8v1jspchgzR7hgs1B1YYicV/32F2dc1MvZ+LzICPy/nLKpvRUWCE7MmqJ2VlbG
9Oqw/u6uou8thDLdA7SYv3Zq6SEYfKgy1AoJEAAuoSsCfIcsgvUfHdXSj3r1IBgNumG3GqzpaQuy
cb6cuL6UC9rySK5zKvPCsVTbjPS9jmqRioys2A5rd/XFZrT6qeHOPcgTD6tA3T6A06oW98Kh7b0G
Mk58Ai4ZaSDSVMguLMWVDNlH3e+XilhQaz35a2PBs+8LoIppzIGft2S3FoLUCw1r9if+pJrl0Su3
dQEUg9fPybQ3gbSPDNEnuDT/+iqnCQ9yIi5Ea9AIU4bMyi6uNCeWxvMFzMqkXPFxiHHA62B2mtmU
evTRuHM4NEvIDZ7Zo4+2CdFLA/cPux3BDwhy/1CPqZWAll5Br5LABCfFm8/Ef7KeMIjOQC5kKQUi
uDZ9N/G/k2QvEQL6n5so17j6mHLEDAq89UqFNW9s9iqxSVUuYNkNh6O/6BPBqe4ZMfS22/LJEBGN
c5Lmc9W0p3DPmcxIKs6xpWLoWosJUr1I7XkTLwRkYkFMWt7yQMNoLDlsY6S/nQiH5lRwJFKEPmLb
Br/BZtZ0aDunGYiZG3cob08MvJ+fXcnuEkSIuZtDkLJY4Uo0mWDcERzhe9ZXL9TzuNOc9v5I2bGU
yBgvwsmU4SOVCnTjV598ogDuFKotGGkbK6qWOWUYW2yjn+ytD4fCHrbrDfGBuDMh0OK/VfCK4QeN
Od+aZubas6JOy2Knkize5Cdx7BlSPSMfXvWuMRkefqSb9jm90yMYrmiyY5Rd0rLJytGjCZhzZhPy
6h/8sCgzNuuK4vdPWAaLMtt+CmVXbIb2QtD75/ZZh991VwPHq5G7l4D/LBjZ9O7MPBqQMOzVRaix
e5yWyzxYLXrvJVGYqNuvsEl2eyC7YBVRQMu4vacPzq4hRJ9mxTL1tU17LRbJ7EjBaMUurewgQIx8
UPMZ141HnFPH7G5YNWW/5Tbdblb7kXFKLVx8VJOag2s51yiyNbUrgr2j8dx1W9Zd8SmOWRtjyVl3
I6SaFngeml2acvnrzrx09P1ERm1q2/SPTPM9dKSGaI2hEplgFV/JeCc5r9zXLBv/4KmaVod8d5jh
Zdwtt/u1lBxHcW07roKOPy1b5mmCugteiCFhg6ZA/pFgDPB4qJuW34yExyT8i0r+0AqE1aWq/5zc
eTSd7teK9E0lzn7ExhcfNLoOXuIyaeMsFW14We9A1zpr/C2+hCNXow6WSxojr+vT1ZvyXC6kgpdA
jsMF41HaV0aLJEFC6fRMWnhTkICLhYFec+X/VwEOnpn6RTocoHsIghQ+oXmOXvPu+O3oIrqWt9Lu
5z1n5ywDcUy6pyTZCrdZNkOabf/m84irK81Vucehukfzgf7KcaefVc0TYqevvA8hf02BoR/TTS9v
YQmKPAa05RdUdE5WTeX5uQOfms52gl1OJWytVpm/HDsfNQM+pEDog6PS2O33nnnp28cIH1toP6sN
fN9WyurWlXkY9kByw0AN9kWyt5Kmbn8Fccy1DXX9rzQrmcAQZwQh3gyvKJx+DZyGwp+ORUjK7s6J
dg5XcoaITS4iowzV5DMHxBQ7Qr33hGGzrdUg/DES5voSmfwrO7NUbXZw9EYPiC2u5OdIzYst8DTc
i0VR1vwAYsXU5Kdf/2JgcwpurROIwMJWLdtWswS+U78CC6ZMxOjyo6UbP6MGVBl+ec1K7pAgiMPt
4dEnFoZLkFzE5doNt1mumPXrfAQhXEZjh/lqrvnFgI09HJXNI2NfVreJ96Z8yaZJbKQHit7dEDjV
+1d6i8XzpZlovy6sm0M7RAK7R8geP3+LIQAdGcI/QJGsmvZaC2QMKZCPHLemJDzz55qK3JvlS5fO
wAwjKn70Rrtky3y+TjtrJqR4p8CwIKpcJNmSrrWUx54EiKevx7V2HOZpgheiWNqOoibi3u2pBCSg
sao5db2UWBFVj2AfzlELo72CxodWGqPNgpPoLKdiIdiukEhl5+fa+zC6SfXI41QwYlyy62fNs+mf
iCPW3jfaICj0QU2tVEgICVL8+vLMJIGtiokYgATizTOXbl5jN1kPXvLCYKxKUu1rPfQAlq7wRuyx
SYmpOYFjwwceBNe20XIFjsoMAvhkIeP6QTrZC/n/p6tVgh5Nw1Exa5nvnXTD3NGvAHugOZN06+ym
WjHl36vetm10aCUbMMpxpuzL+P65KVNGR1gTOAk4kcPySOn+9ML0pHOQ36mnDmuqvggJ10YiTetj
9xZyBhHsv8+4Ggf72gDlMkHe9Yx6oSKHk3qfZiKOq3R5srgZJsxWAA/vBHX/YBpDJoW9yCnCAXB4
ezRDUWL+SQp1An87zd1B9urH8Y6omojmE6Gw9kLchk6ctOtKE3NIZ4Bvtz70aaWatrVLyPPzXGkk
+pAtBnMtrVK595d8OR4AuoR9ZDFu25pdSmZa64lXl/3GQ1z0AmqeaN3zCuk9G3TLwh6/Giy8HjyI
DCmzlcL9e3/iHAaLt3/s4Wrqky0yohohgSsEvBobhmjb2kyvjAo8bEaeuwEEnAMplidR28NvqS3B
5X8qm4sZxR4ko+QvA1aUB3CrjQBK9usjAhmiOXBaxbNwhCqNvOO49D0SaajwJ3V8BssT8eaLRXfT
V56JoTo3aQuVykWrrvUqh/6XooAdYbvj1JZi1bB9byL+fnFp4KKEwGXkMPI1TKE0G3ytV1KRaMut
JR+pILmGItnaaY4prRenClxVCSjn5SlsU2nkf4vebVNd7D8UfEg4XVeMKCXl0gFmFPHCN6641vNL
kr/dy13KZfdnlu+byh3+cAHXy8SycoV89d+08gPSk+B/gKhY1sflzxxYk5L5KZVqZxyxIobgk1S4
U1jUgOklXosGNW3dehi5oKJYWRFo34MnFVAkOaOYXCVnaUBPB+xQZ4u+uG1hgVUQZA8Flm6817UH
piQeyS/vKyoE3LzcslbNcq5XVwv2ULp9Hp6pwhQv5hk37khmDS8VxDvHaD77ssg3yeFer38hhfgJ
HgwnZjyJrNnfbydBlmdAtTcNZTOkJn834VI1ZtBqA5pgT0CNlMke+K39lZ4NMAqmehSyAFJOR27z
GQFMT0U0ZXWJX5gytA0nRmTp801rJceFj0EFyJ3JqQQqVP/URSorYMzC4U5Jp4dQ6FGtPp+Fb1n5
mTFTFft0bJNUX4incX49K9gFVdBJqTbBLd6Ad4L0rZ/Yb7/SiGH3mMl1rYjL+KZ4ISdvyrc+SNKH
zVdN7EC5JYJPvg0SbTG8wgkFALr7L7m2A8agXG84RYTVzkG6pOoSNhsSkJqA/V+P6kplJzeyFPYa
kQzFOzh1ZYndGSNMX1kGNgIfW8AnSTZb0O7tWurbPold9Wi++aPyZMhsHoEgY6pt1Zwwoonrt2bi
Of1YhXehhI9BkHtKp7kmY7SFhkoSVnYzQHtmKBlUG/mHXBRCQPcdyX8hzM05u9R219++FvKrTb6+
wwh6ry5z6T+tpXyV8CII1Lv+fLaT+oT9hj4kipTEjlUjL8YKpzfGyP9sG8mgOQLh+Jum+CLgcRXV
nBK2z/TUK6gPPhNmfe5Q58JhGj9YgRnVVakDXqRMS1Y/gp5aHiNd6UySD5S3LV9ysNYTcnxE5QsC
SvXasNuGsfGjm/feVHkJuyTOOHwMvnjKm30OdefNm+sUgyGw7GLXWO/csyZCD/pr8BzoXeJEDiwl
ppmJP7gIW+e1lLwFf+Ek0a9F7KHF3jCW43aoICICN3qCE8OFmzOg0WlHSC4kcQYTvBo9GBLnr4Om
mnDTSV/3mJli1KCGbNHwag==
`protect end_protected
