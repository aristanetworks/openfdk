--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
XIW9ZSTovzrR5jGvHiuNfox5/s36fRFJiLdaA3ISfjEFnQjUhVbOq478E0mds4Kdjwduy38V03Y6
A/VFUz3QEhNUJXrOyeJYiFX6J5lVEcRtcIF/unr3Q91SGLKcQw3Lf5pGdNe6U5kPHD1FdLF1XVX8
GYIc7Oi2QsVLHEE/78nf2Oxbq5t5caYhe8MuG8HAt+2fHeO3qio49Jj7RY3jnpKCYCblq+bl1ZmU
GeAJYtJ5Wa/u6KWdVhZBl5KrczttHTok/HkEtop6OZAPuiYgtwooYqVT094dIZ+hc9DluAjRMCTJ
5hnlMKmBAinfcH6WmxJplZkbphdt5KwNfA1zbA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="GwQ6wCGIn9v8OxWDzo1If2lfxxc/xdtY3G+vm/ZqD4M="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
DCVDJyf1nZv03HFBW9xhyEksm8ha8yEBfXo8W3DjAy1B0VoRciwjMHolczU7mjTbnfALXc6UCNtz
R976oIWHiH2sMuqz5c4gT7YOaWO0s9KYu9iq9Uom3qsIGpF7cTnqidl+HyVTc8d4DSq0loa/MB8m
nsO4BzB2aYEGEKTgHTOLuOgbepLx8pbb+gBRZ6OZSSKrY07L99pMyG0Iea+9PoX/yymajeWoeuNO
aubF0xXfLY0EqMAAYB4mmKez8YyD0sPXKoTMDJfWIcCfrI8aDHHbjgESl3XjULaVgFSg/SxteQCy
Bs1y+G5nXZOgqyeBKN6mYBkyQj/C1YUseDB8Ww==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="y1oVskINnm4tWRaWJj0Y3YkeeKNTmA4e4VMYdHifmIM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20192)
`protect data_block
x2WQ1Hwp4pJ53R7uUee59fyYOJYx8vKZ+Ti+veY1nfYMnI37oZ7dIBLzeDXWPRTBzh2oTiv8MYTb
fAPE7SlSebIw4xD7L1J5x2HVw7XwmnH1Z9CJuayG+vSH/0ZzLzmOBFSeUOKzRVWzV+zFTgH/LhfP
XN6TNTsA2YYOabl+I5W/tv5izFM8um8gjIVkj+wTzFafyoHoW/Kikmc8GOByvxQlXgLoGJwWWm9+
QuVM/9zubVrne3S27ml8eYBKlV22Tc/A7XkT176YQEkjCW4oaEdMlzt+SZgACN5IBGEIatArwdhi
K2M32KEc6Nw2k8wHxxgdM2wzmjzfn2Xwz4yPgDTpz5AQGlLk/WtgbeVjkal1ag0uwAe92PetktOm
AN2mcEGNsrBsBPC8zhkUaxG53LfUOKbD9bFZdKioU8wwRzMpjjDarnOPBfRqIo1Dfrg3N3/wnrCF
BuBKP9ISHU8/ld+aIXUTiVW+ZU2TJS1f6XiQl5vAjKr0ZPJSgIYVwMwZfIbklqpev2OFROnLdAUK
4VTpUOGLG7gr/KVjyFczKny6QBdnKxUtIakjmVF1k9i3HXTJlDkWmidTvSAxP/6mKecHt8EY9hZR
eCc4KWsEQypZ7nI89O0WKrVZQRC/KiJ7xAeKgWs9Pjgm17LjPXB+sRHztVmDxw/+Gfc0HB/JQDxl
5HUnsOmsFg0Atq1szVbxd4qwnuKuGWF2xiNJFhG5z40IDJ6XuZooMDuGl8xeriLwsHMMrFP5B4QC
0oTr7adqD4XhHVNZcKS9osyOtPUswqlMKM1xW6Wz5dXhmqTfYQQ3Ig+rffZnJ6GvIdpSrIJnyRNl
om8i3EnoRWiEYwsJAGRXb2Ve0+PDPmSexrwMaJFnxCCAKOQEkry5wdTfGk2ReZ0uvJ7VV8nQgpOM
LC7yUjA3/fQDbPWAWa4UpKnANkV+QQsgG2MpNsNhxzUFD0yk8n4N6ANEz+rGBNx4lzGdSmofLwKS
Rt3hwJJ2Ty4zWTAeZSZka7oaGizN7T8R46Ssdj3NNG2I7WrdgjEnsTDXwFsNotb1J2DO2i6mt5Or
BSmZy7qDAONKYwUxLcOA5qwTBY8tv7Gca8ny/5UbewGaXKR/SWyQvDv9RZKNt2BXzheJmLQ4k8ac
0ZjN/14YLFmsa5RzuTgZDFdDApF0blizC1FX/6VqXX/HJIA8y4e1FHmfpL9M6DTQ5DEz5tFQq4Wv
8rJQST4Dg4T4+x1GkTQqVP7dtivkPBvpHRwLWvTGMih5gpZlX6cuHX8kC/X5N70lOt2EHkNGvFQt
nAq80ttGT3fZ3E4Dt076s/PH5Q9dAs6U14ZLCG1MuJDoDNpJsmYGE4rYE54BhMPeLhOBsodC+OT3
stzQWHZlcLM6ukvkZnVh/jCIWdoTsMggqsd7vbm92IEZWlhjN74JTByZ1QQk2NgBWV/ZebEbge5v
mxUW54ke7BpsObD5KmYLJI35i455wK2IHXNe02Gv+UdeD/kUK7uj+93gK/HgLbpYNdZYAeM3HSuk
wk7XKLQ0q+hTid5kHJD0hfXonYA9JA8ZVD+5UljlPxikcqVvv7sVubc4G9QYqi3VwOXhZjbxiTTa
vSnyBPSZyfI1Rf7pVDuseDSrzRD2XF1UDio/6wDVk5ulcRaFaPc4r3zfjqXTbzHMb8n5mmHhHjB+
pRjhXBNs3uWqO9roAItowB/7Q2VkQpIJNnTz0mdX8mNnbzXYBVpQdvTsUJiYxi4ppqmuaaPCPMY5
AqxinGfYmP98jGgEZvBGLc7cpXieES6q9qkNcE5uUPRgvm3gUaAh5IAKc6f7BxqFPgkisVE1WvJg
iFjXlJcmAMvpbTNI26NgfKAVU/KXd9lnX1hEFPDs79WGhOjlvKAoWZISbE8Xt6hBVJLBS4jlSfSY
4R0c/pTph86sN9vXI+atBaIOUoomkOeN9ArACjNq5ZeJutwKEqOj0P77+gaRLvWltg20R8A0FYgw
1CNdm54LR68y3Rj2GrVvG1iEMN6HuUnnD/+vZp0l8xItzLoFOpygfA7Xppz4UiLCDUmlIPWSOu+L
oqSBmywsA9LbTed3svX9JRkAVsbRzdNK9pqLjQgEo0JXFpu2bMd0UI5RqfkTCSYvvqah5ibAJPbO
Sjy2kKE1ClZJOzOuaYrIQXRJdrNLcm686eClzmWCdslxAc4Xq+WzaVMFxZZmxEYesKbgqkGT16Yb
yBnjQWTRaPbAPyXJF9iGFrNQNJ+elEbgjw6K1T+uIwSKE4l+sd6a8LQzj85MZdtcUDNPJDmkjGUY
dJHUgYZUIF1eSkqiLdj1I35jMd0yC2noYvCCdhKS2XfPTWqdfY3Abk+RMjvRQSnV0A3zNMjgKgss
ogCnGL7huAfwgWg6iT38dkv0ppvlaT/pl2TURbArv3m195AmPiXxlVczgcsFfCcdY4XUnH4vzp/x
OR9qtTePswxWrq+wwfsZqmKNpR6C6Ora6fsCZIbNCKoJfBNt8wSashhYFPxe53KrT3kEQ+5qaOug
UwhRgrbfWxGYgqiowFh3Qm2LFgC3lEgLt3u9nGvgTVIkg1ueGc+BChojLO9UdlRqztNwMQgIfXs2
jTTKZ4qWf64ISFuvvws9dryONvysa8KAQprO4ll2TgS9D6aEcJFb7Rh/jQw3I7Nv1225S8H7E8cM
fgOVQ/FU+BnI9fJPYh0YthPtF2qQH1f+NBclgngF0RvTnEOMnCWhTTFinlkx+2Tqwb1ShReT6EY9
Yx3EbbBU9IzXREDTusSDP/mZjkzU8993oH/vobRZMPETmo0OFKiJFa0s6D+Kvu8j0t5jp/U/gPdh
NknwY6ssG0elT5sNRMWj9wE0lShzMPJHyuMCWwwKa/2yxmIkMkwV6E6QJaKegEwxMPW0XsEWz+1i
0DBpttqgiySVeZHiiJnLUyts/t859ZzYkaUqYGF8fkuvg8xcLFltcKTOfWbT2GcuD77OB+eTI7fy
JvsNVOru9XWcl4Rb/BkGVv7PZf5yiWdumQIjRfhHMKmRzZT7c7Mwm3X9Wgpd4g6f8qsSWgvB22JY
z7qIj4ERrd98Y+CQCRy3mA9fy00mga/A0+vLEBCoZaSUuzZCT0R5YOr7g8txLoeiDpajCfWm5pWB
JEd60eoEmCJ3Q5r/2nJ9aIjAXZSR/pWkPda15OMmSj9gy05beci4Q5lfswgdkB4FjjlJn1rEGvGk
nvmkBK0e39n0hC7Nf0mI7yzVVj+KxK/WrTKRMnFAp4WvGZjfGFi1ep4IQMJB0iOX1OiekHrkDCOl
d2Ym4CVUkW2IW5iQk6yCVodREuCzSYgj9sc2y9VVbT27tX4p66tLg7l6VwoB1yrStDkLFKQnuXPY
FAzBrzokVbJo0JY0/9RFstQ3YAEHmXArT8LxKqzh848yfZG+WnwqyhtdAjj+f+GkFmYl0qACj9ys
wIAxh+E40j9JZ2s806Z2L16btLAv8+bagRqiAqTADYGfsNVNHOVBtzEDWusTbiZrCz98ARn4I9UY
7FRpKm9Vxxqm3DlV1fP8gwxNM00+NyuAVEDPCwdmv0MFvhpSTvFDDTRt6QLVF1tj/O0ic2WovF6i
o1RBJMyzcVXceSGRX6obgvxL3fCkX7RLJMu2TNJtHniqYRSFY6o5ePq7XCOfmV0hmqAsJ21EmZ8r
aaBQdsJEf2FwIo2TEJ5e/BAmagVQ/QjhPR9ZeyNiwceq7JB7JmNSBGFfoAAg8uBYYJZ8ZdbRvxj1
Gi2lQm28I8pYnKm2AcmUA+pD8i9uBPdsJyBETcvWtfUlH9JhdEpxobLvjCG8vePEDfrr4WpnqSzo
sEnyAJ0+rLCDeBtJxFPjo/B57/MrSTgrjJqwRWy3WKLt6cmaQmbZHDxnndjiUYPzyFsS41eiQSmw
d1Cvvl+iZxt8St5w4tS8XhYuoNCzgFwxGm73du0NG0Fkj9wZ7V3/95pXU+GbC2svziUj8OTnNzvy
ex0EdJm6XS8iQMDaKs66t/xH7PKhfqEyu+XpCdMitwGPuCPA2Q3+8t8gjoMcdZ9D4+pmBHjwfOxQ
SuIHOQWAUoUZcHjTg9/RJrQxy1SpKH4h5lsCgeg1iG1xGBqG3a/SQsuKBxCY4NWvH8u+BeoLlr9e
d//KbRNpHmX3q5f9DiKKtrhZXp7UM3Lqth04uASNvCJQjGq92AtWwLqZePlMgD18IYdxgwK2lTue
TgXQLVSQWFNOYiVOiAR70cl7SX6CQsMkZ3uwxKLVHH9/BwYOKbVdKhJItUTD9n/DdrLadooxGdUy
qj5oZRFJQSPA8WXmMAu8LZ8nBbxjyDXcgI0SnPoSy2ysqXl98sj97f2bKaVhTYtCRf4iFzaNZAjb
6E91wvU3XgDOzYatj9GHoP9t01yLNViMPHWY84NECkCyL6vnWfTG7Bg0/xY4bAjvfcICMwBC/qOy
sh3o9v96Zn0sOkbx948iKLYem+6/0FDhvNXOiKY8OjhirwnSgRygCZkmBSci+ovxO7TFyml8ensy
V+NGr23T3rlSgChB/o3Ch93hMLhBK9HkE8PoUOAVcmCTyM8GVBB3Cd4CP07SUWl3ZbK3/NqXIHo6
TCZ2fIzN2QNpsQ1M+CPmJtZtHEaOU0QbM4taQiLgvwNEH8vA/w/vq9cnFvIwaExgrk3mavfpGBEM
NzS/CeOBAl+QcVJLqasb3lIXzpw46QxFjSzkSATdA4plvZKz+b3dYyBypoEQe8gUydmM9QPsI4Z4
TQyIKwgBW0ayLI5bTaC2YLB9NfaB4KA9hpF/EsB2ZSCzBQV78uBV7e+z1T5narqZ1aTuvCv3XIYf
tJK3XyqUeCQmwpYWp6Y/Y8pVd+DxypYSg9NbwsICQwQ+VVpHrxyF/pxLXbETIhmXAxc9JnZdEpqS
lZ2ktJJDsUW53y5e40Qgg3hPcYG2KTiUs2QdFI+tpVnpTL9RKxKUPjS3ouBhG4o1qH5e2m5G9TRP
vQQFYBfLvwivKilHvcxqPjLGdyIC1RPP+eBisTe9MOSKxcrXHmPW0+lLz0bL3kNVIwSrATpiGje6
D9OZ6aQUkwTuajAPJl3JmM+KXWE7rsSP2IZLX6l4DqSrR0rQYswNJiHEDIfGzReRenY6EyCFnD3H
kuT3e2iHTmnLgEh+8esQnMgcc9WmCeS12oGT5Xdz2UJLX2FvIwsgLSKWGja8eyoYbmZXV8XavlcU
/SEpXjxNCnA0AnOaz3UpHXWTRxvl89UrtzapShbQm//61YvTnAD3jGcOHVKBA4F1fjAkyYfky2fT
elLG80j4eM//oizUiVagGkROpW2dnUA4tjZFWqSZhdvqb68te8FselAHklw/q/SFyg9m2N/OTiJa
UsanqtoXS5VItLz4XJHv67lA6Kz0B/jqiI04k5aXq9N5Y6txfpfmXzFztLdAtTq3GQ1/4IT9rN0B
4Pvmok8ZGeHo1b642m5nOX0uNP+oQqpwBV+Q848j5Jpr5Fo+1or3gS1/PERqnIyQobsxZfKevvJ6
pYGJB0/I2tAaUhB1N5lTrublIuRy4EE2BuWQe2/cqLami8aQ1LWz9NI29ONpzWCGIoOb2qLj88JY
kgbWaktwM2eIlqiKdIyi08lQfv82Fkk2I+PnWsR8arEOjYwoIiihiDN6Z5EN4hfC+nQznwcK85p0
C93MYbD/UnoBdNyPpU45+aEOPr3ISx2AKMf/56vXuXTyj7XP4SpXeZ/XKPu9TKzsDmbhoO+IOFLh
BLxDBPmaykew5KJxIZ+XOc3kkych4vWAsQWRq8WUmMFuomCS07TnrQ81kqZ/bBbR45Jhs/WbDs67
220dsxjccDj2/d5DCQF6p8LJ0OImCIjuXlBrWcl3VpS35ytYn06tWXGjVz1nt19XxOK194D6T3YA
Ou3OCdEx9vPIO9ZmvbpUjmJzCZ5Eto/TtgLoBjKPyE7bpRbewsoYoS71qSq1QwN0Rj+E3d1XhqeQ
uGxQfp75xkuAtSQVKOFjnPZ3cpJb+fxB8usphTbX1Yw2QO3zsl1Q12PbA+i2rnuiLio1wvunABsh
XRuTPCG38ZkXf56eeGu0iAiJA345V3y2t9nx63i9SbeAJEZRgXU6J0OU7jAJvE7ecuFevwAf8aeb
7b98s4yrb8eY4GUt8KUSrAdzmyily2FaDNZEmx7WOzt6WXAroUat3kBBvt5DenYbhSfr1ysFbefQ
WP7pYKgsq2hWTKqSnMgG/N9NH2mPcvdrvgtCPqphFwmKQVva75klIjbZ1iO/2ZPYnY2qXnwmMX/O
ggBBnskNm7sMPDyZsHEP/Eeucf3thCYER4uamxYLJ/RkjmWa6+qM94gJmO/sAk//0QdK1GdLmTeU
bIbiQzkML2ZLAlSHV36A0IgGvCUFuC+vGv7HrC29hdgdWGeAmAVeOV9RDzpZG9JniLDzqhosq3fi
3QIEefs3sI6mX8HGzl5SaEG9v9rObzEgXoH9CjTGNQ/QZUBKtVbYIcGVzyKvG0qJPdw+tRaA0HLV
0in3Jb/ZLTO9uj2yRHJFHfylfzjFigfZn3livi+ypUVcOmqrtgiFieb5sa/e+xaVWgqPzcsAWb/D
qBfQkgR7DZCX5QqHira5QlOac6Cf1OoJ3Rmo48gUjmL5+JLCo3uHUbK1H6EON0djvciwV+Bz02Nq
9ggTeNxWIfMhX/MgceApDIQCT/RnhWw/8m8oXhkUaG28/YfxRAOCaoO4sU15j+RWKHoOkYgZcNJk
SimjPhqnTxIOV47DXtn8IzDzKQTOnUhtKvU8SGS0c7LFqX2Dt1/P1pe6QqabfpWr1SVG5hkoHuYF
Uxp022/CZMTpQT6amVhSXj+HjD8yy0Fm+WOHrt4i2Q9c6EDjmOmnLbO7qxA39BquWMkosHaKsFl8
VkkuxhjyO9yzcEZEdAKp3Gy9ixK/fD1niuUCrZhgx3o93a3ekOXMaUFAqQfQhrdzM0X8IEgRHF2H
2zQoD1JnCdL3VJcp9491EEHlZLuibZjcdEhk91Rdc9YCdc8zpTv9aEV+Aw7Y8lXHA1maaIcFrkVB
CT+ykg2r+i2g+HWBqQG1rdsyfZpzDHgZHK5XDXWhenCyJc+MLgvFd5vDGe8UqDeY7UpY2GX3+oy2
MBN7Nx3AdXe4mD1QqRVC8WE4Iau/rJC5NAUHTGVST8h6luGXgvIf6JGN2f+wtOeXyLQun19Stvp6
I/dBmGC2lL321pupMLHuHTU7N12LiU4vFXruACkpZZ5bR/Gk0L/KtnQh8NCgUcvt9BlyeAkhK6Nv
IJmSSJcZCj1IJkPWUOBjznB60tXpLj1fOwCfN5SCtaePHv2l7ZaBbOF34qCkFrf9HdJk+9YsdpG/
iIIntCIdYYTV0iMeDgq/73xLqaSRfR1WQ09dAta+2lhVdfKNI62+j7WFKrw4evgcoQy5DHQuAzOB
U8LxQRa+Q+AwdJj/+Q8ehKf6fu43jdLuSTJQscytK8oZ0hFEIuIcBSLl2JAG/UGqQ9OJ9x29R0DY
qz1RRkkQ5KZ3XywdfpuneMw1/oJEvBL6jkywaXV1iVWKJNargJbkUpvhGA+vzoTNpUHf+HNEP9RR
NqyN5GBXNh08/CEyCxu6vSqvvSaoUvPsUPc23TIfFzONYBGSeUMoZ+azXexh7yyUvjGb28XfwgcK
tOSZhYCheMOL6rch2C1WdYehhL8m3PKZb9gCM6ZCYGL0wrQF3eWYGRu1gkXh8tYwOokh7ELz2Zjo
FE+tqV57QfTa9x0vlJ0rI+J1sdfQ+oSbzfQf/HP2mccyFjRp5e2SjPycapSqSSCKWubbQq83hwA/
LAFD+DRGuz5XSH22iEkTqM1Yy5Bc64y1/aNyODLDZnok9r9PChcfGo6mSwJa28fGNjA3hjyc/TY+
3Y8ifi6/byoOeT234cdVkEeJTKhoS0U7TO1rctG8JiF0BFWnQRVaIvdst0XiW+EWtgiFT5V2TfwF
kOzsm2+/FHIWIMY91ANavx01QTnSe2S8dadTVpwebC45qnNZP1aRLhZvwCOMsh/D7WGUny8wd2z3
TaP1zVaIfFzaNJk7f3/eBX8GGd+XsRz+X2f7HUHP53l4wPanPlgB7VTN8/FQ3E8HuEu8Kq0+RTRL
4jv6dwWicGKHuSUFffQri0sS0PvQXEMi9TpJ2hHS0Eg6Nw6Mwk7VPgpfLhShI7dYkc/yyQ2K5lIB
HXOuN+QRN+QXdV6tOHbOw9ZU8t6S8iLo0CT0UjRfAkseRQig9ZpuFFCO2A9ImXgG/u8uW4dMZ38n
vKGdjhYCJoOMk7KOBCdhSn+5l7wDEhgAFdswIXX0oYGG4MN9ozhtzJ/NNKKHZkDxjXjRwb1QJ312
oHJ7ZRY7Tb3lNaMUJv86AXiD+sOlkVU4pbMAnMr38HDRu8znSG+Ca4LdeHS58eYhwABuByYvu5AO
fghqspKT3cJQ20h7LsSPxrw35Qm7SXEge/77w4moeyeP3XeddgS3t03BEWbrl+BWVVKHzHh+m+FR
RQPEG1yuSx/4nV3V1+8XAIbYknCeeM1tpNeobHCfaGpin8In0wmQJ5shdBg8zHMCjceFbp65eZ2X
xAEYqbOF1FMDdSVQqaavhFgkPoBZHbolGnjrRWNpylE5d8+f08jG8x883tCAtP0H+c3CP+s6dSEP
b//WKZi1QeHeBiYNDAIWuQCtD2dMeuUstFSCtRzUoYb8rl/NDeuxJ/ph7EhVkuLm4OUUDm57aAZl
e5cuyiyGhNyMd/juTiF5r3BkgJY0bDgmyzxZESZYCpdAE+O8sMf/s52YA60SS2uXXfM/l6fCVbQF
9ginUSo8UX+MKCyqfxd9rmBgN0yIf359tBQHigK9KiBsggQAl9dUL3Knp9BllJAX4cug7M8DID5d
ybn25ElAQRAbwhQYpi9YJOxwFW7/zQLZmrJg3oj10tZGp6b4/9ahAl+2xOuOvkiYF++8IRTA4IAB
XhOTSLocvm+XddE0RPz4/YKjprSRe6doUAODiZYXH+ZEvwfKvavhzmT5+bAS3URrWtHFGXfKH0/S
w4lSKXN/Lw6inBlhFvvAEg2O7fmhlLL4rBXQQ3FLSI/Kquyz7ZJZuQLISDF+3dvdkfpCnqWHV20a
bttlaLSCFEQc5GwbKNjBB2Rw5vEsYZWJnKvkiFSaIGRXaxq+MSMXekLJnlwSkR6OG8G9PaGC8Y/n
0Nsplj3R9mKWUq7+TiUztPeGW0Nl47YPFl9K3gfTC81lM2jd1UhmoC87rR/03Zo7kq2CpEBaBz+V
qsVpiAbPWUVZ1cFxdR6XCK89sjNMLbzvJFAtERf/boxmtKE/BiLLKyI2SnPVF5U1o42Pl5GMNdAr
tHS15Mweq1z36DSBWm+qmnopyA+BnbjhFO5le0wYZcPZts20ZJpEFp2D3u3fwkB+CiXOLXM19yII
PNh6jjsuETBmjVXCAyq55M5B1/FWuu2e8QiT5j7yu9SmpKqddjRC1AfjZZIfYN1qyrzway88IkYX
GChkVzxNIQ/2Xo+qTSqhmi1zNVgLvI3pzMGfKL/uyS2fffVA3Tj6WYEeggPt3JBcizdKX6TH09y+
H6aiXB9yzSWGzynu4WID5eYmWW+ugvTxibJOARpBwfcKa/90d7nbdqBikOBxnoPJnH7czhbLa8Lm
RuS3RDY1WEe4tiSO0P90DCvMJhSPEo439o3YjVv/ixJfJlDlOX14327ghaSUuWqbmV++xE+GgO7b
onmIAHPAD7nW6qvzMs0vr/nMd6jqfr5n3eRewNpbEW85h/PHT7ayX/JWgMiL7HCRV1+H5xHbsVom
HRNjENlBW/qiqGrFIbwot2ezivySyF4FIEPl8iupvstbwg5a7lmzu2LKqlZ6O3BVVGVDyik2YpEM
ebf/HER3UL/GwledRygmEr8T6rh9RK/SHYu8fHLhAgEDmFFCI2URz/5TwAZWqMawlxbX4e9N7niB
IUQ5BiQACyb5/RcX2/LMMGHSSWHt0zqCWUsOFI/J/6JHiojWjGXtXHQGXUOYd26g/xiYyVO327El
w3i9A7VYnfkb4HZAWQzk8icFGqorfSPM7Hui8kLyNmYeFW4KhxyyAtRnhk9UItvzwNiu14xuhGUC
Y+7wfKTAb/IHeMIzuwFCf3KVvtuO6EAa53fZKYjPa5iUjetsFOILAIlSyYjufyK7xvVcaeBPEkj/
CymPvBJGAX2QLt/3T8vXJexp3hNnFyqPmc9H0iVk7H5cAh63GhujKVHz894r+68Q9EdqK5DOdFLF
TVvH4SLgIfg+t9ykAIQdfQhPsa97K9xEk885pQUiJYdUkO1CB3Zj2XG8GujoaBokbBan5bYSQsay
UQE04pDKRPjUi/XZxtkBXhMJDb2IP1k91LahLOi2tJJoUVvDeCs2YBi2JW+21waYqBOHCf1On+BS
1INWCTmghJbelHmTSqjSJM3KtqqUY7Z6Z8SZBaEgWrGxQiyHvpbp86QIw2nV6SurOPchUjFknYsb
ldhStQ8M9DSVlDy+47bffBtIOUcWtIDeGp6Ze8wPEx13kV7VnzSbp2gitbTD4VYX+EttTg7E9T+h
HMXm4OAYFxO0mznbF+mXHUuo2LFcKkIUnUIoNkFGuULT1njRdq2Hntfj06k/22Skc5tfz5PecEAj
aNCPJTfBJgGPMdxFOf03e9aRfms4NE3/ryWw55p01QCvN3ek6c4Lo9mzmd9xJjOiCnLsXl+3O72+
gOBGEcsWPP70CvHzsBhaC47jekHl963EcMifYwx9VLvac4MJYYHZlPV65GQ9IUO8+YnUC7B0NWjg
OQvhKnKrH3gj5+rPow166o3LBBD1bOxjRT0MRIm2sk7yEp1opgfWDTUz7M+gifW3OrTuUfOwK7aM
j9Zmzcqfp68O8KmVEBY89hk5Dx2CkGBxE/LX77T8c08OMu89+j5UgQrCuqGYv0VB7FM9QFd026Ng
5GfVYMxOc1rSo3SoWMa8ai5Swjndhw/tlH/1f+YQVlndVe03rgPDy2B97G2vxq77izrVT1gZKuk4
jSSlKWNvntS/RqCoI3uDxPCdVuhGFtKQ9U8cw0ukS5qg0y1fro1VrsWsoOAs5YeVIBxgYoyKG6AV
yzr553trJ7eDvel0yZxnTIZYLw1GZJKuXNBP1qQnJDytLR+iwwN+PD6wbTJwx9RlHih13qiTankj
MpePuVTUjYZFVekMsBViL6pISSztyYg3mKrkt7vV9P3IKhr8RKni4HZNtsnFqOYOCQc/I5tj98eY
EeRFzWNlF6DZeDtKyyRLlTLk8iU9C7NzP9CthReXqTa8bNUkVPHPmMazcfPcYLquX1lzVdRnNUdT
5YsDp4GWzKzyrQUH1nRQEpQjJX93tB7ayJWQjZDsuGZFI1gJYjWM54ETCEiciAho6BXi+xbZMz5F
OqpGvi0zvKHY6a8I1TyqXNaAXfp9r1VMw5qgfZEyBEb8A27v4LdpmCDDxky20ENt6bGhrQiWw87W
La6SPw/VN9PmBWWfi+zXIM3dnBAJ/NObIGmjWlF3FVlTJWBIb+uDMpJBCTlzM65SlXp4FYIczRlb
fX/Tg53ZVUMoV+gGKq5qVFABI8pxWNjf6/wEQaleay2Hdlt5ds9UYmtXTyl2AMJj5yHkMNqFHAqx
Db6oKDY4Og1KHikcxNKwVDhEHKSYXbV2ALLeFHtl1RzfdJcDwTylHQ5bNSrJgpNvL0uVF+kZfVeK
iArMdyA7awxgVKlRKxYX/ZBnmBeTRfAW9QHNWTKtJeKeARixogUNop9jdLQaiHEYBN2PPYKQT6T7
8XUEHaowFWAkDK8FbX1mcVi3sVphZN+LbrxHYsL3Y7WgqXtcrbAlqm6VXQD6gQxVlfEgczqjpDJ+
hnAKNAq1S9gVr/KCAoXLtxwRA2Qx+g9MmJTWr/jRlVxNHXoNlP5x3/smPHUHHb07iujyMPpNgH3H
tuMlmBtzPjXNNH9+ZBby/7KdgzLgGK3amBPo1j/aQyieg7+eKKy3ORX/5rSItRXvUxjYQX0ydjBv
v2Sva+A4VScUSttnRkVPhuBE5HUSdSyMnVU88U9ql9sxUsUgKoDyQn5GFTlTpmmf63RNOtxlWYEP
A+QnThK4i5iCejbqWiGej685K3/C6ENuD9Hyt0wU4sMArneFbO12tRidPIkKC95kO07Zpb4pDBqJ
byDKUsWNvqpGMSB0prrEjbfs/g9KjZb/FcvbfITaaQtD+raiuA5jaZKkF0Zgoyar6zRBDnP/xr2+
zkuuIzCK5yMgsjnrldYlTcrRvulwNozsD2tQWrX85VoQidZyg7zF691rMHS6rpRWNLTNg/kI+aE9
jnZdsFtv1Or3S9dMtdPWCluuzimRQaaXnep3Y6ohMWUxOhVpDRP0m8sUd8OFd2IxPLQeiTU5Bdr1
8Hn16PV4md+LREIhhUo/4/+IeEv0+5sQ+79HGzHzDqGX8bprz9XLFYjkixTrKSWznXE7C4dkb1II
QHUKuNx2aZc8rTCcPemNhdbV4rEMq4AI6pazB/QGZMvtcFtbCPbFF+8foIigDbZ0o+WGgpgsr00r
Mv74AHwPCDwPYcua1DBCrNClVeb7Ug65tyO3kmMDH5UawxgUyjesYHoLvCXnu8p1zGgexRUk2IH0
+grRzN67jUfg4EQRJXCv7FPl7d8GdRI6AFbvBoo5E2PVNVP+ym8pVhUZVZdJiHjInooSPHOkjObi
Zz09eUHU8eX5JnMKLfjqFa6whunKM8ptoKIp8OfBloQ660CZ7vgbU9bc/XLOu1Pb+4plFa32upY2
f/0NKOohUF64zQ0LZd0JE0K6XlhV+FL+25dBkybGK2lSz9FnxMftMax7zj0Czf2NN/s46vASdWy3
hZvyHYMvnvEQtPONTUhuhS0WtGcRO8ZnZahoAobgYDckjFM8JqnkNjwiWNtM9auUFeyzwsvdlbxV
z5cb6Xs6JXGnwKPvdY+TgqBG20KdjfWQ3B5zgyfqreyVAqrEGIJ3gSh92uupKkaIHJkrorudEmSy
+YEHLEAHh4vmsiyDFgidMKa/N+KXzAvUIv83Yj8pCiv+GOUHMBdEF4qF+T2L2GEZht2ZcAGdvc11
ke80zDcDQkN7Az+cQiC0rOMiIDX20L70DrnchJTF2iczODzTqk8oFyugUaUcqHjpvoRTwjQLbCzI
jIbLJ5BdfBOmxxiDeBrVGfPhUUdQGYnDaZLJiZHpap7enUuKYTAJcpk+BOnqKfOQY6zZNUhPY4Jw
PHauxNcFoUFNK1CYwiYZyiYGhGmoOuynoxnSp9U/PhSwz4qGtqJvycDY8eysB3tV9hAkxZK/qSrW
fdWXenbjEaxmiwxmP59mZcmVyXKNHIFDin6FAKPrYVLPOf37dUNoViPSzOcoBpTWAljFq7dh/kXB
ggvNANCM54MwpoYhkydZuV+sJUgRnNFBey+hmni56QaYvMNEhJpn6FY/jbkWP0Z22LCYCat59j/5
8aOG1tZnjdkN7WKJ3T+c4SKuyCNcuufNf0v7vevYZfuUOUtNXzpoeTp0VBPlcCUyc6OGMttNXXkF
BuYGHXJfoFcUatPRcN+g3gwvzYYJbuI6nWBZjpC1IjG32WK3ZifKU/moDF3NlI4M/opSi6t65ns8
LvmAO/sG7p8WGTs7PEqkArWK94iMluu0cGsoneuNkPyDNkg2Z62I7SPyCeEVLh2JdjZFhp1ah10v
x3IZ1UP3qqHbYEEMoIEo5Al4EKJKeJjJthS2uhncWvMxlPGeONI5sRN7IS/0nnVyIWW5HLzeEJTb
vsJPly2LRmqaxAs1GKnXQ1B8zXvA8lKdybrFN8QePi8J5LBlPsyOecOV2/iAH0s4GGtvPuqbo/I0
v9Up2EI3hZ+U6mX93QkMJPNVShEvmPVY8z08nfM1m9Xp/l+TpT64OTNhhlZbdOecGUUD1PIxsbFv
Ia6wpcBi8nigepFAD75CNSuMotUQgP6PSHo+nH++larwNiwkD19ruqpUCyMMSjjoqqCzltotHPE3
IqnztgIMhbLDrpjZAVWrarGf7bnjxw0TUmsuanfDuUK3AnHexMtYRLDBrP643ZSo3z0Sm41tAcUv
S/Zc3QWLLp2gBEn+aL1uoA1V7t+YfuryhkiOp784K5cT0veyhLu9YASni0IFwEvkWXy66gevg1+I
R42KW+Ds9mEagzn2Zw7d1RLWpda4nTBWt4wYIbfcCY4PnM5zpQ1qLp9D8JjjJgbgNdZrAYs112i2
jQq/2VEl30AA8nAHwW+/2e8cFFjY4MUFOcYcM6V+lIsBo+K1Gx97NI8SqpNcykOa4aaJpQLcpPC0
+XCmYYuujDxBXAl3SiOjNIBc506HBg0Iru11gPLc+M4pIFfDaJeTyBzhEv7IEKIxMMc8Dw4id2O3
yhfTKHViPznaYyWRokELNC4lJy5im5RmSXQ0SxEw1ivyVg3weLLUUmP42pH7OTklYvRMoveadMZg
J/KiERb0GgzuYa2/OuW0RLpgZktvyNDw26Iq0SicKn3t/KChbuAtzKi0oAGVNjhWTBaW7BMs+Q+c
EYXRQwHY4NUfYrAcI53ecdk3/iqw/XgAixI2pGZCGqodbahRnU9cgLb8gy459vqvK6CaIC1DCnZW
GyIKuAD6C8bor/WPS/amnv/GYYtQAI1TOD5XQBa8vknqaZrZWMmIuqIbli2sq+PyjaekmR+UIe2x
j6CV+XGlfRwX4ADD2KVJNl5s64Pk48087CkJ6cqOC3I+vcPGSfzgKB7hxX83PcEkQPtgacg2Jw5t
JMvws+4Ca5ChVhDi/AFMw5/Aa0DxAdxY5nuk1SD8kKRnaXZ73pnjUXeAfmQ2ZFprtaXd7rjBZedh
0Wmd7EjgNZjfk86wNle1gYF7d0l8KwVbs/gw4QkSXP3YKwyvj1Y/GJHRpPYV5UqkkT/sjj8fQ7Mc
7wnLyNgXgxRuNfV/lViXzIMqObxIisbjrSnI2cpLvddMyScnBcMIDAxsWq2hVyRyUkr/L5gKYclr
ogF07eVu70baoIuPQ6c0evnYMMlbtlqEiL+pZkEpBoDa8srZQnQK8C47nufvqMaKErDWfYc2SXXH
l/uXY399ag60Jp++b46yIp+Q984PgbgcYiMroMtzwUtFioPnR13GHe1hdOM7W7pTRpPDTBoN76EG
BcDXqMb+cLuXYqTRaP79ChAmCt0/F7dg0SULq54hpeiYnM0z4Ruxrg9aAU2l9L5/0JpnDNJPe1Re
s36MebL2tiOvr90cNeBECBrwk7cdu0bnUnCRYHjCgkJO2/PJlLRsKK9y3bokqL/oDmGZeHbuUkm0
CxkMusvZJeUFek+b65ARBLbEbu2+T19hKHwLC5uAL0LZTD+XttuksPLw2FPYnsCeGy815UyYtKsZ
wmdBFdLLkCkOIaBeCBDALg40/gnJKeVlBozvu1Jpp91kf9x+4PIYTk/1z4DzOLFmyaWx/i0dN6Be
/QOA/TR0LOHo4BZamGq16Lu5oRVpjpkLc6nWPJaHAUAQwf5GYnZDSXu202l+MQYDhxbP8a4q+dmF
y+yzX+jlqykXJc1Pi0aHWR7Q2OdFV1HLg073eAdJYN3hYRANEFJGOscAFfw82KfeQKuP7Nx0BHhB
BW4P/psijNwwXOH3s8PwkS1P0GBUz058HHnXYTv9JezY52qU68dknoAr7wbuktMxI3OiGc4buyto
WucoysDfhsT0g97pUrp4CiDchXcZZWjpjguw7Ea9dn0o6XeyApRGbgSR88EG5yrykBOmpb6ZqMLe
iMwq6Puwt7sckjJReyD0zJ1ohV8kzTl1BtlWK+z6LfwXUWS8TMdW8hyrnV0pP1zSlFd6XQHUZTG+
Aky6pZ2Br9caZfesN1xAhGOhlXX5ZHFMVnH2beF9AWd5rcpKYrPhSq5U8qQwPmmcllIF84TSRIuB
kg5coOR/JW97GvPWxAKI2CSmJF4uzlxmVnkce6OiI3hX7uu9wfM342aqZ4C83769m/dk3d6vLFct
j2bZIvx3AvCb6nRFuyKqgotJ3rKw17AtrA2oV3HL+OH7XcmREoCB31Bi2wv8thtqtHPA8i+vfFXc
Mk+q+LSyP/ct8PCCuQGwJWGFNCn7PkgF3+/MlDWVDY+og5iwIYgjY+QDD1XB7OpwR+IzschFQUle
Lg+qBKPJUUFYnnDoqtAEm4o5bP86PM+osbffQ9cb9S3Ew+R3ycbB0QT7+1oeIRFtT+5Kkdb5iZ0T
pe8AwXBOPYyk3aUwxJ972OVMVLTcI67OJGLJ5XiyCeJPpLPITz9yfoffalBm7uytljhoeauMngoL
Orr+UmYGJf5zeOh1YnX8sREGMvmFR1wgfQZFhVJCzYZooATZoakexdLd/PMFZL2ILL/Q+Vm6uTqx
YnVves+vs0gahthRzk5VJkXVY9CkVdgUdcXDbYZoqKnsuLavqlsrS2d7ArpMfPtFQxLi0GJFOyPF
waWMWTx2YaDGn7uGxqD8It4/6/XaJnXtYRf8hCaSVaxzSCrfEqh4EToFXDKYGScEZrjZuaEfjbbw
MRXACfyASvCAaEw4YopzynmmnAKl2Wj7W5MucNlhqhHMUC6T0VVEeykfYdCdcRvhzkdTHS1JepWm
32j3TmlJHJUe4KFyR6ynZQ5+vG3inYZCa080EgEWRVjIfb0Odh6zPr5Ye2myah2HO9UGOSPytslx
t2d1EcsYxVdHMQAqiRDiXqIzJBddDjlYxXayLm/pHKpmoitMo8wWiMgF1xheoHnoLN5XeJf2SWpm
D+1yep5EGPsW44tD20Bqf6bcqPuDvkH5rHdNmWDjvAMocEn+6O7+ckVAts6cGGGOHjFs8NwMi9Us
24s1wLbGKB0Ykwll/p4zdpb42G880KJ25gaxJN2om5NWddq3uQf7AMUfm7xKQFqZk6ZedCpxfV3S
JWcmuguHPmICdFQcqdeIov+fdhhkHsGvNZaiMwwaB/5e3ZlwcWB3dCrGDx+spNIqjd47Pf4VxDHV
fS3adJcYHR/qy+mko16CxFvF/H51VoSi2rvTFSb6TMrpTBuciufWeL+JKs/oTOCBtfOoXsDLn7gN
TOo3EgxEOwGBQ1lkmopIgKU2LCuW1eAX7mPSGiUAl9UstgPAVcgu2um0NKm+0AjXv9S5f7NsZiG6
YH1arzgz1KvuIg1Ow1e0z7lTplKa3/SS1Na5RjTvt9bRLty89ARAQjz8ny10iuWZW94ucGyw0Uwf
R/yK9GuU0cE9qk2McaZodOC76pU9oEH1ROdqnA6VNmxm7gNpl03Hi0J6RK6n86khhp48M6wExtma
GPqQ1nCIq8uq/A3v+Lh2GoXHN+rFSYVr79F4iQHCsoZlhaedINiqAaNQuKW4KdMTr6s8MmrSum+P
JiZJQb1poHaU4U12bq9TT9fqOgcQCiMVop9EKxVI+hByfI5TuQeAeG6A6rpE4xdvfZhuYuUtehLo
Znn3jvNo4uOCD074b2K89+Jhr0vqWz4rlfO2uJ6lCIR/7/8jtkKgnQDE8yCEdBaZnDE4BZX3oAE9
Q2eo2Fn2Aa0BQmfdUMqh6bGNpOR8sCjq/h6Ah9SnyHRP0gggjQUjsHHlOKvQ60F/mXXlvTlbHLH7
PG23n9FYCXbVoyzQkxAGqdYWXoeUdGezsgGyAtQ7+g6YBVX91d5aarEUkvYTHuMaWZP5EuNzIZYO
MoLt4n/25wdGfu5ZHr4qJ6rwmREsFKa/SbveHPiXQ3Ureh9aTxyoekhZpTOUP2xnwgLCx3EyqLhi
8LwqR/DlEcoUGEvZJr7D6MWbPczFtyHVwFRCbqvmMSErYRVxzhEpIwzhszgmbZUseYQrvlatJ7NE
El4btfTkE7LgO2vqzNJyyoQwDE4GKKhX4q7DheUDWXgoPdMqtqm+kwrKymnA0WrMQh8Tpv3JR6+k
vyvyzwZ56i5NwwjNqZKpBXeB19qQvJrdZCPDyEALSIrzNfxjt539xskk8zu+bGrZ1vuxIT3Ld1UR
XgB8bjFeDxSR9N9y5TvtreJZn8MwBPmYBBmJIb3F70m9p5zKEQiBmBt8QjVHUz2lVm/eAtSirnt2
b1oJXAGWwdG5Ik78q8Ii+ji9W/NxtmMCF84fEVi3pzXEPTzw9/uuFlQFCKdlxtNUqX2JiZlDmr6y
HmsbnP+OTNXs+g33tEcpnT+fAZbKyz4bRln/a++icAukZyOZ3l1qqbFXbcrlf3nFkhFem+S8hH7i
QMEb+Sra23Ko8h/nuf22nFQooz3Hdbskc1jHhyh3wTmV4YvMSsLewOwwItHbQPCo5tBKxItVC25Z
jembxcup5OY9MgWwlEK2SVFXjL/uMiTYsieDWiG8oJi/HU/gdVgRNWGx6ObrxEoQGv7RV7mGeom4
tuDTyIdz2ZRihZKOdEPPYeFD8wgygIR9pdT4HgDEMN0pz56ctqfox8pzaqorCVrHTubSJeTEfslV
CrlRyvftVcTsqdF3KSiipJGGWI1y5GiVGHithSVdJwSiBTFyZTVFooggRf23PMRgrWG7yMG3TJ7V
1cTSSisWiR6tX1y0ICzzZO/+vizRyZD0oHfODD+dB+Qd2tCltQFsYa40KipxgGY0fqODHWh75ryT
11aih4j8aRwH9BbGH7HJSDaQ6zAYtVjih62fqA+LTNwDOG01+Y3YXTkEUaiAWvc4uAzQXA4Ru02C
ipFMuMcbfRjIuh/wOMtsON9dD1XmldAAC3fE0MJM4zxzcFVMdBds/ZzDVytl7JTy3AOjAnEAExzI
xZpfEtF+hHI/VvX+Ngy5WzHD0FF78XO8f/KhXgSo8XecTCtDhrVw/7z5m1AHQY4cG3ELQVvvKXin
DSlhPPto68szx6Tk/+fK+2ldkgFGzsL4GzxpejmpUU/SvAnqHBi1RhgNQi75UAXOFbOiBcRppqTC
Qcmv2XV4EaTy/prax1Z5D1FjvduK/DG8MiWvjNTK4CS4M0+lH3HtLf18yNNCvCC04Iyhf2JgbWYr
7nEIz0LO6cReVrBgtwqlReGs/EBWPKYOOGqvOYMfwvrz9fn8C0t/vJGGuq3rtla+x/uHjp0hZMll
zh3gW034daqgqoR7Aavg5UlHSWvK9SFBnWPTYQcG985oPBwt6vsn5Tte7tI4jNqUq1g5gqnSvj1T
xPpDdFHgCBYv9DZGwDDf9t39xCFRzX0AKsCmq2hW+jmjOjTeQ+bFfA5qFsVPffRaJcOGN2WVKH7H
1ZZG9eb5VJ3jlqnLv1z5DB8mR5yNcD+8Uoty6i5imRgggZ+TeCi/ZF1GfS8+U2cl6x1WGqFscc0A
y5tqyPvlPQlAYCyPPxL/wKmR8qS6OwwnP0kLtNam9b5JkgWeCF2t8VB/EL3J0rBs1Fqk3ML+i1lu
ublLFrnKsHukRpDCZ3cfmk71A77+Qld84T/SheNqX271yThDlaMtQgVfy6v7RWK7zZlamXHrz1eE
RCcc28ROjqbE0D0WECVN1ibO2Qxpxmu3m20o3QOIMvoebSPnJ+L4WYZwzcwp1RmCd+rrnhxbq4xT
lCCnMMMTAxd0ym6A2wUenpT2NyE21YrvaxhToL9d3KQKeG2DzW68j1AxBmqVh69mr39P6/zA7sdE
Vd9jWGwCgQleqUDp8MgAOxTrv6QSgqLixUIVFOZrqKWhH+MLW6AaKz9FyjD4dFaRT44FvjjLCia2
T66RhsaRrOv2jtbuglr/Zby2/ZGWx16LFZk8VGbpQWURAV/809WYU37+HPbE7OrGcJkYwWqonm3E
14yDCTLRnsrBShI0vS0OcUEUKYZCo4EdoFWaHoeRobQiJeFeQwmMigBvT0anpNmJoD4ZgcbmLobs
1PBcp1WaD8jkyuX2ZFBnzu0ZO+hhkbK0/j4iSQTLU3vfK1cri6oqXKm2m0X6iGHDdLZpFv7ImUaW
p9GV9LfyzI/RJaCpA5i56Ufdm5Ye1DZ/1Q8f5ZIRbJpW0pkPkRM4bUFkmWypONpuJAO+tWBe35Bs
DflySrA9Bgy9UdfPi6+6I6PUYZiWzUWJ4G9bHtxo80ekN+WGT4DfZOMcdw+rpKZw9v/+rLg5evRw
4x3J4EC78bclkucDYG/IGiv2dPmu8UKq1FwvdgtB364JVYhKGGQda/o83TpGrA3IeP9CPhy3c0z8
74hLuqsgqzujqeWpd8Wv7ynZO9kkBACbRhbwQrp6a8eR+u6shY+NS/W9DqfvDkADDw7TgcEgyhqy
EsWEUN5Ue77l1aGaTBW+jRHs9JVjE42ZrRI2aD3ZHhAR9uD++p4Vh7xrqsCg2E2rckJTmGjqf8yE
TfLVixRCP9xid5j3nI7xJB4gZNHpQ4TmrjMGU0w+SO/FHQOUSPf6xImexYBLpje0wqJHvcmgR1jb
hTU+pCy/7li0TM+hp5/Rhzrab7ecrgQVfR97IyBECdwu8wKN1HvfHn2PZOqGZyWwS7vCt1yewBet
i9W0FRSiHIYZ278cDv4qw8gma0oxPYsnbh3kSjopLurmlMIEEbzn23izgUP11IeNTuhj8118ceef
ZPtbo6vocOlGhJyHRrtUx+QJHhW8KU9VqFYrIwQQEjNK/H6t9RPUEk2G5og8OPMeJsOEA5SqghoK
236u8Fs5qnJ1h9p193r8m9E/Vj4h/nnFWQPz9IFTQnWjIBpsoqLNwLPE+e0V4tg1kSEN79fWdEMY
tvMJnQ5ggtrFiqLgLP7p5UOGl9q7/jRWbXI+fAAXI/43BmuzEronnaeslL5nTbbh6n4fXCB/LKRr
guBA8GPTENuEjppEcc9xVmty4PM75GQpSf6d/6/V+8M3Psb2kJVcMpVPN5uk4tO0bJxCYu6ckai7
MWPNIgLSsxBHol4wRgbubqswo6CjCkujdBrrLMk1vNN826jUBqxB4tUmg6do+OnXs/EiF8sZTZMW
PYrVGvZDc7HrytKRqT4Ephg0eE+W6jO1mQnLMn3u8OPyFxfygVkVTE0ZsDU2AqTYwKxRI0OFUp5T
Tipp+ZKz2lyKNfarvgcIm0EUwZxTmYvD12MUFvuhpj4ezKwiETWbhLTs+uYsiole6fYdxWM9AAY8
U0l1WSRxG2et510DR8tAzAaHSdQVpFf4ybqdh5JFMIdbNeZLbRaRj19qBCkia0gQYUeA+K43hRDD
D4dUfck2L2LYuvhAdEdX6W6ZGgE1ro0mYSA1e87HKYC0IuDAFqLFrkOVzA5sLMCcikRgjeU3YxTC
y05rOtEM/Dddt7SfdynSP+eHb5p3rjMJ5EwtKpENPLO+8VNhJsB94By6h0bEgDK9dHqYcwnVDROe
Mqw+6rCGisOfJAwN5RntgVV8zXbZ3erPgQNJTE/y1hqMRBshh9thfhROv2b0r/Ks4qxMCPMULFia
988apzqL86VKjPnqIRoRN4Pkn/QTtnWLEy1Qm1i+TfyoVGkP1haONW741eSIALRsmaDuRqJ8LHIf
9US9MGFb6ajb1K3ZbzlP0uamsySjB0Km3p1rPcnAlkYkoYh32b8yGU6aoBAP60X99VO88tWB/+R8
83nR96+6eC3pXLV92sWllpzqjNBVub6EjrVx7B6DsscgmJvDmfV7ldz3camfG7EapDJuFG7ZO4la
3FxyBUtQXwBQwtNGoZqFC8R0YhzHb7UHm+ExV+iFhEmrk8tkmKysADDQ+lyYFXnzI2Bo3E+EZr/0
pEjjnCip6jirvTz3qJWyxPagfbtYiaLobp4kHWKNbn3sb6KQBhSXTf/S7S1CGDU+2pdFoipaVohU
qTnEYBPGaUa8gCr/yb+roj0njbfADEWIWThBzJlkroz8VAfEo0rCrZhqsARU4tZJF2nfQIWt+fVU
sI33bcphtse1ORbTYNrPT5rpPBogUizcUmopTDPt8LnUx/lh5TA2l0xQy0mAzjeLFQuXhda/MS7U
r3mNeAEwJNhFnWFX6JN1JVHMRXab9gBtM0tVhd4thiVWtWw5Icftr8yRfHTdTGOLK4XzaO3eOrXH
fJ+g3mUAUf54LRDv6zcV5ggkkRh7CfSSSy18sBzhCPFujgDa6ZCt5vlhPb0tX68MwWxlWCIXTXt8
faE2iA2XsedqyTO+crpuC0thhn+wtox+7Ws+gyj5fjkYbnA6yR2zu04l8/1UPdYKQIG9b6+kpXq8
6d68qwZdZv0hEiVPgOTi4s8J0ZJe0Wgz0XI6eSw8LIDmxyFEMQSbDtBKMSqAf706LL44Re631UxO
wE+6oHFGIvRth8bh19b+cR0U1TqEK5/aRS2ta6tt0o84jH5rGL4SUzHNPbRZv/Pww3FxKCPSrmcF
/0zhAvNqDS+lkdFuuC3VxKlgDqTq90/a+StXpdcHzZnppYEu0uFyLrSkfFP31Tstm8Tm3OuTjjxG
LFC4rEHp2o0vwfzqLUVDIlRc0WbdboHDOPpplZXTtbwrD2EPCks1vpvp7WCCHnGZV9CNpWIgsW3S
4sVzu4Icjfp8f8aaaOjwTz7XprBRjmPWffUSR8NzqgOZghXhl9gZQlbkjcyXt6wuHHCsxYtwDvsY
ghekHsKzOiuiYQeIRKEOORkl9QAy8egj922VeIrDaUtcoxq3u/WgydQTJtPOIp0oNsF6XZjjZR1V
0FDzLhz5vRWfW6dRi0jKOxQWMxMrKXh3hIHOtHjF7qI2WvkvKhFmdTzFtTXOjasS7/N56WyJeqDa
Ao83k3tJcGNE3YWgoEQcP+nmXwR7Z4XqxF/5ZjMifHUd3vQ/BQd+29mwUpD1RBgEvRXAlHf/ndZa
RQDOY3rs18BGsTp8wh+Sa5f9lqJpv37wh6V7OQL02U8vNOYBpTx9GDFe5xVgdCBZUCml5KwuMfvL
P4Zklv6dFdfgiqAkKZS+asTz66eGHbE9CGkjHwKnknyAlTz7Uy/YdpIhBO2/pVShbnw8GlqWNKPk
trRvdHz8KplIdTKnOysrNacozPzEIql5/HqD6I+NioNkUHeZxGNHejT8Oha3b+365wpzOTV8z/rX
zy5xI67SBp7crqEfiarx8uMc4iB5yYQ8eKt2/lKQKTAlrMl8oDtUL4pKkj0d5n1or6N+a4fDMTB4
tgw8ickybMcWBWjeOqSPlMHDtJjvUc0CBosuchyh0rBxZITinvj6CSIW27mtBCgbZ7VF/AdrZjhq
y234pD/BR4HhroNEtqvNB5jxnRhmJIX7eD1mkXYEsMVhQPk8l5mLiryRpcx3NekASpR+TEHH+Ej0
+WiBxBjZelPZ3s3RGt+9x8iG1jI61YlLI9A4i6fz1y0JHMuaoZUfRjNnLsYRjZh9a4CeLhLxmLg1
3QIoRk+H9/mNkyyNCJWA4dp3qtSQDjJU/hLYsjq6bQowxjCVghP5fSg/Byjz/vmRoVh8Kp0QgsrA
HapPjToj/4eFeOrNGzui8sRe/HCRwWGHXL4rpa5X+hgYvvJ7ykdACnUNJijXcIgxc81QXBiU1Afe
Zu4NhjmEYsWxKcdFYjp6f4HO0Gy/MT2dnZWVZd7EjuvrnGjzeYoKRygOE9DYTt14Q6I4waJRcxpj
7rVeIMYdy9WtNyHMKilVpM/vI8y8URuczykaNvRZ1lpStKuSL56e2IOGgyR0g7bSW1FOhM5z4Cqj
oEUVXU7b03b2PEsvQVd257w1lv7bEQLUJA8opnjtaw/kCIa+778CE9mgdKOt8ITukJAFWrMGjb51
4s4qbeQNJh/3MouzHoDlOlD+VhxNZXaFVNGMGbFk4CAqu975UD+zNoER6/aLbQZnxCnrE3KzgXSI
HNoI3qTeqbrIqWBxRKdtYJ9CLRubvUaY1W9A7mqluUFYtPEgVPkUYlYmQmhaBVPc/AqjboJaPRJo
2fhrUusn5oNrZmxsTfNUyN4SERIoos3+zxnCTbOKVb2J3ZLYOd1N0y0CSvHYYpRA1JTM+VtJAJgP
imlAgu6a5/wXX4r9b2vquzR1DKFPvfqb1VXzae5nUTuCkHncMPOLewQZgvB73J9Ob0Ey1mZFS7MT
JShOsYJpVU+V/WUVmi8RnC3dql/eIU5IHzmK2h3xg50yWuvzbnY1FsS66Fq+WIeud4oHnglMAEDy
gq5JcSTKx3CQLNQZ3M/+Zqt82ChcbD7jwblpB92BdK7VwUsGHJBrAsRtHtU/LRhP8ks7XiYMpHps
PZq5QpflG4nD+dDH3h+waS87z+bCo02j//+vqbVvYdNunaxw8t783ULLsqnxXAWadoSSsG/1eQpi
TpIyXvNpDHBWiCyzo0la6SOWUnFIVwKxTWPta6st2dGNq9x5xGBs1Y1dC9V+t2rSXi3EqJQo9dKa
bJFyAOCNjJhRxM8wwNsOQnf7PbJrKqqKO+GstrDJbNzPyy4aLj9WPRjKD2XUxqpIoUXFv7iFKoEg
0gfDWm9z0B8ek/XKlBXk+3r4KyQc3N+GvFZ3iZkOadzdYmqx5Ymngd85ayEDrc7/tXyrSwj3ODPC
RYjmFK7zlTlOcn/Yt09wtFAud4fP+rrSWth7VNeaVgveYXeYnL0EWdSXTtjHWsdWO7R/qCP0UsaF
MdO4muV0Pf88O+/Me4rCdl99bsO6URXU+tnR4fXH/GFCIfF7lmVtVBsKLTaCspQ0Ix5DimjVI7e7
QP1xLa9osWd4yVF+vfJ2ZshyjY5NBjyoSsjuuo0vqaJFZW7JO9OvxutmLyujLJqBUlAZp/qoAkoi
4BaajnWWQQudqDhertPttLGDI8sWbQ00oD/uQLN/1OJNYwghREiLVxG2B3X8thYXmPwnEA30b2Vy
1IO/cQUNCD3fIa/8qW0YRJx1wt1MTnTZlojXHUkmVhvu6paP7tEcB064cU9n9OiCCZ2EATxPOO4G
8VQYQ+BI6Taol6H29GAU0m3BqGfBcGM9P35+hSbFVte2JpJy955KHz33u42WR7e91loviqA2kqCR
FWc8qSYCdixzWaA9bPEhU/9IhPgwpz5mbz1JdQhdzbWejCu3GkIO9cCQnRpCPzkduc0yHZcJgMH6
Pgdb9Xfn/Ny6uypoxWnckFeWryZIj6BRPg9ksbebjbZ5VwYqzKc0UmIkzysDN0P0lwhq2rHVzEl2
LAxg16wxqlOGeQJ/nSPcAwV4LN1yL+bdxAFT9wxYesS0BBbniJgL2isVyM6zFV8l4gF2uVC9TMdE
ZEV7qXOn9qLPvHWL42wxTo8UOaFoCGL9Bfg2lluAMw+mEQjREGR524jhJkS8O21yw+SX0W8hTYsz
eifz9Xw5IjI84Ox7KeOF/bpOB13opYFwpG8ehxN0pheHKy0CuTootmBS36lJhClRpHRURSQmX5dc
qn6cgcrkhG9eOkmZPdRnvGDfUObpriW394IJN6/LL8Si8oDALLuOT60jtXMig7tb2tkBeVidGaEl
5yWu+1NYjcHW0fgD4yPQezKXv0LWREDWtZUy8s7KmmehYSJvdj1c9TYo6Hwv550Se3GiD5Sy9n71
kR6oruBVsAuCoEOKFtmpmAVkKGjOLJRs8ukcmPhBwpohMteY8WXNKg1AzBzjvjPeXE9bdFcvWSyY
BwAUP3YoN5D96griyi6mcFVA/MGJJDTgXMBesQYZuScJ6sjOuRFMQEY269UB6JaetxLMi/pDuO4P
a6IaFNbnKinXfCr4y/J2lzQnla1GXhLYZwAS1ceGcdI/wyi0J/OoWwkZsjxS369iNYRi8nU+BizS
DmelRoW0rJvk7CP5gZ44MfHyA46gH6s2uJsjjminPbN6MPJs51pyL+nyx3sJGvZP5NXjoWpkOElM
LZT7WMMVBSPBJw+xEpUrOP0cN8Ej2bnQ1iEOaaakQ3jar2BSh86Va+53sJJ9YAahyGEt6ArVitXs
fNv2xO2laGLyVLOdgVN5uiPf2bNvreauL3M2NQ3pdzC4lD0kpkyOJh/17TeCUX7dazVl6XFz/kH4
ItCBpi819QCGiwwRVarkVgIjS0dbdeKeahsEFRS98GsNN9PQETZ/GZMZKDYdqBIkNuZ/plXyU5PC
hQtntxhIA1uWK5ykmwB1mJ8UySWJShyTKUs/H8b65JxOwdIYNNmWBUw/a9h4Mptwg+9MjNOGuLup
WjixW2rDiqcyvP+gSTxquBzsThLGNDPDUOblfqT8VHZlONq1vZucOrgvfrH4pSfKSyDtULpMPniT
aHpf93cgOiL97peCS+opfvdwmJ59Uh/mQGa6GJjYWX36HNiD7NT2q2lgZajrx2Fwrrxgg2rzeNYa
7qj9O4pL46mmpVvSQ/OgOTHnZA+fceKxk8mi7/fBT8tlSVJdQNvfSeseGP4FJ1x9gZLFwMSHNVUX
9kBBenwKY7qXd92TpMF7cuX7w3SNzN67AYezV+m+qsIz+Ykajuz5pn541IEsum86XaRDdANzRpXK
0gDklwhUET5RzaeHzgvQRV21q/V5+IuNUXU6xMIC5Hn9wmeJ8NjDPF0vtERMJc653HrExBLi8fPs
2CnWVhIyzXZoRq48Qfu+8LugSSInqaYv8sHjse8QgENEm5glQ7SBNtjd6fyik+dqdl5nwAeGEwIL
2Q08tsFL/5JDvq0Mzaa0qwMvH7kH4g4zEb+bEtskuSc9Rr5rYvAnxDhELT3TIYO+cv3wxoOvudUJ
vIqKxYju/wDTZ1EjyzG3B7yUVYHm+Y5gOPC1Gw3Xuo6m5N5kuuYxKFQ2cQFkdzGnbrtUetqKcZ+e
4DpA7f+urt3UvQBTLt7ACnXKr6eu4cIhcWs5qE8bqDdsUTBMFNJkFl4e4rvCFGhnbrPrQQApNdl6
8C3vodhI5zufCWsSHA/Duc+qysXz9LJ9A3bbURSPgn66dxAEu/0YD9VtRDTzGMl1rkOaZ1qBc9dd
MPLN4yODg/yCQhH3TRyfXhZ0FSiJzE35eO+0h+LX8R2nhpWE6r0L1mHSxBeXL+91LfyzHYQuJM7h
yJgbGLwS7B83OWZn5zGh9O1kI1PEm4t1W2ejY/1StRzfR0FaIYctyD7qlVeCaMrwBrBlcRL/U9Y4
k5VhVDRnp/BGnzVXiP7eYF3h98d7g10hOD+nYstZQzkpEO1tNQ/O2fF7VVQ1Qgw1ZyGYVXbltnCz
kzdSG8ah3k10/0Z8kSDhHDBgwdbWCnqWYqEGce2eCoJvsV3ctSawtPPk8DVAGSRx23QZeenmhL0g
Z0+zlstVYhbrPdVigp8=
`protect end_protected
