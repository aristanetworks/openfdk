--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
hCOiIL5FfsUfmRLuQV0BqlnO6zGTJ61eu8JQrcoDBfOe3zMjRTpvq4n0ESSQo38jIl5uOufAWYlz
Me9J5D+ycfai8mhzuFEUd2rQ4SAvTh7UcbbgiN79MwA/xoKgFxxXMuTnVJv2Oeq8rDkgw/03nLDv
uoXpQCEYezKz1fWaFXds/iQr3R+Hfn/B33jJumPbtsIVTaLE2NtQddiWS9pEqSt53sNYMIk/4MgC
lVOJX4K2R6dBaWGGPZQ0mY9NdF1C1M8ThLJrN+5CuoMV2j1yn/54wM4nXBS2hnC3mr1AHOdegtOO
IgZae9M+RIhT/iRLDrPhGs531HgRV6QLSdg0OA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="K66spO5ViXvzAKFB5ZJIYmJ2U40Yz2inFWzY8lRohh8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
L7u43RmFcEeFqH7TPjeH87Euoi+PP8OD2cH95XZ5enQFgf5yonWeysIrFp8TnaNJBacvzNf1cuSp
kQ4GYAthLK8aov/GLdlAR53Nf7cOSRs7QJc5PSpYsUB5GY/+qTO383UcVkO6DQN/MUPqqp3V6MC6
DWF2DL9iySiciUl98cJtb2+Qntj8S84PI9maQ5j/xe3voBKwjyeX6GUNL2v/GJCSF9imScamtRJt
NK4+y7E9OHi6Es2BujM4UOO2Bc3aBPBV/ECpMJsFBuJwiiFJE5xP5F9qPR4LiJNRP/t0KRwNNjNm
JAroDu0MVYN/6Vo8bwePDAWCWarLTVhrePKfLw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="/P1Y5Sp9UZ8EHicMiVJtrOuzzDpg2w3GFC9XdDY2a78="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2080)
`protect data_block
HGUrggQ7jPOi1B8pV+2A1t0Ngkbg1jynF0R6rMF2okleRUo3OL8EOvCKrxFdkAZto8nGS4e3uOxf
2bAtV7/HhBTMWFrtCje1hbU13I+2YmZPKltZwuso1oE7QO2pKr+uxMY0bOKzvRgCaq/bAVbldRbe
C4Cmo1dhE0epJtrcM/g7leO/H1lQI4YrSWYRU264FOITY6VICsvap+UWV3zLJe4gxAcFqqKVe2XB
IDCLxrugzAuuH1furI3tgsOvNir/o8H7oRi9hvAP1JbAh0WNjNOL1rsZWrF2pFdKNm2nOool/hu9
sV2FHNJuwR81B/TOJoZsxr/uOPgPvkA8qb5x9lYY28VPKsUm6Aqg+R4y6KGSDTFApBNFj/ipN851
N6Q00Vbz7vCUj+x9/45dcz4yCEKdSdK90+xKDDlxkxCmCEDsDv+RroyYTLgErDmTbowwvAnVqjxZ
fDqTWL1/nk1CIqApcWdCWE+tILX3bLPrWpJqMjF0ryhlNcdsQEMg99o51VTnfuR8WIx1MBrO1KOd
iM6TAdWSO76o5lAH5DFnzz2A9FC6rHW6AKdpp/02QoHiwzPQP2C/r2QGtxTVDjwr6gGFPg+INwTs
GXxLcf99mYuYpw+A1dGt1dmjsIWYJ9zzJNbNk+HrDZdTo2FeFGjZJLbCYdX+9BA4SBFYsGV6lz+K
iIEJEzNaYJszgD8NlHqVmeH73+WJgcIvI1adEN/V2N325IdFsxwPyeLew6wRPSsfdvLs+/QvKDqa
LuSKyB8JEbNV406bA1DTHZzzUqGVlyVAp1iQRPLo+56ArUN0AyhpGKsObmpRERysCnD+r5c9Zh+r
Ee4UCmLR84mrINwOipyYbnKja9GeUzQ9BqcBk9UP6+43LkxzFguigIycGQRe0weuDfFmK3wKwAmW
CpnwJlGIvcyASp+6tA7StzxiG9peipKAUKwDfsTdyOBjJHQYpgOyYdEOe+coHW0yw73w+QUzK4dJ
g/T9BlTdpf+XUG527CWs1JpkxpBT6zEtDCWPcAi0SlO1/mSWo8+9KZzNb4Uk1aEy4gH151Q5wL/V
VUpHijpgMlpIkqYZflWukw1XjjJMcuPnGRQn4YBb2CGT4J9lJpBurUe/nJDof+9cXq4cvk0ZWDjx
LOigbqY7bDwf59XF0GLAcocxsHpthRaqAXY+HQCET9yibkTRdJ2FClSLG5vX6xgMoZZYnXfsL8Zm
gC2gxvrSgDlTz0//DSRFBQmkgrAfF2LQtk3Tg4DRoT4lvjjONWXJLnPiAwxAk3i9c0dB/J2FCo5+
lfi7Ce3FGeJ+Y8uyyCAztbrtIu2ZiEIPE3qXeed1YK62ij9S9ScjbW2TSg1gbg7/a1GMYgAlk7N6
ZdPX3YU0IeJiJyIbOVvADLpBwPP1bk0O0zub2rDzH0UYZDpqD+uFBcYsq6sRggUCZtZI2VvC96no
hGmaUA3MS+/7qjod0OyGbjol6SaNviGsme9i0MhL0e/0RowBKFgQ+H3la+xO+KBuU1NJvq3tQ/ET
vFmzDrVuEq+bdFyY/HYXZ+GtGj3l34SauzCNQvvesiBI37j3fQ7t5Ex8rg/BeyEnfAl0ohpIIBPi
cL7ORMlt0xu1BxomQZwrdlUs0ZVQW1CE9A+CHpiBw21uF3Amp+RbotrG87fL/Eag3AngO459Z7wN
H+Gx0gXy6qqaswpnlRkgGvx/9719AwB3vrv2szul2XUtHHBMq/bGG0WMxH5jNotwFJakeFqLXqWb
3hyfsaIH6ttqdCXPomhcNXvF+SCFXMwqy0Tn2ezvw0e6BYtvLQWVLoSKDupr5tjvym16ipgJZ1y+
/y6pYV83pGLh4G/JI6P6Qm2qCAq4BANVGXXaDhh/uoRbwSVUZnX47/pqQHn31vYeBaXMKPbDZoyZ
fDd0WPNiKJ9h/mEDVtZ9+ESalAEdmTCgXYVSX1zaNlIIdPtq/wxnu7wsRzcYqRlHjIjlY9crii6a
/VXsn9KffJ4KRhsXiZc2t75HGr/ekZek5FpmDT5+cEUPhFpzMwrOPZIr5cmEKdoxKcnHP8H79YLd
q6d2Dyupbx2UZ7pPgXdhp/nQRnjUb759T1Qc9vXEfln4+u3StGqf8JlLOLuGRnKa098yvj+oRTDO
dx6biuZrN79/uwzn9yov9qnvcwvIWJzXu8ot2YI2osqYtUYW3lK/Pi4c+pKauw6MBIqNCnUw+/Xy
3mB+7FSh0M5lZWqyH/hx4gaEXOR+46YANwvfC9n/eOXHKo3LIxj+AUPXIgRg2AHssJMSBlsM4UeX
hc/vqcxEBkp8AICYYSpXtn3ILZXakRosww4H8qzsKjMOdz6UV8aKh0UA1GeSEwW0Zhgd7XD+Z3eH
H+tmNjuPOKf66U75in8Gj8uhC2H6TVxTcP4NXiJ3XtQ9xd2bpX9g9eUPY2M1nvNGF0rOFROJhHZX
81cl5oiC5Ifd1IVP3oL0DCs1DylpimM4TmdASuuUKPq+mQ2jek36rx1oE8gkkNJznq8mBawHH1AB
bnxeTV+qNatq5VdtGlZFdMG9vJJmXewIjvF4ymKYuNTS/Q6H+UT12M/pTQBNxbczaOBVsIGTXsal
bMgHLJ91RRqjO3e4yx5OdSN4rwCIkaZJ7RatcmUcw7rJCbhoIOIO1KrPZHDntH4VpgpkuBhgvpRr
sxIdA0Fpzm0q10UGCU2LS4MtL9H0h/87Jjz2fc4khynmdjeNAjIVDRyM+lVssK2jAtL29cFbunHR
GFHMFvNlh7tkgeRRNi8u5A1rsePzwNFhRoqjCg==
`protect end_protected
