--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
RqQIhv7Dj0EwtHNNurEEOcC+MqbGsPanOdzT0DqIQGyXRNDEGR9pxSFfSiYA1aurfbg07tF+pytL
hXnca3Aq8XrbXkjPS/oiMVagiwkE6UPye2hCoyWyXJW/ofnKFKk29Mduv8Tpcft0U9NIyiPhspEi
rJMjs8SAnHcrYm8qeY5fSCz1aNnWyxoWsMWJbdwEvuXZXTTcDK7/Kc3aFPTqJ6Xqd2lrLmCm/bxJ
+HqV1qHvEyx3iG+rlmtq/fzUiXMimb3N5WWH6pApqp7+nkdDXWc7b10c6J+iQD1b1E2yBFEMGZrR
IsmHWXV92upsIIahZDSvY+TSc2KropD1lQVzJg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="zLHaBgdewui3j3QVqhgPeda5z5uCZUz14XrCb+FdlPQ="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
l+hiSvbPwFHD+3qxuxddK0id+NUp/ccaQ7ym34zK5mr0VjqVDm3PutZk8+PjMj679fslNZlKpjtR
z1m4+nKLW/a9BaZSs3bl0IzrjD2cQP/2+ar4B6jnOrKyXFYpkTb0uoaXnprKhhr7480EJUK4x7U+
quFfsCKBBjPGVRI5XyykbKuHQN3Y3Opdl59mBS/lBZp/KhM49Atm089jGFFEPMEXE+0TUC2mza+8
bwdW400rIPiKwgBXW8rLwytflljpJyPatrV+c3t0iTLGuoaut4Hped28uTnizRzslAR9AcQsceQm
+ESglvUiHhl6ubat1Pg+d5GZCZowcE7eVqBo3Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="bctXnDIL3Lgg81YzOE1Z/mnb4pagytgqPCDVACCc7p4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4672)
`protect data_block
xfTkN9HRfobKHvJ+Y8RGjKJPM19AZKJ+FHLtXtFTpCpYRHnM6Vz9lsiJciSzoRN6sJUwnIWw+XdZ
8bpZ6S2L7euP0hiNfmWgC5++wBo/q5Umv/Y+EwUlzfoSfDjTuWAgMsfgG5glgkYi0skQxbyI6IJ3
KkrceYCY9G6xiQDJHcU0VQBL8Fr+zeEp7VuqcfAvzfhtjcp4apJ+tRWp/aa8Bh7oqnQQq/0pQueZ
OXsEFaaxnp1nuxc6gw+8NjZUu0W4VbSVTdRg5Y+jyDfJT04Gp5LqyLv/gF+5ec8OvGNGO0Pmdnul
QP6wp7qYAv9uvVAg9J+B1fPDy2ObmzfrUJxd8Di+Wz1g3NkcePdstJwNwI5/r9sofcD0blIwW3NS
rLqYNi/5//vx3uW6VUnM99AZqykRV/IX0p6Ynh7MnVxSyoy8Yo2c1DUhqPoCUJfmC0s7/8sBQ9BW
j+hoPUHguijDiH9GCG3/vmgtp11qiZdRIIQDAmGCF8gke2EGBaFK47mLDszqN41rOjf1vomiUiFw
aMzcfxT0rob5NAOA8mjsOpCyp4HBYYCb5wY7SahSchYw6GZ45jPWghY7oIxy+2GB/AVUL8bf7L2m
PNRIuT1STJM8MqNPiQCfCuuAJr4tOLtUV0yhhQZba5VZmzk+yBiEqLP0qmeOS2K5JqV8V5IKZVYj
AVskvO5T/r1pQhkWhH4Elq0Gu/mM/Em6lPVI7bil2sheUuB6CuXGQL/L0lmysqgz/htR3Rq6mB4I
Oa/+7aKSbhsRCsF1MIgL9dZo0pEtJsjyQ311b/XCFCJxZNWu/6/olTygkgqLYpS4D9cooNTpl0Q6
niEW5lUbPgK08isNKLstN/Ns2nF6YG5x3aChVKv+KkDAdXYKAu4vwnll6ZDLYVDo5zL1UAUIPP3t
RWLo5VxAQGFCX74oIC3AsI5VC+WFqw67M3QOeRCSLSHBa3xrkrZQ/dTKEwf/CYsPy5Ot7Kpslvni
5R/oXRtriNGEEYs87JzCFVmycBNo6nRhxboW0i5Ryph8XMIoufhGnzkVI98oTU4aMrFUUMFrr7Uf
io8ztpedKFYSJQfXLux/5j2kzhlpidoLMnMoIYp+s2CMf3SBw4Y8sXWOUGudekmGfv/QqZIJopUh
RkpNZEk4uhLFO1z2hPal5dGjP94VgEoR5Mo/nGfdht1d6rBQHdr1GaOnYv9R1K8KPbFEI4Omjz5n
P3weolnoYgPb7LpejGTFgJ+itplTPo82/OjW0pEsz0ZPxx9rp8JkFOqCPMmA0txFLeC7Z2MmwjDI
VrlGE0SzbaZwjG1IAvw19FlOCsZPFjI3qaLizdWj/nyBiOxEsqxju0uoT4wzhoiE5+oLaVtvw3Sr
C590LQarUISIaek+FbT6yvyE3ATjoqdjjGBlY7wlflmBLdC8CiYc2Uk4CFBfN3kG0i+2A6RLRExN
HraFaA3+TNEA/UjYM7FGz0ayur+t8Iv3BCIe6mBwx3j6GM/hOsE5KB3Ndy6sBrrLiN6aeTp5rGuJ
TBBG8sOxGFZ2zaW/V2fBJR60ZC23VoRR9G1HJReDcbRsXJMLOonNI+s3KRk/MdddHLrmFoRwxkrR
vUVZh9iMGz0YJ8TiRWfHZD63nmSKc5sBQbCMw3vxiFEnYRuRSS9iZzOtMzq/QBo8lb6fLD2HtbLP
u60iXUdwDOooUe9A220S91CHDe5d4wCDMWAszlwnWmTj6ooKH6V6MVd3wr3fnkKdfzyBwwGDi2iV
DlTraPxze9EJsZDLUsbYJY/c1KdwFXogwNP6hbz+nDSGqmWv8jC/Pr0zTkiZH/ZoIV22Ultj6Mq9
BaYpOo7sb1pRcfhejJ43UgXhZL38h6byFRJ6rF1K1jmXxgegU6mEX6uPt7Yg1ZhxgS2aVNC8w1nn
qnB98EXrt5CUudvlxZeLmsosu4yLQCUTHbTyLvuhX75ZuaUTIxHowOVxt7bIakMK/gB1uIPQHRzX
cYt00FilgfPdbaGzVbBebRVUwtfCae6TV9alT4Pj1t8yeOKgH8uUSBnwy70cRsoh2CkTKIbqXtgT
BlWsS8kUKGcDXu4PZNK0g6lbdujmWCsBXo/yqCkDgWehm3kJ8W0PNzIor+0Y5q3CfJxpw2XXSkbs
oYbDdCZHE9cABEvYmNWt46jLfbBA9abMP0yqCyiZ9p1zaNienz9JLGpaCL2YSn5wKV98W7PVxmoH
C7rBn+EcMeT1ULFKPqNZ7LnleEH5e4BBTBz5KiWZh4sgiMnVVcOGseBmGRHO8QJ7+fuX5tPwVL6G
fPejrbGVLnjBFaWTM3kAqfxtwPHsYijbLsmJP0dvutSJXyvXqvBtWAVLM8ZoOYYvXIt9UgJTsb5k
lEJJxDFWA4qHlg+q9IC8v2ukCORqf2kkw7I0tH4q07IYFvhK0u84JsUtWoES7W1cUa/Ojbh9qfyV
a/P7GMA3ZKHx+QUYbYUEvxW7jW2bz+5FW26hPd/bCXLtkydTroY7UVdFi+6bEeyd1x8nbuR/42Hp
oivOyOzUFwSXdMJKEcK7/iju6qzqOIqFjarNPyEjoMlyQ1QTZGHQuk42W5yJBlqh77W9h2irS7rM
w3wN7Nn+Mh3uSZkJDGDl6Sa0pO0Rh7AnYuB6jty+EopXTLBEaFx2tbq4bu2j8QcvkegfqCecw4b1
d46T53ecOcZcHzNOFb9vF6I9bDJoXGs7uwfL0rQdNXeaTvQdPoqABBcYatT+Ur4DFNxypGTjPH93
ULLLxkhIJVUHVhUF1lTBCjDwVNVJRwrugtvX+xwURPlHfYR2R/VARswcWMf5miSzQoXda6nQljva
rJ3uWD3i0zyB5MKpNsmm/0+J8HlhMmhXY14N+GPrRxSgl5WcwV4NCW6/JQzkTj1MM+rmqZ1vy5n/
GV+0CEDd/p2bJF1HG/2Dtgrw5nkuglI7S5EIk9C7wEDRrrhnLH5jw4f/2GUDm+qNgbHNG1AjHZFn
Mlj7FUQPyO6eoz80XwcpMPG0y56K7KNvryC0RVzDj1gNicrceOVld6b16kbO6pwikqnWndjOHYK9
LIUUhu6zJlR4rqElyyERm0h6DpQA9KRJQBgfQUkk7rkHMaq+Eb3fTV8xX/CnI80JrVSLS5DeCRFe
z9y8lk68SEE/AZgAplvg5ELX7SUWztSegYsYVTDiSOiV4Z+AvCUHADz0kFgEVUT6M5XNQK9R4Y/B
1PxLg5Z90ushzuQv9U/8v3gwT7kb+J2JmPFhktbzsGe5oarIuOH+qIe405u69Mt1vdE2/c/v6ouL
wJPYX1OU68DooTa/jn3k4vRrOFda6EFzVsK81tYT4U9Wd7oY/jY3mwtztYAciwYH1DQY3BSYUtc9
71rG1sXIcaiV+mTlj2Fi4lOY/nRU6o8lHH1dZdSE5nLrVtShDoroh649imfSG8e3F04AQvt7Se2B
EC/DWG57++uBMf2gYNfDjJXu3GnoSNoVkVhz9Wa+Um36wVFOuUSqZHmYb4421C/bkbH/kUvGbJ7u
WOUs0ed++AWVH+tGOmIMpKtWGcJOoX7QyvIUy/oyTe85Azzjh1diHjmq8vDKwmz8a+2C/qdl9oWF
4P37cTMOX4q3jZ/c2Yql5nezouu+WQiZdc/Bv4uzPOKDaRx5zFr78yqpmL4H6EHHimLrGBG14RIk
QWPSY9x0+Y4r5reVpbpk2icOIDvts9rWxgEK/zycqWAG5+pKx0n+eUXao+GeJ5GS4hcWJ2xYtGMk
HPPWcNpLk9aFeQOdmcnPWj5AFJj3RM+2QHPa6oUloogWaYvYGwmdjImWjrl+J7UxajPmgMEtaLUp
rfpFESrpbI8/LD4fCSq2CzT9tio9GsMAe7R/gqBR1yqF/e5qL4t10AjZ++J+UuYzDdaWsrrmVy9t
5pbgy+Fp6reThizOjBS+KpAxI79+zu4YJNHehFgyp8eB63w3LO7YUIv9LCQG9/lMf7HHDGKbdOnu
fLb+FQNP0KF8YR3nwgKFYBFidwzfM4X03SvABG/REs3/SFuoBr2EQ4GbaZqxwbaQRWJJv6xUF+rH
K472UucZ3H/5xiypbz0bBtTlHx29qw6ekVPLPh5QLT8Dcdtay5Mt9RJh1XcyG4mHxo5dYALm6cDW
/275kVoXFFxcAGJEN54dNQtqcIxI1L1A0V3NRpTDqKDyQAJGUtkygSOYkvYt8B0oiCvCxXslaf28
6AQLaxA6mpdRgbmIf0Z97qKHDgjBMaeBkBfuW6VyqFQ/8abyqT2FEofCymnf1xTcIoRhziGmR+DT
SrTbP/gswLsgWZFR2aPsxW2R6LxNKVNhqb4GzaYoAQurhb7jbn+nVXFniqp9nbV8/KevPBKnQiNm
c/daHoBLQSL3qeV/RFD0nMYbDfRtZDBRLmu+AxKmdabpWIcvhvqh8izmcxCaTuPJEJZtU0xUM/5p
sqpqDdW6M9H54UmY4xIMiYbGmmxU5QdVPnsTk+b9y180GnHHD+CXW+s1G0ZoyOejrH37Oz8RnYMn
4fb2V27lH/5Q+WAsLExVCwX59F1NMNUMb1OnKXxRQmqkA4ZLT4n2NojF96WND+cnviZn5s+NQs/8
0FJ41Egz9lF2rXMAJ2yJxBm1nKLMzuKvdd74ca68UJqoVKMZY+p/QKYOakFuQ1qD6DEcOGTvCg/l
jUtjWLJA/M6g/+sv2lhFodk+/JhF705H+PUq1SzmXcfUSQev7pPLR4MdGJempXCs6GC4i5Imp9MR
2SmuaxyiS9xj0PV6x0IpdNO0C8WO+4+YwTMW8lEPRKzWH8Tyb8NtDj+Z49lMSdByBsNJRVyKMI2/
d0BtEMOer2yrrLzjVAzrCRa39uNBZzPceRUlaKb4YXBDIXqu/PLWYMq0wloE+crIQuzy1l17N54w
8imRMoxewLNg52jPtr5r+EHSAgIEfisF9BomTf4+QatXTrgQOca5zURB6XhsKprMUOyr0llu2V3Z
PshDzxblny6e0ne7qLdqUitWr/XpsIueSE4yZmBnmJ3B9p+F3LabGvMzEpaEWUhMhZJyXdv5sJtM
y+oFQbWvt56qEjC18yV8RDz68zvfDC7TElCWwmWxVCA/12s09ZcPVhx3XnzabdNB0VxVbWRV0o/l
JZCuwRMueynR1hePU/4qmlMy3tzeFeKQ06ZZHhet//qx7I78phUP69Dy9lzIumhJ20EGM/L6DUKv
MH8TeVPKN761AB65t2nRktl0Q8uN/1nCEvSPM8kqRW1eDKthNf1JWTlasnwzRli1d+CL0GfkRD22
n026mVtOhpoY4A3oh7sZITjuUGEGHt9qPyqtzcdGSwLQxPVfZQ0tQmyTVwO0YjAuwEMU3WfO+5oq
l7gbsmqoE6eBZYOq83Qag7fSO9eWnbEKF3mT6+B04dh7TYmTa39rBAo0vDSGiwdAbQHLo/ojLaBv
v5QbXCwMuKGm8I2GzkSTF1SEXbcdd/6s/0/UMV8GSjy/1AifLO+MNxsQBdPVW1UhJYAdo78HfzAB
2H68G9MNaHj4IGWDSV7n8Zt81bBS1FioY+ezQyGkN502NrMa8434oI9JhP3AOC1bDsJ0ijsZj9HG
zBGET55gCAkQlb7xSBuNq0Z9wp4AUyL/ICNIbd+wBfa2jtKwvWBNqtBZfqXvgSPwXzWKiUJGKPb1
TUO8UT9j/kJCjZG065FCQazShmR/ZiNIMve0ZlujzOdjupTfHq3vGqBWN8lh07tMxT+9STNXFDy4
i73tGEEMwPmF4tJ21E6XyfMwYZeT4EWVroOJxdx+J0IkWUFy0pITzrbMR5Vy2v0tFbgFKt1wzz3u
c6Xg5VkYt1gTDcU6D8Qd4M0x02ZE9RiP9nQedIV1fn/jg1IpwAu5Vp1NbEbpFUxqpL0YQHGDPZBP
rb8ukz6kpcpOHhHrauKvWf9LrBQMJn04VeizOlra/msDNDu6oNkYYPlTVxbhMMCHld8QnMcbFbGw
DpS3sFJtnIMEBNePnibOHsF43HlNjCf4o51q5tSl68krdWGt3fNq67iTTNhfWc6q+eZzo/7OKdkw
Ixevfu7Zgtr9634jGLTuONTojVrImnkspgNQ495yKIk6YrpIhPW9LoMfwY3TvMvn4FhV0O0j4cgj
+ZlNAm7ZnYB1GcMfdQmPUh8f6FtiE3cJWnergtMlKHE5XbrRAXQZRVTsQIUJuNLbiRlhbVnScDpP
rqxAuT4Pew+MSRME+bFaQP7LQScAD+P06FwcoQVWwbLyfzrtX0I41ct0d+rm+T8/6c05wwRvBA==
`protect end_protected
