--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
CV9poKgcOZsZxoUzwW8kGLL9OJlqsrQ+4ES+E6iLp2ChpjCqFDBTdCgwnAng62JpALGohyMYxdqi
KLmX6nkMg3RLdz5fW8vquM3wENNmNw5VfPGpr7qJ5URc2yr0u44MpkSMX5NIF8K4+WCLp1kyoufB
ZjwHlTz8gE77BFLfzS51JoXidVvj2c2hc/bBQGnk+Xqd1OaaIE5rV6c3bl/iqqkLgd7RRtgQFHr2
wDXIMsA3itrwcYroH7sYknbkHzNcPq9bZKN2QywUGCBPdMIiWlu+cBjdAuYg6MEL9wCLfW3NQMWS
GRHAFqrQlfIqjdajurA+HgDZH8qTBvhwKeyXew==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Bwo5KyJMBND0Mqlv04Y+H7F26eKvF08JIPm5VTQOaKQ="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
TPtmJGVy4ETuR7JWKk6zuTQqL/t4TXruSgDaS6ZXWVpqTNX/Qi2e+A4d/1a2ZraHSy6+dqLo6TGu
wPDcYtPKVa5vFcDlJaThWUqriwkYfrZ6KF2+WLO7Cph/fgPUE9R2GoMGD4DBvFj5cUqhEo7O2BHX
tyZ1ocjfNefzQWaClqSM8JLwxugc6F5rtuksPJZP86kYxOEbMgYcQjQf2PzA+3ezLr9HQ8yissyK
iGyKMKb5SL/nrRijbki00zKRzCNRYTl7QCbGcgky0xdyyL8QqYyHfAAJ1sCmxT/VmWUy5HTFuiQn
YH+DtuyJsvLQlu1nsnBsIK4gZUXGmPptXgQjaQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="JeHTTn0G0w5YlDGCf7dFn7jN2fhiygva9X2tbi4TjbY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10448)
`protect data_block
x+/AFxSoFgMvzxIdbQg5Vqbf4sY2q4kQmq6HnVXqcOhDANEoKodPWMjHwkZVsbukjFn5+OXRsL1y
fjoxgYf+xOXeLtz3XXnzcy4PRJhAI9v7lS+TWxTp4Yy6szW/t+ruG8vtMPUn9p0td7pXfq/nyS/A
kbddXOMltUh/isOBXjk0nBO3Of60Tdv7sKFscf1jLycCLpqKYLwKc6RfLdEr1r0J9uFfdzsdemGj
x8RWsoiK1VjVEUseQLQoKnhmg9fy1uIpjlDywQgujIKKsDe4eRnC6Ba5myAQ2poVNrVKcLtHXsZ4
Sll7t8tUITTYP6nNXkGpPdgiQ68V4riyWaxQI45j2Ii6MTWaxMlVna4HPedsoD3Hgm6jGtUnBqP5
hoPmHZtZ86ieJXbb0V1hvish3VfxMyfo7ynFVpg7yF5pB/oRadavwhTAu6iZFeLme8zof6HoS4+4
+ls9mXBhed0IiXt1N2Anu7s5AxIqmDLT72mXEs6KobT/eaIIBMRizwjV1xD0shxtH6SLnsrLe/2L
DI+kd/cNDqrwhMJlbRVfKh+Il2hghQiRD9jslrojoJrdnzgt/n1jzfj+FNl692+0Hvrmw7wWFC7a
Ra92KapEBMr6Ma1IghQryh/rCIUN0DlBpvRLzwu3b2OL9rRc5Z0VFpInv5glc1fPC5EfC0LJ2vF8
GFiTBat5/M3grbtDdoDkCGTmALcnbGgChHSxm9jbGXfN4R0g7P6BFVk+aq0R3ROB0EdfV1uQ+rue
Ox96glnzfyR0hyyYq/cer+XIsVhnjD3h9S3+x5Fs3nLhgAQyPVqejqEgNwgTPC3FEDxUUx3CNAty
seZmRJRV4ibaYzS0rX0lUIt21byoIgDzZsKNGA2BVdCKkOCS1yRM2YUZ8GzzWql8+E2mOCUj7T+n
PLL52kvinDIXufXXSjFLlx3h0LHp90jhFys+bLPY8CIyRtv/yX5pZwrYD+Nm3WKEB1D+OHzaaErG
a57eRpM6wT7pnpyhEYIFaKRp32jtfI3U22uOFXiMjUP2I1OBqquIIgoe5XkmVYho+VBZgUwsH0bD
ATFDdI583+OE/2QT09SVCd7H0pAJSpaYbZR+bAW+6UDL6XmOP3YcBZRqrX04AP/+l/PKL2bLK2R3
338K/DJvxfM86o2ACXKCiSpeLzyq9vFTCZLo15IniXKoCeIs2xXxLG47I/8GdHVQKQC3yaCDfHwy
oiWGeUfBDtqXJU6VJbHpBMZUQVDddXFt/JIerXJrfz1z4TYIYCF0DgDc+mpyo2or+cX9iN3LRmPc
p7DPfdRKXH3pymSKcP0McjQ4dC0zh5oi33Pshm1MfJTTQAA4nvA/5R9Sga1P4x4A5c3o1j9Uv89H
dlsMLypxEg3O5k9UNSpZjVERYBFQEWvIF6rYlNIk5vlxcOF3dEPSvtIUAagTwG+YE+igqsOQi2MO
vIhqxNJcw9vF7OqHP08+o01yZk0w4qVdGNZJ3mWBc8mEnr8ijuNFsJxPXNpeAqg4YVFTJhsJOq5q
EF2UFRamXNNgqJJj0FIYYbcMB7duh/yOMs1d7Shy590VW45t7jfspCY2opqPQOl5TIeeH/a7BZQy
3cxe4GcChEmiIsV8eZgxM0WLpdXVBFnfrjMsrt38ONIze3vwTwn1ikVRhPNiITUPrdcsUd+qixUd
jVwmgIkDieYBJvWnRKNiBkHg5hn+7oN+5Gx6AyKYYGupH0LkyuXfZslJd7kCUoygoz9D6j1JieQ9
Xd+Z2V68UTb1g0InUmkqw7KdZ4QZxMp5gAqIT2GpXPKJwX3/29FhIcefCbzyjWZpl7pzsN8IMYbn
UVF7V5ViQvXMY1nJRos9I9U7nfDVubrWHt9IoOxbfmq0M1V7vUvFXQbTzPIpewpEcBEbchO3yH4V
yQAlrPtucyQnue7b8SOm515q0sMMKDsSEKOmeaVRMxVeYbXXbOtBAAoCdTbVAr3T7X8WNMzEBmrr
q55sIOa1IRv4mzBc9yxGuq3g8KJfV6dKoPU4FqFL7KdgtlNJpY8kTVEIXN2VF9dAq3sa7hDe5Dtm
otS5edIjqMiF5tDTAeAz1FhK/V31gFkBWQwFQvp9qF3WWUjv/gcBUulHG76b9mP8nf2HsNllztQk
oxojGCA4mK2/Enwblxnp/2mHbNPYlzDcQ2qr7fBQlC9KkLHbeQ8XCEzytuGynInjmT8rRqR0DiyD
qBp0bpbBhUovKF/zr+D2tHN4Fr0ouxLch/UcPsi8+kfd96znSV6Zi9M7/XPlZ84pRUV9zUmDsBYj
OhwQQnJccquNekqI/3/jY+GnFLHBXNHh3edwpzavehLBqeCCE6ueqoE+Ifgp7prANQFyo/KOXEih
pbOY59b+TdlUZRXT+wZBpWfrRTWGbDiSGy7lkCBiP3q9ryq6NJcOaPfH/Uu0SHw0f2whXjWUvBqo
7UtM0kFAVblbPbGopDzkYt3D6SH8lcf3y7IW2YNEXyb4Rd66Ib611NK6a2P/x80/spQ64AKUQC56
4/fBqNMSIXVf+szSDS3RZmpm03yikNP/+Gbmy9JEsPjksfwaQACijBvxA6JFuD/vB1W4IvdqLziF
Wmy/MtBYG0zIEbywlecBtHlawTzbwccQ3gFMwAd+ZUG4YhpNysLLeBX0k+BE2EfTdJLzrzq+a7gM
ld0VuGK7/JDFAACuwygL2oG0ihT4fEluC78/MSr0uv3GQt6WSwxftFvpqWi8tAyESbRwlfidGsfz
3fVwKJy5xg+v483lEVXNykye4hQyWUpmliCsOULZdGRpHuSPWnOByZlxhQR2TjxhavdcORchPYZ3
bZbPq4nj3Y8Je+VJsgKtHF5OlsxrBopnWUAdi2qCd6G31HBSnVHrlbWwcWLBwgTCv7SgQcG46tSW
INZOBaS79kgefK75JNZvmjeZcNbX3BDQx7zvEr+WFRn6XbCsom0ANRM63A/6PqpfhdgvN3NdCkr9
oWUB4VBAtjQM6fJV3uBS+xyDjRttLb9YAwW1lZ4SISDQwZ+KAkdW/gCDA69yBeoxIgqrgs4ZB8V0
ZNhxkIfARnQtmT2BfQT+aZS33uI43F3BOMifrQd/YDB6YSWgTiGol9jQPyBFUFUjmIT73+tlWWHl
MkMlsyh8dGg/YMz8rroKwU8AQy9ZioZpKiekv2vYQcz/5EOcp1fyQs0bEtq8/gYo7OcgpZl2ze8u
o7QSCbkO0OCjnGgn2c0MDAhIS0YfmHZDZAvR3goH5txwSSO1J7EPmwmKhoUtMQszRwk20Z6EmdVD
XVZwFb2K01Hh0cj8oCQ6OyJl+yKCSHpfShcbJ1n04ryuaY1vJt5nD6Z0XhRK4fo+qC+mzdvARgQa
wozFBRxNSbY9Gs8Z4bWhbJ5scgwpPFJ/MbcFaCnCBGaIpWhpMqGB0lIfxi3QXJO0AVRLzUoPmO5I
s2lAVWGqmJqeenvl9fCa5CiMptk13vI0xh3KXTx487B1xEA5EmtBWQTXkdE4bdl8a3okcyDUVYev
4ceeR/99rp2+HIyLPzrMpB1OeK8NuJ4fuGN0LEzgQHri+2bL687MQqa8yR7zsahzBnbsuyvh1zTp
6TBk6FkG/mNqGYWeiG5o4NGNbw7EbRvg35M9Jw1rF7oke2trrX7eGJUI8PvGKpdtNiKIpOqRQAs5
1R2Og0ffJ5ydoAj8eJUEP+S4ZeVY3fxVflPfIGdyEtUHT3gY9sMRWc52bptr4walQ3cUj7w8LNcX
ByPcWtxSx1qIGFopI9UtU2sJSiG/0KGeIVBedWUtzVZL31hkG39Sjx+1671SNxtsSJV6cWsHP/OI
J/PQbA00L1gwbXA/CVXTFx471a3zcGvHkxddPTVLUyRdS0ybYNUoGkpipOpbVh0Cu1hbDbWkZHLM
2FLMM4v36Kz4lYITYy0rk0Ju6VIL48YPdxTlyFCYv0hNDIbDkRTHYCSxSmtWGGFrmYBzclOO9fKh
eN9XPCqf5s07adpaqeCK0xxaCBkagWcTqD2BeqOtidpDuyff4187nhor26pPZ7gwRiIQ2DRPGdSV
ukYVqPgfiqsAWSxKDBtNcUN0pNvAWQn56Rk0mlgkDpfPeM5KOHN9cAfOvXvEBtA/mGxgVRBr0wz9
UbFla/dMXqYEMAAw+SHuVLU1IramyM6/57jNPqxCdrsXb3Iw8t9pnY5fd87RTS6h1hy64uXKOyEM
1szoKgdquGkXsa43yQa28hbbACKYKqmmNk/Cw2AtxE9y3xrl5Gcf9wA/3bMMKo7WAN6KNLAifLEq
WFRUqaK52h6bLIa3F5TCC8F9kf+a84/3uSlseOMW11e6Jjk13g90clLCvhQ20nftnvBHYunlCJPG
QyrEHkmKXIdefKexSZ8FKlMTDRawkIueqRdL2lFkqIeFHwDf7pvcDSDH1DO5rdzhDqjcaJXm+gNv
PflbZUHt4cLIHOqHhPTEq54HaMed94v3UUdHefhgQGG+u+XGUd+VFA/SN8T3LaIgMs/BNsAnYTY5
Xh2sBwwmwLBMLIc31Z1o8m5bhQXCjodM0v/JZV/DkJBPQ9zdRnYM5T75v1fWuEYzGDe3bhumgfqS
SA+MoHRjWE39zzh0O5LE74JSnWxnh4BskyimkAhy7p8OwyCqbSJPYn2TlCnAVJnIZgLc6BCnbcZM
voTbXt4l1E2TlL7kmx+kU4qNQhqXfY53KTLHXbHnrs204O18P2Cp3pkWGllGTCBJmib3i+zoKPbM
NRW6wsGDgvxWPE2lvt7wJtnUNabRwFx3TpXquuntTDoxPVG5IO0p4hpNK4nWlfvmqMTNd7icXCCJ
MaHDYA1qumDfS2hmeuBu1aZNAMVFX1kmnR1Jy+ANVIDJ70kRPGfh3qO5XondekEJ61Yl4Rq4Sx9x
DmhE7QL1ddSoWdLce5M+Ag1S+u6PYbA1tx3Kj9gmhoGeG32tALYe77hbNIvy4PfvmT5CksqeiGJe
UBXN0Fjtkt/EPBVKC1Z7BXfA2OEye8n6D46C5VdF7lVRtKNpU3aW3zXnCSBl5YKkQEvBTAX1qJ+Q
18c1+bEeLDZmVmAISxe1S7jofwbSZb515ySoXr5j9DhJsS0uRJWO46yzuJsbEyhGvp0vfr6JbhWh
SfiaouIti0GosarrT7WXN9SNEvLUuSuNNc/QiB5H7kkhAHZhAKaoDBAkI5wjxLQPZiNtS+bbE7Lm
zCONlZegEg/LUX/5THlEROUBGlYpqc3XZbnyeXa922Oj1O2tiOzdjfOFfDvAr4du5sJBjYFuIYAY
BFW2450Uq0oxsjpTK5KGNAtBXKC6tAg6HRCF1KwMAC1DzoOSfGEOt+Ixyti4om2fybYueuIn3Op5
DFjldFTapQ8vXsByi5TzH6B/04RX/cxG1ZtBYTP2GK06PeIfKYkR23T+xBkKTcosxLN4mvXxFlw3
YrANnEQhnbyUZP1f2vlE6cgthiYttMDTt0duKE6feVsUsdXHSiw6xcMt9U6VU+A/TzFkWYrsLkij
aW8ar5tvg9F81FauyKl23cAzWaUqCVYWw3TV+TneGbN6Y2mp6ZDnzugdcoxpVUBpuR8+UkbsP+pw
qKKB47RQU7kRcBoLSUqCB1rH+J3z1ZXd4KgqHn8EdToBz+dOyUgWdgegB8ipeZU/g/LS6Mv/Xg/Y
WbLwQXEOGosqDCnSGEEz1OMeDkk3UytXIyCXoNbvnIEfL6wTm3/PrmXbHZvg3IxYcgZ/aUxQZPeI
3V9/b/UE9abGp1lJ7wjwrQCKfqnhiZFHKNsd1Snm8UPtIbRNs99KDU5BtpTCExHBcQ9fI8A8dKqY
GBP7BYQALtAl9vhNgo7WPgcXt1RA68APOStGlATHTThagHHiuuG66A7K7lQnYcJk2WMVe/IkIRUA
EivN4Dv5IbIj5qOp81DzmF/IYOL0hn2HCpDlTZ8tdhPWz4l9Fzyh3vz88yKJUGVc3HP/PU9Puan2
4Leb5PMfXPIEjnl9lY2SQyrP+Cgt6XRGefCVRqsq+I9lSu6AkQphO3/d6IA9LQWn5PfljyLod7sk
h5vNJc7ViTzYNtdbo6Ubn6QwQX5pN9xGYv5WrgwbhYjCIo9RuDFWcM07yTXaU8fb5gTQMRSFwyrb
D3cShl7FGFhWdaT7JPKxCy41GOn92n482kFITquQlui0XUANE7YeMnkfct3cOurWkTq9YFzQxsJh
58gB+YSZMBMqUdUusLd3PZzHylqRaptH9i0kMPRxvohqF3AszubzgXQDc1o+S7Nupgh1tKwfHegL
1GQnN1f/V6vB2SUJJVPhO5YWvsivu3KP/s01bf2+JXwgx4tiU5OAW46Ugq+VKrKu3xK7TBWxF/KP
NvRGjyLaNe4XJLXbryirrVp2sipACwjgLaApkVT4CmyfshPBBKcl6PAU8hfue0jINPcNQmfc2UDF
YuhNGsKvSw1z0iuD9J+cFsBHpXCBfQ//0duYEAN7kLNlD0L07wChLpMxf6DZ/ObVgDu5VIvIGahd
ZporWZ0D3KGeG4BEFmlXIDayXX2Bsbrn7ocMHV0PvZjwRxDDBEPMHzIraGce7I/8Po0E3f++xcxa
/FYlrrxeDtLaeUjwBBAueYDJbf05jBdaK7DslfjsnqLAUK48EakSXbqIc4Fzc+V45vvWS7wQai5r
xSCZzezAJOudamM4Nck0YjjpXU0McUKdtB56S6s7AnJ+nR0DnhNbLfpbCxcEpv3x9KmayH3CTua6
wVpyMraH9UDbMVvXgG6dFEeDtrRL9BXNx93ybVgnXInvRbPdMxG9xYWKyrAfhWJSZJNTJ5Xif64Q
tXxiPS0UVtdHca2wdqDND/CF2aS/SfBfUR3fxPuUfdAOhUckefxDxmX2YNztmbLdiCSZFAyDgjUT
iJbjX9TXvLRVrt8mbU1eEP94ASl8zeJ4H9XkNPQIZmtEfzuEfE+i2mC34+hcWYQg05SWm+7TOWFf
6Qt1OFZHcfKaQtFVbK7xNvN18bYZrl0K4p1Cmfy99IDj9oxpgFheZbqfruHPscllgMiyNIxoU7aJ
1BeG1x1Z/iKNp6xvRje8JcddWZ0nw5RkTVALJ0d6E7IyDr+bNDuXbo4TfUeW5UsxODwzICU7FIS9
jZnviTKzE6AVALZxOfwvmcNFkoHVdDQk56cXeXXZNnY+f16CpPYHNt05642MDNgpm2M4oEY7VdAf
jg2LyGIiSLpBGm9JTWCYWv8Z9uLxzmkOiP56+dTmw1Vh3N0zTLbw9W35RnQAPb+ujy4f1EQJIDYf
8ngdCVJ1As56zFnUc+ku8bjhYhIFBW5FJMDyn+Me9BaUE8amxEonoHO5eIgSG/mcdr0LL6hHKodg
8v5z6t2EMYLJfwISDzT6KuL682Is6xOnfI/RURzH+qj2wBMBEwFFC3wdpy3ay3h48RZcBPxZ4SvT
7KObOUAoIEt9boJaO/0hq+tfvSfxI/8bx/0HxkRy7LMnOPviEsNt2hmUePNDXsqAk9Xy3RNp44Gc
p2kiZM7I2sVbCnhvrOp3yf4PcaTB5daDHaeKBC3rW+U9Mr0ICvcNc1FfwsSVh5NDXo9E08gNZ8xT
hKF4caLLoKdUhhr6zz4ZdCAks7apUyOpekHXFPro/uN76quVCdLX0nUu/UbQNfHDkDTF0OQVH+ns
6RA0AGg2gpAKjtR7BCTRJPToaLKjxky8lyWuCpK8gc1CGHGge0pjWdRdVhOtQ+H0J+2nb73FfsHl
yBzYHKuHqZzJfvE1V6FnrLqOGcMDWt02GIYbxWn531rtXx2j2voK2d0wgFlOqmSbSn6l8/fsNeff
C39GO+JeMwIQObHbiNRpFiHByTBYIQzSgOOIwcB3yqTI5NYql9Ceo6XnVfq9hSs7meKzosMO8u7Q
+dhTZUjIGek0CuEv2YdJXPutnUCQnTlb/6SaV3yhcZaBJIYFM0wyon2d9V5ro8inyOYZbWcLaumR
aHPKiESY+cv7NinAmMdWwVuwIGR7DQ8r5Yv+S9W1ZlM1omMBnrIfqhbymAOi2exxUi7iYzPyji2e
E92rb/bLErJTKQbi+l6MyAcCFRSwz2+ZsU7ZF42sSgeF9nXrj4jAJ5AqrIaO7W9jS2E6wr4sOL7c
WWGfNQqt3LsOXGFfUgLmuPMhbw27BBx84vHAHfH0GHytD6LseonsnjYuoLSYVuT+5lob41lgTYd5
i1eqA3ld3X8Xbf6EzZn7VG4Ui6W4xfZ9ngBovwcljx+pG/IbyYwNtb7Osc0aODmNB6Ym0yZo89Ni
u8FKaNoY0xtH2GKChWDhgFvUNpYERpsE4Z5ImVH/r/8LcOzRBr+HNb/kqwijxKrdgbAycYTALgaM
yiONP9d0JayR1/vq8z8TXsM/CpENxEagHZ4hqYJMl9Rgrx0kFhwqz36O4XwRShhf9sjzK3zODuEN
BFZQkK9gaa+4QpoWktaCfAXGwejWG3XlfBbDjRIh1UvmvoGplYMUcWAVOpH18A0pc7b5SXOwMgyb
y5UtnHQZIOl78RzOh0QjyV/OTzKaXr6Tq/rVRSYxbE6UpurwhOMH7dLkEMc2jtMrf7XBHl3uwUB/
DdQlzEbJufF+uDWF0E3UWx5ea2j+zZ/y2HMYG+ffZ0lTFwhltncN1Trq1IJzKissePTx7Lqc3DI3
M+vH+Jn2xWh/O63HWPGtwo5XQiM6mlD1fZ/z6fDaSv2tM+v0Wqp8htjc0NnR1a9BM/iUIK8t7gr3
myKpXagNycvmUL3gmo46BreQ6zg2vl4+ob/1a78FhQPZ+dNsmSp7vNXwiL192HEFvNDO92GqrxwX
Vrvtmj6OTY2KxvqT8wD9T1VK80VGgVnlS2BWMSaQFVyDZ8OzpojoalYzalsOI2yZvY8yK0nNNGhq
aNutN9444u0pgF50bttRBBRf+J1DOMFP2fERd/alEHrfAxI+89/QGAfZru21LJHjGkt/hSX3wO2z
LclTKE8MWYZFbSdchMTq1Eb6g81zobgy4+S5dLNTQJxrUUeNtXh2vDUVxaZfCQ9L7rOK3UqCgN5k
DNyCMkRkweTXk4qQ+BH9CC/y/8Gtm4wJKC0IuJIkT2oRiBpqPufar7pJMFyH+I23Cpvghk0gayK6
jCjR91FDR1HHZbWTTw4e+N9Uo27Pryu0AZcBpWq/XZgKLMlrV5Mrv0oEvTv0U+AJwFmOJisZpzn2
9TGv3aOCpUBeKLovJtLDScaqFxvMOUQ6SpeEYpxE8Zg2K2HtD0iQXCaFhBxqPqpw7ktkbJc4G8wu
OsDrAqTHtd4doLou+pX9ktTjkBGyrLyHEsHsYcXWlu+MRYyx9NETsx/h/C/oFLL3e9nV0NdMfNGE
Zqj+/Y+JXS5f104WDRgmg9kWhMCdhDvjI3Eg1l4vfEc2PrmoYk3KxvxSlqgrLypIXeNQrbcuRwBm
Wi2Va/30iFn8OQotuPd8mOGoUgTSBsyvRfioz+NGOJXPROJ+moEH0CXHd3vQO4chGhOr9N8w33BW
vnA0apfQjf1OvcshvAKYfdINTUmSPF6ERyE09yv4z67o4dy5innCdakSAb43L9KBc/gMh3/pqSaY
Qor4+i7MxWdJYMJmZsYJYPw8liKRPvSSEM+szd0iWtpBhfUHBBY1IjdoM9kWhJGZ3zhf0XIzoT2b
w9BPHRohhh4jiSRSdpUDebxDiJ2oZQagEPr2LFPYXtk2W1/QA6WV2v+0E+UhdryM3QUjf3JWkIul
VPqzVoFQ69oFCnH0ZCFKykMXWX6gbtKky7aUNnqbcnRacZEVoscjkuoiQ0RTzrcuJ4uG3xEc0Oc4
lIuW5KHtVhL0WoMIaVycI6o5jxpXWBvDNsNRFZTao7pqWSzr3Lp5d5UkjOYGLBJT+gtgroFYgRy0
/Wh50ZiErvpMUeM0q9Wig+ymw+yOqnI8MtL3d0frMvGXn3tB8NeR5Gi+kgmKr+C/wxkYMM2B9RTr
rAaT2tsEjT8QvYEx5BF74Nv5H9QOyeanVfx1N1XXxvA9VbzMNzXJZBQChj1UB25e/4oXaoA9HCoi
CC+pqZ0JfbLVNa36wSfkgOzdvp2Zb/DWduCGeXMDJJhkch4e4IBd+b3/bXANVp/I6DLzBLyFQb93
s6ZcOsiAMzJ9p1QgJr4PQk8BFoalowawzd9enQ9437yRwo/n2nC/ue7ZzDS4l/0rxICaitefAtaH
hmMoJ9HPxdm4YDSlaINfHXpx7KD87Z40t+kq90+me5Jm1itFErWdQOi49O8QazXn7T7sXuD2S2Xr
LE62T+vxzcRHCKFT9jN1BrRzMYim00TVLFJELADbdco8Q552GlyocueCOh++RBVSl+/bhWQKt87j
XGm5SsUgg65zrkJTssayaS0+6TJvMrNaNyHYzhWyn/sq3yPbUxZnvl97s+gZw71QDiRn8MGH7rM/
sGnqjbnry4Q42Chwa6BK+LcVeHCR2O3kAexHPLni6js1RvIfL9E/SXjJ6xtXZXLI9O4WGVrHKEhP
YFUFJSK+sU0saR/7e5hyNbPbRRZkLP40O5MycN88qXfsqG7xN6kchH2f9RYx3hbm6guk0h4LpSU2
ZKIKvUZQKZJOCKzxnkvnrk2QEN/vJwjiVnb8JZ9vNwa5VkjMzH1h0yqy27FMz0tAgBcPt8V5msrS
p5+K5rZgWpvzNTywcBq/v0DYqvQ4Ed6++cX3N39iHQisCFR9O2XcC2cDyChU7OK7Oifzq+CtmKX1
v3h7cFokW+bMx7DHh8wZvJt8x+/+Toi5/LyswkXa5On9k6TinSZf9t9mTTB0uPHgCoH1YEX7cM8R
Cu/XTKHJHPSSZoc8uQ1p/6yKfaM2G6l/moqa7EBZd4u0Dy/GjjbCGKXmZQrryglFvgyZqiyu/47f
wt4qa+Ls4/5MoA692ZrX54tY3XUwQXug/+/h2ntc/u/J7d0ZATHDRVSV9QulQ6Ysi/8hCmdDnlFf
/qe1XVo0MUPIQcQlwWtfya91u9EgWMThL/CvORBUY+InPt12MemtVtsPpjzm3xFMegpKSycK2/kA
clSewDAvfh0u6w1Bi4EmCn+Ka/Kv1hF+av4/d0q1CKVYGSb4sRKUF2CsjthefSnMQ80RpmsxXbM+
nEPuJxea5mB6pxQDIeRgTKAhiM68er+trvv9xI8oJPhO9NCB9DEQBkpVb0/amprY+5rNTcTMGk5H
9oDWHzjaXgvnEeyMGgKo2hHshYwcmEXY43UUM6QTheMWW8jTw3s4lGStHcq6+3OaQS7CjZdaUZ0f
+UwkNOwu7KL4abRD+POdWvgvPPNdnwoBmZltGi1YwC1nCddRCDMd9xeQXW0csor+CH/4vHRtTlKh
QeSuDpTXqyI5eleaK5u2QgoB1AvNlPqIQiD0/pXCfuMjzdpOgUMO5TQ2IkjDJ4EZ+QdtMu7ZlQa+
KthjUiFkKkmLII7ynIAqcr99aAwbV/7hRUXSPrXJeVxUYEf/3YjiTryvzN5N8/tNrq1OO5Kqnz3D
68rxWSGYf//iUMV1Q+8mchJnz4mPTDoyDB96GqZPizBbum2oFy9WaP1IsMmSxcJhx9kINrkn909A
X5rwZNhL4Ms8ptr7CoXgxUeidmYqzCgQ2N/cld5KStQlzHcbl9IzdPg18izDcokh84CqC76hQWwt
hApSRV2rjZJiFCTK2sAJQGfzZ0GB0RNq+1xwwTNWbtVO+z0HgN4k2GL0B5Wizgv5lr776yTTULmP
ABQLD8VcNs6U3Y/T7wmASQRPBncqNceS9DC/SJG7eKWO5I/hwrtimKXEman3WU6ldcyw8qu38UKF
UEZejTikhzRT6pdEsRiLF/sxxfq/ftXr7xETp+UP7lg9cU0g+Bp71d62pQUG8Yt/p6mbIuV/H4xF
d0fWeIQFipB9jXgti5QF49E8gVE/DaKqzTgCyKwr3UvyVovcuOtuU9sMdzLIaaQGlen1vtvngDrc
kd1RvhLEEzhboDSAzfFLSNiMwYwLj3po1JrrsiMnHUR+HZx2ilI5iTLnELGusark8FIDww5qjHNj
HR4dHuYtY21yUqqvrmBHGo6tqeA+QSd3+jvC/L7wZKc6z4vaeHarjQL96Zb7a1gy8R2eNI24G9lU
BRLU8C0Dco6uZKgrwFfE0kJRW2ItHEL51GGMzDcOcdSONqvpKYCas61XmBJTxWxOM2ILLYEpTtlL
hCEhK/lI0w+i5bt2Nuc/IrHVpgCAQF2yRnNk3nU9j+wGNpFS8uMPZWBlw8lAEMxOWI4AI4aGopoF
BlfeTg/potRGJbWfxtjE4UK0vb5C34VSErUliUqmAixX7JceHaGf4z3dwagRBoZZFgjHmnQMO9hI
8xoyArVpzU0vCfqfmxPWilPbkPF4CV3jpPeP4J3p7SSCZPVb+I4fKxJBQ2G/ZX7GDlkld7Pb5vx0
DLsdZ3JKcLB1paTgxQU0hxBan95iuakG2lWQuBb2sLtPkwQ/3vT2deuorW5VMul0Vk6uIb7m6qZ5
MDbyv0IMOwo519YUz10ZXWX4CYilqU6syDcCOFdvz8z657mIUN0Py1USij+/nDG4JK1m7E3Dd4MP
P+o9c91Sx14GmTVUM5NEZICzTj4Ki4vDsdjc5as/YjQMtk3kPSu8f+GzViJtT2JfVxhCHCsY9Oij
9NOcQCemY0oqSfpkBh6DwvQwqJkLsTuM/st5pjuRAZsVyoaOCRMB1/TvwOE+LzBY5jjjp7G3uZEA
/eg5CkX/LeDsGtC9TFwzuD/EUmT23mWWTSyYJb7Qav9wK7bNmRKeZx3rYsHfk7RMlxeaEyr2UMh+
OoJ5MPbEeTmrboki+7on12Qd2R/SMoqnSNW0IF88vDvsTv+Q/Q6OUE3BTIbRPijqVO+YIN0ZJIc5
Bt4gDFd7wARBW7sQdZrrZJ47ta93pjbmuZ6+ROGYaDFWWA4QNaXfasXDLNq6Q6HgAJRjwoLlD5N0
/GNQ2WEGJVVikaZscjFSy8P9hEtcBYDDCd8ABNlQs5RjET0hHQIHvDTzgHHoNLFNtT6Poapxc//2
zp8UNoKhpkPJUBTPVhuaZjO1U2/2wnS8grf8a7g1U9rwRZ/9OFjZjCaURLAHXsi/zcSmfC0gOz3L
1pkHUvVOXFu8OsOIrd+0YNCRbx9/bZ3UJK8aQUotHfTS+mD0YxKHIDEe5cbglkg/DzvDZFLEOUVT
J9+EmEcLn/lW2kac2fBaRCbOk3mhPOUG6hnTHl1dKH3/uuwGw++l/P+sUNUTDgHIdPcyehEcmmtv
plM0PwA1MDpl+cZORU9o+Ug6ukqCF1bZQupkqIRluK7QMTiSIXC9vbMMJmUE33HuxoPRsWvI/lF9
s1LZgzzOhHOFKBFCkJsLJkLZ9NEWRYbX3w9Vdf69L7aMyTQ43auXG5LlQS1eNS0Z41eZ5wRzb5Cb
8AL3htlzjRCYJ56aTNNBpfaZ5Ep+FXXoQA4iymuoa2HlKi9IbX4edG/tXQahIaam6/f6jghidl9E
GWaY4ZUkcm1/l3OlXmy4aa178NO+bXjsyTkV/mPmhZL1BuTVnZM4SFTyDk9+Z86BoFFLrFZeTNHq
dKJ14vgXBM8u634dLQd7It04YgMSOvmpuIv80280Ug31WWtwThdIUphoZr5uG2XuCZ0AkCVj84i5
TOQFn8mzlkh84JFYlt/Zm8cGJ+Y0QzA7QrYEKsF5zpbfI3w6rC81l/o+q5n99VPGm/uvpxm6BV19
P7MplkkuEMNtGDm9tNNVHOiLAouLpoz+KZ7TXxP5QR9nR11aNjlAua8WOBgV6dvYkpEaRKh197gn
ClF8oJ32Dv0cMPz9p6q7wZAxCsjlWe+5no/z77dR8h+gsajePotDfe//icj674LoTQoI4O5l3z/Q
kMZ0VkJ0UBmCrePAXOSeePlWR7T1WZpEaTuqr0GvrD7XS1TGp8FM4CV2gxYheHsr2onggmPlq0i2
Vv+JOfdGQRVnw+ErsMfQFidabEYFiCCt8rsEcLKXJwmMULVCq6QgYImrlHFNQcM+WmUm35BVwFPB
FPSoNw73wM9sOhHpBt7HUXc=
`protect end_protected
