--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Ps2x6xrF1MiOXgPfCAf6gSm1ki0/6G5rKLcsDxaNmRiPR6X1xZtE9BOno1nBdyQFjPSJQp5FYlQ2
kLqLUHpIPuSOzlfJZYWK9k7PQPQMrhwYjy3rENBYFC6fxcgqFHGXNh/M+thavo2oWbeb4I45Rugu
+P1+0Q6R37cFSWJqyRwryAHZkDLVXtRU8TZGkyAP8wObEqkYwfz0pilxKBnyEDKyvUwL3BRFOzjs
JfI7Y8DbsoDQl0tPPPYLSLyvnm7i0oP/cComiNkSxSt/3WkbKvdqcpPJ9JpDVN5+LjSfq7KhiXDL
jUOihrIuzSzn8Wxhc2azzTwxzS949HJWqzpCwA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="jlfHS/Vdh1loRHtYVBSQO795bahl6b9owLN64Bl/s1k="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
RPhM5lb2ziGKb8ItDXQosL/+V5a0SHqZ7iSNMRsqjn9+OxDNr281YpbRX5oxXn9ELkzTtSnFrTqw
fTBprYis56HX/mofrdpcXogYdljOnxyp0RUg/6ZDcmcmuNrR3uHDP0xRS1qhaJm+x7g6e7S+g09q
KIQMj/zRq29I36ANDRMpuza9qLPk+1h2eXrnjhDVcc3+tGkbYm6xrW3CURUnDHX6eoC6PjIRmx2i
ID7o9CuC5EK5uB3mmEO0bpPa8F18ZxAkcy3acC3hYhs5Z0cQWXlgx904z2PB02mfsmwTCJqGpIgG
ZVXY9kcdHfXSzjlBCq4MWiN6n20wwuqklBzHhw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="eXilqFo7LvGPTtFzb/9Gcdn481N3jMKCR1a9bl+LfAA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6624)
`protect data_block
3Qf4QFuqJCqXwhMCk5/petdbMzDzMgPXRkRU5kmp0WUmy84glzgIMHdEcezn/93waHXtTAJXHccg
pk5pPsgqVH+e6t6TgUJBuKw6db3VfUpQyp4tiQO7/42ITMT4gqchnl+/expLhtRTUafPvZumbfiF
Ck4iWdQKOcGfAxbGoyEP3x0WB2NGAu3DynlUSrQ9rr1BU8tv2gNUHZe0oirgX2tbIzQmy7RsQwIy
6pOTB6j1FMswZdOvsl1mx4+SdmRBSWzpos3TcD0P8pFLyOh08EuWCItkFlSv29uV+evQZv3QOaYK
C8JHbSr0NbllhbInHVIUxCtmcuv+er6Ed2W2qydM89lZFYpvYRKBqhHrc40RmavDXs6fQHqj7eYu
qH9L5wW92lYy6wDJeM0zdUZtXixYS4+ze2/JafrlQ0yNMhET2/1Um2SqJvsv9ZSpgZoHaQfKz2SQ
OkcyAKPK1Pk02b2dlYlYzEDNk8ScNeJLjxm6RbAuG+2sG2WSTJZmQ6cUZmv9IJjygT1Zr2N30QlT
6zYPzrIf05aU3wL25BGCGdgvL6hCpa2lLQA2bpRCtmvlGGXpOY6AErwlTvy2pgEga0FM36PQzapW
BMC1ks4koPg//A/zN0c31iQfS/UAUsS/t6JpNG7+74b9fjH+s445g9Yd9dnN/PzA2FFh4e2/ExFc
Qj4ew1s/VRorbNOLY8OYp6aOG2lb4ytNrWB+5mo9nrJzrRCzblgYa2eSOV5rqrOTa6kmWSzW7ZMF
neBRxPc8uS6m4Um5w/tXWK0qfES1AVvMN2O0A76Idj3pW4WCJIWkUxPAh1lCESlRCpeGDgTkMLaC
uj+UfK7q0NFYhSYpG3T8Kjzhk5aAt2YzRVs4sCaZqTUIUIOYVJ0NYkmvDY5WS4O+F+Sye3gthHqZ
xHcCfuYbw3xYgn9ZTphOONrYSe25sR8IfbPjZO+hEHA4ax7VsuxPfkNi00WzNqUFt9feqTeaL15U
1yAatCdeQnMaqGkbvnYfT2e1b8Ewh85WaWIL0r0zhMeb25RYjgHHmUfcD1hLcaI3P4IzYoPwgNnq
MFhYnnOVTOBv1rXqXrsTKjyI0CEfqCwCdDTHdWheeF5nWtZNXGNDVf5TQOnTGFWFkeBOLmHfkuDB
VGBaDsn5MT4HtqS3u5DabLsR2GD+/a0cpPyMGX3uhNVkP4PVR3ckl9Bl4VL6gL9UuNgdU7NpNwJR
SVHUWUVvU2+hfupPYA/GkhJzlECCtDUxfBovM33+d6JymMw80gCj64PPRn3NPvSzOlDdzBThrHt+
3CtMM9eML8XiCqiqh35HRRsimvBhr9msOJwEIIq1GSsHPITbrvKu+pgi3lAh4kYZmYqf799E/0Dl
IZTy8gG54LUKs6OzVK9r6O8heFhl2EtDycNTlTytAHJI/MadvFBGDuIg8zRuIs/BK23wPWeEmV0C
Kzjm+pGR02S5NQfWMHzKgf8ApKYVohWLzYUhPFuFwdPubBVdgXp0JavkOmA3yviefBcW6MMfvvci
gHYGGIap/kp6d7BQtr2vl9JusFI6hAH05NvU/oI5LeJZgPVXoqdzy4ZGEVDHdhNYp+z9vz5DzwEi
6zIpFEDvVoxzOygK2n2p13S6PByZm2FlSTzbABBJ79w0HMIRDOSvSags0Rrngk86264GCvPK/UUu
/YThEYdru8qtOVHJLf9naTvBIiwJjmk2E9ZT0+DRgDapNwG6QTojw6DyT8ddooy5g7fT2mctpmXV
VWxu6iC7yW/7f2yyqkl2j2YxhXe0BDkMJUqFXz0XP6ojM4MRBWodGDhOqBkOOR4xfrZPaH8BjK9/
5rJuQWWgthr/bNb5SxnVEs9k5uNxMSpP4A64cwSj34Lb4WHjmqtsI4AnYcL/72xZfZzrBnV+GAYK
6bk+TqrCw6NE19NEPjB/IN95BnMgPwgyBgL/fpoiQw8NfoYnbIHZXgbuFnlmLajKiJwTfPTgz3fm
X04hZvl04QEY5XT0ouNoBizRAh9Wkqr3+nAabupazEWqvnA3L2t7mytYFVuz+dRD23bf+v9EFBTZ
98yG5ir0KApzGfhpF0wNQ8J5Bfb7/CaYy4u2iNMOXV2TwnUQlkw7tAd5pouOKoApWCIAGLoWTCHN
hWlf6J7Ijrym8EUp6Bm/4gR/GkkUYh/crHBYDivnUcVag49IPOOoNu76ww77qApUIchIp/JMBnSO
iF+pz+Nm36FJRYNIS7VDSB9gJF4mpiNoO7coUXk+dpcJDYLKMOBQtA8EMrN6WU04uNw3pAQ5IFbF
UtaF40Dm7civmJjijWwwsgoji0HuUNtxNHA7dIvx5INap6drJ50FntZlJFQWv2CrF2i/8B7qBDve
D12yP4tiFPrPIFEOqgRS1CMTj7BTRKldTihtmYe+EPfTkvLXOE9XmmPbRSL42LAHcvOQwMPY1flr
tTyFvZ2KXSS2BQCLXNRmZZ2o51WAtMlnPmvxfzEnQhErTPAWcFgtFkAA+xhw980XTd3L02Gmf/AS
sedyShPz8dHuJU/gsXAnCmPUywfDtuXmB5GolNfftBKdTsq3oB8O6ZoXrmvnUXB/P8lc6zcAyw2E
2CrZe4yR5u1eRmEiN+32wszDIwDjQ+fJ/yiQK3xB22VxHsGSeYX6XEzSC3UuBuxydkhup7p1UujV
zF3agB6PFCytLmjnFSlMBFNOOmtvPEM0VYBZNrBtLz/K1uDTbgKwuItrKC2Q34lafmJt0Zxj79Jf
72SdpL9zxVsykvlVFygUfjGmrojxzvSUx7+uwzuESRDEsS0UwhkwCqc/+hX8DlN4F0eb+LqKDp6S
ZJIba1Xw3zmA1KKDfIHwUtmEyLv9nZ8F9nxNUk3HYaMWBVmecFQRqabcFp+TTUzEmsqUU48Q+DhY
y/qyM6zCZsCuObHfgKBXyrFYLo/BQwLTWTyd4g479V/sNTDkbQeTn3iKVHYfuGJ+4nZ5mIp6WwCo
id02AqaEaWRfcN7tj0veUgV/q6oL/hjG7DOOWuVYu6yIONeZ/FNPera+nYcpirrLsCRKCONS8PrD
RxCS0qklINhiZNR2fBwCTqygMK2TgDaZuwtqbZ0PHyP0NYoRxd4swbKQeLPjSYuu80sHro1wFZ2N
SZ4kKURZyNedQXCRd4AMRbr/nzCJZieIoadml4wbeSyR126bspFA/q6gS+8ZmxQzsMEY2eM9GeMj
PrOvetflWFP3V1POwxkA4U8M+6k3o8KnsE3BOoX7mlg/ceYdny5uAgn5TZqRdY30gLQYthO90lHa
iixY0j7IpAsDGPO54OAezsQYf7uZhS76TCc5j9ctA6hsHT9JsdiLmrL8NOBwnABcH53mvTDYj8tT
MvudlXy+9BjGhj/6nRUVRFNkXW0n3NDKPeSHmzBGm3TpxN5CsDBhZHx67c7nHFZOw27cSBlPUq/+
eZ+WLNwSMHpDUL0OQ+dqm//G5N0g9SZxF84T0Qoe/ktgRZCuUuZ1v1Lve2AVGzinp3F+vck2ggcz
tv87bI+IvI1cjc/vt/pETeKG+kEB5zo+EBL/x+YA6mcsOMBPC9jXw+tHMqBMRoKnI1/cUg8y9t3z
KZJ+nPnrBPxk3P+NVZwvN/m8njjTNBH+ub7jBapmplP0ngsE4rw86vcbKBRnnxvWrCmOgdF+rLQU
FjZ7zk5IsEIawlCbYRJEOyz3sHKuErQ6x6LtocP8Lx9cjvyT3Fp4IlCtzMyXdkLfnHPjAdRBR3qV
OwdLT3xrauw05ffY41lC92TlwCUOJi+UJDrdB4iRgeafVEKmAvqP/+ogS6N2ShIdtL6J614iCfsK
vsOjgqyQjm3+ZG4RpLCFalw2wbAtW2oWThRHss0Juor22nEf9ISPdNJ1GPn2GhnF+2JaIky+3Dnr
RVqIkrDPFcg73CWQoN+I57cHIoOBUAkoH7xKqySKKb5DZ/OmyFbH7ASmunpbOKLjeohAcq79llbQ
yxvVszvEqNpyDgpiFkslkXXjX9wFcPfDnKC42AB7GBxAMpCWUWI0sCi5+zPP9P0HwvLZSrQi4Joi
kYmRIj+cl4RS3edGuoThM869jXddhvO+78de9pcI7NmSkNpRo2D+DIuPeTHlH0vnmv5PD1nH+xFP
TFJRaROGGYt/T1wxZCVxV4ADOIPPksviUvuVziLBo10wslnW6f4URNMXrXkCLLG1g221C4OqgJeq
tfOVTuPeGq+9J2V1/dFBpHcbtPb+An+oRyHAgBM9axkyuwGg4EgoeBxrMHi/bCdsBmWNct6sK6wk
JTERRGG8LkoLaUkm+8lrmj37u7DtPsGQvqpr7FWJCmtLDfko2/sgLrcRaLG9JSRquwt30lLYRhL2
3Jub5K/8DOo27XrVPvWXWCbhXTmOaCfkjl2+7xjRiHksdx9y0EGKKBn/N1sWqTkTwAmTOwUBX6fi
cPeFwkE4RRzTIrMhmIz0YP5DykENFfJ7MY8Kq1rAuqs9MZR6eWxgNe9ZQXRvAGPMSJ2w4b00EmVl
7Q0+gbLoLCRx0OaxzP2XH4DrhLGZw4ZlAwxhLEpdu8v/VFBB3cJFRAbKOvCZ2uA9Os3IQShxNrnq
atX4BB1dRomJYrMBq2TLibsu+BiGlkbp0Zexl5DDkrfWK0FzzyXCwZoiamQUxjzaUsYKAVMNVC97
m8u+bEN0TEOivw+OkxPoUk6xTJWDh6ck/91TCgsh+ola2a48H5h5NQqnZ7TpzaQOqOiaHrdU+eb1
+GpHhjykh6mu3qMn4EY0fP9fp0qdL6TUtx+Wv2rrjpEATPa4H6AkhVYG/2/UuDi5UKRKV7SB6UkK
F1uWCylfGrv9ZgackqQPovmEppDfN3d/u8Q/U+zBdsltsiYAVw1VKL+Ib9VSyaQFe58QAaCw+1+0
s2suBlXio3hClr6r67kJDLfiFVDNf7w6phrMfrwqkLeA9VBdcUlMp3YPVKCNqcNaS95DF2dcUEgr
VE11Ql5gE9QMoZyr/wmTB3+s2ClzO9VMDynk4JlW50JMhgYVenw4jZluBQSyQsNOSq5bSZHi2mRM
qnDKSA7h4EiCSQxT6GFQ2dB6dPnDFTMTljc4KIz6kLy5JB2BYdRSTCWhtxSiTeZuPj/R6C7qKPqq
iL1PTAkPAGhW0lf+XBINafD2eHwh7t9//2rQ1lYl4Ih2LR3KCLU7h+ek8qoJh2RDTU9e3YQTUvXX
BAYntUohcQVUo2QHwwNkgnz+7Ry+zToiGpZRsgD/RG0HTeMwvTam3zMwAYdVOPJRelI0eXIZDK3W
FO4jct+fi0A84X9TEDa3J+VhffwNQTSTdrxviGysidyhrQUfVZua3n2S0tLEZlNcA5+YW8fi1s/r
QJ+wAlHQGZnhe+dUDiu9EKAPvYX7euSpTQuVv+FSnXDuJGlzczHr/4Lm1YfOi1JpAJFJsvr8Zi34
PiBF6ddVo1nrBynmf0eXzki90LjhKQkPAzUS0NhfEmWLEZz9hYmrDS0YTaCyFv+t1SiV+C+vfROH
8f1cb8BhNH/Te7/exvPjuJqk6jJ62nVakRPSFOdf80lfZHgDbd8uq4ipliqyqQJ/HjfecgywpaJ6
Leadz8+DUmIyRqxuP8flMG2vgWhp4hkHFki3ZNjrSHd03wKz1BMKe7XiVgPq9ord6rUIah74hZG4
LPrmL6CSNHiVpue7Mo36bKt7hIEFjlqdN+Y0iQIP6iRFZfAGsdUzNgeqKdNa/CEgztKND2wCFhhz
AJmcbWr/ceRKKFfnZNGmJl8wT2sQaLCtXP4Nr9g8HJW7MN/r7GwCL5W5Y2DwGKwySAhJotuO/d/2
ucsf9qsO/aDUp9ydLLhUv7o1WIDpq746B0nB5kqWiGWRN9dnHBK9hahrb07U/7a5A7FUVva7fie+
r5MQw8IXLCWg1dnhHc0W/jMTQI8v9e/ID6o7UKYPpQq2OL1K/cYrIKkEUScOYqf+owXjgy7Y3+zf
l5gK9nkOS4XaeWY6oGHpLjMdE2+JIohyc7HCu1+ulBYN8iGsl2PIZaffhoNiDDmBAhuvp2/NcirR
zN34mCSpnXCm42j7kBS1XuWb3NZFdnK1sQmxuFVTGvy1kG2Yal0tPbWf1PVrts16ZvTCwq3shQaC
S0hBuaTefVvzaYG6C5PEhlappvVlEI2wxXOlO6yvPARqO6GRR1cf/JOnqRhr93wxmqynoLsG92wC
/oOYcwf7j5ecx+hB4MuM9SfzZ1wb9p8BW+EcsSTDgcgTZkbx5WwC6B1zYs0bcRVXmMG+nLL9dXob
YGtDo3d5eWKXQ30uCcgAdtRgu25EH1y22xXtRybRSmoBPgVaGoywBd3ckpIm9MreLTaAJ4znESXy
f43D/YMQhQvdGr21BsQ+42TpSRUtPyXB9e9RS6dhbqWp9nVkdAfCmKL5apa7WtLXMZhdAcUyWBQd
oNqLZrXR/3GzXjpPm98RI9tamhfRYwTSJj3fzrBbcnrkbuEax4tQ3Et6RDmFKE2yvgeZNRyXTPZK
ISrdDUO0Ft6OalFKyT5fy6eAxf0peysNqBj8iDNZvGnNeO5ylTG9ZFmvkcomflcVZm7ZlxwV2eLg
ndHIdp3KP3ECDZKuflBqVlQS+MXung3RUEgJLX8g07QoypnZ8MzQ4ClA7ZCQIqQsdtvP7maH0a11
Kw7LkS3bO5FHBc9zDZM0XVRBSeONRrQ2Q81F90bDRpPVj6R4vf7Ti7cmrAxuX2KPGAO42bxMXPO6
m+lukrxRclCYCBhiqOg2j4dMbL5PuN0G7kAvOtYYe+Y0CzjW83AKikKBWtvdQIpgxNMk/CvSmRwo
jDv9Y13hqoCD7d+7TAhgfhaMI/N2F7jt1edF9cj4AMyj9qEnLQjlY939WJ1ppP9cMC1jPumzN8Iw
l5tmWKGHU2mscAS4jTGsmlscGvrQk8G+btGXVpjAUY+pKHN/xXinIXAWMmticFxarc2xpwLY6T+7
ZN4WDdW9jMqODf1eSVLj1EFegytgWFNnqKWv9ZbD00+5WC2yL3BbDmAePdphfQXZceAyqzJ2c2KQ
QuqDVbytbilkIi0w5GQJsfeatgbsk/iW7SmTkFLm0y+lynNZIVlmF0mInqoguX8YaDfte8Ez5dv9
JECv3lPyzqsJYL3aoXzoDCMYYOlIECjx76htPHhzGvPVqYVxkEjBKkSKtVtogSwOXhoga7fNGeqH
Us5eIB+h6dJVK842LqQUmV5O/6C8EXKjLgKGV04I+COvhPGzcuVEr0F8z7TjvJsTeQVAvsiK53eb
ybIQxQg0Q9tpI+fl+wP2VLQaI0CxyFr6r4++PmTGlnxhSXQ6LccWJdOJ+5KwjDv6LEZg0RHETBzH
AjfFLGbhJ+lkKI2Nl/YTqRgohlEJRP/gZ4/yg+lvR/g5sBihCw5afkvM8Y7C426++6s0PmbwHTKV
j1vBf5dehJESCCUuYGbCICxiiNzrCjjyeaggkGJiyH2UCwOdnUYOegey8XxBBKtf4c1/ES+BACHv
U3W4HnqsgoryXbCXFy5yThFJCim+xmcYjQ7Bc4Y23X0tbdtyb4yyAmv6nXvZjhAgNlzW0du3QUtf
vybY7wttdMCyIDEt6XhKpFvyRZylSlYhN/0JZ42hVaFxhwbv5ynghEYPASHk/NfTYeFz3qAjCCs1
atMe3Za8E0YXYvSVCpqhiONvyR8sl14ypU19Y8CGIfw+IvQpgpVanxhxYD8g0Ao/8MCjVryVmPb2
67JvAzxieTZA1U2R0oxS27iRuYQ4D3rskf/ZidYmjjuWM8rbdj7GuXUSG1BeSBHt3nzGPyyC2D2A
We/JP95cOiawM5Jw0P1a+tOEx2QFQ/FGw0stz78wynPy0w4IfLrTbEKtu83voGIhpxhJeD9eDJLq
f5bhW/y+7pkIhNeAJ7/JbG/hdYUYsKto2S6sSAhsOAZJWFDS95gOfNeENGTp3qrYI1lThtBMTzBx
PJP6Ow5F11sDtd+tUGu4sqt02f8DY84xZUnu7Ef8+DUqeRulQShsk1o1QFfW9SlpEFZb65SuCYGX
NSt7zrL0ZbUpYoiN6OuJa0K6nfHcZ7YdWXjIkFtwE7AL3TEQgMJY25TsUDRwAl1t7EUmsXRJ8gWA
zNL8Y+GKfOYIVRCxpnyjLF6W9qguWByieYw/UguAT0Cdj4X1O0nBEC9PHsGadol/X8N+8GTZb27L
yefeUNRBmUlL40Q5yPTxtFRNILdWcO3/dl8QoHkfPuAGntUDW2yLLJbO7TxvMOyNnZYwYsAwOAE0
VVRq1Fqqq9CFo1XWuO9fe7yJxfmdFwulapMgILRgZb0hD8gVi5t/OKBI1l76NnllPCGeXyQsPM9Y
nJNJ349/sS98YgYwklUmlOZp5eL0iQzGjsEsqgqjNUbIYqRrK+105390jnXONSvT2h/aH1Z8VVKS
Lv4bgHHCScgmYadjwoSn6Ite5SC8ec7KDDfwmiYkr9+8Tyt/zd1We3JFq46uV5exSvBQtYkjO7JZ
H2JWQNYGH5dD1zhm7je/T1TvLrp6VBrRQ/VIhMg6G2HPBKX7BaJ9s5gNpeeYwfLVSIgvoEObAvYs
Q/jRFEIMGX/DB6UeYcCH7lZTjVX2vSAIitXfWdTTImgN9E9ieRDk/7KFThkcvdIi0qFLldiy+UMm
WktMBN4ErdlgrV+tb1UYnlGR7hOVwAS0P0lIu3SU4oD2lJ5Z6g9RHn0kPskugM2RBIBpF5ozCVXs
D7N/r2fgVoEJtosQSHSkBi8uybIx/qIQAvnp5KoJczRImX592NG8S2udjGdi+g4zeuLZ5MO7Wfaq
daOM37YU3Bt/IaN9swhF3rIP+kHpZxPvsgGhwejgtyWHQbu0PY9alrr6EsyicJaUjVYuK/O1dXiG
AYS3vZmAT3a6Wx3M
`protect end_protected
