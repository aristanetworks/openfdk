--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
R+PI9V9nClrePePuE/4fKdSqGyxryKEDmDU6ja4mtzlEZfSv1enx0n/+AspCGtmCV0e2/MGOVgwz
/JL/XhA2DwIzv0mNTlYeuRPBiyoJLciFIOCLzsZMOj/vofTNKDcBlqYK/Ij0MY9PH2VwlEUgKHTa
hJ/NFTzI6o8f/Os8lC/ts/G76JzTp1LTA5zLmJ+GFWM8WbMzyRBJGNwCt3egIzcf6l3kruIxt0Gs
jv5rR54C6bPeBLt0vabeAXvN7NlX7AYDLh3TnZE4ChEZq/9oscIoE29M8jZjz3SRHg0JdyHhsFaT
vldrFpZej/3BNBuK5J9j8TGR5vY31pbeQ/UQGg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="EogfA69cTwCL2pggE7FaJQNy5N2+SPvbUv2uKpWiVCE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
hKmd1yPY+DWl8SRIu9SDi4cwBcQl0o1gZ3E8iUK7Q0+/xaawyCXLPOrSsFzKpYjV5E+gAltJfpVg
DrIxbtYTszUrcBNAGeBGzBEYqRrvwV2OBlXMYizE4x+C4pGjppDWOXmFaa3Sa+91uZ63SujgVNOu
WerMdYKGIs4XRMSXKODx0Q3DTnJmnCT1XmO08u/t9J5C4kHfrWe1h1oErXghz+bIuuOhTq6WpzBT
gVE3PtYPnhVyjjhu31zSUHwMt897qg1FAR3aN8mXO1awEMMaGrPxK4T+WAh/lnJCkVF1ooV3Uel7
xQ9zZx/hBzhDQrCO0iENDYKSLpJm43QuQGH15g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="zUhAZoDXB6swoWcoxXAh6tAxiQ+oJmIiC77GtP021MY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34720)
`protect data_block
WoPNDi06gknuTexgykZ6tWeBouv7WO3IULcFedaTep5PYwAnu0RBUwLWo1eDdA8F90QhFcE6nLsU
0iz9lh+07rMz56NiGSjyYDveBiPAR4Z2Q5eOzK7/FDSuAlFzur9pz0MAAU7aqVdKnDbFGX/ttGb+
O7kZzbvpPtL2aLtfxCbjPXnJDQ4Vp+lbJphUxEJJMhKKiifdPRYTWoGmiMnfjjTF344dvo2vWdUl
ZKEjQQdGYe6fk2EFIOFS3e600TTioR/zJiYT0hFByVQL/wYrL1CS0PsdsdODT6vPkjTWF6UQu4St
B2iw27ifqzbSJbSiqwa84GxLhnaOQFNTJzR2n+vUeXb/jHdYJs8CeoeqrVwgx0ph8j+VnUqbeJss
V9V/4Ky8Ihm2HxHNqv4lIoTY7VYT/HEbtu4gzW9kcphHdOrEfivyX75r5wB1c/VZr0N5T+ZxMZlk
5sPm3IR90gFgB9qgljsPj1JnN5/TdSK1NXqq4BVal/8jupgZZG6fAyZm/xlulbUKa9bqpHbOQzJI
wGIx7OouUlXBgkoFbctrIDfUQCtdSPd0CFvJBdQ6R5HNqFlYaoIzcM2NLZHqAtOHewAXnwZr1tRU
aO9lnodiCGjzY7ynXUYUADscYaf0RGshZoR1VXiRxYUqoKyPw9+OFm4UJ99A+p6/dYP5fMZv2kiC
CjHQ9npA4lY2LcFurx2o9DoDL7UVOBTDBF03pUnyjt0JdSvNpyzeydfPHxRGjsF06FVl4/5u1U9/
CE1EtkpICn/JOABuvppIZnDq55t35M6SHctCNJRLEktGXVCbrxbRbejFye0rT6XJUuymM66HtrPm
4VzbxCPknoJF2sVKdBYrqmYXpjLIxRuXu0gSgnm+q1I26ErHCWJthsIHGYSy02iZOw43w+C30E5Y
uHiHgDkh8CtynZBYK4G5+M4Ks7zJi+8Us26ABZ8MbASpIJflFZeQdn3+UhiXF8cXoGdbEAJ1mDtQ
epPAr0ln5eJo0vAoiVnEtePztlxh3vHRkzuKsdMiGYEu2D0LZtmHw9/UOqrwMWD05aSI22UBca5C
VJF7Dm6uUSodFmb3tqs3ht0aVAvOM/PezT/OsUa6RB9IQxBJNgH/hpwO951g4NVOCrlcI95BQYNv
U4FZ47wsnmtOwxehmrylDz1os9F5JRT+k1R/VG1RkTrgG4UzT0Xbq0Z9/EKDm9UF6oxIZh2HINHb
1mdlcf0yqxM7lIw7WBwbfP8f1FFz1lFUKNWCn4OU4QcnHTOyc8nGUTAuukCxkWnVdvVKuctxCN/X
nsqvzHVC/vCpJ4dWu6poZw1NaIsTSBF/CvsHmhPFReDtz6frNLU43L6Mz/c4VHQ19Fizj056Y8Uf
PsEq+9sNV0FNE3PzA5fxSKvXxyC/909mSzRfCroLNlfo0kZ+8DcWRJRs81XOJ936TM0unnsyociH
Z2YW6SbDFKXyZQ9V4Elmax/9es2rMfOyEB4K+MwPD/rtd9W1onx4xiG/kruUuqRyaaxGypBpe27x
fCXcKqgI4aRDcSEcYvpFegX6kTJpM+iW3v+YMHedDVB3SkZCBP4awcs81iyUtDIVXY8qxwa26+5k
SZ1nn7rjAFevbpGfU8JO4e/UgGKrhQCe4o6Tk+hNRXp/ZKc83RCOsqyxH3YPhXtuDs1oSU35IkdJ
waz4iu/fasYwL8/CO1nMkWLuGvSxJu7y6KRJfHlUxh+GW7dOTLW5s0R8p2wmN4ia9LCkklTNHUlO
OxnZ+nU6tJY/7OCyoh36dSTOqMOu2fox9HgUEX4SW1Ec6pCPrEeOtEfRbGkcPLeI3xLwEF7NAmQD
FegthQvaQbWkW3V3PWJ7qwVXGCrF86A1/WI2fXuKKsu+z4yrlgk9lKtlrNW5uH2Nxq6lSl3XMxiN
t6pdxCUWHykrh/Wkc9zwyZMJxHJ2DVBDnYnn/pnydCuqz4MHApeheGyZJsrIlEdPq7x+7LHem6/i
MnSPiioFiP8Ql+FOMNDDZjkKok7LA3fklMjN9raEfFUKYLoI5gNS/hwgFCFvg1Jkn0eck+x1e78C
rqma7vOqdOhMmZ1EvyAx6ixSyg+Ka7kAxOZ9lss42HonhVqzYpx8jEgdnTtS6az0Vc1e4PeIOF0D
8BSs3uagCTUrrEstNkMCN75pXTF5srBs5LNPsPy0x7xA5rsqSIniF9kNha1HonIAPlKLiY/Mt6Ol
GaFrH1Ma+DXl76IzHmaHXogR5qbCYyE6PQAf4UNeLtahO0Ks1XyHg9RVXyvrVIjTEzuL6HUjD1Yf
750R6QPIKsGWoj4ZoyjNeM+iSKEaw9QHoPIvMxoOqAL8EaqTCBtDuyEmBKbd4tDPFsDM3l+hviWE
uz557peJy5M+8LIWbFn2EpVd3CuyJxM2er1hxYXbR0cvPe00yU8nWYwqB24lZr7UNgTjy5IMbAkW
r3WalF0LnxApYPszggNzdcjyPg/XqWsgVLRUd/lkqxVA7637xQsx33G9TdnlTuOQ7fTn20+ZgKOX
rY62X9QEmBzYX7aZmINJgW1X/GFwFOMe449p3jlTJTCHBxMo+xwsn3fqOT+aQOwqtj3Hf3vjA77g
Bmrfl65EdKvr0ybH/5axfp+lVGW3lebbPf8redA+FjVkujU2PDiE+0n2w8qsdqUj79mlAINwSk3P
id9BxrXBeqPkPDUVlJRUqOPPowOzZn+xRWEPzW8E2dhnD0GEyziDCbJVpOnCCm44Cx0O7dyz+85Y
rq6vtCoFEDEnNSjB0q6GskcIDipsjywJbOnqF9NmyNIPtFUBLqemNUOO0pBL+WX3dSPJe+a2BElD
JyjAKPSFSVeRbka0S0DoW0/NrBJFV/t1h9LMICPZGC6zSU04rFwi16ijtB0S9k8yJ5ItgEZHnBjK
W4APfaBC75sQh1ZKnVOMKryuTq4UPFbVmKvPOoEHs3M1Ior5tq6kdFmMIo9esE3i+MJHfMhn4fBF
OAfiFsm71ksbLvsRF9PTGCtV6Ew07D+w+I1pICx/p+8hmH+f1Vjik7WZI56xZJ5DnjkfKrrRp9HI
SoDQYmhni7WhboeCbEBtZyNuOOZener8T78MJ5vYtnLi/spxvlHTiixnRtrUog8x8oldokQ6qnp7
6KgXyM8JI3zNiSRdfvAiVXn93lJwnbolUgOr3UgrhHEqC1zkLnqPthmE59vCH3f0BMzYZfcWkJh3
MhcWIptC3MTU4dhCLKRC0HQgA/VAx7g4QCm41/TkX4EoqTwNGfk1pMe5AP7DQ4WpIsuR4nPkqeF1
dJz1Ow/S/FsA23SyFWfaRxqpFgrgFeRSF5YLZHf0Pm7mEJ37rxSULMiox2kSxxRwZEChDO8TKhJh
kRHPJExzePKzQdbJJmBy7X/FN6a/X0YLOFyxI2MC3eNWFMqDuR7FYL8MzyNao+mHtQj1Ct0PkMtF
4uTRfAxvQTh7rTA6TcGCc6Bbs7YzZR0QSVnDZv/fNxC0V3wjebMTciNeF29yFM9ipT8nxeuq5UTs
kICGpY1/QR9lHMQAnSM8YvQq25gS+JHCpZt4+hLgBiFHOYP7bIY3B2WtevReWoDLytw4soY0TAEh
cgBON/aFosoGkTouDRxEpyAp54qeJnHg31G6sEntNDmP9vZBjoOrMG6rGAimBNrzDBs/zfoe/mSi
nVKo6W4ZU7JCu5No/iSffhcoEZEdddIbByVVKizmxf3PuJ1kAMVCRgNMOAqvoUZHEipP/84JoXt/
41v7mwvTK878CKwS43iZ8vyjQzxg6R0yDQuSkjKsBIA2BpDkrGN0xzM7l250AB0g7G8SYib9ecZn
fkAN18e7Tt6j8fl266+Z8/zawJSsA6c+aQ6JLfGUIQhtPpZown7PDeG6TokUC8xJQrtCDlgsSSzP
mtkHf/4OczX6dfK7eF6Ue6njbEeAxEEt5mWnbEsGA3u84py2FoP/ibWbQqpG7MXB8xIeUErq2xuL
Mrn8Ox41T8N0wqeb+VkwBkWmMfVsveD/BaICCZee8/P1zgJOGsV+9OYQhOvDJkmqQUC8IpegYtiX
yTlKTCmAUnnPUhdIutX9vE1IV7XcXkVdTSYXwnwmnzj/gg+GKY89g0PhjcMTywzXeUXXy+piOKuo
7vnmTloufFfHCnJGAF8Y/Q0gSyYI7xMvWVlqEj7tQaYkznYoOC7RUPVf8apAMNkPmVA/X01qfGFF
5Oefw3fgO+iXZ2/ESDg//ZGC/bTVkEhkEvOSKWH396vtE2B0W3dCLRw8Xrxo4Crhas7XZW9CeNkZ
ssi9+9OfHMpJrCeY06XeijUTHNJzc21XZqaQMURDK+drNSOSSsnaKTCwrDJzL3gKA/HhhkeiDFBW
H146FtN+Rwub/z1s70BiWwwdFEmSZmar0UlhMS+HDBRXBLW+zGoYiN5+0evSEKtH1LrScbRDUG+V
kIMLsnDkswV1/LC6HAxjaQy4NWvBn8Tl6eMfaVZrDaDUgWC5/ujaM2qMiHZzyJiixCFEzPNIzshx
vL/BxOfj4lgC5BRh08NPuZGH9PYTEa+JGapqS8JnQJ+VL0tw2zN5fZDZk3Wu2DrjbUEJjLDYDjyw
paLuZqJ2KyQ0oEfdxVLbsjmZQmKoDYpd9VHOtJTXo/nBqv1k9XCC3HhmXeWHnSKlU9IZZgmSk1Y9
N0p6SOzzfD5kdA4p+bvVkaUtu1qe/BWMMG5HE5D7NKG/s3p4YxyB1hzKfbzb94D+yrITDuawPoqA
zSBEC9eirn1LiZb3K8FRM/z4oiHI1WI5hoblOXIWIlEW+rX0j6GTUe06SrE71QYLeTtleXih9jax
0QOKynXWhQmmqQ6WKkhj6hcDkxYthtSCwc2ZOBgHaa0M2HmWH/eC7m+IiDMOJipR0MJKl2UqndwG
3BuJaaNMWj9UY0hDbgSbbxLIPijLCEHy4GOQbnYpK6G75etzmrq3legrW2ke7ThHAnwi2/cM6C5p
Yy5zt7oP4XDf6XOXGoKR4dq7v1/Cvh515//Kd49YT7KAfH3JgXatkuykKrQ9dgIHrCZj5MIeKqIq
btP+xBvKk5cUC2N1ZpnKeWyqGknLb2qW6P0nNerMLJPM15BIq8bkB08NQcg4peb7Di6vXdqhcHtG
po6G/UWOFJzA92TMoQLaM95DbacQDWvy1a/mNbIyoTHcTQtwO0y5G+suI8pMDCJYgVHmBI9Jgj3N
FlbwIBDGeXLW66Llt5SfT6QDe+Oqlbz/6JZMa16HJo1uHuUvsJcOgqSGTzw6BLgk1eSOh0eNC+Hk
KCTVMm3QAG8Isl4sFPQQxkTVMoV1lNpZjmzHI3unWNREsYpesVixkwRp74tKTqD45Hq4Y0wTf/k9
JQG1afj0tMCJr/hgJ4cDv609GukCeMH3Qb+M3UDb8pxwbLj3y1MR9mnMVZKgCZueimXl7N30/9zC
DFXszgVSPJWxqDSdROi91ocOKueZjP4trtVZ/q1Ov5bJvoLPGm1IIGDmjmDdg3HB38dp0Gm543dA
0CwVy82OnMlXWhqSi7uk9QEXVQnpZOnQCIYZiabAjb+Np7DOv2zw9iJ8h7HN7lJDYaAtHT2Lh4m7
8DPM1f61tL7+igNqqErvZUvZxdCTqZtpc1BUMuridr0lVRcvkrwPpnakRmqk7JznX5xfY0NnxWqz
VOhcgzDzd4uuAb9xW+NEZBtctZ9HtghojlLi3OSJ4zPCo6KJ/W/wDmpeGSK+ke4jKKr5qms6MfNk
fAdK1+TvFWfjNXYhhQbpjztwArWPAN5hY2ypz8sLl0gj6vZL9G+yA8/9Js2N0+/4RVBT73dqLI4H
1R6bjcSM8fAumvbSgBdoOs5U4gEBNEscywUPz0fodO5i/c0CpfKrzib2oSOtp3AIDIflOEPKvzHD
UcHuAg1ur176GYwJ7eqq8Yydy9z9ORkKMhyiiSh51HLoSiCEwVi7F35iOMQzOyMM2jyTrGlTOa8R
jOX3dLNtgg/2AlXJMvv4RuJJmMslUjUq3hHwphxYBKBfpkmBSOSEKnpAU/Yd0QgWVSYmgD8ZEgom
SRTgV8o1+ly7cM8dR9Twd0tX+G7vPxy/JmxHFouGoY4lc339zTZkEJV28MmZ12boCYxz6YaQgbTH
IXM98Uzd6K4bNTa9uhYN1rOQtG459/aG5cWMpoqKvSE9WL47MGfsIaEQPlnt45wF3FgdxGf47rsQ
4cE9YwVM9Ec3LAPZSSlFQ5Z4byF37X1LNyWAmexqx+jvLoJZ4hJKADEDLqXZMfLaiB8QOemm08oB
2uz+EVPVDuEggZCE0RwF08YhnpZy6cn5o/rm/RsmCEGIlstQMnCSEGvhTXXQElGWOOYqbvxdGAKE
FPwpdo3uPgxkCodZWxCT1rGTvO7EbeYTzruJUDQ6er+JjTRC5bylB/wTnu4VR7eYRoLT9nDBSDfo
5KSOT5PPNAzT2HfJfhHmcZJvXTRYqCBpFYcctBju5ff0IrETunDARH9UIdiT5094lwvo2Vpg5A54
IbJ1BIUP/6j6pUng8E50dpvnqLYEZkNJ3Ei5ybMmIoWaGwfU5TjytrlPQKklMMeAG6Qp7Ceth39+
dElLD/omKWpLL/xUs3yGySEUBPthb6Ttz6k1McfG/0ypUsDzBxv0wXjMd4KvAOXELJ4bLSgN79D1
a/JATEUtLBTEeFcVRR4JRbL6mH103qG91cRSv7kMuNEbO+VyGbvBoLCDNgUDhL8HCDqoATfrmNXp
y3q7fzif+BuCiSKH6BF1Pho0v5eYgHh/H7UKfvSFopYI1JaZ5twgbcuCwwQiXgZcKLWF0/PmUo9+
ng0Zf0RoGXXb9vTzRXh75+ejBnLg789UpsVC/UU0/1w/Up+DiX7asE4MGl/TXLrp1CD5EvLd4D+Z
w8bfcu3WO0pxf9sDS/na1hnYSq6oGZBzHmgvnCjTGEZ4I5F6x57CM9fXgf8pU53ti8alOv96TVJ6
DMbcClA0vEVz1mGZJRc8mknKwZIcdNHLGsojjpXJXWTpVwKD6gfKEBpWMqQoaHsukIy48/y0F96B
IYN2rPy1s1uBwwlotWzdYfc6qcHrsqjAaRCl0fCEA+YYPcl4JBNDk4bnQHXvucTRNT+o3tK+Nejh
Dr+Nr1hNnnUDiiTyg1t1icAeZM+lf958KtSr9UIs/xo60Mt9g5Xxc79tZEAiGAQwmZB+jX1Jd2WG
2XMwfqsAgpPyUBi/+mqHNpTqyMR86pClOS34wymSml1QAuCfEOfWInq5K+ZbG+PIh8TW//2l79Sa
7luAWDZ8K2xlgPd7G6iEOlkl4yLlKPOT80clskZc06N+WlowJ41Q0lPvo+6QWWWbi0lCoeWBaR+H
9zFZDIa3hvgQ7VQZE4lzmvdDaQMGnWTgowZ3wxDd13kKqzlzHyGNPScJt8Zh9BX2wm5D3/sR/8G2
hQJQgoJua83OfytJxjkg7QqCE3B5G/Ofaexd2Ewg0Ox/lsi9LtsK/B0WtNgswo1cvIVEhVRRMqSD
gJW9DbBJKeZ7XkHspyHR39ynl058r2mmX7uhMCiSM6XAhxzFchmZd75hRgnU8S3xhFthKPA7Ig4p
FXIeE8pZO7ApPIzc+x7TdIGnKApE8E2U7USKpbPD0cRcDiHvBi16tbojYd98EbdJjc/IAQrGs47b
ie2twy4z+9etXZzQ0A01CgwcU2CefQ3saGTcZYORX2xWHGuKSb4Vt1KaOQxli9AvQxDL4FLi/cgI
8DnufAC4JQRtrkzQ5TqKj+/xyRI8xrJqaPh5XCWXRKitbIwR4AvXqVjbsXYK1RDVTgybBe67mvy1
8/Kztv+7cKa+eP4nf8s6jPM2v395p82ZSsl270S43IZGX5bgDiLnj4/S1HDqipQMTuR8tPUvMEpG
jV/Edqu7qFcbGCq76CHyv0yNcFeMC8SC9ADK2eJKcVpFq8RZZaGyzqpFwRI0848inhuPaC7vZr9e
cv+07EdpBzLQQxg7PpRDYDiJdfItNr1jBKrZV9kQ/m/a3QDWcetflx8CIFOquSQt6x/1YJlFvDHS
8ILxE353kdeo1EJOE75xwSCQwiR/DjyKM9RPu1ZwNYMvNd8v40pUBZoYPVcIZNlyb5FDQm8YCvof
PbPWAdvyeatH9dWz6MeaNp3PofJa98/CcRU5U69/RP0FiqK+DlCtwEf8W7MFHJlcy6FQRE34pqW4
9dgulL/BXm5jJ3wn+wLo2Hyje7aP0Y2vA/5UsXWbD4YKmkzXPvK/F8WXUImrPBLFAZPTeChJ8OXE
imYutdyhE3gPYl/9ekMjmsP6E/pFrp7W9WKNMLJxSncljMkknL7zzrVVMYUezNTXbFJsfpNCQ12E
g2rk7+CsYzTMMPCvGvjM40QewYR0xkcjd+lrZZIqoJRvRqjPusPbhLMe6KcxGdM7IUgolS/mK2i0
yMM3tUmiemJ9xZb74+ebvFydxMKEKB3mwf9MkpwdEsDLQtnfTUUIIqHKuf0qhIhHlW4T4YQtRCqN
V6QyGexHQHyaiAuuFJNAzM1ObDHkl9w5wU5OLG6Hc/nQ53WsA5uf3DmktC9hKGnIDuowrhJOQAsy
1qO5TuV4510yUYJGMlODIe+S6LJTpU8KA5nXTbGZHTkyjM8rGbd2pCw5LSQu92NkUeGlsg0bb9HV
e4dTskj02dY+kWIlGeR4/8aN9AnuQ+VXHgihIWcOIbr2PtYes9dp3/5LSxcR72O7Hj1uC1vEDY0G
lSbQNT4zTW4kesOCRff5m9IOjlnE8OibON2KTmEP++SmAZ5r6+HH77yebh6CrQykDdZjHlwoJzQy
vNpf2IY0wJrXxyjlEm0eT0q63UCACI0RoH+dwxAB4Na/T+bM63x0/Y/A4tv069JHZZ9zMflVrSr0
RKjlYvmOD1mfCbw1E7OgXPHAoqcB16Au5+Do9zAZOYi1xcsVgI65nihE/a9cM5BmBbBBOx1P85oJ
J//406sVK+XrDPL3vRZJdXnWaOYuZAnotNVmfMPRnD2urrAFZwYou8iLT5zXyFzXvY4mIaW5UpcB
5WYyAcRWvULcC1hLHWs9XqbH7aJwTWOTGWpCwKWgHAJwOusLfNB7OrMKcu9IZ7NQ57GTkQw3R+LP
5k+F2wcjiPHt8C4wCQpaWYDgZURhCdh1F/P+bB0I+YkxJzvuXy3SHppVmr0vLarEzCZergwp0p7/
Mh+WyiSnyNnk6zCd2gAo4ixpPA85xIrK0yQAQaKdCgkgHmTeHzH23fF2cS2Mt9gxFLkpRSUFn4gy
ldU4HGt40hfrMHABOwTC6iv44Dh4N+9sc1N3NCXWyciKaNM4OcxRQRQDvVG83E61pAGe1pDUsnit
1CMpcdHNJxPkG9De7VkQrkKwiwNrTzk1E+r83bwcmD7gNIEdJ/9gmwHr+KN5/HxuLeepdWDJruLG
OFG8/1337EROkqEGsM9WLzVDvOhUqZa67kS/WRFyGUkvu5EWWqP1AoyYpk6g4ZwKdXk72myHBVDJ
TnN+zi33w0kCJ6BXqFfGsBRFQ1moZb12jU0IMRPwCjqw5TVWmDJ4Y8s4JBm6Kr0mZo60DTIKw7TO
Kzf1890XMWujNKb5aUI1vgczjVZlXFM6Lg+UzcaZg9yMYx/gzduiuzH/EMJ+F7VXn7pKFMYuoxJc
RP5hLzDzGqTMk9H7hyk+9N/p79HV5NbIiMdC87AoDI52hisX+9S2CPVNWPj+yaSAImowCEq99Kqm
WmMXaT+edYo2S9xk1/nWr3SM1hZdZFlwJREcGtNo6g7ayQyyPzNvgRXnUIfaE4uoKZZp2lI2uVqL
Jfzg6ckNOgyuZ0wyFW6KdqfxKq/mAvwZDB3bw/adH3S21KLm4lQeTROE3aORaSw4oX8DdTvHbUZ6
cDuAit/eVXfsgPnq9H3SNItDPX+oStqigDQlU1RGCcCJ1LXV11lQrs3e3EBoat1yqUreqPE7eoHP
oaFHqAnS7T9UWA4l6VaFWosEfozRlZA47o8OlDk3EmGMxmr+KhEOGwQOFA5cphF7Oj3C2QdYOuzq
Z0BpU3v04zOVJwGIS3Jj9rAtCxt2M6fGRNCQJtqz3x9s90MVk5XoMVg67BPRE/Lx96nZ6IB49uNv
64HeazuYEikgfLJNQS4/q/x3Fo64EDrQwc16oN7IRRA+CUnSPy74ueuWVokzo8KHOQ0Ly/LFMosC
H69Lcl4uHxApOIoTGIZ2T2mGGwH8c6zPZij33csMiV+mon4E8R6aaVCo3qWx2y3wYuStV09NK6dN
CSTJnNgL89qNiC2BZQHYwLxK9Ioc0CejSCzuixRB89e/f7FLRlLYGnXCrCGWQLqlmp5BQjDC4kIG
UUW4LpJiyeTpTmUtH7BaLkGUCcq/Raz4QwP7NXH8lpZKxu5HGvjdSNB+rcdbiy3bpPTjl96h9hbg
PfGf13ibHvvSAt8ZunSH7hIzp8wMsIDO5/iUCgVlykKovj23f+iJQqLfLFEVYaL6c0ju5Hk446QW
lS2syMug4L9WMdFfZYon/jZMqkXPhismLob6favbIiIZ9aTCK8hEB8JNXd09GxFsnqJfvkIYcFjO
ruJBZUXngWa+RYAX6uJfRCrFsvwutJRVAHnbero9ECIRtMCaAZrNNMLKXaZyIZXH3UIe2tKbQOXD
xe6mYfc02S80Eszrg6SPq6dv/5F+HS5AgfAwY+3IkKuRjT/KuU5oDTrTTlKbX5CBf+0BgpHAZuJV
1rafyBUnRIkXqoDUaz1i6w8yFsAzch5xka6kwFRLTjY1Wu8VKBVEz0CZjNkx3AWrpuUroW3yqZFB
kUnhFxvHSiiPw6cMy8I0ephFT+GjYc661fVBtmZz6Z1lv0XpWzJ5+6Ja7+f97SKbwRNUEsIDQxMt
1joME6rDD3D5Wzq/XSiM6Gq19oHD25XVzkZRMzAei3d9tO4odiU+4xHm9Jtiua8PXpCO4ilPJ7aS
+TU86XjAonw7b7wh/g02SIGE12vubJHYKW8U0pi+zZyxGn7SESG9HlY4WFi1kA3Zxs0araAhW4La
rp3zLWdnzi9v4u1neJr1zWNAzI2K9kCezsIJB4YM3RKQdaGUUFzSAjFYp9DlqrnIWI/VO6Bcnw/C
JPlSAmAuiwRRi+soyE5Krns4/enuNN7Maj82hoDtYaqwgnr/736yAoSEsiAug0NqJDaN8x5ClNm+
ySuiBeQZDl5rRrkF/HGGY8HOzDhhqD/Ohadpo5xBf24Fiwh4/WIm/03u+Su51gZz1XRbNa5rkXjH
jOqwH40Ev2Qh+B56Q7nt3Bf8HJUQ04yz1e+CnuENJxvGmJHVG1Elo0NXWaNN0xL8fIoG+bLMsj60
2vFkWOQJDAhJTtWJ/0hKJyPtpfEqwoOIRy9I0jD1bHpLZz3HHbsbLctoSunr7R2oQsSIdRmZdZdE
wlu0T4bgHghDmxbHj6O5/MkLYF1lLmDAxwLZ7IRONGCkeeBgaoANgt/nUcs1ryj679AQSfWRO1VR
iPxl/rWgzdT6DQhCF6JbjoCOpw75CeRROPxKPtZ335RfAJOtoh4iteb0PyT8mAk+z+dZ44zpT860
eGZWsrb6tNHdx6ufhpMBOn8rHRxIuM2rNpFOYZmg00n760ItJ8zzDGS6VMDOBlVqe1jQGRLHSfU6
489Q02AyZYKIQTicAhjMywZxi0PlwY1J2BQqv1f+gWkgSYlon6FDBXkOZcf0Bzys7IyzrMkkMv/g
DVu0QE+9FAafqofjaVpGK5JSl/HpoTvoHh8fzsZwrzua12+rNHC3PzC3evQ13w/IbKYhHpSOOsij
nZZt8wC2Vs9F4j48W5WQwFIIyU61DQJxpbBc+7U4aAKCdQtu1rc8ABChbt3k36S8oifTdcqCpooE
mKNg/VQEGSaNNjdE/jiGcOwSnxuvTNtjKDxvPdZvDo4EYig7goiqA49xZUzC5e+P6pzRAbdUWbGT
G+b9cAIEAirtm1eCTzfKGZDpdBP6Okn0yd1k8C8NdeGmkjbEhtjncHNaijBbSrT1BjbV7qgrgkbk
qmUuaaQy4FDYbm1HQYfY1za235BU9gTJUGfrX2HUQAaSJ2dKlmXHdPL2qFSvgVi7HAbUNj6h+lUV
V8yynU0z398JTM6uKeEuAHa4tnHgsrpiMwMsfHEWDh8sN7GOjNja2IqC4OxBPRfRqTpWGlXZ2Oot
FNTg4aKDYOHfxAzw++AIftn0DrsyVD0oxrultgatWKST6KKHsJgB9oProhe0xXsF88DkAZI41hqk
Y4cTchPQtfWf8HdZ29OrkxKB3N4+FE9xDbqW2GpZNG0pX4WhuRrHnWU60DAcIxjQ49Oxf7w+RGBH
gJX1sMq5qGzdDhwSHpX0RQ7hGXCG/PfA71RI/VUcI3/FYgm2QVXzT8+3wKczwWcU7h6qPHzeJfuQ
YXjDQYm+qsXgUmLqIGIoX2OsJ6kbmUMAHtPCImLPSB+WjOGKqJG5ZlxDfFfLxgJZr8pIeFC+YHZx
zLUcL1zBivAaneS0cdMmIHLEQQ9TTelrSgNpY6vJU+nNpGxMmMqJrcGB3AkaObpIisp4js9ydzv7
ds+h59e8F3mSjVeaz9JIac3Q+2H8BdcLCMgxHD0Fd3wbWF/QZD/PhlqrDWICENAtPJy2c1S3LtSI
gS3iVyNEBameXiPZp0fu7d++hZToUOLjQsrRmD5E4pwlGpe9boaiHa4spKYdj8XAv1R+q+zEbIww
9XuJQWjldMjHwh9LoBoWfq+Psj3KMX/prp/NlryEbd8GnZRty7UT9vGlElIHcF7jWEtjmHWl9iZF
tDls8ygqI6XgKpS6kGw3QrBNxqGXucBfnDis/zsojCTyf3I7UOXcCUg/8g0EAmOzUn+ZLl3UrSFa
5jMjuRFamalGzAPfTVBEIEmL3QldV/orqpFVueP6AnA6fryyJvcYbR/rTQ2p7OH9bKbguhUDgdpU
jGKurWzOEvD1Rq3M6iCHAyr48QptXZb8qx/n2vS2xsT84no4tmcWAkv+tPrAar4vuBCbx0vrqu7u
uxSUlAUXH2GogD1ZufkcbzDGAotJjLCBdGk6Eg4KcILhjqc18rMSGBrCB9P5C9SNClMudj5yt+K8
iSmvsyryTjGCv3OHV7q4qkqmfht7o5DFLRmh4lHWoXncXpkkLYouLeLovixcfOEKW9uVPkOZpcc6
iipTUME3K97Q58/rbFr+73wgsydpAOY9StT4uwTk+uYi4ZDy7hGltldY2LSL1kafjor961in7Twh
x9DmJiF/Vr7Nb+/kGuHmunacnu8NvvdyujPiqEIa1XUMiycrnhgn+EeyEwPHN8S9YVrcPIdWeBkS
L1OkrilSqz7TJBxgK/xoecOFYsl8BHnG7uh+GqQ0Fjz6u6YcHlGucQqw/EQ7v1g7/WZRm72BAQdp
m1v8FB5ICl8cKDGDlkmDNXv39VNpFYXBKzBfF/Y+x+roEDdkv97yAmya4Bg1zwvebwQyVCqkbMCl
YcM+/GNgrYKzxxd5xo2EQtbaybmqN8XBDO7TV/vbXXlzrBdpWCb5gUrzcpDinDLvOq6tfCEomCbM
JNA0pKWavlVuUCQ7eaj8kOGxGIUPc7RfWG/y+BGZhW1+0ESSYLhFUN4/5sAsrsDhPoHz7lUj7CPp
DbcHVPoUsK3N+s/9o0jHx31Oprsay+da4qE3+WOZ6XFR3CRjn3oOrfkQcfdjlYjp+52kN0+tgvQq
mANzelYcX5mh8WrMmhlXROOF2UnEYFOu2zEtbj6sVkOVYMP2XabFXUM1TozwEzS67ivVcRaHNHzu
ye4l24PaKpAU/5Ja7HXcLeGv77kRSDPr9p6yygwIYtm3rYNSxaJDqTS9d3dTq//iT7VRZBnmAGyS
D5IVx/UCIJpoBjOHpGCQAP4uSehP/KVi3kRU0D6ivw0YgoU32vI5++E6jsO9DS8bERVQEObp8lhn
fmeHHiOJ7Uq7o8LFlOcitQUd5oRtlkNmyRCWxnGAjrc0dDcTu0+l8PZHbunCfmKMDY1u74OCKuMD
H798lP+bvKDLteuI1z0SRHTZ+OZysmIZemvCp7hwpPkPk505rWdOrsh+AkREF6J515XnMKbcd7GK
W2oXVmm1lz+8z2kg2/SQG+YseSxzLwFljblcZAj8wdBylUxMHyHKIhGYbZbJryzM/a6MbvXCT3MV
O77nHS3CInLbP83d3TRIipHYuNN22CpEF1qsvDn+kmrySFzEDJJqfc2W59zvF0tkJSmsu444/O8j
IhvLSzZisISzc1I18vf3LA7b6PsPcCvkB0thbZVrUNCdRlUTCZtpglcg6elOOsXWR3V0DrIDo7wM
Omjvo2VSvHQ9h7uc5QUYByY7h1cczuJbN/BIO5U9I3Vjfbjh7pPNQOBPbeGtPtJvHo6h225ROJum
eTtHKDGiHlgkYN+lBlHIxZjtxGc0CtbRzO/uKp0KKXHbJODmmzNaBtCHBg+5mqMWwr5H4bQf+Vh8
RysvZMkpxCjJURRM3OB71bu4yVFYOrSLethFl2Ms5Fhk2nDOerF+va7VSIMeIMkZ6ld9nsrhg+kK
f29hD5WCF3Xs8qV5y1w27xtdmJJ86HTcEdAmaBzALaL0Z/Yfm+G1kxGQqYigt17w9ql8ApnEWON3
g/RRbWqFsEVlXbTdF7Bs8XpemZJoBM2dPjvDSu+CIbGQVetaXKAt9vudsrhAmw01LpxzUcnR3DB0
+8mpFUCI750GJ0sZRdUoMG2918MvaIORsT4HJLmzSAj9EuqCP4EgOt1bCBABodvNhxOE9qGQpjNN
CQMUUYPHDmVImkIvhNxQi9aoRjOh5WTfecSSXi5Rb39WRtQYn/berYXvXYKHwc1UD/lEXC2dhFQj
fUNSGWpvnFOd+PZ3oh5KBIngzzSVUxf+aRAYGrQlQrWPOQSPdHCIaXGN5yEgR2bVLHdtXwcuYQVL
wjgMnykORsVRqVpbQiplrDApn4pWqscULwtfoQ/KXY5I6OpBAXCVWisesr26g98vYcaQyqoPfDUC
yquDF0gXEAhpzzQLQRvMTTGfA/D/tSvVEX4qfIHkeUbbkEFY3JciHKE2JokYM0CuMGXkfkp8pIo6
nKsxcGR65tqzox4oKWl17MalQ8lc0wWKiVPb1xeT00m8h3OUNYh0DGIos+8k5+66j9KqVVSeN5Oc
vkavtDOPUR9Zn3Jer0ccK08eQe3ECi/6ZG1148Z7D1DT9eBds+cNtBmY9gCIVV8Yrn+Zwttwc40K
+bhtKvxet/XeN+HGOGzWjYjdBFUf6ESqFXLd2h4a2KCCEaaWVhBM3SP/+ARtv4ZAaGyQXCLF5BOc
DOfyapeUbmVnmMIZAETIzBL0EgZlvAFTYFosK7JmNGeKNMcv8xWQVwLCVudH4Gfc6I0+EFgdsYD/
8M0J9jdU3iqO3dMvlN0ZhkcJCiPkE4KPZbRNOKcxxM8o9crfXcXwaf2cfdFCQ6KwpFUDsg3OkIPU
oJ5KXKGoyZpLJEoe0SoA92all5c5qz/K3dGmaX6k0BC/HgkuvEq5xCKyiNT6sBlQt9sSo8ULN9Uh
McddDiLTXEnZC1WZiQ8OjtJxk6h8ad/cOpV1r5FZ4He0Dimkf8qnU9p4f8FEg7P8MRCBsjBgJovP
4nKFPPIEbzhKDrt/F71GPV0K0bSREv9/e6D78N4ktvMK/6LhM+nnxXwjfCvsKpPjQM7N6wNWqtnY
nhtCPeWImh5gvAVZebCVoEaKucy1/y80tWMLbLMLqZGMS5LQtSxpMde9JOEQb6EJeKnb79CjMFrz
hieNoEexx60pRnPCCBtUGFISSBXfodZp+P8x0jt+c5SzCpxm5hgar9/UMu1bYiu7FwIYaHwtDYSZ
o9FiLaCz//+qDfPH28s5R9iaXEoxiBKICRXcy41xNwBQGqh1CNf3942REamTArqEVfiVgKDM5avi
fnJvIb7F6tXfXzWGl9Bx4EvzkxeTQuY2FL7FfLCPRCKtZxsIKkXaCCUFbqAI2RzyEXLT/yredq/i
4AlbmLBH8I7M+ruSTHzZfVrqA48qIPIjwWa6QLYICPfRBshov8w2dbPLpIuxM3q7E5S/YcES5pUQ
QJ0dL9SeCnOLJVZ7RG/ush60o1iZvPTWDBDyOOhOMEWHa+U9IMHt+e6/hgRauyBs34U54o+IzLrs
GEmZ+wOysEWDRqXMZGFdDEGIn0CJp5q3yInwYinRpmXF1LGES6rutK4jw6h0rBnmh0xYncYRPTga
oQj7TKVVJqL1iBezXu9I5pcayquzo2gWXhxvrveW8eIrvqQ/llU5EqApfG+GUjnP8igKWkRZ9Gaq
e7EOxed/r4PNWXi/q6xe1SnybEb1+UC+vcdR+dPgyG/WT4tdLsFnmsydmkr6d1MZGveBlL0UJbta
lpLxJBXpyInG5Su6IJlPdkOD8UubMNC9MJYyB+jowE0TZQNkPudYoe1TSPLRuu7H0jdqLmGgKzzD
KHY6hME8Q4rDBzzYMoY4nDHHwNPpkf/qw2weXpbTqRnYseyHUFrscReIvCUNf0e4ABd5gJ0MezGr
W50Pt0iKGlGk850pKK8Xcy36j1mDGEG8geXWbIG35ALdgCcoUCHLrtdVJ7IlUWJ1TtjpwC/UY7k8
Dqj7QElRAhjd+63PDbaUWO0+EVsOaduckdH7xeuVODAzTf4qtn9Zv3HPXT3xZ5fI+8zmp00sMuTq
h/YR7l32TPb8XyeY08NOoiIBkL4AbeMFvpV/9fadzWqrdfECJhP3BGMcb7c8mVHQ/COOt1cHde+J
6ptoFYCY5myTEJKTwZizwJnXfvIz3hQ9gygYbVwI8wZh5aWdkCmIlTl4j4nkESlPJKwzlg1aIpls
nMJICFuoxvtZhCE7v96PmqnNClo+i1l7/s476EZM7XfAe2zlrt5SSeXzN005qR7NV4LEdm9xlvZW
54OSLjbUnRwd30BE62HGUBcH3JTPz3s9KSRTXO/lqmpy2r4ht9SYwxP8Y0JxDpl8UDVUnzDcLhxQ
F17N5lu2JQh5uiiwYvbpJgh10MxEjiyHpiyd8jAmeNTFsKreSMV8N4v5Dfud1wdrifkuLAaTlmKm
PIw2PG59mlJjDjt9kZcCg+Zyg9wR1rGI6Gu3SXbeeBz+ln/DJ5zChjty6yYkPrDJA+LuICleLdcn
KVGXMubQ7pyJmPakh6f04k858tBq+7+kEV7OUsuJfYffDRygNNDeMroVj4JuaeP/hr8M71QeVyDx
aey4fcoST0GDM6sH7g8I/5gu7NCX5k9XiwoXtwI7nu4gkfT5bnwCb64HoqObqUgnvWeqqASAyV+3
QN3iW9D8raYcXhuk0ZWcREaJ2NWHytr3zvotdVAygBw6BEVPYpb58BlbFx718q1YpnbbIPNG1Kvw
UiJ68gxgBZxMXl8j+t2M5lcztxXS50f5vsmrirvR4TcWW7N1g120KjGpa0Qg+sPaOtAcUGekHD9E
CMtA29H3JaB8smi2SxmRGtgcnLbsisZ9JxLyAflvX9xiFm2h7fTJ99Hl57rP6rewotJ5pX0VBvna
HrwfZl8M5A4NsFsg1fqxbBYaUtkZSPLDG880Ki3O8KwqYeR70wVQhY6dygmp8RG3kJ9t6EGo5KIM
CnBk/bIs9E/iY1ZJU3OM2riVl+7bT7AE8tKwFfT0IerN0zFpJ7Kw0cAuRD/b2N/hfTs8O/X/c+uv
Ebrct6eWTf7EEqRCFuDoMgw2zQx+/0fqe0tzGjS24rBzxLiwCgY7ojuV6tWsMOlc7Dhwov1OITT5
pFL/9KCkGA1NHU77pmvhFj50RNYJ/ClwvvvYXP7BWdkG/siBJ9Byoni3ZFzz+Y/4vzuqIhkxKFtM
8pXMGYcrTIFW6tN3BvQxTK41jxj0bxCeTT2CjyXZFtm1tCTwAfNR0pBxDHUrLX/qwSjQUB5cTstp
VRt5yZ0wGSw00UphuCqcWQIiLTfVOMn9b+0a1GjCh7OmEkh0K69uORaem52Z6S7svLV1nF1765VR
oxyd5kL1ahYP+M70i60hqdxofgXYPAt4J7VML6Cr2PWhUrf4ruMahyJyjx/yW5Or5U2zV13a3lX4
Ld0STssuuDowwVEvp3ZJSDPrPCZAczw+36B5ogXIv0JTBSkYwzWHAFrnDrNSibEGF1gFQhJwmlTX
8uwjVgCxfIwWv9R6gjrCX6gOeBjeHVPROJzbP1NPKXADScq1lecl9n7ZollpmlCZA5i/6BS1nAaW
8QK0RZThOgpJfYfyH0bFz6hQ0EcOMMsA1yU2yv0uvID+q4vaGcjwZ1o/rRfP3VlojJ4WG8qwWqjq
soX25g9tPMcqHqIZGqtlnZqGQSSm7/7HChV92eB0I0tIDRjIOsCbZbwdAZJzSZwptchOPTNIWotU
YUU9rV3SLzszcMdS+jbDD10dBjiTkuJ2q2lgUKNKCt5Xv9Ye5NRa3lREObZUKF5I+/7OKyawooMl
YGfw/GCZt3l8NWZ8sgWxi8OQA9AhQMSKOamjvx5Bd3vlK/DX4WsT7w5JdE8ZzkBINIb62KUXrzLm
QTQFMYmCsuTJii3dgo+XxSNHZyZ4dA2ZwFyfz3jVtyJKOIQkMLjKUu35R1TyzgvB4c9zeEuz1LZX
I1Dxe4pZxNAIXkvGhPwVD671Zef6H1VTd8SE301/6eyCtROzifVeSNht8D08w7CIlsWNiJfzH3SJ
BMJfeptSTXq/u0cq7ScSMJL4ARwyo61+i/JLwsqvfxVu4H9SmkE5ruNZaoMXrjz1I8EPoSivBVuz
D53Z8dyselkAVC6OSwcMwQm8t78+XRikKX+UIqR6ljMKaRRDpsV1oSwir8sBuPhsnggmCBVW+unH
vOOMXbeexu46PzYcwJ4lB/FkAZZKUwrJ+PSJpviytWIKNoqJa+GWwOugbziY0MveBn1kkWUz5TXM
DLjQuiLA6tshL3j+duI5Kjp56satAH9BwlVH+uxX6/OWEy+1fdbp63uXQ/IKls6xxHrXrxUUcOX8
F6nf4SslnI+hD0A4WxUTKCFkUleppYH742dmmaFFb3Dismwu6D0Hw0dtxwlzfGCh1wH2+WpwoWkP
Wkn0Ft6VIvaCTXJuZ6DG3aW9LTqUy+aZmI9e3ZTfpbhD0D1Nq++C6S9O87a5kWQMs4J6Ae88bV36
LoYkMz07NKA4nms0fYm3EGyuQH2jXg2+QM51nvgt1d5X3mc3aNRnjw071N/QY2cD++2Mph+M9ECy
9HojTSJUunfYEnoY3IgegCevRRqC4ROLr+4TSTac9wHYknJhyfKp8O2V2sgyG3dmpTK4DFWbquch
NqmyP746Eo6S/4Gv90TGFwdU3xU4aego6imeHmkaZV68cYfZx/fjUXXo5WmnVKq47t+29f0Ob0Nr
h+jXTW3vDbBn4kz5Gc0wiTF1nyqdsOPnLcYZwKygUaB3FFVLFR1Su6H0YCs4iewYQMPi/4n/XNwV
A8ETrauYGt9kcp44WqcJyuoCKb3N2NwEa1h8vbG+0nxogrbZT+z8Ss5WbIaRV0Cedf1cxYH657sI
xcP3U8glqTlU7GRqcAkYFVdcBmNLrgTjELRxGSs1Pyk7Z57AXnctVwJjmaqaZZz3fIFTryLhUwzd
q4MrZHlMoVGp4Yop44ZlrRjVZrolyt67nYA5e1MAoOdEjTnuLSyODKrDNesPr/7yaLKtpEeF1LXV
TmIEfXXFzRJaF/hxs1uQfLttN4K2eiz15wFQi4i0wQvtKso9tn1ks6Tqsmywyy0ty52ZI0WG5CL4
D+1h9ibx5goqJKNpjhx5FkUAYQ9bj127NfWI0eBeIt9Try8DbBuwG5kwSvLVoVRGwFmIc61Tg/U6
Xpk03bDLlM+A8GCV94aHWHohLtvnmbzBbHfCXiNoo1ma64O0GtLhTN2TYNLPvSB0bl5OE3KEyX4y
d7hR7miqCsfPavB9ZfqcQtkMeUimeIhDl5VCzle8NGe4cRZKj79XYxHYIeL9W0FkVUxGLMi1/xT/
t1sLJiALudR5LHZ+Nu+HHStE5nLkU5z0zbok+Nf0oN9DFh5oJMlztGZHbjzF6HhiWYTmFtBvMh53
/cLfdtvwJxjcndN3Y+3Qq1t2p8s36DYGlOQTfyYxlgUIbLEPAiW37acur8XG2/8nA8Ux7hfs6hw+
zs5B8iwzCGkiVMScVCmvuFfiBKV+C0EMwss21DKctub5KlDzolekYFURp8BvDhA01Az3YavF1yRw
MQarH7i97v227trebxqkNvX2nV3UXEtkVs8XzqSoxeHg5ULzJN+Iyjq+h+pp7l1H14zJfNrj6dEA
aJlft1zQBfnBxy7oqUFp9xEwBWGl4GdX92GZc9ySHDAFQJ6YsTzaZWtVdHb4RbbfufiT9QGR/ekK
omVF9dR44za08abSbPknSd7ZXnpCNcnZMrnnmNTiPf4eij22mODKHa9LRY4JoY65MMoM93W/GOss
CyAZuEYVxCgIj48+4aas6hTPPXL4tqqeD7e8SaXsA6L+9TqIJ58deEoFtQzTOrFIAAZWPNg0er0X
dxJCretKp53KmagjULyc44anlwmCmrD4wEuXiu4GTdenRy0yPxa1kOIAnJg364HhvUcN1KEK+H9c
ekPGsnKmITosY/ntT50/oiwzp2N4uHAKcPju1t7d/2CZZ42lyHfJAsf6ukeCL4T2n6zTo8hmNjCO
aQIK36Z8uoqetEsHe54iq4ja+6WLtdrMPEFkS9Fto1qQkBHtrT1KvsIt2Vxh0LHg2XBoIk40k/6L
uTWlV6T/SeidXkypgVj49rL39rPZTpm3anF6TPhfJ9DTmkdSuJ7SOVhpchBaEXZiMJfqqGWYTcj6
cYBPX0v7COo0mjpbujtwkTqzTzyolWVAG+6kZatryTfCyCI4HvHb8gn0E4QGXSf0Km9oAvZllbJi
c/LGSitTxXJRf4YIWsYWVY+yUFyHfPToFYizMXuqmVR/PX02B3KmRcASGp1Ds5RTX7Vauk/OtYfA
SZejeOFJxX2yY6Fk8TGq6PzVRbm3zFZ+psU2pqWu/HIlEZf3QvyLtumbypSrgGe+MhzbK4D74gQU
jweoXqvS0nOJRIh/J9lkxCYQA4uJyfGLtZUNB7vrOwDGcMJrZ6tSGoUL+LLEGyCaHzgUv0eiwSO9
dIWMn5QVbJIbGpXFhHUkchp8IbDlcyJS8+3DuvP+OUdfl7L4pqvhHQUs8X63et4ZS/1qyuF4Hsag
uO8s94I+22JCbafyje+JdLFQINozFVyIV9LcfLw3h9hMfHlr/e62ETRIdeDvTdXnr6yKZpwJJ2z0
SghB8xHQIKt7O6wB+pxOlM6XaPPLyjy76qSa3oGPFQeaayu8wQvMqhYrVg/Rfmbewg9VP/9kaO49
nEOuW/sVcy2y+AjRWkdHJQJXyOeqDLhUMvnGPPkLJca3qvmOTKUoR4kft7hkzVNQVkPZcwkFJSE3
JHm74cXSP1q15xiVrQSF8ZUoiUuqs5SWyx7BUSePwqB0DSNC0eZgQ3fAQi8Xeha0tXd4UdyqD4d2
Z0CKXpIQevwsOUgoewYZIfoj3qBVSODE/eFufqTlNmXCumpgXBA//qilKQ3MCU8/kizCTaaeW5O4
gEUuXQt/FbnVlDbmGmFbuAJrSMTvvjIBUAkvcnHkiUpLV24WNp3V+T2iZ2x7rCT5o4r01bZxcw8e
P2we+o9gl+Bs37DiSSH+3QaU/coSB2uYQq6t/NQoaof4awjTQRATXLAyzaMRHkk9LEs9sVl2V9Ir
OjvBLvCaa+xLuJFVs/TSupH6o3I38a948gvJrASXahizX0h7IGNwx5bLwShtq+qRYVapTF1MwIYZ
R34Cb6t7D7aAZEo+9uo7Ck+lyy2D/h27MoE4+OdI8BTD6Jbt5Br22AgpE6ThJ7mmWzqtc6cefQJM
qFlNx5rV/MEg4P3OmdYIWG+VrITM4nzyyXTtCvrFTq5TZI53+my7jtUlRq+zgv9kYux7izbKQenK
Aemf7Zzvqm1wQJIaTsj2GuCjtQ/1Y+dPwNenJWy122mGdxXUndWy+QWqrz1zuJCb3DjAHqGY59w2
zL1Pm9NVm+AoCoGmsVuSvC6uWg6esUeEZYyC5ah4M6Y34AnBl1Ipak3vGckwI5BBXaX5Nspec5rd
s3z28/JE/WBq698njE3wU/3O92aFkJoMxLbImgivYT4wb/V8CuLc3qyUGiu8GniTRIdXhJBRlMS7
DU7tGzYpGZ9FFZORF74NxKhzhuQS4rkPtAQogQ87qiQtnhu6Sj7ujzZEOfXpUzmfa+VqHHdiW/AC
gqEVIZurvy8IeeRcsRYyQUY5dozTVnnC583EVDtNef+2YmWS4BrpA74xW/9rAk3xB1XGp4eLtXly
9rAWlruEyFd9yQa3YQdXso10viklV7SlAcQCJ8yVXcYHUvVHAkDOGWI+UKhnlS14E/abNydsKhEy
TU6aZHne6ZoxD0uLi5fM5nofrF94tcwR7FtZXdXDXrrP/BBRiVQtA0Sxrqshc4wZw64UAWk9TF/K
5HCHcGOYN6gSAgy5VDpvyYVeMayxoTAMkDJnvld9VNoNRkPbWExaTmVCpOzmGWqdxXWhUISs9yBx
kYYhLPEDfiB4liKI0ahPGaRteNyfZfjSdh+H02fnQvlhma9/uXGravrnY6tlaLUTDNR1t7xHYIf8
X0N1ZQLOn3g6BmURXLfZ0n8CUs0ct2aKnHBGPepnqkyDRl07GssqyrXPvFHt0vWuDoz6s9/r5HFm
SWYYMFpPqmdpgcIw0V9hqznp8sjZABVLkbnuXHWFmMfJ/sANukS5c/8csQ20G5ba6FQ9M68vUR2b
guUGEgN8F9amF845z2c9De/jndsodXwfejEe5qw3iW/GyqQVSjQoHsM4k4BoSWIHEz18H70MNa4Z
Q0DZ3yQLT6fVe3YLF8vbEqO460CqoktOC0odFpnw8KrM8tIZScQfkjvlcVj+70w/5iL5cWjwMhNC
aE6SuxiElXxINsVivuFUusrrv1k2Xg049iFIKmlxziojDPi4be4F48NawYiM1Yuw6swKJfVtQj8+
eyjTlSZm6fMaYA5JrlaMiMS18ajzuWXq1P3AX/Cs+BkOZElsmymEQRxsFwaBthCOl4miWvYCNlyb
jlont2HEh5iCOziny3g3cIssjNUpFR8+NwZ2nN8zb2otm1mX91+EkFAu1iNwlXCd1XTKvsimpAN7
XP+MQsbiMX1d+RYK+Ohbp1+a4L68+7xLJDZe+ES+v6M7RNeG29UT17ZFbFnzQTcAvc7gYQsMV6X8
y8V71Pu5txc5mRfhjM6ulcXjSSJ07DP+Hkej2yPLDalICweI8xGGhTVX8ZAcUYVPJHCejo9o70YA
olrgrGRlOQwsArjw9slgMOB+EF+xVFlky7svQr4Q43YktPTPt4rEtkKyzdmmRQamQmDnZXcwEWN3
AvMXZh1/EDEYbnNY0XM4hJxG8lzMCoun9aKe6MPqdonRetJyKAXs7M6qEe+eXbnJyA9MKz4ey53T
hxlc9M2ptNeOy8us+E6F9TtWB8ECrpisKkti9EwJmxRt2KszAwm93NqyMR2ASbfSs84+kJtoiCQL
iDUm+cv83BK/aJ9vzS2Oruzge6a10vLPCi/K5rrb99vYJhmKbDwhVzKntz8bMfd86s73b+x+cqlc
eaXmOX+vEAZLFdwpJa8/2efZ2/C8FeVbjW2nNjk7iSJ6OqMNZcaTr2nQ8u09x1gC075kwhOZ7f77
Id2XecPYujXovuAUaZ5SHQg/Mfc3ilM0/17eZebCNOgfzdVXiciZB/Gyb9ipR2kozGcDuEc4t1nS
jklXVkstj7sOkALSSxUCyPOZ+u/jJm3ERZcBPBFrvYlRdLytM7PJXjSA1oKMCkMCJiJ0NLZgPR0O
JmfW28XYzfzl28pNy6aWAc7Vhb/tSRVbFsEuOLXcniBN8BBurCN1yKGfPi1ZyEL8slE5RysickFR
nbRWZeI2nL38V+4SHXedScH6BSl0+UsPVwTlEdGp7/wjs7InFxpz3CSSGlLzDkHx1awFfFOQ+faD
Y2RFqk/ij3hb1fFGRS+PT/SVTq3n8l+2AxNMpz3XCp8jIJkcn+QoxGtKjZEt2/X3hGgLCN/LMxDm
TNPqa/T7Vf4IIXCKa9UgpPzusPs+J9FnxtnD9JF44NmB2U1anPDum71u9QN5lWJglfhbKRp6xoEl
yrqa89IswtESGdZLFStuE707FaEcHo7YkLTFyDAdtcUOAmnAoNHifVlXUF4eoeeY/fhMnc8jm6Yr
ra/hlBu0DIYwKOzuYtXWfXi+gUeuje8pFPcGDNK4aqRBpP9ml44ym0MNCU1C/bOpCJOtpv39Ttfk
gmUkFvn6vIbEN4GMaF5UYGyzVVLjv07+/eMRCnH2yuKYsDS4H/qDlDx1UhxTuOW3khVqjEwjf7Dn
t5/0MRgrAqCPP70qPYzUZ9AjKsATIsMA8SZqKHDDJjhKUHvFiPM61cXT+OnOCw2cI6zEHzlz5bTy
cgBXj/EIgZ2NSUYHw5i/LXKOM92sds8q9xq6aghM9QJPigr2JDG618AGWGU6VQa3zaeLnCJb8rBQ
PIFEGHuSdxDHcukvwd1oJfPzwW6hrStR4mZ95iXBIBdDkW7A68Kp60lZG/5LvpKJJgNAh1zQEFgK
StBU1fY8WayVDpE0KsAI39oZwhEg53Q2pbdZkvjapGiQTyHzJuUrzCA73YeFrM4HcoBXLkqUL9Ms
BS2L1H23FkWnB96M4sFduUTECEwSiIvOsM5ovd43mQ+gF3QZxRlixYnRPiFImNMy9IzYesADKwiI
kjI3SgHenKf/uEjQT/OVf3lbGQdkYDtV90yYLADCrVF2UH/aP8njKlzeITlGzSSHshdBVLdaKKxu
9dILhlFxkUnKW96jdasUVZ9jJPIxfK7XydSVF078nz/aZ/m5EVdfgRxY6/rBjdM5AYmfkOylvJ8H
C0oKa1voUlTuOSy5Sgcfkpvj5CSQsNSBymml6SgK6sJvRUN2wJZPeC85AfvgikuA/h2dA3Cp/55r
0qvF5kXKpdyjl7lOscwsvQR0Md6EN2WtmGmfvaZ805pQk0SXOD/ZtJ2jjRlIVqnSMmQNSXHvkbEL
3j2bJrOy3hlbIF0Oz1sPvl8wAMyA4pW494y2u7y253VA2Z4jSyuRSzVBt9YdqzMqaWFaM8MLSmrt
l3bEdGrlB5KHiR0A/AWVYeqRfjTao8+PIjAgmOsrMzU61u5YcKSpVQ0HriaLe37bq2v1G/8oBMFG
Fc+M+GYp95EVV1H0ZAi0a+scT7ZsioYTrQO+2/nC+qyXTn/qQ2a/quUCGzaWHlhfOPvNgtCORx+8
qsGYlGOGRejdFwn9e12M28u3oItVCkhXInJKRszaq5coXs4OHig983fx2SUUuigmvcaRYwp6PzK/
lWTi8sSphVZ2LNWoC8cYl4jgykFoOAfR05bSVD9p5ly8GMThqjs59p9aEQ8UqTabqkldTyMf+ttU
dezgEY33DjTKs93KlJ4xC8n5FuolBLWcf4VHOGnw5Q8Xn+5lkXmiepRNIB9nPBToHF1s4kN189S5
ovVtOtZNVDTwTL3Zjlmo8d8by37Av54L2+JjryODaCEmRr4We+dUVz/EhZ0fHQp45edpaV/6rWD1
HaUxeY21FQbh4L+9ZsvQG2K7iXz07aqgaGAsCFqfV6x4MQ2ogfYB8fLvI1hdqYatIwQuZxLI0Q1a
qv2PQTmDlNc8SHiUQstL5uGg1njyAjXeidZySbfi0i4HlX0BfuR+PgV/2+O/mVQq3ZAwcyGp4TMp
yVadf3VIGlbS3HIKbbv+7oxJa0ks4q3KSn1EfwXuMXi98osNUwcjIv3Y7U25Ek84F+JY/ZptcUem
FEhdqfiLJjKOrb78kKwpHYtvGZo9iel0Wh8C0B/E9aotjHY6uE/VUP6Zrdsnqk/E3ZA8kr8OTCBX
wU2l4mlQHHBRmO69KQywEVnW0Ybvdp3lteG97c4eiGKIMsEI7CZqQ5g71B62ae0Krh484E+j1Gov
nkXVPdQcnpitCX5sSvI+jV8wk0y18kdRdvTjiquqzkKmicHJ9ZMsXA4y0ludmmAQ68wa3Ac5PzAA
KmrNH2sfR9c+64T/oEriJMomddloD7AK9jyc//reULtSQz1Edm2Xwyy+lXAV1H/Hpl6AuMve631U
OuidiKG7oZO/0ICCc7e8Tr8h0TRabRlL5bWlrZzLVb06biV36bwdoowdzSYxNzWcqUxdRQnwjD4r
SoSV6HCzUMLbndMpU54avFpS1ftDucR/EKuF79ocrDOWAHC5B7rQ6zK+pARCR9WkelfYzF7hpOAW
XhVCLkzyBzNpPfv4U2sov6AZwdRm9kXJPt9qC801qfoso1+YtRccwiLA67kfpAcnHCqvdOQFjr47
wkZak84ClVAqaxR0/1QkZoob3hh6ihPBoY8qaFJwkLUqvAeAiEbvnlawJXolDNrvd1xrKxV3SLkP
I8n6KoVWPO+7tEF/5UUPlWpdjzBzvfwU59Hf3NOmj6RxMiTAdvS03UnHAVHBv3TPMGyle+HsGLbu
DoNQ5QHLCNBnpQM40GtR6sEYkRxPvh8p0McSFA9BbGdCUu3Qj2WR3KPiXusPHKhyg8hofkVESWri
JZqYOaiLjyjsru6WBT9MoSia6/KqDzK4xEUjNF0QjSm9bXmEozKFxw+VUbp/UrqaBTO2h2Vsnfv1
PclRE1iOhnlkEo8onoKxVaswKxtlV+jGLmrhQIkm0I26ONCK7dnyhRgCXWtQ30ZK8LXsgkRdV4tD
C4Zbee0FEZo11fXzUOo53jMSCxTJeFX9g9C80nMaXFQH4Q4mQqL3CvmrAxao5rtwwb5JFDbGXAco
8ZqCwS/ckkLr4HsZdq0fVKYTu+RiKytXbPtMKK9M/NUB34EroPfeInKUkpwXSZ51874D13K7m5Dc
FI/Adv1Pb2ZbnaMwl/+0P7y24jlJTvAby0C3wUfaeSB6KWd0hm+2YiBINEtM10M8jEk5ipf5P0bw
EVKsbur7T0EMSiIvhdcdutInuX5bqAKBvo2ye5kGKmg98+h14dTzNXqyMwGff2+As0tyk23EHwMe
eIEZEN7cqV3c2rq5iDStA9O6ZzMqOcGhgIT8kPIrFQ+UovBT2D5eaJXfmdopt/Dh1uXR8CBHXXFQ
fu/0bQlErLHr1gCJUL31eZOW4v/sJZlyS3KDVVTthqKP3WJ9EYh2DF09t03JAmDNeoNQMQT2DzAk
DQ40sScI2EEqVeKGrAfIqkidtt/CxATzY/KCEIUct33zEczjtI/ihQ9IQ4t9mh+ZL1YuaBpVXfQj
M3qAfWDP1ZS2zlLBuaNvTtpozhPd+g/Tgt1WGvYpEQQ5d7KT1bPn+kQxm4oBf61OrQms0xECqTqL
QY7W9cXRHTTARjhSp0bqDoBazEJvgjPlyrY17JBT8kgynw0Ekub5RappXFuUj3hxHYq5wcfR2awt
tGJXLUpnIcUZ/CyQ1mvjjAfKCmKQEVm0MuRAd1BMMppFYskr4XnvuF/KYNYWW5+Fn5fiZ+92wbPN
GtScfvideSgJ2t+b63UZfWXzQ2CoLtX0cnnsmYD13YoN7khshz0oXV1vHTmRMh+cMqFA95Mch1Qx
iSghAyxPnYidY5AUsuRrrnWG0bBhkEuWS2SCIBS+tYi6zGSGhJWBa93ZLi/CuST3Xl7ErgAJaOYM
0i12nzNjUiG8Q9phDT5lJoKaCEN/0CMuFHcoeizSdziUYmRh0ybIdxd1EN0k8E5+Nvc4TZPAi0nl
pUo55fat31h8xA2wYSKVEbnVBbehR3jP/WhFd1rOmzQbuMJGcc+zf7yEKWR+v/TanffiE9lCrXYG
fN1s84UEpgIL3luz5qheJiJqXx8lrzSBJiUOxWclO9xV834Kl7Mrk/vzP2PsKiesIBKKady7lNK1
WOGk1PnxFO/gg7l4KlePK3qYpSqFvqwMLcOsoG9oeH7E4XG0RHxLKfa6tNy3LEEe4ngw5nepZ4sp
IVGEH+YCC1GLXhMOJgnrOxNSPeSqB6dYwjRbW28oPGeROMAmP6TpSRDk5qTbWmFiPqdBBRJSc77o
JMV1QZJluLMyQXcKyRx5w8X15wakTonPNv2GqlPXwBw07+ds0ulKBiOtfTNZgp52Gtj50lFlXEib
k0I6EhiJZn3lvrlGJWwD0dkUoVtGmDzijD51X318dxHe3pde6ezQZGjbmp4MHcYWZZTsQWv3tcyl
utsCoscybrB/43HFoiW7Z9CvDWSDGyLhQUoMK1m3XIKwoqKm/J64D5QZTguScq0khUsS9iXI0BIL
Lkw95+99/tHQ+kSEAoL+n4ezGYt65HKaoLnvVzlbroGDAwwUUgodwj3EWafNNN3blzVhuqveLRD3
YcAM5OT2FKJDzjX/p8eStGo1HA2BYyTMFTZ44ICIWnez3uCH7vQULvKTw8UrGE7zrLdS/znWiuh0
NDDT7H4Wm/a7qu/xLuhOHxu6iKpx8ZDeMka7Q2xm0R1K4DNtONtvbXcApx6NydkgF816qal9rQQ1
lO/Cvqgp0MRSp+Mi2qW8Xv5e8c32pNDjL56FN1IEpph+XKM7rt0T9L6n6Kb6c5s+VzHihINb5FUV
RCbZtzkGN1bTSV0nRFoTt2JwfA2T9DerHON/GEqiA5nqLfiTySJWVwnvKnNRXbFaoW/OKmvomx5e
I+vbBBbj1H6rGqtOk2qUO/l9YQJEAwtv38PJQgCJJZFlfyupirllS2QaJX9DjHjgrKioFU9or7bL
76pCpDQkdNTvcw2uAha4WWRWxhNEzbqxKKYPxRrYytZI9HggcIYGpSQbogGWGkWXeMoU1EF+pTzF
PfCWKlFQMbMYpTirFnm/2soyhax/JOrRbqkVGhkd961pRGFBwGkCHeM5h20caWKNv04AjGn/4YTk
QNTw/J7qRWDhyalv+W1Pen7VsSDFx6JjL1YadqRnISeYOP7VQLKgeU21lzraki5OErPi+xuYuDAl
0VzvRugnSQrMIMbzVQtlVpHmo9+hKbTLrrahvqo0brpGx/z/83C3Yv2BFMlN+8Htr8L/MDEa8mb0
U0KeUD7a59ftmmj4qfnVNJVxO+w2mlOUyJs9+dNE24DnGaaqn6FIgH3CsAqbHtI6YN6rvcAfIy5A
OGTTj+CvnDGTZNArzbaSK8pWH4pEhe2YFmUTKSMoa5+N5AduG27QG2vdqmGoCzknrzj8wIOX2oDa
J0CqVw7CUBIlo/EYxRzHRornUyHHfhYPuhXzISev79oyZBGmrAy6erkt478mOT6VqvH0++X+eMUZ
XbAJrM8DmOqtk4/LjAYe5WPJUn6yYo7BguVAzq9Zn/AYAZCEYi4+JVm9Zk+pfeD5OtcdVm0T7j1C
e4ch7jxoJEpnXeQI7lxT6b0TQJKN9VMgWYjmZd+BPfMPq/a4HRhFrXP6+RgS9GkModorz8HZ8aPd
hVqdzCa5tEjUL5i7xD23dw8Avh/pJbSHxatIcIgcjnqV2eUF4pw0HGg9iOLDz/dv1j3W14mVZznQ
zn2oO4gFxLs27xP+4jLib3dUhptr0x49JMwYKLrt4HMqObBp1kVimJg01PPWi3NoItlutj4YXjDu
KJRdBhmd1dYtI90jkhbBMc2mIQJ9L/NJu4T7MiSdLVq2/Armia7KhmY7OJAQbfOYJv16sd7fRj6l
Og+OGlPj2tIxi6tvRyA4TIoRi5WlXAuJeBcg0fp5/BUvsxJXujW684vPLm6QqE4ZBu33GnUJMHrh
7YmzJ+HYw9IlbWHo/XMArJVxdnbW65q9hqmZekBnwBlntamxlQO09qCMaUG6w7p5fiNhfoppmxjd
/MVDYjKEb9b5E6j1sIgHW6VlslZlpT8SmAnctWKCUxBXD2Q5e4VAo+M0N/Q6vphJHMgr2WNwkG2u
K4UO0DRxRis8eAyL2e54zEXqbfbDBjxxaqCW/JvEFXzZNL6l3ppn0z6tBp/0fWqRq8wwk0R6qSc4
ZpN4xeVgqq5OuSYA2WZ6CBYwy13j4tG2ai52pFgnd/2KjS6uKU6LUuuyYw4s9qmLOhp24Ar9XtW4
jJo8+R1T+uvKTqdUb+pENxQLieYsvYO0JEFxqRXwe9o694R8nq6FcdJ84DR+2DkxGGHYHEBd7UwF
Mt1Xxl0SomJHnfgb/69OZG8dQdnjwLXNFEm8Oc1rX5wh/jTwjeH4RTn20SizeDxBFpIU54vDO9lI
wAC/vRHpQcp7qINq3Jk4E8A5UWQ3LLeqqEhaWHx0/CBbW7LpIzym4EQ2wF5TBwaXQ8/4cXdky5jm
j0pg+ynEgzon4Tn/Swfa+XZ5OL+SJXlrFCj1ztEw9DqsRw2AngWhUhpqWacrxThYfkTdEwQQxsDT
0onxZqRzT8hhcRcehZe+/DHIA2gb1HBDbsL1TTwfPnYR8FnvLThgaqNIrY564DQhCg9h8769plA/
T9cOr0Y4h2JNodMXCuB5yzocn9NhD5dCB9vmDzPt3/oxw1f47i04CRQb4etUKFRYUobEs4RudmDL
EY5zhL5ItRaTcyqMji0R0qIKbsWWtOMiAq3qqXYmSxpeH8fAz0I7IhzQURMH1EdytS8ojdltRJ7x
Qpg6Sqoyb3+MtB0XrOnbJ/9rhfNXZN6L/ms6Ok5rKZ1fR5rY8ZiezndJ237adBOUQoymXXY0WitE
RpXTIPrcJ+FT4L667fUvKJ9NsuZ+ArhK+jNq3zbSm+oNUZfP2oj1HCfmVRWZT5FviQU/VKUZp8h4
gGCV6J0vdQLoQK/UFqAXjGhUl+skQXO3k1UanwrwXQSW9AjkKXgUUQY3yMWnyc3OEp1K6CR5YK/A
GVaSp/39zCD1Xg16Kng8XhRiZlwnRrTZg8/sroywdvKi0ezAkXNiJZai8bIS310GtCi3+rI7P+aS
s+gUAh1Q8M7AURg1R9Tg075ZovauvEGsMDV66PjnPiWrHp9LgeUwRPdi3+fWHnqePNKnWw5SrUib
zRKi6gx/wPCkQ7Ddb+dIXeRwWTxVAqOIl6EYlG7EbgK0hGJ7v/GZ/pB/W59eOUsVXpjxtPlBDV3Y
M3Le6Lu57WtVQ0nPCVyMBp8uvTnIzddvgdCYyacVGKlJ02S7WYE342r2lMGLnA4YfHkOVTudCau4
jok5lRMpPfpb+LNUmPglCEdJds/RotDSh9zgLpSxeaecJZRsaaQtY95cnfsRPzhp5ZsPbUjUvlT3
34sYL/1Xxij6LyYv2+/KT/rxLHWqlBggyIt0g658svaZdJpGsJc0+DObM7VS8kUk/1W7li+AgH7y
f94TzpTj00X4JC0rNlDRGNb+qrAHibR7/7tWvunjG2BsvY+QZcuUMHjwoAMzJQQ6ZYsEhYUM7hT1
KaCddQU3O5Q/ugraXNqWIAOVHJkYOsG1fEbFK84D9HHH8ocTz4eLLg4qnczsO+OEreDaNc5gxP35
TeUwmT6TIk5E7TITbXzovEfaQp8Z/dd0af4hkWXygcZ5/UFVl1DpC1e5MlBKBp8WgeeJh7AEwifC
5WiXxevrXPpjQETDggKuESZrTNTqZVUaNBIKY64vyYdXGjFhPM23T1CLW61+UVSyOSAkMUXKIAP+
bUtitEcQWtBwgaE0PiHN/rKcshiARlHlj8pobSoGNt9+fxUkBQzmureDNPExfsAPWrbcHpFAb1Te
ZcGXcCnwPF7xpJiztKZlqd9D7OiU21v6Pl43mk+qFrgRxRCRSy0n2cyfm5TPS4Dw+YBU7qDpPwP+
ocj3qFrjSZgLksV0nws4mmypHGEzK7dfAzYNwtAxKz6y1of66+HoMG9sAtbQsDLdh/4ok2Rh/GDH
uqF0JLmYylMyuhoe23ORxFwfQ2tUpvK0Be3tbXnwiLpJsHdweBPVCX/CACXHU2Eu3uzpOzjzbcYl
vpFngZL49UlTH5tuj6SVPVPvdhaQ+hFAgtvbOX2zrLC2KveDeTZHGN4w1Sr3zP+KBAcAZy5JZDty
YgSqgYh1Sp18sI0FTakuNLa3LGUzIUFl2jgPSj6Dg5wJeB8NjGk2piyYQTAq+qClUJ1mpOIjNEQz
kPsJ+JJlo3UneEzy+b8rVFHGNhqUXeMXR0Zrk6FdbWkvWMrmU0RmEkg4Mf26+gMtf2OhYNvcacyZ
33pjNfoNsTyPcZH+1xfhSMI+xj7Lnix3tOYrGIBi/sQ7M4pvbCxf1g7kSp77/PRMsTcK/9/hGM61
Hmt50nohJ4Hy5L8NMYTdIhfNwZID46Fxv7EzSLRcLG3PMjSUy8W97svytCuPcOU8qvzRRhW+U+DT
xtrQeMHaD7ZaKBFusaFqAxCBQoC3dOKti6fb4r7NgemcsWkYVbZnhXagErSyCsFOeW2x7Pq1qZgc
gF/pMZ8JYUlDjqRKjqjJgJ/78wc5ZGo2tOFhDQ14yLhgsL3GRT2XtVAEhRQvbi8f0Muh2pecHiuS
YO5DsiH6VV2JEvu+7Q8b80/0XxBaiyHokEoDk+rMYJQ3ITxuYIj1GGGz9RjbQu7W3A7C5jmBpO7d
/sDHVaBesd8jMDN+iZv6c960lRT9sevyiP4lQAAa2YQ5qpSdvu6+6h9YUflYAU3bulaVdrEhTszq
OMQA552mLo6hyM1uE31kQUAKm+dI+oE1BYuFBhIiEQy17QvqvqNletyvbNzGQXy4qJxrL2W9yrmg
CRCDi1IEVf6VmmmxhPHmiRSqxQeN5FuN6IxnaqDkoKMUmB2Ti2ibJGYdK1G5SSPsXyPG7mPdr6Xj
b2zTtNDAVYQqJ1HnYT2AiY2Pt213PeNgkCFG5A0+C5g/ICbaEnXR5zxVpHUGsrl3+Ce0sHInvpgi
OKXVRsk/5N8FTqkYpAJeiOByTz5Be58/w3VvjfoBitV8PyhUGe3tK9ne9/lGMT93nXt1OhwUUcMG
0Axcz1EjWq7lO1ZuCIuHIzIpuAdOW+ytG6tXukPoR6QAi133wZRBeN2U0bQp2ucH/4/OUf18rgR+
l2YkdJziXLcjYxz48tKb5X/7uAIgzOcHJmSR+FAf8EtuGxiJuwJkbUzMKmg/nm/KBoPgx4uv3X84
jO0yETCiC4VsGWQROkE9aT4XegYwfc4LdoX6dtverYzgJa6RDwJqyAdp1DShf1cFYJ42wiBopXgI
XkU4a06v9ktYGFfnhUGOVFfusMUB8eYap94Sl9i9IxBGquo+VjGKPkJM2hfKC4dwo87ryHvu9XdG
Kx6LG/AnjrVE5plwzhjR/3TYjOgqWqx9cWRL7ZYItRz5l+IeqGSfvXxAplpkliuuAdwT7DkvjsMN
n7qgzhHBdWtkUG/utLU72kODqzGCENXXrdg6aYBcbTqW0DoiK2tLLFRfXb22ikUJ1cgJeNsZy7/o
BzrZ3WNcMxUjU75hlP7bjtKImtpDsiMPl8EaZJp2PCh4bY6oD8ghS/vY85dvFwNtso795ADGnK9v
mp9sGwDxyMeox7FCkxHDwQubyPxX2VEIZshsUCYGysYTBcqgzMmDGVdIwhsRUsJ63Qaft1988Ppi
NAqa9oYeXvuJsVOAZ4S0a9ZAqWLDlbFa5sUgB7GD/bpPC2EVbDwtNdYGvHairTHerICuhxBzBZKx
C91O2JlITU8VqYziyvJCAQuojSh6JiqRY+WUYtK8jIQ1DVsVYhnwBqJT+0wV4IsakNk3j4jK1m4i
QwlOAQifFWzZAtcR9RKqxdv2q+EfFBrzIycJsQdp8rgoizZ7HEPyAWeG8hBlXftNv+Vo0NDuYqA/
4nRgdUWJahXq6IJp0Gt8CERAaLrhRN5dOi+IQmjqzYDBaYHlQCniQc1FT9IZw48gFcmJhE9rehD0
KVLqgQLrlz0uOY+bCa5F7QVSThrXowyL5rPQ3jucshyZXkqKeRVwjl7drHqKh48RrDiEcl/1RSwP
17JyOEskMieI/aI0oWMcULcvLDb0D+/h/EbEr9a2Dk2bCv1QWHCky9EZT2iZahxT0t+S1+b4FqoN
s20QgnLKEu4BlT7f4PxN4kKro3ahaROJJg3uChpaHF/Fiaji+nJ06ObkcLcftl0cnVbAc/810fgU
BT5AZa6D/SOba+M/s/H3FgZ1Z9hBceCct/Rmvm9wNKTopUJ0LScXEj0HU5HGGMolFHRkQ5q9xAqL
y/ZNWYf21R2z6Yk4Q6jc3nnSMT+AO61Th9kuK8ajq7/G4/lHA+3OB3l3ljn48JXaoml+sjQtq4sP
DWINpw8uMXOgI619n+ttAG4F2Sy75USKE07Wrqk1oNJ26GMeD3BkZWPPUHy7fD5lXoNO0kCSenDg
cEaBWcuX5w9C8C6wJFypOsVwoSoJYpHB3kOfRVzWN8rBRah9l0wDWe0WE4GMYHXcsngwTxRHcddP
W3COpG/TJ2D+SEhPDCV73kPNi0HlePerAkb+LLOkLRXBQX4ATecjFPo5VkKRfB3NVyMrj8/J7w4q
ze/cXieDletFamoiStme87bdo/CpbeF0pJfjxjpkJerdBidPyzMSmFWCc8JJGaA4l1ud2i0cKqXT
r6cQgtr+874Z4dtXLAmIrq3TCTqkGDWIlTFBuyLqyxBD6fFQprdFYJdRooThzR+mf9mkxGpf3rIh
WJ+Z8VhAa6QTs7mg4B29lp8ytuCfBklvWTfTXk2rt+AnmK7J/7Ic9gkeMJ9LCYdfY6EHdIlHCg0T
gzTTB4vaKwfTVBkef2HOplSdbjlTkosmUQ6YCS0Js1gz2bwuZyiWrdjJ1b+Ghjxwx95XhyFogAbl
jGv7v7aqipbu4/mU1quYxqxv80Er1zQXrjMUAt8gqF+5+BWHzrzGoPI46aoPJa3QQ4xeU7G1K1fe
/L0jhcF49NO2DGvQR1i+lGZ7f/0h/zhvnIbN1V+MeBJCRAq7r+pyRjq280ZNY1cxxZholSTMXbKw
7TPziu0rQiKJrlhX4ooHcJB9Fzf3wzV3JWMKId6Gf7yz3EdNgTRzCEAYJe6zKNmB9fWfwwOQorCQ
T1VQPW6x+OCUIe3DtmQZf2oG7+NOHrShTalr6UhFwn9Ya3H+sD/zqKWdKsHM9v4c13i/HCtU93v+
kwFxbN6LZtYENK5yRA5PujtFagGcyoP6KSQ8JoSPqvLf4mueaGfTnQJgHrmyQgFZoDdocRQchh9Q
uh9BNO8aD2+1g9SWX9b2Ys3B3x/q7tYkwqi3C+9P9tCyr/WEUSgoWptIhKr43LUim1fICqC5xMe4
gGKHXcXLM9Rmag9DGsOhigHV5JKo2VYO40JpzEc4w6z59mGTYmoPp5E0aFVo2IFhIleRj7T8flWY
Fu465aU4MekFRIzuLnV0apXfUSBvqrsXnHJEuph2RJrYRNYTo6FXAAapSYjZZS1W5is2docyUqMD
F04ZZTmnLHBttMc2Sm43zTRnMCogKaacQd8bbSdnDq8L+7j4pUeDHFOwfsiX4+uc/sMOVw2Wt9iD
249ty2P97K5Cv/mzC7Wt27Zi9puVeXhgvuQib7phYd6qVZoYAtE3mu8a+ncUu+a5tQT4yFQ4FbUP
tzw6O1jE7PmqP/o3p5xyU84iGBHjmFYG73m/dCYJ4U9K4AG+jjGjgyRHvPXcQNinghAe6EbxyJLY
ahRdYCaJpxiQ/reueEUNyBscrK98tF91P/vg9AZOFdDEzfjUoQ5c0I2G5FRR2d2+tGmdMPo9Z8bj
f8pRG32bdSy/k1zsB8V8ivk8PXR5SzABEfSk19BiaRlA+iKRyOZYk+db1d7XdOTwqR3dJO/Q9cpD
gXrbtg1Qn566MDvnOIpOerQ2dSdVsbB5kzqHUsN6hPmQHa8oGVKByt3wP/iopQ+p83MyFK8Wa9RJ
u1K66/ZTKW2IDlhdMxByop6JkCv5KL2+EGQi2o7CaqXODLz56zpF7euEjrR6vrPo5tCxovoeObJz
e8GrvfXmUwDT1r2kHUQIXLX78LYVmsoP1krnZ6rfv/SdMYCvQIyhIsR2fsRjjK3ilh/szGn7dWDs
TYk4dwGvTZe3z/ryv9IuqegxXbnGTQPf8YpmyDQxwvF0hBGOaN/BkVJMkenJMIJyUostzAhgCLrt
ivcn/mNCuQmjwR5iag8/z8MtwuPBfwafw3hQG+HzzeUZb5oSsyBDatw8uIJZyLDC7D7+fsPlzthY
GYBzRmh0EX01vwglw3LQC1slinbMAa4XgLnkobwl5bdnF3nbszQFiF8T7ZPmjAH5/grrIpU1sJlv
/EOWN+HeScBDALRZbk+ujY34hhvAJQnnETPQ5Z0S/tl154YF1FUQnz5LIXrBwIb7yKX19ebm+xpa
qQc97KeE4q4psXExXHsumzni+lVRgROkGNY/vFT07vHbnUVrnsiErbGlRh+pMWeE12OKj41Rmjk7
hjIE9IzEpplPYI5YEduvGXcyRb+EkL0WQy4txF/xYteaq/3YyAJhBqHcbdK5YYOC9OaUUNs6nm8b
PGzBee30cTtHRuT5UnRRasL7qjnLkOE79QIDDCXsFMFudEgjQ3sIPpD2Jx6mxGCYXXHwJaNzSIQg
MImU2f9VqPIq+yl8+Q9/mo2bx2K+Xc11WnxXc8Ip0k58aOs1g5Chou1C/Ju1S9pQ+Qn0uva3PxZw
Z9rAj97ZTB64ETv/99yR2Dti+7TBvtATZN9MPU5BCzK3wbZJdKI4OPfGPGNkiitOr6M4RMFpFA3x
lZHOoev3iLgLu1BlNIsY9wtpH2rlOqPRNPvlWAnz/UxwqIrI6jhWBCNvakIVkqsFvURST1Xk5A83
p1+eImmAN+QcdBCRMPFaVpWmHOqVNoIIaUqM+MoElyGbAXhOZ7YgibmujaFTk1ZY/WrInMejjh5l
t3vSgxW13VSHBBgA0QhRg0iM6eSnADE0mtCuRfYFqs6RQ+YlxpgNu70G1tXSbV2IlkhD3CkUiQkW
0JBODxTxhlzqFGqVODiGWjQeYynkBZJ+DcvMdIJGpOvSR+AzeVbCS+Lp7WOWbcFlXjj/Bvj6uKUi
B3hVW8Pq3UXispdKZL6TEPyP2VMBkTctg2M6uUbiThCVFvAJ9DXGXqHBgNsV/450tks2FcbaQSsl
IMwtRP7ZjlWPnoGUHkQ2TaBta3AEdgCEby91CjBER1jEd8ywD38uAO3gpm8wbRKRytIRkyNtNqze
Dxuls9gSLFgmdQR8lVuZYlxP9ezcQrbIT4/g8XAZUieigK2IvCvlQrbAqoyf3orSnatHM7fY56dm
N4MbfJpFUFWMOobWbAcY68IlX+Ua6zKDMdoKE+A1oxMMgCLhgH4GT99XgFcgqwwO/4VqEe+REpct
uYVH7ECjmQPFZsoK2EHH4tLxcBB8kfPXzKZh02qRg4ksa6nH6K63ULrOavcJ7I7lqNNT2JxMlv18
SD8HoufHegXuedb2zXfsiS2vpf3L/odiVFZhBuxTAzsrmR0VyeMeuSwId2FDlV3JltQEFi3ealOJ
7RIC3cwq7+tb2V7wjT9/Zhcg/ltE05LE1xLA4sHLUtiP8nU4I3FXxHcs6V9qjhnYPa65bqU++iWy
2v8QQ6L2Qr7YBPBD/HwETblEDxMDkeGTnzviqDwvi8nHlGwuRxaO3FW2IkbLV2aleAaGWojviHPm
8E/4Fvn4TxNY1TwsKXEBLFeMyoXZuoIL2vMbFFWTG/P41Gs4KSKZr+MNNLe5vztGL+I2TNjwWnJs
m8/V6aIWuS7m4ybQma1Hs5WfoRe4de3fZVVl3XxRld6om+88I6dkzETgcN5u4n3qQ/NzXkmq1GeX
vb/2hvZFGFOoHgItIczRyCBWeViQg3YQkzDN8D9+bsyuyAA9UGuNCDuRbWz+r8vaoaVVsl8BV+5S
HiO9tJc1R9Up13kzCe8/Efx1n7XBkndlMZ3QVyCktToQZO5LRx427L3/XcV/ARceS35JPQmLC33r
NhaDtbxK1WmOz1iVhyoJSsBv9jck3MPHS2rAJUtEsBM5cU6mmbtDPnM8iMgbt//O0o+dUFXtt3y3
BbSjsfOkAnUT8wh45wf5USvIguoG15ER5sq0I4ZsfR4YzOaWioxmSVtA8AEtSitgENAZZNRoG/Xx
dasoz04Mz248dHFZjTS7eyzapAyDpPrzaT2f0taKUaxpIpibi/gQGJIt6t2C6O1VLQ1vv8jRGn5K
1uvN5UYzW6UYVmZxAASqdcPhCFrWbC9mOHjCsOAAZ+xxsm0xaKwjts9vMixWlp/kJsyAmRhtoV6j
+Sd/XcU3yx4xBYyIa64gzmfUPC25ww0+IHcloUhTq04FvGlqJS+jasoTxsHMKsVue+RTC1kWb7yb
2f/2L04XakdTta5O9LWFRGQvpdg4fBcmEqif3RYhXmHXtWXTBCdENSks3tRy2spGJEQ1NyodSC52
LBvoZHsUk7qnd7POyMOSZYO7hmfxWoYyGK//ZBjv1ReFBSPYuQVsisPDiikupj6qXl3VoC0Fa2Ny
ISRvb4IlC9TSZNwLH3ENt85IGdEsE2L0cBQxoBVHqzLH63aTRn+u1bdyoMrTmEzmIZbU+HEhXjNA
oSoPUMcH0tmL+oQ/s1KypQ/3RkPwHYGaN3TAYi7H6OSDGzz0kB8QK98yB70qY6o/4FvF/Y2iltOM
aJidrZc74OQYrFiQgsJc3EG4B+aTTcBstA92fOpHfnR82jz26234xZhCbjPehuoccn1asD4Hr76Q
bVka7th3ymmeiXY3fCAA6RolB1Uh0DJaq52qSeqkAaXnNs4vr83zYH+tYT3QCRJbnEv2mP0vvGyt
IpVtQZupA7q7KiPtlmoWRZ/XNLnxC5H9uHeJ9M4GBcd02dXk8d0v+7KRmQlgldjbOm9mFumYsCEM
FOq7BTvDNAP4KU80xH/737znT+GAWYC+qj0n/H2dBjnUTeNHb6MizYVwB2MlqZzf7HDxG7fvsUBy
IPDrVSQwUojjncNgvAy/D0K4mIBcwf8NOdryTraUGBBbC8rdj8eALXHcNp3D88GZo/oiEX1yN3uZ
AuYibqRnrWBM8KZEW5idmVFDgRPVobHmEaDuowRzhA70InCfeeQNrFZNt9NLbGWDSYYk9N8vcAQw
frIl6ls/tnbDWgD3e3DNePB2WCYJF6DjJJfRIh1i6+K8syvFzHPYMUFkgShGVSKF6da6Ams1UpLV
RHyOoOCwzdcGL2Zu2U6RJk2kmD/u6kSJ+mNhyTEMwndFi3VWZn4cQ/unjiBax/7BBNCIG3ZaAf3+
7Kf6JiXgywvjOoLv12sbFqZwICVRJaxbBp9OEK53oC5lhOGO/YHumDo4xqoZIFj7VvFGWqbQOc/l
iwyQak5l9Qg8uq23OVxc11FwSxUe7/w19X0q05bXLIhYS5skr8HqnsrzMGKCxVsLRFNwTn1Hsc0c
0wWUlzV4KLgspDnNz0U4FiNGittboB3pX6FxuZb5hZTsrxWHbeJxixL8do4rWgOQghykxvBEf61W
o5B50mMvWZwQ8/JWi/FWFgjOKI6Lh0+czZ63HD+xErNu0GE7xaayjaqMG5x2d2mBEWnSwTr2ZdV8
pSd3IZJcU+eFBljyfdYnLy1OXcU7wEVoIYoqwPIaslUQHG+MyCJJAf8lk5vC9R6QwfYEnEybVLtd
tW+xRQSMTH9R4QUYc4h2y19cG2EEnPtMpPhtkJJ0RicuB2saOdAe7wGtmXN4BqkMq0yulA9BqR0R
syFXJPIr38Z/unyJEJRSqTQHAstEtE4w1gE6AAkOQt0rd4HIHNSYBhed9hVsF4D3vWzDhJibswam
lpAfS5d7M+r/ULzZqZ8aAIlf8oPBSDd1OxaME5uiRakyO7VANQ6hFbJXjDBZDsgL4lenMTzK/DHY
9S0fbigGplYcmtBF3KBuAoSFagKoOyPSHDbg8V4dP8c2oj4aG+DTauFaKpVoxuft0glB+rI/iToa
dGD2m1qmAgCv3Q03Eh2vVcY7OYQP8gfQtMKgZxwfOI91PrMKQP3e3KWZLoin2GOi2YhMRLqI4H17
uk6ICj/5rb1qpZVe+bbmu3DchzuZCtuXqvTWZW5w+/gDMlLERCSrGICgprdp7PRohAIdYyYG6SzD
QodDhxikZ4uxKBu8B5HJPr/PgRSkU6sKxJOasnl1s1il+0WgLBCUWHb+lEgTdwBNKgPtEtPVcNtT
OzxGeEhdu5p/hCfffZ5G5ggh8clSvsyUauvCy0kWArCYDgvNqo7INeic9ukKbMi7yDgen73AnKh6
YOxTA7JdboPtkFSWqtHRlxIyBgtkFbW7cyqbbSg1dDR530Qa2T8KVt/EWsVBli/t1P80XS6VPG2x
QT/kVXbgr8Lb3b0h81JquDNiwNkPsaYxa6OX120ts1L9W7Tg3WVWALhc42AbSAbqB3fTHQf/I3KT
X8Qwd/ibkzKz4D7BVuNFfaXxu0jJBEAt12vQRmezdgUpvyi1b9KOp2cMl9WsrmsGGgNvbfJvvzcT
GIDLurrd0akdsvFBFiLYJnv9GSE5UNaDiX8pmoqOyiSy34Gglr+748NC2ftKDEKeUg+FsOIDB2JI
4Au0wKGC7nfQdJOhbMtabiNY6Fk5S10XO+EaWyrqYbOs5g6nWthBbNNntXIFRaazUooNb3iP4NuH
JM08yXZSK6/zIhp6sReln//qrJsQb4p9YbIFBd3Mk1aZGYcb1jH+n2bclEWfj07r9Mr+1B/a+bYv
h1glT97y4fjrxEqIqUJlYklfAwgrGJhc/sIHJKZBWmlCEUpnNImBfcdTuhLxg6GQQK1pIncBYEz9
Qoa+ssjwJmcuEbDXcXsGzwc8ZJW6zx+DyXvgoQToWKvKY+XzheH8YU2CxbT0BK4t7TT3i1v9+GgO
up4qDFHcclUvT9CnMM9WeW6qdPTFtzc3YHKlpI9wTm9bCU+xLlaiV3SkRktDF5g7Sep+UODnASmS
YkQZSz/Enq4W1LThSaMWXIc6B2dTfmlvUDyodUTztm3quLQxxIjVJTHcwrgTWNgSKh4wTCuHthoI
s4TX39sVQY9b+lT37tBEYi5kdcXfIgZHnCYWT5Dn368AEJ5po5VtDFtTC8yHP9eR206RiuWEwHHZ
Vvx5AjyQcrDWOtW/DcgX0R00OQ6djQNFTCc7kaxBS+3yCsQ2m1RXWwbs90AqiR032eRrWQmy/EJj
CFk77+bYpXvM0yQMc8t0KCnnAxbyrn8z18rehoQ3nvQ+4XI9R9IbbUk3QpTb4SvEf4hoRAG9QV0x
2M6Ef15uz34dB3E8f+O4f55K6cKsbQ812r6UouHVBIAsJc/wxTFMmcU3ghQxs/E0GZJRULGurd37
/twAVcPsgpsupzLEBa2MUV7Cz9OoCtLOD5+u1NLumgDCDCY4eg6uVRmP4VZ3XXD+vF8zpuhAM/Zn
zJT3IOslnmb/3i3xN5tOfUSaS1BCiKgacF1TWaUzNFV54rFx9v+0ofKcLe1MGm7rYe8OUN43sFfo
U8jT9s1d0rN+WrM6ciucQEcfqXH8CrTAUTrrcLzuSZ0pi0ONM9bV7F8J3XumoHXL6ywg6nEymPgX
Z0/6sIxYNa3hG+q81IyI38xYJK35TAN8yRUwFDPkiElN2Djd73q9au+Js50/hIHU3hcrkQ2uH+tI
sqqg+ErXFBEnIdept27ZRONSuHedyoLfNRuMuFD670foDyQck4G4wq050VuhDUrE2j0kGQ3QESQa
OzgJQWVXir3KmGpmvuDkHOsw0Y5mAE5laBy+AkC4OG2Cz/JQfCf6U9X7OB20/+tzmU8BHORB1Xi5
u5+RGFp07f9CeEVGjIvbQ523VRGJeenjU9RzkmvJQZ5026rIyIpY1pWtK76APm0e6jX4tZRcSO+I
n5I3TO4MfP3K/FPeDtPThmCMgO+w3HL7tjVyJv1lXwOiDCbtohNkKCErxpXVHVoYrvn+lEDh3LuA
QSTYRmp7G33qayBDUU1PgdEH0weUztjLXBklGlbSWERn6DZfP4HERkg9ygmIQlVe2NCNKW2WQjbE
LbPE3R1JrnuXmVAMvcKI1puMeql9gdqgWCwgEdocBkAUov68LxlYrVCwJ3pda2DUAOgylQo7zcGE
j4xtniYh16XmDkulOL2VLfMtiSs6YgjA/eF+z81FWJuiKVooxBshBIDT5KixqE2QpILBdCsYOoBb
o2h703Gruwl613VCMazgIyLHYj2sqzicWjiMwbb8vxOx87BitsZfnUlJ3pbmAmNsfd/dfoRdE2bo
7FbQGE+CHa6PBLa0KPBzcvh9RShjeYkpsWyg9uu99o9NuQmGdqAdem22lyWuzyhjyEcVVr/4+H4L
1GWvnNQKKPVbTJqHn5wX8qMj74TvomPxnr0tqfxm/1X7UrnrlIHaTUfMIOxeMVVyK/ilAGtdS4H1
JFq5lCQcM0CVkAm5fU3mNaFLZstktXT+R7HzThNn9r5saQmBuF1eHwHSCT2vEDxSoXJIs4UW+8ea
xGoonVLM3hiwf5MmFWhJ5ksh2r21ZfkBbprN3aGG85yr3VKmSZ9Co3i6PPvNZf/8nFe1PEimiY5n
0W5fIAIQsWZQBv0yP7EwF9fKgX0fK5g/CJPu8JmP+ITMMPzwQ+dQ1spC1Mg2JO5/Ke9FeHSzOqMz
OiN3ynjWqiNeZdzNBb7sCzmZi/6KVyJOMluk46sg3OBrSydVOWEXZUS0Jbl00VmlsK31lQ/AdfkX
Zudm9ZwIDYTPd7e3e3I1r/KtO2xQ8WiMM69wGQ9z2xh/fwcCn+8F3SoWjB0rTc3BUYtF9Yi2HxMV
u8/gRrg3LLfp71dhTtWWx+zD9bMYEe4jm5uKPd8LTbwTcXrGvT/wMns+7phc4MJ0NZZ9wU9wXq/g
PzivkVPw3pftcRMvj4ITIUsfOLvB3OKklQ+yDMtIwbH3NjxxUCd3r0DFqMLc4pvK/MmigLiZfkox
TL4CE2r8h7i9hLkSLklvcTexu4Xm1qbkHvPve+RTC+1oCSkYo1mSlplmnTDYpqmif5HwbN3boS4X
sTjNwMU3+ectzfpQ8d0TxFpeZopMoY4Iln3ekG5V2AVxWylmb31+59c60dtGXQPeJqeI49N/f0Rn
SAPXfUiA9mmtpYI0jv5pW3uRAT/HaagJBsqIZnbI31Yxw29h1UiG1zAbmYi9MoL70Z1sqKhYC/vJ
UOk54HTJZxTUnJISsiZlymcnSyG/Oo1EyL/C4GToKUHaDQUdu43+ojwiKbn134t6JIdZtD3ZemKn
A+Cx8Drf3Ol33DvZMEIWbB7BtDCSH7hrSJplDdBdTg3cj6QFf2JG1YuwpRsnv25m6/XQ4X8OEhW5
HDiH9LBPLqlJHkUzfTMwjyVHZ66wqKwCoIYBvcyfeCoQiNCcz5hDv2Rli6vPxcxj+4QiHGoSGRWP
fl4/adhidT3hjXtB+SGR919LugSCpMTzdHW+BP+Xo/FiwG0VGJLetpNmKtdk8AK6oQaOxOiiDRm7
Uhq7bscNWxiiJrG++reO7mskwzMV3/lwKDth7VrOxkO8MlGqI4DmNsqcgZtlmnB0aYHAiER0yh/B
NCtpIsKQPa5buGIp9MU0LtESy2IhhtG3CLFEMSoVc/jnLYfI5SeBNSrV4CT3fm2E8F1obAgyR31e
/3i5Fxv/HsrqGp+VAJTy04KVcCJSlNQGy1ubGxDvy+AJ50UA3clTU+v6AQzFrKLzOUpWNzw5asgt
WR7HsnCHZK8sR1aVcjsMknwm8r6z4VJmP02lMYqPXwxbVB6+5PxnPNPntt4OHmnu+Pl5ZfQ9fwQ1
6H3AXh7F7AWLUfP/qgmAoxJ4hTsTgQfazDy5cgLIxi3vXKXszNrhuugIM5UDehxqXFHqu2OhxkHb
rKxqGnC94i9ed1mAepMO2SST1MF6DBk7BDy2pzdao1HH5Vbfrok8/WZJTsU1azl4jvGlICD2CHI+
8ZoFF+/r2nH17UrSBySJ04VU77vPsTBBB60nL2KpOHcG7HzL/FUoAdlL5Rh7MfcROPCSRBiqfpvc
txuCcb2unEz15BnxPtvNzWpJLhsRylWxr6F0E9VyHICn9iWEQe+H4Mc0XIXonr0ZMhFOpzXWwC+0
Gey62tuwMXqEz+Z4YDQ7E5Z0BvYvT94rauHH07hd7TZq41jKufJvdYYFtq6TsYvdTsPlzHtin2xw
oMIX958ejPo2+fVhkKNMHkHd1c9dgWRxLYMhir4UnHyBiTuIToYc1m0LZEXwn7h9xfSloyS9DUoT
0f/8qBcHqIHFeCSCMuO0jxZwgJcyVwhWlh1/eSq3ld7VzZkvEpDuWnSjBE9hZM3kHNESog9Fr7o1
q7q9uUJzmlvsNAzpHu5uu+XPK8e+aqD2hNdzYUB3b2HjdZr9VRwaWvm9ZIsWzJ9NP0M45OHC4vfQ
bvdMr5Qw6zOlgUopq+YqTM5bAyfoz11Q16DfxT2LtzNG5gD/ylzS7UDPE9lWxfmFIDD2xts+xKRj
U0pbQZwrEW5tpslFxSMKRaATjcgbz0RpTIswgxsEoawkyo77bcfSZKnxxGPWRsf/QHEMs7zFFXC1
SAqAes6MgZfns2db5Ff9m469zxu2XKL0kpwbaXajwX1kyYh4csuebBLJPNDsNWTubhxczWUrZldh
GCouaJh+87G9U078pfV1PwO6D3h3fBzoe2/8o8xr0hpC5SDG3XxiW/R4SwN4YVNwh+XLoeO4/tJZ
xzE44ITugUcE6u1OUwiL9dSSWJPtxjynmbPz6zhlysOSfiigCpJuK+K9k1j7eM3mlVUluS2Rdagl
iXgRR0rR0rCP18uEDCKQ+iGQGXgISuO6E+7/rMJCkbblj/jzeAfg1La5qbwj6epAOMSQ65q5csZ/
E1BsCS3JMOYfV20wW5PMblmZTNJp6hzOKhlDcglpd7FQSBguiXVwUjpZF9znK4uU+1a0nSX/MM+P
4TwiOMh+tG9AOz2JzB2pJtXZd6qbWTbijkCID1NWNCcERQ8I1McPkZCpyv1aesI8tbzs2Tt9dvjJ
CrPWDZABeGsxlWViUdtponytgfWaou20ZbSBBTFzD/EeF/Y8O9v7g8eGc0ghyeJQemXaNz6baI6i
qJ6T9uGEh4/L7jrDDNuuZs+KkS2HzeIVek0K+9Ux5Amx9lcqO7aTGHW3q5smw8VfH39rmMit+UmM
nKLJF4taXc1x/He1034yK6eph62ZeIzb9qsL2nPtuhqvflcTRuDH8NWESUaNlIQkLbvhsyD06ExZ
Lw0lzWejCdzE0yAstXJaLzTcHydVoRNXBTLgPvFH+2Rs8jiiYu98N4DdFIY/juiMcx6NaufADA1a
bAlydaDYSErpMxJNw26Np7Q5WiTTpOixXmpaV3XAqGYIcPcTxgt/uvBf6vyVif9Ve6DCmYBgqPW6
IEGBwJY/dR52yiHUDwGbZwG84/7c3S/ubNEtrnQ+P3JiqCMkOee40vclf/WiU4+CJ26b/vGCX910
zf4oIlvp+63s5qoI3nbR8nWm8MxkOk5fH1Ee7E3TB5jx64GAWq98kR9vM6dvw2he+K+RlPRtSLvd
Dhgb9ziNxHvP0SQwchzIVlwi1lEHix11q5PiXaCBsxWNPNWUNpd22ltPHsVDVlzQCKG4WCUArXE5
tEJFIoko8Hbct22Taq0kuhIi4Svb3rowD+9iOejGfrJX9MeFu3b9pmJ6cNlWdpWSxXd6HQCFw8Az
fkFWOH/jQ1lyvzjCC1L8qaX+ol0WkljJ0S2BIyqk8llVJLvUWVcZY69ud6rSnQJWy33YmDLFDt8H
niGRQwXSdx/saCESVaR0r1iQ9KiqKzpK67lYvT+MhyBvmM6wKmTHb4IVZLp74X8CfmOvWFpsXKn5
HANIsBol1lAquQku9sZKvY0/Dailf/YSy/cV+P4i5k+je3mWJ5KmMI3vqtteKd0exgU4pH89ZDuW
eqNCE8lu3zqB0i2I2RqgISTo8l9EgHJEefGoE1FbqiyVPvIBOSDQOVutNJXYd/LdbyhIHeN4S1Ye
G+JROTbwT+iIFd3AnlvQzUgq2Vo20MvNXgJHUlcIWEsgZbx6ylY1fgLLlmi6aB7sHRHeZgkg2ehr
Zb5VCn94R4TCcuRqSct648h6StoE38epkDweWpV38QRRXxkhsr6mUqiWfF86eWTsOdXbfrCuQtwk
c1/kNgT5yNokGBOyJ1UKaZeTtTXaqU6LG6JrFnz2TGJ71ukLkWi7HG1TbJqvtcjwKqS3epVrU33j
ZbD39Sz7HKQe6qDOwet0E7PRmma7pXqYjbokBLhhPw95TW0riWvU6E9+9YCh8ayp78agUvH258+y
7IMzQ8Ik7qZkA2qp1qHIvcwOV0w1uIL+amlTXiD171SORKw2wMMevf5FHKDWJ8y4JFRKQwletP9u
N61nA4EwUxnpJexuHv2DVcr1dk37vmnVrzG/zPizbib6VYqUbBwX/SkCxZFQuIHv9X48nPta8t0a
GM0K6p8FxIO7a2obJZsm4I2CXT9Hf7N4J8Br714Dj02u65Gu1amY8loplATa3n+IsFGBzOlJhOCW
AKs27j8KytJrX9jna9WVyIaXqTnb9hp2pxROH5ZwXySGPfnKNZuOiHEEjrKY9Zct5qtzK6driY8a
EtS0QvENROXaIK5aP5Pdx94/r7D52Z4C3zkw56k6iO2He4yq2XSAYKlMVZfiJF1zgCcHiWl4svHb
T/PTKZetBA==
`protect end_protected
