--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
WVZKltK6sISmm5i5f5726btzxg2Un0rkhuUuHuP7pws+QeV3TKHcu2fsJMB5y0FExYR+VZyEIajG
v/XOomtF+s2EZNJzu6lOzFpQ8u0uABejCApy/YjQC5o8HMg2G2IIYrAe87XtiAEobnRpUnMP6dZq
Sm+4cqyG6jxE6dlL+W0BZ5YV/OO0bB39F2roCvYfv4R6zjJPzFx3CsWL0zxz1CJch7aJ3+oL+7Zy
xLwpHzN/BYzPAmKFxasLgN/IJ5rZuqiIv7coNJL/6aBRBDzW5k4n3QtIAlawm/1NgVFTqfdYiZ8k
jRi47qqUYdpX0GwFQ90dtX/89dBI+AwJcClO2A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Kbi05RtnnjO2X6/UcTjR6/p8YFGn+Yw/TAPVSDDxNEU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
gtV5oNTDFzUQqGRJBeoWEdYy7H3hutBEQ1f8d80Q8Jdc0Y3SFMYNYmoY4lqcSgeb8rULNwmnJjNP
CI5N+YOgcL/0UMFbCkNeOEIl3/tLrEw9eQ4phaBwkCRzON/u9yaXT317a/EHbkIxmMZoYDQgE0jB
1zVI9Jmuv42JqaMhm26EFC9SpWZYLAYubRRR7thjrfPOJXIw+Uv6AD+Qn7uBD5d7B9ef6VVhD8rq
glZGWE7msft43gUyO1rEw5c8MvndGZdCGr6cKYfKPJr3S16y+E+sP0kJkZVhiEAokBuGHDPlk/Wc
MYHvUoHALAQnhMzGcuFZWTmMp+HKpNM4vXUovQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="k8XvqRpUJrgfrkufg/sZlk4KzUnm+izhWyTE/vD5bXY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2464)
`protect data_block
HBO4+doiyL0r9rNI7QDJm7LK33js9RqCJQTkT+I5as7L8R4opVK8kpxYmJiOOGyKl1KwLyVlNp4x
X7pN+FiSxWQiE4YN6FkAHK/uZe7iQ5sDpBwlBOpw2uGlvcBWQNV8nxDilXrJMcgsQBDIYaA3RP4+
bT1z+VYxrRzQg2RK9U6pWj3gxjUYerM3Wmes/mCOkPplZ79yZHNa2ACEZnfIJ9135bO73DeIT1xn
hLV+AL/8FdARq7FPFRcxfEbtaU5vk2ZPUt3beC1woh2B545ErpvtGCoRrSJjXz1mEghMCfKn4gPU
bZ7A+9Q+POdQCWkKHhzuzLoVJHqvNlH1ET+aEEJg3Qqdn/CoQxEu5JMV2O1Zt9BGM73mOwtHnJjp
rcZ0edppXE5cKXs6+9zT+d5NHUKNKZGYQXTx7E2fGNATeXOar2lPLFnvatAczmLJZwmIHQypWz8X
toCcsjGRsqpA7T9SsV2nOL/LohQkI9e0TVxUMAGmgLHisqq8PzexXo+BiHTn4g/1QYXDY4iFC+M7
RJqIYAONg2KSiBnqSPrb/JDYKMgUT5FTO6pbqaoqLrRr5yRBhy56MjsMz12x3Ct1AQcErwwrc8CH
JX/t3b9phCb8JpQ56ieWeL3hL3xRgOal1qGPN+wUWYb2c4gpIq3zaVa5qOaAzihvwNaDQ9KkMKJP
UzV1ndRTjGYwaQKV4/CGxhCIMFpUjEd9HctOhZfk5+wbMpXW4ox2bwBfVkPsRZhMrXTbSvlTI5rr
DM3b9XCV5vByXdH+0m4JnlUoPHYcoU2Dr/eZ67wyCUqpI5iv3033RBZGiqw+88H1p99eMOdQr3Oi
jYw+k7p2qAD899kTDwFhmmZJDMwYqMLzNBMFOC52Dnx2pMqVxynLJ9+aGInS6G78ES/7jLZ6+8J7
0F5x5nm1JpTrSmK7azvxsXT753pd+dGcbHtLzswKvOeBi1Cz38DonB86ThlWPKSEamKFDBfJpuN5
x61KbWfrQrABF6L1qruwi0aC8Of1x3ViIwJ4V0Th3x0qy68Z+0jMHqz2h0PQ9aBF3iAsI6kdFvm5
yyDxsBaHqVIwYZxUj1TCxsQI05HB6Ep7FZ0MMiP0Q2CvceCch0gzzkdr9h+BB7eQi2GrJ+bs/EIt
94PeV+c0ylr2w8ERhTGJgd+BkMTJfRG/gC3QUdhZXewbKLd0VG0WiB7eMkK6P9D4Fg3QmlKqxsQE
SDFSTLjDlL62L0E6eW8FeuJFGNgpyv9b7zTb9Zj3AzD4BjdsjElVVVrYn/LAXVZoXNIBn09AyxIl
5qBb77i3WinSczwYrYtsjw57M7HUT3h1pagVno4Tifbc0oB9RMfgDH1DW/j3YeDjAu9rcWsu5yIB
O85BJbJ0O5L2IpLM+AMMvZsxDUiOkP3r/Mtv1xPFJo/NZsf0sQxlXDtmQHDrWM0YcxOdnUKNCoqG
PVxs57JM/xwLabuyC0qc6z05N/dK61+RRCvm1uxXJPsevaltBcMPdUIdalHP8l570p9DrQN8ZtDL
NqQPrPiE/5Djb+IbKr5CRnWiOJRs8uEI4Q8d6NY58V4womORvOca8VmENiALQq/JHk8235rx2duy
RMb3VcQf/lA5HjLg68pjkTUre32T4+bn9xqQoYg5fl24TWmh9brlvRQTBkxPAdpu4UTHSpJXLANT
3n9duuj8CjwLNDeqhk1SSc6kyvA7zrBL+4jrW+KHns4ayeu1WamiolE4uWYfwH8sKTDAgxoYKnY3
clkvxhCGZIsb9iiCsZyCgtxhdAGojTxplTvEwjU71j+GOJw9KEUFCjyG1mbHUirs9GaQAG5sQsdv
3Sv/yWhGBWhvdcbJh0QA0GPz+PDWMp+zXNu0Xy24dIiMlo2vvLBT1DOaNy2NvRZ59Oy5xk8TF8MO
UgKIANJ4iyUsQZ7hEihJlhI8VcEIKHTI7030PJmkQJnN/yw6xpO35hppUKeYF6ifU1nBMXkKZKK5
SSrEKgivqnPvzbkKqsLqb8ENKKvD4j6Vl6waYUgpFKtVdeyB1idqma9fEkoTgbkDWfeFBTyCjFe/
9AzhOpifzQKzliqPHPalTaPWfMiu4M14iyYWFervaV0QbhYue4MZjTfsuTEkvJ0MdvqiTVwCEV1E
muqa8911UMv9wz11PUny73TU8+hE5SExibfINMJpxk6JwrrkjbMZhFNrMyOW4QFVCnVJF8EOu6ft
FCksQbXdU7WHUft3oBnScbuOMPdRt0Eg2nhkGamPuJ3++VMpclURw9Tx1eCnpZSPZSVfkG1rtUzf
LkEu9OOm7xzhhQkAXg2//t0bcVb6rRiNWEihCT7SQmh4hKu+Mp7YSpPkqqOWfWRJYOpZDJHEAFgM
6E1+/PyD7HLVHaKEBhOIK2sxW0e17C4uNxx291Tg0sG+6gffOVahaRmQ3EMUxtHk6QCqXtf43H98
lYtmsKHtJiGdTMzdfGDWO7dHwo24o1aIEPte/waEfnK0yw6VZdfDcGqPLqAMHmBpOv1rOE79CEry
k3ITFsXdbwlT75T5lH/MpzCTo747NYan+7t5KvKdNbah6NIOu2Z5aPOF1hfJ+/e1BxtQ2AOwXVw0
UYLyxp0zCJ4m/V9RUg3aTkTlHA5WY2ih21UP0eS3A5LUxE9p0kKdsSCGu83lPUPas7JfADSz98MM
I2dT3EbHeqnxtvKNc2IC3AUOjBubCzAz/rmuNpPYFfbU7GNWC483gnddZLcda3SJMLQJVLEpnL7j
BZtPnphAx2GppTnEjZq9JUxDgn7sJbDDJXutdtgW+lnCfkJFh39hQW2ia0HpV2aAqI/HCBa8uSPH
7QtNFeiNmLqzifv9E5sWR6e5igMU/29kGojbcIf48Jg6jFAvMzA/4OTtZTVQIkIvEzsuU1f7+8wb
9FM47apPV3+R4/vkqZjMN4CYhtUK6IgtJC8UjNsCcDtfHlVHHIon8Q6kUAjTzQ3ESwj95nELp49U
5SjxyUiUHc9Qu6iteFM34PfoXUnrW0MIBaLRSJq76E/tmYhgofc7NXocXTbSkIS6GDx8nnxc85hh
CClVWdkZfQWc8wMnU/APxSafH+pegBIA5WwA7Twts1tan17euNFXVG0yv2Si7iaMo7sBkENIvyDY
ohkuqTrJehXbXQ84SU7r6VaAHRz2si3C5bLQQQMl1y2CSGMma4YH8k++Mp8yzncF72wR8t5pQx/o
+TSgaiSw7BlZKbY5CgmgUSCQ5JY9O8gvHYDbMh8fc9dFa/XU8AUjEGBYGFhLQC7Yhk1F0W6LtBHJ
pL2kYFFqO4tdSjSxtw==
`protect end_protected
