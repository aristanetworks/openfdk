--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
DbDnCF3DCebGFs+7i75uSfVcaH6ZUH42ZCs/Fp6R+56qXrpd/R7/NL+loLaOc1X5WDEe3Svz+ztz
X7/HE6KN+EvIibWsjmlAEmoXyjSBm2IsvHzT7STK4AXJuJtC0Y0Yd4XbyJf5aQxnet4ZpRYaPK14
IGinPdedWTDabCJFhY4k7sMkWh4B6/jofvdAontt2G1iTUBbG0s4UduG5eIIYfy7s5zY17Q6dWje
i+2jKxFEVy7oTS/8Ir9C5g6rHYYwtPycTfAZ+wYSUvqb8LknhfIRlCF16O9pZfQYukiCfQaAxVvG
HA6+rTg0tbVtk3e0uOkoOwngVQZlmswH2dkv1Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="kU6rRwpXX0b2+XRsjfiosTwYEZI1c8mb/PhtHOfLNr8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
inIAPmbpRINvMS+kEzpdHI+F0EFXuZ6RPnWlyshIEp6cReZQ0mJo7/AbFcUECroGN6iyhVq5GtdI
nVFWJFK3d2NgWJgg7+nKUEydg14E2p06PCKB8tTHYoYaIdql3Wxh2LI/J0Vrx8PDqdRIN0PrGgxK
EnUOKD3phLVLIOFcm5LKlxU5fegE+iwuhJHvjNOoSLVsanaA2hRCudp8ETIsl9k374UQatMZW7G/
5jfPzv8rnmPZwdLI4Kjdmbt2x8SZMy2+2rdVSGDg119GqxWc2bfsvQGMHcXBGLYnliRdBPw1EmUZ
lirQl6Yy3LprmgixTCZhe0UQuAqxsbZxuPSQ2g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="NyHXF/U/dkYe2iuRwhP8eK9vH/xxE6T0VOHoVsxJzYM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2720)
`protect data_block
vFV4nG25pQtYdlpxy+LMSZQT6ibSIC6l0VHWEE416zUtGW5HmM3wTlGY018hsWpV/lm4cOCKo6+X
mM/0CLEkoFBOFp6aGSLVZWswuZjm5BG1qwFRnoIMxLqOdnhHrYO7WPpsfh1uJlxPFYVCLWWaXx9G
hzSfGsK9iVDZ5X7vBVpAT8ljPbVXOqFgVmKXyN0oBGKR9rejPnwktw2RD2eUJjW6hENlgmclbUui
KT3aHX1qPRytFS2JZFL4nkNfEAXj5IFZImGUYjMQllLfGEyBGyFd+h3povpbxcEEvFcASDkG1oRF
fn1Ry7ypidE8hXYisfMShyudJa3Pup3YpSVFeMueg0y8/sAWmwrIS3vpicLOUd5Ly2gBneO6l58G
hMY1GZwyjbefCaRwtwPgyvK6Bc/DoDPm+ax//h2QlPskEs0cuu1txqOHCejawXHSCWaQiKBt8vBo
2COeZZ57DR67xdIAgAW/+uBZ1PHws2DcvOYi5UqY6yRTOD4Xx1Gpm25qnwfIh63m9J+IAHOrt9ho
EPfrkKFR5yqg3n7nnNcn/EeTKXEVo0VqvFGnZtrPxCvK6IUS18bIOzkNkDQWFrcePnon6RsVObNC
GwF+5GgsSGG7vfJpZ7ARwm/ZX4DqdYdXf06iWBsZcifwynYUmilwjZhkmruINGhi6ByPEQPq0z5W
yW2Uuy19KNco/c6D1rCK8GCgl/SCugOLZpSmjpOgCrxNK2GQMp6WJfEuzqSRFa1EK7nTeftdoMks
9cayXJD4qxSjHoqr1VGyrQSmhfoOqd+vn3QBTMKQGXMl/UsPT/RLu6qHegMytLl2/4keMuXy9hb6
rE19MwDeGdTaPUgUIXNv+rwJtLDWsigJ8E8Yr7pDQ6zKvsj8s3xw8KZovDjyAn+J8SBX98giTO3h
m4jwAhGCc+fB2FYH5qP3yUD5teFoukJHG6XM4RHt4EF1+kxk4Md71R9IPz50fbYbxtmQh9CJj5cc
IbHFqRRN2lja52GGyfq+xRyP5WzVMtuMPkkjg+c3LJBUovJoyKUAsIZMWnT7ovLIYkzWOFBeKzvK
dUx6/F5gFZbza/X8MzWw0kS4HebLIqF/MX3jyI+dOI4dHoxzPqqaG+YJzrKf+XIyyPJs3DzWGW82
6IZ/qOPz3Tj3Oe3u7ttvi3MBuw0vHDrNex0sg8JCumqMeopvC1Z2kOKErk0NeAnK+H64A+3hr/Ci
8CaOeWHWFF6BrDg/9NdMYtk3U7Ga/gdfzARlo8T0GptODzAHWq9ZTForloJGuHHbUsO2WVv+ZACU
KJqYiPeVhpI/TmR9KUUUhtrSxNODq1NI2xF3cT/Iiodde3XU5PajJlnuVIRvz3cUzgtzG0rcsbbB
UcXVZE7n75UeXARne8glROyE1ivj5G2BlYKFAogASOpachEYO6fiVE/qpPwdDcmYnqa4mcM0aj17
Bhx5l8NHa2rDmdeorjqMMka4aIpmRzvLn4AkyN6hQQwjRhNidcmEoGOlBkgzvt5PDQdCeJJ0k6qS
uiVVm4fBRFzmPdz1i1oGS/VNeNWh/fsTrH03SSHCrS7f8a4fi/3V7xUalE9u28wnxlDOwKl8AQYs
4/MbWCAiwRBfoNsRBiuIl7A3NLffWaBSfRbTUVZ2YXEivOayUfO0qwKXZB/kHK2b210pxuE9C2Qc
E8VD6qfDA3D33F36NyIox7mVPQVj3jKWIFq16HT19tm4nSgs1kXrjbiRHpMRxv+IynZDB5EMwEFZ
5idIhRzXQTzAJe1tredZOIJWkdWKRwzxgrpgzqWP6ODj92phmtiinfCa8vRiCV/BbzkT83bhS40i
74E+1Qp6YM8JagBA/pogqBvtouBUVqzKKqOyflt/vXkGb9Iy3ZBLT8J7BxIusNuoq9zho4/ycDSR
w5AcW8jLWDdPhQnqdek6LWwS/GwO+LaCf31DJ3OMbm0/UIe8tQ7d0WjaZnq2BJguWNt7N4q6+mFV
zUzgwIiwmQh6UKXHvI4S0/DpRkIdqnFDyl4xzJby3mJ8QGagJFFfXpoUGiqYvlXxCnZh/TuKH0US
sWTHhqwe2dLZeYzQdLwmCDErv8Xx4Cu6RMDpIFdZnJPrpQQfoK/rhClPZQEvEOR9/rcyp8T6jXFn
3zfx6pV8ie/ucar9phI/g0fdpk/gQBFwqw8tTr7xy6aDdStPsAWUxaFhw5JulhQ9Ld+dfypjttw8
cqfEYslSeWTISUvdAYLf6q/6X7zqX6D6l/xAGjfRdX4iOS3pnbDNEZ5C8lpHyRDGl+0zU1FqkVMs
YSXHzMhBKdkiB6mhOnfTGYrhuWtpIfFIqF1P3KjixwT1kFoMG3DfFzKk02JrWevACjikkOZpGYpr
NgB2uxv7/1CGVLKh6NFddQ8pokq6DkoYUNHb0aN6SExtbt/HWWejTkpMekqQqisrVilruOVtqtov
ZO4GgoFvt37JHlRplfYncdlLrF/1k3Ppr6AnYrK/08wY+KQaw6BKroSqSD12y12UfxNzi9bIJ+6D
bn3mZmjTCLcBAvfw5hD3aLRUXWebCFjy1+rsICHW91h6m0RcunW/9iRahhQgAYCCWPWEB7H6AObT
Fv6cm7beZskS+LSM3YaycHP9pvvPWgFd+UuslURdTxwDX11yxg5UiUTJhoOr3KCaIByy/pdOivua
U5dBPZ9JAZ6S4+Lb4bcruMbWaNIqaZr5fhfI0KIVAxImxFBXkaTjduYTdcvYNGx16B1sIqjaCPQl
GkPCHP95lYMqxF85bQo38xkdACPxLivtIOGJhcEhZ0ORjDQkoagyHpr2hrBEpyhLdhSrX8pMCIUS
u21NEv2iXkt2nZFqOwz2J8tWLYC6p+D1fv6Fughrf8vDb595/6yai228N3bC15ggWG3oPdI1cWak
Fgad1LzBWja4+4kwRKid/DDXFz1zAD65gLORSJmqOP20ktt2ZdT9FAVu4ghjku2GgecS0EXbC22v
GOtI+rZZUqhD0HzKd7G1NFLvjmqf1aFY/w//kQluw8yY57JMVEWQwAo1u+RAij9dlUbCU/dyVzIh
bCekoJINgnqqYQE3OQm0y5xnomQKIrGEyqR1ML28DWHtOy7m7jn2wav4KzdIueJ7q1i2dsuRMCro
TkCRvv1m52KQNmSARpiNwW1jTNU98QqJ5DLiKBSm0AJldGEoIPYdWsh1h+jFFg+UVm3cv6DhkqiH
5ABVaX27jEVgZvVhI/TS07SxvW791+bSue2kBssFISfAPW4tLk9GMMJFyV/0LStbsgeyyaLDVZzX
kU6UW7Ci2Nipgy2o4ceflt+lypurU9rRmhlPHkcLQ5QG+jk1XXPmF5T9zu1vrj0wX8nIvOMXZxJV
w+GJK8Ete4PPM4z2ngKghd6dW3NrvHrgY2bf/PtkD5rS3Iul302sgyZVzsVMDYr5SeHUtzhRPysH
bWdDzqWbgwD5bKOBg/gySjAl/oDzxAaRtKmpLR+2uVhtwye/rg/k2wqorneOCIf5Yd0qv+4HbOGm
YpY04UJvkhYFrP1eCcEKI0trWBUmOWZI0PZ6CVhLAFf7EJMTI6L6J/4yjjfzU8duIhWjW6H2myI1
wXtXa5PSb+0bSalPto/VVIEVHE6pLkbc9g0L6i8Rw4Yw2q3sUik4eJk=
`protect end_protected
