--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
ZeywI4XKAfjeGcHTcJZu1RUI6cTCBGz5Inon8/trMkQUpwcTxkuhBQKv6hYx3hiOOtaN+s/zHFW2
8aHPJ5QcVXi3tGGxIgJHlwg0cLNV8H/LKJ6WiGPXwkIUufpzoSxm3o1ZHIis04dK7fw/CijLXGKo
tgu+WmF/w+k2owomTG5s3Uc3D3zsLtoE/+I41n41J9GsEEcKYRwiz8bKCgMBdElhg5PDhi7msxe/
ktujWSughLIEZ63WnTjV7IXKhNFg7zrBHiC9bS5O01hZWAYo3j4+ZF1wC/ojccpjBVX4apbjRNjv
aQDkZfC/Mn/+Z9UzcQkoJRuYcW3n4jc4IGA7YA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="i3ofl//gzqvJVfleRxQq/7YAHlNCRpifAQf09UbuBCI="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
SJpi2DxocaOCncmX+7qitgET6XHXjurFQpMTRqhfDyTNeA84Ccnc6xFEpWe7PUeo2KD2lHkwXpPk
71C0fBwDCS2+JzOLt6oZN98Tlga0IVwDWydfGalRuZrxes4Rm3TYmzuObECYoIYV7tWjj4GWizuT
EOiRS6Q6N65sibr+baiTMODM3X7rP+sYl13ta5SCEq1sfonDauAB2Z2YJAUK9mWpMoIbRQIahwBs
wQCRHjLBCPyzt/5op++fWI7ATUviduurB2GteI9MtOPXtwARg6szAShRqMQZNb8S600fUgs4NKQv
gYtow8qhi9sF8p9n1cJiLw3TQJNYvS1f6S6NgQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="uF5eq2X34qV34ZwkWZsHSo4WRHwIl9Fmv0jABHxUM0Q="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6704)
`protect data_block
DNMf7Sxe9y/2ODOsNZ5+/xSnm+OjeOHmoZo6ipKEQYtL3QC545nopQH/yLSu84pQ0JjE38supU4X
CsYI101siRFCIh59NRfDONOltoY2DsBFJsI6VFqDT2XARw2pO0YvmFliAJoLrWS2xzTpWER8zfV0
wBD2ROYNW50JTTc8nji1Z3ZEP+gC4+2j6DrpsomB0WxwiU7PniqR+Wl5MxlCClatWFBkUdFE7HX6
sTwKmuzPwbupxZosNhK9avd8tctwbS88Mz5Qnnw0Hzk8ItRQF9Nw/PGgV2bVPb4J5b3ctaF/BMsb
Ca2kqxzppFe1ferkatkYYkrX9usVhy4KtZbXlNbBTba9sMcApN3ksGvRyQBZv7+mi3JYIi188l1v
45ofqWncYEK7bxw+m1GH5fKPVSycolVl/st3aR+xpyIr2HyZYxP96kkaLN7Nmau+neHEwdxKL9tU
g9JNFJ9ENVWNlE+Im/g8jgAjVa/VwdQtm6Vo/rYSEyvVcf37BlyBH2zaz8vJz5sXRwJ5MXofTng6
3oIcQslsGxZdimOcNxE0CMDC+eJ7mTYc5+SlnKtXGBWVMKkhI9tRdXLAJzqnOvvz/bqzDJ6nWkAF
kYSrCJrDwU7BWU3haXPQFEZ09e/vJYWuCpcSCLTk/z1BgkZqovj2CdNA50iu4f2DD3SnN9MWESiI
q35GoMC7Aj4z3oFYeUOCPlLU9VomE2psyxhvQMh61Cfb4x/W7Hi7iVQP9JtUCtWh1WXu/r221EO0
RmWe3GiK0FhcLB+QOVBxaqgJ4/2U9hT8/+DAKiQRtCPsGlXJ9is8wMq67As78xOK5illR8Ir6Shr
hcB3Xxi8u9CV4xcScpKoektSYteW8+PUH03YYQx/CYcLg/2NLBpTEhTu5DNiW7BfOzVCufTRnN7O
8NE3m6Cj0VcOO5pfYM2N+0vo+86lmSDtfXkbr1GHPkCXbxBPj8UVDtLeZY0MmyzXjBKEGukmE+lM
gP+OfBPIPKuZMqX5yhJZ4bTRvHa4Qd8NF3mBJgb9OftYHSfF3sxuBHuInkZU/kqVPALGLqvPZawK
S6knla7BT4JmCa9GVvXHN1goGgynI3wW2/TcWKvqp/lc28zg+wG0PspPzhZOL9SZ3dHqMNDKewrx
DG3gd9zJtP4Vhtz71gYor3CdklGrupBgffXWG0/+hAF0aV0eR+35r3J5GdTtiluASsWSxLUEFJ/y
m9f3hI/kSWLMEuDTgV3BfjGtcKL/n1D5hbw1T5H/FuHeY8kiVyRxNW+ALGsyEqHSD/asc6XTum7T
Vd+0FO6GsFLmqQZLA9FWZq/U3NvDmBZE/3DC9aYpqhKbgAHuqBn3NGS02iDKzoBxlpS/Mbqby7Z4
R8k7egtnAQKkYAPkSlNxqlGJft4KLkvlxxNjStpysa5XhZ2XSHEzgUThl1zXWrjTzwZdCJZTA/pY
VdLI/VHWMNCbKiBqfdqlA5oynqQ4iApS5Tap8m5fVtpbPHFlTdYkqqdKMk3Yw+7CasOdxlXwHXxt
XdNg1eBe3FvHFaYVLYVOEwoyTHDuVz9bCLi3/UIX2rM+ZkeDMV1Aj8LON3p4WZtDnC+Aot6obUmH
DR/PVzhJx9ELK8f7KFjSRQfx1bvTHTnLLdDj4tJONBdFIyN1yfb6S9Erw01LBBPIQzslWyDpvrgt
nAXcWv4sahuP0C9ELykfCvd/Ais5FP43twMlhfv+A7jtLwY/38eLu7VWtKQRjWjHfwKRzNmBTpQX
f9dO5s3M2lce2+UntcpAMp7mHQP7ZPxIy98j99bDMI6vocoJblTKWcdef6za78mU5NkTgplRtshw
M+CAJYRZLDCWOjv7uVO8wRDxVoQXbedBsaSdegiwiwQgTf2sf6cmujtTPw4orr2m4P6pxf+IorBT
LtwRJQoDT+1hhPstSU6xh+ouFvYmvFRmDS4Xf21s0CCT6SmGsA/R0X9hN+ukEW41kf/+mXsx1WJT
veKiVtAabxrdnoksPn/n1Qq1ArabHOdHdUV0Kpf2ubmEsqhjAS6qSb+ewNzFSNfrf7x0sGwnRJeH
KgK3dB5zjbWDn+q3S9EQ80h4XptE8PpVYiTXk3KaC4x7OpviXU8/QHTYUSQGq7riIW2JSSS+Gk2d
J7TvrRRJH1lGi+5qUHgy9SKOknaL7b1l+91V9M20cwhfqbPzlzL7YK+byySeO8tNItyMXfM0N0qF
l2Rw13CtTYpsqGF38bbMFWdagnKtkwudnbu0PbpIe2iT0VNzLFSwy0sYQC3oR7xi/MOzl2EHLthm
ZezVHl+ZMvKNs3qQ+9ulJQtC8ynpJieYor9ibCjeL/n4YoYsgbScd/ObphltLlGlGg4k4SRx7opo
TtPZeEegYKpO/DQeWK7924zg2j+Jnezeidp/NLolPfvLxrYAQ9NAfP//iT9ZPnv6DOKcaoP/lKT7
Jc4OyywLQhLgh1XUr/e2RGqJW+zotsRwVV57FMt6UBkDNVYFAJ4TXwdMwXsE5lDaC6MIoXaPKBI8
atGskssoU/kRnkXhGr8IxwrmF4oWIvQGvk99dyDNMAGwz7hGPMWyfisjRo+iMUoU9gKEGjFBkEnx
5cBIn/ZDPNuIqL2GANPkgrpyGmJCkgWruZWOzTiOk2PgvPLMzsrX74U05WDsHoQGx8b7rDu/USvC
moJXwvi8KFOJstQ+7SO7TzkIj+ynBquX7CQtGCenNukKcygtzTeAmiSRjiVzweH7z+5v49gzpYkF
++FZCKoidRjgbHpQnTw0KMTX5HqVCpwlvP3/JGXb1l/2GcA91GaaxKsBhJogmtRcJfK1tbnPfb5C
UhmTAT0Vg5RIl7Cs7L/snT77pR/SaWe4SMOagsLAlQucuFiTyprwS52quZDhaJyHd3O7U0iiIzVC
qflTx6x5G3p9w+iIFtxMTI6cMaoxbltDVIuauLydGO9eEGqWHLr2k4024zWXPdQKgGM0vfzOpXKA
2EsxblleCECJ8GLWEtc/Rn7Ol2at29fqVeH6EihABuiZs5e+dvOCiNMskoW+P4++St7zbnQPgG17
V4Y0X9NCMWw3IEAja3DpRsFBW/QUcl5uQM3371Z4sgVSz/8EZ7vs/XLbZTLfYUjAkMp8mUmGQ4wB
AMi5D/H4vmcfOW9SVJeAxdApwyhgS/Ny0VhE89UFFIdUqpvhPqaYjkBZUk1RqIMIJQniGiQWvmwS
a+9XO+Y/qbTqBYJYfW8fyggbC4VdXIqXCBEnxvvItHotE95hnimtdyovtopw/o1unn0w/RHjKceH
gkBdC1sLSNz/x2q2zM+yJHgBqC/tLJR5WWD8nAlGfcFMZsctCJV+NyGBcKzp9Iskq0gpGGntJgFM
4xXLQfwwWNsTFxADR+mTcvM/beMpiKeu2aAjI2t8bSzJH9XAlGICBUfElC7ia4pEjXHtCqu7Z4Jo
G7PesPRuEGIBYSRp3YHnSGKgc7iIVMoVSjbDY7uhAIPQtUEltCC6Yv+XfwpdlmvqLXSlyLaHTXdV
GuOVTOwao5wURFVLMkpGHq/ZRvdST7pt98dMyvxINV94q6osaaUVyOB5mzqPSF/rrffa6VUuMIrl
rpuShVa+oiY2w8BjSCDpYng/IbWMrDKw98Rx0y5R+QMyVBbG5S4BC8nMLq/Br6x9nIrPnNqnQhj3
9yajoJ68ZrHG5N6232YOpmr2t0h/s5UzZf+MXuB/FIrtMETXMezCcvVwCLWCEie/TMbcir1XElLq
xfvaqofrz6kTv36XPSx5y9vocuQbxw6wDSdMv3gggLBKpHiTy2wD0bkML7jHOouYPhLnm+zBRu+J
FKn4Je40rYv+BcpI3mF/MNSGp1ZPqAljUt8Bo8LaO/b2NgMFkQjCtPtC5CVZbiyrZBt97XBMdGpS
vpkuQansl6I6yjxeUSZC03X1KB8YIk3V6Kl8BwDW6PWsYsijD0RRIPykZb7te2A2Oskbt2sgoLxV
wNg9Y8sK1ye9xTyqDK1Jw7hEH743d18/ptkUtQuy1g7hVBSkdRtKR5QXI430XcNT3oTVvUQsjp04
gfI59DdmSfoMU1O3NCDTMXSYXhRSbLx896d8DkXG1YlmzneMbAG8afLCcIYzv+ksZYbNbHGyVVpL
t/q2gDcyF9ZMmDYt++13PbtBJ0mbjR0fr7m7Cbo2RIQef4fmwR+oY1OT5APhCRLA5OrqP0ZvcFZ/
mSL0QV4AKfXveCe7Amt3me/eXkKZmRN4I7IEbTQpmsOLW0vOzH4KyHESS4bEORbEGMcuu2NJmjC2
fzU0FXrF20Z+7Zf8z+kwC9DHGcnhsF16fZvMGU+pFg1c+zDR4TkAC8shUTGIHvEPi6TQ3TPr12Oh
z5kH9OzyC8JPowR53WiPT4fXFiRxVVVdF7CpIYUV3KQ/89Xh3NRH/I6ZFnQQrUzJNMP2ICC1J4gN
Z3Iy5jZUh2q5d0dTlgT+jGYij/06q0FCfF52K9rI4bTY/NTTb6Hw/bHz9l3KPzfA6KzyfFaTfiB/
AoI7QddNx0jnAfcvhVIsqr8EbIZF/18GxI8dabZ9S1NhmvSdvCj0c7TJFyaXbJ5Jr5MFuzoW/9uT
Lee1Ux17pIV5WyUvBOhlG0ffiQ/j0zB68ZNSNKJ16YMBCpWSCwgOokFJ2G8tdoVu2tqVzbAgNaNo
oRcLg98CN0BBPxUY+GvE4pDBjcvcDFka17rIP4txoZI3OibFpNyy5scnpCIJ8D2WEzfn1Kxa7Il7
okYPCLtS7parImpG6DFKd6eCYvmuZb4l276S+WmX2fbaidr1muwsY+EgifOFjd9R6VoJH0vqFqlT
++vACu4yQgjsHi3Yu2EY6mYq/eIH2UqFiJVgjitHKxPj0PfsYSNbpVif6n36glGH/U2A+1s+TouK
KzapHbM+AAFaVrDdR1RULPDCZtQq4fkILRfW+KojK6r+ytgl2m+gImjctzfcw6/rGSarpzw/79Wo
2N7zMWzpS6792i0mCMCz+0DtKXHfgSIDcNWkPKQAdN84cEDNtuBG7Vi9bQs1GPUDV/9RM9Q99KnQ
lXbI+XCBbkO1bLVri0oJH4b39/Qb3fhuz9uBkKEvZBCAShqCJv8/8+AP8hofjTh7VZ2nUXUnbBF1
3yThkcJIdZvUEwkMEBxoy/l5ZJ8Gn+7azIDiKKiG7P3AmUgChNgWHwaFt9hN0Un2LDtRgSEDA8SD
JBj5aN9RhyuDsulmu7X7sxqwxEswmLzIihUIQPMkD3Rlci7Oq501r0K8pKYjtvqf0uK3GS26iFcm
EBnKLK7d7ZyrLcf8FHTialSJssqOrEXxkTAeV1b2I/7EB5i3jOp/22OQfVc3cJMqIcnjuGO4CJsf
YHukRvp5AL+yCMkfKQAromCtQfsaKKOTbOuvVtTCod8Ftx7NHxYW8ty3bGdH1sYAvCahXFWjek50
DVKflDi3i0TGz6BpE2/X0RZHxhjVF0OR756XRckUDeZ7SwLnkSFKjx/o24iMSvUArz82MQ6FU93t
8wvAszmgxfx8LflNdzXA4Yp8wQg5g4iQCX8eb8/lM+geh0ZGEFuuNd5tm1rP/z179uwpo53EDa00
9G0G2OkM4ZCV357oJ5OaCNI5sMvi7XBsg2jEHx0GwWasZpndAeWU64xvtIrlEDl/MV5ONcLr/ovO
39srNVfMFG9Oh/NM2S4larcFUp0whg0NVmA0gMw2pzL14y5870VpJ1wsINfW8ODuPG2ExLgtfDW2
qT8+Pq6SIn0ccs+nDnhjvBxtAlnkoLc7pIIvfUdHTt7jX0fi5mxhko0rM5PGTaVzVRRtfRBXliPK
KD6w+yiML/lWQa+uPHL9g6MVUjptEnRBOIuOROjJxS15jPtYE+L0lUgevcddXqn4Nj83V7fOP44k
drKfNG/7+yGjo/S5KPtzFjmbXzT0YsJZPTbut06HlIgugM//PMdf1Z0SxuL960sACbIW/AGUqrYd
R1lHA7+Alt2pcgMs34Z6WSsuYZLlYQkTjWDcmKpNSKcsPcSQ40bmh3EytBvSe0e7+GNKMoLK8LP6
yn0V+zT/YcV8KEUVp8XP7ccTwS4K/Sjs9MYwoJcXJlMnqo1GYeUDmlxG08O3jSxUAfYVG7emBoSv
Te0snF9oF18Tk5WIYIWiX5B9l0YIVzXraVAAbyfa95dOJhYSzzckgSuSdgjeKVc2x8Ss/HipGHJU
py55jiGhKPutFD6HSTNshxw1yf1ZnAGJ1h1qmq4PJDeitz7tR87me6rMg4kLl5MbMXC0v7M8szVv
9cMHCwWDODmKkU3z7+KfKlpj8YdpDF5SkbLZwBTS8IhpW8Ovj0tPiLHxlMC+11oP8pNqPBMM4dPF
1hqUWXSQXc2TStqLKWpTFpDzTUcyNgVT7MUH1HmPK5cKYAOmzybaXZo/LSLe+J66dQ44ghzBKXKk
UCgVbTyigSfr5Gb2jYdoLN3nwwVD726FeD6CAr2U7oqUxAlvk99L4OvNR+e0XOMA+RfG8/0frMy8
Q9LzNTusxqxT0uU21OxKdYN2nGScdCNMREnM5fLtO2xjS+ZjOoI+pen4g9Zeu3ZodVxc0H5bp/AH
mKRzawUNBmLTiTzD4iW5R6Rlk98ZAGl4TxhcqYNUSmFU+YKRp3hFuvi57NZNdxqVQl49sPPY1JW7
RAnQiMoRl3LM8Mgg4TdFCerRpXQARvIzuGSbsrMWQv0i/CLzIwJ4fXdTn1J3wZ0U6E7mDW7Sd2Ua
W/Qfimy524yVQTrVTeWo5BsEHdhcr/kGpv8+NsuB4AEnjLrU7Wl3QRcRKEPRw3ralulpT+zNtewb
2ReM7ukQh9gdUOfFwblkPXVYOKDIjy3c5/sXtUJn+ebPQDCo4O66q2zoY+HV1hs1lD766AvqcgQN
VmLgNtPsgZpzPDgTVCzIAo55f6iTLjPIvMjDKu1+b8pM4/2eKKAA/2K0jamuvBtc+tk9417i3ewy
UP+a8ZE/KVLJlwfUFisMPhnrOg/M9b3crw3s91riTxqp0YBplUT9Kv/1MyDLVJQdgymKuwuXR1AZ
qjY5w9vBxelF6K5fXob07a52j4aBNK4bhyHYRv6HsPikOiIPGVQYmns2cYlv4c2HTIhO82V7rdS6
NYeo9r7od5kJWFY17wKcchSTopqs5L0GadBy2sP5Y4KBU+kPpv2+XHEV2TN5rvw4uPpQ/FGXzQnL
DMJ2WFVdQHUVqE9bVwpDbHNIZmfISHKzq+EEsBMn2Ts1WKmS2GuDQ10xATeVQEomriytHW+M7xhy
BHBsHn59vvOJwxkt6wNsYO32AonY8Aad4TTcge0vHMFTg4YRhVpcfcc6UYCSjvStD8YUdlaDavVI
DVxUFfxZm6uhfT6wCb5xPdba3dzFSUx27MC4e0RcOb0Eqz3FmBe6gHnGUoFK7vjff8qftZj1r0V3
JfFd/uDX7REt7x+6jPxq/A7zYRyDqYx2OrrFIlEOcBifGbU8goxmWw6cfh3MUNRoaqmbGgG6b6Fl
1qFyZywElIJNnTfarfX/ORkgGsuOisC/NPsHzYBF01mezvRjkx8GAdNlTqH/5dXlvI6dLJ4mZTdt
c2iUJwao3JJmd+g0udDQ6Q5YOHmT2yGMv/ro/3CxbXcZyADyaLeAEPByYSqsmTCyvKGmdWG4/ueM
juzkCan8GV50L4aLDCfJX85yvzqt7zZgMqg067kqiIRAmI+A0e+HnP5PIh1q7PB+4zHIDVaL1Snd
IXVZGAx817iWrv66HZLRKFkjZUG67jZbR+iL3JQrsJuWSbnr7JiqZyNI+seHZBoNWaMhsJ4PoACZ
B98TJvONUNmscQfHoCeuh2JJd8WHRG68JY0PIEjrjvZiQu+OsD2/NkuqtZOQ3qU0gAhJR6oJWiKP
orj9qGClEjtts9IywGcMjxxPE4zIikoOy3NJKKy5reTEt1x+sSk+Vv+yE4/5ze31cGsb0aXZMuCL
pFyyPIj+ps455kmsc/NFt4GTgInQJeFz5pRoiqPiQAvVVAJ2r39kioZfpGM4qyyEdpUedOIj8+SR
E0IlWZtDWI6ybjxiDKGuTfGK0L1nL0s8MW4TIBucwXnxt1/Mq12A50G5ZPo8btc0yOqU5xLAwyMo
P7mNiwhsd/KIsfrVtghUuPyJU61P+plsgzG6zWQdlVT+eUtUbeR7fQvaQUpXLbu5vbBk7Tu6/CS3
vbFqrC6//BTpyAIsLzN2oqYlmK1jdPTENSxf8EmkRGlMMQYz0zAV3AGArGtX+K4IiMyoZBBhWlrD
1nELqGdFXFUxosGZDr1LOa8rhCdiTThY03GVRCPLT8oOCkstMALtkwuauI5eVLayL3bErxz0oBws
dhboXonJxQsWu7KqMC1wLW2AaPR/ItNcNQkJFdih0o+jC4GXKkdTU8kBlf/anMfCX6hqXwcnxjt5
6et/QuwMSOV3vIRBTcABeHsBxS9j8vXiBO/BFvxtprPAGtr8i8xgfBYHLDa4ef+CmaSraFDDvRs3
ozMNe4PhrEQRyvIAsbCpvPGE9OAHRuswOo4qFqynOm7n3hU0EMouACtj5jLu8uBeA/8vgcXXelyp
JqNMDW53APQOcMF17/5OerDxhBTYkfrw5ces+TmMdomGZWgJwh5z/CJjmMkstyyK1I99w/8MVb4H
W8E83Pn3dm8F5tYQ6nf5v6FgxJqFJsu0XXNZq85UM/QhFr98adImJ+yJqoLE00rLpuJiFvMgBr7J
BgLIMKvBiORtKB/DL9I+MqQXxvSgtZcGGgW9sVfeVtew9iyUN07kmh3R5P4A52bUscohg66SsMBD
MpVu8/RDAbmYcEXW9QCaicM9n23qovneC7M2LZpOqKe5/+OiZttTxOymREVL+tilYVO1gNO4OTnp
0I/xhn01hM20k+Pxeua6goWe20eG0nnH0ApXkgLxsgM9zowD7CnHUTb15U7kFi/PWb+/N7mmDUM1
koolTQv7fCpljr4ExI6eAruw9nCXjTPa6GH+9jmtoWPuVeY=
`protect end_protected
