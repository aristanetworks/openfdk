--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
oJGy+puYue82gD3ynio1x2OKpnoNtYpBIVtI+nQCn40I4eb/G8dKlRdCrHhMkkAyFwI8rzVWhE3t
qY6d+mfrnGluY5ycYxiS0CPfGbidjj2EBxLdVbtDPvOjK5mbQOLNiOgQadCNk9LK/Giw6MXZlGZe
2CcrYRXVxGL55BFSv1Mz76KtsfFW6TeXv87eaknACI9kUvqHf8WIJ7oSHtrCl0QjszG9RX7lqbi9
4LeJo4lhuh8GiZMkh1uf7M+Aqflz1SoJ3gWi+RCWweD6SmjQynzUequtu9Aw84mzfvsGD33Jxgo4
RSiJNMM8SueJcRxoVqrdbI997WWno/C/gT+sAA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Lpglsi0tBKulZSkk6grBDD/0WKIjBPqTIHuBHjk59MA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
DHq/tX7oKAbaA8/1f4ikVIwG0X66ut7MF3/Tqli3r5aLSqCaf+soIyV58EpsAsyO8YGbP+G+L8To
GatVxQwXneM5ORLvg2zpfjHoKi+lZKImdsqQIEMNzpPAaD2C1rhRNFSNhRsHB7vMf5z4nn0x93EE
jryqAHlN/h89h+dhGOjXQ76S9SgA6NU+3/j++cPk/zb+PKxLakMGW22AGtmOO88gQ9JEWb/zUBPW
XGI1bJ8JLzE5GhHVCzicRbaLhz4MwSQhc0mCxbT27ukjxx/3pxoYRcZ8dglr7Ck28HV+gUy/MwtL
m2pC4UVVP4tJDMEu+A00xApd8XOUXOVfUbcPlA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="3YacBw4haSoGp78UDY2NxFlpMawzrP3y4/yWxYhJb7U="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 68352)
`protect data_block
ALaGo/4gy40YZ2eqg6PM6YyvOczigFh0mp8HXOQGrzmF0h8kZN4T2Qs1XzUTkC5PW2bpeUiqdUy0
7/GP/hb6gKaPvT+oprW6014NnE0f/moOkZjy8OWeEErjOMbi48IOWziomUIiMdWBC7ljwpfS+5Sh
WChMlaBm2fdTwu5vU/M5BEqsnSX/Bfb71vP5g41IVtSuUF2GuATC1IaEIMVtID/hRqOf9UBdH4bv
OP2sKBStEVCJUQavrtQjAgUl91FAlMzWzYX/P5yq+P+jO7/Slbj/YHsP9PLrfff+DaRlMtDjoJMd
r8k4yjdYw1wISoyc9dDCmLEd8H3jJXVVLtBFl2+f8SCSB5CFgon2/iU8umYnUUb6IP0w1M0EjfSN
6cXE+NBoKQ4zsINoeUCtNlix4VauYVJDvnjBWJNs9Evim1zcH75CyiY1ZpKIsKuCILrHxbGlTyph
UssN5C/KbZkulGuM98sf2/h+0gQXLXTQAs5T5wJqMoBI+A7Q1l+mPFswTXcu9mKSN1po52WhpgLh
IXgaXueTS9e1FsKKVCzweewnwocJy4oBe2czLoGDlGOXiU4nksx6FCcOjedNvlYVu0MKoB1hj2mQ
7x4ctJwPcxw7fXlusrF42gaoVitN95qI6l2ic3Hsp+fy8cnps4YPOCPxiYZtpJNrG89i+3ZrWZ/D
zPBi8qfzscNOgO7jf1N2pH6qh08kk4zWqYSPNr5LCh5DBxBDLt85rCR5W8Fy97vb305IK+kiPpVw
on11EnitUIlAYeh8O0rp95mDZjLg1WKyaO68K5f8LeAKY9P5Yg3qYgyKfbJL47xcOJSPA9e88zNc
betH6HevbD375Y+cPpN9Sa489wXAq3SovfoH5BkOXgMOZ/G73Yni8VMnSpsSRlaZoOwDlPWbB/yK
EVsk8xgFok7WGJRlVe2vIOSyvjwv+C8hBNUtXrVJ3q6u80bWwHTTWiiw7UwbY9VE6ZVTgqXN3y/Z
X6x2jr5LHEipksN73iGOpVpNDbnVqlaQ0jwv/QWbAQyzaTVckFnxXh34flgwDJzCrgHhCLUSmnoh
vn/yH/LMZFdbDg+qpmw68sJMqvT8MltAYFbSSuzHBZWIoBf4qWzPTAK86d+giLQ3vSf12yIrdgu7
R68IVEjpYUowvSHUEItYUYjrlSNYGyO/kWEdpzPY2mm47IK1MMdVqUJONYC1gktaa2KBJnl7G//f
RbtNakB8E4Epks7NxqkfMCsbiQKxr8jlQ8tBVmiWyuEk233JfJWNn1NBLCKMn1pFJ51BcDk/GMfC
Y0bzpxclcfj7syj+67DxQhhIjfCyohMqNy9taBeJVv3EQ42qeFhC8AYXtxh+cEUrOpkTjM1Fe09b
NlwJNYp+kbedef/bDuqbImGCaWGW44urfDqS3R74w+jsnV5phP2Xr8+CuW2v9lDHtA8nweUDgKe4
f/yihdasOarLUAk7lgn6tWrQPGs03bHcnjOLT+lh2ncwzT45Hmmksz8TB0gchh5oTU73wD71MOe4
gQdLZNZmZf+d8buwfpuyeFPHStmxNtgoWiAkKNmGYqtv996HRXEnlKgdQ3PdiHF/5jZjwUeCRTG9
SWHvq1JjHTplpylRFzfqIJ36AE7jjRqA+CzIgwhiSnfNhU3UvMlQP6HiZUcyzHTz6GlvmD5SnWEX
dV4jVt8dpHkMh1h3Ppef/F3XsiBWKAq8tMyTP9IWXZfqdf5ooAlDPL3qT9S7QzAq9H6lmP/cdicP
lDlyhoAqWwN37dPMeQatwAogRxDtDQS1eyrmWULmoE38mGA2Bg3bCaOvftVnvH39uhJv3Ix7Tor8
yBMUt9wOeXNuEEYXspIe0gNLV1zOXuAPTximj666Axcq+Py225hWnqAx5WepGGMIMHW7dyOMj2zM
9jdz1UpFJRjTYmOCZ8ysYzE/8GBNrd2/coT8+GI89s3tA3+x8K59uyhygtRG4Q/kI1iBVncjP4d/
mGdQiWlKU10GdS5kBhGDtQlhyO1P6spfQy9wtC70ckyq1zQmBxpTvDx5qPMa85iXm7bm/nieJ2Jx
JtFRbLg8NLOWfQPjZvSiRDs4AsdlynJPEA26JGKfTJfg96HtKujZkxNCQsVLTixYmyPn5pNE0HEl
ZSIsZv3RTKqjParaojyNEkCbyU8SK/7qapoZwF3vqgaM0iamrFU9xf8w6jOuENNt8QLjS+ljFkNx
nCHdP4SDJ6Ehj9y1EO+Q2MRG3GoAAgj3rmYubE26992Q+gHrNZAZovhOw7ZWfrp55eW7itUHiMFr
ynUMiAh7aYhyCQjfVIVIEK0nDqSQ5e6HeA53NduTDHdY1W2u170uyTVyZeNrsC/Ziz8Ur/LhV1ky
VNh4vGFrCCihn/U/0bqO1AmI1pslMchl8bUi4TeP8dQw7xysWooA42Zp2AEgc8YLC5qNiSNPA+Zu
DwB1hNPFfcLVj0RhWP5HoyTUdUre7dzNzdERHPG9hbHU070e1nXebJbrQBYGbiNzQQBtG5kbuVtT
zETbImxl56AHzjUmAfScACEJWwzSP4C3Y5bW+1wjHJy0X08VstLcqVv783cw53zdBDN3wXNO6RsV
NOOPvimPdotDGEPOW3GVDI32GOPeJP9FCSHy7rJ37YC4O4rnvkQGEezDWqm1jSNhGn6YooDQF0t+
RpYF/HXYjm9yQixwuyzpqC3IEM1fPN/5wuUVGGPK78tP4ptAPqvFEr5S4+sYP5OeE0wGtdDF/4ti
Cis8MukgopkOzLbW+4eIQVMo4vcAD8fsufInhSIPBRMk31533WLRJi5m/kebpjC44I5AZIq4dY/Z
W/vUJ/j0qL+iXWjsTKaBUhUPVBhHbfsMSg38M+dRFVTfPMNUBon7FWv1xPOmc/9pQlttAFfAWbDV
IfOuwDmv7Q7EKXiN5FOKvI1dLahPQhhjzZtTgpG2D+IxZClda+OIFQcJfs+4zASOaeBSqvBx8e7g
Wf43B2E8HLh35c+FRDVr/nbBDrwai2T0YCz+240nFBIWGe3aW1rU20Kq8is1wn9GMkShoL5CcQ4/
r5CK2PExkcKAFJL7pVj1O2m8grze5iAgTv2UR6plQxxtssksuuvrwdiPVuK7BgrAgfRXZHxJxLMD
vTL3rdttyCvrJOtKMgCJIv+j1iPjyckcf3aLhWu93dWsrAMXDCGp2ZdMIjHvx5DrvEy9qngNBQJ1
GmkcWBsMXoa6JVAaX8HO7Xme/tVhIJIOlo6RYuZrgx+iFFhN6sNi73/E4XfPgCGb7rzMUkvrwIfZ
GVryRoa9WtVSYiDWKaNX/Pr1NiWH8hHCdQiqCS49Jxt4D0DSk6uw+S1+0WkDe44K54bwrAJmf73t
mAHPVvzuM+Iw0WcygOnoYFemMgh2TVTOb3Tb6uF6n4ou/hTrDcwG7CG87zt+TNihvIU14kF/5AzS
9qMU6pdzSB0zlGKu+haOPKi81M31BTsPSjizpPnAOtbpxVR5yiBYI+gCKDRL6Ib3/KQRVGY/9NyS
jDC+opInxOJqvDMvfVgxzjiGRNXggn78ZMYNPa6soywD2EX4Hrn3HUBq4dnxFOpVDvkDtnYT+1Zl
6mGVIy1Q9FTy2CjLxVLHrAspZj2kaaAZ9grQems294MN8RMY3DSH5tfPYomDawFMKZQTD5JSm4Xc
tgiuwogwJfJS2stkhL59Bkdhpq418CcXJJ9m6axBx0P5HQeH/cvUKapAFhIEILehOj2rme811VxR
YGV5qB8lD7Dg3iVHgH8HPef44z+MpEZQRcvWTsq/rwgC5a7BO1DO1irJyYYy5vHgTmRkljH+ZusM
nF7jN1zTBH1Z5x/Yuez1GINFtNpVI8lp/ugjxEogZ1QFbj1jQWnMb2tddGLHhYTzyHVIAX897swm
s/wsvZQMnqqoi4IKaQx4IH6gupQOVTPDLkxpLzXTLrHBc/wWwqLP2wXN1fyWZFZ4qUY8BB+B6nUx
DEtaoMWCn7tA1950WBa56ADbNdv+7gR5m4sCrCpbS15nDtGvKasColLZMLwhABrOOjTzYfnT0H7s
m0Xb+9sMO59dYsCP8WbM5Vl839jSHaXhtefCoZiLPR6A2UDtMit3AqeMMTAAbNqur/xd0ccAwAYn
c5kxg4U2kQwJtERoEMMQV++5MqHWMSDKdzSWHGIyyXluOByfC8ctIZOjaP7QIKdWeIYEsq6PV5QZ
5p28BLtzZcjmkHdgOblBVV5Ik4w/p/xo7ZxSHm9BDAcKhjsT2KHLE29zRdS++O/F2rIuuVvs63F7
8r9nCXUxLqjAUcPMHV2jm/voFX+dEb8cFzu/EquahOLsNkP724vY7FvquKd2ELCMpib5IHpH7Z/2
yPVQuaqASwhqtV0GMNK0kQGViAMFDdpLFJQm4eSMvgO3+w1a8d7+Qgv4UQ/VyPkIm72XkdAfMYPb
dX4OKQnu9kvnjfWKW09pBskB3It9STSfN3x14L8eHH8LjhlDENWNo1+Xl2//8htWiYFY1M0gHNy0
tlnyBXGb+JJH6yZsVB/bQjK3MTYL1tECY5Zr+uuOIAwamMfbrezGyBMKqAhrBdryttjVzUezRQWO
fqNE/kX7I2E3qHp0dEryLYPxS0jLner3UOO/5givPPZLsfk5h4vIUdrFu9gVeY+Jp+pLynzJPu1B
DqJZSfwazgeXwwYMor1bJt5VcDl8LNybsWK3MDgPJ4ZsFplNzUvcD04LQcmKmk+p7yKjx5IOTdmb
NkOLQ5d9Qb8zevDhHikgC2lGr0jfMq8L8Qca3aJGHArpOKY9BXLi4T42JlHfUOMFbTyqxlBKSngi
q0my6LvEq2NmllxddeH+7V2kqgj86pYbJkPRAjTL2jMAD6L/MCgbGKb92iIy1PuxWrg/Sp1zEjB3
n8D0TyMcH9BxIxBjTMzlNmbvn4iIKgoEjGur7arm2MvgQagClMtHXLlIbSxLjBC6Lyca3ff1iXZu
U8kiAjzLN+y0tkHv04vlzHwh/HPwhhmTc+nKL4IIYGngIrU+nB9q8QVByIN5Wgb2nRhRNyJ2M7uE
DCpVqFiKu9/oPxOgli7zpMuAPtJ+UjU/h7NWuNpGvEuoRf7wlssFkPbgoth5h5iCvO0zuqLefwR2
tUKU9xGNZDhnZOI4zmIWYeumlRF0OtlKyTISzNI/5rAUEVrpb6hqc2DbQZjWeXdXSXSkEmRu0rP1
1q6KX0/KvOFNSistarCwKHx3ePgeQ2JDwex643XqEJUOLGyZRzgtgrmbVD+RNQuDRFbC98jIxkX6
43lekALph6Kor3Xltt2+3C514+xzHJv844UinXx07aQyuFQX6t1tFnqDin8qOpdB3tC7Xl6dIKCW
v9C+LZz9HDVFVdcxF7xmclnqTweLS5VKweFxE7An2mWhVoCdJv7JsJsrgKOj/pdYarJSph0NnJSS
3sK1yeSzw93iT9jvDkQooVT0A51PXkXsFhTZsHAud7+Z5Ek3CoDtL/H9Irtqq102lPuqT3uubPnH
WoET2BBci4Pod8L/TkorpXFIlsp4/zx9Vg9AImMs06Ni4tS5HZt8JjubQ39l+mZvW6XpF5JG5BWr
5mXpANxaGVUi2aQ34McnmBv6k22gpUXRth3HjDhNyzJ4PnLFANKihZlGhtILq4AJGNUP0+V7LNEU
/5L4EkhQuxY32IZmBGu19FtgIMVkcX9Y4bpSRzzchQqA18ZvXeoffxtxlWPjZZeWhPiFNNfg5VD3
fXmKFXW7W2Nwxx2AAkJK2RGdAVezMIrmWeuJ5j+upWh02yXHitYPvS0YY/omULJ4VEnOXIyDp8+6
RaxNTEbfIyJSJ3rOHd8oLcjt8TDzu/bKKB4Aj7AvehWAt0DJE6hltb329iAOK+Fksq3j8OgTDRAy
qTGqnFTbNwZenjuJIyI0/GVxT6FknVH6eCoMRjBiS1KuckCuhMfHs+gOIXP7dqY5+2ahG4VPglvd
qXn3wlzeXGxwvdmoqH/KOdA+XaqJxy13T8mtROooZtqmOEg/i/8BQV/o2id4GqSCWyJV4P4OV39m
n2vow9LjxGA3+F6yOpLaIbZCTrdxvY/beoduL38KXeheHbt0ZFSPXyGvwNXxjq3ydvCgJJQzXUHC
REoSLTo5Cax7UAVumfO0l0DjZciMgXVnR4DpTjhhbcg5zWyMUYWRzr9FnGSQyh2fTso3xPUbzyYX
cmKDCGsippYTPHYhabKYGU1yuZEL7bvsisA1bRsNDr3o44is/kARVhTGOIHT5AYU1WabxDUEdgGQ
yn90B9waZtB86wTBllx+5NeuNyRswUSEBAE4qGDc/tUcrbaqVcemF9iX+VYJZOzzL+TqK83Xo7Uy
g2uKaTi6ifPjW3TR4kYRRDsgA7v9oJcS/9Os5Z2xfwhR0NLVMuymjj7Y7nHn/ciD786y01ffEYtw
WwL2kSobEfxO+UbZsTJ8bse12ETeT0RZPqb/6yka4OJvN3C/F/Dj58AHFzNUiNBQBXLRx6dqmKI9
VdhFInUmUWJRVzrWgvH8nsXpBucolGmk46PPfZgthIOKhEZnwL9ISg77sD7Fk1PEaF+tpHx08K10
OAhDKU4LTV7oqUZSpY4Ms6+YeLxgHLzdE1U6oTaG6/FOQcDDoXnZdHiU0eJQTom1sdyqAuaVBXnk
86TlO1EzzrvRwcRK8Jpc92ljmQMaG1knsPtmm51JbtOlTEaVftHdSPqEMekJjdKi1vz3t32HfBH3
xfR5PaffJrfPt1H0GRYRA9hLMPpydeP3klVyRrQ4KxPQUNaZ1WDTKi1QiLwmqUrADzhCmDfirKVD
gijYzoE9zW/P7aIE02R00MIVIY8EG+bKgkQMdJtFrxwKtyYSE0MCsjIyzm+MWDJFjMNV/XklE3I0
R7kdyUVyW3jgPchSQtJuxPx254km5eHl4/PpAckZU88TeTK8VSRV9N+nBI7gDFCRIeFQboU9jLKn
Uz3N540JdTGCsCllTvU/SLnNkjiWmQ+IqyiTpTcbqMflG3OpfjX/5Ztvx5QrLeN+uZ6quektW2DW
a2b6Nio063gJS6Z25RUedUo1mHcPrwHg75yp37AS+aYL9rT5T+V0WfWZL5T7DsBEu8cBafPacQYU
3yvmmHJLc5p41nulDNIl0Uf32SnTqjZeaTJjM0rq8upnZ0gFEBtdg53fv1apUj29U6xehiXAsKbe
ocvTT73Gi9OiT6dFWVOYcSYvcu1u0XIZYUIIkr9laYOOYfv5GP9N2oW4xwXSBN8xEYwwNAtm8ZYi
Xs8a4tXEaviwSBd80Ejzirtdjh0xN3HKZthA9SSGjUwFbTWTN0OwDtZXTxX2QdQLs+khzcFgC3n6
yBD6O/uAyLzxzN1F1NA6zuTw2WpAI0Ls6/iSIHsgIr/3aarJqJBylbMLlTga24Fn1Xjubk/YZt+4
rVS3Qv+8A41zfoBebx0mm8IF79Gpm+ciFQ2ZbLCdE1GT8+DLw7fmzmPSDn2St0xhkhrs11CiKhw9
AI8lDoAtBIZch062rwraW/tYbUuI2M9jQ6Pt/CK9j+0Edo8S0BKvanPU2fOsOisanhvld6Jeh2Ak
8c24BvMeU2FJ5ne8XiNHnMbgc0e5RV5DVp7ji6m/w3Y1VBdM/noazInJD0eyzX4IATCD7oEUAFMF
WOVpWD6N/4dMOv5DSeMDjvx4IxAuGwqXf/nolPnMebJoSpmdD1jTKsY80lDP7OE9K8K/tzyvnBE7
DST7XVxkIogkEIsmSPp8n4uCuCUtYz2h1o7t0E6OO7K+BY+Umrrdd2CgTokpaCBO7gUYjJT3GHD3
w3sERvB5UAqbAz0ur1q+YohZjBgIX/DJC8+xNyK4MNRGoDm8arqeAlrv+pUnDfW3G2hSYs90RK1k
H04G2h/kLM7zl0saSTuzxF+GCISKI0wCQG1d7cb6FJKqD+jQ37p51/43PQhij/U8esabSPoQWkJL
Hxs53FKNNH3imzSLkvZeArExfGLwB6c+ZN8b3mWKDaMS3ylRd/MPNB7dSGsOv9vAmEi4jJY1sl3N
VtXOBoRmoP7zq5WAoGBf3EWJ2f/ok7MuoAFtdFuRXaRzWiz5VzFdXTWhUpZ54vR9Bo8XiCxphoNW
ZDaecu3R28otaEtuelBY/irs2CKV8NKr+vOhB3MO21kyrNtqFdsmkwJ6AqhLdvfV2W1hGhD/YfLH
cJxF8fDJ3S6FsH5+1ee6lzIFYlXfvgj84n3XqOW6k1A/CfXF0Sd6mEkeLCbVXIQ06XlzYWJqnEEI
iCBYZ3l8UL+VpP1gpYI0Y6Av1ROdAkVNfWpDW3uOEVmUyWilXqa4UlygSx+yTkUIh9uMlMsIG/6r
rliher/kqyZDGKK+5OJQ1AAfgHP9UIK04jKU3CpyRr91dfQxoUt9Ej7oC1w7TEtOWD/O/xxR1UK0
T319L+bcQbG5rGO2ydUHBPxG4znIdGNc7eG9YGsky6w0DAR6Q2IX3GaysoJsAv7W28f6jNrlMvyb
dKVp9B7y8YWBxO6UZG7WlIhzMAwwn8Y834gc/yZysc7ykHXRtPyjlVBNuNZ7QBEHy7xSWfKeGKT1
Jk2bpQ1NH2NTBDmZ1yiLNuFYD/NR7aM5JoQNN2Xnh5yYdtMl7tnWk7z6UueTAjaqCUOpoXoB7Ncu
vE4kymEhAZzK7fv2VF58ukZPImS9Oe5KUEBsMu/bi12si6OhawQbwSdCyRUhM62jndaV+jFr0Ynf
M/SR65H0ylg4ohoNZD5sYGIYRjUrEjPcb/2XxtoY5GVelXGEP4a+vVBJfEGTtz8FWop8x4cby4u2
o/WBVACmwOwufyC2/CGMLcSQal8wDaM2D59QOhJUw+hGfQRmrUO5fXftVTTBsccosraRNbbE4cVD
k3mljCEkvZYNitdiBSeriCV+cpMzyoXmOqA52PdSme1VUhEm16DDWvn8AxbV3Er/TeiowGeYkoB6
BOucrlYZnA7dn4UpJ4LjHGMC6ZATMtfJzJIkCeyWhM9Ko8euPAjQmZQo3i5DhW6O76Z4looQ2qqe
l4IT22JfmGxKoI+PizcY8rwC/efce9nliizzubLv/H0NX1eAlv7er4DQa/W/Hbzm4jUFxdEVztF6
CbJ4Xc701KPmRjGsBQLbnAqEwfdH1GG/i1JPjLsayCnQDRtXt/MyjFtNIHbHki0/BJEwGTOL0pVg
eDNKyhuWJRWGzD5C5BUVceqWTPsQGv2ybc6r1+Z/ttSlqOSZBfNJtOcWhYSX8KWkOWXrrFjOQrdp
SVgblAIyi5DtQS3J5ZnUMNEOOxXfI31FEkSdnD/Dif32epdyIAndB7doITaHrYFA1Amv3uy/cDf8
eINzFeJ5WrzyTY8r1E4XupBv6HEKpCgYx/6sHt26sKeYlt2mUpVtq0hED2r9WUPLkR1he4LzCaGl
C4vYJde8c5uny10LG3hCVWRwkn6jYywJ4IR2qMP71CrhCydSfc+FSwo/FjJ9gjmpIDMRvIGo0M4K
9cn5gBPVyVDOnlKeJf7d3c4hMTdT3WTRRrAcAiyTjPJU45N0NV8IIMM5+boj+ePf8wk6ViZTQol6
yqhKGUtAOErjmvdQf866xnoSnV4C2diYKeSe5VW4UfwQBFupg22KC8LABcmimZJmiSIfMSnZ+NRb
HdZQm2uo1+jXh+No/nbTBAzBcKKolHOaDAyX4oDhgcN84wjYLd/tTYmpwzmhR/SqQ9+cXNgVD/Fn
3vWmcNFlu9osB+acteYmPtdQsLEkLw5dC+0fpriUUQXpG2MXhPkHA0iv8l0EnoZilSn7j1Y3+Xwc
8JtJuuwtWrXlAQ7J85VWsuUaMeIUfxvbxVrZSPE0p/ItmC9+zJRG+aa1mfENhSWh8Dj54avBXb6M
cLLZJyNLRIzWIq+QYVGxMEgxXP3QjbvXhw0zzlzfHsfCkEoy7pg3ZanV5LAmB92MsaQcl+HSAJr0
rzN6s00wMSaxdrQtSusL1jPFW7dmsnu1qVwnJLy5xGuTzC9WFW5KfPtw3m9iwXi8xqkXm3UWoriG
wqfLxEThkKP2JwG8e4rn9r8ucx8qrfrPkmwxvhQ7u5c9o36tzb+EIVXSW6LS+KSGeNXnr+QC4TF9
9XdJC0X7ir+IvMRfSqi1O2YanHxkd5CEPYy/FvirQK4BHPY6HGfoClhpyqsuXlCEHHooAycsA3lq
sMqKwcR/uk8hQUq9FdHVTgMQsXlOUeuyeivDLoZlMsNm1pGvuxHIYx0wIwPY+Lg9Da+QrMWl79Y0
sl4Vn6vBtJ8ni7tIZG54F81lmO3qtp7CFJEwXCU7uyA/vQUyI++33sMruKnZKUPA66yOhjdRks5H
enDmfdDtG10MoIx8ZVzM9OlX0N7Gv41JuX8xY+xaylGbSWQaGrPYFORYB7fX8Ihcy5GM/dxK29c3
4LmORMNnwruo2qSQ4P2dgNxIunYK3jFQTKOHtz1JWHjouXlJMPMJVSaDdfngFRoTOITQ1T5qq/ff
f5mlfJND1PbKs/gjQtQyAjD9ALonZZ34HoEmIJpQgaZsd1MOXVrQm8Dar9v1l39e2cXOZqgCybDH
RH1P1leKowKTT7N+g+XcXbwjtT425mB+QrWndbBVlwvkS3ZusdICD/qROUrM9ONxAIMwlrSOyldk
qujAuQAb7vn85dS1B0N5mww+r8NyIYDInetF9C4G1cTqNQJ0MlfKfFVYmeU+I0hhRhg0711i7piQ
0WXAr/m9y+2KeLUzW7KWmxlQwIR2mQogWz7BOeqi81UIETUSAJDxXodwDtUNqgBcF/qX6m1OTurI
2gYaeVGLTDIuYwW4zL7POjsxHRYo8zpgAM1XT48Ockx/5OOzyEYwghyBPxNIoazuz3Bi17r1YWB3
oXVfC6LGjzh7VXe+tFrqqHb+mHhkeFyz7ygSCqT8WsYm7fUJIACLo2OOq9JJEOWaFZlBaxMJ6XUi
B1akyJJAwWXK9Ja11T4OVk4F8HgvbhtrcJXO9WEwkfqnvvZT2UA49r41b5wQOG4/YJShA9/HMtR3
sbX3uaxZ0ANo3+LxIoYAssQB4p1TOzPWSr2XtySdR5gtNVTeYfYbV0GHxyj1gyFAblLLNFum6d3R
19ZmhPytw1J1KUgS9nnyzDIWKOcyoldiJVlM8UHGweJTrbM1bRyLglRbgFfjLnE3ShlGjhVKrWo+
cWC9gxGMeyRtjlcSqMHWWFWFxgwut4wRJtYquOcgsjMgAfnFaYhsz6PCr3Ar3Ugy2ZB18NrUBFoM
tFtRmDb9vG28JpIZepz7sslIcKaKgfcMQONf/lS5S8U57+aizUjTA37X/bHJa6M7vqqcjM5JyIhN
yzkZ6LFEQnpMxQLuN4do9YlhU2r/3lTYCP18g47mqwkFupRjgQUHZ6AC67/t18x4ploXsTuSUPag
FFF3DhCahxzbJb+xfvE8ox3nraMYg5m5n/Mg3t5ABu+2y6mc8aUkauFkRBflrtRCQooQ9R23xjUZ
2LzQSAOIpsA2bvLE+c5G6ETHhXiHvY83IEkdiACV+be4F4dbdnLlhdSYDRPGrh3lv2ZInKO86MtL
vBUQcDWVRRAn0LLNSoXV5eRWzocUFbs2qR5X7SvPwa4kqaGMqbJRPF3ZUCBgOvudY+deVbBRHkSK
CKfTOkLnb19CqBdEu3okPzSvyrTCUqf0+AOEj5Gw80WerZtrl49SkZ7EZycOrcfs/J3wkkcamG8T
a4784IT2KtN4WCjaH80tQXWkmKxcoFcZkviOZ7N9UPwKnx5mX5Bxd2KyfxHE4nyZVrMCO5ojNkQR
fXQZMtS0S5EwiqdMvCbvECNzYnfhm4ju1Si171aqHV4vmYa7o9tqMeN4JU1ZdQkJfhz8Cwsv4RSU
EXWmNn+/ELznZzTkHYp/qjL4Ej1pPSAtimD+I2Y72RfksLj5HTXWAkcZv6E0cLeZs8oCc3euAeB+
0xp/lGAgkxcdvAzcycmsMBK/bdHn8FtPNucVMrZ0CqxX1Kp7Faqb+0jRyP6QqybdcEOrs1aHkF0V
ep9XYO4wnOCpX0FoYnzABxUymNdNzkWPnmhCT1Ptus/QbH3lb1xbiv32Y7k0aOZOiD+bUq6Akj9F
lYJFSiiWPo/B7/1qewwFIGP6qncemcgqSQl42UJ6EV6ze0twI3SurjhKfw5cWVM9QGedRJdfcjJ7
JfuwRxfMmh8tAqte5NCh7zdHvtr1+d16GOiynZpLbAO0NpCyTmK/F8r89HDytxw8pesd1hq/5lYq
P/S1flO5126FTkNHo83iv8X9TYrIUpnRBhhk9EpCusxlYPRrssn5c7gqUiagv34zifAp0a2kyuHB
VWj0mkVK3EhIU17yWJ3t0NqjPJeOkQXNFV9c5VgpHC/YZP3jvmtKz3md283l7OoGu/GRtBqb4dhe
WDTDqRAJxYXhK6YN+5JJw/voAeiDbLry8c67sEuaGvVRAdr3/El8SG4MNrRFjOyUfLy646gHAM1+
ZAK0CFFnd/B7PzmJN3I6WgFxHwb2xylTyIu+isRO+L9+SGqHRq5Pl2oz8YUSglCC5HjZ3zJviRgt
IgO1kl6+9BG0wOkMtEd/O9Ui/nRtHr1ZWZ8Ym6goGAZTccNSwJw1n3zwyL/YYmGTeq6y07SOzHeN
O81xAG/JhFTesmLJAms3Ge3vYCiiEeb/5lzWnaVcYo3JY65leMSX4Nn6bUie90JO1SaglUuZ3CPo
f7UsN56t5/lGbF4BvSv0G2EkBfRbR6S6f9G5L64t+joXEADoyLEBO7GjEzYulMUL8zbPu5cPIflL
o8UMBnLmCUsOB82Fg2Io6AabYpQx8L6CjEfVz2djI5+NmRPttMzJ6NvpQfcT7Q9CXIpTGjcsN4bs
+Mi+HnTAVCOIhF2cMgB/VEn6L6ByERSzA9ZchOsJ660qCf+GUWNmSlhcwzyiKQHfq46lMdjUQ48o
GXjjSYm0bo2O03e7uWHYcHvdMx9ulmK5AG7I759qilFTg5t5+h/V95NltPWWrJEVZr8Kw+4QUxby
xrCPwk5vVk5W/LJ5fdStyCZdvTrnGWkVbpPHfOlgrRS4x+1LFFlogOUdcrcQU927syvVoc4Ig2xU
YLuhIKcNO+xY/+F0oZfKjaOgLkWYBJHNP6pYjjpmSKKFyBIOw/9qj/jbDatY8lmmLjQsOUWG2K63
SKJOZqYdicwGJKwcz7io0BpRW+V3LWxNC356sQu8fJTxKRgckdF+no2h5S2MGt7EmhGcWWc7cqiF
Bvdx+wUi5YA+IvWdzx+CWNn/TCYal/eMKfWQltzelojuZ5O9D+LMoA3606mT2BH03QA5ianaCXkg
Z72Os+QMSGd/uYTbWcBizOco1xfXYS38PVQZiw7LPpnkN3IdGETToy19Z13TuZyztqmWuKEFOBHF
J6phhGL/CScigJSePnt0p5fS1Y6B0MKGRXdAeixsbv3J/npjKe/kPKnBUOJQHDGq58JQY5GQRnbE
Bu7ZhuWJWO1nudCGM/zFftyQFxg6crtbPXt/6P2p9tXVR4LYfyr/zD3+WDHLZhwSIx6ygQLzz5mv
MkuzYW4ZNDUMSD7AzrW42L6k+FWQiwe4pBQyt090c6NBI3O2YgosPJXMHOIT0ub+LAt77gOKIUZ5
QxGFCMFg+qfF5MNjfLPoUpyWOD7rPiCI5E+UOG8gAZqSXH9yFMFl1YnKL4oJhLwAMGCx9y29Bkmb
n/z6m6mvHRaRhxkYuo9T0w8IG/RSUXr20DGYCtGtsQ1vVRTzJMiFdpxuQNlQ4U7qGKNuLlDyfx6t
HN8jFJq9lYlQdlk7AF13xLWpbPbWln3JpeyYe6KANu0JSuy+XjRXmCBmpS24B0ATMSQvRX6OoUOV
aGzRslMs6iVmCBrHHNb3hLBsHXravYM1JCMXOp2zxzJEtBaRbHlCiW61GFZj12JXjg+4BotjL6z5
UVGZntUzJRCg5ZfFB3W9fIH+vcik/UuGPj1BUigh4Cc8VtJ6bHjDST7HnnZ2r32xzbUlnpypJ+G4
4ms2mFLJxCNnn1AcYoyi0X9pzfdaKkmY6mB/seFiPKdr0Aw+mVWXnpfKJALYFPIM255RQiyrg29e
LZbmrFqWAbQ1lW6i8ABjhgS8tQAvJGLh1JsgLIatp9rvGCzvUuH5+2PXui/tNtqVPSP6VgSm2RJ3
0Sx14SXc07Oj5oSOtYGJX4aVmbC5TImSG/fe8kCz27nIHRGjdK6r+Snu1WflttscmBGOdWWDmABZ
bwHNIkEgGYRCqpxbFk5MaDKcq52KndH+g9ljU/+QsZ8S8VP2oX8v63gtQPnOIGyfFFQpf1QkF+WH
3XeCbwjCfcWV1P9aOnf+jpVjN/jVqfHFJ/GCpmRsC6jwQgHgjL99B9aLMKgBLxIR3uxKSMnr0f4X
UE3TZI6m7+xtNEUAAPmao3pnZ43J2paeWMyAjImEh9kxQ0fkZGv7Vi2Vs5Ya/C39eCrmab5UfpwN
y7KWZZhns8aGddTBOufMzl9ymHImGHQ9UEPQ9w8hBPlZ3oodjZpsLPc8od5nm/cREq5R1odnju5o
CPMMGedU1aajImZIa0AztvJFZz0U4zvUegwzFCPiLcvaEas7KsPeGw4DYiHnYmPcPjujFgMSH4zR
ULcNZfL9OCPf5kDpVluDy1cTBG/tRqNbcT0Pn/Ph1vuda9PQmHjlRKxum/W+4KsEzQRx9Z68AXII
JSLh21Z946dhf/DF/Gcz89HXPY6qNzGzQ5liBzMyUH/lL8yPWndmnrzVPJhdcliBK578atAS8CN5
GNpg4uVSSvDUDwMbz1KYYw3OLUhQ117lz5E/zwpQK1xO2szMxqDXmTi/zSWSAtl1E3JjEFSwbavl
yBojto1bIeYcG1BobT4Cfd42SZae9xR8gUl0n5wXkusEhtcJBDDLKST9uLRqJGHhgwcl/oudsZ+1
RNwZDTSycZR1s8RMyArsW3lArNgtGla0IV+70hvE9juNzhgYBFAAgBs+5tAXCKSTQOsguCiv2rb/
UDJZl0fK/jqcV0zq6cOJQP90/paGjibAFhQguhH698wLCeq3OPswwaMYQQga7+E6riJrial9oEG8
2hwC0BCIK83h78VwdV5tYn47oFyTUxY6ohriUrsIBF8QwgmXU6y4+hzq7lL8riRnzL3i4UJs6S5z
jPUiJ4B0BpznqC7iiP5UYRbaoBKkZGVQUgnBgNj6JzxQaz9b7ok09AbwHQdowfIKoIeVdb1jaJ/F
WtT3ZQ+lLf1h1Owfj0bLlsKRijMOLwD9Yc16PK5Rl+5+wgSzE7LMIBV4FCWtLNcH/RGvOQmkIDwB
KwZ2GFi9vBvvsdT+v+vua8JnqNY8gHU+8QNTaCd7wmLE0PkZ3FFTutavbAUAFnPWcegPMOA3cJ+z
GAXT59FV35bZItn6UQI8NtSzCu3P6Ki3bAT5kw5ISMyKbrAvOhtmMW1kMuxnlbo+ZLnDplFQMSfp
MNI9O/WehMgOjaP3xAf3cHM/q9rLdQ/twzTkt3/D0VDUXlF/4dM3M8K7yWLjjtcV8CGqoWlJL9NF
US9rS3+lxemWecjlUpAiqRjhmdlJn6ZPY6qYkBxzWCCyeWMe4YfMMgTR25gzfGCpkPo7kNTZgNtN
rm4/IKC8bIWtz8LcjgJ5UQa0qNO4Ww1s+tO1SrkGHW13oPqYvEPGwx0kMtXfkzIOPpxKcfWkzS9n
0Im4NFbc0Hbqr5NYTsZjdDq/jQg6sxc8LDMYCZmXLy28H5T0iEB1N8c7WPvRV/6tfIndCdNu9PKr
rud27nDCcRee9A3v1oYk9UzoKj1GRbj1c6/6mHto2S9EptpZg6wToA3B60F9JeXEdoum8YFMBKVQ
9f19HvaD0BQZdmsBJDWdoFcQDHBQtCSNztJcpCxMiE2P3nxBI3MySml5cO6nS28bQAkxWKQ0/kVA
mLEsO7tUN1CWO6q41ebO8gU7Iv7pPBDX4z3Wfwm62eHAU0KvZWcBYv6945JbUAH0fl+39e01CHqF
qsyw4FAHBhaRvNh0eZSPL6yYkX5Fzz4T1bBOL7CwGVOdoh0uOiQCz7g8nkYNjPKlzdDF2A1ugXhn
lxaIjSLyJTC24clNKN0mOJJy75oSe2MKfDeLFTLEij/54ciP2AX2uBI5tGGV3ZXM+6sQhDUzjjir
UBOZlfVQm4x8mdVnszGyfwcP2bYEl1v00d4ckMUipzaP/DxDMK66jqfXZDbi7NhpA0tnoNHOI6vB
SXjoYxB9HcAbyThrgp0J2IRD0zd3JNHY1NgGLMkxMB8ACg7suJxc05G0/3wvr2t8tBeYO7zQW0sp
FbdKyEuHDqN+RSUeKfieR4morv9cBNN7vgF0AJu9ZpChDEJMsCYaQU4+HSHU6/kKg7jzLOhYuOyo
NOuIBnk530OK/jVsAT8LI/IQU9hnPJSV2fYTsR4sqWrKLl21T3x2DSWU1S4bV8aupDue7sNmE0bG
G7tKq/MdiazeKbIwnBQ/wyBZjvMx/r3qxZpay0uR9okaA3mhNLym8ZdA9jeGKd3tFUUlzSkAIz25
y+hLnpzZ1S1jIafY4n1rYtYr+UoowaOhWE7eRDKs8OFPGpNpJ3rc/dRnUkMwfptxzFPxi5/RtoA7
eo3o2kGZfnsqQCos/urgP0uVFZRvKnTLXIfEWsdhsFpHCUDisbmFy87RDioHXNfmWaxeTnxpZ2FH
NLLyIu1X+zGzRyvhABxmXjLQxVgIIxF884/VkJ9p82VbYed/h2vi4EoM+lZ1U/58XSy67Eyukd8N
QcMMNSf+I4HMd/h1eiBpAfbgOhngILzi9Zi02tGqk39V+vUlmDMw2vjDZ1wtKzrjAz0ewSJw1Ui6
XFVvcs+ZoD3osctWXYa+WQ/YUbWCVB/ypzMjob0Qhl6BcbXZbVmZG6tzRRwbMwEjf+JEVH3BTh9M
BslX5SX6mqeUz+wrsgTlOXTI0iS+2M3+nnRWfXdhtKqwN+6mtF18Lxmjr7xVm2jbABEwcjCVqsOG
k2Rcpg9eICg8aT3Zz+JiQHKaBihklKOMCk59GZ2ch8DMOX4j68EZGgUoR6ef0N6ircTFbR20Qa0q
RsiSZffQnOFpln4t932imZ2eg5qSRFrFBSSUtVingrzHvbKf5XP0ElYdNoxbNY9nFb7sLfqfpaYa
oUIp9F/P7m2C9Z/nguJeuozp/eVBIp1XAN8VRlWDkntpWsYdokKUhXUtY4Gc7sKebD4H4eRCZ6WS
j3ynNoLQl0/25nih+WXzaI6M6Lc8AOSRtTD44c4zy+XHkLVvUjJs3QVLRyeh4vMaFVlXKDDRLyZd
nu4L2IgHuomRFHDqY5wZ8wuEXiGbWkq9vJFc+54GCRBbLoc8J3/PkDMUKSjnkUvcmJ+FeR+oLUCX
63TvML0i1JMq9QOKkCn4h9UcHcCuDmp2Fuf2OjHbMo9+Z5PUi0O6JJEUvF5IRCgcPqN/MuTUAVbn
h7td2PNUQMDnSfhIJndzxMB8dMwCybwfzhgGGgn25Ul5VTN7C2euSDdWw9cf30yrZmNXMpJRmH55
LrLGJ9x3MWkGlYJkEmwAQilVJsjlNwlAJbMPHyt4sNHbsuFRf37nDuSSgh1+WdFsvFyYEoKTm53k
Cez5C2nq8QIBvL7nEhqVclSrhPAJmVoR8uzQ5rBRETGV72p0Moi+NNsmrBB/D06rFzp9GGmoIevi
4N5NbT19p44kQjszy0pk6muB/8S3UKgw3Q/y8b5G2j8YXFL/erGkri1jMM7RA3NYxnoETUdD/iV8
BIQa9WdqNZoeAko+LWzD3mJiJbQAR6mmri9GuhE5m3OG8PC1EtzDHO6C2ClF6lUU23P0kNPeSjGT
LNkMpJWWOP2EpQhzdpCEqhbyyxeqqnBiFkVKCqTZH4U1NKXzYnqXKV26Oqv4c+Kn66wulniar2wx
HV1bnXip0z034drrwSD/7ECkSPr/Yzzfznrdnvce48LbogE7qggy2JD9FnyLHRDNy9qiZc0XLYYH
sfyb+jmhitgYwKh8jvHl+LUV3Ie2ed0f0nZXS9Iwu5JOZfKIx5jF4epCSnspYVa4I9UbyGcIAIqU
L6mCmX7sv/cleJv4xyL/6cfD9371F4SYCBvUQSS3cbfKWG5p9XxNjTEMrwlkticEistyreKzGaEe
a0VWtOtHZi6+tmpngX5FniA82+N3izkJqajZL2lH2wvzsoeyy2nuuhuVcpk9UrL+cNwqgHqgqg4b
BXJVZEjJG63fy8mio7hG7A67ffhIT4Gdcl7m0mbdfm3jfnLm6EbNAyid6dIUgGmYsdMYiLhOlEVE
5ud+ePN9viRTcN9X7VFWKp2XAxtlSPr44gR6qAU6IHUhB6I3OqHmJHBTZz+HFaMiJ3tkJh2c7UkV
BQrOp/Ab/jxzs4qYZUPAtFtmpNugz32TW+8Gp69JkLKH2mwscB3UhduFeCAsdVOzoVP31hWbVdzn
cD9GaK8KWSm6ozLJRWHZOnrGWHdbqs+nsyO4H1lrhoHtEly34H0n4beKjJWgs5EI+GqqZ/DgsSgy
d45FUNOlnLW1Szumm6tY1cLbb+SM7VLWVx6RtbvzMZ0Akt5C9VMvbPh6Nh+A+856n9oU40zEbBGg
X4kY3WAWWTDM+hnEZWLHsSxM0XW6Kvt8ffHzO3pbIA8EwO1nrfaDGf9J1XMj2k/YRkhzxVZXzoYh
WFtTm/4plp2pn9chLRgPab9k8ELfOpAQko8V4WaQv5fTOUckqX+y4kqnjZJrZeLpK2N3+nOZGrbh
F/SLVtddBevDaQeRKXxh6vuDbJjreKG8RdISQUzobc1/N1Qjr35ITX785I3LMSd03vva6fE5VveK
tQC44LOHafH7aYZI/gOhMsJW+gLOZsO4YFMNjmuwJT1zx6EUq1D/L0nDkzv/1ysq+FQRiFd+Vr06
aUFuYFID4WARrjrqYFY/jxff8zV5iz9xq1iIfJmZuSu4KYbFO4fribD0MAlXcCjkIsRhxONL/7iW
Gi7fHraRQvofE9J54NxlSV/hNEFC5hbFmOBYuj57adpz2erVRzdmBWERXSPe3gE2qwULgdDohevr
oLCENpmGLtRh5k+EyTXoc59f2i9sHRaquE7cIHNGAAs6hqqcGwcRNyF35/o+/eKZ7CLujMOat2eV
3V3t8hU8ntKrrGyHMwaS8BaBt1JkVcaUoalKGZ95IQH0JXuod8OXOsZVRenkgmpVnuU6FE4K4oZK
RG1i4ztBuYpH0QkxIBYWF4XarPvcrdxXEQ3pzE/5tY6kxt2RLpa7+Vi6ye64eeMa7Hwifu+ebwgP
I4ot2k37lC8t1gnOW56Ic60rQ54Vk49S46Nq3/mDkSf2nNVNVAFMTGGkVXdF3Sh7PkZ23wnHAaaM
c9Zy6rQZa/xe/Zb0CtWwd/BxcWMYmK2McQD4Oz6jwf7EeJJHTMbeCa+yhmHQx1Y6/MY3MLSafxnl
/ji9Z5+jSb6+aG2vSUi/RgxSg0RTlU2Iy9ALIt88GnwiQWQQCk4ZD2P1cCaHnlGEuAp3Ea9MiQX8
TSUW/D6k2+5Nva/XBhDl7cqlC4kRK9jnGis4myUo5Ux+UcuVUo7xCw5f4oFrnf2yObqCJaCC60iW
HIIbHuyzRXPKS+F51VvWeT6g87DbfAjz298ktN7xdEX7lyX26GtAiSAdpUk7WA5hJuxRWi6FKzRk
LflBjLJSUO8rRk+ARs49/Str6uh3vrniP+Httgr3JORs353BkZEeltTQkC5mpNopQ4GI2HVDQvim
GmFEzayYvhWUm5gzpYaPCnU0Yl3ZTuQfUja8IwyAqTqpf8BFBZvNRYWm/RsQkrzrCNL61x3bMYLu
E8ojgyygFB/k319KMQPM8HrkTbAlFJOymHsP2wnFRVTuBpuWeq3QvRGd8PXyT3bN4j/RiwCeT8LL
HMnQvuE9T7dBhK4EDop2HILmXs2wNq8UehxL3Edo/BsXSsQpg0pFvLr5IaAlkPKm5HaCf4LmqUM7
BoDUiMhCTeKcfJx5xwIDfXk8IST/NuYKpUDp87bnHE5+uYYj5frq1rwriTz0ytqkcOTX9lK21DvC
JCAYVZUH0p+NjN5pospaQ+y3A91KjTbsw4rBWaZwFR2JwdR69BmPruowGr3usRjd2oDaZVGFjEt/
APsKh+iE5GHV1uCKc+MiogF8LrpRyqW26fruFKMmknpmnQMlxxECqr+pvNG5202AMEKNjd9jl6gL
eek21gkIojoCPRQMv2pn6NvpKCFT5ywZkfcUZmiJXnADBZWNhkxv8o8w42zkz9vVdY1JZFEyPS84
qkvGLEOKMU2oiZkW6RZdRURz3YYrlireokSyHEoDK6tBwqbKKNddLiVh4JOEzL5fVBURYFg+Ei/f
acvvEdV9F3bBrcFJwQ5TzzmzPdpbizL07eWt20XtcHNVWWhz4hoshze3L4K8KoQbMb0IOQyCxyLl
nrYM1srBzzv2wwNd447wGSrUBs1uUNjQowS3507UKe+i0nC6bx8rx/bUwGhCj2JHw9Wymn2MWHSx
v8oc1XTHo52KXhhXYLWPd4KuY0zs3oShS+AWB1G4CqDpdwLovFOPNSlU7nKVDJWMx00XJHIbrKyp
2ykDVnmhCfRSZyw1yrd4N38tKBVGd4GSac83HvC/ss0dDpA1XcmtyKUJqtnNQtuKU83mMwir6g1O
a4WWU4KlwtwAIgEBYna+Ba/nytuZ3AHa6HimTQeBBLmOgXjtUrb/ErK6rHj2eP/27cE3LTwdV5Ai
zc3XjnqTs6E87l4qLPxPPT6i1bN8Z9weYAC7BpUpckTHF51LI5qyXU5/2XJVio8Ppd+48LLg7xh+
jbCff4eB4YgN6JH1yNFzpkv94MPioyCK+9rQTu+Kd0lR/5VMXioms58ce7CnvBBaRkuIEETM3UP6
A53o4VMmhpjo3XDXVU2N/lCMTHpfaQ3Mi6+pQfp3+0FachHukdodZXWujnHnv2hKFJhQAUkTIUyg
gr/9dIJE6Chz63DXFdbWVZZq5RL3jgrFq5+XbFLEBPBDqAsHosnE1T364JdZwHfVvSZXLJpx/fc7
wLQZUSN/cGjLNJOZJI3hJKPiP8uRI7DHfuSpIOLl0ncXr6cZCTM+NY5gjz0thN+qZzPwgu2srxHE
zRzjJpEQ7DmHeHgia9OYmHG34zLUmFCC2wPbpHQ6QE3iV5j/6vsUgWLdZMAcvHFiGzXRuCsnljLu
LYgo4TbdX9ModDULght0jQnbX4IN0+X6EWtaW+uRfwziIqEJ69DQlecJN0Go4m4fCKhcFtWoSlo/
ldDzdNlu1WLcStFcf9b4Wb+lA/3TG9av9rxYhDpJBIJsDI+0IiOsmKdF2k6oxGfCx8XvSwKzCXu+
9+uRfKjlK+1kD7U6WiDjNFQmsZ4dVaA62nU6DEr1NM/O1+AY+NEyr7O9H776ppmrsd2C5NgKC6ox
AP8QI4vrKi4QSz1N7/QwzQZuxSXOSQwHWg71t4wko4yK//86dftEBJm2kYojCOcykkVedxGsN2/R
vPH0mi7tLj2WCnCMzjOAQylTNd0a0B+0NFeg/rMUOv6105Kh1+ywZwZXwjWxbtJlmgOXV6eSkpXq
EkNv/VzAER/NsR4qmd9Y9Q2O2aRSMaLY/YO5zpPVAanXQ+AP5XcDAb0BC5JMTuu7lxTpFvYz0bkc
1B35bjJxfz4KNwDks8svwvAvvrzp8GX9dw5VMYqQTAxe1DZpiad5rq/3QZOcSE/scbUTRiCI3MT3
EJ0XbtZVL6P7rrKuzy9yupBCsL2SppsThoedQ1Ir1GaH3rpSrphBN8G3I2jNlGjszE9etkxk845A
CzHBhkQwSyOSobvbpeFwNmB1X7wvRh/nVfvClkCKaYW1Adpa9FD94gBLeGut6UTLNz5sj5aNSBFC
jQeFFsUs3Gp4895B7QMDtTTSTk1nYNC01CNekB7+S9KpHfaVOXdoxmtuV6QO3rEZeOcwWRo5vIv2
I5tQmaQKnIcCJxD7BkkavnWgw6jtnimAAYBgjmYXJYOiubptGf3yomjCKLav4kHpSpwi/4gu9C6a
hRz3gtms5aSO4KStIY0/ev4LHyr3bkRa1EyRgKh9CMjfOHaFE/bs4umXwrF8U3YBTIp1hEjjiQoH
KeMnWBSQMA4/5j0zvmAv91IB0n9Hjz11LPtQCMI36Gjxmgj00uUuUK9pGjVfO3BFnwp7y0iqn4s9
aCpjJ2is1+/XV+KN+3o6eE/K9fmAzSfKOTUAsM3ErA1pTIoT+PWoF5JesdKXWyT9WtLHL8Zc66XJ
YM6c/ic1SnoXU7IjFd0xihLgcGCkLpz6SgYtQrTxL66R4wZZtrskrqXXluTjA/R24yKueBRlPArN
4/WdNIr4n02Cz+0v/k4ZVg5y+WT4rvkCwTNa3ln4KPlG/kkOp3lV2szc5MRmOFCjcD16gw+EIrMb
W1GfD4q7Z0sWTN+tEUzOSh1U2PovhF6cKURHyC15qv48rsIOhJne85TqV7mEBxh9dzH5awXgtPVY
NQfWG5vhoa3/r7oPY57RG37CAKLkldzqXnMI072i3depyvgvNQKQrhC5kIADGJw+94WLxic7Sr4w
HpeMzsMQlRH3+KLJtvrig2Md3Dtmw/x0rvyzyn8ikVM+groa2b5G6GIxgT+Z/p1QpGB4/NXleXxR
j7CIMeCapVxjlsXwIZyp8KuWvZY7M4ecgmyCW7Lg0WNBDarkiTxTyUfyuIG29EJqKJOsjfEDMmA1
G5smVlIu3/iYqnK4Q+5RkaMljfzaB6jy6jk93oABWm5oSwKMY4ava3EcWKofxfztcMNpqfD9T72V
h9yTuAe9v0yC23D7wh2R5q2syrEgrkL+DzrTTfuXai+k1+7QBez/rAeK9xNwJ+RF/jGpKxUTFZgA
tZoat6xHV00c+cNlb6gQSPGRFdWV4Ap4GYZwCahZaaCgsAndIsA0TMVOOnAdwz7jcFQ92c/8odM9
T07zIX5+D6Gj/TBUJqtYX2c3zokeDZttSij3HMhJC4pUgnHBeMArHyQUcirpfKLXP+Ny/yrruH9A
wOwmBwRbGMmlYGKZ2Ee0bdbUuq2Vzas5L/9DHh6sL+WvCW+ifg7i71Och0Hsslad/3lAaynK9FZx
WRBc5r/0My2bRCgicSP8g78IT4bzK9nKprMY3MBH2qJA1m9X34t7+Nb+vSHLtD3yfsgWZrBaK6rx
e01fK0vQW1ftpLxOstJJj4UofObGboK02ed5fi4bWLFY9NBqgOmiv1NRgkw5JYvJMh5khxpXr4fI
JEmtIpGYsmRVgBAuiOV8/QH7FTHd1fagg9UV33LtKdq0NSLG/Pwgga7faDqOtBY+9NBsdRr5o3X7
X/R0WFeiacli0WkulBd9qsh62SaC52nhC2ZztYXp1rk5dHuJ72LRDf0cZ9IQU2snHFxTXmE42P0A
WoDj3vmf80WancRPO4tobldOvqGPitrU1a4hs/yIBilc3FOZ4i8+Lk31qF4LGp24hJ8wBRX1AHKx
XIXVhbMIHJGaOsgNDEIb5HjHLOJHUIq8qsF7S/IKaU0DuIrkV449vrHxdT+sv/PQ0U3t6sJ0/VDk
yg/ZTUvpFXOHOkDCLqhqiRcwJRd0c8IeaRlSwxr7hL9NAMmxeB07ECkNH7xITd+a2DwsDEULc7jR
MMIDGxqDE0jVSqt1uufqFlFjvl1ZT2j7XxUvAmJzudfZLKhclwBIXMbdQ0x+Ost9pHrPn03KI2eo
+p1tVfTd8AzTEE9jw9wN3P3RxJLmILYDRk3oez26W6cewD7EO+T6k/zOPHS/cH8QAqn7/XFNA8K5
1FezTzAEXj/LZ3W2iKZwaTYaX2d+vLqqJTOvlYjBmL9QOxbMMj65flAn/bt31XtQK+badCPOiCPv
S6RvWSClx0oUzsyTBhf/UM6C7dRVhdPqUU59++GKx0rgZRD5Xdv8jPjcrd66KDIZjkuJc3oGYKgt
Tf9VItF/7JYOpo22K6lJW0MRtxVpcl4Iz2/dQF13tnemer6IhEHrKKN/RI9y9FrG/CMy43TFTz1h
nhGEj5YAz2HPPSgLoOa94AHffuWoWq7oG9qx7MD1p5o6c2fTpm2URt/Dd/kF5CJQLQXz9JGL2ObU
QMRUQJ9HfQhpm6QerZeudsQGUiWN9bnJD09rwUjR5vkD5WQFnVuSCzAMn+LGKuX2Ic/HIprGzhUJ
busKN2xyI0Uo0rwKxd8MnIvXSs/R9u5o5OkTXhgfN7TMXKJgin9R0y6EvwNZNbAoPh6rk0E3N8OG
Bkhng9ARyOQS3VBNkOGyh8Pa/a2GhBuLYo9gfG0Fo4OeeYDMyzl/kjWxWRu8p5cJCyoEtB/37+EG
ZU6AsdVfjh2llnpHcOdN/dztP0qLB8Yr7dPXl3DNUpqjo1+HXvrHNw1EV2Sby0LrfS5i1gS/P8h6
d1uZBrYs4J5j3Jb0mXpII7QieOJY/zj0AtQkEIpNfdOjSA/Oi2qhX/QAatlikUHjSi5wm5Odhzm7
0aR1ifCW5qKQZ4e3MP981ndR35anKnI006iqyvDEPqmgfg9+YdxLSxzJ0nYQAUC5yrcZRXY/KGEk
Ld4T4NenQFeb4LWiaikL+pyBsEqIF79GJAbW5ujQJSO8O7Dr2s392lEjt8LgLP3EIN9j3RzN8Rul
CwvyZTHkB8Yb3QvzWhVy2w24/MxJYf7q8VXOKEZaiM0YabCaOG/Ps4Qt1tVIv8amQhZE2GWDFjtO
YqWDkqSlZu4ce6Sl4QBBNyXbyHVqYBVpCjnxD/lebBM0QMWrcO1/+zaQVwIgKqFVDUEKPu5BDS2W
btoJqcBA1S+X4x3SesCelPMEvTq0FH0zbMOBPb9MQufLU/zvcUBrPqxCJVsxJLKuwE/4jloC/27T
p5TOoH2/nm+F6ayISW5l+aIa9104gA/vKdV85mTjAFPRrXPEWsbv2BKDCwAs8Z0ySBbectdfpqQf
lzKvrDAjsnpJnuCu3G+f7JTlsEA0Rnbm/IG5jWhHFPGvjmwr0ToykTqmi/Rpuq0xw9qV/WaFMRUT
Z3LpTF0tgjwvMao5Jf15CUVavg7sVyKIFfTZ37jlrydlXZBHomOW6qzV3Zbih0GLCi2O0oTu19Kb
9vt84wvs0bJDwB1X1q/+fF0RKw/NSIjXXTcK/j7z4O2RKLx5cESRR8pT79NQFPYRTJ8adNChz3gv
FQApu8f9un1tgFb+gyZMgUthvWHIWPLI6gS4knxy/W4VKFkHkyhSI6cssT+a9fzz8CKphNnWYMoJ
EJTmf/boFfcJNZZaV5DyXnEb2JTyGYQn61QdZk8i3zXFk1S6/EDSvSHHuYiNHrvzxYt8fOVEy+lG
MBpxGJHTeGMvIvlsHYPGWMf+AEqWiBJFflUEc2PztMy2AAMGHEUR41dheufUVQYy9+0JCOmhIFKZ
4CK0+9/vmu6tAdRLoVP3yVEiilnm30BZigvldJrQetrM1A+MnU/rXcGOMYVsz5Y4v/PCz6bpvPuR
+NFBP1hZkZmwvOuTf/YFlgshbwHS1iG8ZnNw2taxynkwy9h09fYiwX7BUlLeDZN88Dqg15bQcqIP
zmSarnOSuIhSzz6VxvOfkM5Fgepe2/weRP/79fLId0+zzmnpUdJ26Ha5lib5elZ9GGWYUcvhc2+I
xp1LOeYpqWL6Lea4IEvFnG0qRMYH1p25cTOOP/5UYmF9XLhCw3X6pFIP/DOPDNcnqGzVBUYEseX+
a3y0uMrAgqIoE12xFreAbcbF4c/nrn5G1m890gRh4hHHf2RrTavZN5injRn5obxDHZuE+V5DUUok
02DYdGijVihckC/qVdUoGrherlCjY5TWABylZe77pD49pYo804UkBMD0iS6ouHBR794mejp1fVQ9
3aQruzMw3/Gm03Mt/CPJycIAyCGrtQostaE6ANHyhSB+KgFzUoK4fB10GdsqM7PgYes8wKzMYnOi
NryAFQ2e0oKdKfxpiulES9WQwKYt/oFiuSLM8xQ26AolOXPYHv2q6wH9xWCUwj4R/sm7zYBU0Ig2
l2MJMJc0qQjSASdmW0mjI6RxyQbUVRWZe4HFBMAshtbHdYVkoa9gRzybIDp/lwIz3ZPX/u8P7M4L
eiT4jFifGdU3x88vb3ba08687DpKCuPKUYl5rL2LHuPH+dVoHZa6uamp9i88g8DDAJcon0vdXAbZ
H58CmolMd5HQvKdiZYTHRwU/4ay/kI+BYDjg9o2bjFzbg2P45e8IyOUOrjd+7C/OYa/91cHZvNWX
CBj7GlCwGvJ/F/rIQtFG1QXUDGDDa1R+pu0itw2MHoejEycexHal27DltwHrGCkMzJ+darcXVXVL
OYOFki4uUPhPT/hcRCzWi3PPu8a8JcrPLm6KnsbSYLoFzhYa7SaG6amYBDzmX5TwzGw4p4JL1V9u
NHpQapYufW3mhZRIjZ74UEaUNZoqBpmCu0zA5Nw72/3zbly9grTY/nYwtfBavENwxXpidSpynixk
dNEVsonfFAcZEBFKTIsPIRMJStyNjCuNhPi/aITlqYPB++KYa6v8uHUQl0kYpaz6UPqXOaPNW+Od
jvKW8lStz4UKplHn3igI2Uu+hI2TXyQq23fibNWRt4pUVwW7aK0fqRHwVmw0vcnZcMydp6orbnPa
eIyPiVnxhfDkn7wzL1IFE8Jy+piNyeMraW0Yc0grVlrvV0h3aBqOC2f0BOOW0PAlD0MSejGbEKy3
20Z+vtL/g2kywfUuuxQqqaS2lPYwHYE+TqWntjldc+BJsBpxN+tDKLcuPPNLsy5DbwZbaqfPoBi2
4E2I4xCHG2Q17smJNz3SnH/GfKplpVlytcTOSLWk1SZBfFRIcMD6ojPXgem2yR2pYlt3gAVyXr3s
Ied7nG6aV3nZmqliIiEugSSlecyDyhB8FRn3HYmj+jNX/HrfDNE126ce75HXW1pA+6YbL2C5mCVa
OZjyCXQIb5L0rZzCaxfMkl59jsTl5QamMQuIlpAmQyO1cRoWImTVLHynZnnpcEgexv/cbr8F+t17
9i2y4N4omq4sYjNUvmXLGfCrThbvJ83JmirdjWtfnISHryz9DFOLIKHyo7nVgSxXbzqVqUT4mKAp
Fm7CL53rDoBhIznAj0JxYGhcL8Rdnu2rZB5Da0iTJ9G04ViBebgn5XQLWYXlEZqCp8ik9boADohO
hb+hgaVgHTIzn0si94mhGaBtHrx7MALWMjCT3O9iFeVrSA2EKWYggU4AI4o6IQBvTml3YUZwzSRm
P8U7MduilNZOauomF+9+vaBa9DFUfeHNwhwpkmCHpihQXlP9oAAuONfBJfzd3QxnrgEvropCYx3f
P+0AvojdJ3sroChQbFycwq/d0UWOelEOV7Yc8BIJ4JKZmJuF6IGhCTRQKKsi3aHfiqM9mgtykFLv
t3BlObHPMJ1Mlu2JWSkW9TVaIqkABpG3gIZRrE7F/2HW8E3rTR+WDEC2eGtYwK5F0nQr3yRS7gQR
xmBjjPVdDpTCxpphz6m7QsFgEyX/yosW9eM5yTX1DGiGIrFMUiHoNGuYUEghrVUVG6BwLujKL0cs
is6zEtB4HHi7/YmRI/f8burnITP8Q6HcviO8RLugaWpEqwil4q/xW6yaW6DR0Y32dhJ0povuMXAQ
xqYRsbLll5Dj140bfu7VwtaYgOrcnQnxZiybhshGx7dhg575PpcWn9tXM5pQZ1QwFT9+cjy6HhXx
C1v7W5lB+7tknqdsnUlfB1B8yBu9x1WXVVAK0VK9nmVXbqzTxfBaQ+FJnWOfUeNAQe/axfYfzHq9
ad/dQhXlYC7cq52OuSD1sauNgXqKhYdFOCGIa12PmfYpRBNZFo7U7OM2omW3LF4/etd1+B6DFxT9
nw4IGAjht8vQvLwVw00M5YS8naErako6IugjQaD+LfxoQcIh5yL3Q3sSu7auDI2FN7Q9ouXhNnDw
ovN6WeCs15ZCz5CT5lbFXTFWo1cWPHOOKzFoVwe6CEzZgUijFe5jX8vo3Q4azUyPDOQKkhhuncRq
AL+UTQqlLKNSjFj5HIaDOnf9uTDOEWPDCAM5VqL2qDdO7kr9FDTdUviqjqDPwSLR75KpmjMaQvf/
SqKXqpHWSV5n9qKhlA4Z9Wp+BVK9KDNcLLaVFK9aPD68G/jnYt9vYJmRkf2qmC2LUhvf+ypGMnXs
Lp/Lh9XLiTUsg74get/PxRY8yQ0CXlKG2r/2IESTSL5iByLtm3xU73t484YgwlAFoo42JKFFeijG
ojAGXb7pNL+dBAcj98C25ozJgrMmNKEx+v363PuqI7b3AdqehtnFb/wvxp3QnCrSS0VVnD24/d9M
bdcbB7Lb2vQJqYNOgh572dHksSl+X+EYa+etBmHjaOB8g6UT3bQylWu8bIlgnP36g6wR3TDlJneS
620dqi2+5WtHB+ahERMWWYlA5YdKygxnY1g4qePOtTSeIxgTC1ieQtbOYf36VE+E1dZGAuCp1ruZ
RJP78QyPxOkMz8Bpq6yFKtbdQNzJq7Z6ewVPSZuS1o8eEgVbEGiaLKsDP4EM65Dx6pUvD3c+AZXQ
DBgcIIdqXEP5mQm2T54/e4Qe1QfebhpeVR05ACXwvrc/Rb/ohmwjLBYdaEJhT6eU2ZGrB5xnJ4hb
+N5yTPaJK1DYXo0LeRxu1WSMnxMez063kiIfv287iLJseXaD2Z1+O4fYcqwmRRZ1bmnUC+mIPRaz
AqSV1yM6yPX+T1LRIy2RYNpwU4pj3JtAPUAx9a8JJaS8irkWJ2PUVYF/0B8IhEzyLht4vcr//3Y0
3PbmeNpsnrxekU8QEqW0Q5z+tCtlSe0l1tIsw4yoxOUU5UxMdlMRuParP8BeqsN9QbHX+XNUINzY
yMFEIoys4OQSp60OKRyTxQRhirXPeMYWrzM926wzG55EENw0GccI7tw0ZuD/fFTY3no4h2lwn+Cz
/hkuufqqIxBS4tgYBSuFLBxKJ3t1k0j/NPFRKtXwioguZ8YdtLIEnoJ7IX4fq3W8mJkD1hVwW2nz
IxrF/7W/KuGRfD0QjKEMTEsjtabCiiWyZxdgOLtPnFpJJ1o9ng7p3SCpQOwY/a7zaBaea3755mVI
zun5+LOXQiki1MTSsW5QCP+zBRLnhpOWp5rkxDs2rdgiejf4y9Lwuf78QQXqbyGABEGaA69nc9MZ
CDd874WMkQQ2NUAri2RTkeWdf3SEt9+mL5lVCuL3QMYonzkENxeG1v0QAW3i9quvixoIZMIejYbc
81nEOp9aWQNBibuNfDkYiYnUxchFhdvYNmuLdyiDOeOABK1VR903U6ka5PkyKMySWpZZOQv7j073
WHOaYZMRPlhZJZJ87m4bIxJHzZWk1gyNOegeBi6oP1YVnOJXoA02ZIonFKnBdzE10Rv9k2vz2N8p
Ps15eDtweyVTUshhuGuCXdseLs8hQH18AicV7ZvjPUyBaWnIPa/ugNwxInxpViGkknGXaGW9z539
aAMTg8vQ990RcO7/gahVTODa2AInsWujgx0hpLAY/346GnegQy3YUtqy1o5yFHRx5UeWns7SHDhl
AE+9SORUSo5LQOz2KZ01w+IjDERA3CFcfgsQaaaVD00boTb86hf9eYwT+3Au2qmQhhMhvuJVaCl1
i9NKAimkkDXy78e83EjtAQB9ftfCAANfp/K9iVOPajOhU3E3/STMpy5jS4honPf7VPCU3PPNLnpZ
xxtTZXlhqQ/xsO+h88yTNhM7KMHZNuqXySkRimL/AeuRYXajR3O3++W48SEA/jz3f+BGq8gj4vVn
6BkdsgrWB4F8F3kqRhyffXbsPdCrmrmZrxzORgVa9bcfbcmikYq11tAqDzsmcsgwd/w0wpA7muTj
6qHh0oJDiYXnM4AqpHFDfXMZ5JU3pIZjpJrsrl81Uu3kj5pDnA8swnkAi5JLkLTRG/Wk0D2WE2co
MNLiz56/qbVZltX+Eyxyf4H/1tDnTW6WCY19+FKZpsntz1ct+Rj9v/83V88aNR/bO/FNYmKgb43k
L7vExGvJUj/eGZo90kIBCvGjeCmfbWLjOLkyJc2oFZkHKG+LtL1fM9dDOv4S5Nu6rKwQILwLlLtE
WC+OFQzjTUdiC/CdaBB364z093MtprVXr0P7oaJ/J6GRyO9qCjd3mAjDgrDAn1YNNBPNi1vMEPy+
FskDDh25bWUOrkgCOaIvNIEtg4U2ZqLdDeWg1G1Sl3mnKyoCQua+nVJVN4S5HR7ns9MAU2zXQ0yN
sxhHuMHX8cyBVLpg3rCJ8kQzjNqi0gUdEDqPt0mFI+IdE68k75NPYCd3DOmtfcSgUIwGg79aboSN
i930gtKFIM8O9WrKNXwsGmYtM5UiAj4u6NNPGc+H1jU6O3QREYDNP559XhkoJaJx6hb8dNxe80+H
BBK4XbxvXPrUKMVGjCK9pQMO0Mt21QIxvaDBcAVNaZNjn/3TlF2BzgSex6WMkAsxBzpXqeddQbT8
V+5JZxe98uzF/kJEitmXv+8BtfOauH0H8ANiSpy5FrP39ZELm/CfHdkRBvNOz64wS5X+oi22241G
5zgUjH7sk/QNtjmQSj9A7PBDMgMhNL+VijM1WJnWg18bcUCQVpShIz7Er1/CBpjwXITvbQ4EAXEa
XyrBLB70fq3/qkPS90E79JRaH8ekgWBe8BaG9TBemsI7NtWU5qyKLnRGMqIJjUw8D4Q2nq/2YV6/
vMb/+vHe8RV8vH5mwr9COjvAaUETJheGVFhT2tAIlV/t7P2q7M2m0wHf3LT8erdf+0ccGn+i61TO
QLSxTGGAYT88saVOWi95avkjRp6D5d4jaxTVutrm2/ufxaI5m3MfhBuxgHO6zjsZTQH4Fw07DgrH
M++hosjkqCh59bzZDQR7xCWz+NbQnVxt8lpOddbkb0zMemZJLjR/LlMsy21e51p36oOz29INbpXO
QjEE5J7QfzHneZzUVwQYqRxubNpmsz223VgNDx1+d0rAtQ/F7wl/s0IPLe9tuOw1RkbfFAlV+A+G
hkDJ/PpD6iWHVLnfhwooTaNuTe1DvgicDS8T7e8UWfHvgm65WxZv0IeqgSmLhZRujEva4+PpOczi
kminsqOR/acoDlZ4pCe8Aw1jzXX2zsNrX9XoGntb93ylCGfMMIMoiFQ6q5eeMjKtuoaXpJynV/P2
uJee+3S+zHcCJGmYla4M4q7SXzMoa/Bh0EJP6PeV320D+sXMfJNiE1UCHx43ixFT9QsMStVyYMbq
FbF7nU9I3TPJ60gbYPQXjSwHP46vz4+FZEzIt3RwcJqQJi27QdTH7JVrLxvLitvjMWBOueTC7vgJ
fsBc0JvU9OxUiFMFLe/2nui75z2ftIMvrz14Yi0hN8pvmWqOGVv5m2M4/xIW6JvgGNgAfAaez1ag
PBI5YxKtGeqEvmpj7DnpALyZNuAMtN/z5p3l1/1DsTN0vHA/XkmoUfYjAsiYiWqY2bWY6b5QXA7m
1IPhqpALn8fYiyIQQEfysfAnApI7wqtrpyGYuHd73gX4xdLT6cQayr1CKcEbhu+/4Kq6j4FJDbz2
FyMGQGvhhG6IJi1RgwjO9ezsTjJneTQ8lIXaFAoQFy0gPqXtLjIwzpQjCsDv2oNLJpK8G1BGkca1
9nZTl6/25bxosj+PEdvwtf+O/eO9RqrqyGA6Tmxcm3bgYmuNhLhbikClRzLzy6JboUWwu4eGAaSl
x+1PZ6DU+ux3ZwmepLRwfu/7uoMXuTuQPHfyL17aj5eHsYlAs4/DWlzzB71S3OLw2GCwYv63eHJR
TlvnKzW/tloW7IxnpYNwLTsw9SpxkYFHvXUnr0HCNVZkGtlgpY6bGGSxQV/ejloandb7ARSWDLQ7
MxdK9OpNMl3L/4y4nJCKuCVe+bfcNNbOaBgXJOJrygTc5PBp/yJANtB1ss6HhvwvCUI6q3+/r+vm
J4poYwIBin5RfeJtaBh6nPNbmhZyj5Lzz2cDnAiS0HvoL5Bxbqt3b0adZpDNxzTDzQqbTY95WMdz
caVnvrYeSmahC5qI4pdMwHx49cXtfYB36igY52EyK7S3U/LrzTpD0W5SXyIVTFnQys0+qFNGLauR
mLHvdkh9bDh+JE0JsBx5hwCPitGjRhUz8RECjuXTlAC7ifKjIUoNeXPSYM/qjFZTCtHp8SQYPX6L
0vx0tgheVoKcsf//kMZUyJ33ccUoFqzCwAIjpneHlMOY5ZCVjUWX6yNypoQLtmjUiZ6584jb+FsA
imX2f3u2EWopNLK0c0yOtpkGydOVEjx6/GqrztOJlnPTROZJ/Obc6wt0aD+tUxspFPf57ytbcc3j
XsIcD4rnm65bBsp8LjnL1lZu5UKrpnF4zSeoBpFp+7KXhMNClgzncDMmDsb9OhvxHmaw2RngcLMb
R76XaZp7zG2W9+3GOkZMH+tXXddrRkZCJZEpbNS+L39EO495kkGNndLMAfP3ucsi+5agDH3ExfKX
GQUKHAz8JQBNjGhIVKx8Y24qj848I8ZVXqS6kw414Q3Zn0gbLnoUq+RxCwXZugRuc+hyMDCklSKA
aY9PF6CWaQoSGeQJrQhK3rqKKwEzPe5g4qIIQoFs99TIHJTdHiXJiAQjgoezaiFerRHQo4lNclNp
H/wm7hSKTojtMH0XC0YVtp/7L4NBx1kxzB1MNtbO3VnoTTLz8+HG46Gk+91Z0b8jgjp3qiN3Htc2
vG8MmsiZ/ePLmVNT1d883sPk7Qgt1fT4JCgcFiCMRmFlaWOEGlbcSkHExmY6nhfB48So6+5nN1AK
IQcQROUFdW81g2NcbNl3Lz9tYyR8z0CzphVmWcKQ8e+/R3yyfchurXksqPlVZ5bpdkQiRWwM8qQ7
JJLsr5JjkH1Xd0RdNtW+OGWItty11Y1MVO1FsBAcDS4buKsjYBxVq7CyH10o7ZrlYmbpzMoxCnYt
IS+HEmBhx+JkpxEPoxt12/qUjXMADVsuOTG+JFC+od3xDUe3i29v3xSjOlhTER6WvvINkh+WsUoO
gu4WVmOjBdYicAgAGgI0mG7gDVjHpPcJfvANti4i2mM6LaXd1PR4IQp9ZRy8C7h2BZRb37fDHtlQ
bOHHJgh7Futqfht5bmnRG0f/UmEyCxvySpq+p7WBGcCHskYnGcRzt5wPhuc3cFPrxrr7YECcEYNU
Lykc5Jmkx/uIwoZ5non4x6B2WZCiKIRvIBUIYw51iQs/I45PNSNVAC/joXicrATQfRDfjRzU6S85
0kI8Yiy9o8T0/ZpeMAGlbHjSidwtOD9rhSZwC27REz//jWydwqRVbQpTOSPswFa1h5w4LjecnPio
fnjqqZl/THobR+B0F1oCUJfk/DhMk8GxAJP+Wi+5sTOZsh5pU2/pGn/xMKZuwe7zmDx3+druTKJR
YFokmCsE9WFRLVvbywTgF0ubA6nJmHsbdWXqUOAtjAShm1GIu+UlSuL6ruMj/XRXmK6E8NY7R4ig
/vyyBI35Z3314aj8Lri1+PMllIxC0HlbgbLAwWpN/2jGyS9Ihz8gw42jBR8duV54/bOtjq2AlUPl
IldzKfsrnSUf1bn9e83V6sB5LVV/8Vpk9TB7MuKy2lGWfiouPK/GtX64ufqMr3OwUwVUcbr9QlMU
zYhm7gxuHjYiASaC10qfRx7gK9PEnPnIJFJTRPFwliHvRv7BSA5h3IxFvQi+gc1KyGqsnObwh8W8
SL61uIzga7nPYb4lPWdMw65Ap9WzySJDrBd7t8S40Mc5sBDhydXJtgm2YQyS2i3+MImBR65Q8Grx
0QtP05J08rha2LOPc1aj7jV3k8uXZA/Z+wzQlwLZ28dohDRrV3xAfkCK8J2AJ95kT81tDMgjcPqX
gXASHyFnt8SDJDCQ4UgybTUGK4OMLFUoEWJQV/RVXHoJfPi1DHnz0ax+TQ0jZI+VPW9s7aARSJji
T80jy3emyUVM+0HO2Z23aJAGStJ5CV+9STvojgowzX6fSdI97siV9dvDiCCJvLfXmFObQWreGViO
XXtkOOaTOxDDGI4pamdjfWL1Rq8N8ngZuIlg54279A1DNl98hpdzigsSgumnIuMJv4vl+wRO8o0k
SJL9TFSEApGolcveroR7SQIFPWg7zYzXv+CJqkcvQCQnlLkdagytdVAhBCKiWmYDPSIi/l/0f43y
wqCNX/KuT3RqpveSWNO/16PwpWydfLrPBhOmBB+lgRYzHkZFTMWUh+8UHt1iA84scTWGAkUjg4rW
I3vjIwYikO4QMmTS4tKKPH2vkgVn0wWZTij3Qmk61X4rYl9bgo/wudkkmrguFwrwHBaopOW0v2Sv
k85nvP26QiqJk2+7GzCmebOrCVh7cPgYx52dwuPTZyO7ca0FnWyEDOE1HAwdewv4aiigC0yuFkZE
63Xf/qrw4h51im1XwDU1rA1z3UTE7Na5mGpeUxafMuCbMAGQCtq+kJPi2X50Y7uKcVdJ1J4qN4j+
34gLTIuLlYTqVwsVEIaZ+5TZRJGmFR+xlAyZ7SLPM64CFveiBoNKKFZ4oydS4IBjsRsKqpccQzix
DA2ZONSZDJ+SabgY6M0fKlL6AQ11ON3FX82oA2OZiXpzcC+FjK+A+J9d8tsGtZCmAIkHFAq7QP1j
fZ001HlXfWPupF0oYvlBP3KNRpXceZUzGiP6x3TgBwqjatA0X/vn9T1tA19AaaMHXm0qvgYKtF5z
mSV6jvODILbll3cEaTwqxsJ7BlB+GVlABcGzJRbAM1MfShFzq9UdITyWFVAiLnKSLIAJYLHMtys6
qgSmyFAH8EeThjjn8Uc2d3xyZ05eKfoY6xVTdzcdbWYS+ZAObm+PUt6Isunq69MLQ9fup+I2df0B
PEqqKKP1Xnl5EWXW1X8mcXhsJfYOB/4P9CoF7bgYaje0aBMIg9DezANBwJkt35xpqzwFZm42wbFb
BUE4bOl3BdKuXCs+pZESSeyZcI6a3t3h+gbiSNCEKPrVTlFt2BJWs9xUeCefHoY4+kVGpvTnfM3P
XzAkV7LWKS4X+iJmqS/hSpTL2id1h1LfvwuuKP1XAw3KUDydIU0BmXZv/wCWqGnambLB+wnCSmuB
hxubzmgpUzcZsbfglp0xt7hpGvetkFudXGcy8BWxVsinx4VkIbN7bdQXRxc50c40t0JCsObDSUyu
hX5kS06rM5uCk7/5fTL0v4h9cQG98t3p6JVOUb97LKbWQgQWoRI+9ktW3mTjIvqvqkJ/XojFX30F
wKfhSDiBPaagAMys55EZ8PCiBRffGFGg5grl7RBS0/rJbNmiyYuRI0Zqbd3mTrId+a3a3L7OuOKj
u1b3Era+uhtyQIv/GZMOMes5bN+2KdA0pdHPv9zH2cFINRpml4/w7IUiN9M/sLt0lmby36mhjov7
dhWYUULFCG1oq7GclAv+UbbZT5v7cBbNU4vS9GEDawlU6hS4uMsAD/Ii2HIRmySGKtLoi9FcAal/
9B97BFEWJ2Fk2f4dlkwtapBOQ6cKiHLb1P/Qrw1KWQ7kbmsDCFX6mRLsZwDt+eFYoirvIJjoFlRF
S3TzsXrQtnTwHf4BoDHnH3DBEgeu1ETEoflAaUHjfIRLCtQ6vjiXXdfKBom3EL4AydAxW4MLr4Kj
RzLIJVoM3ctHAK4Y/GA4c5rKVWXmqrV7XaUGWxhh9TFeo4vh9eW72yI7dOu8XYHQTSaVzIliaiuA
pyBfQpVvtd/+AN2tTV3bxg/Uuvp/8U3YIX5xt0IQKKR0NXyjbO1GWudt8pc8p0dYf8U2BuRy1QFt
L1o6IvJMIY57DAjAt/OMwwtfsqJLv7caFfKYQKmOmt1SsRDiJ0/fvFJcS0QKEXUcxICYrhCcy1nh
lJopM+KaOWkx7CD1zIED5NQtxkXIKPNUxNRfYvrHs+CCh5PCtjR4rIq4F9lKZdzW/Wzt2hA6vj5o
O4IyxNczXBr5qX93928NVnwcGd5SDUFXchL8LX06fN7p2KT8iIXifJN58aWFu2W1I01pwPaUQz6s
qBYxvchNoGjgH0Ecn4MoM/J328BSAl8RgeWdtUI8e6DcS2H1Owq3l13Oo0nyN2TTmIkHAYucWpXQ
ntd3Y1Ge0KToqBTj12BTJetIlYdpkOAtDz9TYRnKdYCDm4Ksw8eiXiD1F2XxGTZD+/YDoAHpOhN/
hURX3CJNS/sH6ExekRzyAKDD7U57b8GfchTWA1jehSSSCm8ehHFBBYU0srnMRwGIAuiyi8GzHlCz
nBIYA8WnoggxCFaoNwT/E3HlqTX60mnKjbFIB13Cj1Qh4ud7ubH9kEt7zSNhyuE2SOur0RYDF8IR
SIsYEb3cZUX/Gv7HBv490dLbkn0nlAOiUTa/zpEMnzsMV2fNN1bvaA6hQst+37p9wDwLzqFHGTE3
qq0LejV5jd++UtKJGDqeIhlWTTGP1vge24VgIJBoldVSqZAgiIC29WIuAgUooDkXfwZbSQdnuzm6
fSFugItVsn3zpN3wBQ8W80WQEgDGvCAuQElr2KPKunBIZXVVG0vhuT4Dd1x5m4B5rJ+stYiBg15s
qIqoReOBVT79xkJp+rGzOiEJ0+8blAbgZ+DW7doPItvaAMvTZTgBbfcCoCtZYqoWD6UDS2JFAg7/
cxZhviQ1kIUPqTLBD0HygbWswncKS0ja6GNcT76MoWy5ptINAxOlvY+2gCb1qFUX84+GNwuQrmlo
ddguAFMidqyEkDUgmvg0ivGJhuvQr56CYaHhnoqJNyAyicuGxJfleqMeUNAKLFkD4+HienT0mamk
jJ49ou30W4hHSYkKLuSJL2ZtRDSdV0yyJyN7AdX0LX5w3KMu6FM6IOy8juwHmclXuy+WyJaDacyz
TjqVB/F4knO+8PnrEsSfp30qelq/nd7E9eA1mdzV29Cth9UKhRSSg14vKSxwlQ8KarR1jjx61R33
2VRudA76NHukdUpULF3fV6iOK6zOTIf1yMm3j3a6KDt3kYEGgTU4sv36JUq1gr9JIgWWIUaNUV5m
bCmpBH8llGV0UPgza+t8UgETVygMupdQixiY3KO7kBjGHUGyQ54CB4S7T0rBxFEyNDOgEz4Uf6O6
VFh7EN3eeAmc532GId1pTI7gZvS3XAtFVRXB6rhjqi7xun5hIC9wxkP1IvX+wvpAYaf350YImPl0
EZzywdsBUjCuXBFqMH6ktxCZoFOG70HO3PIJvb/6l4dWyQjZdFWSSvmohFrNeWh8hROnl2BbucFn
JzYbH/xmTf1LLQ5C2p0cxFp9D5eB6rdIZ9xrEHo1+HCaAeL9ad19xnjOzcfHu7i8rdJNrJLRjaIU
sF0NzC85pcU0S9bM8Yq3nuO0HoQKbIe3v4m/B8eJJadk6Y81REHTcOmr7sGADBZOyFdRlZa/an3D
2+E9N9x5bH0H3aJBN/M6axKL3f53Fux9xw8WRp0gs/qc9BM4iLRTOBeARCqWSJley/G69w0XVe22
Q1BYSSnAp597erwL0a7u3+gRibfAw/CAmR+s9T/VQTVeFSoRx0YrZ2UHd86RjKrF5wkGuKsLT2j6
OdjVaVZaj13FF64+9YMSWzjBYQBZ6Ow3Xy6KaxIWtpb12aMDKhsuKat4C09cuZ4dsO5y7my5+bGX
ZvtZZZFsF1Gaiak7zG0s5bnbh1orYp+nkfzRn/CXT/5PSS21lYisbKqeeCbot0jzswj9Pl5evauG
ov4yoInKvG5vhAwASPYgjpDVv1zHtIi+fq4xuX2Mp5cD3V6XgFXtEkvHrHNSyWsz8mc0B+7TOjT3
wgGXJ67CuUIa6dh/mbisVvMxYPX2mt+whhq9n46SvdIEoEEhAivZ0/a6hIKUgTWtHFqFNB6NEURJ
OvO8Xg5OICUbPPU+o6SkNxrKo/2e8xYvAYGLT+LU2vCCGzfr93SZG/hOfZwak6pYOtOUXhFisE1z
IDGQP+3L3vTmP4QDe4NZo+Wbtfj1AtkwZnaby/8CV5STXYVu6zGdmtKqu+xaIwFtjXzW99Tq1AmX
qYbUx7J8LuACn9nHyl4d1RihG066PyrXbGEYMq7/Xe6ooxE/Jg2M+Wihwff+H3sQ4voQkNZeO4Ge
TXx9uvvIGbDxz4Y6mKeHyMhI8iKMZLVz3QVqL/2FwiVpEOuSxc6VTVxhxT4MolAn2MCvgf5VQm1z
6caEVfCtzcGnqq+uD4WtRXRVKrKoYXjB+t+Lby2NQ4zwkZRomReihT+BnfO2/WHO7e6Z21hePpM4
hiQ7ta9saHAn5MfxEFcOLgNLPJlJDW/DS4d5fqXXVOgcVvwAPPx36KA0njCR/Wz7UNK/qoWcTkKt
WYNCMc/mKNo2wP62XslPDm2DHztDHjdqETZga9OMjwq3+qPf2CpWQ87YUa2goqT5uX+OtwnY+iON
Vrml/GkZCRzuFZb/UNAqVs+pNSRkqAJ7/fG9EL6bpg5wuv+I48PpnwsjCwfnz0BD4T/CwNbP3UBS
za4Ij+8iHD2cB22iE9mhds2a6Nv9YDZWLYXBg0y1xoZOVsexEoOSgZDXQw3xBhyWeGcycA28NLQg
BtUORIbSL3zG6ExnuK+JQrAbcMFGfHucAuoZRtVIQOIYjBBkJwgosObFkAoYZcc4QHe3N5TQG/ta
baldijLnrZ03htgSTUfEP2zhovW62AjJ7EQuv5wgU6v/x48ipdB0BiUKnRig5YhLI2br64AmP2F9
GXBRbGUQDrQEMVlCaOJVSQVvAoNMZS9GChGVhqyQ7ljBLVaUqzOR3Lq2jLsDev9u7sBFHHa2wUSJ
nYhy/gSGr1lx2eZ9Fo9tedjeknaYNmjaOik2P8t0TxKXsTZZVmoow5N37NZ+uRg1EAAJw32MY5IY
mBRxwk0+Y1WpLr80/kFFaUsaexcosp1QRK4NkVxkzC+6AWFnBYt2sdSEMD1Fr8gLcvO6LHMFUS1M
pC4oJL8UMiu/WjaOc79rzFU5Qm0foycfMK5MldMBmhbHvBXHVHx1MbhaOkrU+mauzh3zenheUuhm
ZLHPEr0hnoRL7C7iyPIHyS2ZBAETG9b1yZxbppwyiOc9D2epk2ooS6Y5j3UPQD0x9BvtDkzmZBdo
mFna0NdwgWD/2S6ra6PVl8N/B7WT4JuksMsCaKKDgHYQOKtzFnHd+VxOfzEC3bzd80tcFdOuHiQs
I0xJ8HtF5Z17S4sb715Hgw3iZuem2+ePiyrvho8pmPwUQg7GPOg2ZVx79q7PaK17Nr3zhqiNwAZw
UshU2hG1s2VtMm/BHe4FKkHid0gDUA4fxGGrMjRJv1SmGkbb/rqetAinYYtY42LCMiptjNfrCAga
tZsA7ntRLhTHa+x2yNKZfs+1MO0DflSOeXpSn6lNLheKBEpiac7lGB4ZnkCLd9McogMv8y8jcXkN
5Hi0OWCNdnDSNN6P8L4MPhZsT6cGacdgYdVo76rf55MauK1ynNrbedKeiEVk6smwi49f0xMF7x2H
SBb4qzhSx4b4Vo3suOoQ3IEHTm+mQY4shtUzOLJMVxT/hvOkGh+HHJRMb1TNRLifz9adKQIZpvwb
tMh+dxYtrrjhPBbOp82IAr0u4U9cjfqd77TnwM5GyLxpJ40AUgse/bIbFiB2IkTrTwqoavDKOwcM
HHudXVCUiMdFhRLLDjnqkalyBXn9wZR8Hycc1DB2S/EaObz/Yhqa0zpjbTpbTpCiQkmjzI/6LHMi
P2YeMziXQnQayjvNzokUldAIm+fhDTAz1ZhON55xS6Na5w5jOyjixy3vdPtVChKAH3QwL3kzokeH
2e6kp1JSw/Jco5HPR+CUYjrXMBBxtB+lpUKDiZrcqYSfxdofr+0VKDZb7ExkXp1FO8R798aRvJ/p
s2JBGKHTLdTOhaIXutAlfEUYyiP/7XvkclEkoQoQDHGuJw6tmf/tzcSTqhtWnDyU0Bfomzjm93xo
URwE8t7zWgKvZu2KmZVayQ25OJHyYwJXsxxWNrM5FaxLuK3mhw5UrfUEXIHzJavzQ5mMXvetLlXR
YuEP2m5u2sm8hHILtqoZdyTsUkXEKxpegp2O6L8G45wRNavIMmnsOI8BRh3t+jfWApRBOZbpUIpk
/8QdmPiBd/8v4Tn/4QBvqevonrACBdrTqXtaXd6gACKBI6juQKK9Y8Lwqsbecpaj7Tnt+3k7gJHD
TydU225mlEFPG3WXN27KrHnzru67b33hpgQqagjX2G8Ih8jvXyzKKpQIPUiqe0+Sgm+zEMFYYbay
dTERUaboLUCsNWEHcXQnKB6ZlFhtHFZwaRC/yt+dpymDg26pz6A9hzveX5pLDzHowBNXQzeKWfTL
biKNwN0IMp/c5aKAuNSESPhdZ/vrMbocvXQRaGvZRp8+G/2eXSnmw4ouMQlzw+oHwh2IwzTNBwdk
Vk45L4Vfr9djEviPt5RxfvkzfMiSGWlk//XFyAP39mMTcUt4uWkRflh90or8df8JjdIGNE9cEcZ4
poLOzQzPszZ6ozl2I5ZS+2H815d4U43FValet4qirsIs9Lq3xIov+wzQKTA9J5V1WhMCScx8OFd7
rRJG/tRm0UoQ6jbFNhMSbdBMwJZhxLkLZ7c8BNP3VfYFbGa0GRebfCoN5eScHP/LxB15dxRMShdg
5L9N1tW4OVIHvGyRlQC32YhzWS0JDIo0/PJhdoyxkhorbvq6vVVS6d68+R5Uc5YXRZRQWeCQTxEC
2zxHeiWCYLYZi1nCK8fP0PVVjzG6DjVbYA86fIz+5FyMbnrlK77ZxN+PmVNHgt9hjDPj8XMJyL+G
QHheE3unZ4vK+I77IJeKkyVshJ8F+TLxyKhfnvstp7WZhyzBBiMz03eDIfEwz7u6L7YuwbcTh/01
d1/8vwdDEAnnO55YsIEsd6xmum/BctEbOYYK+NGpbe/luMH8RB7pzBRb9EC7/V3sbQ0XxjlfQezH
G62I/SvWDPOjKaIrs2PNXOq9j8Vgpkohqe8K5fROj5wI9oOfBeNeOgLN72tALjjPlVJG8vV9MkDb
pc3p923/umodlK59IfgbYMaMdEE1hI4pMoyljjmK5nIkZ0h0idKMNG48o3u+0w59bRFXk3rAlBvv
snnV5HIEfbxmRVKJ5qQFj+zGzBS1nUC8NZzz0AHi/IQd5IyQuC/fvxNG8UXJ13W+LySBBInPMqhj
Y18vExiLDUnaNbD/fv1O6zOsw2qr3b8xxlXHxAmoPQbeI9OpJuuFi5SJSF4gNhd7vsA45hZ9KrU9
Tm0pGuecORVc/MTqJiQ8C+8D/9loxm3p3bV4ZMCRuCQCskWcullC2cdUUO2ptyJp4in1MErWUNkY
E1svXlL50rJOhbiqW3YCanOz4f106gsbTU9Q2JUud01RKwZNe8NYj5XMcq6Wdg1DJnd40lTGDgw4
d2nOkrd0w+peeea1ex9Lty2vp+6GqbJmwepEMoL2uFls0fFZRKSIXsSW9bGkCOiNZ/tpn7Yu4iDo
qIR1jZhd1GbMQc9XBShIrIInLbg43D5UexLT5jLAHYCYDs7oVLW4rkiozXKIEAg2teGNQByV6WUc
Zsvg371dEZ1AfoGhttRBRjlbPO/ghAMYjXc8u1QJAc1C3UdtziAiZkM/8QDR7XcA8FnOa9vbh2bH
mJ3tZ9Buoxa7N9Roiu9aT91YjLpFK9dQK/TMHNVin7adX8/BU7fYhC7xC/cV2fbnScDlxLK4SrMt
aadbTUVEiPQEwmj8uBr2nexnRl3d73yZHUsx+xsPEp3GQ4j7Uvh+4yzPK+nLV9Deg3IsMwU+sCvq
WeJYA4aOSNyf1+5roR9tftD58ed0KNdbyMUNk0LMrB9arBmT//Gs9c4VYHCTtD/GE3k1Iq3Rm4HX
YdFkNNXQXLAwmvsGCXr/IexqFf2H5QIrbaYhdG1jrDzJe73EEfEXGwGbpYhGW38MG44Sd0mvDRON
EZlPT5an//Gl9rAuB/UXQyCx2KS6GXi8K4FLfpbMGV0HSgIarjEj9y574O/ooLZ5rNmKT6SGc8/N
xVNcppoy5vz11yvbMcBks6LjZMu3+hmyrMYRbx4rJ7YBkpoNSXo3DHauN8Ol8NCTFArTKp7+p1O+
sMSmrkPHeyjb+9R6yQ286DAaEDhXOo3PWP049XBF8ctGe1qI1DVjugjV4l3ENphLJrQcrqoowt94
PV/grt2Dz3WxUoEokgG8PvHLdvLDbReXIachtvdwaS7KDcQj2DZOza54ztpZydzt5RyrukugROE9
jADTWObacm99sAIWyZD1fe1o/UgVppmJXuFm6thyudgHgp7TMm3h+ZYQES//Ie/8Q4wGws6yzwcr
O3zQCzyjnE46CkvGf2PIpMpi1Xz7+21VPi5NVhxaMEPyC5AgyNxIVRfmqF3AaCWnNhDz4iRkd5ql
mp9Q1L5sSXwZGnBaQMDmaJsdT9HnxH1gc0dRTXM+A/v8erzPjRJ2Uh9btv4djowYaDAQG66R0y1P
9SWKMasFxUMOOLEbpiqMt4KOci11Wlzo8VkAoRcNAk9DeDQDAcrnwLOHXd70SGO1BZ/Y/cWaVQIX
MQdZruvD1fItReLKItHx0ddWyFN9THWHn4Mskhy4j2bGmlT2xm4xm67yW8m7VLXj5Tq1sBb0716U
X9CFEOQjiVZOpwLsAQeEB7eO7dwbqhbvQRU5kNurRm4ZBSMOzhtOFf5OVWuPHRD6GG/XLaJdXi4X
nd+4FFWEi33UXtHuX2EWRIbidtiFMsYFrQW5qyfAdTSPkB3ojkpGpjU64IU72oNHR7lWybxG65z7
YHO94RbBQzElMMMNHrscHX7HaD9yhCkP/xgWoGamevOc2b+Fb36rsCWvCK+hqwycBLA468ow6Fyq
1fj+xFUQ+69q3TJKHzCQ6hUudrsVrUYtZWGmm3Pmw6eyGvw8WMm0l8d2z0E0hUFpmSS75p25rRu7
ii3yqxeKe/N5Pl2dKGF4wcmxwSh4QGROyzrH964Fs9X4fOFd8wIrR8a6uwKmf0e+QudcN4DBeFHK
gXfCZzvuGLyme+lbaW7QtTMd1OkS7WVmtWFqElHJMpdw/WkzQdC6OWrmeqQjaMCkIabCrNrL/b8k
TnsHdYUANIv9X/YgEo+6R4nxg7jF6ZPlkQRtIMX2i/AQl8hQRK9XnVt/JFqfBStnEoj94BoVmwG6
P5DkX57mYYLMPvQOpcvqBT/LlRXNxSqT7ANJJqteJAwuPd7DyWqjRKlSdSukpqmYovruCUKLD6b0
7TVyaCtzyvZmsOrDRxj04mMMypqjxd1VB74Ny9uicL6qpLF33YLD88IDAbPMU/EsIQJSsAy31wZ3
sNBM1ZCWLTdvwGJMipa2Wq26XUoeP1IhCS8kp+IHQ6EkDAgjcb5ahosN5pJBj7mFq1GhbUQ2BD6s
GJwtuEL3gahYDrgS1xPgruj3dyxiKwrUYBFlnDEEzfzzPXY7RxYIxBdNY8xqKx+sYw08g86PMGWy
nIdmPzTG/Ee+FzffdDmvQlGGaSEKB098NIU+vRZlwAEAQQU3Adw9Cy/iNn0B0Z00ZLBaL+rC5n8B
29tBDh0NmHWhMxzYeY93eFE2+QJIvgk/TLRtKoO6/ZjHsEkCEoi1heNZHcaYxpWdQP2aLev3EZ5X
LSUe4p1Pu8gKK3mRwR1dDLKb11zZdtR02tjL83IAYO47OExgkvne+DMjE+NME01aPXH5onkR7FVc
NMrxmsCquSvcB0Fryso4gy0A9OxtBzUkWS+fcgLH6vP+GKpPZ1S9fdR30gKaYMPVNOnnRYo8Lrq/
mMDJlXVjtOUrI/TDYZHhyW93SAD60IvFnOA1Y+qtawkucTlVTIilub0+dozcEwEr6ghWJeJjz4ik
9NTFmR/H+oy8Mrbnvk7IzbT/8f3Cs8etGe+7UrO6oG1tVmj0YhMnZpaXF5ugCmT8vxSuBTd4PhBO
PVGauo0YND2M4I74uzFbwDGdW2P41u+tt8a99AhK7mqkHB+NiwWOJRhOarwttLkLCEZwYklaNZpa
vjv8KVX5IGsxHzpU48Q/SZrpKpaakRI4uOj4mFqktG13VNX997LZOaQ96iLxaT0QY0q9rKoRCFQi
8mcRscEyZiSI0IJ248jdyiFDwdYFzky3zUY7V+kADXbU1/FMiZWX6oP9b8cN07tDmtM9X0YRoAFM
F86iZcD8I+E54LXvSjU25EClOMJKAWslJgRVHRgkltf0tHH99ljm6aUWa1EyclbjON5nTTywUZpR
yKp0ZuJ37euJc3U45/AGzd+TsDah9wIToLCoQjKoWGfAZDDafmu/ZphfioddOFBvSV5s2o87IzTD
rmpLXBGbrBzIqMzn7Cxljj/bTXkIU3w8ATmBMrRJxmiPwDOBmvhmZPnsHzWoy0pQmensSpIFUCNz
MVwvg2C38jRvLa72GCgGXvXls4XuPjYHMAL16C8JNuBbWjJwK8zXojxfpxvcgf5Ut08nlsSwyFu5
4uSdDflgO4MuN7wRytQ+SEhx2E/eOWC5DAdjDiUo9KX3v4wBc4MCICDCnFhshTj1ksc1gaZk5riZ
JTy05QuU6vNxsdz4Wjyt59zo4l7Zjser2GHxg9UFbrAQvO2yTMANbML5bT/DswFJYZtaWn4w2ekN
tbdyoK4nFmaoUKUjx8SmqgbamO4lxjwbrvXrSkdIUZMnAPBiCbtVXjIYfYxnF/wUFytVXJtNXByH
dgvWk4vKHStclhbWzMZEWd8gMfJiqGbxDeCDujFtfl5XGFnBQ1GG/HKLgYzmC2umhWb8sN9erjoT
9VVYMaMf/8VNTXitkvsj9REqme0oZNUtK4up1tr5ckIQMDXFWiviIQOOHudIohkWjvPx1kPXgf7U
FtByWJCDp+rOlNxrhbY9+/gzvLYMibz/qVUruz5Csl9byLZ7f5oQz8xWwYeSuVukW5gr5jnvFVGq
03xamIu/TAHEPhdhuUz355qqLzgpUr+f3PEqAc1vgor/Uq0bbZGcuZTodPl7kNFhmbLrSZEdiYJk
lnGwH1ZbZikUlsGv3YHfZXnvJrEkXPwSvRbOfchcVEEbZnhlLhLTONM2P6IhoejS/HD6Uj9/cCiS
PQjNNFn4Y0D6S5gxqvvghbb2rSuQI11DtVZG9wfNkOKUn7NdPqwN/Ql4f0/2TwjLSGG2aN3h6rPL
vElYGafIPBWsafHQnUwVL96KNOc/8/b21YXc8v2H609We7SANj5QC7RrwCcutnyXer+KJZXv6fXr
ItlxHJCscbFW1duSAaaH60tv9SAcEdvfrzv7KbFBDvYgncQKc8IWqvu6Qd6QzQ3mkxrYmB+xIPjJ
QJTDONWWpOhDeZ0QvtoOG5ndAiH1ufkKOgsgv7KrnQ8JoQf/Fo9d5VaIXHfog0rkECfHpVoJOq+u
CjeQMcdeYUY6YWfw2fdrF6pXi/Z72IdhfhMO1jSTt4L/Aw05F5qdy+C+pDeZlES2AUOisUyH+gNM
aIL0KQgcGGcWz6n85hPy27LZmyY4oDy2NLOJ/Icg7mpNWAU1W2Hcylw8KE61/IKZxZsmSLPqVhhg
mAseZLIgMsStz4EWVrJ407BrpbejV3gUElSEjDdD8zxjxvm6NI0azwW4QSP8pJ8GEfz/vlGVoKNZ
dxN/wZ9nVPoPttoGuBn8fronC6WXsxyN2DOwMF/HtmpJhRJ5JdqeLPhiRdOQgyXtVEJlsFgeHRRp
LNa01/uo+nA1s2sZClEuDoXNzTM6U/XIYRxifUmmCBsqHrcct+0nJU72aJowkvSVWY+n2GPJz8pv
//2pwoB4F7ORiqre+ATaflVRz6u7VO8+tZcsyq6wp+wlTU9Xxpg086qFZOjAG1s1JHCmjk6F3bL5
NZBwfT5k8iYjdT2gDfJ5x78o6FwsRaLC9pns8KAgS9t2wXgbXOdkQw6fDHvyK4KxzW8XUmOaE5S6
cxvwSfpS78NNySMTfxS1AzbGtnSFcS5wfdl53KpTThe4hZkNWgA4NzQvfsZ4WaMSP9z7dmJgfGMn
7RcwZN1J3l4l4nvuPyycYuzbp6ZVy3fMBkMdjRqWw7v0xXR64c98S6WzwCvQlzJOCe7Es0gVS2xJ
HpCl210kOuvcbUz0HQ0kEJF1I2BnH+EaIHcw50osQC/2jgfEvkajQ53l5IaiZyGX5pDfbxLq2tC+
SNZzL++nGSJviQCUa1zuMvm5AH7bILIDFPSzsL14m6FNudjHmpiM8jjhxi/c6E/jzmjBK3sohiQk
LtySTSJ5RtFsMB6/IiSLd7PUi4pstRN+YZs7jLZUAhPY4XDZEdLX0VpPUyeMNfpCPZRjbWlI3Zas
+nn0bb1Zw5H9oeFBrqGhfpGfH6z+actndYeqWH/XtpTVclqWxHGNJkNJ57PUIuTkk2GPt27ozjY4
IHSR+ZbV4fhm5II7FyevT4N5Y95QzdG6IuJKb7brjbzZHaO/ujTruSub63Mk5356htjg6D+UrIQv
OTtpRpbCENizgnfS30K1WMkZy/QOlHJiLvybnlG1ntPAQ/MSh+QMiBNzOiHTAdnHpRrnLzufduIf
RRMDVi1qxdTmGNSCKEYsSoaEr8vFMow5K+5V3QL4yRzVp1GXIAw0kVZCqHCuyRaxP2Vlcz3Vd4Cw
E0Qz8T6Eei/AXgbjBEfJ1hhNI/m4wI37i3BIwr3gXQmd9ojtnAZFLmLN8ik5q8EGcI5nDiixu7vv
eWiVtL2l/OuH/yhMpCYF5k47VR+MYYLRlzUi2mvb/Bo104TYlsO7NgHcANhsNnhtXrGomOzJ1SDN
FdCHN0ebDIzlZucY2wUrJJ5/lnU4vDD0Po+S7OFjFwcvqvvV7gZWW0KLex13+I3f4Oq3qZ8G3y6h
ZOdnfKLWzcb/Boqp5UNIv88V1P19ztH/SMER10jaXFrqz0r8YqQYmsCUmQT1VNdIxBYBAQ2gapBY
Vgzee+1emPJiqL5pK583zv/m2j6nwv4v12YU2WPzgINoc7PKFtcobnVD6aoIeu2gkk+SVrikey2a
Ru+HOthSjSQYXC2miUpFyE8zl1Kb/hTdLTzeAcoLYzvAx4EKj1QTp40yuIzgZvl7JxTpQKpTnAp6
p/+7MTXkotUOAZqaiBgpBq2O4oyu0CsvVgcRIvaBs7cZgNnA+vmI2LkVJBhIHKyTKt5riayN+0p/
+ymzsZW/6NYQCV/hT0yf0R7WoIP3WZDEPgG2lGLe6Hk5+7c8gsayFXNseRducUpisehwzRrBf/iA
9Y7+21ViWNVcAmRO1rNmwm9e14tVHOu9K+CLl4yUHA2UgMDpcZyBTZiJHYEGHTtJhV1vlMe5tSzG
haXlzKkEgofMwozPGotTzl8qzBDFXLtLI2wgYX2c5eGRmrGzyK5cIF2jrIXfddW/TxOrW/yQ211y
567/tHJAnNparl+kBMBJVyYy9AlbAMy1k3mn+Wj5p/5rkK/TYXTr8BxFmfskoAEiQRc4usppjX2y
ODgDQBJ21vzn400nt7ltQbOG3BMdoovkKEUfMTGijsG7O2IGDzWeK5OzaBQ2P/mnxKR29U8aNtLm
epoUcvpbCj5vJTrj5tA8FLffSs9mvaDU/tN6bXIP0xLBl4nrT+UPtter/2LT8JFHsxckuQ9UUu6s
TuvJUIxna5BFfWQDQf/Rh3JOLfqddGA2zByZPtDmD3Kv4UJbh8Hfvq+9vf7sttiibZhM06V6SB4C
3ruU2GrxmaesO2QPYAtW1Bv8reYwCh3XMWcUisPJNI4cNihDFk2F7z5NzCU4JHg0uh2NPXKWZaQL
rCQ3ib/Q7gGu1Vcz/4GwM7zWop5RaZfY3dYq14fbPUKYUpS2rw5YLGrXea7/ckCaDz3mul/TErQl
9FeycXWcSzHMFp9yw64PM3Uycxn1o1COtHm3La7hvHMxLvf9Wyt3/U4ilaYz5qQkDn4yHeWRkd1f
/iDvaKuF68fRp4z9Q/t7zb2gh3odvbp4PfC9CyfNFuwL7DX3QlzNfDk9ztIJegje4NFYJjESYSsk
1KHkA/o+OCY5Ql1bRxhY1P9k06wYnod256/ryLppjCeD6Hb9taCXlZJiayMQ9UU03qWVuG5C0hmz
jJArq+kpV9BMTur/Xs5tDxcEcfL3Q20skT0mpuY2ERBExbVngvXA+tajuxVtVnOE132t/RC4Fsdw
qPJdyyBloMWjSFGqIehWjIKGxW8fX8KCLowF6JWTo1T5CufxlYUg8b8UpE7WAeia8vzCa/GVv9Fz
7A8MtL48Gxh8TXN1Xn136cMRljblKKOBHM+YwKlgfHvOt2O9flZsFBQy2BcqglEHOlxHjhq4sNGI
rj83MjDBZWH4ORJn3tGlyHyE+Tu72/SHGM7XWzb52KP17gB8D8T+89BLiBBlQs5+fmYpSPPaHoAK
k/quTpndcOr5S93TM5eP9GUyAjlxcJINIssOrjnpJdw6BXLhTrhxQJDcdtH1X/RtlXgtRIOvrjVR
q+JL0C0sUK2w3Qg6RdPzZb8sOuykPaoSDDBA6QqAMC2VlMF4j4a53Y2gUFg5eVY+m/WXEPJjyqOb
QR1Joyvt3Ijp3FMKHOA2hFHVTrkKcAIiIME13mOhbTJm4JngXHppY/3QfUQMAgT7oq9xeMcgy/pv
Wfikgu+RWYCtLysv+lpv9oLtfkkUzuLhNd3XsPaPqUWTler6w3IRGWgWWasVzMt9QbW3Hzloau2r
QKr7MCBbk3O0hdrWiHR8a/u262veJ05cwcp94MVQDa1skI0hCQgfb3d5lFhoDQjqRU+NVRMMSEHk
C6BVU0HA6fytCGOtVw/S45U946++OEyWD6L4E7liFlH/7e2ClIQ8swLNKytbwmpEtKoOUpMjUPC2
Zh4GBxg5PsvurXwGB3UUij/3LKabTXcJZV+kaNCbSbbCIdNO+uQ8vR9Fajf9kdjx+qrQ8PY4LOkz
LCmuUcYj0pwr3pIPFyUdWJNExAtCMkxL/d7AkKo3HB8bM9gz+eOGykryvPCBO7uwnUcCF++4r2Sl
Q8PD4M+KkbLAX1iVtNRm/VmvaTJy4s2f0/MwwPUiMOmDpvtcUMwlfDqRHiCgSPCS91J1QVTMoaNQ
SHiwF95qQ2Wj0J5G/XxoQ9fy1N1LlH2IY+PJlLsoT4uL8dBe+5em/d75Dw++pod7OQx4iF8mKrcG
bshWhEAk1PGizD6CXeNGnTOfh2yao/Sgt1Q9+drveItSbdPkeve1MmBWQrLAhpZZ0X+yJ5IUYh9A
24ui4XOpSEgLviprYGR0tI1Mam349mPfX7sMMXf7+qlD+xyL0VFA94ISrimNuBMImxqUUtPKeJJg
HX+ufa2TkNKRvNhER0CJ4qxFNmlwbeaKPFQy6DSl9w9oF5hZ4xrMT4v1kBfPfQH4K0O4OZ26jMFQ
qa0/PCjwodxlIe1PYwWn/0vMCmTAOGVWwbno4UnvW8OPP/BTnUE7pUMoKgxIY8moYsNQ6BT8Nqds
SkejsxMsfWko/gAWaEzEW4PtoBtsHhKaBb1q8p1rxkvIUxca2Afw1hDkXc8P/QCG4lHYziDTI8qu
+qnhcAOgkqGteUanudbUuByqgY70WKGzJ6B7UbsVYTqBAcqnxhzNqPOHeAJJe+97gQiR28DqFr1P
+t+yjR1lArNinervQseXuoB+LfNw31Cunpl3MUk6dmV+4sckbuEj5hVjZg+oT45/xev7zT8ZdFnk
ga3yLTRPKUfeUJLlBUD6KpGFTX6c1LdBkWl5FZKY/SOWtKUsAQ1tKs2ityizC3S3KXP6uKD5ndmT
fXclxDxMiJEyDxgyzJcFXTElAiL6yXhJmPRD9kfv3ZG0+gL5qM+UNT0uTmou8ERax9fK4BE078JE
nAjk8cC44ItHahs+s9Snp2LdISfN5Q9HWtcIYtVH9X3sxHW7ee617otKCIWvYWs0X3bKZNnkQM0k
s2CamG3xtHeAFsOxwfqjMzvM7A9kjSIYRnR6bRPo2LteH47IFGkrHeE7FY7/C1VLVtloV6u/K7Pa
k0VSwjcwTMlfe0Ecol+/VUoNf7CIHIbOf8U4rbKevzUxOUHdanJrIZCStrpYWoApdMmo0lhk93mg
3OmZgc4oKX3E/o9NtMXtDpxsQHiDmHOK9TAQ76vmgiOZ1T6r0/V0mZYLrxwkdkUKl4bOHeLu8JTo
oJBRvUA7dkxgQyW6RrTEPOh2leuaRBHbxYKbdOMH2GPpV0p397MR42WyGRHx6zt9jDLw+KzM12sD
X4ZnuA0BRNXi8W4qMueUsjE0RUP28nhgGl+fESrtPbhhEIlkHjW77VYQrha6CXXEqXp2Tep34Y8M
nY3+yGfGl2062rZvIXjwFkAei25F4JaI+fGSPUNMz7R6YiQULMcxcjQtJSLy10PrsmVG1rVkcUWA
jPYxHrU54H6apuJ0CUa1h/iBgxgGqKzdK3CarZ7yXtyEOtJhn1uGEWuB0yLFIzrgc5UKgp0XSmIB
rgYTrCgjmXdEC5Ls11Hqlj7aiItRNXHxkaU5L4q7nDrrtb0pr05vWDY39gAEbRkgxQma9JL7PSgE
/Pr5lZuq9NY+uU5roSEXEUnfvxMlEc8PLqRUsO2axr+9cIjPqDn8j2Wpt9Czp+aHOlbZKFQ7NEdQ
E1qR71v4/uBScxsAa/YLGupp0kzQmWkSMy4p5nyhO+Qd9A0qBb2axvRoTSJ+dRiTZXpepzaON0pn
qbAT/6la/3TzqF4ZOKRXIyP0CjsdXYmO7e4boLmmQ4m2x8WQVWR6QhsHR6K8G4EpVHU9K1s0pQVr
BZDVbOJVIESHMy4lNOnPQBo9nx/mJ1WPz87VJeL7OD8bN1dmFf5WldCGsfjWonLEneBuomD8j92c
+HV4I0OWCBKEUlThXeCxd8rbpmD+jKBHHUXv1gUxFyB0GCvbY8K1rFTfZ7pcBx87afgpJq6yx0u1
XmQtiK1mwgUOTBViSxZJbnGRsefZXYDq8RisMf12irfY7kC1GK643BNj3Jb8Nz8uuSwk/9lO0YTq
/oeYL48aOPp3MaGhaLGcGEmLnMeh6oh/iG2e7rOFLEDTCKwycBeYVbNzWixDh0KvVs9FWKIkyRNe
z3h0MZF/rgRdy05Ve2E6GLynzoBdC1cX2Vfz5m7pSRm2opNpp213Dmkj0wfUuNEM5jIlloSDeYBI
8j54mhxJeJlRcFtimBAU/MlYuA8p91fbw0uMkvvzUVprzJnlfC8d4FqIvL1UDIkwJor2E94CRKqq
nBL/h/PgnGrrreBT9UF4E/25D2UTHXF9jA+Xghb5w7SOrIbYN0KSPylo/mPiA/jQRJygFA2Yu6k1
MwKxEfrsmTiGqAgBNHeDPxflpI5qUrtLulrtcVVhRZr+OdETy/GhYBTrsb6isZpAmEX/UgUzHAC6
RZRRFcN3EIV49Wj1P9uivDFL24tcCwnZnUNqEXsA5uBMJfXxkCoL6TUVe8I5KD7tZ3jPd1KDqlte
QtHwET8ugiy2eAjEq8R23Ip/AHUY9H0NUDFvcSGPz6PIJolUOlpG4eVrfTc2rItfT2NdGrWiOfgE
7y3gjodNdZkjst/+r2onZWbVHM1PUpEAIdaTOTBKyFHti3UJlQJkfkfEW6e97+57jLDItbfxcUJq
TfoEPvZBXdv5at4griS0f4Bee2zP2YgifByrPwW286Ovi8VvihWD+CNjcw57zU1uFHLYALShSFHv
i8wFzhFm4Yn6vasJcppP2R2kw1gUndDCKiRL1Vi4EFAlTpgAVRQte61Ipjag+ckANsbGLfUzqge8
ZdSdyOQWRrOLdVTHnUiPYnRIh/6YqJmvFBTHs4IrPREu6+qLvm1c0W6FEgZEvXh4hlU4OekoD/od
M/k0QdiYP+sx7gguGymskaHVa0T1hr/DoxTMbF66IaQg0B2Eu8YXJ2rJ/ULoR5A/oU/Fx7jWENyI
mJn9TYLNdlcCWVUCgNzPsK/13dP0Uymxbqr0Wa5XMIFFa2ZiWWiDR2Xw0tyjSZPoBb9pNmfM6ErF
oOSdvWM6ICWGk+SXim+7ewDXC5J1Av6G7WS2GeEmUqVe7nOyP97YqI8OlcRFSgvmYoP9RWjxc86S
6ul+5gU1aaA5O+JSKGD3qghBCL57zScTxnCIrIWhMZh96mi5NcW5I24s2B6Fjfr55nwEI/DeBLI4
g/QP+RUqKcIKPwbFLxT8w+nskfE/DoQXxZNjvxHbhYrgi04IRXQdevl2wD0dBVBAhA3OFs9yArDd
vo04t4ks51HtPtCC5tDnX101V3ab9EbN5sWdIGBDG7tA51ltQVi9e8CUwgqGI6uPKEukiO08KeGx
zgKnCVKBbdn2UnqJNeqWDcYX4OiPiu91mBuXSzfbwA0gXW7I5cSiE7Ds0m+58Fq6v9vtpSIzkOHh
2+l4qBtfDigCtY/e+V32FKIiFbL/cgDfKkcaA5Ri9oetSIAVQTdYy8W/7SeJeOXYZdsy54YhnyHf
f+kjgY4jY1it3mg0hQXaKsVwqxOCpKnr8GZbdY0RlBFGCxfjB22ho3bdnzYRlERIV2sQh93jevug
fHR1qFQQCRJK0AoGbnf4wUEVVHQ3QxVIH4B6sMwlePcnuD8vojte0uGPRhns3/uEVF2bj765qWvs
HxTDWRLXGvIJhBQp7szhL2k6AE4bT9SE4hqZavI/69/Dg1mwKGq0sn4dWbTgkU5f07eUGmvzxOLD
v0ZM8zekcL5ElHNa1hNSnliE0cSMZp3tSSnQYMkpWxIeyS9eGe44FwJ8RTPa1Kbct8F1rVZEMVkx
JS2WBu1VM7FVWjL0MrKqUtCkS7EF818dz/OaDTr+VDF2bJVKUinAo7M0mD2zOma1dbK2FB4LcKmI
8ZcBOdD/hGg59EIfwQGubuDbNlWOT3/keeWBlhghoht1l9AJNNcTnWIvRmd3kPpr8ATJlR257ExP
fbYSCDOhG/6locXjeg8YVCyRSeaVQxc+ygWpM3nSJS7/+B+SOjn+1o8XDkGx48pQo4cT0Fw3TqC+
Lz6FyDBnNf/bWrHE15CGW7D52p7iRDaKODe2oeWF0boseT2NtPlkRUn/TIcks8KzlUeexPfk027W
MuLGPNLOnrhA0qxNShqEkwl5VILv+WAAB/EWrjpMD4oFZOiTn0bZJg7euF384F5ji0t+JWFKURty
rPVRWO5GGfRmYW9JuNj9zGD8Jd4tgCPIHqmMiAnhauuYDCpANKFfsCeEFFUldWJUmJfksOGN9Vib
RVPzbL8NcQz4OyEuCqSqq3BWVureacPJxLxbSXMGLJIwCTYOQVUXZ5PSfV3YDOrDp/rSjo6l+/mX
zXk6PVVzN5Bsl5JVcho+NGr8Hik6e8T8uzn9d2JOCvE8Fydmis3zR6UmQ99zgb8V2TNk11Tau2fg
ZhYKxtQipgK8kjNx1wUlxfttJHPlY2fpT2AogD4niWBBf3A6fcXpmtVf3wmztFoEdUMH/kaJf2D5
uCHWnTy4OFR15DzcO98kV1NZa08gcOudVJfDYuxREWTjv9xSVylrRTyVMb1x/3k6s1qwnO8F8Yue
Q073G+dHphLEau3jJznUrc3c9MT8lhY1Ds0LUVkBt9288Wly7DDDUrQuDLCN1i/kmyJY5c+fxbfZ
2N+mff+HO/+7MTBHUt9HaefRKojHlwkXDD7Zfzls8/AECKEgSSOiGPc2hb03X2xIe2xYWNhGZKDo
qAwJfF+M2p81gGlsz8YKWnYmnigrREDqHjC7zDf2+oUa6IfrAEc81Nsez+yUIOfWOPC2J+EvS44M
uszy+aHMkhfBrVxL++5g+AL0kEdQ9EEql5OkZb31xofKONiNpWkAafJk62bs/C4eVCmr6cJeAbrF
Ih69tJaVwqaiV8UZLaHDPDhq9PNF4Pvz8QWRGTswBkFWLm6LkFyulhdGMSeLga8xeelVwvOUODGl
lXJRgT/5e/wAnAjh+L0VShPy4ViKcDYowu6gaqscxT38b5iSqJa6kFUz6XGOuCZkMYj3rlSIv2Ua
CvbT9Y5hcd+LWXpuXuBtpGlWfh2kCyXIWDcWCPrfMFERhW+MiNNahrraQbBdzOTv+GKnm7ZHgEcL
g7rtf68Q7by//vQpXWRmtFIhXIe4E4ESBLXCUU+eS+qIrZcb5NLNaD+V7d6vuD3VUUg9DQuqiYmr
tM3WkpmGRYlBbUOSD6iqyX/UaAzPYQfjzqDmCISDuWr4rE8lm02FvJ+t+9hs0h0r7v+3jLzPfv86
B2u3FiLvokxK4KTnCAlF6Kd98HsxFSuNNxha3nIMEQYgkhqWiopCchZt1minVs4rEUNLTxP8DHSJ
T4TZpncAj6uqKrYOevKFJg25tfBkLG/jcT6WiBlHRP5Zi3zWWk41AJmxIu5IZGxzbHNKxcKm3Y83
7AVcEIkm3o9CZ1ETW+L5um3n2AhHKQZ5SHx2KjyAabotAYOgRxbcoaIEwb/IUOcN5dO6uiQwhVdK
NlbVuhtkW+jBNEiA7KCA7/0qeXMqSTy1oBVxYIZn86KPDaYYwSKhErHdWnq3meAxAxtLuv3SHOB1
x8MKpYpZKqrspimlIKkQWnjen0EAXh54wx9mUTkPjOZhG29oJpAC92yDYPfQCd/f3SY7uYtqJCsL
RD9sIdNpYGth63QxKhT36NbN2FH2DMSTavh3OQnpcOl4Z2ETLIZt/O7Bgl/DTkkVylnddDjUmttj
xRtr5pxo0ZBzPSXMcTu8kBCIgIYuA+QkLQEY9++ch49ZLvLmAHsgQNbJTUI7L0O0ahcb+W6yBVsk
kgrWcSW6PK/rXfdlKKFSpi5zGVwqoM1v2lwyDDoXxVCi3Rr/VNnI7qOwoPqM5bWOl91EYk1rsmWH
AMyvD0ceU6aQ4dgHwpoqb3TQGqiGvpD9lmY/RYSIl2OloLdS9/JM71D0aP+Osf16kTfsz57bmxrv
y+uu+ToHtZiTT+1Ug+aPhf6cVuf3xfFexER9fXP47wAWRZQiciGug/vUTIHLCFPBF0VwTbxedBVG
AC23DIdl4WqmXnqHyHhQDy1KhNOll63UAC3U33MragVTwNawP2oxxXzFN0B9q2DNSInlXQLvmlIi
/T+ebdlXH7jL+2lvcB8vs1ukwpz1Qv8kmH/IvJp+Q/J3/uYLcH9l0Up8sduezdywM0lhe/T3rriC
wz9mJig3lcLQzzYNioFzpr5pS+txadBrBwmUMStk3fEVeqDYxliTaimnHl8LwCxpHGInkHm5FP0y
1UkweiHkEkyrQoyOXl8Xb7L1GtI7xLn/Brietmlqf+hMUehMq6osv27uwxYmlbdCfDP3LoXINIyQ
Y9vVkgGVjfFy1oMmGGj9mVkIMzRoa1JV3/HjT2SwA5kO0ypcEFNlyQUhSjeqC1osvflVoUyC0zbj
daJvwlJJ1+gtXxkKLJPgkB+/nFcfI9wvu3x2i5OJx2mqUWdND6Wdcwgw4YN1qeRwklXRP4rt+hte
BK0rVYBIuep5XMoX3uUR6O7PB+Y42TGi6zVaMcTVF/KNP+3XFAzwJJyugyq7J/mFnajxjZpHugr+
bI1oMTo0abV5KW8jX9OVmjfyl4bIenWMjcOrnxYj1OD0m1dwz9kkfSqzLI1WXBxy3OFQoVmwZ8JP
XtXCctH0SM/4M/g84LYJx7Bbm2HTyw1EbRXvbz8s5ZgGiNE73nzXD4jnQfTyQfwBfCAClOShYQCh
wKh9O+uA7Dy7ZZeYD1tptyO6cSB378GfaGVY+qu/FU4TQ0IzSYU3RXkbygIsvSQ0uwF3wI75adqV
c3e7Yzpd59+7HftdMa+iAZZlZKv0wQbqKky6F5YjyEC6IcfSrtVZYvKTHIei8ELNJnCp29r9+3Kx
0YY54hkHTrck1Yi8FR8lDOu6SRj5thfJrnfqyTRr7lTkUtAjM76WOFevHfGqIXmnng0HYwpwnCVu
WwMwuXIRGfNEaqLOkwvKGuzdGWTvS22jjlQll9Um+pTO9HSYzl9E82kjNzJUNHTbUyVdChH0k03c
I96Vha6DA13IWTd1iOyvyWFwGIJCwtRr6DROWf2lCp6z2kdWC/XeUnjuHPF9s/FYXLCc4ly+O2xd
IV/GNJG8ltmwQBgHQyDPgNJg0SGGUwsFUSeXMInWOtXCOFXTuBErC4L87994BBKaXqYFHpYvyJa9
TA7laHGKB9AWlhnuktAU7Yu7t787lJtcTZfPfJeKWyR6D/aAbq8z4dPSk6hi4nUvZVdYM8xhkMIv
13mk22A4rjzGOmXH8oP+gdONmeK4msCI1l48yGNQ6cSL0aTszoRhkj+vzzvsj71S9mUEgNNuwhDI
Ru/Jesuv5kENkKvulud3DR6CfuDrQPlPU5hC7Fr6RGcauPXbooPrYRapupVrPNTH3wjHr9amQePg
IArj/wFrnm8PNhp0TJAdX3PTmR5Rs1zZonh9KMA0AQlbcaXHuoVYnjo7u0D5sdiP0h7/ymROO+Ii
y8TepDFLuam5fTP1khcJ9ftEURhuYgRoeEWlq3vvu4LGjD0rufUemnC0XcP0uu/+6uzYTAr5bUlu
MHDouX4+/gPVQ7qlhVS+rvlfFBaZhH7TyhdK5b+VtqkFF9x6RkMnGKxgP4Dh83douXbS79oKqshM
ek3FCG1uuWLcZMtQONzY0WXRs2sDRsS4q5CjourUaX4/Nuho0qf41dhODzMizCqL2KqoDbQp8h8r
e24xXBd6IuvPm6R66B5zWisMmA3c2iD3EDFGtHDw7Zo+opd6l0eeoRf5Q65Pw/hhLJoHenAJ3z3W
ttWZU290zN/DKRv378wWdvwsTZdZ1Wwg+I2PLNP8X9H+rceQLkoC99QyMLOXS9uUVoX1yOOX2JVF
Rad+2Ad38jKA1slC9vEIjQfIkqOE1dTBFoHN8lWXFqkLwPkZ7f+tiNU/ZSHCN2DSY5uMNbSOZScU
I/7qFjt5f8XUBJY+Db9a5hVzEaKFvcTGT1Tw+U6Ex7Hxiy0CdItcTZY5qvbHKriSQuC+oGqPzOSY
kBSljoPYoZPS4tM23xm4YCstp6lOvM2q0F8VUDCjSCTouSMGkoTuv7T2k17ctZAfpHvzyUIlmpUd
Y1b5HO7ZXXbdOg1pYmIvPMPBKfdpw9KwtZnOOl1BUvRy3S6N6ccwk2zO2N7W4vwSR/BIn2DH7qdZ
kPtQVMiRLgXLP3Wxop1TbTjQltqmZ17s9K2rZ9+3TR8I1v8fvvcGhyHyqbhKmW5V6dpSrUlJdSNR
ZOvK7e1PakWZyczBt0UmCwLUmhgt79xLTskBhd/G8SaktKWw5aN6pqdwFxiLMr8mBA+dwDacvla/
iHP1Y3raQVPgcBUqeOphEcV8x2VZ9gKT0Q3Y1Yit8emlGNaTAzHz/QrybajFiLzPQY8w8DyVkIlc
S2V0Lc0RPiRJNSJE9lKz8Z4xaspsUtQpcWFmahkOP+jeOAnu45qRp2IR89EWSuVga0L+qqyNbBWO
6wYcsZOT7tmLaR/rG656H4E3al4Uou6PIFTX4EQv6xLLGh+ZQcGWsen4Amm1uxIeMJY8lsg12lzt
lb7TQsH9hQSv0s2wnQz/kOtqVVbKPdIl3bkgVF3FtImmAx4z1had6ksP6UwB47MGzZEpiJ6TkT4R
YclOf9PX9Dfdbt/fJ+eVSAbF94JmFwVs/9sh5U8/6Un0X5ykuqPSbjqtm5zeVJqW3W6IutWQstHV
nUSiGyWYOzE/TmdvYgB7/i5AkZR2zvK03SJWMXJSWtPRLZP/lQJKGmklZqjhyTrapWuAGSZca/8w
KI1bCzl2hZFAA3nsv8uO2uuSOFcEQYGhcVXZRL0p5arY675NdjsQP8r5kxQ6swJUzdKkNzhxOuRk
MFh0OtJBER4hsfz6C9sE61ClNvjC2OxgQ52ltn6GZgP4jsWiSbvKTSQ+1sXlHdE/uVySvB8dIm8C
ljKkgXMeNG695PIiL4yuVJZLuan/Z+xpgem3QeSAK/PpbR/ss+qiNW1Rzuw/dBGTTVpYxpePqpNs
6zkkHc/wLV3349Q7REHffKvGCrxPBuJM2Y2QJW53EzBmY7CM2QKs62iM6TxixLBkYVGCJu8leozj
dxN41QXGLT+hQrY0Ldkjc1EIXvc/VIkVpRpLnbU1TQwZUkM5GiEkPVUlo0gzn7u5rbwmb7CjJ7lt
MSi+Z4JRFkFq2LKQSHc1yysrfjoSZ+83dlIbprzMR0Rz3dCzx6lglcjD+5hopyPDxylDYstG0c8y
Z3CvbeqrZsncKC9+tUQwQDuAEE/szGptkyR8jWYAbHhTzYd/NZM+wMjAiSy8cDgSDjwe+t7d619Q
8WxE0rK/rzbgO7eX3ylMBuG1cxxwX+eWRYqVjgvCHlDKtv3mevH3mFm8IaF7+9Kldw+zgxy1LSM6
IXzffQby37zNymQ69aVxunSJyTxPCp7Iv/DSg2y4IhxCIqUGB9+Cmt5LHvFzipaHbsukRD2luW3t
mI+V2/lQp1pcguSEHrfV4bbELR/PFV+UnJmhLzoSP+R6UXnmZorDGGw/oRwHRuWuViYQ7NVaSH64
MOaFAf4nvxfNyLk9epohRUXZMqN0SCghWRUdPE6Su6Z8iboHkJ3EmqPAB2lWoxfnMPV8icac079U
Keo/OctYqLcx/8Cabi0ZNKqY33ElZDTRzwO0oZZ9Ne56/5uGsDrXgTv1vwVFt0ywxDap/DFOc+G+
fRn4OGakXf/y7CemVoGiK/b/TFLDBXvaX9AHkuFEoAlS8A8pxt/JoKOtQJO+UMpd1qqH4mdaB4nB
rTw8EhSiN5DfHr6qdwK8Dy6dn2r+RSDSQd0p06WXm2Zj3E+ILtgdtEb3Acsf3vBb5hN4Lz/AqRb8
QRmppc+wMWXloTvtnhG92mp3XDA0g75W0GlJVfb+WkntFJBIkjQxCv2cbDWpx76ILFaaD+bj1wGE
f7oJnSMIfFHN1rLrIR6GpWqTpOf2jspRmYAv6pcGVLHpiZ7HvtYI/oeQmswFj1w3xnKoo3V1NDLu
GQ8cfT2hhiJ1UyuBoMisbwMDaI2M/e3L5YJ5q70hZ3dx9kpkoXhw1kaI4YuuvfoLW+K2Wr/QdtUY
JHUX4JhP3fGDlhFAtlFn+j7yAlAOE+u4hHsNfzMU9Fd4urhXULTpfN+6tyu6AEIT5oDgM0P0GR7O
XqL0P/JGdVfVkmigfOyFXgiBse+L+iKODe1+OLhZ+G01A/yWEcOV4Qh4QGickNPkwVqE6VAoJOaD
2UZQawrxPhd1xUuDTei4LF7tnNfW5FXa/t0Q3wLavMjHyoepOGR9u/Pi6IMyOg8y+lUjRfSbBHGF
itT085JBJBW/SI+QdDW9vxioKuLon4/KiA3BJE8EtuhTgwotIpF0RcEhcQf89hwlKAcMNizl1e8c
nFU6snw/oUmJlU3BpVMYiHdX997LwYsIeO2tY0ctV1jqFbqoVNIHj4H0o/7zqPlnU6YH0MhZF3GB
qIubBL8xxA5Jl7fhKPaQm2jRxmIYOeUtC3F+wlC+A13YUHw+ErJf+O7P+IqBhq7h0b4c4N6+Dww3
ReTKqJckTQ2+zYpLYPTRUgHP+25+YQc9B8lTXWwCZjpGd0gUuMS/yO8EU8+lKVBwiZSo/XseeEnD
IpqJ5xFAcQ+VZmjqzaTu9wgzI/o+QflAo0FjmQ/PnzTZ0Udqej6t2Ow1MIXY+F1ExEKr3+M4/5MO
ph7P0unhrDKkAm0+efqY+XWyXRK4dzX5DOd281mvIJ3GvS77ZMzICcYWSJY4mhihSXvenosYGtKT
1J01hMQbQFAgzpPVOGIZeo7HZs3D1BOSMLw7J2/MMgAvjPjkrqMTB5eWV8gjwU5i6AqGZgWINLju
RD/CIpzQJYAlwsAADxFb/jd0s7MJLTCPycfLCeuuUfdSmbS6h3cE8Tg8IE2+73jFRHJ1TMdDEp8D
cUIPAmJgRozPaQ2l+y+OR900nsPmHzGLhKASGuMGp2vHMLGH8N7t77JX3nhwamIhehvFvC9NYJ5H
VbkoSRucTwasjEa9CJdddnntrFCCfXAgx5NY2is47kr6Umz0q2efx6g1ViUel7t5KYQ42hNfQI8x
dWXEjbUQtdycTxtUELde04KQRzj/LbHgSHJsz1yHxDQ04zn5i5mpilrX3NSfBWo01WWt5m6oz/m0
6EdyNpSfQUgCibJ80TPU3o9AW3FWg9317+IQnHGOa+cnervVV/vsxZq+6/ueZ8Bq3OwzCe4PvIeu
1vBcVIoeQz3zuJadu0Y3Y96DhWX17t+X8uVDLEfkcIEb183kwIl+wP9tuWyHkCLCMf69BJ3a8aR/
lJwcE4oTniQEa6G/fsG6CdI7o2csR+cj1A87iQLGyN3ryhXjrK0EMRxGND6ufGR+n9/YAd/QPgsS
RzR6DeNhX3XAsGSUwzNZQKZyZ3k2EXJYbemc08uMqEOo6OM/Yt3UmaxzzCxyyjPrUcpRu7GSMKxm
ckTBNtw+iacM2wC7Jf2Pu3dN3vuT/9jsmkPbEE49y+Cwhx5m8V+0kEGm4al+f/rGZe0iOqUT+dK5
90QvNB3xTiIQkJeSork6Q8lfvpiyim5RfWmM+yv8e85QcVUOPfyh/wwjeWu8NQDSNdAy5I3EmIQm
Z+BfDaV1GdeEoD8a9AYQwNOfkAXiMLH7dPzaXz7Gv0EOc5lnPv0yzsckdmPmBS5j91lprVgHOQRd
S0rddoUzq50xnQHETzwxN6PvFm22B7wKtGj5VGQXrcIZNo0i+9YHlim/v4tteKHktYaD8vJ2lV8a
kis9O23r+3brfNR4gLSYvVzyUKMfjf7NaFux53KNUyvnpoK8d3n2S6HFvAwABtUiFe3rNWi/auV1
aMBpC6EhUd0SXPIwXgH9slCrG1mFdLIf0/Pq4HZyLJoEHFeENbbM2lco30/xjzoOQrJytgZx+Ccf
MeCp4XKdD81aXWCMfckeBnDzXCa8u/+QtfTucO/qwEhdr6oLU7v47j33AG471roc3YN5rCH/iKJo
xSsFDrUBhO1qzYb1auxcGIeoa3Ef/EaaLs0ARgm/gSDK44OFWOpM5G0hAsDUTI5JOVSgt11d7mLM
GG3+TVy5qvWMDvVbk+Z3qBCepEyaEUNG8j4oa78r3bym10GUZq+e4ny/7/r3zTEz8r2UY13mAuTV
ycU8HcMNuJKA2d78URtKFB1e910xMeSEHLl9uD6FBJ9e7ucG6yln3DvOGpAUsbwdvVY4EH7H6Pgc
0Uh5mnWdoyeOVWYyBzc1JgQHlqXkqhtkrmPUs7hPBzTas9TsnifY70K6eKwvMaQmh10W0EB1lfPU
eJjzTcKPJKOQNpEkmOnHpqwjvC1oQCmKgBL+7txhwJZtd5i4zLeLlUcaHkZTCFizeO86sNAWUUN8
5Je3CRL+6AswLoojSB4nScnKwfsJZzuDFHXPRBLVQ0ayjHheu8eUdvy56rtC+LP86tSj9JesXz4I
WRfytwpm4u8fj4+pRA9k9Q1bSjP9KFGBWDVCk104iaT9RPTWqNcZxfFRpzsJmcH3I4FnTUg4vNt2
b14T3g1B/aWqOa4eKI3IBwWAW71NpNUgV0WI9mQlxQcN51Gidw85xBfiOTFyTOY1XmnIRv40HuAZ
sC/0I6YI8OM0kW5PdWWoy2qv1nOJGPccVJnbfJSLFL0KQLqnpXWpSpYUKLO6h9SK88cyDbWO7khn
TxFQmpbmPBiwhHqWqTOzVdxnDAqCD1D0UwrWct3dsPOy3FW96dINY1TVWG+ZuCVv7HdoPMLd7qqm
3CcZ06wOCTyuwkdyspp52vnrQwRDz96xSXhkRuIi6yCdofwLrkf6LwXH28igq/CYfqQP+QSJw7rU
rBc3DxFFrrxa7pECVNvYq1gkRejYDTwebpxbm28z/Ng3rikuB3jsz/LOCLVW33xYP8PGwxNKJuPO
erLuusm9jpS7RcbF9a9nKFxwKctZwtO9XKNKWpUyr6AtAI8sRfTxvIGZFn505nRyxsGhwfP5d3qb
aTcrANsg2ZssMgzulXyxEwguI19ZglY9hjnUxK/c8N3TFc0PqbKTz2I6/9eHDyktaoAhVMlgwEwW
p1G5GR3H176irO9GBNSVOaXbfKrzzcrWZ2AxPWImvgZYuYIl9l7oQc2RwWTfTs2Vc2VAca+zrVQl
9T51nVsn0WyDzVGKoGqCZvBGUAwROvpF86DVJD4lmF8iOpDZ3k/+34plIVmM1pR012GhP+mOsa6f
Sj1VvinbbUKW8OhuearUdoZE6IG41NHlqVLpbyJZ4VQQC4OLdWIPbY6oOtDmapRJEMtj4U2njU1V
WPqEtY8YJ/kyTya5aTmH8vIHJdqAxb42HB/mKLBH0iECaSFsFkkwSI0vewYLhIl90LwICjHwOx+w
Sw6qcCl4K97yHoDShocHGYuq9sx5LUDytVRy18K2FqGi0vDNg8rFPPRiw5Ytffg3HaN8WB/EnpG7
8SD3ZHfcdsTtUhJeiAE44/28adt3kYcldtLjqGPh5lVsqkLbcdUt5tIT4VGmRUScq/e+Y1N7cWXn
4IJxppSkIcq9APOCAk8YyAmDOJwXzsGq5lSS8+iHGQUUaTHlOHBR7GITlKH7xAiXc9JcvpOi31Wk
GSnWdnY790N+Q8K5lvVOoD+LnhpYAM3I5iqhYKKGvmJsuAi3pPUkyPIjMZkab/i7WSTdVhL/Ati7
aWZZVd6n8WReV8XDlWgY6df0t4nKw4vZFz/fTrgDhbaUExbjCD8jVgfUIbQRa19DLftV0JWDd1Cy
7Pou4VGqYT9ME7jAzN6q4iZ/qBX3IcOriQjrg1JHkeUrUIcx9uzAhtspXXc4kuyHHPcVZPdDJQeb
wDJYe76UtlvLwWwWDtiTvow3qdnOwJk56+y5dD8x/+qA6Vcohk8HhBompb0N9UF5ke32A4OshIzz
QouF6wl1VotXE8FhdvQZLhzJqFYg2uaf5rwmOLNaRtRcYaxsy+/Faa8t+JvAjUbiXuvcxGZeO757
O4l++ldFar/Z1hsLq81bz4njLuo0VsLkcw+5TIBldd3J9CH0EBi+OiupPMKp3KkF/DSOcq35Rgto
joDSQ58oym2z7FhzQu5xPWdmOhtYod3Gt8U2dyw8M8XUa4JYtcQfFmQ54M/+D41+kRRT23s9AfJ9
dDKbp5pCLo7bQSOHHERZDuZBtQ4VZch7Rlth/tCqZsL3LgZK9fu0zmeNIU7Y0jlcwbXyUffK25oR
xK+2DluLOH1MZnjh46k/he8WQMsdPbXYlSs/yZhKXKNKLaxQjzT1lkMAm9c3ijBifyTceYKT9RJW
2wj4qZInRA5eGL+fpg3n7Bm7D1uBOC3kgO9NXaS5QR43tXx3gjMBlCfpeSMi9pYjvC+4vTkPt87F
79WolItXQ4u7wQWRmkdVsXgm7jhguNO80xeaO7jMg7pWsmITCXlRsO08gNXjy04zuIhw7xtX6bkC
gwJQ77JOAxtIuQWzjWLFEmBVQJxPmlgBe6TaJ2tBzapwggIe7dNZKFGjPjccmJzlLXHGG+PBsS8h
XX3kVwMToBLTqyLnDO1FzBcj5XreRChIqWF+Ks4mCd7kM0MKsAeTSEpqJmX/UniF9jkZMiIm7Dnf
lXWtDvOvnfJi1y8y1KeAIC8PtKaCfhmKGCvAo7JqgJogN6mss70L+XYiezMQOnxUPn7jyjDmyQGR
JszNzggH8ZlFsX+yX1sXnT8qxsaJl6xxyOXobpL9uglV/ayJGCekkVuwRWpLhoKmDjeKBdOTRb9h
rxJ1sPmA1TJtHbpHQPw+QzTTi5GyjcBmczvWE1Ua2y1CGGVWYTZpYsJkb8mFMDyiDAdDFcS1nQ1B
oLg82h51XHprpKa32WWMYFuw2toMp3dWhzjm0vkKVKie68X9L5m6gYShM4LCGv1UUQaavS7qMJs5
3wzb9KeEdLHYCieBdGLVw/vfS7+SkUyTqpyjWuym0yvFdSEZEvvy/NXWpO+ASKvEktcaEQyoIC4c
eQehAM3SVpLGLvHOhzsnH2J35OFtfQjNzsJGNjavxjyQ3O+qnzcRIl8uEJkZWkpEFHbTn3rdFSPO
D6gu2efnMp6Y//weOQcwIdr3VZyC2Rgl0Z2sXPfrpE2ZpVkgAUbTpnjWhu97WvUrhqBKn8kBNAWv
CBuEjDSAeuK0nYG6BYOJU4EhL3jRRwbEHRji7mexJyra0Uvf2uwwF8Fgp302XAPyYA2qAZNzlsO7
qdZ5aJLcf9xNqLshuUeCd3wsfVDwNOMgXHTdiJYWbYmuVDXWzar453AX0j+vhCCs6cG2CXFQNlm2
j5oVXEz1vbwVGenY2GsIyp1l2QuN8P0lFTQndqMXwlDeEstJXRiAuoRgh3PYmJj1p7ZmU8Qukvm1
VsLxhS5vaf+BkNvJUwTu04p/Wyj2hTTTgIji+LFNyZJKsp2sl7QngoRa2+fUGZ90jMth1i96Yl2M
MPz4Yh4GYYPxeZE5rDE1GcxZlKw7C7RPTiPWOECCZ5KIAiu8spxw2CePIRLCeNqFEOHthsDIcM3M
M3DugRzj0bE42LavyunCveH6qZdrrbMh/SZq3L/XuyM89a0Vta2aSt11shjndnmhG/dEgeCBnfnR
Ub+URMRZroVYq5vgj9YFlWci++ThXcUCHu/J43zru4DFghUblVO4/enl1Tcfy5LdUmQJGxA/+4a5
gfeU7MfQEn7CfE/T5anawGBUnOa4/pSM/NRZ7Q9RfaGazD2CygkYc1OIDpItl+Te+HzXMZJgZpTJ
+PVT1wlCdCOReVTuG2e+FNekfnxoQwD7O2HCkajR1Eh4chmD0VpewFr20XuzxG72z3b0eeNy2Z5D
W9pjiGhzdaifa3yw113a+H9jFIzoPyYbEfRz32zHumiBHrCiiY2mUhGLSuQEEMgvBDzOpGLaIfle
LnR/IVvmXf6eBO9Pkq5W52onad5r6b22L9uniyMIvNOlF5qRCuuhL2+zQZWFihaSjASmQlMi12GC
d6sbBHHQ13gAQthNaVTIHSsQ/oDpDTQjI5lUoJjsz7vpE8UIpwk8WcqZJz0DUyiQ3PK8N4Ly7/ib
1hufV0SMzQgnmbVkPH8EvX0ArI5U4xw19je6o150ArmIH8SfrF33kYauk0UF4HqX421nruTR4XYT
dDgX/xrHfNCLfM1/X5/tgh8DpynngTFE3opDY9qIQwLBtZug4bYzZ3NMEaqGjz7Ezv3vVTC6QZCL
9x14cF6RMe5E30KvaWq7wvbdFGYSQXLzg+HQBssiF9OvKiRG1RRgfRVhpfFameS/0vGTcI7VdT73
FEwDwzFeAF/QsRX1R+jz0mnkCdB+5egkhxT4wA+GjreI6rrTL+acTcp6J4Bl90pkmw8BwUWXoedz
RVo2K1sJxwX8k9YkEMVuqZKCLN53SLBbTq1nHfJqrMd7vA4SttH+8Fd72cMRX1CBpQIYLTeXC31p
6DoiseowbrtPTo8soxEFtNCF11+Vo19TkwghkqZUPsg4UnzezP91cmGngeEZrwqBKAJ+EAyUkjM1
Dhg3qQvosdJ4MiitE1MRDuxwEQtq+2c+875WhxIWX9+xjOtf+c6i8ywaoBw6O723bY3iA5+j8ID0
4TsG0QUxOFBRvV57jDi063hZXzq6E+tI1FP/9ZOE0ral1kE7VyhmYHhhgZRuZCHmjwZOdiI6ru9X
SOS8pzKlVcFdmxDldX00PlxitNFwepc1w+PqM4vKeX6BVDVDw/mZbFT0N2nQVfjqRWCNhM0Y7g7z
exW/oxH0D5Rvf7tq//RZAu6BdMBCeM2YZ40JC3LIgq9clUTs8KP1DCnWG/XGIMjCmZrWxjbIbOc5
Qrvsumn9MlCi68L7rdCkST+AL9sIwW+hHvCN6v0XTcek8MZTTBDxIf0Ugno8qF1ad1Zdf2aGih19
pkn99vs/NRuvdEs8BtcT+qhIsAOpOtpQ7B3ndm69/2HCuD0jLz/Tr+oP969NmjED1nyWi3XXngLR
Qij+THTD+hMb0geG0BpY5I124ixG52mBpM5ny9++2L9JlKPDLsGPlQX1xS27fqSfMT6+scrE1QH4
SKhvB98UEevMujUNSPOyDHCCSez3mEL57v+Koo8W12BLQATaUfcqug+mxPbca2KjoCsR2vHb5uyr
IMYtU7u776QjGFkFBxsej9ttr7X+LR9nahzV6iNY7xWOF3FMMWS7TuHpxMRmrLk1XNLBpAp1iEqg
BNA19fpxgwB/gyeye1CHMIVx0JY5ItcATgbeAecisMu97frnWJR4A7K8cSvj+MhMcDgj/PMlhUG2
HFM4UbarF7IYwAG3MTkU7z209b1GCFg/tAGIAgFInfGFPru0rIx/TIM0S/dAT+6c/JiB3dqDrjgR
3DuldmXZPwCUT3cs5LnDhx3wPqyF1vw6slFZwUBT/7LhB7X+Sv4AL03H/H8q9lzvkhuzPX8gWJyb
0tcdtQJaELUsQeDXaoS0fRVp0P68Z1zmPGFKRdzug3MJYFKtSvS1915V/puXl6WEw5Kw71kFveqQ
OWlxC77ZPLcJ4eaqfkZL0+QS7MEYvziLjPFKYkxRpP44Rc5Gq4SSwqtUAn69X4ulfNR7R7XEzdqe
tVrGH1bQxLaYHttgN5DPS71Gh93+0ySKguuhdyAbNwnwRVWwyS1gXpPSblZFPBWaopGzb+mk/r02
ikxJJ/rw1ET2kJyRm7BMSE21gCgOiLhrL62w5rl2Tm5hBd5Ldrp0THsRh07w+akZkaG0KaFwSnTT
Rk2F/I5rohOkC+L9tLoEKdX66LmHlJrzphERj5nklJJBycWAz0zMz+N4kk0Y6B1z6/avmlC/RZHB
lnqVC4mYIO4nN1BEV3gHTU421PQBO4URwKvHsaTpHmYijPJiCUxBwMaFPj/1drxe+BYOA1S5z67K
CXTXqngjI3ymcDaRB0PSC6DJFGJA4giU6k2mRobusQMEoiu47Py02IxVP1sDXxLAeHeIqxl24SvZ
37a55b6r9u/FI1tKOCVD1Yue0mep4zLBlV2322RRcLBwwkP66lA2o7iLx/XpWlAUA1iAPZBZUERq
KsJI0DgpRte32mSRCirSXwRUBweuVZZC9FeUepPoQoMG3G3DK9x4t3heyQ0DqnrX3r1I6oJV4avq
1Tld6pszUFVlnTg5y+m1kwk/68HneyGYr4Yr12Cn+U8ABzDyT+30C3tEhHThx2D7B82Jn8s7aUzv
dGy6e0jqKGEsB81UDie18MX3R9XQRDPijFM0/2fRLLigA4eDe2fdewyQ5Axej6yi1ZUh+P1ryHy1
3lqk354p0ujYwfSkY/yK7GyslX3VS55CvWLt56E/ISRhEiFeRTplM+WYGJvZKHVUXzkvIia6dVRh
QFyMJJx2CDOzmAeeoIrYHIeOtQdZHDE1FushoFYD12qLi+N58DI5M/LjOaxBWPASttC7Huq2GfuD
0NhoPLz6u9vV+PQ9pVByjpEvI9hFeEpbRUhV5p/6jp2dyBfwT4O4WivYVZLcuCSf6JXTOevLxo/j
kDjouMHcWhCWzpqNSWf5i+7zB9c5c3wf4t+r84NMDAxmUjhhYEjgB6dvqqCl5CD/SHXmVZzyRojW
xeLJvj3zXS2QyV6sgarG/fqmUg/0ijzmmPwvKpRi4T7TtTkK7cDPDdBk/IbUZ8tWM9slSeGL/0Fv
ikBZAhM6cJEoZyxlhsS26Q1Fu0ixghklcT+SDao+AOq45sWVOuWGJa1o/w5GE5407tY1ttDKV7Na
W44YKAoiDYKb6Ceb/2kr63HAtk10uR7pqNOHF1P7ZdyZ2aBIblRisYephaGjkuMgF7yhX1BS461G
jkHQ/p4+6Rl5mkCTvYqcLQ1QojjJKi86JaZAbpwjXqepa+Ir1de6e2pGiq5KICDJjbCu0PqQbzHs
p31yJE7ctVML9MhMS6RqF95EXxqdQkrQJZWMM+7zy/3TGb893f5QzTUt4itKGB1axlop3wafx4B7
+ZIEOXGm43zQCVqAElm99mwzxOg4IeNMLVsSp2MhVmF00kTORmktmVv2Ohvpz0sxgYlHRXMVQp3N
u7NR6bwFgGdwqzrDhTPRt5BsiUrYKTu+iInrx0liOl7s9wFMv/+OMABQenoa4sn/JJcuIjyfQrr/
3BcR03I/AKeF7aY1HOPYnbP+ZFCVwQ7ipq+pgPautjC2y4Y5TxwwKURsYQ7D1hwd0TrzAd+vy2fi
H2/o4FLzdUf9UlKEk1tZOjPYIdXOdgP9PTjoycKRqLW4ekTIkEL/2w/vpCKzw/lQNo9Ax8dr0v/N
3wt3jA41wxivWCHGwwuCy4uuDbYkHotLAzRBgZMihvfjVqusUW++81sRDJfPNSHuiAdRMYQKUQff
NYF8147Y2qKlOinnbcm30kdKCR9x6TbvvM4+vsqUPdV5wXVMWTB/Jh6uHvC2xKuiso/D+hAVWA7V
oCon2HXdqFedyYHWBVOIogzwaWiHVAVM1c6X96CChj+xygjDkMJn3fjOpVog6nHDww/ZvO5PChMp
WadlPEF/wmZzARBagrPfbeTBhPQbg7dnqY9wWokgUWzf8lW67if3zaQ4w42xdPzObrmyVFXUgYNx
qGqLQM8IfWlJBdsBbJKzuYf/oO91Ro/Il0Vy1//wFQxBS936+RKggXq5sEBTT9L3otKJzkHzitms
Y69UizLnC3gW7P43oH+cIioHwrfweEjxh3fsuKzDi3vF9sJFp4hmrHa8z8mP6cam55yThJNUZBru
sGQ6R4AhQEUMqwUG8I/D8qCJGSrcMWIu9kdAq/6K27OyKH7+I4PPyF08rzf3ti7FTTaqPkj+4zTf
yJcPG6It4dQw5VH1HmLSdXwqCm7thmzQQhZTEXudHK4pDcdjSAcBQ8nF4H3H3BP5A2d99ICRYamM
eAWEOmcVamceeiVz360+49unFA/r8X+GKHR8WeuqSBBaduHWFRWqvTsKb6i4gSKznFDQlfHY2oO5
foSpuZoOve0ZUxNup/YnwEM12WKd6IgauhK9fZ7Bw9kLmowwM9ggRpuKSalri72bmQtH7rGwZdNt
7wVw16R7wLfAsmrNoiHtQ5NrfI8DafnHT7snU7ueq1KKw1tzM3OS9TbsbtyzaM8mmlIL+B7ITU0v
7sNCTrsaK89eG4NNrjaEMMbPXg5zf0dhL2nIv+tCpH7GeLOU99bY1j4cr/sgaVOUk1E98wk/B/D+
hIHz4/iBscykFx9YH3eLouzKEly8TooCF0tAKmXg88d6TLV75wzjfozlpUt60COjZRwSZFqHJM42
ONXvBKMA+HLZM/y18sXzaMrCI03G813CqDbM9OzNewOTawIRf5aG3pFHDEFqzlln0NuuY/aviG3F
cfJb3CE70xab/gyzcEQedVuYUFNs1KSdNXnH0CXzeg4Xyp6l1lxe4LDjYu5MvR0P0gLL5t9y5IHb
xhxuiBwrolOEo7eqwe+GynbfLNh2DscSx8nTqT2n0yzEyFb2yOHX960hpZ3qyrXCnL3s8pui7RGU
ibfTH1OUNn7lbVfIZhoJTQyw95jCsmt3mNf/Gk0wANx8Vjsd82UkUixSOshkDLREoZU6X2aXgK/x
OcVdOcO6qBonGL/JDH8TwwdKKG6/z9dbDsGbT9z/gpEv2qU4mi3V93mJ6MNokQY6+SyvSFpoFwVe
f/QfZ697lJh2ID41D9TvluxJrGaH6gGT3PNJ5wyTYSYGKnDVX3qEUQr+WH0RCzGi4YCCIfN7fvgQ
J1fR64esPjucX8X2e/wj3Bg0JH3DiqR8/s9rJ/B5AblCepSObd/st8xXj+jStbHtw7Ja10ISz7P6
VB2yTsMz5BucvD6+DAKLGWsVtJr86NzaCFjnhYRENlY/RVacNq6sBzsOaWlD0OnK2MHdW1gRAvU4
ap/qvlWkTBs0iBOlGhK91XNZJ21h4cfeMvwQi7CUMOxZc3rZQ62jNt7H8E3oVtxSowpVLsJnkbp5
tLNqjGp1jg11OEIWrx/WmT+LO3gbw58Pwg7HcvodMR/6s8lSI7ren9PuocbCba4NgDYVFvflOqqI
rCBv8Ch5vJmorZyPCMsimrgcTr24Lt5dafyCms2qKvzGFWd4ThNbKl9hjbL+raRlpSAGLWnmeP7D
JGCBC8QP9Jc+pYEjewC9nq+JYgrXAobsZ7zINzRATYGwk0E8sQ8V2KGCe5sbx039UaQsgQzIMfSm
f3hq4gtcf8x4M6HNNopGjhhaL0Iuf+gvtMg/cg0UPyk/8giqQo0snYmTQP2Eo/VF7lqTaMZeClHi
6SI8hsz/zSfb86BNLJtSAHRtaAjfwDaepkC0BB71vwMXafTbyqjETY7sNs0F6nmmhDrXk6xwi+oJ
q8X1BtE54fasgzsY/lrO14oeCasB+ID5F2045mQB5AlA65AKMmA9xhmRpUBjNoBgAOTCaaOPn7sA
D6I8IZdjfDqcQkODuN5TLm/oAVo1UWhuY/Aa9uyNJyThCO576DVDnaK1cT+WopyGTkmllDqdZgiL
3BuR5YyMwTJxlCKlffBYhfKFpVaE/GY3BbBfE6hFUhRploMtwXCeQ0EpdhrXL2DAT89WLTg0Vxd4
Vn0mLCyzagaiYTSLi18QmTwj6w44u+pu1zgAzcoZ88J/0KQCVI7mosAylKtOlxZcwKF769oS8BiH
JQqIGmLqTNRtBDpY089LuCICagdCTecOCuHIKFTYv9VpiU0Xt1H8Iwj82nN0h5QAMYZTx0OJn/1b
n/Az09lKS2AUo74EO3V37s2L6qhIIw78nJjG12vFjZVFZJFoJWA8eHAX2wjyzRperMxurggfrjCp
XbWZaEr2lE3S2Kq3xjCf6/oasnQ0FoTyWXQE3iSFh7qN/Z93GPoBx440TZFY4v5z/OB4wYZfxzFT
kdodteic4UUBOnhZSLqtUYCBsg+JvRI5lYwKFxyiw10TwUEcaCQTJU1DbLlTsykS/nnf0lMCR7Pg
NYJkkPfWfM687wkDIIXHcqSdi4tw8JPZVBYSpdqWHxz0ZOZ9Ui3s5sFslbOMOjN0Fv3IEZknN9gf
j14O9MWhelN8q+lvhBiLmYMxHA7b9fr1GMGeZ7Z5xpnCIZwJWOJmXzdr8vdSd0mAGMWxmT8+UPjT
6yTNolJL2j3UcXTNrRfTnND14YEBtyTHvd13nkobmgEk7QJzw1te5sFywfAysJXohtqTWH1kbieU
LxcfQrekVwmT9N+4IKtSMxm2jGKg96RcJRiyvK+QCG2lIQohVxyzEas5Aag6WgbL5znlojf4aOQ7
Rj+3nUL+q/12QFRjCtjYjxrufgrkOQp8/AWwc4bJBNsHOYqU4nAQqa01dPF0rbCAjYmuF6Pbxwrn
v2cH9RQLd2hQeK3POo5Ym7oltxdw65NMzWZj9lkouxZ9rl9BW9193S3ZQuPkcSHDSg25TQ42koR5
1ndmw5+qdItwx4/fhnrKG+WPSv9Ec8Edu01wS575q9mDWiXSLvEza3E6JlueW/IhmA65kybGjgHu
n0km9d+m5sHOS0ds053XprpxdiKaAc+ghxaSqWfNCPKXKLd2xpt0GmrBg3iynZcfupffWju6hlYR
LpQ/6542bol4R+i7HxrHrpDxKunMsbKcf4ityjv2ifwZS+ealVkXqjMh2MFnIb8tIxZL6bAFrbO4
p73VM9vwVYyPa0O2Hkuv4rfF5ZzLwWlwEzQyphqyyzmQXm1VrLVy3/T8fyFl3cViPGY+zq4PE03J
z9rmrzCFSZGczbGcmj5Jd83cGK7Aj0NXEZSAZQbfipoE2PJEE2cGuegwMktfJtM1SUukYR3q1G2J
BQsxd3a7yyw2Te4ivFQ7K2KORZiK4MnwvxcQBaw0hTLTwJUCUdWNI5CZdn/U2+f6nOTroC0m4OOv
PZ6j7oXTTlabpA9DRF+xgpdMl6pS/DL5vc+h00fT7ipBKQjj0AnfMv4GWAtIbAVJbAPVt7Nqyg1H
gb6jPiIy6I02MhwY0ZAQ+VXU9aa3BXXGiJVD1nq3ZSzFVDNJf7isGqF8R6/EH6NOsQHdBV7xrejY
HlQ7LrhmyiwTWLu63+4RxWz3S9+hRCkLC7Pge2jfB8lpbAu4l0D0RW8QQP/Wk7KTTLMPAGVPu5Ky
OGQ1Anl3MpeqwpP/eiCFk6N0glAwIueGwu+A8ZgEBDC6ussvFd69GWfe2apbI/f9JBXE/9V2SPnw
vyKgbsMyTo3JlCpGLKkC6kQwbqbHFvXqAZc/2ErFcdsjNSSVPC1itvBURFMmSER6A/mcpW8JB7Dj
UFjLOFjozF9YG185uOd9eiG+lhthG1sTWtLtIABZpBUVZkOjUivxTQJwRVHN2BdobZTgAp3ixd0T
1qttUq4MyyBfiPX6P3+XYnahK7RIP/pXto3tPyF31siu8aw9aK2isdCfCBL0gtiK/79sBfRE3Gca
DW+QX4PHgoHxfTPY11NS8v39khv7sQwEU7blMiU9WIc87h0yuAqiXC7FzvcVio1DKRvix6Zc7wmg
DwFkVW9IwFPWTj+CDqlO5Bh95FZLRdZbpVEfbsDLPd7epnuS5Afp25YWNVszLInEoSGht2ltnLtf
Rh3tnLmSf/ueoaAw93PUTLN+f7bGYDa7ramCAQInWd2CogvR4CLRnVjS0PwMMAF/Wi5XWn7dl3sG
2V4myWVQOjnzfaj4bE+FRbyUjOc8v7JWA3CVAAiVxPAOJ3cOzWT3sTUUjsldDOQxy1KUDO6xy7Kc
sPfLaqzsBHyJ/u+ploeP7b14LtSnAEVJSNNYnQuByGWuZVX7YohR3VBpEtl/3JnmhbFb3wNTsWQv
ktK7qWfcummeUB4hYdcq6QSIYgLM+fgK2Fh5uuMUjeOqe8w6kU+ldl4l4sIpkBaHMQCmZGZ2Sd8N
dfPhN4UphBH3ES5rmLi00QWz+QdLQU5DtxwW0LBGY6cvwSP38j7Kfl+wx3RL6diuxPM8rVyHDD9x
M8dXVu0o5aT40SCqSEmh1ZmVxSJPlXdx7e/0obLEUTXjTXeBT+fcOgClKszKxGB6Erc5rPxh7eBK
uyhxNjn1dJx+O1Wzg5PhFRDTtmzuTmcQ+bnfiEoYE++5ffMCQLqO5TBOZYqcQ/H1kf7u9AhDgHuG
kMlNqXfuGh07KkP3rtJnN0J40smgLdUASbkSmqQKEOejEW8N4ABY3NqZSqtYg8q+6zlcODKcHXDU
wNHX+OxOxP0Gy+mZeSGI5GCh4vuEsODa3Q6QgXTmlhs21D4e6/6JRMt5usBvOnxOJ5X15ejRHhcx
5s5z14iOBe52PzTh+NXr2WXiNrg0iajW0W7FjPvJOK7C7H1+ZwMvtR3EccCo4/TbMXwhBvknM1eq
vdyE6eoeOsBqp1JBskGt2oYaaI6X+l4+1Yfcq5AjxwZF4tW11Y++ZwX/j09tHbErL53TIAiYsMt/
cXryBY44uH8WRnsgjnpszM9hB+zILIyxqFozZVnuRysYYFgHhkXwzQndFl77XIL9rzPl+j3jxsmv
bxh3dJGZ5/JL9k4yxWaOxUsqNTeRBZ6BAxWBp3AI8FC1JwmpmownDjm7lqkJevXg5DYfVTvCC/Mo
xa7Nas9FRI47lYv5ZfQD9tHqvyuRK6CtjdSde3G+GS8hDgYpSuQJx8v1Np8LLSrvRetLtbhdxDKH
rjvv0RwdE59vGr+Am2VaEC9qhzPagLvfAckkGdPo0JhOZHqN4T1zIANe5ANAca9fd+pSWTH06udS
atBGEfnJLEi6c53L/pB2k+BpY9Uh5tUdEp5ezY6TOFCbt1kIRxMK+xdAHTKELvWxp8twQkiwrCRM
NgFF5usWoWy+ujg2RCxd+id1/KoNRV7c272lDA2k0z+SIqwBtKxqScUDfNIbPqvZWV5entljtK4F
Mm/HEllKvf6jULwivwe6jWPY5zzYn54EsC2WxX7df/pr/NvhgwLX+AsNgr+ExO3cGD3gQh2XLGUG
Up85C7J9qftDQMEYpq5f65YY2cU4Y9+5tzLIsh6RX7Hblx2yBrgjMCpb2mSzjiVdRAQnH9phpIwG
FZITi80iKClCTYT1btWIrdH0xHXBpdTpq+8xaW87UtMM6gb8T4Am01cW9+iTjrMgXDKrx36NnCqG
Cv89izEGyEnlTSsDtXMVEOc7WRj3D6XK74M6mHUDn9eflf/PsQ9uxhh1+kjKHkfaYPKhm4UJiEvu
LaSpHw4vtMhcAXVogZa7WijZTfWk7mMz1CBwA7a1JMRU9hsWuugUe9JliLBMJAw3qvQW8FE4hlIh
xtPAYoJE4mOVKrvJujGZfDOs+SnTP7e6fTuVy8/DoIwiDKUj4Gk+mEsBB7z1OcY6i+4zsYVgwCrK
pkt3N7cPPXH6vkiOkzApwcjBaVOb1tI4swh6QX3qv3sSG0gBu+XeGJfW2EqywkC4pNoqh27JyTXk
1RptIP/zR82QU/ZMzaGoiswEbGcsKcQx5ZHWcJirEizsQ9Nqvh8ZXQ1RTutz29k4OanyRrgqgMQ5
77mE8FTFKfdKZ8Sm06qS5xj9GdOTVABHGoEF7bT73lL1qXkiVBtP8lhrWpBHOxblV//j2G1+Eec2
gh2Qc31sRSD/iIV+2UDyWeExlviVp9eZR1NbR/3L/o7fWnfPYFrWk2evwrwjWn9iik07ML1UGAqD
kT6QFI/uvQuetc/BqVj7YFkq3GMZ7CuOspLTV10ocjBNLR1KWwZjU5zq6RDobeEipSh1MqLmgRi0
7x4O47M7Xeuubx/ebEu5EnpjfiCYZ+oLPlr80pYFFmHZX3M02eFNf4LDc3sZ2M8uWmssrnNRvein
k36xKUnHtg4k6v8vj4XmLZHtFs5lcDA/cWfT81NF0Dv2SkG6SYyIo1pFBi5Jkzo/mIlfAXYCoyNG
l5llCyZItP/Z22DbtEtQpcdMhm6RIQe/yz5jt0+RXaqtJt+bVD6tXD/AMFEutyGTNqkEwfTThkD/
jhrU+wXrG6hY3Ma4TqqMBBHqg//RGWQUMINfNdzo4OGmugBm8WG/yLDNjRZD2fXWr8teTjdDeE+n
rnS4G9ajwhsvWX8sXY3Z4WRH58J9kvMl8yCGw01gxlox2C1AhbQtH7kd9HW47FGm+TF0UA+licvJ
ModXAEn7zLby/h4HMggby3vOAEo3+KntD6oEOLyBG7L2BX42KJQzF+wlhvD6QChPJRU7HCUggVqx
zdbTlG5UHVaWidWWCZmlk8N6K/and6Szz3DaEFJ3/lW4k4Z1Qa75l4uABm6Oco3Ri6jf2y4DULu5
8SJcu2xd7qAa/Bi2EErkZRRdDQKJiDkuAAteyi12jnovwUVuBl8Ce3avXVPNtMPbXqTBF5+N32Ut
A0UAY0HtGOyqnswjGwR6OwD6adb5Nawgz4wpZ7gIrsdb+M2Mev09683V4JRPmB6KCCVvDF2qhL20
MKTeq/oBwIIOdxP7tRVfs4pK2U9lAobdsEqxcPwLoe17314+JHxNfWFtGPai5fvfdXNh1KovKP7S
EQiMHiuk+KY407O/Rde072htKDw/keMh3yqeL+wCZFGxWJpPZbEkIoTJJUI9qBVmkIUIDiaBU179
Tp8N7Z1fCplvZN98YaOq+yAp4XHI9BJ/wCenb69V3nzkOIEEaCoQ/L0NaqT47awdN8Z6n9gx9AI/
iklygbVY+v+vSp6beX4On3PFG1LLyyHR+UPCUloLl6gmp6jelLp+kE9lyKldWzkO0lNe8c7NIWHx
qKxk4jnhebFPfsnYGyQA2k3eJMk9ABj1V3JhEoHMaZzP+QWmaprtb8SIBBoIXrPaNoBiXUAtmfIZ
J5JdiM6boDjK9N1g0NCIYlQ7a1IEFA0xXXa4BZRKdDRDIFM2NPiDy2mxd8a4GzxFZc4nTx/3lMfa
ao2txcIein8kG8ZOaZIn4mUOH+2IXySUutLmxlWpCYT8s2ynqyAEFzZhWj5fuen3pASBnBVjpZVv
uZieKWUVl48G8476EqMncwMsuTssW/6Ziz4dID+XCjqXQto63SFTN6P9kBROHxjMw1X7TrjObtBs
zOlafRAZfVBLKzOwewcF/H9w8HRGmFrP63VJUuTiL4tSABXIPAAdGzcLpI9Ef05Hc9AClT1EeDjE
OgkocOOv/s0AkFR5Q1pwcBAxrkRvrnULJP2vn6km7z2tBGK9a0WZqwbujlZXpOhfS5haC0vrXe4W
oXgqxzyOR2OZ0OGilxxJ6h1n343yILo2qfnUsVbBtI186sCjcgWUZa9+tCPM87IqEF/Cjxs9eUFR
PvuiXQ8DRzHdEAeua8IaOhSI3iAADR/FF1tE6Zlq5V563Rm29v05hf18aA6o3YZ9sVn91e9Py7X7
8ylxcHlPP1dZufoAvdAPBuL4PvMmLP9bs0oDS3xGtaLnK+QQArqjECllFMFMmiZR1UcOMNcdmmRY
peSOlqQI538PNII4WwDWkilmfFpHuKrjti2K0OisVoKOjIG85DhvH3vG5HRo8BjemcBTpkxCOYdN
CVAbGQzh6D24BxQF9WnVHWag7nEqOe2fEdIPOChFvKLsMSKtcdLDU2MnJs+aDMzD0L1CF3yEtkqB
Ek83jsv9nvf4IHhRNhXUee9Eri06V29KyMLX3wAP0F+i6Z56RWcC5oGozYNfXbO0Xs4hJqJzAVRJ
7S2UrXBC24+3dY2gZuQfjvTefVM+eug2rULBy/G09RKtGBv+qgO1yf44NJEp510g88Wx/WSiLaDp
/iyhEU8akRRGpbW4zuUwZegLfw9X+QqgyIqJ4arhnAyWbuVaajChFaT4kZilCYXT+D1GvJh74DmS
9rxCFMb9MfgRlqERsz9zOvFJKyw8zXtoWdcwS2zZbPkXPk8Ku2yF680fQl6xfWerbA05JXoR4Snw
0Im0D+nOzfLcM8qHyOLqQuU7P1k/rSmQ0yREORZ54j68dl5FgaSIJuZqygQrAnoyJ9fyhHP6CqL1
mYCQ4Pwa85OblZZ3VQSgfZemBlNuF49akavgUMINGbxtOcyACF9fBKfJkpMYzDkc9itL0kcRPATS
PNdx35aOrrKUOu3JvKmeZXecX0tLzbSsQmjlgjzuxuseCXyRx/xKp/XE4FYIcRSQQuneHI9vncsj
uMDZow2gNRbWVBpQWoLMlzXbuDl5LGZh7xbQYNY9ZAy0EpwPZb6hryQlTMEFiikCisTblGfIDnj+
6QUmrChj3HD/Ul419D1rmUK7rnDArGzTDczXXOgRG1ZcrmG6jkaZBcD4MBMk1uQud6HylkYe/gUd
5r636yDkeJsVYymq5XyNnrWQ4v8lwblcWuHYZ5qWnvtMyKD5lxAXVB+uhNtdyYqKqDHN1rbh8ad4
aRg99CCvfUNYdTy0K1odBoBa54UmPf0UnAchbmYA0HXKMptAHh4ImX4iB5QgxyZXnV362T7WDuAu
dtocBAlFwJ/s9wYgGGiqVFgP38gxaTcPvASvMZVgFwldkBf71N3uQ3w1ho1lBq0q+8NguLmbQIr/
pjJlfZRcZuPMzPkjaomd129EaQxaHJEN4bMnnxUXpbXDTKQLArtMPI8tLZc5uXAvabth9UyU1DVM
16JESnmg723QyHdW2LCEC9cuEHiDGM46SaKKDrh5G+N3CU8rBGRnXAOvzqgUyAG915updf0pDlDz
raKVjn/Z/T+VJRJd0V7t/qN+0P7uXnu1jjv5pG14L42JzQ2uzkvYHkW4DbyaCsIHbX35N8pKNAcc
sZNyqyz43/IRBJ7nXQGo6OiwQPteUuvDg94G6WZW5V0qXgV5kmGjEBtJkvz2MEaXaRr2eMXOv5s9
L/EFf8T5o91AJPMx0f+VEfC46h2vrCwJoPlRdmKb4pASALDlGc0NWPsfKyTS5THOzf3pU+j2yLRp
kC/a8+8pXRuz5vTS6wbfXIeYJqzfe8WhyrSU+f8mv7817NAaasFb9QNHHv6I8/2tVpdni3qkE8JH
0+g8TYzkav+7f368hX46AI0HmJARmYumAIRd6H56I9Eeo0QBh73mTE+DbSCYgSk+PHWkuQmmcd5V
VFB1ZjukdiriQ+m2LatABLXcS5DMpaZn2fp8t5255aYv7q4OkTw3FjXZZl/5PtZz4eQ2Ay5CTzkh
xwV+qVHU7q+/HsJrymklWHgGY7JdO2aGV+L41hAvng+boKrqmEfXYRybwfy/x3/J9cgfn2ToBYni
udtjDotNOW8P+OOjkrgPDIGSoAeeUrhjo6DaHEARsF7ylTg7Jzm0r5os+yuov1amxhA02LFlAEgG
a2bsXXmu5lGnq3efsMXGHOhVCHkAQcglHIbVbE+A7Yxf9eqrK/++5SNOMUHWiUWwO4GHw5D2pas1
RdNbY7KLSYbNR6YbVE1jlKl/sHnqZ9NQuImnvpjDwCuE6hNu80DhaP1WdDs2DxUR1yTNDPGbU/B7
1+Tnjzngqggwh4OSUpKCUJkAhF1mztz390yPIiDNFg6L68mfIBMyDJfGAbf8GN0YmdFr+aTwHBnO
VppXo76Jz7SBWgaQ8YVaavOQjfBbmWoQUdF9YVk+mpPz15Qk23nY1bB1MtRAWQayasF6FyUK9i20
E8VeDDphqbyfLC3v7iNOHtrVxe3VV6u046BPVi/cHli+6oP9cu7JbDPX04652DGN/IB9uaLAilP1
RPlTnuG9jl8NGzy6eDsqyuap3x4CtlHK+GCS8ZFyZiAjrAfp9LBdGdIbYUenj+Y4ayyt35SHe1+Y
m6fXuG/yZutjVQL6DZM3F0z2JeDeSnah0Ye619rNH56sUhaJ54IJhZ0Vs5+19FtMownBWo4J3E7l
3KJm0nRioiuYi8cnB3UyMrAGr0hEdN+atD6gecCJ5etVVRWnzzVDKmgzK0Bo5QN5GCSznuKpek+4
iaD2RdYyLERnohsi59ozmgo6Ufg2wOIUrV+MUC5bgiSpL3AgbmTEDPXiKpDoqXP2t+HKIJSZXT9P
yK5589AU2lQCqR+fIdqyHXvw3qlMV3zkncsKGJXZDLBispO2vtJ5qTWoKnj0xCpe/l3DqhUOda9f
3mp1cyDxjZ2baz/IQWsrHBesqf0Qgmxg2rkW9OMKX9PNkgnN7/mlylYvBAmStkxX2s1zYUnIsl9j
NDSA6vJA+LcRdgjJn6D57R19JdESyTqBR8vjQwR8y9b+/0d8U/w5TwOg6BUqIRsTSeXYkUJbCMt4
UnHhB14cm3GvoBwxs7k6jyZiEQ7J6BNw0v2OeaXu65aIpHzOhaBHsnklyWXYUbh/7riJXqeVZJce
CZ+kvEAokEDixflj/1ZXJJKrAHeMzIFEf6a0H4qton8etWGUYJmjXcHblZL/k/ZWFeOUlSt6tu5F
s7l0sJKA8XbktMnJkAaxMtslhyf3iUfj8hyl9kkk9LIfRoxhaj/mCEtiXLcbQxIuP+SPED8uVdKb
2IFprrwdwSh/ziUo2qsIso/SuHaUH7q1r6Audvx+5/ZcZBZUKC4QXitfYwjs1ZVeMvKztASqg4G1
HLv34e2JrncV+4hYYYp5MpoEtLU6RcW5obpzid13Bx6C9+6EHQsPa0mvFvV6CPDMBYI0yEG+QH4O
+w6E8KbMz12VkCi4Z3m/XeCaXhZl3DFwo0+xRYB0DqII4UJCQKTYcqe+bRVyQGIQsPqpMRScFTU3
sBvHSf6Tj0R8PG9eSyroIOYzMlJCO1EXJ6SMUDzHMJZmc1FtWCKpXmBcEyza20cU9q2uwboIUCCf
XdYhJVFyzql2O/MDY3MITMEHq8ksO9zkCEAGrs27xGZHTnmCv4IHbF7owlTrssXMIkYgvdHdjfEo
EoBvc/hKTTL9qZ4rma8TEEAkjREsFkq/8P7BxftMutsyKi6gGbTNVKNZ0E6W5c2vCL4l9h27/kEL
isjvnezlXsx1IPr50EPmPbStTK+j9FTgzixX0DcERC6d+xvNRiw9xz9PuYliLwjg/uvlDB6uGXGO
pfYmb/yuiJtGRqmJ36tKFWysvMG0RDnJBooDiNxhMZllA9eE5FCPAbT8ui+C1qJBopbciikwoKcx
iFVg1XOepL9KYQ2zOIsmCP5jdEYStHPTN1GpZE6PwHdTCma0j11lhBJUSGZlNC5HcTp9zEBZlovH
TrNK+ttPU9jSzNPdvuLewK+CEX8lVNxoP+ZXFyDpatC2ZYP1e2Y434PjHgQyURi6FAqhSCadaf82
cvKxIXZKH7JIvaVr58zBLDdKtmUSXS1TZMlw1WcejBKMqOq/busBulG1+/rPLG+oodMmeccu2tHJ
yJC7jBU5Up2P040A+dWtnyOx2wsl74uekS7rfLMFhuPKz62vWNjpL6+mHj1As9z0AfLV67iUPbmU
aCCIb6/K0sAI00Pfg6syJog7VXwuaYMyQarJSVZpcVUOcgmEsGBnURa+IM8gsF9rf//guUV9JyFz
sO/pu24TgwVNlIbKber7XhI+oWIJ+vWa74usDtdeeIyBhM7XrrP2SIzpae4srWWoCyNk3FL6u5vU
gXSnBjCqZQDJKFfay3uyU5FLGEkz25c88+OKQTZPjKUS03DMWxrE4T8c/U28qqZY8qogXwEjjo8c
q5CedEeShiiD7PWIA56EwmObA1b33zUHqMVFQfAcWC9nhm3JzEtPbZ6kHAo1x+Kc97DhZKfee68R
8SAp70XWWSf2AMRMszG+hvhkdU79hMNfV8Oz9etK9HJDmyjBzsV1+1dqECsxnf76AK645iP/wxJ8
3muX2tPFNB5aS3v+AvdTJEb7MzSt65b0XzImzzYNfYXFIk3wuCdlDeubT0I/wBckDaiXeQ131asQ
uaGDlJ4eoGNDyRHaPP5pZPsBkbuXWKuAFlxnlCqAGLXgHYflkfm00IABfLH9DZ5fExrlt+v4233y
/mCYPdVLs5gUPY6uxJAQ/lroiuM9FGMxIFYccewepMcyH/CM0aHv9M0zyVwy9VArOb/acXEhErbb
S4tE3DxpLWw2qLpVVwV388b96vOoZHK1LauMm5g0XcbPnH4FA3VI46HPOD/B5sq8M1QrRhEon7Nz
CIs4YR8VnqGC7SY4hxrvY+kpHBNrt6VD/WTlUtoVFLkbWQS0rdiqCVeJkijUzOI6tiNcp2502rTJ
NYNXkJNbhul3YDJVZMVP4uU6IP+liM7GaL3+uyEWFtITNRULs2FT9ePkyUv0q3fxbu+8vCgKlot0
HpizRRW8CclOGP3v5R1u/tVpKj74ouUUE17PxQ9ghYoyEFeaDCEqHr+piG2qp+yZKChB33+in5Co
fvKRdVOs+1cAUimdxeACIiWob8f95mMmepYej92KLizG+iYG53G+X9SrhFfGQ1FCvTq/B6Wurwsp
yT93bPX7cVyayoPq8b/OMVa6t0giVNcpQYKVy5ZpL+g1WpzzhcHougxM6AaeFRK8gYFeR1HAD/MF
wREg6S2F5q1FFCK5Wzabme4f5+3hjXDPug8Da69FqplryJrUyLkIEMqmuJCkqFE5l8V5U9qbVOJJ
GB24zHVwqDkD/rOo/BgD1+Jt+ZSjY6ahi6hAAwb+HQl6/lO4k7NE9p+NZ7AURSaIccohSvS2EmTz
apVl6IM5SMpn4gHn829ET1hxJl+2oU4UnOTh+65pfTqskoSQV+xD8/9D1tMimq+hkY5PlX75RtGZ
VWbF+pBzuZIS9gcaXpy9ioXhEBjmN0HY/cZQgkLSA+240TVchMLp7LqZvDN6tFNY9KIiaTFAjjNe
Zd+OPeeg6IRVIhEqz6WyFvVvVccf58wWbSylFEAy6dhlQe86xxUPYlD6ZEPMWhDuBbc7mTj9Pnij
PNW8vdxb+Xua2+vstkuhW8L64HeYjV1DzUasXzVVd5qCuH74v2CUuGV7R5uVL0hh8uFtQJj/eWrf
jCrVyNhkQRKAAzzcWndt4WdYB1fGyh1FlQz4o6mRB2o6F7GzGZNgQRx1lcd6k/3Pi4qu694G96w3
YBreQf4CVY5KZkyQjvSg8aM7lydfb4azAM49L4S7ROkmSMBlUo2XCd9bqVYnhjUHBp5zhQIl4lD3
cd3YbB5bibLdyhYrE9gJi5FrqWIFWs70wDjtOFL5N8j7oIa1kBNrzR6j68We7Ol2OwexW4zYgdGV
hPqI/CTVuEGZmKw8g4XNR1p5LI7b0dr0/NwRhaykgy2Rq/M5fmjrl34WCsJXB8IBGV2MuJFkxW9a
nomp/KuAemriPQZKmM5JXm3UNeUnKlIxoiGXKSt+CTHdbuOEAThApXVmihTuYbDCXrj14rePPKv6
rxRbd6KIwoDHtIvvzcllusA1VZswckryo4NmnrSuPRIxp2P6/x/Wk2gI6IeJef8zNYHtsBiIreB5
uSU7MPgZ73UKVGb2gwBswrdsYJDNFVnpST6kWf2sZjPgjPKI6dOrejZ627ufgkHDmybBiexkNNlS
L+y/lgPRJz6bLabCsLQh1Ag4aiB67oF71YUTWgPuw4dxePHD/XS+VM2j2gKhOPVD51Nbu5ska+u0
PtutyLclHqwo6oo8lTmJosjPJm3mgUvFEWbCr7Yo6V9PgWjdAJYHC4fNvlNmiIRsCiAO+hTz+m6F
vejAakjzYqdF1anguNffAhqVW3bkRwh6OslBw5uMbJOZSMH9WvQbGIO2kOoTEOovlM1aIJou52H1
roTrjVg95AEobeq4Q6RX/v1zD5QOvqK90mShpCEVPchtPJg3yxsmzb3QUlgZWs5a6GtxWObqP/Oz
9SVbVYNh00H68xQQRDjIhbPt94bM/8Gs5H0cxf4yB9bDQxhu3P2DKdVanZp8tHss4YmzTaVzLaYf
bGwuycQGzO3ejV3wcEp4erYIYjIKnuX0Ughz4E0728gHrjgsdUEmlZTQKNceeV/4QOIdGYuV0gvV
XXSQ4KnWxCqWt46dM5iPN3L7qEF1l7JBFPp7Yyzt+P4rR3gPI2JyT2H6vKU0eJ7/TYDq2bEUJ06z
nqXEJqQjFlCVJnA+uiq57b+3Eo2Z2a/z8bjLinADzY3y16MgaD6NF+t/a6xjla+CJTL3bWi+eGAO
FxQovdy7vfD7D4jA++QKaSO6WwdJKwkjM6MiKqhfhPOmjaDxRk2McpNpwRa4hLjQKHhnd8weJseJ
ndE8MjTpLf7Z537m5hkfGvH8LyH5rDmJkR4WWBWx/Aw3HSClQ67D6Txu+2gTAQOAR2lQZ4LcErh/
avDGdjnCZ8SsKvAPrW6yOJoRv1EJTf9zXQPQo998uyGSF7Ij8UNL+aFww6jQDRSq8pY/XWRRAie9
Pg+r6QjYvXLhEr//9qtIaLIefPYyS71KFV9V7eourAeEauc74O7bTGDPZuPn/qtt8yLVUKGviYQp
ArwmxCtSDGztPyCe9t4hc+XaXTIhhKO6gaPiHJgb4d0jiUspT6sl7yztdtGjBClstmTAaRrOEG0v
ugKGKpYPQ6tA8np3Fi+UAXZe0vh4wGxIH6yrYIXgVmje7084KG8PcsJ57QC+A+bZxTAKzG9dymyy
0wtgTjfXWOnIhiGezZYbGI8NfFsptdQRXifeMB9vDNLdJLr4OOKeODom0i19WfBpNSWQpet2dknc
y4Wdow6oboaMlkhGo4qEdpvDt8xyfbjFI3jDx0PbmHZkTpM304QHT40cQjrQkKT+0YIaTeEWBVAd
SZxqxHfhjBsTj8n8io9Qbr0vCvRcFPegoRU/YlWuqIEuhmxBjnnbo8uIVKz83Z7eE2vq02eZLZef
YwPBb/Lj3l4TsHyMsK9K25O9emUG0QRF0i+cic5Zfssh9TwLmDCBL2IPqui3Ofv+4GSDZLhN8n1B
tXe1OGHemWNhI16xgVxN32f5R53UUDte3e+a80gLO/aFA54FAY9Am6iWNqeYw8K4KiLtfDdozXe5
q4QudBHFD7XHvwhqIZ37YuuRI/NvID+RU0xDsWQRzlEkLwdCclDqQkx2IStZvgGmuMUJ5XLl4L9w
PK/hwxgHtGgrAsTOLwIVCdArlsh7yRq24JZ4dDbhcqg5Y2hqy1tIJkbnO86EvL5OZ+htT+QxrTYX
92BBTGaM79G7drCWFbRG8qedz15sV3928T0KDOTYmzENqwuDYsTq2NH8UV4Q/ACG9YB9vXZnQCUu
BLb2PRks7MtkKvbNt1JayOKxSurbYf6rswWP+J2sBeG/czkQqujq41VrxnAKQ5fa70tNKN+qPc/k
bhkiaLBI3umyN9ty8pzV0XWakyW1RbQsoOhc3RW32tvQdKFWyV9DmV1dbmPyZXend+NQjl8Rc+cV
EPjDNc14F9dXgX0mRb1OTXdOfg3jbUBkxTcuRdmo5r3h123lM8HinUQ7/M6e1NBITBuUtDXlxgKw
0I+1rNSSicTOlkJHXFSorqQ6+LEk6wfOF2thjMNEQvTnLO1yHHHOz2Y4ktULOh9aUtLJih86Ultz
acGcXRAbMvpQs4uDLt4trsO8KsSWAP8+GRzJCf4wvJzeaV4WwfmWMNTbPIBLkmTB20Mj24nuxQiw
qZfi9wqsxLaSAj1MwJBwaBm5BRnMP14hx+g1xGloY/kyeGxfK54lbKuu7FE9RqS2ff0s3cBQ33rw
X3nwVlP/Nlwvj1/aWEQR9vuVPoOiQ5wCnyD/VIhKOCqJc56q+MjF+vnhzUTeAaYR6LdkXtalAHp2
/Ns/R+AvuPXZRTJB8ti9E/jcme9PE6tRqUdnf/cTVjNl4YpVp/WFGbDJRl/qUu4m7jbyTNyBmI8X
5YzN7759jRq8kFsZTvYltWKs32GtO7s/dnHnkIuNeFfXUCkPoS9DcT5c/KG40sG+v76BLHmQw9tM
CO3dM3BAYVZSUPBsAUJOhXiz/rg/7KxRgqL+QiA+x7sAVcpGasxrEJffVJgIY/wN5TXG5hzZri1y
9F+ZxxujnmcnSSNO6BNIJKNYsTg4B5VHJS3uL+24rS31OFIgwndQse36XNJyc85Z651cPcsSZb3s
lSPo9leba/rSPa1GupPFPmEOOdgJlyGc38R6/akemhbTMYYLofw+L6TSVGhbCUgPkwgfaUbt8ZTm
cqOCcL4rCakOVWoaaxJ632pIt4gGij/VI4FlUZJlt+mXbncmgzLBplFmKv43LP2cKVU5coVJ5GLO
SBz2u2cRsj3tCE2c7pvHmpEwJrnYAW74W80iX/weMSlSYuy2fwKwQNQbf3sfJL2yHShA65VXGpXa
QcvCyLVWUc16VhWfYHLuDmFXkAzp97uFuo6Mq94i3GenO5F9LlfGz6dTR0TK2hWMvhBK2zBgngEe
tWvPvJ5xn7dvy+FwjFFh4EsDE0DqU+E9WIcN7mOlDrvE7DNxNbF6NU1lLZ0dNxgx5egmdW3P6HmP
iJvoSKErKwR2ynocOjLyqIoyQPBOSMZ+gqEz91gO/abgIRg07Bagh5/djm7Ax8tIEX0pCjDHQW90
B6BfDGsULAyG8kxDyZbwrcjTUd5xS+8vmH4/A++gbw9FSVHHAwFcFy5YJJr2qDKL1y7qmwSptir0
iiadg7USi2OXFZwy5jA/lGx5xDr6sEZ/+R/wyC3fjkb34dy/ZBEz3aUGBUvX+A31jegKzykB1H8z
egPLjxGhZHbpraFJinvecrHyZSL13AkSjspx/EE2mAiGOdbA7kwfHwEvkbcj6GgoEORmBgq4kiMl
ahwXsvvk0wYojPTaUN84c+47PY/5FioDs7BPBiSkZibWwJoQgnO5On1UAhUcFcqIbqgVGNaApUOU
w23brkxv4Fvv9b2ZEkVF25/ah3m9Hc5VV84lVcvvgBx/nB2Pf2qFvoRRAfS+Z1FnsdrvtiDvmTjy
XdcoZ+4G5U6Lxq109a+VAkYnzgt9eR/fRtCyJMP07TigRHJ4zxRkRg1G5Axa136/8mDFO0/l/Tmg
BBpwhc90s9bvu8PFF2RBo6BnRAIMMCGtCBadRe0Yvl/JmYpckJsJA6d4vzr+/EZ4MggJofJ85Mv+
y6mSfeB9NXjgVE/MbwsiwsA5m4TlwZ4gAabhBGOJ5Udj0xeg4s6yccOmCfM4yvUuTYFECjrK5sNa
3mXlhs5NBHVdtggb4PIn/RHGSKKoK330iXTcBFhGiTPsMfqslP2SrRgAmj0Wm1TK2cGBQhNSL/bk
CGAqhNtxy1lNA/SsdoJxTY+79+Mx16gCXqfN7Ds3AUcfH8XPIgqlruF6J/6xCuDoJU44lpesSmrR
2ifDJt70+1If2EYxwkPS4oSF+u7yd/AZBhBCc5PSaZ7sYyokDRa/yEAMj7Wb7sZo3oaUF6WHkZHo
FcEwgAiHfAx3+60NZMjQFDcWYjVWqs+0rycbhibyUXQcd3Me4n796s9xpqXtur9IGA6ZhcbkVWQ7
WNXuSUpsU/1doSI60KAM+UwvwBxVS6YCr3t3l510jILKkD30rmSEftcHCeA2g9wlTs0MwrrqwM5q
xlQSmw4OLw3eh5a0leho88YZBmFM+LM7mKqnSXPQWyT8d0RgUleMVGS5VeCXz+gx+R0qKvzgCAw+
m4o0jCy5BMa9BJb6fjXQxADYkEm05pz2q/hqZZxSpoPMZo8uxXUr8S6Q/j9nMdWJnRwUzVqlCKOM
2m2uUugCpPlYTe7/6Ibw1AEU0uMu7hHzX4Lgo/w55XUC/NNDseGFodjNN4c1RuZLXkI3gDGRkQW7
JR6xRy9w2043qkkqCuXY+AQtYmOlGfOdE0Kt96DfG5/MlBRiXSUNlELLK5yT8aTkDSrbSMkvucoC
6nEQqw5xvBFnlKYtI926NmHCy/QwbVyr6q3Gh2cFRnYkEwEuSHxzlpAIO6+lBD9hS420zqxllUHD
lhyOTDXbBqbTX+ouaT5cS4UF0c7jqOvBIYOBe4AEAANE6DRy20IDgvN5QWKK8vqn4KiszNKZ3vCs
iDgE3ayg5xH2gzQzD3tnbw4XTY+Ra/GDZ5rE0PVsSk/Z94DWn6HzJO32rUHhurW0XBBV3I+qt3Zp
Xi2raUjEVXGtmB8CqUxjPeKNMLxNhwyJ1hiIFauZrACkVOXsDg5K1vRZOs1dz1N1/qFsjiSaFDDo
6E0KKl7unWElm8iPl+w+GGLyMXopGU+rwBTUnMt0k2+LhJOpyRhdp+NkIYeKXABEthTJMtHi3Otz
zqWhvOjKPvKZrkJv/cX4LbMAAqUzzvu5q4hX5kCl1orRpzeaJ6CL2Ld/sAAoY6C19beM/+Q1GhSU
GF95zeKZMtawfeoau3nX6TkwZJo+rkViugDxOonTl3vg8bnNN/+YYc6tUkHmTsSj0SYpXHtlqWk+
zIN6W+PHMnQaiq9YDOG3fKOZZDfoToIUKP1dd5Xu+Ol4cWbTbmg9qG+k6Ucjqm0sDFz4Fdw69AY+
XDuNVtfHV2BasAeYPzfI4noYnvPq4pGhN7pFScgMEyoNrF0ppOMxEo8vTwcBmYXqEbBH0hMQLOS1
p3Mpolw5624VZm0GC8f3u1iNpK72FI6wt9swCtCdPOULWpiiG2NLO/AEgY8HR80O48Xx6XPINIf5
apMA+iMjAE/656jYjSo1/UOQuy2oAscaIp/nQ5gg/pY4hlphkwgb4qQHaSuvSW0AGuec3bJhhA/Z
n8W+z8RdsrWeMDSo6e+wRwGoC1PepoC9TFM7tkhZ8I30vHf6+V+fqNyQIwqvZP1p7FhwTKLm79wl
jML+QedQsaenMW/N/sCmVt8LY7LkmhGvo7DmIQZ8rzLaSs6Yz5DKsnwHgcq+nkjEAM0V3L0g3bWs
13BvGuDrLwYdu4PluTwkd2igcaaUohWbYkWwDcWanhGFzukU8WnGEu9Saoi3XrUx0Tpqear2Q2Xo
b5lvxCawhjZFtFv1vSFNNhb2hjl9Z01d1asvdxJ1RIlKaE8U70WXyaPBgPlKu+QqtxGJ+00d3Jnu
W+UWYn/YngNhuprCU9rKp1d+1r8oJMD+PoEM+ajdKOqJu5x6S5sjRVEGk8P3zu1pkJrW53qs7AFo
3ohob7rr/A4V4rInXQdWZUeT6PSnV38UAeMLDUjJvHRQiVv6maIre1ylKJkGS46yaGeezbyscmDI
ocLqfcojHaXRLM1O6yHd11R55Hd0wUEQb+s1VpzqiyOtcXR+PdPoxfZbtCycg1Uqb9rt7Bp+ncTX
IWVsXC3IbNiqdtypoh5Yffn4jv9YuJQ9eWxkqjPJt3tksCrMlQyWFvjPwG/sG4NovFZqi8Y5w0MU
U4tJZEkMQ59zf2+DBnBeG/3bg6z5hbIdCdAy8SQDylMsOXvGBDZDkjJgrzMaiEGdQiHMJhMPGnGT
khSlNdw00lIubAWlmExua3w1Wh11fNPs8Ubv0VKR+ZflOQDUuLZ88rrazXDzu55lKXIdpugRg+n6
+3rEOzFZtB+/37gWuG7oXhqyYdo84f7nfoisnQFHJEy7NH2vhs09qLdgufQYSw3lI+abKsKvmKbG
q60oW5CtdgVjMbFoxWMBjA+B5eXHGIRklttH/HXr7hw7+dwIF18jX1YAqvRCI6xizKyhnz+6zr5U
5RENumHYBBcieVK6G+Xlg/Ax3r3vYdWMn8Q7yKH30fykgtT55aXCUvZ1rDdmHEjx712/A0xNizyJ
wCm6My3QX5M9q09iIBlM0V1+Y549LgarF31xfwk9HIjKvTClbRtjrBTFBSFhMr6jvE0Y6wtKGUT/
j9wkPM0cwNL8MHzhJpIYaSt3lUcgdfK63xI5TDEVYwHddjIIh2smcXrmYjq6vfkO0KwXXLVHj4be
ZCKUyrUkksLCVg0zERZz5H5+qMGdQ7/yBAeubcHf4gocAmBw1bGyGDfcXJEwvS6IP49Q9jI/zLHP
e8uIAvNPLU48woHstDv0w+P2g721tUcouMZKN5Xr0XOCBtKxIOUFr19UM++oak9WEhryBzy7qgnY
1Su7giPUqwblMFkCfvVam77wSODjKQs8mDlfHmiJSrimeeypcpT6BhGrgJ/1RTSA6KHiKxvqviws
Ol2rVHWG/Z5WdlC883xbeRwc3Rmv7LNNtrZU6OW77AVv5wGkbHW/loSRrv4XPYghlEfCrFI3d9r9
MtAJAKRVW0NtqmzC6NIX3sJGeDBEC0ug4ncaExJkuU8zFi7Wm3feNN29wgcuJLUR8cPv6zWuYzEM
7exPsAprqF4DGx2QND7t0mGOa/L6jBROAJbtwRnH8Jf+uY30OSLARDGGko3Ev0rCXyVgQnEBvT8H
/OXAb4Habrwg7y2C/xWstDuU7aMHU5j21lM9ygWi+gwi+R47Q2OTmoQ1m7kp5VqJ3EIWHL/AfTwx
tw7G1KPcX0ogOIwLiJj9Xc09PHHyQAbXRB9TYPHrCVsFUzNNZIC6IHhwifz5s8HIIWTTzAvxCF+1
HAXfWlI62RkynNxcShlDd6L1ZxJHLTEJAQ+XdGbD3TxzduMcHtgvEt+/JQVeMGzsaJcwgfO0nhot
EyO2WxYxzgfYjrmbwmtFug7PnZJbKoiLk+QKH7RadH2rpH2Zgbvu51i7ntFhn7Y2Qhn+S7MsSOCe
DFtCWXPVn2yrcG24AF2RoJ7zJoqckCD2EKv5CatU0f9xgwv9578PHBuTHA0KDB+DqDm9XHTNTECt
OBp/Z/Jf0LZF5OntCpGfDi7SU6038u95x3vS/8hbHhJrtqQtMkrBcXhtJrFLk/MJr8E4oPf/G1mL
k7ilPgHxkKoF+8FhD5tRQRelYZUdTHBe6HtVNPukyGPD60PiLf2M/4tJ/NmuyeAV89OCKQyBsUDO
QTvjuyx/kTCYgnhyCIOxxR1MVKnHCGMZIzwps7p4ZD5Y8oENEp0Wu+ipfdTf5DYDcNiO+65fZpM3
xq1qlgNKWhOkQkDMzJNRWuiWI1w8ZKoGWzQcnz985ZVWIv2aK28UMLcA6ZQBgj0jOlcD0hxX0AYj
mVmAgtbMDd3C2Ymeqh24QnzU7ISN30w/jUP8zuQiqCfjxaPPmG5Q1PQ8eK7H//XCgMJUAmDhMK6R
mwUguitjMnKHjaObv57MTyI09UY0tZ6LsxCtiV4JhYKtVzQ5+87z20O8PgWOs3wcqFjjLN+hqkBP
rwt+2Ejo8nMtHdDVQNYj03CY99zdWKE3y3QcnumlmgTGiKV64Rys4kn1xhQh4qoW0g6dSX57mRK7
fAwq7OqKw+9vIPOlmbWw2kPcDps38bK13+Dwds866PcCJde4b2CNHXhO/DD/FXeV1DkyGhfE90tY
NVWtw3XA5p8fIKA72zLvhlfsVPUYKuYMyI+5PnVCDl8mkbD0v2NV15311GjqXmIzjfV7hYIa86j5
ODEQHa+8sj+5UYikHQOtSeO8c4BnH2YidYxXWtUoZa8IIJtVsN0kNSXnNktdRmGKJmw2k4eIirsg
5EEKKIObEcxSHWGA/zNhYJxe4TTPnHpgEshEK3BSaU6lo4lvUnz8k3SUpqf+F6ViYkMj/PF5a+iq
4IaV/yYUqCwVO/SfiuGmsy4sRSx22fIsjPhIWZ+XHJkRA8jmEdmhlR8Bcm1DpnirWSY4X59MoitH
u26Jpfq/GhrIjace0HRy2O5DqMDnszd15thVSFqxYpTfXH4KHb714KOMa1tStgic4n0oa7MH2bJM
1HpT0M2jJwnvFGBChHMiK03ob6kUuzO8FpD/88SySPNDA88aKzGFovcRWjPBcZMEHtMfKgWO+c+e
7crk5TNp+TJFKCo/JIXH1s1IzyLBwiCGf8B6tlKWAthOjtBc5RkGTuGu4LVXr4cL4Xc/l+YUPcDV
HMPH1xrPpTbMYfQV/i2neQGBENyp//xZFm3Y609ykkiZae9FaYin7T/ENLwVCUuZ40igYebFUPO1
GXoM9eVvwPqzcm1ZcMnLFCvcNF4kZTMiPEoWxlTl4RoZ8xgtWpmGCjKpA2mp6jeClh5osZgNtAXS
Z2SMyfoa18HqKua88jloui+l66wBNuYdqhgLUguU3F/271wAgX+Go1P0YBN4QjkrGClFym5GdZSu
Tg1sTRsV8SIop9u8/S7dLCYG8G/WANgVqLlBdhPUrxrnBaIxDUS1lf+rSmwrKdvgo8uelR+GpyzP
5OmUCYwp9mkDGcSH1v/ddUf+unXX6tK+ONNOQZHxF7OhtOoDn7rg9B1WtnWIRP4xczHZtt6Ow1G2
egp2yQYEtWDLjimLZh9fSKVVRqDza01xHyRNjOnK7zYnCyen8oK12HecXgbK3C/xcCed9FaSUSaA
w0nft5beZmXQ/bBQ3H/7M1QEAj5wJJvI9Zp1t8OHsSgDxKNbojuvTqNgxkhHQ0NyrNz2BCQ+6ZLJ
wPE2JrWki682eqFw3hfYANyI6p9QG3pk5DvTTA4GWg2JkSZvPQwsNwwTqYyU4ML2I2Nn+k7NzhkR
MyDlHVYrCAlN0bC9X50gqNQ6Kz4TkG6RHsVVkeqpSk7z3Odv8mC3CiVVu7T7oLzc5gN1NetPZ8+r
UrCRstFKiTCMyO8PqN+67r76SWLuvlOqpH/v6m3TPpcX1i8Fi03eJacMnvfMSo/xZTd6WIwtN4Xc
gaJv7U//1Bba8i1qf2K3AcST1VUdJhb2V8GRW6KrIWHO0041xYGFpAmQneAdQCPiuKy+PgWzmyhR
JZnEpyDtF27Kd1G9yaIlcjDsRcomqCKyX9eSkvJGAHs19xQym5Cu+UB2DQywsBE6UqgjKUlpWWHt
8fy1PxUgvGdpAEbxSGgG//vgoUZ0MtIjupqN3nxEwTnNvmCmeIvSCkZbTQgAMKP2SOn/kxxmPihV
uylsBU4TBjY3lD8d/qlrVTruhfrDoXvQQ/g9kOMqUx1PpnoIr7QhmkX/DGpQod88AFp4MQHSmOdd
ZPf3Ll6Q/aOhL0HQFYWTobPpQ/M8ptQFKEc9SL7QmAI/hrFb2GPGoY7OdIAygBS4hPAzJwaEGMBr
iUf/1IDoULDr4rdv701ttGnCZE5XEbtStazJ+cNYhh3riYlh792peQyn8zdvYev+qHZUuvJOq+wA
9Hd1B6X7yUvrR24iJ+3U7h9ce7Md5LT1BT8hFrmOF9hfJRBt+5aksKcICLe9ift9VwfCN4SgYjUv
JmmqWsOYizl4
`protect end_protected
