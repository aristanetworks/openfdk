--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
ZdBqi++Ph9hpgB6XXJtkh9WIFWVcNZ+iyFONQblK1ZhcojWGroFKU/Yy4g3rD4JWLH42tGdHbfgJ
A31QJyMAWsuCoHfl2vTDliu5IHy8XYDUgseniyvR2SbFiyohbyq0IRo1wxSLonJxaTr72dBWtYAf
tuZW7K8W6a52QC4l9KBDVFCm3yWhUO0+oLZHTFuw25z20mQ8JU9IdrEXShhjEG9czXItKo7PUvcc
lrIIDY8TcMjXBijkml+DfqAt0NflwTiSfoNNCn3TSAj4UmSYbZ8v/QerCO1OFWU3wKfluCUCpsh5
6PozXUazdc1Y4mCpwCCrbxKOgvRrKUbYLWiCdw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="SPXpS1ijXcBWgaXCw+5tHJb4ToCVV4u2hYyD2DjJoX0="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
JG7zU55C7chQq6JPFxaMRUFsN8r4KR2PdEHGG4KVYH5yK1vWF6+/rqk0Rfy+lOnbEFD3EglGxwmt
4NVZwsciir5LSLww3iBdFfcZq2h29HifbRQ4RifQVPYO3k6ACcgs2HLZsr1gxKS8Ke+03L33YTS+
mF/6JpPwuaROb+uHq+lrUU6AmeTZADrsyk/dsBFd1/8x3DA8Cqap2vRxqy7zx+PHmm+55Ma+P1aK
fkcQA++fTKERbTfC5H7v6ZoxhEkv7HoKSFSfm6ZDkQEAim4Lu8NsywLtW7srQ7TISURy0hNwiAuT
mTJpD9bkJEF4xN2+AHcBZJPV204cc0BOqHbVFA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="4iTXBpMh5FJEc9ucU97nQTA/STnrg7dh7V6Z5BMr1dE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4672)
`protect data_block
ZNxWMSAiNb5aXe9mAoSBtFfC9t1dCGdlGXCGw+Ffy74I/wjSpVO5J0DojrV1jqN4g+p9muEGsU4+
oNXa5MlMm+V+OP+slpydoAsd5ZTOIhJSU7YIU0xCDQHfRhbBZ5ElSYMmy6VD/rARWprHMt6PAFd1
2u1wZRopvoxa37H5uwpuuk+yToaNrbBSwgJ3XI5xJfCruVQAbXkPgGVPP4Pv38EYh6lDJ0VnVwja
x6Q4QurAoCx5TuyWdxysxkLHnBcNi0TvjzHo3fi7rk/1dJnuFEcRCgomnjeMt+huz1GQYGL2ONHf
bdzvb2QaNMc0J4D5HAKSGymOj5MnSGZhOsLU5zuN6f/H6Yif+liXfzkOtS/mhyTNnCT+rCet8azU
ryUEoizGKVFdQIBC7NjmBP0vTqw2B9J3bKwV7cf8ZuClqSuJ59zDP7DiSSTgBYb7SVcmaYeZvfAV
l1AEyHYTlgeYuNBLYp+Sq6yau7W0TobYAcuQrsDdfyJuOpZJFgchQNCUHD+DI4RnN9S8UjNfJAiQ
pgWQ9oV4VdlHzyZZatWEMPRjfwkvM02bFj3ZIFnc99PcUPoJuABQr98KOa3T+h03nQTb0urLzrox
TrzE6DovkFFERh/NUaEGMgzhOAfXDxFeE8SXdUdTAKSs+SY3GXjguv7oT51/odEFVTCU1Brdg4MM
UNz01sSz54iIiYZY3DttEp4nRxd1v0gLAUycQgCN6SY6emW/eIgLfP/CWa0YLRhf99fRRQhVPxGJ
ul2Z/AHxe4BX9fxtX8+UZGB9GUsJCSzmD+yJzylw8v+48sqY7TuJA1IGFZCJBVz9nV2951lWnRDE
as4n8i18qrB74HDsLHmBaBURpEvxqTri66KN1tdshcAklX2GkXt93NBGG1ILT7z3jRX8IZpVe24P
HqseKxP0hM8SX85nDSvy8GAWUZjEi74/liwuBuxYfzqf4k/nMrV73aGb9mFHI+YboNzoF9xVVhhF
yubYei5IV9n2JPCaOgBWjDy1WNXUancbQasoqYjltNpzUycIbm+ZTwandpZQRQktJsdvyj89MHJJ
eH5M+zOOFIs0a9tMu9mk+2EyrvZapW8YWSsGyi7/nhyasuuMUWM5IPYDBTz16fgzOpxi4LxryeEE
RITa+i31gdOYnJYX+/++tu7LubEzyFORjYl/ddjMfWzsi0dh4P2qVXhROun4bw+odrurFOJiWT2/
oaxjzUUTjZGmBEoWjQl/M3ER4CZhbUO6Y7ZtrR4D6bXkpKgfvVDpWMewxC593mlK+tuwf3S9WgkX
fe9tOflzOO0o1eXdS0jFwArRUWKF3efMgdiH1+SH4vREYty6gKoHWBDCdJ29fh304Yybxp1skSb4
JAmvnV9cKle1huJMUyK7OM7qw1IYgZ4SuE9kyT6MV0pOxdW0T/Z8E6PMrGTNvvr4STKoPi7Yyft6
olPgFwVkKXpSKHQb5zvMSGpmb/mP1bg9DUlWjUMOH+YCh71W0d5J32XmkVEplRJdcGXr0IZiSd0P
maHOZS00EEf9IqLaMHR4oRUNpwd+4M+NiutLy3QIQrAaU4cXpngEb2vl2W/lw/+8IGP9+tn9L1eY
ZG6rXyObcnlCc0EWfkpVRbWSWq0gaLnm+og4S/feAP0e4Ov7UEVkfjpzRdYwYuWHQiG+qi2CsA2e
g1pVIZjXpw2hZF1xpiBMPrN+tD3Iq51LkRlGHgxUdSxFpQVV8XhysXLodBIcn/3mcyaF07yxIj0c
/+x1kuYRFB9HKDScE9GX+fmorNLU0DZhejawA8BphUcH9PG+fDAPqA2E85rtAd/evBrCRMoCPvez
yyungjcxEX5rkHGRrZDqf7JQdZV4ps4ydpvqXENoaZZmrarL5Ejgn1LnRk1HQCmennYkY2d9ZK0A
0eYYXDpFey82R8GieMtkJ3jV24eps1BzzQliR6pt4IE2AqXpi8CWCb/UoI/7P124M8tEEB+NdQoo
iJ0u3fdgV0Mq9t8YKxb+n61ZpJwrrHTgharYYN+1XkpG3T84Z5c/Xi4dr/5kz4pWziBRLV1eIVa/
51+ABuuEBiCFoKZnH/3D5/P59xRwW9mftVw0KmXv+Vl1wltlWQUi1HemQZS7hd0CnhfMjBbKGwrG
NDY12CWVsjwfmISQq0USqMq5qHquIl73QlsBAIHXXbKXszZ7E0bMbLyitVrxJttsrq19rDo5G/MY
X8tBluWtvl7Yl0C+Nbqrfvs0rix/KMMLvhXpzJfzDTF/gg9CLWpFTXUi6AEjcX5c7waGR6PH/yU1
Zok+D1r96NrfJyv6pGw8xD2BSzlSDhbO7iTz5BVWBha2WePuEYcsHkIA9/Fpen/Z+ODU4UDUFQRC
xKAd+sl/YMMtx1zsanlM2rYIvKWBzQbgwBDaSngQC9jl4HtDJC6ZTQce0HJbLcJticpNeqaQ996y
V9/kRWT9CXgv7ti+WNNzY2wJH2bVQJLhwsRbc219nmsBRjKTVydLqEcBv5yeS1GgCDme0dqDhF5U
lxzsuY6gTk8dBnTCGEsRiNLFs1/Du8vE86392+3lLtARGjI6IP+zUa4WkxUW2RZHX+I84kC6qlCJ
nRYWg58b4eErsLnQDf7audf+sR0ct2YjiPfIxZCvoETnRYQ9KnoBopxRcmxMOh78uWdZA/3Cg7jJ
nOuI3Ey5CutYeweLvn4ho/5HPCyB0WBdlIMtKxQVGN6AzsfSVjwNX42DgXqG8H8UG9x+u2Ly15eN
JnvcHvVyuICKznmHaSS6m/Efa4Sk62eZCEseFLUpsxD0bmAonqznYZs7tkEApIiN4vh45a4Ze1Iw
6iNFjnISmrD3kcbhQuUzxPAzIfZA/zbhqhnmEIutJ3qIaGl3OPD3XhUGiyYAZRuAtTuaX/2DV5n5
sfzFSOsYGO01EuPon9Pq7vhyBmMt/FZmP7ictvwRFiugGp9G5SW/OgQrTR7Xgqwznfeoo6++BAZ/
q+24D02dORHEvi6sKFFLBWo9WrEmRe5m6Wi603/1VIXEm1N0z8SxEK6rN4nfBMsOOanWB8LnJP94
ehooktM7Stcrz0etfVZKQqKK0txeDgNK1uPll0BeuFVE8zTxIfnTMZdKt+Q5bksAuucFt1a8sqaZ
SKMCJ4PZLTNGb7gHzvQLI4KyPxzefvHs0Y4sIP7p4sRvY+gQKEcnI3eaMvzsd6gM43/iEc7oYKWK
X32q+ddqskwFiDemapXrZJzzeAA0foHZmZyadJFLPdLTWjx37JEO6g2rmsP8NiphPUebvUALyLFu
j3kLwN5sAal5WTw25F3ElvGatAXH0qq/s3cH8OKueqb6KaH3C5MwiBlQfpHTVXXG1xuFaN8+uQO/
nNfaGizX1Q4eO5KFiE8hIitMupPZIRZ4mXzaRNlrpectFmE9j0mg1fSE60iAoOIC+oqPdvHF+B9B
8Rwd+/arKCLPztyDgxdJswiaZhxDVHu5mxn5GNOIqzqRpMsYsL5/MqOMFKV1bxp3qCo2c2hT3haO
hxMyKVIOLztpmW56WiNzFLRSPEhqpbSVr1OskflIGQWA2RdXQngUTpEnG6U23Bht+tmzaxppv3kz
N5T/ZXeTPOEu/98eqquLHCeb/zMrlzM54PcAnhlEfR1NIvwVukV1248YZFONmf+ea+75nTpNK2rp
tC60OPCaEkBe39eDwMjzHSAptycExLwU/hmcoMoKrPS9NfhPkoHnhUTclanPtI8I7r36PQl+lWkZ
h0oldUnbl911F+WNVrI6RYFBNhmOlY8DIel8w7TnXDpY1PAlwLdre4JtewHds4MtYV1Mt72a0//p
lbVijw7Wvcse80m/lBIXd3G2QB4tuOTuX7jC8P5wWjk/sv0+5kqHNibU94JKVSxSremAJ+g+zYtY
vqOL7K+kE1DGNIsW35ZY0O8utQbrKUiO6Vdg8q9BAredLMzqgDfAuMADYcx+vcIaRmocVz3o/AJt
UZhudIo6d6EmDkiQyz6tQxnohALoVt8COhJouAKxW4zkbOhYvYJJoTwyWbNiUglmodEmj8H/e1uj
JfLV61undaaKStTfYqwxuO2ZAfQT4/RygA33Er4K01wiHwRKlBwZgypw90YhXVc8FxZS1kJLx+yN
6Wz3ufMm7ESGhH86pTo7YqrSIhLZkrGmkQmjWrkEra/TUDkMpzXdGTNMdYXFIW/o9YNihrX4C+wF
BTbyAYgA9QaBs8Ya/qOC2gvXjVG7u1FT6DvSdoIw787g02+A3ABtn2hxYkFVrPADChTDKdgSGTQJ
/7luTodcFXcRRAifqrVB/zUaXQOcknb87z2Usb7qooi/mMNF3/HEXwQBfQIJpQNt0O+wwwGgGhNs
bI3t2yGr4rRDxuBkS/gYdTwoga99nS/1TwNBXWD/OwDtlnTCbz1GTY1gPLg/B3fIk2o2SyUWEHgc
T0Z/PL860ndg3nYKBLdhevxnkCgTtUo+Fz4OWrj9g33JFubre6DxIL+ph1v21zOO4offIQombOKU
raPMLzkXzcv7SopH7mm858nKLkP7t0xSwxNvL5a8OaZi6Jwlu9eWwCmM/K2ga7O/GlUzUBWJq0z+
FBK4Qx3e3X3S7GY9xHJtU8X8CeSCQidlBsKEwk+VN2SrhpOF15b3P2V2H4FfgdqQyNbCrxEgS5Mz
Xt7eFYJ4CmWUoxtpKhVmSHcbZosoVDRqYpmQ4V54oTD8YhVvOuShQ6e/4AbtTeuMBqNWNnHNvfWM
h/oMx504OZqUSnKfxt9cW+W/rmIaBeBIUXcLoS0jvHVirFEWZEcU0WtwBL/SSUwW9qCy6ZpFPdtd
GtjeRdgidUSELn3PaSNwi/LB5KuAXvBDkDP7ImkmpDa/QsMEsYcG+0OS71/hTh/IsHK0LcCol8m1
sdY2ngeoKrXH5miXV7FIRPTuabCZKYiWa7hj33LT+A2NF/EwbjaBrEHqMTo/AFyDpNvF+MRtByqF
nsNP3HF6XLqYmVtoNKue+3i5pQEGReorSdLYax+TOrf+KDnPG+Cok1sMq7PyF1uryMvRu+bmGwmw
jDPsvMXJknrzZ5VquYGR2AnsTcfkEKVAYUaPB8hECKrs3ukmSRSvaLuCZAc/YVB/q5gJIm/0Vc3U
5DKR1GGMf3GvwfDkmEiAldMsnxczMZSAl0bWBaWbl7/BC0WZssSVZ49g/CZM86X7tgv9RWCL28pD
38Bg8g5KOwVCHWdVyGWLprcXGrLf1GwUwDHwkBm52vVijlKNcTwvwf2TGzHQYZ3NV5kNZFQ0V+de
M+Ffl2weOHKvAIIawDnip8yQ2CK/GKOBX+6rfG13/Y1r22q+d6J+DkVhkvJErWHEPDOrn07urriA
ru2dHKUswtY3VRaGrtRwDVUoVdGlUJdIg7A0RWgLzr2u1DqJmzGZ4KSpysdX9LleYkTwOewrkTUN
jpl7g9pBdkkSnVNjl/lqaZnQ4muPjOFGb5cEah5iCDywmSd+BEMZtAdMpnFJriPbvzivvPHisDRU
NCtEZVICayLMPVp9kp1vIffqrdHoMtnwJqK39EJPOX0VBNQc1ISos+zdr1trZLILxJiI2JErg1/w
gyiLpPKmhvtpcKe6IyBnUnD5jASNQex6v8SBQ2Oj8d6q3jDWGWGuw8Zoj1Vn+zcK289sETPr3PhY
zG0KUKaSuSR6t+4R3c8PYWEeJIjD50WkqkDVsB1PP1nHR3xYDWbVYwZD//J4BWyqKy1pVVhjfa8/
l/FP5tH8W1zt/Py6T4bbxT0TLuRHECo473UVEVOwoTF8QmM+VoXeQwgkRoLULf+C1oOby1zXmfdt
2DE7Vk+wc9+bBgpuA1a3iDnvf/TscF200WX5ln/IKZy7GCEI7yveHKqEao+u822SuH2Odc78FM+x
00rPPDiEbU0N/HHqIjWbTYa5vTv30jC+ECUrS3YU8bFb4pbzRmdLd8BhsXUS3uRUdvAx5L5JGLGn
9VlLXQIJhZmRV4G8DM4eGp63IPnz11r1wmRf0+v4PceL5OZjcwlE5PpHUVFV2u2cc6DNwWLd0ZRm
GPfQ/D1atVwMpCo14oNtPOdC5ngDBy5DBhTjHWvTtXONRDcvAYLoGyJPu6drIDXCyiOCMb9hRO0u
qkccPmL9kuM+IxlVSy8EVWU+VH2ZYp7SagEwnNfZzj51AIxz1mOiGEvcT1deomX3FOAXw/nuM/CQ
oJY735bwWZRviTlTWodS1+BrfZ9hmt6+emhjpXl7UyDY5OInwCsz9pwFxGZdu5Z+xYjlASdd6w==
`protect end_protected
