--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
FQ/FfzYnNq83C1wR7yF/cinMLnY+sXJ5U2H+cIl87kV8Vh6vr6BngMtrca8ZagOSq6ez5fk9GwTc
Xy2H9GbOBowjuagv5Mnp5uI34aS95EV/CKzb58oK1I9r4cb4Hiunm8JbiTGcpqA3IZiNvZRaGkgR
RdIITEGLOQmYtwJ8MVFpOruTdbPnLSA5hyEODAAKD7ZGdLhvZcmAXdkDAu7xwi4zTpYpI8R2hNDr
ud8yZkcDRoP395Qh3KFkm1rCToPtD+lKQS1AoHRrOH7JH2CJ/5WGeA/A738FTUt5QaydjzZqtGV3
DpmACGQS2bqFlOwFcIR2R/TTf6N7yPE9T6jFUg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="qndEYjcq3luKVosFzOjczkEHhL3CxQIFuw5rpfDiGXc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
rRrQ2Y2RGAGq5Xe38lZqwufNLMTo3CHdm6sworFMNdMCY9poSGpIxyj+ZD/kPJFgnl1gs810BHez
Gc+I7PYQfjo9tOOLQGKYQfOA5a+ZufonRnYUsvl6LNp1/RZBkarhn7aMa9rzrniPUVJAfbooud+V
/O47KnBZfm36nBsfw7zKZtOoPBX2e9ixVwqU49i4HBmFjQmsai9BTb1/w5dLCtEHVwn9tT3I0vOQ
p/5j1aPZWZC+INT3rUqjAfLWCQoEXeHtyfM00fP83I7hSAKcP1d5Zp1ZZgZqg0nDB2of6SqvtdPj
NR7NxbY5JNov5EXV6ghVkuiAbOlqBaKBBW8a7g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="mb0W+DPHR6D2oZcuAI4AwVI+0aKx/xCc3UzGy2eoSEo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2864)
`protect data_block
eVmDXQVgw1nJnxxSjhtedAjQD8Ny6VaO+dxNKfE3+ISz3wJLFV4OWqC5brELgYHyKP+aCMqWXPxZ
fnQKrJR8X4Sghsed3p76Oh5zJJ4fALNP0o1/QnSs6Q/gqcGyHqGGPuRh+FcqqNzWjstqC7K1byZf
8A6aTfmy4m5UBdlv4DAugcxSRtFyBO5mMio07xgovg1d2I7juohXoM7jNbAFGOVH8bKQJvhF3HzM
K6KI9FsCvAnDYp8fXY0Lw5p/b91vl5AwlcUMKH3dxybasRJn8wsVHyyvPTeW/yJOaXp3XmWJlz4n
BYaa+SN02+Pfa8tuI7bnKw1b/1QG5cVj32hcvQ/eMdFEE+s4dXjfA93jGHLRIWCprumKEYgjYqc6
FKRvZFWWq+ybMB2ptC1NHp8vvj5s0nt8GFEAGx6QfzuENySjJpCLsr7AhIiSSZvNkDXKpIEq76dm
9sYnh2dKLCEuwD6U5Ugw0EvLqUO7gHMszYtO2G4wcG/shqe+PYaR/wJNsdhl+232JjGeurWeve92
MqTqOpSnFmLz4C4P6iYDvqWasDlk3cCQsL0k0eRj+tAiCnb2Git3vdx7szmVtnsQarkd53ncmRLT
GmKc4nnznXCY32A5c7LobofFCbWyftjGifdaPQi/6/b+l8wnmicoCdbu+Co/kzqatQAjR075+f62
FsDyautSZcOushZbQCCWk9n3GtVbWC3AMezR5H31pJwHz1uWbdytsoS0p9xIlY38tkOGmwUxJD9D
AZa+/tYZMUePVoyZ9M1FCQ9RAlnjaJClc6e5CLs9nf4NTJMt4hb6eCR+xWCt+wZ3TceT7T+/IUT7
RE2hMzQpaRz1hK6GsgVPNm2vmcm6rou1qGMfY2V+HS9ANuI3ir1aSCGmaBspQT5KT+iqQ30wlAft
LB+c2bpDXu9SlML5U3ov16QMMuNw3xIdxrDRhpig9/lx1NHMn3Hpxs46uCuvze95Xe8xNObvd6A7
G1j42Qh7wT8aSv8N1pZ/KxgEkZvCd40qwZ/hLPBVZHTbiIkPpj9hSeg48LT+x/9DYaT+owx9aCb0
ncFJTDXdIToF/bIwe2wyqUrX6/mDnjlmRfemwvUYmMEvRX6caK29f1W8JLFyUKnrVCFuwrSGy4g8
CVHsBs113gUGaW2P6eE1eXzoIIs8a6+W6Zp5AoAeCJ1xEbcY3mlCOEwIZ0tci8NDgnuV1Z/Bkk/7
ANsb/c2wxLvaU39aWo0ZABqHQDn2ML0J9mQwVNaPoPw6u+DK+9Vsxh6C3FYs+16cS0ZFiHyyB5r1
4p2SwG8QApfmwINCfPNqF0ml28Cra/NEkhS/tcXpb9/iPPLqwNutcwHhEYNYSAlLUcxc4dPP2KzF
7RtRmrRFEVdhTr7CMYzS1t716LAavsyiuE5wvCZDN/YOJrfOmIc4M9I+vrCLSmqBtV0iPdOr5v0Y
8QBmqgzfy/hIDV3fKUCwdVsel57mjRP9nbTR+YsHx9/8onEVLR72w9uvmaLYZz4cNuXZmi441SWN
DDKh+m2vcaB1xGXmm8BBqB8xbHuC3WGZNV2aXaaLsFqwUImkTkNgebembCl9Dt9oukSGalWzF+jO
5DV+gYMjLZnOGCY8J5nYX976GtMC6X3+o7qCLH8xRGhYLK5Y2H+SCAIsfaPQN3+30inmfsUv24sV
aefOM/fIRa3UOR0VqZXLAN9m1UKZwqvN8U4uW+vFTlYlgMs8BwQOO3TiloZ7H8En7w3Q3m18x8XJ
088NFtn89SK1S+Ajd2inh4E7R3nnYg3csMtdPLQ+zRkpmf/7kQA5cMSy8Db3xS74Hj1VVsXSQmMi
oKW5x7myT/7pVjvtwIIpwtZhrbVohDIIWFHbYt+UPCBoVNDNH3HK6Q3k3VXO5v/fEzj4aYvlFlRL
JBRYdAqrm1pVoeQ9WDb/EWnkriNfwjfj0n7hpTmZFPidKzdYgD7ihcfCfZToFuk64KF0TVF5hM97
duR9ieYriCIRr+ih+3v0CpdxaOv/q/1esuQo7TfrSeSHp4xUz6osxB+l9CGnq9imhW5wp/TL67xH
IlaQJdxUADNDv8ql4jiI26tG7wFFsgNqNdkt0ZB63yNeUknFafGWih/1B053Fhtq1p/0IKVQOxc/
fNHZSLBNHoG5cz6frzDQ0hgp8RIFHBU3nTR97iM2PAEnGPxJpmEBigZtWWjmUNo0uvKFvZTM04w4
W43BKxuhfII5rYFns1BvFa1gAn9uzb8iXxk8rAeimAwyJpqPFdBvbvHhqKImvGZGR7oMbqLwLqOE
VDbIfUheemHb3OnoGuqedtBeE3X9+ujluRcdyOOV0H3D44CdPWJuY8CY2RDb7/CHzrtWfG7fFCRF
YLs5iSTiIPcKqNvqwzL/ntSlLdZIPz69AlYC0sQ+j+wpvr6NUVQTdKarWBLCTrXTLKnX26nnMhf/
bOnNvISOs8TINNuZHvVkkyzDcxm6kOteumacW3paUZ+Xz/Kdq0ZexcOnflfPuiPSgxqnCBdSTlBQ
FgxxeAcY8SXf5lS+yp18y0crEG9ft6J2KsOfzLKsviP0SbU3Uw5VPvyEWMwvxQY3NkUxJWAJKwtR
wGJAAlgkhIK2GDljEyPDZiWDl70Yr6ducq5/bj3FPe0vO18yk7AjkPLUm9JvNyvaKwEXDsQuFeOF
RWZxJ/UHJZFcc0hzEybf1X48M/TAQmyxwOgSFaDfQs2KUFT/0yc2AK1NPL1F4UxMUcHi1a6OUmxZ
M+tFrA+Z2TGL++h4btmugxangxn0km5WRGgCSBDg964nKKVl7oLwoddcfxMdzAPOP554zAmCHDcK
nGrKMRL5TbeliZgGAYbwiIpstIGcAV+WRXAuP4/hwB6gzUAifj5OjLMtqXsBbCM2457ENhfpO94K
6jj4YijSfcq8TneabSWZpqBAdPSDzByWQ72F9QLtxzvZTx5FAFbuZAImJ+pSdmlDHZWqAj3pUeQk
NIEhV0j3bSRUOQyINee3Fds4gEy8YHgy+b3vuTBD/RxwiMESgoZYxFB/Nk3/X4VPkMdbkCNe4Po6
CY37iJksW+/Tv115os1hqtsfRUV8UIIhTc38O4kMAao+EuKbC4d7H9eyYsDVjK8mQKVawjxX4AMo
epWX/0SJ8DU9tf4lqVwIy9dxz9kXyO8Dfyb4v0+/ztZZL0haPecP9xczUWpV2aCCyJMNh6u7x1fe
YrjVIVSSy0fZDF2OACOeNKHYPNTTrpQMQGAJ1OPBL9FoVst3GAEdhy8WuWw0rUHYoI3oDsMWKFs4
90DT0fQ1uhc37HChDQ/ia/3fikcWZ9Sw83rNpSvQH1CSrH5g4QLE/noJygn0vlVsCQKi6vApYkO2
fRVb3mhHxeStOhnKR1ZYEMTuVxgpnFbwWV9Xzz2a3zDa+fAkf2GLOQhgdtlwISrA4atQDBsC0dAc
7mZx4sh0rLEB2Scwhu/N1rEa3km9jyX0REtzKjoA7TboW3b7ejWGM/WRS0S9/gIS5pbi4w/PFjkR
GR3ZGBZIQbn7e6VPueZ/mgrjJswumPjdAflIw5dokHMk2oCNGI8NExZYMRUpzdae+lvIaz5XNbZt
USVtTi+Tciw0/fiXYWED99wpLmejHG+dpPpHAtl9koUEC9O6P0wfqGsrJMI/icLBmZsfsEvIln/s
QX7DBtnKYU59JvIoT1bQcTKq6sXNumTgGIxoBCZ1x+OdPB6rD5wtHYo9r82Rikmfv/kCAo9Ppkdd
GZdmm3Ml0MRV3Bsvhbb6pe4e0mevPnumWOpZfouNScMw+g5j8LRXJAUgdzD+91Ctm3zHpKnKwkGv
/UytchdrzwykxKQLRew=
`protect end_protected
