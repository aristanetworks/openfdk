--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
MzTSECbwwlcrwsJRTx1PD82pmr5xTiMLAeb/VMrhyluGWX8vbq5yNdrbdCO7gsd0O5fMBDcvuhLJ
ekfCjj/+PGImc6xeNQa4P9JYhVlzHoWxeRneXu1ji/rJywN2RpicEk/cO8rhx2ZM01GKPg8O8V6b
UzJD8mmxm16DQC3/zMFTUlwU1P5lzMdVF3itNvYB0r9WsPMxpprUR+YRC1teBcfzP6lld4HwDiN/
Frmjy4zvWAIWE0140JfAcVfR9dltrInCC5o27ayzJkd1x0EnL2u8RmKYtLRHqZKFyd96uyjb9Cyz
fyq3BMiFoJWzLFoBAr9vHEqAABqGm/PF5geeVA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="oB5RDviLz5Br/0GuCUE+R9j8JDwOt3jul78pENGKrNk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
WEiyQI45D2kTUJhirvceZ/ck1vzFX3iHcI+JTem7lSGN4WojLu+WoZAc0Q8WqBdduwjMe69DSK01
ouKfCwG+gR9iRz9Owpe/QTJKunvvEcDQORJ0M8QbNqkzoYWUkYgTMWgKawUCw/Nju0WSvW1a0PhR
hdAlm2CmQIeOe6Vv5V6Q5atGMZoS/XwwWBgUU2RZg4x5EFmfxWdsFG+SuUfAbAxTfgKtDhI483C7
NnqAsM4PJPQG2c/JwaD72NP1IqueOIgECm5Wy0c7crRwVQ5i0VzTfGk/u7syPMtq7mJJDNT/273b
Q191XsAn1RUDg+ry47wUWLewp7FRsIj7l6M05A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="4Q4PxtqTkMca1ZdKMAwh74w/mZ7v2nFefmvlyTfE2XM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10576)
`protect data_block
9pYlYvkVFIib3CEyMBwmysdKhlMrPpTkaZLkekSpo5rxwl706fGNbPpYkDm+0HXTf/5aG+wv/r2A
4LqqAP32AuKmBrL4jQ1pMhyllztqzSeUYY64BJ/IMwpufSx0xlO5iHAZOrJ/+LQcCxeILWWb+whx
9GoBFtYc3Z1H416+SzDPj98O3LG+z8ykcW1nVM7heeTu4TO1giEAnEt2994CNIXiyG1QR/gvNkbo
bMfmldIrxwVY9MNhEkstN8ibnBxjgCccR0iFOAvWs/z4I7+hQe62+DyIggH8qlWAuhCgi2SRKxnE
PfTDD/DvyxgpdWU70jVX7pSO8G/UKCyhf4ZaxCvfhY86/uuj4Fz01d/JizTyqiGauRuQcDZfIQxu
WqCDbtoxExFUqYKwwua6QTWxhEI2tlgXq5x9pBc3klHxTVwHfso6i1p21TYkxM11y+SMxWzWOlTC
CWILcW7iRYJjxX94BLb2CGVQ6E9RshWr6mbaJ7kRuxDz0oAdwMNvwg3he3OWk7KTsOmlDMLx7o2P
yjKkl2U43SIqk5tkFN/msZcGrHNHZmTFRrH5ksQwmbVIeXbm/g80KCKKaKpIcVJLiYFYIre8UHyz
34AMVE3XqTldaxqywo1cr3IDj8MwT8r+hsX8KpujkehtSVBWE5k4gC2wQrtFAwyj/Ck1sPp03X3Q
UrKT2cCHfuOWvSGSSqdXhnwKTM8l6lr9XvkUNMmxBM26BI6XiprjuxPzXYHGw8wZEjUMU7HjmxbM
cFxCPbrdlPPey7TySBdX3kGFX684Mb1kfWreghRCP303I4euGxPrAztiqKxbD6AKGpNTAJ4iSRpY
eSIuTipNbC0t/9ipM+Vfps/VIpFLJg4CI2dAsYAWiBs/czHbctof47IhN3QUT4x3GMrbCQGj5C30
TbC6ODJVxGr949lvxRtlyNR3kwtU052jQtFaERfIk131bOVJ30u2xK+xA3AlJm91aIdjjtgvgvTY
niG1q3fDik0uLfHCT/pHb6YTDgyQRr2VssgAbEXmleNn29p6HDT0gkulFMBrfzmH8YVol/kKDevR
yp4ir6+/KaSMRsWifmH3g2F6HEgbjYpaeLrOd9Yg56omFmNQnV1mUyZ1T5JJTcH28TK86yOLhxKv
VJmNcEyRRlySTUeOBYdtPMYvgLi4AiMS6rbhyAjlKZBAfGuyD290e626I0Wjo8mApYGfXKe+ek2H
uRr7vN17VdaCzGKmzWm2W7cNUgkKVJlrQgkSbIeYZASMOF5SJZkxgef7QQ9SMxbJPZPKnvSgxXN/
zqx7ZAC8FXZnQAimeQML5YQ/9WCNHHnG3PHvD63XcS3hNr6C49Pwg/vHUAY5YHgjdqJmWcsa+59T
yuP9O9krIRb4N+0t/lWqtwdfhupiaiPkVaAY95h0VaOEkjDvhJr1N1KI5cZSAWMp8WtjMIDB5b2y
79vkWWZVMjbplGU8YHVzjesu0RvsfLKiceIiQ30lx7BZn0J2yJ8fQd+QUGofQxOcfdMIohXU+Br3
kJV5cxGQwDl8zDNRpDwJdJmT91qio34HFA4nN0EgzGfcuSiQZhhjG77Z69MInecj9Pler9f/PN/A
czWvAfeSKqBa0S8sMjLghAvPD5WoM7ly3WQLYFqXqQv8YOIa3HMbPuMMdLtxRynZEhRuqtnhlrUa
cSQb4H7Vkb5DzsLtBMoqGJ9/ZSostWUu7w5WuhSc9MZrY87zGKobbF+5qPhwNew3m+15jtqKGmHC
/JVu6rM3ruGFhHoZDmDAa9fzn50CYv1mrFx/gNkzmTtSFinPKBrcCAgazAJTGcTsF07kNeBVgd1P
MMHcwgM4vtFooIU0ZyCtUd8fFPYmqfH0WpC86r0PBPcUpdze/DJSNkHQ+4jN6T95wKuW7d9mhUb0
Z10DVGPj67Q/57ZMXI+NPhilvVYlbNOkAG416shgxo9w89Qs/ppnoqAwwBcTA0s/J5t0gfLtLi20
8f2ujwqP2FbZnB7hRF5rc+KvK6TE/GM/zdGwplepU9lcYqWAeB4aAN0s0LiGGHqlCdj//ew4jNcV
6ettiRTHDyC/1n7aXLr3baG3n8IKs8rvcUOta9x1xvGu11CYzplkLAvlIqPtV+wu002t41HyeGjd
wz5u1UMUYY7SgLEQAo1aqBOG/ZWAv1FV1jKm8EIUP125t/jToRp3PrXi9HI4Rmhe345nAFaRNLuC
dfBS3ZVV5Fht/74vTpJkJjVcmyViHgz07eX0Tcm15pl7dMBAJOPA1ooulidXWR2WGtd7dqeXuP7R
oLL07NWL04csdzNEwxuI7VB/LC4TUp/efw0jmn6GlmQZMm1ABRzDDi3SKSGlaWNeJSsk3kdoFsXE
xAKCgP2i0t0jz4bp9WJcWJhcF86yiKwQ9hEgKJ0Uwyig6AiarUhjy1ZOU51U2L8Sl3UCCl9EfIio
NBwgRoI7DNHSkWPYfDkQipEjQfSbE8ZychbdN46uoudKbACyrula480c9bhAtbZuz4SCto+hi673
tBeh/kPbvFF3KfsQSmzwOVq1t6kf2xrGqjOrX7+b/884VP47sux0A2yNqlropqxTe7IHkQ/NyJBh
GJGhj3pc+0eYdAaW3XHsBIMGX5uhPDlP81/2fmiBvBx/0kybEYEGPk3f2jG2EMB/IcEVORmNz0BP
nSe98i1925U7g0c2Yd8ZVGzmNcPwxWm44hcOEDSVptOORHO87c+StMkRnjcijHjzSfz2J76Ul3et
dl1wXygWNAyGZzDZux6iadNf7FMCi8yOLzUG5fvyOd5M6Zy3J5JK6R8Kbvo9BzzuDeDZMM0Xr/QO
6W5fzYsfmV/dxKMXfd8GC28TvxFf/BDTqS9OHruwR1uhp7SX0pewU0pQywIGgafVHYXJROX8TXhq
pHXgoIBl8U1Dhk3gZlR+AQNeItNU3lEYaC6yTl4LI4+YDhx4B1xMQI85WvIPPaRrjJNRZYlvI34A
1yycXsuRI4keu43goofnT8De71JZocQ7EWErj4bokrRcsSWF3WHkBlUxC2nBxZi2TVJkl1CRtLMm
TYG+cAk4eLtpsJLmAmYk6Z17f/TaLVazXxRW48fGHvgb9cxqAVZ0ExwRIbcDFF5zbXziOaVM+COd
hrtiDvq23aX1kXQQdL8qUepVaWrrANbSPyYNhix5J/v3R0uZgWXLSDUqEa1JgQZIqESVplJ2bU68
HicPmrDq6KZ7hRJfybH2fMKT8xpqfRD1HUOhO0H8N9PnbAXfLmPEQnEb/KKlANsChCn+LJSpY5UP
W7fm00ILRRzNP+lr61RQdMyGAVcXLm62OePERNySq6vfefVLpkCj7JstBH4SuWfw7km+zGlyNZRJ
XNNwIL8e+GDJ+CNCj9PGAl+e4x/7+hGG3gt9BDSfAlnaWoHtPJvWOYFY2vcr04uY8j4DL38yuqT0
vGeMkd0wT9S6LaKkSNgf5O5+SaPZAUsahV4P4n+69jd881vvqgbkKtBpGBvMEyt4ExjA8rJKmLQj
Dw/Om+tJdcunDtpVvciRlYvC6AOsZ6rCEg1xabSFRtgYW7fn8JESvt9g9zjQeMeeo98nUBdYxHIP
mbrqi8kWQYVKkUkbaCeAl1dQcpvrAkt9SYLednjMLc71KsW/QoGgjK+MEuS7wccRSmoKXGTGikhy
NJz5XnuDBKEV9xSqYMuGHE0PIEOi0cYjC213OzJbYLkLZrQw8jdBR8WkZfAeBTU9a0OgLtD0Abi/
zSjOlLGdDsq+o/b1sqZGuMtygVWBDnhEIV/Tx49jkfrpmc4Q0KXC+SUTgNsGreoFLxj4ZY4ocyFy
XM5XiW6Dq13yNMYDTto5mD7GY1FGPzTc6vmraqJqnMV266ECLxMv8FuiTcLtoQjsDhkL8JiMebcm
9vbfUVWQipbT2N3G2TJ+/da370EZJkTyj+RdWvzbeFOMWVCyJJH/frzdyIpKw7/eZWFQsfJz/tbu
aIUjkiCqnqRgl1kP+RMQ7rp9VCI26sv0kECX1QnY6u4eDlu3rrWzaqPp0vYHWON11VKJYHwU5AsG
6EiToW1LXUf5vzpEgHKIKJd7rArO0yTYzXNhWyiskmhGIhoRmN7G1lO4kY1NfiEbJHoW2el4BeGG
SHoE2W+ZO/NMFcahDUT7wsND0tv3hfqPZsFCGU5IDY5nmtv6dzvUQ5ofgnE8PCQGPiLIjijG+wPe
WmCyzn8YmI9rDLNmZuHReGBka1haAUT3HCizLdkVznLhjfYKVGSBgIsPdE9ZDAPqHwFTOXPs+OQj
3Q2Yby5sKhA9M3TOayR3ZGGEtsMaw85fN2MrBeJAQ8PkSjzOqz3V3BIkxHQ4v9PvgF9ZlIJdRX8s
6Ar77O9/ZXgbO/CF0bohmgqH5bdaAxcNLHMWJLQEC9QStrrUbc+hZiSaiIp/WUmflOeGuc9R9eFV
u64W5tgeVAPfG63PHg5ZJVgNugAsUWe2i8HRcC1qocd+wPcVUBZZxjimly3mcbnYldo7C7wL0jEO
/H7NMIn5uJaI5MwrlL+GNyfyJ0uYEECkqWUSendtS26Gt65zEp0MRlc4ZJAatOPtmLXo7CZuVeeh
Za0pfO/Oi44nOTm/xGRVqO3wMiZhuQfWNB/4bbUoIpCo2udtVoy9L3OdyXxwvzMGDt64AG93M37c
Qzr4QAnH5zxTPsX/B+tRLjdQEFaMsKMC12TY/L/itXVkBZcWJHY4hRVaiqKFL7KTvVycp2I2HMyp
QQHLXBWZ8kfbcsPEggAl+ZsQf6VjbGPkEWUCxJ9BPfsLhO/ROUQIYHS2shAvJ1DkvyX2fZ/d774n
jGX0eDEWhGZTMy+XtrNnntN+GN+XGbj8J949KdWXO3VgVYhtUTlyJkTTAW4uzDmWVCUeqvBaSg2U
5JIg7wPSJQC5wnKE6IE6fJsGuAQHwrESZvg/cxhcp9LP6EUB4iDhoJXaDL2neR9tewwq8/jnUwY+
RS3Go9QPUVppWUSSpQahrYHnfYnDZHrJQHW0mq6IuZ0kcNwHOkBzH1TYnsuNIyytyyVLq4MKk6Ty
FctSK4COVOyIgrVgVsF9hWvKKd+QOiHSyPiK9KYtmrKDcPkOTsd7cypdbbgisaB6oFgZhdTSQdTF
MicAWGvR4i0gN8tmEEJQqslntAnYObJAlMeL6H5TiIGRd/IXDsfilUN/To3UgjVnbNKB5xHO1S5U
KUeGKfyHB8l0BTWj9cKqxV4TODmsj8oW5mgr3KWPBgNryrAM0Zonn1Sg6b5mEeBp/qnmYeEbw6/8
GUty+rrsY2s3za/rTpF3cu00Jk0KL3Fz5D9KzLQup75UV1JqSDZ7r7IGG2qjlA/tJ+HRt/RdAOOW
klDsAh2FMmYGnLh50FCFPT0c52atu77PC+foXUoDmj3a/sUlExhC+cjGXmRnt7vwO6lpoUl2EAwL
Huvzztqr0hgzkMpt11FPe6a93yMx0vDj3tjDxc4PplRg0AK6IjmHk15BwrwJjWp2xzsK52arL2W8
MJ9ysUIq+9DYb8IS28cnE3auCKr+eYq616hDrOwM8vOf7GqFn7xsQ4ZZcnwKxe7emp1gfTR0aV0G
BsDyvEnCS0xBKxeAkQNJRcYEpjWNumjRCCQ/puXwZL08LXV4VWpwefv+iY0rusmAmrebRh2B/vtq
3DyU+zHpwjNTsH2McYywb5ZhG0FLos0rvsWEDH01Jmr/4Z24SOUVtUtCe/Ew8KecdgaJhGZ07iVP
N1i52IBgIOSRqKclcGKKe8IHdLRPdjfdHSC/1MeZGbGF3X7Br6scleu6WNnWj6hmlHbst0fpo5MI
nhjcgtaxAJqu4RNzxZBSCOepBl4+H1uVXezCrRo8hH/b1qcSMJ5lZeY1rgXOjhnKXMhuNchmTxGF
V8I2wbPmuIZpezylvBjPFez4sUmTjdbnmdfs5TTjJ3GdKC3xhpGZIOOw217PnMy5dlARiEJqXd2N
HEsYhKM1Hy5GCoiyYsznVHDKeiAWGpb80gfmJoFsBHxBptqgj1nYsszo1fPwUOEhJMmtU30+Fajy
fSVmslbfD/LJSexwu8XApnr2Te4pGbzcnitFz7ltr7Pq9o04xHjMrDMgQ15ms4XSrPb2lI+5VF0n
HgYDx4pji7ZV9aMbfVresrY72BVMNzF2k//y332ELj00DZRZfYymNUn4C1D1tsRrLXjvdKk4b5Cu
vDAHGKOrEOvrSNXmLJrciYtn7SKgJPW+DFAxN7yCnyBS8+6UGPei0a6Js18UPCKh9PFOlbjQzMXw
kvKiBNn3FIMPcJPZ8eP4WKDBHX8zJR+2LuPlT9UQ0se/x3kufOiCwYzNJPciDGseifyXUIzygPnG
St4X63CXNR56ZT3OcSjhv/U3LZ21Xt7WZfopYlWsX8qdkAr5DKGe9ZWdqUdzDShFB4KlCzvTnq9r
YPrWgdW77n3x5EDeZUJ3cmEZVUF9KhbN/HkHmDjEvrOgY+i7RysFq96zrnAv0WAlT9D+bIDn8Lq+
bQJeKASp1X9fv6CmXOw/ZX7NMX15X6akqj1lWsn78HlujPQ4pCYvzg1Aoe0T6jEQ9TIpLwf4Ehb8
KdfomJtLsNs7CrN+Cg0BoukreslY55yAxMrJ998LucQTrVeWE14Yy73eMQczc3TmKGVP9QN3kkaE
hUF4Ul63lYFu/nfUlzzUrFaN9ETY4bpt0N8jXs8gWiY/4SEubDHnkpcc4lJqToSF/ksRKYIf2X4j
lx5WhSrRkndNNFVMczZeAPSRwv5nvqsMEnpqEKM77gIFz9F7RigtYhcTwWMMLVGK1ML5hUP9kOsX
6g6CWxWLgcduCKMsdZmCscIuorXzERbjXdI4fg5iLEbnu6lyoa0VGjvxbiO5JMSRys0StHMBgP+P
aM8dsyFugzN5HuDA1CzQQRqRziIA360Fjtl9BAxdkDN1xVKcoJRY7hSUxMapTQzcVQEtYvtywVaB
Y7Y5vdirt/gMgrNP1a6qQGeNaWpHuIJ3uZZAjZgJg4Dtgh+RHS0hC9gQ42TEHYA+SlIGA5Z0D5SD
kqSX1gDcn0HMsl8I1iPZLZk7xmUrqK9BZmh0ARFC07jS/3n2rtGa39moyxz9p2j4l9AAVBIAq1R/
2VI/g2RQ8J7paddJIQf0E18cxxHfPiAknjHap8Mv4JK7RRGd6MNYc4rb4FvecQu2DrJcCnsh78kW
Jq40l8JytjarLK93VdBtsfuuHyqA7F2jWkIvUpTs3BRfG/ZW+B+YFmcugmrVvJtuBkS/Z5DSkZLm
Ig6MMXXJGVLe3RC2VuDSXWyTws6dmv3N2Jcqyp8VLlCHWkIASb8VkJXjcfqaFSD+9anWQoTnrFiD
XhLjKTttMMHSC/KGOgsf9i0ScO+VD9WpDTZx1/+3c4LFk4e2F88nACoCMiLgVsxx5p2YGvZD4IRM
e8UdAKP1vvDlQoZpn5x8hbZIVrQHg670bXAHznO6UbyZBVm4efScDLd948RA8OARbojVc7Ud53YG
Wckfngucj3aL5P3kV02Vo/iKBWRm1uC+0/qjj0gO8HokTMWhvroIXlF3EFRTmxSaWXvpKBH2Ne6t
g7z/F5ykZrK7lRQy8d34pFQfZvNHtDXj33ZNofJx6xb/tQtNQzjlMVDLVhoSmGVn3CkcmAdJJEkP
wUix7excIWzesuZYf5O1WhIRm1Bg612+oLcx2SoD7pWoBpNJ1AGYMRJJLVOscgMTfJE5NbGWxYOU
jzQd0JwzTBSKWc33bnIsYvMFEGe+SBSjruHVhBjE04iFqT5UGIDzXBfUPP9Cmk//G2s+H2CXh8qR
oObXtaBkK/jjmkopBuTWWzO5fRQlEiV9oYnhOc8xYUfq+JVbe822tTDpsC1sUpaIx/Rgpfbb+IGk
izeTLWMgQovJ2fK80WjJi3IzItrs8DNIQlrAYai+R+mEK+KIjixXXPb+emfi0Er6oJlDTRGdpIgk
wjvcUL1L0pxjbVfZShcmp739T7am7p1DyTfqevJuBh2DDI/fN48jIg7BhWZbZzQ2EojLutikXZpd
Zich8KpRc0090BK/6dmgWwradBMX+6V4C5YU13YGA8MCtc0ndM0uFN2k6mxDnOaja+O2Ucb7W4dk
HA2Q04OHweSvJ7tGq513egM8YyePS89xfqoQx4LX0VrQAfmb3tsvnPGwU8yhFddb09z2osd4jwdu
Csm9NuWq/WlhxBMUDzhM9XXUovCs4Z3LsKxua6BCTY7JbZOex9ZgBHWD50sObuArN5mFP3t2IiVF
ltYuwRWoRIWItuTlnPm0SP2CNq6o7D7Cmo67ANR+DiG6jsWa84dDfJwmNlJHzdxTcXIXO4HH3UMD
oN3vI4NN4qGKf0IPZQ2mvULD1Aq0T0HFiz1U4P3Boe5gMNpQPhighlXN0Wkr9w74f2vjp625s0ty
cKpUdJqKHvZ7Cc033iyjJB1RM1k71MFqAbMF22OR+u6iN8enenjXN60ZaRDcaSrCYAqsz0qu0tBo
zbhRP48Mah6xxaXVQN1dLAIfL+SCoLaNJ+XuyFevpcJqsyomYDsFEmV2v7O4tvlr/E3nWTyGulcP
fF5XyTO85i3mVFp+itLAaLlM75Xa4GW3HNcAkRfWNM2b60gJEHAa03KaT6qaDRP4Q1NwMuvoTjsc
ULiZh5J/B4Ptzwl5rhIRXrynh8PAG7vEz116R0RQzMqhHdEqn1PpiHzED+n0+iMGx+b9j7FUQPqs
m9aP3PrcN6ItTPJTON0pygvhBQwFJz9O7VYxQmBd+FO0BmHq8i/VvKC9er2zsfq/g+YWEmW6m5en
Z9tTLfOcAGR7AvY+bE0PiJyQPKwg0G1OC2+8AuvdYDI12/zopL19c7ijJaEPNT6ukJ8yq66ZAN7g
BMbFm1LzUWe25b1t74HnuIcn+RaqsB/5lTGPJO78++mTUW/GqX5a44zFS9owX7s3G8YSbw1mYKT0
GiA+D1BalgEUQDn+xktr0XRwv4q/06WgoxmDmn04uaeFMXfyIQ/jHI4AbTm62vNYCwQoDfIGG92a
JtXuLkrTT42P2Zgy5R506S2TxNszscvjnHSmKuns/T6qINixlYE35ozTwkM+QEIH0yAtm6O8OXXV
oSjRZ6YaOlRC8vY1tZD09pvCrKMUUQkGSProYj1LwnYAl+do8xPjUebRByWevInl2xz3xysGY3+5
djEeaX0/1wYVIs7cHq3J3MPNM/38F5vlANDX+sVd/EmxOvjJSOuit2vllS6OmMrjCc4DQElnxcRh
jYu5dqmGpG17eaLagxlgBHYNlnctO96f7hb8FjS/rHxKBkwiCpW/L0g40TwDYXqHHHuluIbfVNVe
REubb+I+TUbb0Z/5YiFNKoktWR3f2vwKTEFlrb937buJUJtwelcc3jCsCVpbN5fjGOYW9VbMQIju
NKz1QmVi0vAOG660f2d7IQijeZ5EXHcImkQmDgggegpGRH5qOp3yC6KEShStjogg8eS69PjDDUJL
F+D8gxSccS2uk2rue+Rt8+sodiZ9S+v4t2kxvvaBp9fqBfOdPuPvkfdvU74IctU61YgdHnvIPm8C
A+hrxK+4ZGBOp0vT4wzPqxVXrAiE+6/wZjv09vjLfbAdr78hijfdXvyAI0GqmPYZvcGH0q+3RHZg
wLru2UAZDl/q+tf1gUHnjxMECACYxf+F6njExG90Y8hz9kDxZrw2NDVbwPuYoEs7L8lT3nUkrWSA
aYF+6Z7HPcZvDGPAq/zZ4r34+xwOCJqtZLlc2XWbA92XFjNp4vHGECZc2H5IRilQzf+8Q/mOo3vF
KyksDJ5t6gj0YoErOl0PihdQgQBIqTsSvNY6cqlPlo6JMl+HqL3DFeAEoIigyKuw9+rMg5Ct0Lkb
pSJ5Yqe1itk/ZmcxssbVMFpwSgSF3rPtDC2B9xplreO3JyOJvjkMTrZ7s7QWpPsI24HLkXbnByX1
kOHz7NElQvnvdLzv7kBxqQMqfzZRY12QtQOMrkzqBTvzE4onQ6OcNe3Za2gGu/5Oo4aREgCTlpYD
aqAY5b4kZgExPNFOqk6GqIKXKlcjn46GMr2SwTH8lLj43PD9O5DWY2snw2mhL7WG8XfORAho4sKl
j1qbx0tQji6UNV6r1Tcka/fPft2AFkQ6enhG9gN8tLp7OXmJMN0CNR72qmgfAF3DjS72wJafoTOP
ILH197tek4VDyquCptydpD13CKD09oZKPqevYVkzDIx6OHNFYMB9mkAikZ8jpEt7nvbSXe3sZdJm
1mL06fDZVXifILEcQwzxTIys7Kwj+nzQXGHNtg4fAga83MmRXt8AxUA34S99G94pXNA31XJ20DcA
997Wv35DeGoCZ6xNdpAcKjPu9aIIm+kVSTHG1fw+3hkGIKTPlBhD4+QyhTWFmR+wyo1hjNETZP10
/IkwjwslhHhDRxxVPAHCQPpLEq07MCugl1jrsCn5cFcW6zd8vofc1E9+WxMJ68yYPd0NJuCX2NBE
9HStTco7xgw29oR2D3jWICDsji5zh+Z4Dr6kEDc5UepIZ/Bpo/lYFsV3HEtmeykFcQtj5W3RzqG3
V83F2qh9V4gZAJGcbJg2onLFSso9mfJ1WWvJPma72gR5OgCwrc5oikVouywp6IHma59qk6+xpQx8
qx4rk+kWUelSce0W0RO1+9HluJ6ED94ELMMgEU9nirmXGhNFtz0X4QZuRN68D1s0pE25X9D7y6y9
vKKv+hJBvKHxHETokawKgEi+wwOBBXrZ1Y3M1QjaNdOcHIRnmaH86c6nAkvdFl2vImX16FF8VKoO
xiLpIG5OOx7EXylZzupAfMzWeBZ45wgWmGbXDDSBeqgUZtWt3+IV4LzJw+12h7QqAbdSXJXAF39r
f3nriJxKl0PoV/81tKdGaWjAHOzy7HHYKKZu6FbP5WXOCh3sAPshSfyGB2IWcsnb8YzVs2l+OkNm
Blzpz9wxF4Knz3Yk+Q3BX1BBjPpkkcQ66pK8DVj+CoSh+Sdq5vWhvaFDJW/HCkRkcL2jgTVSLEio
nhL0OzaBPuYrm0zuSiK+w0mmceZkflOkOYnnkhhjXgCByfw76chX3uh+RmSQP+5CovNoqyMKdLDD
dIef2V2dTTJhrlBMxaWgUA6ZjtLP26X8bQATOmtX21sRyW82keZnSPONni5EuWxaj9yK+015erCW
6yok6J6HAICDnAgQ37YnlE/MXyNzAQUIdp/aYIpZ4VMUUPL/ntI+SU3GzWhUm34NA42PBR6yJSm2
/bIxUcXDbnFqNF+XVi7wIBu1FTzRF95K6VqgAcFnjb3wNl5ojqug+sLCXRWNW5xGrKgcktPwIXV6
KNz833b9xEnyYGQCbCdaAWQzUzxaiuv7SrEPEvSMLo57RgDVRM8pc94KD6OLUs9rFVDc8uRuMQqK
kKXjBYmeX9y7JY1QLYRE7NUO59tpBaNe4tU6aICaaQy/v9yuLHCipZwLSYk8TSvR+VM0K+EACgek
qbm7P0LR8/OFLZ3ViknSY9GgI06qGbDa5RUfA3+iUdo5wMtoCWJ4R5G+nxS2O6ORG/c4F4XqASjp
iJScqxQcf3HONRWv+9DH6Ra4TnDLTUDhTXKLlM4cDH9XGaDLAMFt/e25rBpuGfG2Zu3Q8kc3ypiw
97M2h198bk1ua56Rc8gkmC2nWeGT8IjlQmwIFItZYJPwPilRqroaVf5H2JxbBTa/Ww4/VjHlfbOJ
e0hoyX5BUjTeGLemIpgdw1TNS4pGU06GXmMert68OmozJscGDAld6YbEEqS5MkY71qo8HsKwdJkD
BLf+MrqJAP9oT+LQmq0d9k1jdSVdcf5gONeKM2J/C84uLnPIXcIwVic3410bppOuR4McJd3QC3XM
Adf8uNWFQHr+y31mexLqhALzFYk/h0Gg2xVGOqng2Dfv0zaad8XsZNYc2fD14S3m1Xtn9/hd7q3O
A6LqET3pRTFR2A9N8m6Ve74IBWDxNE2W0Nvcfq562qrky/Q+o9uWBT6em3ri/9WXkfZOw624RJQI
ZQFaSxMQVA8W+Ga8u4yvBF+0q5vw+DGkX6aTSk+roRVc1F//hNJb/MQ+gY2lypPq9+eKneCNrBFX
UvqL08bcLAZUQAuUOmOG3po0W4YcZYkCoXTuHzOvp0zbIUsreKuyakeminZjIu5lQ29FHDW//056
113T1hU7sI/wOye85TtFa8thVmUYK9YQh1p4FRcIqK0cDyBV99zGaXA6ntIxqcUklvl0gZ/FWmOQ
a6iiKUBIhTbjDiRMsU4VfJGlqi3ZoekYPP5j373fCQ/BnPuic8p6uJYphnkaa8OzOQcIKRa5iEAE
qtyiKVCd/Txs/a2IgNhYt6a4XIrISLW37z3eP7+d2USlt4ZSIiyfs31GmlARj3cor+mucFT9q+eC
GTg9dxYzZSYg/j54fwXZIeis4snduWS018Cjp3TSg/nuGeQzEX1/Zz9q2IepdViaoScdTHQzcQ+u
zpgL5mjTrU/Goriv8H8YRmM0mWO5WiprQKXYyU3girthRrL8lf/GQb4eBs2RzbD5vn00E9ay0GVp
Mpy2WuerYwp3ZnsoQ53mZ4ZZxu+TaLC+H6m5rU8A9ewtkceGKgjbB5e9Tm0jxzkUlbV8i3dtpXS/
cMBVQFSHL9TwH9kRk+4sS/xewNqy9y8dTIqpANk9a/GykNGWjx8+arx5Ye7TN+QonLmEF9wt/4X5
wjODjxnbNsJiZu1qDQYaDuZIPFJj3egl299HEpEBIBPZ2hbBqplmJVNQdb+XkVgfzteLXrnSArbg
ySIG/AcBPveqHxbR2G8xR80V4o0Fdhm8OHMKAmyVjJ/yABsTN2SzjhwEtnnf5+Fe2QxGNz3M3XdB
VUEu29BfwH6Y6O+yHThfHuK4LheuiGSjCekAQMGS+o9Pjj3wmqucTO7OY09qkRbA7l8wZOPAYmlp
yNchDaATyZcqSNQn52gToK0tjZKvBqyahEW19Ev9Ymk3B5wDjmQeG1yLdwT0YAgOq4SDfb49DNZk
p2pvhidb2XS3gIY6LHDliOkM0s/H4dCYWXMj2D87DXm58Q8q/wTE+wXzLQffM1G+7IbJzVS6tR26
wcIz9e4FA/VuzvTJXbSjtLfoCTKg5c4DbIsQAvQ6NSAFIHLIL1EMwJM7fKMejUyJ4tg7BVLfyoDQ
99s+280txV92H95PgHDv/d5LQD30081GLREsG2L2WaxfYO9dF6JUAOgKe1yiBuHTyXWwGHofzg1w
j73HYFmOQgcCvOotR+UyRkbjPcgyI+lBMB2xnjShb9YDua5hWvUTbuDlQv+nOifu90ZgJNsJgrJ1
IYoKLKEsCKzntG+5Xny5Z94Dab+L55tShp4Mg6056wMZXL8FABZ34wosKnw1O4r68jP4u8yfjQTL
iTahJZSY8eJtDAeu/oBj++zGL5QIj/qukS72pZllHS3JAOPwyLXXlqsz3FiP3Wgf1eujLoM9LD+v
L3bJgsHClUUW3gVTGLRX0JDpbj+BT9vxsLKWh7TUAqxuOskYbJs//xFAAPIdzFUHQRMWcU2lLXxi
7SRll/BDM66aOHXHA/BZLeTUnoo0v+XHy0vj/osEvVIAsz9iW8bh12HTt/UIcxwlMjGHKoCPjIuu
bMA1zobP9OhTNlujGygfiE2WxSoot+NePobn0al3IN4ehqIyoQEja/uJtAHG72AUuoQaHtXnKixd
6rWUg5RAZNH8asqjsPkNn36w85kg9g5/mOVpJ70OSizrZxu/WKXwx14evBcc2PF3xDADi3QLsRBh
AXLASm2UWVYnVeU8jw6SbRzi88B+8iu+02K7xmrEhfegVD9NKfUnxw/Efzjvn9EG3EI3Dt+WleXx
9db6T+JCUVOcIIrsvF1ps5SoXzZtcrXT/wUcbDurmDY14122mFaEU4mK4hil/UE6R7ofiiXcuKav
Zn95NxJSmPTD0PEpHj4r81+IxpKuV6OYXHDtYBOqzl2At/4c4VfvjJfLBxYyBmMPN9FMuTvVE94R
N0M/D2gp8R+tBzZjLyahvWC44BbfjxwzG2F3730gwKlvy5Ij2p1WvnGdKkR3XhOOYG1gUzg0prj9
q3XE3x5bBNouporCFX86w1l0C3+eqsAJgMx9qNvWtwUsYB26KEP2e73a4YBu4x/uBmM6Luv50xyo
3aSCUN9tbT2exgyPO9gLQ1x7oE0GTBJtRzDYUF8hMg==
`protect end_protected
