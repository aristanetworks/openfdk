--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
VZ8lcQoYBWYCFQAbzacAI8PVagNgzX899VYB+Kqb3Iu5pukoQMQUK3Fl1QkvgBXX690eS38JEqhp
cexALgAT0P5ok4d7i4iOL6qhAprlZN4isMM8ipEM8KS5cIsv3s+eoydJY+92O81QZqS4MFJYTnKb
lrObvg0lrZ+O/EYEzqqBWUxCR6QC7it8tZrcKO6dsgRPpUvsUdgiyvzYwltMW9VBdIB2nCXQ3fus
/SNNCta3V8ZE0SKxW7J1ZhjQ/p+lpfJn3OidYgVM4v58YWZARjludq+KeJHZG0bcOqm/8xpvX8TF
KYasgk5hxgDxljg+gpAvBz7TNocrW2Qm5L64DQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="DuCTUxNrmOsja/0qMmYoAGbq7L3WGI5sdiaHazPletQ="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
Ipjb0FV4DcJ3GE++s+qs2nImSF4xq/gCQX+3QwK7EO13dnGNGbMUZ4Rl6DhiK2LlckyActhV1R57
f1YYZuPr4/lqB/srMFsIhbK6DO53PYRkk9cwelk7WfispK3wtOmCxmVa4MMlcFkLMtS94csMZakS
5LyMUSJLhNDKSxUmX4jZn41Br8Rf5/hP59bx4E0Yjho/EjFqv55SBUgYQChSifTsYSBwJ3hu6DPw
9YbLZ/l70QCovEyRnBO2g4UvKuqHCbyUjKHHu9l051jL+5kgjeZJqRfm9vrithFwXFjR9vS7rzzN
dMhrVoS+pAy/o/3RnOP/2rG1jByXZcbSbu0I4g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="/1roFi/1H1jnpeK6I+X8ItxZwUfYmh1RH9Sl+pvCEtk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6080)
`protect data_block
l/vkjPHE9feTsk4QEwP34kmP/L4oHfoKzqtJOXD7+mpYy4vYGvERndlXlUkmWME03mOQ2+QoL5Dk
+lsF69KUkdHr976b8KeGAfUIy+37tgGhwyeBHqcS0AOgU6UzsUn6XA1oZgQMTzKHZ5NuQRNzzIMp
Tbu/VSyId5x4X80K85mXTEM5blNNYYpqmE/JUFNwH3ox2l8A1Pnp/Mqh0XJN1kb/3pWRmhDFz859
/rhLLmGLx7F5liPPDPX44vGba39CmfpHD50TVphSu8P5fE/z5P8NHs7wRGMtQONz5CUXbEYtMtuX
PAjJSoZc0mbb12/5+D+FRkrPYK42ZW/guEAnpoDf7OaXOtAz0+T5FEW7s6nBW+hGP8x9OAW4YZRs
nqzumcULQoqwlWPM86jXfDrnc8p7KrNpqKJR+2YIBpyaOEJW4KyqBOvR3Iwn8dp1wNg9NEsArhl3
9BDM5QbTxVYEUMQiJrqfTlx2xVLu6dzEYpf2IWdBNqkFpTYEIU0PwdiA2C8g01porJskE28kAKJS
lsaH1wziu9peQLpttnRlGA/VF1aMx62Zz0Gn90fZEt/BMr9iiWB2uwT/kiuma3se5moD3dfVyD64
lx7xBWDKPT6RhTuambmjlea4aShTW6speY/oKS/9w0d3DOd84zEYlJ8+tIL6OO3m3cYDkgjxiA5M
aTZE6DvnKLYJQHMyIpnYHYbj64QYABtA3BbZTWsFRsVRel7ocwGaa5U/A1c6ScJU50ktTzGSSqa6
vuokuGugkDXbJibQJH9Wydi116oKUA1UB/9vkuKvKyvO0B050jw9XUlINTCdNcKOdoDqLf50GPJF
Bkj0HndeWAygNKNnPi+LFVt2/Reh1yO1CfDHNEPGe4FeKpg0DFXE+mjBbkzL5IezQfG2xb6BUQRE
YzLWsCfthc7M/60Pxpt+kq3hSb5L26a+WDg/XWnxhBK3yBVU/TL8RdD4j7fF3m8wEgjAKyqHIEs8
M9Ez9P9oZUO62VIUVB9JCUsrcfG6IeE5ylVXrnQTLUoBzsjWbZx89Up+m41aYc7KpmLxrxn5SuGQ
AizylN3yqC4/gRzp9ocLKd14XNS+x7XmCPMKTw/4eLIrbtAUtY++P+COZD8WeEnJUB1AbUcK5tot
aKkmQ2c8VnC8TKG3VvXOrUnvIXo4IbCfB85OsDvCQZCw3j9Vl9l4hz7d9apl8JKzhdMapLjQkP26
NDgy+6/+I9hNoBwB0RgfMmRozmPVHXQjqMvl50Yeb2ceWWdpsH32WMIWE4aGQAJWe5IhlF3PBsac
EGIDK//XAJRONMOLz3Hj8SSwTO0gQ92XtqG5fXsUtyB7hck6ghM/6kQ6DNLmKlWkhK8QgkiIxDDy
vUqdJcxUycgQ8VYUfX/vOxOHI3OIwKpxeCU0UxWSL1vuIMBYHIdLkmC6TBgw09KWMv3uomn7aBXe
WmamESbT+2DATxMnFApkmCdnWaYmMppykAHCz2pvggKY2LTVUi3VLBaCTgy0VO0/np5ZKdVMR+MT
UyrAKcy8UaItz9Hy61x45bZNyEylIvWyvgD45DNeaApuuNtXGvN9f6/yAgmK6UgxioFxdnPtdHB9
b+gS17gL+CokP15c2+0fqF/LIlfQqxEvAjIVqIop0zBrVnE9xZgAlFCsQ/1S2ta/P8t+uCZ7024R
Ql0/WhYwx2QfG+3FaoOYchfzl5a71YtbDUI8sVmgw1VmKZdGB5vByfZZVD2IUqik2uI7BkVrE1u6
4c5vlrqxEvwcHuNm6So5XC5yI4Rz+JnkjIgMt2bRPBCS15Si+Fz5nTTbXPfMZEuTSwaScIZu1qgx
+yl6uecpjnueXAy1xeFCIBeu47Ik+8hIlTCB32gAJdMTk+2mUf/8f1puh+hcDNzjpPWI+vfgiFSZ
N4XycDVr+3D30Sc1RFqzzbhjIxZOfi4IRC0EleVEtxoeTBArwH9H8txf4sZHyNt7wEFleMMHs1oJ
Dq4lu5v6WSfYvtcZuJ/ubq/PSSUtO6wjPKgu2jSjwIdqZ/bYvPyFiWvvWU4Yr1egKEX4UEGaolxh
GU2ZZJtAPrD+JCt+DhRLqMkHwPd2ne/bI78v13hzVGL5mRLZtW9iW1FVf5a0TCJ0LrYPOBjAeZs3
v/KaL+fNG185D4s/xHnGLY+hjvD8G+d/2AUY7FDujbseL6h2aakurH0DwU/zT1Vkxs+7yTZMFNzT
nEVnS4+B1HLqluUvT3hzVbXyTYYCAZhB1VZqVsPubQZOpqd3KC6Z4pcgM0rEu5SL9c1ArNeYBKf3
fIQReAk+ENkVKubqQ4kiewvwCv5a2Uv1Ys7Ss/eTOBkz2D30u3LhSetmF/fm9k+z14xJtjBPD4Go
V9uUOBHT9hNJtM7fM7FBirm6Hilvo8b4krm542+912KIEen7/5xEPHIC7V+QnCE108UFthl5KRC3
0qbwRZQ2iWb/4HEHTgDz4hW0Gz6urUBbE983OM1594yRFJpbuLm0aRhvZrpnkLD+CqgsmTIN++Ju
hysWYPSQTrdRMQOeUcWJa/hu4GD7Qn54CJOCgLpW7ZUPiFXyO2q5el18ceA5n8bI/SdXyekM6LnT
U2JtOnHhqNAJWG6qDZBuCPb6Wv7z5uG5rEfz73SccR0mos7rwYjja08Wj2iFXP/g6lPh9rUiADym
/XCuNrN9iNqPvSF6W7+AtShyeFQb9nZYBkmcoiQ3hz/43kxtlzUjRNUd7fGi6lgJZ+0wpX1aWXMa
YfPBWtUke8O13KD6GRoQYxq4d0bbLSgoj9beA5ES3OG3gzu87T6HpLLHnhD2cGnu+TC3iPw0xjSO
zifJsH7lWFlpBqKi9bh6EBVZ80fNrLQfqaEt+bRNwH6fWoa+Bqlst+mZc551YJApk+VNYjL+jvqQ
zOD+voxytVks8XPNS6jyAqgA5al+Dwe7RY9J5qQ0P/DZOpZZUAya/i7wm2UCiIgG5u5gNGNEUNdS
U3AyJ6NKBEyMpF0cD2Xy6640yocMVXpGhkQMjX+N2bM9KsLt1HFJc2rryKb5HZmasXjXGCxPFEYE
lgohxxlW+dMYSNtW57m1O0J7R40+Fa4hp5kyfO/ywK/PXjRyfwN3sPea+hOruyyHDPhky6ZuLJZF
q67pQUDWxnLRzCwCnawLpwe3hHZwewTDjsUPR89aNbp2PSwKamGcSovXwUQurB7uW53o/CBQZ5GN
BkwbzYUzzc29NusQq/7vP2y25r+flkXj0wM5BNo/DDnhPHQ2baOQl1Es1nHKkLoRN4WVzDF0E+o0
78b4e75vACoCb3uAGnPGBsdsNtBZLfuthRVC4lIQ/0bynwTJMipuHJjc5U8YTx8EwyXXokh8nfbm
yyZdSXJKa1QaTKl/FT384/r+K2pTSLDbHOC7Ai9pvyaF0uEbaTFNoYtgEOo1fu3y/DpNaPKSnckZ
cjXVXxj32MqsCoa+FLvU36XAMFqUJwCjvL7jFyZxNjbJvcp0FYAe3Wr1aTZer+ZkKbe4efAPOffX
q+sEyihMr2vnwECj2ZWvF7xRh8wgLeVrSGzn5SxZ2NHoodauXWP8MC0nqSPcNbN1tk/60ZOyRtvB
EQp6hAv49xBq9YCHlwJONST3iPSS786YNAQ8kcO7aHttDm9vG5lc24Z7OVB8Qqo/OOuX34sqV5Mg
SnsLhPjBgP116BqKnlkvCi0QSIdXiXZRZc/I0oZ/6WzlVOPCDPjnDKbv5aaDe8UwpvXc6xZzDbbI
cngYIMoB5Y4/A88uNujUAw0bGDrdN1Fc24WogElPS22Z7CivGLdgZOJOl/bmfmGY4LQUowRcVuAM
gke/Z7RljkA4raSXf73rQ7TBQBaHtAJWmOy2LIHF6b/LJxUGYohglSyq58EP0mhxSKX0Askid39v
bjHpxsViqNmcu765Xv9whh57+mtYYoNOg29//GKaP21IQ9W9RXlpUdCUlivhzw0hSeTTGnAAno2F
kjCLYG80FEK05CgaVUfR+O82F7LLcctK/QTSWh04c6R7Y5xcLcpne4x8BptliMsG0wKs3ZpsVLpv
7R2jYoblc3kbeXwZIss7IZOqQkvo4FcVsRiXrmHJNSR5hwQkErU3u6I/9RYfCguRy9wBBM8k6HP9
gWIXeKWGDOY9iIXrhN89mStqbPSnoCNelEUX+XTVg6hP+OxLHObLXLVTIz31berk2IS3SEizCOj4
eK3YRJJ8q9m8caVCjTMGhIpDWFdX9qm5TG/F8d8sC0P5/yeXNcvYt1OV7rM+ajgER9aPdpqGDIPk
Mu1CpVeq9VFGIw2p5A6EtchVAHqWbDdwQEyUXHLXjeWTt1WXjVKcqF19055+wDFM8WkUwQOWBDJz
9fdnaPEiQGXKyvJqXBCri8ev28j9g4++sIDmxyM9o6+YpADX50bnNT/xAyVgTYdQboN34pJ/wcZQ
jgYS9KSrCJNYimJbFGIJL/0ia01uS8Eddr4kI0UMdGAEIRHf1l/m9plHmcIylH6iXUZn/2vtzuzP
GH/35lKl8yO6wfBpvHJZMGhiEcHiJ2JE9yYohg6lKzBWTD/2WhfbDZf4VrGk2Kn4Cc2atr49MGTT
h1Wwynyizygxm2Ukzx9TG07v8oG8BnkK1mZ92Iz+h5tVkFL7HQa5Zt/6LA2ak2bm/N3w2tO3l1CF
u0YMidyp40aethAvQZjYa88HUjB7dVz2XRs4Moxe9oI+QbqyFYsQ8DQH3mJ8794IRfxAPEBczU+d
3BdhW+up5TDINYsS9zY+NqBi4mdcLoHMrtLxIl5+09Styn2SFj4xq+RwRDnLkSB+GvdoMiCOn7SL
vzc36GitsX8jsptz3qkB7BzPadhk/2zX2QBzKzcKGyXKEJCy8B1u382VlA0TZDGUa5FF86l8fPRF
FCDvmVaEOepT1ZjIuDLM/QPgq5ugQGyhXntLbENKYBT3sIktlcDO5q3fHeYrXJ1umc5L8tgb9DDp
Po3z29YBeeuUWtRann6/CDsE10IvuiW7mFTLMfU5fm42CXekSC3cVecRO2aS9q7dWhAVMpwQDOZg
bzFk8VRHVK/7qo58pd4S1Q8BlRJ1R3oHo6dKXzUy2tNLZ4xoU/wBIJfs70hmcMFEyp1/D6oA+fYb
6MFNLhlLT0zqe8GNamq9gj7bA89Nu6LLi4YKoCSMqKsqRD00FN4v+eQ8ka80KuPpQdSv283tTRau
oVM4xOTObnINKI9mctQKQ30oHrLxwA3k5UNFw1soi+sl77u0r9++n80nxkmD36fGzDIUKN26tSEG
fRSe9xgO3ixvtbswbI+LJIqrFiHziTKi6ubDPwW51eiZxZkff1y3OglbOM5Y5eHdkYtMoeQ8YiSu
afUrfSl1C28D9LhWd3QWnGrHZMWOaQ9u9CMpQ/GnwthxO5bTHU1X5Ayj68JdCNHFjzY6fiUZlaKc
V3mxvQ/bCMaNUUOUgPoEW3lTgX1s5MgC1nHDxZrhv8To6kYzWGS7l6Uo/FEtRtJ12wSE3i/qQjKt
kJHPpAbbwABHg3FSDBgvCjTgwLE3qDjKUDFDUuKRLqMwXe2u3qnkcyvPV4ZzLFb2a51XOup1J14l
PCgfUppSbA5RhOU/x/Xk+PsA3CWeYcSz7igalO9k+5IY8GZRPizwmoJOWecpSE61VHzAULCKyoZy
AVaRbt+d7eGajiAq8ZnxF4h2ydBhBKXdLioAavB//RH9whLGkKiaFKCLSeBuphIA4QDkafFPnP5z
m9/RP4/fJVv5aL6YgV4DPfYz2m3sFQpv8MSl/9+VPtCy0BjKys6mqgyDn6aAmH0MYDkb+6yyxeOJ
ztN7PF9Z0ePwZK7yLh01cGvokd88jWMVOm2az7ymDFgRG9laEEXTGxrCEBllDzEndcK/lsRrTYLf
FgHEjrcCZVfchZwGIVUXOPOOq2UsKGqywywDo+sIPw1Xd4VyBM3oYk/BcXcjT7GR7BThJqCVEY9J
moqDxDt9vQ9qOwF+WtOOxO79hmxNssnsMbxwdtZqLDepau3eM9MZHiQsM6tFLtC++xKHcxrkPC6L
SIsOWeGQBo/VdtPra2nYEhhyUls+uk/jImS9AiCSzoWf8qhlXUHRSwtj+njGOlItFEDp60qDWmhc
pnW0ukn2QSKV1+USn1j3RjaMn6YwLg2kQhbSXsMMTGeTALAAdcCBsghl5ol8NviJnUgi2EC0vRQI
BBPneY7XsW8Oe9v48gBWw12zBIt+7aoVIm80j5m4wqJoFZ0XRb8PZoEWEnLxtRMaQuR23zRE2Wj8
vRth3YOQtsCasHV0lTC1CB8iWXoFmakcz2w9n503SlNpSc9Ym3Rh+4qzaXoQgA/JlZM74POVbhvv
LWn1c5+unWF3/Ck5NHX6amOv2qrT6jrxKLxidvzJ3+wqrBwxYuyZ8XP68Yn6y6YoEWXy108GfEVE
/BlSTJEuZNvztjfcORMJWABIE+GP/puoqe+PZ519aksYHCmz8CPMr8VTDZ/FIAZ3JjcjjMcSBaJO
8GnlrfHzkZIeKOKfUuuLV1o6EEOD0JDS0Cze46okTOB5aGhIggejzP6dzBNETz9gVNd9pyiVT9qO
t+zTGKAUMTeyc9ux/kG7AmmZRzrNuY98Dh5o0GqiyPWnlaNpY8iF60S6fXMs5e2bq+eJVx6IVjEq
ETWnFN5NsV5HZl1pZ64Y5MhOf6GybnWWNIvMugFweMlQeZVzckZAPeInjH6pLuwqtiunjf8tbQq9
X1+GR3ybMFB3sEeRi6qBpYjfiaNbuElC/NFmznvZm6Sz3bVQi8WgJQRZcufxWKwssVlFRpwOyhvb
DM+I6K409XDdCqFYLtHlEjy3lw3matHEK+2VmKkd8HtEcEf0/8Wg0vvi9Fr1ZwZt2zJRbcz8z/QE
3P/gz2wZKz7YSkiRFheDtc1zIZtD0uXK7Uae/GiXpcDbEcibJMDCSMZEPT3yjC6ldUfpwvKrkpd2
/uw+kMSpPiCz/7UZQFb2UGzCAqn1VYAspqFMgtM+Dq3glHsfspKzb2GmehaWNmS5jaSCStZI31Lr
Jah/j5VYxM+0eT78aNjBTPlVsclzpoRLttKWVbkLpaJsFamNqD5N05abHyMBFiNvE3F1lhO03nDX
xvZZ3e0e2XfNKnkb4kQQI9uJHffq+cjYc47ePmt9F+moRGS5iQ4IA6m4HEQ6fewp97B5heqa1sFf
oKqvdDQ+tUgs03FcICOawDSPjum5Y9fXFAhB0D32IlHrV6UhEXwif1BK6gp8DA0I/6xZSvnandUZ
4CDZTZKTNX57C7I9eDuqEQm44kwPhn8yl4bVeozNoE3XUlKRtfU7Fm6pvySW5TMWfyjLQBBDfqyp
O/ubuoWZ4bLNPQn2BU0weB6iLdMxl9m7Rj108hfW5LIJk6CeFXX+sGxWdJKTBHx5jZTUzEykJJ/A
O+uYeeZlmBe+pslyMGzm0Fyuvhjz+1ySNuOVoLZQ7AjDPzS1hTHesgNR9llgZxOHPv9+/kyTXWyW
PwySjjk7A2jBigw9tGYMfdJ0C80gDeCE+KMi7FudIoZyFgbl8azTqW8se5UmLSmVMeo1E9AOuPul
ALpqLA1TXkNTG57U5vNrJh69Zu8lrv5AlDwml4ulgIWUwkZcD1+5CpztMZAMzZ7/1czHJulLdAVf
IhLM5gOlUeUj5NBQ6JKEz10iR8CiRekeq0s68zbnPmwjmLHONSMwkhaXdJvjCDIKwbkbQ1TVSKhr
gDnbVad4EXNRneiSpKNkY0I+38D7Taz7ToGA6v1casZijx14n4z1dq2n9q6jyVZr+/BsHADr8HrU
fgg6XLd1OmhDAgFmLUEJwCkXGO74T5dNlYZr+qKCs4V9CkNKrV5g8B0AKC90oj9jvYQp/B40EwyI
navcNixjpkg2z7Cr+bAZpFzC6LtD7cUYq0NMyPpm3D7D9TXF+mvnCwOzhLQCxutkRDRs4hnEEe/2
bmBEfa+1mq8u1ZdzqnJoW3dF3P33TrYURHxlpgnEY0uC/N29hD491/k65g9xAV88NwwPS3TceVx1
HmDgHqjdXy5jcq/7wNePA64NQELoCTBxeZAn5hXB4R5IdhEOLg+XTnymJ9LN05PyV3WPj3VRSebS
t5grdzZVCnSU3ZdF8rPuE1oLVwQs9W8IVbnhJANRv0LXRXA4uFA=
`protect end_protected
