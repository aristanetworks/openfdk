--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
DtQ3Fw4d2cyZF2Ht69OAYANavWqxV/HMZG+CfzHL5TLxkeOnUoZiX6Kwmefe1qnGfteorc4POdVo
RkMaIx7b5dGfBpkAsosAk9HpwM+RkCjqgCQWF1szXRZ2tC/Ynfq7Ox1eb7n08NktdRmBgRd71ZME
csOOFoB8EDxVmQpOnq8xxjpTPI2duZJyBeo+LAtysEeuR04S++tgiSc+6JRuclG0K0lMTYE2R5i8
fa4OXnUQH1GLjv0DC1SNlyHCdM+CKTTxN58OyBh6gCowNrTeHB4WhoPkSf0UMqP328BhoIG0Gf1s
6FAZO6M8zwNQZgu/sEE9CjSr77Q9IhINuUdIEw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="0GHjiHMH+qtkGv/jPJOp06lY27y2sYNVP0OjcYo+Ecc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
WT4QA5eClZHmnzCGKfZJzxqbQuWaYFitCB63BNTwiPOLst2noAlQ4jiIvMBVjuRFy0U9sZnki/Wr
YLM1Lybn8Q3HV9s81Z/qzfYihJSvo7jmL1APXQauTKDrjysP9maNoWEEfHsc5UZQ6TANOgfIHQFZ
ud6IK31tAihF3tEnyQRejEjTyWB5ASuxB4+3EjI1TfyisJahyrOLAJACMHqL1BxA2yUUpW3LGRy+
dZftHSinicopEoGyCzkRFEo5QLJr6PXRQQYq6Ud60bIxEILTVG+urBRvJDTGgQyAbmu3wGXJGSv3
2kgrVXuGtILw40SIBi+pKUahRjshfz2mUzbHnQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="zn15FO+p9mwEFZMvkJumpyyW62Gcu2n6OvuzSwBaR3w="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6624)
`protect data_block
VL5pUItz4rg2mnIt+z+HtvzD+056rZqCmWXQOuklovhkkEKV4uNcBzCR6Q9nhCl3KJU7e36oLIXT
xMc2gj32Vi7rJCdtNVNY7ocpAbSVefy8nSO8duBWNCygbylOw3o+d+BWOCiFl7PpXIixXu9vTn1q
J+sWuwaZ15Ky51Ty6jINKxdeZPcVzhpsRJQ38xszFo/utKurk+ioKpcpyV+kw6rQUUHMg5JM84PD
h9jb63qoPg58DRKNv2/2agaDotZuKvaU28nqq2Lrt4U2LlCfxhm/RiUTO6M20bst6QBsM+RO5fiN
4dJU7FArqM0xFI7061r1WY39NXQ9C78m4ZRLlZLFKJFVuUZH2H8pzlJ97wmu6R3H45DeLN9rM9ci
4Z73rQVBzeX21FzNjtfr0IF1US35R1vyjPVkq/ycs0zFJrjlE/8YAoKCka3+muZU6ihSV8s/0f3n
FctLO72F0gsoqD0pUIFWdvyGvGyfLGzaD53AkJlRb4ORAuoHSpvdBHBJNQuvjZ5DZ243ff8LGFxh
WyD36xXCOESuIE8+PJawbXEIkcWH5pT7ez+XzgSgft0mVbmYnCkzNloEgUMOod5oRnmaDIc9YJLr
AnfPZi/cXORbh0irOBDfNS+0rcEM4QkMY7Cnqzw9ODu1xblwLvauKssTZ8uyy8HAxQJ5ww6iB2x6
WztJi3BLnAbYm0FrS/XajBw4ZnpudLsIsFstC40E4VRrmubjcLdok8sPGT2YTf8wc5kVZ40pEHJx
Q3idJYaI9x2VMPei7150tUqfUEAc91jQvyZcUu7rEBWtOAYQg7EFXC8ozWkdpFAetutbSKs9y+fq
HD4X6K8HQRHC6UNaNEvUta0zZMOKHV70D2pfQDte43Se6fheACc20CD/JWBEqmetkTiTcIH95vJp
l9yH5zqaziAIx9B+HZSjHhuNOxrrNRzZJ8xsEZHQYPDd1rGRti9HqyOhASyTTFf0getB/4sHL9xJ
dV1+K8pBPQM9sOJvlwGCD62S0I14MnwsQult+auV9MLd9qVCR4weuaV/U1fq+HlurQtN/ODEfUD/
j5eUQuqdzHn1yg2DNxvEaTjcixWkAx6nvZ+32c1CahMWkOKgp1Z9VcMuXuekW3Yf5owwXt+Wt7E3
a/b+CbB2rz7TvgMZSPEBQ+nQrkOyCgEDQFq3oBT87ZDUG5tqhROLMbmTN/dlH02XsoVhu9/uZnA7
gwLyfDyI+ycYsQPmK25GQbhO0XkyhnS3BRFfzG3h8SKr02VSKGIiXpD/fGhpHTg7ldGuDfugwQ1H
69Rq+d6m3G2ydrwSqY7j8zmMNcRzQPE9yFm9v3ycPvmIsUrbIdSM43eRz2PjJXGobUYGwtCa2jB3
OX32DleOIxR+7kC3Y1Z/857jZ4K47Xg61y7XvI36bsSq7AG9v1BEi6X/i8F+rDdt5eI+vEl+gYJi
E3+UtrU+28xOXy1QpXFTXgGRZnA/YA/BEofUQhPED65HHltBLldf3F6cMZg8f7Gv4BIixY62hjMk
NMZTaej8nrkU37o0KK2sS+/UQ7ckCBEf284P8Zwi+O9kaWchljtHVlOSnF93A/lbmUvA/RI7fCic
vgYYp/bYCs5B+CtbeYs+otMDL635JAkFOHrlzFVrbBhEzxcNJGpNfCcd+lI6NILh5+UzB95jo0bM
vsDxIpgwi0BZpH2BZiw0s3CQWTLAv9ndJV+tNfE0ZduA9bEZR+oEvnS4bDLp8UJFobDrzhW3nlea
nBFt3uDqKM7/bh8QgpQ84zsnWabpOoBFgfAmYw6vmfifBOz7QcL3JPV9NJHCJYsFVEc0Go5M+PRn
YEQNcT47jiIJfFTvOhUX26mS665h0zvSnJqe2LcV8R0fldQGXmpdPGP2kpTCw96I56wf1dc1eIPz
70OPyFjMz66NgcAa6x7Qo58poWlLXhWGsF71EJRpUcYuAN1FMN5TTseomTWA8p/88rK2DlzQZXus
uLZU6+b2akTTpIIc5K01uQuuUmn9sieKkSDGmcPT58m3T/8FX8a9fZQIlpTCJHSfPIjz3xG1TOlU
GHLQVugWWhcGY5TNdBIp/y5aE69m1dDJgaXJYXCf2F/THrhOu23DaOZWM0DetR0e4OTlG4lmuDvJ
gwJf+k4egmIeEwm55Igj0xCYBbsEzZ4k2ZE672+IG9bErDNPG05nEFM/Y6yqtpVxNSVCsfI8RUya
8j+UZhpqGjQjxFvyc6RwEqJzVU0lsbpjFr/r+S08N8N3ZgzlzbJhLeeQV12GrFrdSisswwSxk2m5
eEJzEVW0tty10zT9h1Cg7uUgCgQXALTSZtzis6BafM4CfuNo2we18xFKA0wEx7FuwWcfVM3I+sui
yWC8UCVBJUERjnyAV6RGz2njTOgqVxsSMAGCvVY16xe7MD2ej1DfvOuQg6CDt9xPmyk2BEN4QAHI
jNqQmY+iw4mZhVLHcZW/8hCE+A/0UZ8Mq1t++87Payq2xgegXaDpWdUIiYua0LVONI0p7mkRuUu1
GCtCWbdrEL6/6l/VUnTwSqp/pUDTV4CRtQNIChQ2w4SdFIUEc3REZNF1j5Lh69Ouwc/8Y2lRKIVG
eaKoab8epfedZnkzQ7sArD68q/oW71H0BCflBBQV5EZ1C2M7CtbSVkWo9kNDtVRTGysu5rOerPYX
5wQK6R4hjoJ0fowGYyEJ9ErhcHEouGIYwLuC8XebBNyBRNl7zyqOtiMP7nFa0KyfLBAV/OhNWeTv
uiGnFry/Q15iEluDoLcHrXO1Rf7w1lSCC0eQSoLl9U1qcV6Lx8xv+FknlwwxcQzqiE0ruw5ijCcU
Ntwv0uMWNwyD7i4YpNVyJApCLlC0ri3nKH4w0tpey/EyiMV4V1RghwE+qkMH5lmCGxTysWil9H9+
fPM+kgiU7Fi76/flEThu4OYVu6rTnTQ2J7AlcrfZvCQdHDBOp9mZ4OOOUgCSRyzUNWolO1bVfVgQ
epekNXa5DlF7UrCzJCjYrM6RbHsF7YqzPogqV43n0NGAINQEOICrUs4k114lRFwKS2CF9tRKFFm7
21TXQZPNvaYxcmXcF5PvoApQgmzOiEy/KmqQmCh1mQUS0s8eJos3akDY2EebvQBYPvGxG+McV8ld
rIO4+6whBzpzq3pthnNbFQoXWpML15L2EWVPTKB9974ZNmiZ55MWdYGEWaBIzZCG6WoMkVn9OcuY
nABlYnxHxIilFZ5Nkva4oUqttm/o8/lrF4byX08nnJWnqTjKS/TvNp1eV7fQqIO8d/N9sTFxnlSk
yAGVVQZPEs4oKUm094htX7o1SWWjxLfaP4InNLwYSR8LMf/aT4czlP355tNwRGbRQ6b6K4KNBGiU
s/OxGSZ2qSeZVWk81CaJNHqDqCX7j1hzHOaRtMruaQALYgdBRP4jNYOj64PwYditj5/3QQrtelZG
go+jNIopRsCw0qmXmybsNDLdL2u0Ip4k0ye7mkK6+e4bix9j1hJLOK11V46aQ3DdUHYSpX8HKDX7
2yIT/iMAYSuQPQYSkwWG2QnfjkjwLBEJHZEU9YD06VqETIDDZLqWmO38JZS49gBG2WrGWlsYOySk
AWnNKNe8b4In60EG1Fu7trF5r3+KvyKSqNmJvVRbzBIMnxUNPggZyiTesvRsguIqXOVboQOvzPiV
IdjRPUS22NWl5jwTyKQgt1TUclmdki2zjii5OdFYeq1sgwemi2Dd/VvnPRy2tDNagXgV0w28fMYv
Iwz8bY6Mw78P3N6M650j2DYE7bXcseNIRGUWfTxEQzptX+pHevuhCb5MOt0UJphM2i//E0DRaixt
IG+2jQob8cWnMyUtMHAOE6Ru7E1IRaZgGJlTzE7ZAuXQGYU6fHXUVtvCQFmc06pFRzs69WqQqyWU
qyF7CNG0M3ceoNKZpBdQmNHuRC21STP15s2ZMled/C4/H5/3k+7/DzEwirOAaoEtcZQ705fWh7n4
H56dbSnPCaJWI2TlwfNFirkmnVCDgsKdAmiAVNvT2QBKBu1fzHxcBz3Dp0dbqEUCHtwIA+UQOd2d
JtI1NIzApW70fLvlbnC6oDwNlXkam2OqfgBwDyBYu+bVsALIB+QR88bQFAQ7Zyk2rScLaxVO8vcl
uFVs85Roib3YrErQSnCwr55COH4wPACjZOTlBkDf/BqudS2lVrCPv5zIX8FJNskgmfscp88SW943
AFaUSqyg+rY8GXAxyZUFwvZKNNvJjojGd3HAzQK0F4pJVq+fgRFuzT9+69AJ1N+L4LO31MeNLQze
EQLtKsNzgcGXXV+zvfAj62eGhZlvK+S8/kZsyid69bI2hFE6vkuTR7YQWse6QREdCq7yefl+OlbL
3uo/R1GcnynYG98KwCv4Ln07SrIXDv5Y1pXSFFl+t+4NT+UYqgjSmLI9e4LQ/x3h4GKT53gjb3zc
JUnxyujKLvqXOpBk4NDEduGsiRQxD4Zmt0587AMZjnOF6+DKcWiGKWEnyj5MFGNim9oz/szjRZNT
ruP1EH+qT2xbT/sjAf4EibOZuki4xyrblWRKAgrCnt1Eeob9Q13jbiAstm5BMYfry5RwSw5e7dFt
OFkLyRAHLv8/hmiMFTsqhYxMkoD6iUoacvG6Ivlwi2u1s1mP4ksiGyoMPnd2WRAWXHn0aB6rS3qw
K532uZk2iJIfq+vQ/Lu6MEvJQfCMQQUjODEeNtI4nQFPaUWBCimEoasd1IozKCp+YSoTmKZkozEP
W1qhX+c3JOFiJ4jt+/AwWZ0te79QwmWuueB67hn6TtCvwQ8c9U4MMoRnoUcxrZMN7sEIc7vz0Bj2
wzkyeI9N7eT8LO9Is0AafsQIGIEsUKQxwRN5vs75g93jN7HBgc2rJ1jI1k5GcPGirQkDwnuHYl3G
KZcWXBSyKMG/V6DcVGJSvYFPULv1LwWSjjK1LwpVcJJu79q49PMqXG3Q2CHOogcsVJ2L+r6qPHNl
nWmHmGJFGtp3tb7RwItRgrJquHqrFfgsvAQCI//OClIVJ86GCcnA25HC1c5uPZTqDfrvmvtFddlL
TfBLv2877DxeQjeN4alhzqJF972v2sBzD3nNLzrNOG8Qaom9FgNjiGhQNVzeeM1k5D/yOlbd1Wva
DHHi3byl6yde6AAQfjznoUsjKiuYwodl1ATM6ScF5KLqWYi3CM0/fbKlknd5DFpZj+OVJfFVYGKW
15rFFx8FXMZ2LOEFLQz/mOkE3+Aqz0ndzkc7ubjAqbU8SJwQ+G9hicWQEBZJUnFY+I/bfzq7RUys
43BhRVHE/gt+sIqJP9c8jyI62kN6uLA/WMNvqRgNXyTqvWTH5rjX3r5jCn4tkAKyeahkieo6nYWq
blvV7VOXmcfW/s16+Q/exvKt0mOsvrCFIMpacekU07SMSV95G/JBaZNK7ownCleR6L58H88rSrNx
jl3VB7Ol9EQLHJ3yymqw3nYEuXqU81k5m04o163qZoyi+eI7VxBy2pv58tNy6dtafG3CGi2rAURY
0bw53eXtmXM81kjn5rWEojxRVRH7o26ETaxq3I+lXwW6+mUSAxppgVhxyiF//79iN/Na7+NoazQG
hTZjGtbU5A/YEZwOjTL2+ues5CUQD2MVxCk+qsKY+X08DDh5fBUDp2wxxcXZbBNMNNciNPE1/jo5
2T+DmKEyeNaYWYzuzq0tAFHsuoqwawUHVeYcnJKyVb3dIMDIiCYzdS5siuQfxvVSgBp1N1Z0OgvL
EcVirTgIvv9jttuGXsPhN8icMjsBxzfov/LuTRZaMyhUK9WioCCdl13aA5iuZDX5DtEoIfRDUC0y
VlGVVbbC5LGP7jUKpd/SK2SQxIp/p5O7LPWEzfCRfD8B8fWqFxL/m2hdg4SCJtb/hgpo9mGFwebd
XWheCEsywYdGJrVbnHEacWR212Alhx5mIxDy3Fuof2x3D1gDxuM/IcKLJLJmX1/q+5I7URvxWmq9
dkMp/g4VD3mybLBoEXmeawm6GJD9cxnuzccxKWM7bQ5OeJihIUJP7TNWwcBOANw5eM+wLvCCBs1s
Oo/lkpoXGL+9xv5bRjGFWNXPAKJmVtJGCYbd6LY93e9xfj2CYuac7/CSsZzYEvYb8v0u55GUq1k1
gswkUSstIQDm5TMlfRqKMQJJhS324NFGho0kNsgZjE/5Dgsd8GwpD3tR57p7VpZXIFWaWvtjhy+a
JnNyXGcsPjTc3ANRTMkYzpc4AP8OQD5mh5rtoXnXkKAwOMNIka31K74e5XWY9JDlMpa4kwJPPZUC
EPezT+Kmkt8MYbKSaSX2PAvoUlhzloexZl5WZ+LG6heEXkPQG6Y72WXubuxM9rPQ3Ew4yIrcfNI8
RTn8MVqKe7kwlMvU8omEaRzdjTxbPGqOj5hwOPU4tOwcqwATAz9TySN+gtDth7Al3PaDHsE8gDUC
COStxGigIzpYVaZrA4YXUQgaf9HHmAd0rvPWp0zO0wVVROsG4ALREF1wo4QV+3ZocrNXERn+XbYX
kewg6ngnibBVd9Tcr7BMQsVC7EukkOV1dFBH8QK7KBER9dkuWRZHdwpnMUOzPzD8RseRLIVPEyex
m5iWC11lrUpCU5GimzPPvX3lHcrylEYSWjPtZzS6pLR7hIqZgzOCpOK7mE3tVccKSEng5w/LGChi
6a+PvmUJmMB2c4mAoQ1eRWPtnzzFvHtUEc6gpiN28t9tClqWUAthxXU9eSqAViD2bF3zlLbULX9w
VjMQdcMXg7ZuOT1o2sBfXNeElUYfotzejPtivueGJsIlvjOVVNiRfOWqfr3DY4uSif6SSdy1IHW9
9nkzZgsbAiVQwoez//78mcw0Y3zUo6C7hzPCD8JT/99ukbQ9HhT7rRGhx+/ytpbT7ta+c5+c4PKn
G+feJWzD288PZLP9J41mUuTekg7WFHbcNKhOELr/3yyy/heyPZsXF2bUBd54830vICmvnUF7WnCX
zh2S39d5sOakIw5V3C07nwmVaYH4aUpY5vTee6O6lKxyzub0ptb5PZYSZFJQSQKuQmCIJoxEqhxB
lPeR24GS0ZQhMRaA13Bz08jZfABNe2yt+FzEV+5dy+QIVVROkVAJSsw5SSdiYO+egREUeasebolX
KRXfA16UQCYZGrcV8+UqYbUosN/V7Khyg6xtxCMbw9rB+tuazDRkwG4cMRsGuA2Tg1nD9AgaWp0A
GYmuUMa8yGZwI9i5KAY+MPikHCp1Zes8fo59urLRP4J4JgkZ48Jj8ghrRr5aWuLkKhjjLrHuvgK4
/JtuMmPq5DiedBquTnSwBANg3g5S5zqTs/8kDJyjy7aHYeI0DsWJZDtIGdK0ZfvlLimVaES0Zl8u
palPG+MggrgXOr3HbAMLzozMHS9ywV/N4Vih2/KKESYyctd4zw8AEMz9JkjPS9L3rGU9EpDHaoz9
K9r22ZCZ3nxzidhGQaE45o1xI2uPMmXuBvUOLC221gloXcXX5R5Vg2Kmo2mGZ8xhGg9ZVVLEpnWS
Ae2/zxg2GU9BeQyC1CvVwyGPJgYpbRdPZNrENmG+4DOFtj1OBuMTHMbjgCZrCkrR1Q//SK4w8d99
TShcIU+8hEff7LyExQVkjgIDfe7vQArzKvRHHZlcM0Fu4coXwgeo9mVV6KzdUR9NWITHT06wzYJh
jCS5+8VL4Z8CKj6rRvwb5aE6AIAq3paWr6kPwvKnZ7oMIFkV5m2ZfHwxa2rFldbn9Ux3h6sXMLzN
Sik2BuzGE2+mC8UnkXnbDpH+C+v8ptL+L56PsXUeUbDV4kAC5bpCfe8tKWXHFwH+yp3Rgimq/GCa
AM32HcoZC7GtXoRH1uQI/MovoxN5AAwZeQd1eDDHF20L60Pw/3xaVdVAJMIavKKsv/fQWqiyvkkP
jRdjQIEudqn3c1Tjw1DQTo2f/rRIc81fJimoFzjv41cx6DFiDAalDwGZhmCbDqI0X8lbfjLd6GT/
quDSkOMkznHGJI+U3S+3+R0q9ooP3W+12btp/qOfqOrpFu9u4hEBMAb+dKgKBuwVdPWYRBX1bsw1
4f0ObU2C0I81HhAIwSU1fSjm+yTEgYnjpatWlighmFMyRX/pm1Q7BU4A12CAI3PcTCDKUeV+3aH4
DF8OnCN8IoMtdIMFqLQtCZZq/y0stZVgKS29oPAK1jf7meyTcVNSqmACJIQENL6m6rbe1JHDtQDY
aLMKCnypSqjygoZxgIY4m9WheoJftP9pqXAAOEg8YkJh5zK22D7XWdnbr+5YZqYyg7BWhVZexTuA
CzQlyT68ycgcWafHILk4zN2sXdUag1Z38TkDsw0clPGKgPpPF90DbSLJPPPz8eLuj6JaJWFbMJno
72O79GKDvTalBMa02EAB4gBLpmHVu1PiNWYlqJe4lxzIoOKoW2RwGL3Zh3B8OzwmkwG8TGDYS4WE
othe6DtDbcXYoho5GmPTMyy/ib4ekEZiM4fiYBd1bokFtVLCwARKGLpMj1OJubM/+iYse/ocqZl6
TZVsllXkoSncP4Aw9HsZB1WDscO4szyrfeO9r5ITb9nu7Xg+VDxEmweZehhnJJIvTSAEGTxizV4I
2NwMdyxG6G2oHnO4UckDVmpPDIGgodaqRHsBii9dsBACW/dWYof3+spfd0jFHwxOFqsKaZpF/rF9
QYwjh5I8jglVAXMDZ5etbFB3k+4bPsZU8nijvfmIKRdSCncpjsYUK3DFZhC6yrTDpcDLrp/R1P4H
mHLp55fBuex6JIQMi+FSrPMzHuW8cC+9PFSlsDWgzV6NCGoVQkZIZlqPtEhTwPyPkXcIhMoEzrYb
QB3GS79lKKOo30B+UwKKtEawLGudmt2RMTnr/FjXPWLFmwO91XY22mmSiMqWt9f1zltTAJuBEZBZ
8B0EP0fTmGFb1SsD
`protect end_protected
