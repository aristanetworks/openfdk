--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
k6Y/+Hs6xELNIMYReMMIW3dOeW+U4ihdRh26tGRfhZOB+McD29iwWSpqRMutJsETBLMgzrFCUY0x
e+2HYeZvb0dL07vLOUAd23NT3N2u59VwFsZv2oP1sHqkYALQMCwxx6IEDWZNm/H1taG6JQPFYKcH
TgJUaWOk+yCj03e7ZwZqfIQ+YiqICExDxTbUwtZJpKX78R6zjvwD0FHqSSIJf1OLwzvl4jv5Po0R
pq9S6A+Sl0ZEDtCaCh1PRVelKyEHhb4w1LHYNdgKlTFrPfKfXu9y6sRg1b778jlMEgdWgaPhca3o
kPXTnK3xDr6JRC3CvzONtzzJL6dFD6PuJ/8+ew==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="sI2a6B1Kbw7roA8vVcinO5mmNaA8MsaqGpNPg/Ks4j0="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
ZKQtc0IuqMPZmlzdqFDhdk6TV1HZybNoOFLo2UgX/5K+ClHzCduhRB8Mn/C0/5zc0+3NKMFTV7gX
in7gMTOSUk8sTWjED1Jw9Pebjp3uTSPnTuWwgJ4ecKJ7q4UCICJHOU+j1+qPW4bPQKp6yx59PKBs
b0eMzx1exUiGqSTGHgsnAh8jy+EsC0uWUhDbwzMH1xqmYTCGSSzupNWS9YAK/cqp4yTQfj22p3EL
sQ+UGOt/FhY45RPFvFpZPVqq3dF8GpQN8vExrugaWqqZ0dS9v9ktNIyiK00D//m5T6fH4f7olgTf
NinCzMeoGmdKkM3pNSDgNRvQ6X7J5iNFXZCfEg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="d9vrSTaAKCWf362hD4fU2gD6Mf5vlir4OY7THImZ3w4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2320)
`protect data_block
7YJ0xc0d5FE/Ioo9uIA8XtOdpbEyKoN90OA4wVjkkM/6fJlpYkcJbISSH63E6lWIGnDEPOEJ21IH
Cei/wU037Y1JTxqdo+4nqYJySFrd82sveidPFh798nhFUItPKJT09vXlYXeVqDVm3fkL/+2p7+hN
SpIV40N510Pf1YTaNki3ObmiathkEijbvX07FXByEPFCbopVf1YTOtAxH++ZJ6WTzwNQybpMBmej
+BaW/wqC641NsYWu5bTgmy72WNhHHWLr5IvxbwPwKEsjN8tWR6WqOSlC4yAAOMDEQw+1Io4vFQuG
Mhb5orebUNKDjyoTvmG3V85V24ik6fTqZyNU6bcB/BTuJyj7Hkc70VCqyQ3wptwdfmcOYve4GjXA
+LGpA0C1r/GQGH8Fmb9wTwcuXYp/3AyyeejjcH5PVulwWnZYLs+tHoIET1du6gqJ/3dIZ27lR0zO
gMSJ9wICXbhN4gwtVi5/NRQC5lbzc3GxzQHtSM59tRTitgxLR6vdC/bz8juYLvEyOW+ykVzyfctN
aeyOsTRCPOahNIPF23cxq8N4ljIEd49/w5ic2p2drGwHjjIZxvFmTFLiMr/5yW8Wbur1wsf79gNP
jgRrKgY1njhh++LWLQ00eXA55d1v4bBqZF2VeiOzxmKcyFD+KFP1yTHZ1NkWhJNBaWMgFbCVuaTb
zO0VV/T8cv6eu+J29Z6dsScwTMpOehs5APZsG+FhV5axyGoc/qLIt5f+eyi/9f31L1v+JW9vesZk
nLOlTK6X4LX4j1qulD1CpbXr9zDSfLz8N6S0nN+/vVMTvXui1TnvSf8LRcCwHvum/+OIU0XHzknY
Dk7oXevA+56A0yam8Skhp7P4WDEgyorIxcNAUFE25TmvBHBGfNF0p28EosNu8/pNpjQtTMuDW33O
bzyFW5n8vtLxHFdXmc3TKZhz2Fuul//jbdRkozp3ni0uEJW70qAEqkb+HJXlRc0dLF/VihYQoHtT
AWZGOvfoFIoFEYRAq4mhIi5do6W8/eHLyrWIXO+HoThT4jaUy0PU/H2voDfuUrTi53xhT8cACHAc
/ntUQKxjEHRIaoXE/rGVAaF8HsNj4cxqf40Xj7Rj/f/50HYGXiRb2Aqsgu0QXi4sd25kfLGzEkFi
frzvFgkRtlHQg6A7eEh86+/aCsaFn4fTHGaFJ9E0TdaxCUPHNfRVbx2deHO29zEMcxNw5XtcTu6W
dLaWkgKDg4rwFZEVwwR3hl1h/65O7NOVnlPUPTy6FYaAikVXie5ffx17ECZ3xZcNPuicmRKs6HyP
e/3ERWzFYVRvKFbLDUelwPUIeSpMEXmQWfJgqCYWqrRr3a49gCH2WnjrW2YcIBuxH2j0wXzLvMzX
G8Navvk000vEDijJ5bs29Kig0ey5SGrg2TTsiRqtCYuSIcCLNHrBNtms3ABslnyMNm2R4/MJQIef
TthVC6Or3bGOh2yooqifXd4P0DIVpS3XW3CejuaI2F1Hri54//4Rl+Bp2hTeGnaxrrD2YoxJL8eg
HKs/uurQXsDa7PEGVSIzc0W0zYgKzRjekZoo7pg5qkwwYO/Hbr9QYkxFtIio3V6nHQLhZwu7euvb
pApZsWF1BZrhy9QwstnFGwc1JvArQt1tOYarE6nrV9hciGPt+Hwt81eXWvOFJP3BvZY3smBUsNrJ
QMwa6fGU4q+LrP2s1Rh3iZwKyM4LBraKok2VtxeVOQOxi/47CyjFBZ+hOoqyvgDSrpcuACDLL6oY
n+M0TBWWqG1gosvdLHvbSttxrYYkhVemtHE7QAbT+/PIGF4qthceMnEQas43DjGDyNLLqE5rXVnn
eoSgclM3/NkaINqHLzRqYMHRaHKieNs1ocJdv++n4wMBMCt3Xixz+TbF0ULMfw/u+ET8Ov9AnJwm
W4v/Ld+OhqRGYm+4gpRY0SDnzN1+uXgnEwLlkPrRtmAaTLVKQpL08bm2FNUawG/hku8wLTL/D1D5
nJDCFWgeIdCR4h8VWZrx+P49BFHAFXIH5E9M7Ie0diyr40gpTzWHKAelqWtktBoP92SSw6LgePbl
v0uOXml/OAKtlM1Mp98SIe3dg3dnscbyDza67bajwl+nc3+sOcRnjZIZcwn0Tux883ZUOEjsSZpR
X0bxA5rOTLqtXRHSrrsdQU1CbZxUDvqrZK7Lb4JuKjZoda0Ce7WwElQDANKHWWq4SAm1efWShQkW
tvRBtdoetwl6XH931iOjZ7FAk9I0T+nfMpan8eeXDqrXMV1rI+lsTKCb2gH9l7s+bQ0D3XunHQZg
ERL6sDG5pJGEG/k5Bvzy/VztMsSPxQBowpNNdTjlQmXjRt6qgegilHyseROUmpk0QhmntpiXC5rw
w7FSvDRfMd5HNPnz9R8GoPuAQFJE7hN4GO8CPwIhrjp9qQPWFdzZmHWSyFS1A3PV2SzCOjJfJSSY
DrIfV55w+mc4XbAXAq1OlIvECu970ns30CmszDOqgZH20/vHHiJsaIPD/5K523AZq5sH/c3fjCKB
FMMHwNLVpBn9p0W9Q1ROxBhfHUWsWxUe4YmfckXUHujm/gO9CMIDPqs4pyOszAAm8jd7AktDDMSg
8IgUrFQDeOiJjQ/q8R8OKbemaBdgrbYRcrzF7KOttUc4/2mdDnJjZfLFw7Mxm5On1mW7sgTWLV9U
m6L9dbTAJOtVDy2js1QZIj17Pa03wbrFXt/4oMd+ROBK1r4kOwp84R3neqLKYktXA+TlxN2MDmRL
utXGo7smoUpcULErh1qg1um1DbnGJJF3ApOU7Aa2FB1TcG4ONCpQu3yx/pfBWa1tj55vPMHRYzZx
JsIoTjH032XHWqWWbX1hxixmCSMTVQPz+8aTbl1ePRM/uosQOPyyKcMvajXng1ws6e9/JAjHufdH
fqonfHXkRfsr5AWHWPf9BkrPXHAs0T294eWvdRfBIiGtlVyHum8i8dauHwtVvnTRNk3nCTcpneAR
oiqxWWb0viyP/jnynQlNSkFM6yXTKZoQqLpGGyc09Oz2iuB8p+duQnVC/YIw9p5uNKlAcOjE7URH
Tyx+d46oMqMFHpilL/K+F5bLRrEtimdnP0dUa0ydbaHr8tPjbM1gKw==
`protect end_protected
