--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
fv/ZbXnpJyrlO/tWNghmPaQpQgnblpNdHaiQ//NBNSgafbZSD6vZ8oYM8SpLH2LWJbiSW82yd9Vn
HjH/wXhQ+HCDRMz0xN9Rs9TtDQWhDG6gtXkdb1Rz+/Izn9PuVA9gLYaOLkgBsbs/MV9X+xXnaKbs
XFVE8vXJe35vX3P1o35jpd86TWB5haDvzjywL7SqHvwzRwq8YMP+63IB2YfGw+mDS+auaYFp8Bfb
lWtSGOFNKzHRIB3g+GuZv369DxxsR9ekE0gLiGZpnpxK/q38zQru40/FvN2LK9Dv+0USyf8fLVqY
2uJBOrFi2XY+twGIHlY5xzvVqLWXdp6rOwclIQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="GHWj+EYe6wPPF3/DwEY/vIRroFe6Xm6g05+ydAeftR8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
KItdSFHncLpYilro+pg7t/GKlOKkDGC0w/SViWR/yAVfXHztgASShp6mAffr4t9pJJmcjC1xRB8F
iEhUOmXrcKE5Egroab6MAUsWaY2IHunyZMeFvvsLxxH1fZnKuav3450PS8unnNe2anR/DKyQVRjz
cOgJ1aOa0SS/VvFMpAYKYn+BtAdqCrppqbZekqztkMQhHa94t5nBG5bp1IqdvB3H312BRWFa1rgs
fb3rt+w1sMMSh+wB+gprV1DPzYny34hXGcYiidyH8yuZWqYfcjhB8sxrxKlyKb7855jQRj9NAFS4
LRulS8vrh/EbN3n5V/lCJ4HaItixIG737mH7bA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Ql6SYorpyqXJIXkWngWh2GPtSOuEo0sfIAUbRWZmBHw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2896)
`protect data_block
WPzbn9WWLRAIwu5aQdrhD8UlKVYRbh6vQeyKrNNx6UFc9HW5opOUsZYPpmTAGouYRRWISmXR3kN4
jtdLD7mrL61nL8LGsIkBoo+98sh3JiOuH39psnz2X8hFFKhnVynVr+c9gWDOv3lHpSZj3HTGA7Ot
k3X6zYyYBnN2ltqtKmOg5KPQTjRtoeHkHj9z60K9zCb8UXJ5mX3hHuLIR66DvhwEAEZVd3Lf9uL/
mZCcXhyHwdqU4bSa9sypNeMGXrrEnDf3Yz6YEWH3rfDb7F01nrzpr6nsxUOp7u7Q4BHYy4XFyBIV
jiGMP0VbDqwpIwCu4NT6dXhebuDThI8iH2q+p6fjdgWMa7x30F9gNrq8nLB612UuXXgYsojBt72p
gheEyDcnFODuZ/+y4A71Fy4l/zjBosPp+HI/4xU6xbB2LXceNwsgufzlWoCVYC7SySpgxkmTeRxx
xgi7MygGirSegx1iInOhKg33vyI539a1j66K1Mwc9wQ0/NBaK/lW/IVo+vy6AKxYQkCdRopgUizn
GePMMTOAGOuE0mzuFU2+vnqwSH2mgAISvjNMPGZQvMSdlAexQ0DbVzvsOTeTFLHrPF26L54sqPRR
btavyaceDjULOBi1LHzRBSzFPhn0jh8A/+ifeQdykh6daJX8VD5JGZh/tR74JlW9xuly4G6LgH75
YRNvj2KCjrSEZty88Ulum4VwiZ3p8Dd7ts0uy+JLoz/f/VO6g8UC7lDorDi9fndM7FWgxWd7wXCv
KcPC8piqGhsGnKXHdPGCKC9CaDpId3N0LVK1Fcf+N00/A49HgHtBaIVa3l1qqg7F4Z6W7YTmTlyh
mjmSKE7n5JR6wC0mxMMmnqHGnubeiFVY0UO8n9NywKJ6Gyixb7qRlniR+ibHgkClyqWWwr5YHRSl
+g7oqzzlk8Av0yPG31Wb/jQaR4UdR5z9xTRL+WQW+6qKiacbb9MroH29htJX0XUygZFTu6IIpxBF
ZZAZO1mBjvn2CW/dIOJkUPV4mn7DQj18oOG4wYjzu3GMfamD7UJ37NESpW6cOHzC7LhOi+SUb0t5
xFfYkTORzLjZZCofkIzno1CmwyEQlrqfe2KLjYyn4w97RFQDsqNPy6bVsUwIXMxE+2egvM+r1CU7
fGfQ6hpCeXq9y0GWNZGYhwwXuWwFU4HTcnWxfd7BI+a1sIfobCIDrHeLb0m5hFWfdHI1J/lEYVh6
W7yy7lVWwvNaCssgkadOvvgzzl5UR/7R+EO/X5pOU3Oa1Ko+dyP38B+qCCox8b02SoGdk/DnYc8O
V+bbMnRTBi3Dp7FCY5cknL+6iifvRwj2gsCL9tcry9q1i9exEcngfHvfDzrY7ShCYVET8OdQiDBA
fWcIu76QL8btY8wjq3b1OQOZFmnOaoE9hgNyowe8bX0qVcbBbHiFMW0veErpndEKmEP2lt1D82Ep
eetaqkwxhOCWG6yUzwSDzxKiIsI8OhIptnvfredhCJHJAsAr+/2XGesQ0Pa45WZvgYEttMBIXzfh
vaN8/sy1E6a0WOyxSzOkxLe26dJP8jqnizwyM/TtAB8eMPUCJFz79zO4dRlGO7XMck0tdvSFn9Ad
gRkGcAJQUbK5X+Liugtn6jLYB8v4jyU7p+aFS9+Qz9v2y/bFvQDXeZ8cMtO4DBJOHWtooBHcCLNt
bxg3tELVvqVW9XrSJwMK1eiePvUpPRVLOET8e8Rd/OdSr253+VO4qBA/L2SvMZXHz40vWUiJC3yT
VgPHx3pJlqivKqQ+kL7uDrKXPJqnDuQC3ThTwDTRKfAFWOKjLbDlT2SrQwc47aCFzEDqF6EUKWVZ
r2jqtXVViLIMggLVzgWXFz46dLXnNAJG6sMPX4pvTzUJeTXQVXEfDJAgD1+hmdtbqh2KPfZWn0bg
GDijT6wENm/5z6qJ3R5HTnF9Bts8N1ABG4V2kMcTZ6ioHiA11HAeHz5q79QVc3k0/ADGD30AFi/C
E5Zmf5WbF2d9Zd3YkicOU7ODlDF9O5SJANB9Kyk0gGjS3bELR4Qvk53CkC1fhSgQmLXfVyvMePFo
iYAIcCrlCvSkXfAioLKLW17j/GmClSlRb/k4Orjl4HuzTI3fxMoOOEnGOWk08lmo5axPNhAIbmKW
4L52AG1DAdCrpcjTVsiZRr44YzFz4kCNwEN3ICd1Z7qRy0bUc4RKzbMz2j3LAkohpeyCVk3IwJxD
RmUlniDf0cQv4dEhMIjmMVGL5klbI/tMHXMTT4jtQeitF08SnJlfut9rwpmRHUOe6xC5gZ97LHoh
L/01HDZbPPsUc15rkQyeh5lONTH8q3JvtLTNN1ca0BMEsCV/kXI6NLwtvb/gCJY0Alww19sGqcsn
CW94/uFoviuqYMVmgW1gqm1b5/223uRpA64EQK9NZaDAMFszssIlW/nSQt6wxqCGlDI6z4ahsmgC
Zv45df3DPoYv0oHxs0W2MkXT6wLuxejeYDbrtqkCEzAiSrHRGgVJ0utaohwiL1AtAipyx5UDXewF
LU+XZoFb8nERybfNYik7ohdTElGiW+oNH4+NY/CiuOIKSRLZ1rgwpn7YxtZj1WiPB2HhYXusMXmt
bL0Iy8KSPYgwUVWW8I/1oEwIA097idDfG6qSjZ5N2qloA8M/SyqmwWw+n9/GVxrZ5YRZrMFMpCAP
gMesey7bA4P8zJvBIJ3iPxFr4VRRPku8TreWFay5e1rkUx43ek0cx8BVn6K4Yx7Rgdz2TQrzOmci
tXILTenMoeHKVmKAcMYfa68/x7c8178eZ9ajFTj76uech8MGwpOhl1BCP8Gimi13Z4hYQlQhgT2d
KSjq10+vk2W0xeFQ9ITW0zdjEz/Afm5nbsy+XwXRb3ALzQMecwiTLSgTrgROL7F6gTqluGvO5dBs
jHzB4QLxhv4kStoB9Suwe7W82TjIc73qGPGYqqWfjAKkv2hRkefBFLUm48X2FpHLT/0CiA9ELmaG
494851HKB3sascoZCn6PO1ltJvgrPxeGPqH9FsNPNB0ERziYBx36VDCNWKfMFt0MftRobgaFA8U4
IXv63D86hmnLkBa6xYx16dn6GmNnpkbU1PFTFIlNjFV0cEDNHBdzF/gB1F/I+822f/ZsKLitZ3Yb
crSnZ/Txiiuwq6VTCJjlF/1t++xyZI4i1FcQm9N5QyAoRSbqVLm4S3i74D6gcwv8nhO03PHsrORp
bio+txHiNU+o82SUNGR8rE3JM1hUPGoMKkIClSFhomejI9yfG4OnZoLj+pKpaCdfFNhrPz1phw9F
PhRtHEEmLCA8vmkOSf2mKXq4Maf4yvxaJwNal7v7RYy4I2hmpNUS3j8hKxFVrGd3MJ+WUXkNfgN/
UqYj+6+Ifsn8lhhwF+mC6T4olU4guCO7KgqljWzXNNjzANecpIlO+QwxmOSEdjokMyxoAZ2S7926
cSF9wuJP/R8+y4q3gqaYPZYW6j68psr3D8dcx65MfpNteS8lbDc3gCUCToJoc2Wmx92WKkeqrjuj
9kQQ0laMQoK8q+hm5XllSMcNsFooae1uuvYnZRgyCmooiGgHU0I41lu2a7jCl/Pg+mkU6porUyn5
ZTY7w+eLf9/j3l+3liwcxMsNDl/Z7UFpTChnNO0RGaaVbZyUCwVC4E6s5r9xzNs9HB2cMK8JeUZE
o6OMuYsBo5WjXs8AN6FT+vvNVaqETYciVL15axDnHFmQOgq2IIVb7r2Vn6Lek1tMi2vykW7VXDNG
WYLTWndTEHiSnbodFYgz6649HXPQyzqzKJjB/rXhpXmi1h58+z73h247aa/7pUfgsbHcK84nQp3q
Qd+fJa82CaQFMYxJLL/miKf68IxX1/to3wIZYd28f2tUyiPif2L+QIF/+8IXFA==
`protect end_protected
