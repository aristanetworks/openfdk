--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
cTkstplCNG9bVoUbyIOq6aT34sdRmjNRLWXNIOW4nTK8y4WNUUhJCxbPBYVlE6R37AVPeZDDlJ1I
Wrm2ia9qWgGIJIBUltMpSYxINl8r7Y7FNzzwcxiKJg2CRLi+2P4luzxP4auQrnxFgJtI+PKcka3b
GMxbp3wbFtswI32OCHMttJ/eYAbXT8nDwcZVYgk3qlGAsFX/6IH+XT6nrZ9tb5ByhKcuU67ZOQ00
AsGSM1iSahPyfvTDOhx7FuhSTHZeqp5vAeKZ9X6yoRrfIRu64aDsQHClERGTM23E5b+GT+3W04lc
j3/4UU8xvYhcnby5Ap2upKW0ys5HEtrM3VS0tA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="RdkG/4N2xIRD1t/eGXtbhxVR4J2auffR6v+GX2dIK4g="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
gJOn11Y20wm/CRIjTp/RXhLhfadu6f7m+5jFKlb1rL5ruiVirrwlb/xZBuKnpMFEoFaDceJ0iigv
peLl8a9dO6EtiRTjvCqGrF6XnYgs2CYDyfGf8qMsaHFVkYr+1/J/Ljb7/NvL0k2lHb+tdr+GoDPm
hc5C67kBbye5WfefbO+Gb67BIIpbG8KRPbzKKl7aApKXGkeXiaSQFP9QR894Nv+LSWniYROwfSHU
5feTi1WpKOqPLdhx/FpzdjDur250zMaIj/yWwYWWreN3MJ5xWmlJ+8mvX4fU1O2J5ZgCGks+ILe7
lsgSa1/+8/lhjOhYf2eqHd1oNSIbMVZvHlGiYQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="HKd6icgvlv0ldjxVikzFhZFqkSD//sqGAn5+lKugT+M="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26400)
`protect data_block
6VY3FBhuHjP/XD6z8NFJQ2qzOZWeba3Pfnap/vRtlATlluuHH/ypTjjxpHBAYrxaCHoJz2k0RRF6
qi4Bg0P6f1Q26EhCepyOZK17r/BmCq2/2wNkgkTSnUvfsSZ5e7taDquKm6F1oUgg3twQ3TvwNcRJ
kfLdT/L0njdGDFb0whdPEx1N9tLu4kTZua2pcivRDewqmTIFfMK826arktZ/+Cw5CBoLYvbLfa6M
OQL5vRsGSKAbjr8Ui38JupILZvI+V6Zfv3114a2RNZc1GA0ECPAKlGMcURH9vma2eBaDBqlLz2iv
Pi+/OTtsQFqqCZdGOQ74rerAYRNldHdcTbmrdAKAIUbhYV6fNYz9bXeplhvVFdi+VKj+8/9Vknnj
5+A6NaUxPQGKXngFDeUDokULq1XH+ULiA7HYLT2M1WfG1bL6DJLmOW1iWYWiHk0cgCPu8H7gNnzx
+cUCCrAAlK/vdW+sZ14tCRnUYxK0P76GuD9f1RAZqOx+yxNZuIA8XkVnFlfucfutPE4hwMBXWRKR
Pb1sk2kQmwMYGlShcgJMTh5gCkztnOvqA1LdUXlksbtMEL88IsIEJT2CADtCzsNpQ+NrpeUXTXEK
zwjEsJ9k/LpJnzv0ZVv7nw1SFItIxFB0mrhLj5uoNhzzgkJO5hqLTnnAxSyiwh29jRnhZ/RDl3dU
S/qJEPr9EMk0LCbHfXN5xXZj2xdC5Wl42//Yci1xJ/ScPGPF0HQ6SRdV/CRICl2uAPZNFefMJEoL
hfqtO95QllCcGXjhtOohPgmXG95G8ZfrJvfuJjWQW9GWi4zx5vRS22JsmcL5pqDSq9llLhPvc/wZ
Z3/57csClOAQrDEO+1HQlGzagzXTQ0Z/xxLe+J1v12gX27H8NVwRDaBU0G/b8JT+oqFOUM5SK0tw
UStSUxbXfUPDQMB5ZPsJvqXAlC8s5jsI6qQROpT6+fCXBfz/+uxbJ6VihMhDev6reWGpBYkEvC05
NSwlLrRSiV4Qdf93NH/xrJI/CixLGpCanaTbkzldkTtg7ydIbKwY3luSPmVE2OaKkjNOQ8w+VLki
7oASv8JPa3LSDDF4x/6yG/vpgwn5b6hymD/ox/WKSdmtHEwiJam12XPeray5K3pUYCTNYOHwl/bf
SBlgS8MdkdPitvhVckeVNHJTB60UB5j36ZERsad+WgA2yUGySG2V70rinMwuc3yQ8GIqwkFc1eH4
0ODfVYwCZkl/J5NAD9CFMCzwJxouWkmLZiuW+BvI6sXwoTwApQ7DZxuAbAasSAITIU2DbLo23BV7
QLMZdXc7NNKFMVMDt0tMUXJKbV3mnm5dXB9vPNK1WQ+jRjkWNbGnUXiCLsChIOIFrKieS3zERj+D
kz51R/Xt4ROX2fG8tTItdIlP+QAQu2XIUKT1dkuSZiWpgPdPFEQool13SKVaBoZURpFQTCjEyt/F
BD9/l+Jo70qwxVChqqhpENCT8ZJKWM0qNrGQ6+VqiJhJC7cGknmPJSZgo9XNBRR+SpLBsUzjCIYb
HGqh4b4kQ9Tcd6DXK93CqnYG5OM87JDjtc2Aadvdd9in9bvucd4mirqMgVddZJBYV3s8rXZwU496
uJrrAWdntV/iw+7lgiLKpzJyDCEtGS51ZwIN9k0qHbxbC1i294jrUhJ/O6biXHS2Wv3tqW29gjYv
Tt9wg/5vh2xXQ73gXdeD4p78ytgFzG2gU3AbR92NizbAyl9jGn132YrAGejoWNca/pYv8LYbQWS+
oLOl4ZvzN/gFhJ7o0TzJNMSYq6B90AXBNkrwH4+S2kDWTrVrem0YdIeVKqZW/tPRZYkf69iaRWbo
Cf5KdNAyOICY7CnlYBfJQV6hrr3KlKWLv0s+eFyoKLYBbXxgNfdLSIv6OW/CkaehiQrhgsvTot++
v4XKp27kMYUSV5avW6ttuWypbwQnWw6P/2ibNuXSPYvIevjkt2VmXNGRyt2MHggWWKmGjK/PwMCz
+zOUUvbgnHVgBwRk2LlouLtOjjnuqF91pz3lw/inS0Lxqq45UxRsKuqQFtJIIP0q6E4RW5KOVYdr
J31l4k7/vQBAzJa6bISSRyNJwg9Bj8YI1FLoG7LvA7dk9XHvsFRxyHvzjWYv9MhhbP3FDcmq/UaB
PApJUR+AoUEb8myMCJLNOmJ2uTpqOw762hNQw8hbDKyKQYBXMiJgV9lExzlSu3+UQwwjNNcOpSX8
7//X5ZDoGsxaHAEpfqdwRYUmjywLHuS/87QoKQ9lQysXrN8FVFQX4e49aGeQSUaX/9Wkw7f8WDHk
8c75RkwgE5Tf81eyl+r2dCsvlqQlsM8Ef9hdqq4h+RlGFsKZOl+NcSNelNozMBCJa7XdEBOxT9El
ot2lA2edhazSMzGGp64dWol2weT4APLS0ZaW9oCRlqm2nU8Ym6Xm6/4JQ3J7adSp+81wOPF3YOC0
rbX0PhnwjKE3aStgUv0c1orL3A4wsHQNdQ2up88XIRrTR08JuRWyoOLlfI977hVElwZbaR+mqd1z
xWvrOWn4oAoVfmsn1b93Tg7gWqpK/Y88jTY+8v1dbJrxhCe+bphHarCtpoumWAMR7OV/+52g/Bk2
Ur2uFw8vRjWM4fewNc/QikQdWIyrCQFmpamwGjsOB8qG+vaLxxblTNlIcFjJzXra+mZAeD+vU8mb
EzD7yoPhTGukHyrk37oZ/bEIGjXPb4Z3bgV4CUJ2+wdP53ZNL0GjxCmqeXpVHmHy3SXK7jNttA/R
L0LDsDT56lsWjqR/KhyBrPI2dDu4YAF+hLY985c5raBOt2mSHSn50Ol3Ym371u1pfdMeMy7Ogl5y
2QqCaI66djOCQ3CaqNft/pFzXJatTMDm/PE6MKP/2OZRzKSPHRJoFBtW+olpWyJ4ONhqjgT7Mwyg
+WCv8hUH5kiIoyqtbmnrJ8DDsJxj76vnmW6q4pY5Y5zY3jsX2CaaPw+vVJPCaZowwxEXmfvuxYN+
90mh2hHzKHrEEziqO2NkTWIkChUh4hUUUJgfYH0HBf+C25VJLX63z4MSgjqoevXTsfTeFM0OgnFU
Swh61oXFqGTVKRWcYzF9HUvxciipmn4HK75Nwql3XP5yImqEwNAOt+r+HrA/oBxsncisqpgOL7cY
OgrY3HKCYmrBNtnSOGAVaxGcgO6GLY0mnGgdZDCTEcfgAhSnZ4uzYLAfzoMJaMv/oNmpnXQnDgOZ
X5G4e8WaSMWxcxVsdQXd7UpVP+8h3DYdFCOKi0G1RP7eWNZbJCUn3827UTvkpcRr53v9Rl7HkMNe
Ht/ycLF/+elSlIlWAsvl1/VNeWzQF9Mq0MiMJIG/jhGy77EAp9MgRbkSMMjOA5uDHtSe46k1yJHt
pmMym2CEs+QvUS5Qnch5WlcMK9JmPr9zqYoNzSlOwVoQZ2hRdl6WZoMgnZPHgT1ACZNFfoJuK7Y6
9nf26fTHlMb3pu+xw64A66twNh1mVARdLe9mqmVAFjmrLm6c38UUqg3O4VTpPAGP41DWUnpTd3k9
4CnDIfyvQfPElV7INreKYCucGmQe/QuhndL88Rx1CpWfxoLZEwN+88VMq8ZnPRjSVnNpC9OBbyfQ
zpgWBC6SfTDqbAEW3I1D548xshTBpDLOd9IZvXEcrdQttojctH0FzVasldA5tZkYm3eNBx7ESl9m
8ta8reYtx841nyFiRWOxnCnQyAHX3zJ3mOy/wwg0DWkD+rvhNfa4rCzbaJxYxokDlCYOcm5R6kDd
wtc9xsyuCy4KObxzE7xl5Y7bRVijHXtv/b6ldxvxckP3Pp0NVc6YVfh0vWK0op6UInNwgFiJZx+x
//ayzha+maHddquzr3S5AhSDf1DBjHA2A/e73ZWZ9LxKOOCOPNy6gt1L51lYlYY7q324H0mjBB61
YxO3JwsrWMNzt+ak82v+QnE2gMgrRZ2Co8HX1KcpR9bdURwNl+jhSIppwvncjw14uIyqEgFSxxFc
z0H6Lskwy2GT3f4IcsQB3Sc6Y8tEiRbB6pM39iEBtXNSETbWRiZW0gbDa8Rh8MgU0gww6hE6iyg1
Nu3lZY8Kevl6fw6qmZw4HsBBarYOT6OE0vnVhr+ym2JuRb1d8qcs3/fJ42n/+0hFKXaDJoH6V6IS
kLPDWjmsLlElVv4bYvgC5u7WrOIW3thPNlxYeiR09ej5Y6NrR0prBbd4du3lzu4EhYSuoEwQ8ToN
G9ggPdoB3qyFQZ1eGs/MD+m+y7mgWmc/2cRLo0F9Z5UFkb8OzI0s6d5hpHecZFKIRixQmlpCPkNf
izMGIxCls2Xmef1SwIS1y+oadecf6v5IWLNbCB8kfbyL85sGwPWbF0sSo+oUYwuloCuLGmHLpNSO
7vB9dvGxjmWAPP2YL6MyD29TrTWtIu7aQafG4sGaqGNZ+ei2Nr4zbOF1Y4nvvVoHprM1/lAhdfQ7
GVnNjPifUSs4+eTlDIVzW3Poz+EcB9JDQBqS0T25uCWrOFrfEI8sjiUU2JlDFunnjplQuO1uyJ3+
ppG51Xi7BleIItEMiGO2IQ7BMcSip+ulJ5nsmSSM234T+N43zwwNJVbRveyXQaAEm1h6kRR/4SKA
6VIrzGHW44pFeU2Xqn9Tq7vvw6GKdXVTxFv1T6LfJ/r0HWEHxbUVncfBb8DR5EbguBW6ncw8a7xO
8mpR44SbmtD9JyUgieMmGt+gXqTuuG8YFedGhgMTB8uAkTQ+eCiGJdKA2ju3KVdtNPsJoyKtWZ6f
g2KIATCipzJBToYqPlSf4WyObAw8755sT2wF3Fng+EhFODd2JmkxWnu0+Wp90ftU6qzpoDYyfmHl
QcBBb/yDscUy8P/9SSVZOioj6RqzlLH4bSWruk5cPlNrFW/BEdBeo4etgWmyNRMcuj7RqpmNdJX0
L0z9+PZ2pjsCY3zY8Ao0vpV5hHp9tAUE5wij7YwhIH407jLAwydWllCZfCt12o0kwWU5eTSI1iIq
YXdyeZtM6us0z3W+N5U9Kn1cu5w0ACOBggSypnQbBYRbm5GqFZIi/uHVy1PYh5xL8CWqSzGLgI58
6O0nGW6N3FjHdrInLBGTZPJWvGr4sIQoo5ucLtBHQP9JDYmBes98DoUhB10uNjKC9yDZf2UZwnrW
P0mtOPVnZsrtGt4X9kgzimMRkn7CTRgnDl5bdDj60XYI6gfzVxbg/HJI80u/MZfcnRU/3zhmmBLr
c0/gwCccPae+sSXJiG0X3Qs3/Alva6M+5O+FtEi312cQmn2yzWCEld1bFhmdDOw0VkPWzfTjo4QZ
SkRgseJM1xoDEchy0MibTKIoMF+k7eAw0S3Ux2yVejtUS+B0Sq/D+5lwky6+Y84ZIpGmyF23neRQ
XUjuxIYqqxylMyfgZms5hWORNozsNnpDhkxnLGxC+liRcIEyP8Zc43Z/gAWC/2Kfxvhw5o4Nqjyp
v1RSdrBhCt9wXXj+beHNHLLUBjWZVuuaeScFE6qSYbqWuld+Gnnno960x4mhVNh5TdBUrqLkmacc
Rtr4MwSugvJGB4MC7q73s2gOW8UtrOXnf1OsefhW3kXHuZidL515Uv6tspluVjMCvPAkVo/3t3cg
dVJxo9hrukGcen4+rwrLrBq9zYCmp9Ms71o+72PXk7d2DABV4ePeud2Dh6+jnFnkDr0oQ6coXQCD
v1G4kFZCocYjw1ZnY8BZd/6wjmWXmlicVVgFWjTi79haYeohsOjp3tqW6Lb3Yeo8sVUDkTG+ZDIn
xkUR7QXqt+GZ4e/0rYXfMSflStKzZ2+6vx/nEw4j+7Lm8qqFF/7OxIK1uuv5PN4i/7A3WtZ9zIg8
nNgl9KT6DZ3KDoXQdDIy9JOKEsmoI2U+gIhaIsS0etLtRz64KrD1iZNJjM/EzsOvRdQu8RBLdZ7d
VdU0nR5IgvU0h6EUwOJd+rh0DazY1M9gIS2nN9NCu4VEt1qJpEpY+OAmPhBxVQpSJGBQJ0dr0SP/
wMEGgEU4uamURmdokUwXNDcZ4k9ZTw3i5fIlQjIV+TsgxdQrRGKaItf0Cfw0FpgJtv1lUKCMgYgo
nnKsgf7XJkmGluS70WrfhCvk5otRKUH3XnQWuruphe8T9zZdr31apeS7zGW5tsSd8SU/l96tL6xe
NXyDGL5xjzai8JDOY4J0s1tGwM/KzmbgHevmPLHIBT7oHzmJJmNDyRccKWs07W/jdHz8EmPThFMJ
QZaFXP/uXKvlXKXitPZ1NWwtfy87dNyyw7SHRCglamYPoJtjjK1XUqCXhPqtWQGLBSJLkp2UjgKF
rWWIQLNlpNVl79YZ378csggmF2vu5NEgcfRu3h4Fwmmg/hgGc8lOQgHHNx+AFdRR+4rTd9FKeWGv
fwSCVJ+6Lon1fYJsY/kPv8Z8JAQvDeCFVrdgelyw2M9JKo3Mpv19Wgvm9Htt7JOqYzWfnqNvsDWh
0nyWXVqcPtOZrjjdbSnElYWJSzPDocy0EZ4IOTB3FqqdWVi2EpV4w2pWFQcpYmjutjc04y9QZuiT
/AYlB5gkMbuatt6XYkGr8gM4cn0YFDjVgoFWGVt+mwkfkOYMTCZWFjWtWVOieUh8N2Ro7XOafdAs
t1WFf+59OZ3g76gzsAdYJ30g9C1wVyr11Gz1xMbQ/4z7cfVG74K2MQ+Z5TjjPO1VE9R/20teVKmC
IuQPM0gVKdq23i2vOKPnHH9ksR/NgiZZiIPPpepw2t6KdGnU6aPbixYqW4xx6+Vu0/YQyQCKyJ6s
NzNDHSFI3tOe/ixDw5TF1f5Wc5QpTOVkB21B/Yaf6fQqJp0l/cunZ9pmep+dLyBA7f32EXu/us1i
0A70xA4XPtgA1LclRdYLCgXAlvvxm/a1Gg+YANDL/DIL9fh+SLBa/l0JFFOsNNW/1BBNkxe4KgrA
B1Yz7OTcnomMIgR/grA22JO6s8bWtowkrEr6OFMTx4EkpgC/Z6RkDapzRMePk5UBNEgELRUx0M74
Ri4uUmCp5l6/KhUIJA2riGl/eYEnRwU/OUMMNg+Chog24WS6nSCghUcYXcqd5CtCrxSoQT3QuwBF
tRj50tF6XjTl3qp/qZEonb/0UGDlM0AftfYgYx1+Ns2srRrl6Lbr95KETo6YiB+zl0FET4g/2sJi
55dwfLCsVZaJR+lTrKsRhmMttB0Ni076bTqgu9t9hRoa0fzwItEnBNYyddNroKlVLM5ViSXJq4Qj
Re1fusAHmA7eH+tldiucJJ4XcBNwOjlriC8oVYtnrRVfTojMcc6VuZ/bmJ68VWgWm6mioQ/wbHdC
poGwWs9I9+zm4phbfYL0fR1rgiWgoJ1b7deVxpKpA1ZE1XWXlA6MC+ULo1+gS4edDJ2aUbU+blJW
H2TeR6OeRiYP7kCNLhGLAFvv7w2fUNldzqHMqZ2ce1xqLqcjinmYI09Vj30HOQRQsiGnEP73jHil
qN+0y/L5A3+vBt1G9Ryi7/LQQJh54DhojIWJkmXeJdlBlxl/aEMILwFtO0y2DeybZisMhPdwP3v9
tw99e0pNdUig2Y8xwmq3KjoyaipO3FHfwRkJrpUGF6UYe1iAsLOBk5ts0Se+lsgUjw+mEGOrR3/5
PiDTS5hCUUfAVkRvo8j55M7jf2ZCA6IvdvfgwRg6+AXUipS5+ydhWvzKazZU4ZAuumCef5iQJswd
4Yq9W2eZ3bL2v6IA39Et7cduD4W95pKlKNFRo/mEAxeJElejseIKE+p1PkLOeVVViRHpYA8fFM7P
OGKEILvV+opml+0Tkomf2YPW/gOupiW6Y5Epj/ss0irU+H0PS+H29JZibfOFwq0SKyUH8KQJda3e
PWKwl4cW8d98U0RNgCdXL/9ItesswA3rKDomRrdXGmcN844N26a3TzFQIsN3pECGCKcZM0kNghxy
e6Qb2SQg4LA1Q94QLU0QNRGkKhjebLxRRfJzTQgBCHa55k/Kb+DzkWu+WGvVir0Sj1VN4MAUfZPF
3YhDFQ4x2eBL7DjD2errPyj+DtzJuFdA657johjsVJHZKb50X/+gAasKzE2pJi7LJ64zpFy5pbuo
trVOGxVgsAklugPx5F5JpJzO1YIobzBmuTa6d/EPflMAYnpfJlJB2srP15wpoA8BJTw3OtEo2uKq
ooZOezLtizumNI3+VHSXhSpCa4GRWJR09aZKVKTEvI/qCmproSkjqQGgjdhFdUpKvIo1ZPggJ8Dn
OmhMjfpBh8Gis8R4SkFBqLYz3gj89cOdZfmHVGXaifbQNxV537moCO3ZStWStzDFuDqj0iKVb6u3
FpJCl24qHlBTUfgCFbGPIoxJ59sG0Fm6Ob5jyV6vBNbfhxSYcf+DGFYNQ1TtBditeHVl4M5eZjZ9
/+MjmtyRCarx+IETONsvFIIunQU6AkD7qJLy8UeGUu3lf+HB21hRwrQJdbaiY/JYxpi2PJiQj3Lc
Sniv4D3j3IfHCgN/zHJFQlBBxjUKS2RDxO8sguz9csIQG6qmFiP62t2qxH74NBUdDvp3UlZK6isf
JT8glwDXJEEtEuzt0OL+Z2Be9zhU25ZxFxUhLJVqvk8C4qAmDXC7myVQO2Afbj2PXofCP+o6eGHX
VoyyLkqBgD5XKQVRlekA+KLl7unp6R5M4St2Fh9btHtrCscfJndaFTBm9UjZ47VJQ2SoR2jc1hEq
3pvi822MP84hH2GTMTGR/tAgDg3EMG4AhLtbkxE3RN0W9aelgt8F2hflQUlKj1RdKdbXtRKNEulz
QtfAjHv3woY6GaJE3pFve5Osny+0SVCSogEtLtPAGObrfRj40lj1avdwRT8aj0nqzKbrZLoVs0RT
0iiY3I+Oshi9m/sFVFAUMeBYrsQM+JL6AVTtMT8A/ka8xYichNFE5eXw5twH2R0NvFX98CxfTEqk
xezlyILrF8piVSceBu5wEIlTIE8ptJ+cOXsbogsCxFLpOyXTie0P/KcLfKTDrHemyouHhoqRlbpt
i4O+ZEI9HH6NCmdcK60sKsFXhH54w65o0ZfXKRgCDK1h9bD0U23v9QeiHiTMJxNgdallDNoXqI7l
6aPwA6yTWdZwOiXZYZDfRhBjZ++KA1pNWym0Q+Ryl4k81UwVWO7SCJqO0hrH3PhZdgfCaPQXTi4w
f80XbMHGTJHaG/pBnCOccZW/tB/qRNqkJyC7jhMCy1aws56F+rYjNpmdxqa+4v1SgaCIQOKa4Lpv
sastJcS2Lw4Tx7PF4BBmB0Jg/immiE49jovhJIe9T8ogHjoYOl1/6qxWU4kYLYGkc3N1zhdyEZeD
6MNBLbj4BIq9kxYaCsrFkriaCCN5Ylr3qCKkjDgvGGQzYTVHfZiAc7Y7Ntkk3s/73T1ET69hwLSZ
TE7DO/Q8uH3y3aYNZ/NDu4rdiaipm9qHc/RMp7YSluwVTdQj4rT/oywA4VA3Uu8YJdnQ+uoY4JZ6
ScJudL3G3cpxkm+wvo9nCg05qLljvNIqyevfTF/8WBQ4c2e0z4mMfBMQPZyF2P0aQDCfNM89ff+1
i/6d5gHSJSVKKk1XivvLicEFeA7aJq+pdfqupykCL3Np+WpWMcgP6ZeAkf8Zj0Q8M9+SRPD7sYvL
QtQCz2CJV0hDvmeJqA9K78nu1ws7XbzyaPDbKiXmt2RFy12T4nqcu9RJEFtbOGJ7GYENuMLhv5k/
M9BsKT31DiK/zqev1AkWtdF4RZ1nZiotjm7Nf1S2rv00aVAsgqDwmc2xCfMMf/v7tryHDoHW+lde
uXOOn9qiSJVLKqKQQxnR8h3DLrC0jNy9su3R7bdCj0Yalc8TcElNXDrU3mi+4r8DbMZ2tTAy0HnR
jqftfvMoUyey9xnrLmmb87JPl++gQk0McVQC9AOme9g7xhzsK1qQblQ+1/WhP06WQC/0lAeYxk2H
Nmbguw/nZafBvF5476Z6r7k6KFkaJUeJrnxU7x25pjyM2D97sKAqTc5ga+96Vnokzpg7xNIrX6xr
+vwysMr0Fts0VLkkpsY5fB4PJPIzc0dz+RkpUNTTSSGB65usMUehbFXexQYpSj0UU3kLk5CPHOzR
2jFuoo18XoWV7BMUx7eM3X37ZqB80PU/uq+uWQZcRs7S1zdMEBNw+zKWD05StBZ4AAPrhHNsNQlk
9f5p07ryA3L2sPbgNYvzRckdNAnaZKpLByOdNdnxChhXKDqZ4g7bIgfuMfLyMlCzmOHUAgdK4wIN
QLoUztCGtZ34vNibcJZ+KdhOmXwwr2pFhKP6zff5s+Q2G1ZU4YkpUwU5KUnzs4m2SoyImFbX+Ng6
6mWkS/HzyGK0w9u++bZTGaoY0URDAbEnLQ1YxMfP3gNrkz2t5WqMXFR3Rko9bgTJTGasVBPOr+Z4
NgNspwgPXRMW+SzEvugC4WP92ncG+nglEx+Gugad/3R2E4anUSz1VFVW2vDiSB7DrC8sMWmHSRNy
cU9sojHzvPfMaOirW/pHPgEpFDrgSjT3lXnSCDqpK6G1UfxOz+CuCVUpLUjaZ9QeaVDn3xGEAvmn
cGWImu2WjGXE4rDAKshVdSErKqy8OPE9Wb1VCSAh6Q9ree24wuC98Ew9JZ2CO+IVH4wJpHdJXWz+
EO0WDrcmScsHqrb1A8Fqy1SQeBw3jOvImvIjgXiT7i48upop7u3s/b8u0y865MxG3ybsXcRu9h1a
cN2sYTs7AQz1Fh6Grk3t1DUDMEZELeL3O67uEnQkwWF7zDi5RLUetxAU9GZpTajZ+qrRKj4KnOFX
muvZKWm9M+YhnIxjQ9SoBt/lJo+kuLXg1kZYL6RMUQJexXqiiPYvOeMslIz8687oYzG54pfdDWhC
RrJWh7TXlDBKGLZ38H8Ge5ZE83fLhQjAo6cmIklnoRVbbRHK1DCt9c2rGlkzpcN8I1Iq1faZ+Uw+
N0vUKNInQmBgT9bGsI9ejwmTyucFwtUrXGQyOqq3qgvlYjUiP9nomRcKvZ6h7QG5l+33r6zMmZR0
SrIG9xS7l3XvLV58M+XmOQl5RCblGdwH1fKGm6CRg/kiWnHnzsNmUEuh6radMyISVQYJA71x9J7r
kSINHbRalCvYnAS00S2TdNg+TDr9b6Lc+bUbGzu7iCYwRhb4ivxj34IK5VHPqNHfdmDeNapOXIZ9
W3bydqulm4RQr8qdbvJlJvZM5as5zYRwxqzAZ3pfR+ML2vnBTM9xRlXk0JZ+mT/polg9LLmK5Qnx
2TrPhSUmoRTJfifT/UrM8RvDjtX1CFis8t3bnNmjAFmxz1+WLEsr4aFbJtmhsoYKd0FR7cMh1AJG
3p81ogCBwSSLcnm6NGYK1EnXiHMuT7IvKFu6inTqzpf1nuigZybHUy5LfjgxEY3MkK7LtloSLuXN
cvl3ZHnAe7a9EaeXhiQw9SuvUe9QvmnHBzpLwQVT1Pki/GrCGSDBUnHE+t94xAH6O5pzhK38whx+
8spvmCsTQ7b8LedNd6ALLdWLTZIy6MO791SKOlQVroZ8xCYxPygtYHhRWHbtUyyvxaz72mOMzB+e
ui+HiFmH4wq1uwwHvmrdRPnopkiUYHg85e7s1vJXsRlE6RGP1PZrAUR5yXLAH4xHk30IWqvoO/AC
1fJxYjtTBlK8kZGzKtugmqPupIsUGcfq6t+y+Bi4mUC3tjvuhEc9Icy3DGcGRO8EhJzUomaeKsyl
VnAhjvfV68T4TN6NXje39ihfIfnzLzSm5ZiOvFnHq8PsFY89ZCYEw1bGHDB5fuaV/Nxu33md5gdE
Ax77XGFoI9agGYpjovMT8u8GESGiJ3IZ9wKBmyNEJIf8Mevkb/BIBcJQp3ZGXHLllXk23MpA1FQy
f/RPIc5yTqIDBpdyEEVIiVIQi0uPEY2kUPKco0zuhctc6dgH3RyyYhgX5P1Y8s6GDtGnNKy+3Qj9
/DBc0+cIX1/HZB3djv+LppzceCDgDfKth2VuaXBM3CkMdN3/VIWLJUfu9T6VF0xkhDGwQgZjPrz7
QBqAV99SFjiuiV1zLWzSsfTp/uut3y9iEKY5ndpAlgy969BWsC9QpOwSdfJK0cVEKcG/lisaiShj
B0I0tY1Lk0flCXwRq5ECx+3htxvnLjaswRddpqtxIlTDjCqlnNHiDLNDRloqOspcljvro5xtpp8H
l4WzpBhYFaoQvlqtM9lqAuH9ffSZKp9NrnL6bfr0e2opdjzArn5p5MLVVS0K+ABzLDE17LKGHImW
ZPtt0Ydlewuxy1bZj26kzD42zoSndAS/mHX2gR5PDL1Ln4wfSWp+HBTmQEINmfqkj+iHltAyP2Pm
gampfsX5wmbJaE6jau5R9ns4J/sG/VApVXTrhRSp1WZMUaFH87YnO0tn6ja9YkPQOjikNt/lFGkT
0hFI+mnAQpK7rkNaYqtnGcxs4fmxgAPslHjgjF7Y1ZS9tkHGLO63JbszbQWdBIUXveHzB58JFsRE
uDqH0MQcvbtekp4qQ7RZTAnZf8XkxsjXDBpn9Bu2tnEcdpJV+YcyvsZaasK9G554rnQUumF4JdSg
wKZ4LF4aiC3Y+3b9h5sS6O01CexbfIA6Q8bzq2b7xETuyieiTZMERpRJX8Izm9Rqe8pA50F2DgeW
gcsZd/9cyT+T6R9QOT5vOIX6Yj3lZWrQ7DBAk9aL9OPLovDPhNylhtBX+kDfCQrLSeTpSAXto7bF
tamW6Vj7R3KeZDa7AqyV3aXBLtrxxLmQieCLMCVulxY2PtUy1+pWJDwuXIEmbFJAB7bowBVu13Ii
5wakH+by1Cu/09nepv1r4Pl1HeK7Vvdxs7hq6fUwtsvmbJ4bB9JiQYZsY9EJ5u2sEl+pnfuGS47F
GSbn7EGdHJTxSDP9IQ9ijd+wbLPJFQXVLvW7Q8MaxdvCb74zDBzM6EdWDjjK1AKO0ybS33YkDXE4
CkizqgVBkb4K2jjhMi5vvtN7G6muq7xv1IPhGAddPpCpECFiFleMth4XZOt4Pda0AbuxQU1rqkT+
ifI1P8WNN/iIzR8ZTyamOW0VGLqNguBaPcJ67RJuaV1IsYESnryEsWxQet8Re+0eUqDxH8c+FCKf
SP03AAgg20kPsYZYF+VbXLm0HVeOVi9XmC74WAeDyZY6d9dLsl54Md1/xtOagnETRxW3j2o5zlsI
8cH1QHHdyYZLPrhVqzUtjUgcT+mloYpNsWjSiI0pF2ruAoSN02UtCrezQKUaeQy+RFRjgpacRew9
gSO2qDKsU3owXVRuArbIhpTEnbnd9KfT0ALzx5ylVTJC8pbtOBPk5w3P/Bkk1FOlt5a+i4e36HG6
hhIOGwN68Vwr99UR/ssq8gFoZ1jO24yZdysJRa76pfq4tywgtMOjL25qAx1uPuVeL5HyeV8u5DYE
TbvMup0OQl2Za/UUHWkyTsqfpcVvQWP1DiAnuDRLeQXNozdVk5tbvtcVN963NJHHnRSyhQ78T9Co
2n1VO9C8abDINQiMLaIUw/TSgdJm7eqzhIXME1YMAfbKGC7E9DDHKxPWMxUCRKXWXPnghLcZmGSx
7zgwLkAaTbXosA7d4epv+xDPU9AyRrtDrZiwhtP/0rKYWojHAExDcvFjT/EfJ4TygQzKtr0Eark0
nNmlY87d7WcBg9npDQcu4plkUuGJJLHlCmRUkmAL2Dx+yQjVnTciK243UbhfcBJavYKzD32mfwIY
rLO9rL611mSAEHA7TtEP3/YEDQmfP8Fr542Yuy1Gf9AmwN9Tdqd/FVipqid3yCRar+I0Vnnbcmle
f7V2ScezO1DFLmoi8fewgIFYl9FwfUiao7OR2fa1/r4i/Tj29tQlyrAeFd6ys/2m+VC2NuNxJ389
XNLKhJg4GqEw1ESVglOm3nio3tPJ1oFRkmTGz+ze0scN8sDb1toS4kT7juv1y0JnfFuzEYI1lDMz
phHxTdsWA7BWhP+o4rd2FvAWp7YyM0etIhl7lKcPg4ofJnxM5gCqmh1mMljwqPNPVhDvOGUHGsRk
oA+uiURxsLlv6eqA9TDparzMYgQ4Jz/T9TymltQNsmeMma/VESYp5SJJPO2X47M+24MgNTLKmLEI
xa0kIgx9eA4fFdGgo41qTDdRXLMhy6+7BivyEy+CgH3uVgUz6R7Qcp8TzNFvkYINKKViVvmxArPy
hTPohp0HzOluJFmvC4z7nKb3nd51TiN3PSygh1VW+FhYjgM++4cp6g2ZNmCyo7j+imeZmYsTEvP9
b7nXQHcPt6w4B6xG1I+ahiiiM0S7hdbl38Wj7D4gsyEoEyhv3VMm/Q3hF4Et7E2PaKLCpuyzZyIy
xEh465asa7KG2TG1Y8gYsxV1YH5S++fuL7ROUG9VXsSj1fEgCMS2I385BV6Kk1OU6F3lMhNEohj/
iwA7zXKnCnziyBIQxf6TQCENAytW/YfSvL/nb29ERzC4KShH153V0xG6SLdPRC/Dvl5mI9A5cpTz
kmhnP2O4Xl3h1AuRA5OaTc+YMlq+uZgNlcvWGyT2bROSmDNrDue8UY06NbNRZq0VGs8CUrRxQM/m
SkIHx+dv3pTt4kbaYX4yzT2PQZXfvijBoAyPHgQuAh8OPRqcjZCvCd1ZRarkMuxf6PFhtzM1gwLO
FTfaW2w5FHOdqYBBYVtjduIfOUFvWaXKDpbCGu3oblyLV5EW8V1hFK0uZIUF/3mkq0cLUjqE4l+E
+XgeGpfwk0NSUf2WhgtjXgSW887zydUfrHmcJimHkdT9d2Mauu4YhwAJXM3Jawhb3f1ReESEgfEr
1eNLBe2ucRB4Q6Gi/dsblHzxYvLDH1rYmpQ8QnKeySeDXl5DxQ2dWWiRAv8f0Md1ihqxTRofg3Vb
3YrjaeDrQyfcgSqDQLHwMoGwIS9Po9+w3m5kwYObhZbltPvUa/QqYps6YWdi+TELOaWF4/b8Sr1/
48yNor9WAkrDuRP2olqkWveJbZKngsLVqBbqpxvGwKp26NglV80eVlLAeZmdEeB3hs+ovtjb4crt
pDsVmG6PcLHr1NAaw1Sj2wfskzg7v3wNwZNBYjm2+cYWUnX5IWpfbqkKCQi8lw7TvaQyGwiqogAi
LSKrckF+w7cJGPmIH5B6jaX+JQo3mCiJbj9Yl0hwLIcf7G5rX9fHlFMRj9Au3LimwJxDaDp3jHkV
ZZ/rSCEOHfr01rZ9F/i9KRHRC1Ax/pYO4UpbYKut9u4IG91Hjzy4qZln+XroDuhWJPGUahBrsPVI
F6sg5ULgfql2xw+6a4qa/XcY0f/CWlW/jrFkjdVkh6k7OonVur/85aWcidX7yDll5+T3CJ9wj9nt
V5TD5JhB5LMZWPShU+ADysXx76SxoqNBhLaOiimeJvVGVh2LGrQU1JRrs+jhkzUC2qOFNCIsAMPK
gNNxpqzU3X0FniLx15TMIXwCe13lytBFpRHzAkoAUbliuEYagX5mYHLchwxTJ04tYXRpkMWUm7nl
qjYQak03aba5XGOnaGLYmfvLTu0pwQ2PClkBwRo4h1UTGXBsqxAtE0qoWwxwuoYLYm2taz5zH+PF
MlFRDDFdc6Yd7RHpv3GRUB6EYq7Sydlv+cBIzZkICJNcViRfO6wN1SKoNJvidjifbeWUgoRIY6xe
yD4Q75VKabb7XwzROO3cxzwzUlF86KKFzL3r50RnnDkgeduet8efMvTtrVxvx2x4c+9szbYGXXTL
AlC/wEOVDxuJ845SCZsw/Z8puSw1gl8jHOKfKWBlLrOEbets/PvNpoIvfCVkJnzf8pusL31TeZ7v
6z2eU9cMgvKrh+DGr2RyP0bEasaoiiJ9oYCryxS8qEEYkL+R5mc5EYN3dPew/vK/8o8Ndk4k0p14
JIE8YjrpXwLCIimM4TWOxtD9QcI7AZCC6Dar3GUGx7BuTJolZ+CHvRS0ccztSQI00il46c8aOAvL
Mi5xM4NUcBbToFt5aSJSD/k8bfC8x2xUrz98Bzyf1mSv+rtlmfFFjO9ZOXB/jAvb5dP50rVnm4RG
/wPYlhxj+N6VKkA/XXIRf+ru+FwdOzaIbNUyHvdYhnPBqOHqZnuWV1Yb/RAWk5g49aasXkkwg27z
N9WZFiffIs9T7IJLmN0pP038YsJaQ+0ub6lL5JGvUzbGjLuCw9GvzOK65Bo4KOS4RFjoDHAXm2bJ
6WlkH7VyGyEppFy0xd3GcqMLUtRdcDsdTjwrfOjppqFvdZ+C2aX26MP6pA+KzSUl06zXQKQdbQsK
8EdUCnQp7UHmmCAY1EMzWIjdUAKXAfPNuZSIPnzU5K4CzjkhDmYCk74h1xmORsdVJ44e4Mrq6U2Y
08BDNJKniT2CQr0Em4pagsb73XCuMgtjEgl0JYvrtd9ohtVwZ3OK/VfYfSH4toctEkQq0sc4ErwG
xxKsXcBWmEF6luPAO5Yj3rIuc9EO4gTb197bqk1xdXlfj13vGVnZfNRF/iaVH2psthP8KH74e5Oo
yjSFr6XwHYztFT9RCoIlAKbAyr1q8s/7n0hHZaJEvWBNmoAT4Jw/ib7sk4KT5jEslDuOfMR7NHjr
RMb7ZwAAzRv/yDTCrz39ntqe/g6Zo4BTuPo64bN/vZSk5wQoZQFoZ23vlQEE9SP1g3Z5S1Ezoz91
PPs53Rok+QiT+ffvdxoBLllKB7qHGNzvUw+l1aIjO3f2JszP4OtftUPgiTgKW7NqN7BrZrHUVru+
fmOnv5xpreDv1n2OjlLs0d4Mne6wKnYZ2g3waNmZxpEOmoMBQlOct45wfDdSYbXm2oD5plXrStwx
5DZ/dEP9BJABw+f/L+etF+hjR7Ojmg0e3Aug2aAt4B2DOu/4HMV9+qfxful0iRdRqBN3wHMNvGJF
nCNAPOpv44FWQSlbq9VDE0ty2O8ssDYHFSEAY1x+OS6XMcdvx0129/mZBYUkKdCHdqUqRXVJFFEG
h7Lk4aVYnRWYgOnQnoxiIl0PHUgPFRxEkuzYc+cbRe6F0rxjbcIQVk2napRZbR8so5+qRXCClQmx
gxsLep9kuYtLWmwcbXm3L5WvZ+/MAiWvlOKsd4ZmBadBcTtzU9o764t1Yn+F+yo1/3nWQ58GlY0N
iVt51GRaKnOKp71UZ4ZtInXdrah5d8P0vidJ9NoElR9k83Vu/HhUG+EqEqearJ86kjljadR163TV
ErbKglguCt9kQNEQs0FfrtwMNnbWzg1UXpuxEpcOoKA/F2ho8SJioZbnwIcYUQOHWrl3kNK2XpRG
dt6jkgwZMnVLSpLAmq8o8nuS84B6C55VJSV9JFPGdFVuXxFSFIzdQwn9AutXwmuaHFTw2tG34D9j
jtJiGFEvaNEsszXgwxlrZIhWw7XjW4CRmm7ZXXKZ8dlyv0ngiQEEB1DyaPsJ0Fp9Fn5cteFiMRxU
rMHzDGfuo9HYgSmzpDkvY7RR5Jl0DPLU6C1mYXUCUukGlQZlFXlAHJsnq82kib5pqszI8Q9RQ2vM
y4/YWoLuNHf2eJVdwi/Sw0d3hIYDSsozsXGYzu24l5vlW1dD0/GnbNJotBLJM4v9iuR1DsBpmMEN
jvGuKVRgR3XGfZ2vA4Gww1YtoQc+BrPasE+0b7z6wJ+I4RnJW8qdyggCN+T3ovJ8oS0J6KBHEr3T
B4H43+zB93hSbGLfBE4bl2vseNawHNhA3ThHVPExLQPIwclPXFUPFxhvPqy+td4WVxwZtb6PbpBr
DAzbUfXjqHItDedOEJiSEvMQzIzX8Vse2Id3EogSac25zirJDQh7q7OwmSXF1fQux7ED04/wstkv
uVaLJV3QLBmvbl6XJIrDscnyxCgOeLQPTSu8yP100y9mYrF8mIm4MR526mx3oBpcNN7Vz8jwoZp5
3fZjY14XAJkB1hFY8P47gSMaqpAntMiKlS+0jicNKSK+IploS+WQ5aOTdDH9iQyvBw+PeeA1zyvs
E0IXl8KjjxVWvs5Xud+FCVWpQeORse1QnyRg/etGIS8LHsew1xeiFhKW0aMPwk7xIwkk0Z1D2yoJ
bOrNeMJ2G84NzykkxP5+7zk0Yw5HQD+Qll49gk9AyyYCejXQCbFt9p8FmPYFi7ejWQmoYvCRKubh
pMIAjeLcLoR5pBxVQbyYf0Lnewi/VELPqbVX9GG9QHeAX3PWSyxCLtksnZ1gVMxWwGr5jsRhG17E
q9ZOTrOK/7X5gvdneyZPYiAM1CLBviB+t4CMvRStoOuu3lQYX8UK5Ab9+og51USmk/9YNQ+lN/qK
PfoYEEMfLOsNcQnzZaJygGHjWntg0sEHZjKSI0fEexSZn7aP4eIgI91CNeKn8GeqhXyz6SHLPaUF
BgO9gl4xLjooPy8pz4ceZNCCV8tTbeuGqzosK+PLCk9ec4bns2VA1/8pM7WnREndu/AIa8fzU+8K
X13zWCOy1u2QV93yteWHyFOMFsv3DpxBG77NI5QLQv7W42lGj+f0if0lofqaT1MiCti4ZHFiZOxV
EY3eIb5wfOEYKs+7s8JStUvdrO+ijJipUQEMpqfmz2+6CCsDQ/tyFgL7QGk2tlLLn5Qso5Ujnxcb
Ew9LyUvVvjkhGEOBPUco8eafKt927ndWQ2NPa/fig7DV7basckDzvnkxlLSBCDA0btqY5xq4TTxY
yvpKaQcmBPd6Q8TJMuINcQoccoWfMGvCvwxnlK498p0UKSmYPcV7zfbGJTaMT+7G17n+Sz0HNsKg
rYAvXs9RNiz/twfqUTmau62S/qAKUCCKUN9q1acAStGimxS6l+4ySicXGZcWG397S4VNF3nUtkJK
mslfoLBdpEBKuws5ix+OmxgorkJP6KK03rW0kwQjGxS/jjyXKQaoIA9H0t8vWLmMHXT+Fa2fJH1k
QcKa+Ys4xCM0Z1MsSFWIjtiAefBx3yktji3EhO30yIYxHXtBnAG7tSJWoKPtNSKo3MwrqfVvAQFv
4nipO1M7nVBq1Zv1xe1dCBzTJvWyoh9NY8NrgjuryPgzeFjD+2KSyDleulSWvOopLs3XJesNwZ4R
2vXfscrKYIlNlGdMC8q5Bti1KHaabuPR0+aCKW6jvRpkLLO+943ruMjtqArCa3M2lpj8ZKy1CgYx
S8pX5JpbbdJG5p58oIMOTjy7XojE6R5BYs2jMtad4IH0cQ2Jx76b+Hgxdi5VegCM9Gwzu/mwbCWx
X1YaqJ1sbi10jORJZx/6BJFIBHDJpE8wJCk9g+xLIwHNqiz+AFP6F1HBHTWqkYmHTMWSxogmE4dl
o/JaRHYn4x7hXLpz33PV+MGjlL1wGmcGI81BB56NqQrhHGn7Tg+OVtHHYNXkpMmqkWqWXrsGt/vB
gyD+QXZZCdXkB+pml0VvciKjbGReGcm3BoZ0RHjvwoMET2W6yjUPM4CK8uzNPpu/xE9oKvyOt6Ip
KP6s7Xen0sKrEb2EZfbypy7TP5FzqdHw0OAffl4C1tIUMCgooK+px2Qgsfy/1H0z6Zk1E3oXq8u3
HtwMClsbGRmpqmLwc7IOJeC4nZUoQDAwBTJDrd0aHKvR/iuZ31Z34oVxBM4j+QakNN5UJHqWrRr1
5BCReO4mua08N8dx6u13P+15koqaNt2tF941h2m6eZt+H5oVb+/inR47rTbAcO8LaaJy0F5Mqtfx
l+fVRc8zaqXbHAGJra7HtgjPkydKPP5wOFgd0kZdUpP0ZhrjcYS40GUWdirqlr5DnP140i6PHLWu
aVQ+bvFjwn8+8fRjRgX29xaL93lkYch5Fsg4jkK4YaOEAUN8qkSbHq6dY0WRydAJRxpGLJI48voN
yy6WFssYlzkHCCihN6Irf6HGW1DV0oznsJGD2Q3KzMpcxU/BO9vakwRisdflWJYdYTu3+OIf+plL
+oXsL2s+hXjALi2AmpFB7QFGKz9VDUNDyuSxjJHGST3GhpC4oTCKrHZouaCBrKliTD4UkvFE+opb
5ifiigbx8S5aXeB8fd2z0XIM7H2BlaB2Am7rcGxDvu91MUNTovrOQu27k3KHlVuFgSCuB9i9PSCE
x+GNXvzWojk2Ds05QY/oLMwcpjWy7/ngTk+oq48JORRY4MSJPlMVwUhcLxVdNQ+8stIPLcYsvRvW
0V6mJOaJpU5l5pOdHLRDdRnVivyLBz+m+WMxQtDs6cwtm2HROA9fCJ8c7qTdZPLRE34pOxhT3cJG
BzYoHcqV7t99HJBEd3t52ctqo5e9LBTkcz88dh/Z6BaraEySlpDyuXBPiFhciUTUnNMUOMag9jAi
9bPaQmIr6pS/g5xsezI1Q1wAjUsdpmkCN0m66FWv2LCTQqM3twuPIw2+iVwDbM9+8bdidY5tlMpt
fZfKgg6e4gZgRpMTAaoV5z5CxdrxlQzA51RLC90VCLAEJtXnrFaymaZhOk+S0oFeDvPCQTbxjznc
RY9LUcUeeHmIHg5EScUdm6UEPF61PBkNisSeIV6cvRmYC+DYx54JS/AlLd3/DMlXccRZSo9Obu5/
MOly9RjpY+fLMrh3MRQGQ90vasfXIrfCog6qwFNpBZPyWZJci/nNiVm87u9nbNVHgfYI7M57JWNH
Wy36ddOwQg/7c12dr0LhQsrgSX/GqYnxkUqfuskMBUYyzadkaUNKA7gMv0+TSYTj+NuXNxodLoiI
P6vH0036sir3DJFCSJ2Qg7Mki+GjWu3bPvFcdWAsowV1Zw0NzoVB8vdVJsAF1RHmKSx6eVS4fU7j
4cKB7HWKJBTXHGZPnP5/Dbj7u95mN7PpUPPBfs3y2XpPROcoCSs1yOrjlwl39Z8aej7L84Vw9Tlj
vKcCo3tbgBobAcfABTWcj38BKzBv7erFjJyXz8uG0pCJ2LmjQkARyR43/E1Lx9wiHGRx0psOTwj5
uk+trEo+L6SSws0H7DQJFVKW54xj4p/baLaFDOJhIjc/hScw0//CeBH/cziSNsQHPqEwCDCmYv6N
Qte5xoHNG8ebSxaEWgzl6LmGvqAXESoS0iCBp3rpG5WevqS3CY9nBMb/pSpHjdA6d4BIe3ygn0QX
TzzbbTL5H8UHxS8DQFxujwseuQZXS1F3EV7KsejuKd9TgggvydocYO5Z2dcekH3M3Otl2uHDliCg
HFAe9uP3aYfMdYmOhQUU02VzejMlLwSo9ZGUEVoWe8/sVl+2BOgzgxbhm4ge6g9zUBVN2Iu/VueS
nH4zhnoltbFvujZOcv8ZiICQ5L+3dwOEzbeceyFSvgTPSXLwwEktxqmOk8g4Iippu8GhIXUI8VqZ
ZspfDHhBpex9IMTyLc1oxBOkCLsoCOHc05u9XD2p84ll5BchHa8VEJHV49S6cczHmW6wMgD2moye
LVMtPKgi2yIQrAGQrg38Ir3bfTB3xxtShbGbxlvcIS3Y3rFEX6fuCGHk1hor5eaW87cR9va4aCGj
9ehoTjZwpEqgLpqgmYQad8adNYSS2xQ91iG3GaTk/OjGWm+Lvgxr9jga4M6esFsciDoMbYW+/XBG
B5nXxsx/qGNArVZA2zhgHEeumkcfZkv30HvLMOiqafEFXqvU4DQ6tBSH4ocIQcN+oO9+Sebw8FTX
GtSVJxkCQ7497WtH1lR5Gbj+Qi5q3gjY0zE8w/GLtTWpFuNT2GnBxsyDZaKe2eaOUsvBX0lnQYN2
f+QaDNXEkv0+PWiHgZ05F0brVl1wgbEEQstIZ3+6pKvgadrrRAFpNFidTuDq3htvDclU3Vv+gAh6
PFxUtw0jhC4PFpn+1R6xxrenyFkHhOFQmEcVkSz2ptgNgP0zGc2/S6J502UfvjeYkl0ADIipJQMP
TZCjZWgUBHCrSiD9Que/bsY1w33q/SIc7Ul+X8UhLe6eLptB5Z81af0e4eCfPb/tn1/nTKB946cW
/VDC+3UlkZmDdTvnZQIAKX5QzdpqR2bPmXiINdRDXKrpKb4vk9h05NWNod9ssyZcPnnMMsWEGTGN
E7J9jLDjmsV7xMQ+dLf6qTMLOL2JfwnXPWEMWLCgb/oI0CUiu974XXgz5DX9e1KWsnu6v4Huowuu
UlrwagV7MfcusIagZqWNw2mC4ZTADHhei/eI10tWGXYNXNEFz3LloJqmgfcaHcD8RtFBwIufcNVX
Wl+DKQIjjJA9/XE/4qVV9l19ZucPLSG/lOjZH5O/DPsddJY6y7CvqcGFc9tGEgY7qb5EunZfegc5
0Jvsig9CD9I4UyRhBYwSkg6O8bpv+BlkC/WdUi5xAetIf7cybiX8QnV0vHzeInLoSNIGcvRxYyPn
ZRvPS2m0YnCPzdupFSIZ2D4pwoAc937tg/vlTqsgNR9K08Z43YGO2i7yFdViYnyI/L5dyAbEenYv
DY/oTd/eckANMtwHYa/yPPKnK5UW5LmPTYMC4DEkKya+jImze50duNcrJzxhDUB5gqIvaWRac8Nd
3VkFbeymctKwDNcSbCcL37zZlCbfQJIZCyutMSCP8jfpTnps9uaHJhGVIGWLx8gM2ikj07TlaCU6
S4hSrnIVjsieuclxCQimSevMIwRPNKEyMsWdeYdBdeztP+nJVEwrmmldedz1obUjRTJikTvk7t6U
A42Ix3JeF0nUKJ8ifOHCUOFlAwaDiIvbrfSqy1grqNTHgCb3sgLLmfLOrjlsHiyYJulkdL+hos/0
I72yI4aZfBmjbuO0O4Ql2K6h2KTRZr2NwYQLCAvD4uZ84ZFddJRY5KKCl7TvU8PC2Qh+oNN2Om0k
m8Ngv8OxNxNMUSoZ2S1LP5r2Vc2/dqMIGesUxP84Nxr+XTakVBc2rfFruv6AX6m1etL8SH1ix1K9
cFZRwq3gA82xLGfjmv+2mFYo0V+L+iHh4DnBD5uVnV8c3G9uke5w7F7Ir6ep8T28s1yskgkHlnBf
tLh8Vg6B6UACer/y5Amv/7da+wiLDAqipQOxmJpvxYn42YtqBgdK43v1zugolQFwBLVLPsnIu9MZ
JEDNQOMrGXasEWQeQ4z+hQw+RO1s0M4BNkwElQW1NZhoa3+DQnMm4RGxRA9fbdd/qts+/P4lFsMq
a6wAouDiKhGhXtYWq1sK5ZKOwAejcjtEZo9iH4vtNBD/SwiWhCGFZSIE0rUO0tn75FMlgD3zFmgk
AqEyA45681Gpz26P4WRf6zHKz6zckbQtzNR8JYsljMo+VgCQ325Yt6ucjp3HfbFUVk/cMx5Bbx1g
Y1DrAKkYOxG3n220mYAEyMN/4u/PeA10BYuRhcG5KnbGAUwEi1F1IOrsJiIr3gEqgXq9yLeaVs0p
S5T+w7CJ5YoE24mbEPhiZA5la9bXFvpvSXrAF0zEWwxr4i8HGHPEznc+3MUe3nMURXWD0T5Ahdft
T7j+oc6J73F/iUPJyFRXoINJh69z7I5TVOBYK9ejHH31kDlv84TZW+hx6tx9GrS6d0jW9lyLbkdC
zyvi2zfDtJDaNK3SPd3+wuMNF3afY3EDjpmhtOBeZebqETrJkBrbW6G1uIXjf1vmdvcnwuN6j7ds
NQjeBq3GoAqvUbkAooGxalv4Z6+oB8/7NpCCvDq6YPpTO3+ELMJGr8peQZcAAyRrKMfI0yMGTUCR
Q0CqFsAPnT2t7rPVTmVIR6kgax141uGGXNkRkWYyd5B5RKKr606CY6RO6rQckgDD27sBsslMINWM
iYAjX+UjeLynPX9Ws2WCVooSucCYoNGKn0TZqpjPkctOxh8PFd/yqCgW2yA9EKtvGyo7YGFsRhxf
C4V8yjH0GEC91NSKRAaT5n9Xq8bNgJJmzCjs3Upqe6LCG7xB8glu1ZCwE0m7/8vKiYtcZoMF5p3X
dr/cHVoVh9xxOODnW3/+ZgQu+z1xEpCwo5do2yNwvVqq9+gZNxFLN91gmQn2FLC+RJnGJbnGx9WG
6jTjtgAmtTEoQqgOzLCwJZHTzJzhhUIIlWf5Dm6OIvOEI2wRLl0/wQjJgfMZGTPHdEpjpnSBl5gW
0Df7gF4pbvdbJbz1gPgv83FXJ03bk8S7ZUDfRVOpxt4IrswRVloBIZAoZYi4070T0gmtgMPWd2fy
/wCSJjWwk7WzeS1MjoN+k+NIB+yQYSgILF8tkjv4p3TLCJC5XoTG7HttVu5NoQbgRg5BU5gi7Ylb
s/b3QeeWjGxi7CHnz0xTaVvJVXVRYd1tUFQajMynYMXdKDPbn6/Hv00K4e0Kh9Jy73jyxE72hiIj
03j4Q7d6aobfbdmlOeKiOsALbPsgtHvgmnxbfZ5Wo9xSzTU8X5fD6VoLmjh0r/c7ik7RUW6w21Oo
sgqBkvauZKXeVZ4VQ4MmO7uivG+XCuMsgeUUM54VnZ5aSdeioGwZ5nagZv4bxWo/DbmJk9RIzsLG
Yl9T3QMCjlVdCbWqmJyg1WUEyf/23c7pLRU4DVAkHtpHsmmKyNPz/DDkw528K8jJVtf0erBSLAQf
phU7UkAABI3LjX4vAh0EHOGV1iHAXYjl/xP6nS3zmN257YabB+jy5WcgR6zI79tHy8S9NqAGYwN6
AfCTSaw2hhBCLDQy95tMugUgGSk37AhEiDrOn7xPDZXwAGUi2cXHFGHiykOhDJwwx/W4q9jweOiw
HGriWLhYs17n9GFnYn0iAhbQ7TP2Cpjogx4lA+D33mJ+Id6ZFnwtWjGssatlkzryzq64QZCV+4KT
/GluCB81tKcIB4xwE9VGUNx+74YQdQMfIxANcEs8qf4bBRLjFvGrQec16AzqqJHAaHM9pebHFtgA
U0U4ij0hlDdkoQ5F8NioFCo7QjjBV+DhY83Kl19p5Tj6oijBXj4rTPjNlHuJG91dp7rOfc0aW07U
JszH8o5yr56QaI/uy1jIQAFtjR9KVuZMfBPK0I4NO9rkAnxU/9YgrRzP70MEIUrxLDacSI7obxFE
LE55QMWkzeY0XgUDvxQDvBOeHjWjDgxjD5LhPbSpiwAG5zHwq89bHAzoHJwq4r2UQi2hsfM+uJBk
Pn53ecAEeCAOQKoDta/uBtivIEw6OT2mtm3LxA51FTwMtJBB3IOmtb6XI5fKrcecO3067oz03I17
dN7Jcxc1Iakd3fhbXAbhutCOnswzaL8dWaC4g/fO2+Y073BWN/+ZvXM9VzRWsL//nMdgnsTmBJcp
1Zk9wkTHE4YB9ti9tUWdCD/P4+1/fwugQBRgTJNSh/i4gda9DPE7PgPwtH1GemPZJqY3rjQpV1EG
7dXT9ToFh0vXK/TeWaM6OjrCEiYoUXVCT9tm5rqkYYJTCSg9rv5rMwexYiicSN9Fjfhza8rf3N9L
xj1/aPNLZoGdlwOrqmKSPSPb13QB77CXajM3TYloRFhMoxM80XfV8oSQP53JYjGYnJkAgGv/JW5H
jqjqwQM3gbD5DGKFe4FKR/+2LlGSeb7cHLeiUX1fZ2L3Mxzv2/gjVEcm2wIpbC6AmDQ0zrGt6INq
v53Lt9v0fTeLeohMBeb0vTfRurm/NqFURgQ2mJvG3GHwXHmHvchy2yc8wG7MW2U7DuJ7S6Z/BlVu
kp41ajAShAHnZKZQiYAoiQBASBf3qNx3tDJ0b6MkqusE2V3sAu4koo16l4oRrRe6pC9kDWGdboFu
PPIS37mNQ3bTncPTV9ViCtLgjLjKa7HUqiDVHmjvGHTZN5clY27bnHm74DjyJjJnkC+CQJuT7Z7F
rI5f6yzfsXTmNZ6DerurBQqg0LodutLLFqCn3EvuV8DdV5mquMlp47fcllVaYyubl+chZe7DPP99
SB1llVOLfBE9vJHG3j0zt+zmbFA6y9jQceljm7+p25MeEUy0FU3d1HW3oki8PNgMc3Vhab9L6Bnc
Y7ekf2Z9dvbc83c5m1nApnqTJFKOm6FkJ0Gc/24VJuccfiZtr20pN/Oj8ArPTspfI6QpQGpvrNC0
HCuYxy8HsSMRn1CJtL6da2CZH8bm7AgMKcTrfyM/gcW6bhJijSYN5A6S8cjM77v5PMsYXljSVyAg
nktRfWHgW6B3OZ3vb8ItNm10ga2rgyDUAGCIqPkZQfefUnWD5lS9A+beVqJrb7tPrgs/nApqkSNu
eXa2KREcEj60LBOlZbNBItNNNYUhmL273gLHe51l3cV3sdPw1mDUH+QsoLikwp1pFG3pZdvvzF4k
NlutrItecXH6hqYUlnex3jxrFl3HPw6fLRmm8+B+OQwOUPf7in3kjh7B+KA9Wtn7jz9n1CiYjWFL
A1ICeNcnZK1YT7GDxInnKlRSZcP5nt3dvY8h27sa1max+/z0Md6VbzXfMrAXPytvGqDvtwNEavTC
KOYs7C+JQtcxIFkfhylgHv+9xCNyk8Ksc5QuzVvbNhphre3c4KyEQjbRNyCs3ZMM3i6y7mDtbtqi
eAT2Z8J+QGdeHD8ugK8rhjQqVFmnlXipUVPOhy0VZioOYXcyc7v7jsA5MNVvC3nGjWqRAa9XyLG8
uIqMi2abIIdyL6ASZ30QwIP8ZBAfC6t11ghhvwPquIZRZqJA3iCa1fJVHCu/Bk0iw+dOL2lPTsBt
nPQhTMj0UMLUsJS7KJxlHZ8GyiO52Y4AuSU1M+vMUumXLhoTOoBwS4bjimgkP3++CibFV71CJX5J
d5CPqiuq1+kN1zfhMMwWO1mIi7i0qjH9atbUtGRUdn+ri+yAgwL6Q/4DQZUzklzmMHgYt8ohqGSv
z8WEHm2Hc3jVgeK8w4TTUXboBhmddRrkbnR6O9OOxpDxQIK9GjbM7EoLdxCWd0FVeBu8epB9Fx5I
+l2v7+IY9/t+lk1IfGglRnJ97bnBJkbjGDMOi+97ZBRoYAmpamKX1L5jqlWpYh0q2GbD0hENPAE1
GUWsvf4J4ZVLckwyoj9/wGHT4GCOcBvXctFXUXroIyYhFL3Me5erG3flVUilt8vCzpVZurb+hSZW
ZI9oAlmTrogvhiD9D+ugqlUcAitLA62WuZ5e5Nh8r/jaEGHw0ll/QUJNjRzla2OtgqO9YtkgD3Wm
r06kLCLzkIKEmVNzp1Wen+1t9Y5xdigbe4EiA0MNJBfdFMqgpPzaDR79NxtW7jYe00YpTrFDs8Ma
Fn02BWerr1+0A/MGkpgIcZLVfI9PdKYWD3WpOOzFsR7HJCJHfTBD8ninLgIVvZRdemZ65xdXnXz6
VtxEwfw4BRgs4DjznYW8hDLWBAeG9YBK3RVaqf+Z7MV5X6RQgzfenIYvJZGHlfgXTogRAS4qAjsU
5N1ymbXTurkWw99pbqd8mGb+7Uqua5/DhJAhcDiCnRfNJtjtMytFhJ0j3Eyr/vT1oygXzPEDqK7j
IJgkZG86pOfeDksigb6mC3t1/Oa6YWTBS8I53ayhnuq42N4ddNWx3JGaCZDszkDT0pruj+/FDh+4
uu2MnzIZtJqlLAPRlnWA+xP8rD+W0PV/zrtiWJqqXMuwst8CM8A021fXhLopdbYpa9WEUjBdoQlW
LvJPDvdUBFuc8wRc7134B5+2ubds93LlU0oR2mcRPe1Ljdd5AVAtlMvO9F63NWdBBaLfY7ba31t+
3G3w//sNXIklenEuMhF0RgB1iAJWLr0OOHv6/Q8+vctSw27psjH8f6+ZnNLg5qgPm0eZpNQaqXa8
b2RAxzxw2So/7BWSykfep33t82e40IzqBgRXxdkA+MFYnslYIUDyiJP4FN04I7eFFe3/NrDSsYy7
aEy5O3OQ6CHznHY+R6g8zyVB36e0FfSFoFIKGTxLdzFL+wY/TTXQX/7H0FGHASdLllOlMVFxyMbs
YjuRQS5L5ddoRK9rSrzTCy2c9np2zxpweGJUV7/G2EemC5/MbrnEmi/tQj6FaUHQDwRkloTeT1Ti
+RB8+cTQb+mK9APJLKbj0Hv5CAPLtsLsftFZAuBJcyyiOEGDUQfbrlfOb8tG5uhrHSlgWLqLgndp
S8UiXAkf4blSOY/lvAzgecISPpsloOzBA05VJ7bIoM8t4sUYNGopxxGXYUfN7PbaDWPrdLlGILFU
xkm6s1hqdICEcMsVkEUfM+kTAksZ888Xpgihs4k8p5+RYX9Fb0Wlkkl1rcZYMv6J3dJsjsoE+ZhT
zFumec8+CAJDNXvVqFPWVZIqcMwqs4viIvuA4VJnNpwzu+Gdcvz6Qo5krO37l0I/2db3O5S5a0bi
JDOZAwRSMdWZ/a/EzPpmrzg5EOeRDEoznv3DOIL6bNMcY0KU3gD6ALjn4kK2Wx5ilMKs57ojVy6u
5wSc+oB2T/p0XbcfU+qlbJfFizref42ZUl+xm+j4S1J++H/YnWEbZ+605N278BEKpMXyzqFGCw1G
BQvvfg3ICY/5dpewdTK3hGC/WJXzK7EjoYo4HJIlKi0GG4Era1kVkz2w4Q75Tzw6TH/jon+mTdoe
lbL8YQeEEfFgJ/B1H6m5ktLQl3CEZf9MsxjW09skglOAsv5pFWt83h5VhcLKiLrkMwarDfVRfkZA
syZr3VAoASjAJYkVAbdj+mZs0QjwUdNGU3RyoeskJjrDEqm8DvFuco/+6bzhBtjmaTFnq20TewFM
6l013jNBgzsm97GQOP8uSEbCpoiJg8H4BGgxRelv2uqgTAgiRxz1OZoNEdAStAjEdHkfoQ4NO4Fo
Yjd7L1m4qNvMzwU/gTBEvpNxVV9e43dTmtXDSIjPiU7hl0ZX9BpulEqPeO9Y06boylZmmBvFpB/t
QkgOAL/Ip//N9k0pAoO6X3EC14CnKHrglccjCg33iHZIUOAtupFOogwpL+T5vJ8StJAKQ4zXjMsz
1dAP8DWM2Zdo0G1MVvaCuZ78hc4gfAenA5azyca3dh6fUww86kWwfaOPtT8sTFKUAB2y7b5SKsqV
lh4O8ga4QxwXH5NCeLHJiLdvfDo3INbWivPiCTpUxUrqcDQVpHYxH+tILZIPgLauKx6lfb3DIO1j
aXUna4LOBWRCF0NDBAFEwSGJld88wRhGpImrwvhLF/hEtrj3JyEj/c5UsPL+2frTikCbBkMz2GkX
6Jxy8w/QIctB0Nd2vtEPRUECqHVwfLBNUUdnUIEaq+XBgaN9vLLiUFt7hW7u90s74a1gtv1Ch/0s
sdvqkfjVcXw3TM/QYdy6r/TSgGgEVNvQXsN7PnQBENd1g4TsdHGij2tTgvvjzuZA6U4uOzk9h5pG
HFix/iyhGlFYzm9k68YIN5nPdukl5ih3OtAr0wlzgIhviGZiBk105srk923AjWg6cPV7iHzGVv3x
IDqXC+85+IymAS9GHhvgjYYSXQBDxvAi4UT8j+WTrlDBCACTbM0CuVUCPbwPMFFWoRjduo/OSjNn
D81Jznzb8CQ+/35qUD3JwIHUgYuSYOjP2I88dOh+0M2BQuQs2uMsP4vlvHPCejLry3rOPqBfVfSe
AkBtuNipP+ekcKh7J5acafyZQY5z9zGhhI8bDKRFtGFjTf431am6cphtfU8caxGZU/mEoS/yARsb
FM3dyvVbfRpB6l1xGmB/1gpmXZ2oc0KXyBk5i+YMAFg2buZ185u0lwPuM//drvlNgSHw9QQfzGZA
4KivDia4SkivPanQmnE65bHd6BqSMLZMp+bS5ogjySaTIb9raDq2bzO5mcUpKpskFolQlYlTqDNS
C9k9cNvhIBX5ktVBTyn7gFk2X1TRSrEfgu5wbpnySrrGifVP8qfqWrNTuKyhDK6U37lpIEa3qvFk
lo3D39m3WI1wDRtm7n6iPRVQobm+SyAPSm2fyeohHmE6a50UFbDj9LkLBW/XgRuf37BdMnSKH0Md
UI0TdPrxC4KNuM67aHrG0WLVGeTVUuy7yaFxT56xvGtIqNFgXh15WtHKslKCUkQx1K5JBiY7zP9Z
/JxtUCeLC4M6NPS6Wat19WdpdYzbHttl1PtjNXleb019oYoXGOyMTPslzoANjpUGvRekKpi5kcoj
RtMjEKZspp1sb4bPqvsRbrE4k4luYhZHP0FHhAgSy+p/xrSzqxHTrfs6vdgViDcn6pgx0tHIY0js
jlSaxi6zDgv+9U0+VwKkxAWlAbwhLrgUAzDByeSD9fijzHuaeNXkCsU0TBQugMKoyoK+hLh1IviB
+cQx7gvFzaciTNRQW0jRZda6Ul1sORWTN9jtFHjHOzQydqDZxm+CJr1rCGbY8NTDlaNvYVPuKuul
6hC0ItItuycp/kcOvJXoW4X+7ex9Yi5xijS2qqsl0dLzTlbn7jd+n8lUeNNGsX2QT5/HHBH+3Nmv
E7ERFnk7IRbnN2hTT69+8FSRODTkr0oQ7yOtQ0Pcmf8BCKNg5DLUNx2kP6HKE0AHiWf85EjzxT0d
t2IZv403eb9ZPVFw9EKXpo3WrSakQAXj7pf9IcJ2HvtGJbIxOn2CE40pnIOHr3XVZ5EMHvFBRMxo
cOQgtWTEE3dFDmbaP/rXtGoTv5Q7Mv6AGK17oRYgVNmTR3YC6I1hZI+7TFovFAnlGPRaWqIVbtdr
eNFKLB/fgJ58MMrGFsSa2GlYWnk3Uz5dOHl5s99kwsypdoTEqH5yhM3uo7A4sVU8h3wqtiBjYDPj
qMVuGBkF8U6MF6eAe0KlLy6cJqLOBVgU0sLKoFIuFF1TXPP4rCSWFrA/aLcgX95X/wfE8pH25xHa
Ug2BxuThNU0ZBFRbzLmcPSV4SU9gQMFGsJelbGpl7+jvBxy1CWX8dBOvEa6R9DWv3sGYprRUU2l+
EqsebkzBayjrlEAWwaXASPxiDrpgCHGp11kY8kB/Y35sOHK8MlHrRBg1t3c9Td3SNNLBI2ICPWZx
51E+Y5+nnWHqYBCXnYYE1rZNOAuWCZPW5T5y+G9RA1dng074i7vMK2yGczJS8tS/0VFLYTDpM/8/
9aJWiBZ4MJdwKPMaXPl/y3YM2NdRncsRDfHKsYgDzj6f4gMqBNMbnVbEKr9X4NUc/3XqB2nfGH7j
oRMzjyxcKoFqdtdDL0Si6cV9gaIb0oMdzboFflImh4zzyT7fAo19nEl1zGz263ZFDaiBum0lmKnZ
1JoPLQ8qnrQduKwksgNGqvXUPC/s3f/leDSB4AOpxv2hWNB1SMzK8eErNgwrbPXTPoaG2C7cGHJh
xc14gSXRTFM1b5VvwSqC6IY6l1GLvGQ/m1ChboH0nQjBvi4K2cJEg60UdSO6v/xGk4QmV7mOHdpm
0Lr8M4eSmLqHuEPDyliB1i5gVavaWzE9x2TIFK1bZTqADIpMUbDA/0v2nDRPZT3ld/e/8ewPzx8X
6knE/uIBjFUElQRPBuWo73AlO1F1edASn6uG762zpgUlB6YXLpZsz3cGJxveKnMYATz0QyLSYTJc
rd8XYWSfAIZRqRXpkbjmMOrvOCDtIqS7ce5YSDcJiFX6ZM9B4bG6eSOCQCJA7znXaaOCryABakwt
JD6Kfl9TSpbsZNkrs3t9F/WawXhH6KKW72ez+FJFpB3Vmigf9Tn29JZeqH/7y78mb26BUvVY/UOE
4WhtL7N3Dhlla4TetzQ2PkoTKN6sYh4gLHPXPjtoRQ+/9fVucmp/UGUQ6Yy1SXz0KQv/mPc1mW/U
agFm3D4bP/NNP4xB+GrP6T1lqp9aFDNB/sQZVmLXFW6XvdRnmsmLBqi1d4Jev8MwA7jlU4P/5aMh
9PR8CBkAnxvBicqYBrcYJkg1D4Afwly/xK/YjtxjaQS8ladqi2cQpuuQPsNjIdRR3Ni32FdJVKI9
FuGLin+UJ2vBMBZ7Oosc328GC49xK1pfQSWsKjQpTkDk+epy9CV5T96FQlFMn3DxhOqQCop+30Cb
9A5Kad1FPfuAPJIpSpdgbygwOtLdY+J/NZzQB6RP+7nAZDqM7vgjjU+qBX3cuxUdx7klD3TLcMMP
e+NCcfdlNeBOtefahhqj51Ov33/Ka4O0VdKel/NcLOxagox7ozTMzlIDmBPfD5i/K478AOOptNLM
q41HbuCJE5Uyv5bnN5f88N9POyvUE9z+ChMrjP2v17FBYNr5rzXjjSS4FN6m/UE0p/OktgGJZ9Il
rZOHwYl2p4Ag9KZFdPL1HzFouSY5fkvtaE+FJoJe80/1ka2i7IR0hz7sbdwyaKObl6j8guPDpPLD
yufsTEez3nFNqXQaFyUTAdUqgheqS9BYMHOnHkCP9bRWVoD9k+36gEkHsF16TOJ4IpMiIJE/AKMm
FyjUc2lgPh4kReOv57/n3WhUECKluPwNyl4HqS5q8r1LVLAR8iTQ2ZSPdWepsQ1UN1QzdcMvlSJm
ZYIb/8mEfv6QWKqxRcZvb5wRwXdK26mWi7eAiurL/4CM35VMdG9EgVX2Cjq30Vh/Aw+XdD3SuCvM
cppqkjtM+kLFGVXenVAZK+GMBcfinWWhpploG1HhxFbsecWl86Bum0fv78ZTlfiX2VMKBFt8j7K6
IHiZOgfAUTtvjq2tJ33OLDetlIHjyy82dWyRExlu4OwTNQFJ+PQswb2s7vvT9tt60A1okqB9wkjD
oo60XVY9TxIgDBwyvC6TAe/N8WDeor2MmfjaqqOz9G0Ii23GlkHXC8/JQDAthaAbJBcPXIZ1BYYa
f1ivxAw+rMaaRWjP6qSqD0K/jUVpuQaOkRW+lVfr1idqHaRyXLJrI8B+DBlbRQnBT5TEZpRelduv
UVmyCoSPEqO5+8vEEM4J6inQ4+u9fd6TIl9dJbYWPLc0SbJ2z5PeAjyrvGyZVHiGpDr2J/47N0EY
2BGg2hqUGr/ALgytjJmULPF3D+zXFlQJis2rB5PcJ4ZLEOA9yC16cWqeqCU3gHTaNY1rV7JL2Sjp
VlvgFT+YsVvTWR7rdd1XeaWAxIdhys9UienCUrsXwnpwSLAUofuM4Xw9jBPvJSXhmzB2a0bLnylI
9OGhJ1X4yqENC9s1BUxufOWin9G1v7FnOO3K9u1slVhlIEBIwHpA54RnTrJDR7EEucjtyY+zTSu1
0061PDT59zymat/bJ+8hZ8uv9lVBBCE7Skt/VPjM6i74wuS5YAsh9QfTri0GbBPNvt1ihfCbG2xC
h2+UokCCgIBQekvEKsMkSnUyRAdlaCLo8CPrXUNKnK1VR+evbpi5RjtOZtwluK1pDXjFTAAwEKYN
8a8alKbGDbruc4zBJ0GJzo3vJ0M7rxgMw/uyORa++awtIDz4UE5dlll4sbS0fcAW3kjQlOddvXec
W0QQevG52mAyEMA2uJ3xi2CKj9lKkZ6/CKnPD0eRYh1pmyWf7+AUZXZ+N1XcwaQepOZBIsPJwPAW
ziadbIWHDNeVWOlOhjRMdGsJLpUmS7zwm5SSpy0KYpekrmPpLQD8JcodmeWYbDySv2IrCbpCe/ji
d5bFpRG9BRxITAfv8YQMv6/MSmiVi6c/myvi9CN0PV18DMXmhCzOm/I7DhUS3Bix0Cre2fcPyL1h
77k1ECh4kbi4Mf6XqHNCA7QICpuaCUcSLEySbNiovdKVh8cS30TlkJKHIc0000gs7PRLdLNYsR0A
uJFH8Q1/ZYUmquWrfnTYpA8wZ855y/gf8u69fO6d7e/StKVWdbcbPZI8jrKSr72KitNiTJkpQRS9
jxSa663p7a4gTE2sNbxofa2nfGhtVU1cWRrivD1g1YlarOcROwthF7QhJdhuQXcQlAxSR6sQi1GW
q5mSzZ+m0D3aCjWVv3Qy3XkYmiyOTapGDTPuehnRYJNmFfIzGp/xvfGwxkT2So+/sAJOijq/oqg8
s1o+BQzowsgVJ1ZnABoVM6OLkrDmUhcxfPhXj/iuKfNpcfRiAC1IVgzy95BVT9BPlYiT0HeszpoU
t4Tk4RmMP8nE6Xg1CXSdxSP94VOrYBLxXdQNSj7z2P9+RObFwl8BJzrtt+ToAIqC/beb1J3QN3tB
Bw+NH+4oo4zTTS8qyRdC+8iALpblZuN8O0l0lTHGWWSZTknKDfDhxBW/hEHUmHNHD9shplyhB2dH
o28mdFt191e0BG6XpnPMq0bQkUCw5MgObzHpIdvPTlHGE0BPQDLx0evYKWAv9BaVopu/2jEPaQEo
nUROXySRpGhoUHrHak764ltiYX5kl9PidSC3SvqRCCdUrt8mzyMsKenGwt5Xkod10mVTtePr4PN2
D0zqzC3AsVLuXaGccOtsig4GRiIy1q3mTxd9v9ZVzcgoC3XUDjx158P1ZzsRd/ZEeNvxoBQLOMP2
DAtOpJB9ukCggm3XEt3B8lF45fpesmWJPV6KoXiSND9FU0Vxr1NuN8N8i5lKN7OfPMTlW8mZ2T+H
yKk51O00/n34PrAM79z6hsdFmwsgbu0hhFN0VOH/hDUfA5ovpuP6s3afPGROW6SM0IZ0fovJSt89
r+xZGSRU6uOMcxYGcpypXmBuuzObUuyPWxo5+1gKroKlK66P7wPNDNEdbrxx6GJ1R1lGDNEtLiki
nYWTXqi98EAMHwwTOo8PxBxc6QilvXaBH43y4brfZNFJGVb6+Grq45GyVSjTxR2eJ+Ah4gP3un2C
fD+uWN095fBa4M3aaVai3YlJu3Ut/ZOlOfoAIseZBvzL1wuWztaM+b9qqkCzYrZzREOI+qFSMXcr
DXYsIc73b+SwB3qMEj4yQ2j4hg20IC6BvZ7403j2yKvnR1+g/Mqd9mTs4+ExLdYbAekDx+IfMMeO
WhJuu77c3Z2pm2/+ACYyBWQmX6tAdEPnsuFrGRcLg3XZXA2dswy6REE9YwxhcGS6gNGtLcru4JNf
bdvz7FmhumVKcZT1D+O+vtlUMGi9qUt45rjd0DkgesJuo4dZjjxNT+mxe68Lxu/GkMN9dYfeOp7P
LQnX9whdLM0zGv7tFu1OpO3kFAp5HQlSrtDzmZap2hNH+FEiSlBc8CqYVk+GUD9q5lrDDGeGUEHV
rGXn+rFpe4g5+EHtberArbMkZ+ET7dWNM4J9/La30ihnWC/OLiWF8CK60ZfyQZeC0EJd6/nVUge2
mWsH8Ou+29XEhQdQhQIs9p29bZsuADQL3aBGcwTHreVL4OT80FlqYtCxW0vCG7Y0zL9+XtZX6vDe
pu0Sk9+EEfmUsSm27DRI/bfW8w5Wr/CpplXBHAeO8ttY1SbWXK5Syo1FL1f4byegUoJxAIVuxkWJ
TE+F3yV4H+WqwFdCmuR36DJpt5FhvYmBA23EOknJxqM2LusX++S3pZ8fskIQ1pp48mJVE0kkLFK/
WB/wEMObeVXjmhFISSBf2aReMPQlaZCZ2TB+Tu4WT86/xFjAHsDhPcXGoybJiZ9qd2ZnsD7gEZi8
OOhBq6gdWI0kl5pVl15SC3+JUiU4hL6aZhJKHH7aPQva6aTb0GMi3j33Bvt3aSO1kv+zDpqqmWJW
NKc18ghKGG1g/4PC22/MS9Yq5KaNxJ99CNniC0AkUricnTF5sEHiv4mYYF37tiqZXffeE5LiMpAV
AQ6C4blVZ2/xl4PwY54wdV1YvSN6j5VPEz0DGkkcyUt4ADnJuENv62gsK7THfNdBBIsZKKFfFrXl
YD6LWIJBzOaGf9d5vfxY7lVdJVkd3sPcChuDWQvOTGfWtd2BDXp2QQnzkw0ypmlep3Aobe4daBTb
5u3xeohYux948Q5fuWexK/VRjK6E7rFotCixLVBsdY7Gtf3dfm+BNaTd21MPGkRymHr3blcM8XEl
GYZmiH3bRCl247frEfEYE7WkiA40lqHvwYr1K62UVQ9uJzps9XjdZrCfVIrPk3NGpwLAZVtlNlM7
APdj/jJJtpJA
`protect end_protected
