--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
HSTrKuZbkkLTVScIHE2JkHqaMUj7WIekaBxU1hikDFBGa5B55pvnMrYeMEFHLVBWzgiTFedB2/kR
eJqA+dXJSfLCBPhO7HAJgw4HDJKN1+goWXG1BeRI7232mp0taXmIU1aOGaDWheP6JPRI9N35MeKR
ytXTuEJ5rwDDjq+bI0Cd4S1jh9teoRQoEFXa+ptpLjHVzZjW2rR7vodVq537NdoxOLxx3C6KzGNG
VJIaYKwatVlOlyTdHvcGlw213f/Ab/2Q7mT72amFN3KbNlU9jIMgvFkke+75UFm5s25NP+NAHCL/
fXKTPUNbdyBhBZiibd7RM1b7QxWXUxfSYsuREg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="9KaKJhHYmmOEPFoPXCEqgwZteEiwWy290Q9jd7FTUTw="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
Segyk/ytHDhP0wuzfPfM71ExkvSZJ2aNe+jC0GhTdcKbrr+WNbYxmY4DAOHbvLIinqIZhOAhjVS9
9AgiNUaqgMZ50nWUK/v8vC1A9nWnceK21Sb66bk6Ar4zcLSTbnyynj+viFUhuYyZIUVRo0ifbL6Y
hA0DhIB1yVmrIbAp/EaXZpqoeQ1VyDOCtfEZFgQdFhi+PjzC/+fmihQ1JhYrOqqcH925hHW+NOT1
pPTz7+9qermvZbDdfu3AvRO/iBqBjqPEmxfje0Q6bXOzuCOzb3Fwsnp1YCVnaA7gZLTjRdeipqBr
qf7b2nZn9J0KE1fKEOWEZNV+MAdrWiZSv8UNTA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Cgbl4ACHTNUfeIedrO2Kedxwhs7O0X8BQRESxKunMi0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20528)
`protect data_block
WQaYChxomx+KdlrtMbfwhFWqrRzyt0ONjTJfjFm5fzQmXLyHnEuFTO2J37A6figU7LfjptDgWH+P
WNhKHGVVmjYqOWzJHVSACab74+ZX00sj+CNr/S2RrKcxCW2I2v/2HYzqRzX0Xqnxiem5FFEeo1Pa
9OyrfCDE79lO7BFuyB7LihSA4bvGyPdI2n04WjjbnV/GhCuLeOh2OIZmbcV08oI6NEZ7qEg3U1CZ
m+mvLuIO8dF6jPk7d9JjfHTFgPzv4qpibDZVXMec1vrCsjep6QXhFafCf2HB7dxanYO47QAoqkDr
D2Z5iO+yrp/nPDNlYgs2RBA7op42zaFQmGrEvtTYaopuN2KoRaC21B4ILX+fKjFltVWdvD+2Sg7O
QQ4xC8NVdiBATl9d5DsgI4KfXnBAGKMVCr6Z0+CpzwZ9Fh1G7RSKonpgw8vDjBfuJIovq2Ro74i1
2pF70z76NPqa+J8cJZgKAGDM4614GVZ8zcF39ehAHFcLdH9UMvXFtcRJu/bBtsukVdpl+7mdNinl
sCrpzdtyLZAyTsAsuRQ5lFVE99Zj+jVXySGPjRq0Yfx0k0htCpUx2MDFexd2eYB15fV0YUtwlG2V
lahIIZfSrDriSYGZ4NULXzH7BtVvLjZSRMR1Nb4DhnhJJAI7XnPdX2tUh2KdjyFoDDT7aQGfcjkg
BTp/HQcQWPQiclP0N7IBrsoA66UuLGsebenyPm+1hz0OQUk2TyNwt6rTWEWajpFPX6jab7dIif25
G5y5YsY+psUwET9R7FsXYofBFf32Bv1Icv4WLxFxJ7n7QEdnsbIpJdqDsNuFxQp5Y+i8Oy6hgm8a
8WoIwTZInnr6Ec3CLG3O1xB0Fxu9AuW8+/KARf5KlA1V2EHSi8jE0zIHvAKAuCbMO5RUmY8h+FSP
uexTV26M6fcM/Eyf4/Gmv+Orz9CcEQGpH1qq7IH3nslROevKzlpK2sbLsIOyrHN0ELwZx0oVL5Zx
+NPnUCRDPoCYoPYtJBLW7N97cfnx+h7Ik7Uq/iYPs+3xxY5q60wWrsG9IZH24TKFgbCMgLDhfLuw
51kf5sX2K0uW1SnByvUXRGNDqgeSeg6+qif0K5X74D9mgKa89iXBwVnBvhexEfFHV2IzrMYdX0oM
5SqciMulZPs4pPpSKCCyeFAO76xMLDc3991OVZdFciKxk77MGFuvhOIS+pISOD+B7Rty+f+0+PEA
67JRinKzL7dnhbIOW2YPWdj5I3cOayYShnI6l3Fk+BkgO+mZcGcxDUN/Q56/+84IF62/JXEMv8uN
gw4YUPXK2AnWdV6n4xtSL1UwmCN0d/nlQocJaKpowh43Uu+NF0cz0D1yhHvTjGkCsfZYyrhwLePU
Fx3joruCVk7bhurqznAdGHHU5DQet25MbB6WG3RQxVWEfGX+I74hDkAUc7f+pLMhs8vojWZ7nW7d
5XtS8Jm1PPZlGJoSZAdJb/4chLsPTx9ZXKcS03gMd0f6l3n0UkHqR7cMDyJ6X+zuNJj/wEqBLvVF
B6Q1kuiqimViBq+E5qlrvpaZXj20DvwRr4qlf9IQfojzmyr6HrfopVv96rYBvfMTVcq8ETNb9IBu
ghwCK9qE4dYSSBBMW+YEw7l+OKIjFerz5Btmw0DI6OtFDhquGKT1DZSMQTFshwMWF5h8B/3obWiH
vQBVGM6GkhC7Ashx/cqzVvkakZHwg5rxnskyqgbDjndBOMYmYBcHY8Q6hXbvCfxLfojOJerXcuE5
Ptf7PdpvJVGe9OeneMMJMubWZzI7+KuALmVGVx25jyVfVIkS4dFqegBqT9X11leRGrhiqn1g6Vg+
4BzxPmdAsqJHufEETNa0bbjZcIFkxZMiiV4l03+zzRi6Cg7gGRIDAcKkAvUT2RH6MejyfjO5RDNZ
W1k8+IuKOEwY3bJTg2HqO9N1YgHSKa3agFea3IcvePSskuhE2Qa2Nw9L3GkB1nNx14T7A5n2ZZue
fl1pfq6zrJRCglfL4QGqDjYlXQDfJZu0Eaaj8eiRM7hJuUxUY5p8DX1HmfEH8slTXQet7KmeTVZf
UfD9/yNjogd72kOq/4XFVzNmFRH5ESA4+7CXqzvAgKhNCd2aAUeEKl5/2B2Dz08QjotgNAYijpeO
HA1YTRASz2RzgRBr4F15W5KlDpoFQ+j76aMDuYUQFyIeu28NuflIQK1vPwTosyWoySEtP/bNm8mC
H5earRUcMgiWB4xnJw/UjR1wwvjLhVa4YSeM4uwBMMR/FcrhRL3E1MBwkmBm6HeeAm/D1a0n1nQ6
pzG3riwd1f47+q/qTgekK0vx0RTlTl7gG0Ifmv9S4/YqKWc5cWfGJuiGLcOd+4PJ65KWq5asU8iY
Ec8JZO7VBqYeJZDcOZwCkVnFUOGaQSE/2s3LYK/7qDXq+OQ18y319kR+0SCzf+PVfkCE/TbvjFr0
zk9ImdGFGXQIRezgRQ5SeQYjEh+NaWKNtikyQjUCClz05oOqk1ZED/LYoFO8ROf00VZKg5znsplP
OnFQLnMGJpzX6jFAJiMwr/cxxWFwZEDya7WKrtfPImWpHuF9uR7R+4QJt968aAoo535w0ydruQn7
/1MYa/ypn7bPeMpFyy8K8vFCV00ZAr8slQbB1wMosO2F3q5H78dW1By/mlwl9pEs8qMXDnXTK/ed
0THGccL//pC+rUlqq9dyO+H0c4ouGNc1ntQdZCUAgRIGFGgFYCMEm60CUXJPH3RRHo0i2H4NDO9o
1CdjCz2TDJbe65bKJ2GdaIIF9kiWaoqp1ev4TdZl+x2gIn7ukVRdC6hxiK939AwaTFqFAxaKbd+T
a54nXCCpqRWXvZlBC7RA43gtJ0E/flgYe01fgA7PkYX8x8AIFeSD4rWY/cKIHaiBVMUMVQWWrqRv
v6DVuYhHJvh2bCTU+r+4HtXIr78Zi1VbX4GKZq/ZAvJbHXGzqNow27O+nXoL/u3GgtBcs12KhvUw
mf6OZDqTRJtsGNhnsjVmIK88IqvClmEq7Bnhg9eYMsGVV2dNIBwzx2ZOkU1fbvz3h2AkWSisxAIj
oEbkOVAjxXwlHHiSMtxg2BoT7Ng9ePFv3PaUhKipFTbCjnICU/oKVstQMQLPoPPpB7W2Tsm1aiZZ
F/1JOGPsNm4eMftBmZ6ivXTLNt86+XiudH6dfHR3hv43ywNGK8SeSohjZSuAOKJ4OHHncw5SGPMJ
UHuiLCzQQkeM2J0v96IYwDIZPGQIvhHIXga1DauNgCXGV6QKGmPMfffJ5LaKZlMT4DDNf6b4qvMf
lEM8TE7STp7oTBjef/RaLvRZD0cjK8tC5+VYnvQva3qynrXOSTA4yIxSOfWx2shPw1wumhJIweLQ
VSrr5VLL4qe/FwmY3iSFdLO04zXHwgCa3dGYiHaOouY9PZmmJ6oMPCWsDA3bbQqFBarhpOehgEhe
yMT7Jq3hx2WBoN5LoZfbjPVihOpJltqWCQb9QgvRd4iXSw8/KMPS0Ixp8HdHhr5fOAAv1FZi78WM
ax80jUAjjVB5EWqFZv/JXbm6GDuf9Y1Y4AfLKMlDyCZ3P3VDEXaNmNZkZp77zxyblNgKLP3VwGKC
n0xdCRqWrriOg9KhC7oIx2bPqukwh7y1KpTWbbUpPo+VYV4SzTzZKPJVVik5Ho6a0b3gfGAbaspZ
S5IQr/T6Qq2fxIhCJqT/mxhOC+05VKHkQbQoXuoeaBO9JZ7s3AwCGBAA2RJdUyDCJc6ewGUZzYcy
I4jvz3BiUTViW6NrYI5hzORVeAmfb1NM4flvtBJ+mhJztoSxT9ELr1EUHwjGkRyeArakiQECr8dK
exfkNwlYlt2SUcdCEC9Yaj//M13uAKQP4jKQ21spDpO6y4TfAyFkVU5LWsQ4OgrQeTDTaeTjSpa/
GkGEkwcGj2fKvpNbYVBmDOAbyn/sfwHc/JBvm6Fl6F4DHPhtArYAu2chFNdwUxv0DMuh/8hekh/y
wqQHy4raxNRf2lpdlGRCxQFSbm3l5z2gt1XPF0BmthF9HWTLJ2syTqTqmYPDNnCkyP7ahL8XaK78
TEX7I/WPL+mJfCYKoriBF6+8LUjo59XfGoHv2FLZ5An0oAKz/NL6Wjx2L+/GgutgPhLtIvbR9zPN
Zuf4eT0FLk8Vhu7/wW4zpwghSVT+0bC5/nvSWYdoiG7dLAY8JD2h/6TPnT3nKhjT1iftiLf4So89
hBboSuBbQfqK5nNV/4WhWOk+ZvWMmn+oVjZhI9FMI3Em46QVcf/19NyIA2Rj297XChdFnOSCjPyu
ssLYxeQFNwBj0WFw6X0Rh6Jo4KVAyIbA4pLZDcYFg42pDBnODWKk9SDZzzJpz7gQcx6pCH3/2Yt3
NHvrZYNYSGicPnkQoGA1GE1vWx634VX/gb6zLLwm+Z3giylrkaK1QZPM/2TTP677oSxwv3Ku+mzj
RuxPSgDifaZPw/nAGfVctE6eTPWfCsUXUjRd+++MRA9uC1LdtJH/3uclnZeG0Gv8qBC2r1Hksalb
BNgIirbooVtQWyaJqdWk2W50EpN2CamuTpRXqqXU8kEnEYl5HtRbmCFaGV8nbhdw8NsKdfmhiE02
aBnv4CbS6oZgCzAj2lCom1HFPOEuzgSXvEumnHGxjyqGtprlF96bkLPAVqAxTwXNWBPS2tshdHN6
7KAyke/nUxDfnvPBdyGZvQbqSo6svd5fdRIA7Kirdf9i5ghJ5MxMAlB2XMFfxyM3IhVLvf2oVMm6
fyllCVfcUHPyKs4I7dpnsx1BY/PeYmIwbGnB5lTqwo4D4/4gPzpihSBRo0Oc8lGd6fCxA2SueGuH
X1vr6r7l1NRC8CFenNqLWhI9TVyHnNrTWvvUSNga1IfsYfGI6oT82sYrmLZZAbDEAi/6A5v0Ra+f
1c1rHqstEHckYaM9fNwsvI31y7GRH1aM3p/3RqeNgwDXi3NW0/ftxk7uvXiCBVZKGZZRCASTF+Ej
dQCWpGDDhAG1C3VJRKQqyxQLYdiar87S0Rcfvaps0We2UMeaoJvUjdDmbN4zQ3DCkWuwKXogMdbK
KgfscdNzF2ImTAmffTFaS9UkHo17nUR0wN+x1QT02sVA768l0fceFdHOLv+CNYevDFomVTwJiH9G
QN9HrXKvH7pLSXZ5CMM3/iWbCjfRZUvRbvEetLBbm4rLfjHnc3zc2ZVxQ8uV5rcMPEd6NUyWIkXf
uNfK1G/RW8WcV3InJzLY9Akf/DK4ZPbZfxHFgKe+6gIx9/rNUwEuEBa5PhDMW65nNcIawuEa6btG
ckdJAh+trTLs1Tv4AA3pW8Nlc+0l6l4v/TPGUY2qu6jzEvV/OdLrwg0KyBcZp56Kaqq6naiCDEKw
wdHffD7XMRsk+NnS+VyM8XlgykJyH63FOqjMlElFR/4FWwBDzD5YCOSjnMKQGShqkskfawLzqEOv
ST73UCUDuPgWWhIBCChCTYQmCh9ZTQluMEjTIkdQS5gsH0DiAKj1Fq+R00Ev7W+KBctifBGRmzAH
r7ZeA3gNZXfL42z1LI+BNUoxK/kEL10jgt0izbL35cBQyspP9fATC+VnYX72oCMtOOgnLk5+Bkw7
bgaVwJP5wB9KD3UjjPBxVe6Rd7GFiJ0JB4z9UddCltCRpbPtp74LUuHVBMYXPuTUWYC+8HKe44yr
QroUoqCGj13wJBrv7/DyTiK7jIQnKSdAjWbkYO1r07JnPlvVbMIghr+rsmwWOwKs2QuukMp11irA
dk4AA3oaYk4BLUpMXw5mkaFzCZ7dsOb7EpxU3tCYbT9mj1Bz0HP+L1pIiViyuuip8fOCUgKN8gBa
df495y6/+3GVBMMamELjrXaMj8VpNnp5CapbxvE5oJs6CufMZmfKuI2eVVJ9kacsi2Dk7J3OaDML
XD8ixTT+7fSLom1tQT9zwDpaJw1Li+arAK/pQHmP/L67KTnWP44XNReyP43pvy/NfOx/XYK9/eC0
dx1r3UMAy7Q3o0Cu/cAgtVV0aP3E/F3sU9rP9grGhdLJaL40PC4EC0TxD9QBZQu7hhWMOti4Dno6
Z0uOFm/+M2+x+IUcNJn82cqPlun+7VYLC01bimel966nEcWyG0VEvUAtIu/UzQC0ihxEiFFxmw40
XiJ3z2fwase6l4niZ9HY+Ncgno00tpxWVWTRyk2qwbsYfcBZ6zfGknNdBYlgycmzR2kXCEsEo86H
GA1t6SNMBYH7CjG3TvuYUEfWvGFXY7sVzfOCt/ofpDdectquFg9HzZFtNwctEgILjbvvlC4kaFvm
/A6YwjM85kYPf9HOm8s80BfHgN/ooyXMsuqdHD7QocFF3cdRTXfXoK93CWF/V91A0o97olTTsyDb
2l7kwn/2jU5nWK/fte6Az6q6U/FbaPvXj3wteBPpyqxd7KBIKDPs/CBCxXs7/ajA4Xl2l+eTha+m
2uNv+ShN/4k4VCo2H35ncFqYgT9NhrwQZ8qhnbJgeSumqYX+rRfiXBR/RrOzdkGT+y6E+vTdotca
03hJl3krUQq9aSRnLxA7QtIkkXozBHdvu3bnOpfEAoCMU2gWoyDf4B3QY9wIcWtkvoBP6EDlyhpU
YeEXet4njE2aS6O/ZQQ/U07Dcm1RQ8BQoHYwns8F8D+mP7ZWT3kaVeHGtmGjzsspX7oloqdUmTBh
Qe6A0xUdZupg1cTeq8f/EA5R239zgLOzzNga7TQ0ZVoW9HQJDxICXSpuxmZ37l79Wy1SnQJafQPe
rCyI8+c98NjXSoWSry3CjDK93P1dyWVFCN8NJKutjPZc8OqgvSRJUZwtjNvP1UKwc6IasKcInoc4
NMk4Rw/pgscktX9oqbfb/3aiIwBwHZSI7hGw3g2joZ+uHWPnQToJFNWeftTPgXOFDPdGPMKl89qz
7/k3P6h07lC0zQmCI+AgKjxLaUf7f7/CKQU8wQFMNGSgIpJ5FpEuHfdHbU7wi/AKtKrxNpD7UlP4
InbbkdaKxg/Ati8YzwT89odSrLwCTHiqUXrfHqCbQ/7eORqrEfJI0l19T/5EFbMiWUKSfEW6IpCH
6OItiNIJ0iG5vFtOoVDkRhArmXRmgruopJQxstJm2SZmDeu0T2cCZGkb9GSBN8O2wqIBK/Bt+ydO
hBTXCQaTeGp2MtE6ymoGsTF7tCRwRCCAKOUWykn76nC8XJ5HpzldOyN8Qe1Lf992Zq49SjZnlYlI
1ilIScr8TUKfVDv9T2+yTHcrcEIiPYmYNWtCPOpN/EiPkFGXPzvJC1q14zVncA7yFbgGGEuikQi8
hmrzwQEdpojHZN6X3VapQCwHrdqXATcgIzoF7FsBrt0niGDYG8h67FsDeJq1itWEL+n4L0uq9KXH
gMgtRs8+YkBf29lopjCX/2ba1U/ZnNwZDgcqQ8lpnPfYk3qLTCu0TzALfAfPOTbQDGO2yy16SLK9
/DTX3FaRO+xl2KKntY81u0w+fPPasJWN1XxBl8Z3Hce94xudZJCEE+OGMyqyqnbq8DWDeJpBoViq
5Ba//ENrCnfnbmOjJ25t9HeE9gBdF0GmFBkIgwLmnf30q/V9hRh6iO0Fi7ELsm/qY7EMGLGNaseW
DmR/KZVn65zOpaX9d/kDX3VlIdsBbJHSOMPDPiWDninlFxVX6Dgee6AouFlLrT0yDdR8mXL/g0RN
KiIHkVqzEm1MDaSPUpvBdNGTUfSttSgYrD0Xk75VmlBzFIulzBRtNUSx79cqzg8TbMSMI0JkSTRI
9udLgcVJLksqHoz/9rAFW9e28m/gcBxl18VWPW+PEEvjsvzIUwn4sS5pFKXgGHeYhJjcypDCsrtU
zN/U9HOPKX/16hmSFVfADkgALDGuu04pticqKJBGM/PcftUTJEdZd5HqbXkjUfaA8QUja+dU67nS
/TIH4eHd9dqQaalrmP9dt7tiZIXzmjirNtgHSEIV7UcJoH8CUG2Cou5OgRSpL0ndkZ3MDJ2o8NHK
FPzgvu3Otux4egniMlzo3OAYnujIR0LQ92Ldv4VEEzmRstjdABBJ9OQHIuHHKR7SCHR3Sme83Nng
XaS7wS4THB9sR/NhTnvamEa+3E09UA+TK9bbyAbcvFEVcK7vK8wbYbQFNNuYJsZMO0+OJ8blmZ5k
HoKhcve3n0XHyNZCfZF1IULY73c0GE2liNFuFqu4MgdUzU85M+XgR4IW5vEamlheeoWfLSssSI+u
DTrqBW8EhWtV6+3n39ELFZr73Q5uVgDdeU0u6VHAoQ/tMzOwfAkbOPynfKEwPV4UpICzO9EGkM4b
KnaAYClY/q4CQTCIP3TKpNKa23fqotqErLR4vacx4dh7dr4fOE8ekeFsXE9HFMWmwA3YxFDnDWBJ
jsV0vBK7JugmzuWUccLOIzlytqCfYmhTb457Hy6Py7f/yCt1n2hcec9yZI/BXv8bKw8iEdPUTHgG
d6YfYAczstAA4+cRzOvnT1EFy9L4nunA2plkQpXfd2gCHjUo0Ec4jVoQ5Ihgcd00KJSge+2KDflU
eELdqt15KrwPoMBcKJ7SpiM0BLW5N6JnSK9Y4bQ5NZqUhBrQigNMeZhU7WLsKExwFRIuMkvnNHTo
fomxgissZ77dOM3EZI2lbnU1YjOmLGwi2qC9Xwo9+CO8LSGYYba45cwmYs8TFubICQ9UUuyXONK+
R9ROiYhUwkzlRBHdTqadnp9PF7xltwbtzOSl1259Wz9AV8+njBcQGOZIyeGEOoTYX5Ok0rN1KxgE
8wjh5ovdPmWy7ppxY3k/RvQfftzzY1kUoVmWp24/L9Jp4CrValc8JVhKWZcR8sWDnFUw6DGfy9+J
2SAuhbRO0cDGTgEuxTXyECcebv2D849MSD5CpgxHPwsP9vqxnoRc5occcbcvomfgiyWtBCELagxb
MHgT66hO0wRBpk/oowJ7MccSUYXZKPJMDj4vBWvjAA/T9PvHzyNn4olQLDkx+J7gnhkGq1zMKaF6
y+dh7xTXdZzhxDk2lcXarWB0229UyafWFDTn3Ff45+xeKrZmh5oWnv5VvXIpgGrQ34vcuvysYJ0x
+mB4LkRzMM0zbrxNbGUK+ikDOHusD9u7D3fz/owrRrBBoBBA/ELdVy2eAMuSNBbd/SLE8x5hmV3t
J2P6SrOPRxFttULPV4mXTN84bmweApnNuOqITKrEi7ADF2IEnVdtwg4YF0AFB90FWWa3tfDIFu1g
oOZnbYXzKc++Kpq1zd20of3sjrqWY8pBI/K82EGhi3C99w+y8iDkIb8hhts8zafES50ThpzqmNGB
f08bKgylII3URrgBP9T5jcqF/yiygvGxTX8pXTKKZreZT22YTVNesVT54EdoNAiQcWuxQ0oky0iz
57lSdO+ZANOj0Wctzg7qzbMfGSW/6rajjYXGyDpYrPBKUSVI1E65dDxay86oMG0gg+6T3hktrENI
p6reaJy3L0agzRap+i/DKZmIGYMEEXvpudq0QKL1PQdR71dFpb9CBNwWzwRwrylxRf/Wr2wRmBa9
OSKIzeUeQ5PN5pPNKbZE5C/Nfg2dUXajBEbTmE5qdduc3Grbvokpunx0SyXkMTQo+nJZu4KQnQf/
DBmizE2uJxHiToBjFayctgOJ2DF9tCmjUxK3LXxXBnlh2iBOPhvrFgmveekWGUdr50dVzmQK2caC
SmWLtTVbbrSBsVPt9rZb3PyaiQCi+AwhgBhvsEWqcOlJsedL1v4cL+C/09E3krnYD4FFyaL8My6S
XlbdqkTgca6fJ90V35XjHTujWuFQ6mfqEAr60FYkK2Gp5jP/5bY0BtqJKKXSXnl03tu67iHuJqMV
fNs+hZsScIBSbgEsBeSkUnjTHts/aw1W24O1/1w79J3pVAyaKpfbkFNo+m1nFgaqbsimNbZAhmRU
s+Zyd+fyWXL13wzTZ7AjTCyOq8bPcGLUqEKYHwyzI7t/6S7zo/efvGQ7p+yPLjnxvl8l7B7yoF1N
d5IrUbxxqzmKsRMy95cn3wxglMDJJDUGMPA0HSagCo3FgV5QBGZfk1uD0c4tVE0hUL8XVoijIx4P
ilipWKo91zVrHh400gz35HrPhdbXKZJKkGFQ2PQUF/hoqPGkNlZUieNLpyxQdFxb52bR23He0Tqo
2zcruP+SzaDkZ9uLcgicm0SJblEt/jkEGg0n6/CDWLLeP6qy8WtF02W1vPKfBgR/nmEfZznZ0TMh
G385/dMx2bsAzuZDHfrE9d7xZggJQboS4bzuJ4mbhKJE80n84vC7usDsyYnAswwQm0bVzYWv5a1Y
h8qf3gXUJuiO+f73PEYjurQ1V+J1Bi0WEMpLK9sA33QRoXl9aUVAq+xdP95b6HpQ8/m/knrmzmHC
s1ak/65ic6vKaDQySNIZ7PaGDuB3EcTL21nOq9B39+5MjBRjMRJlbcKtp0Lys5cEzAjUT+Dzyq1f
/fypBQ/gYfAII51rGHFCj0F/7/ANaY/UQ19WtyX0OR4akuFlVcCh5d3pTay02wmOx9vcu5RV93qL
v7MaEJlDgi63GnA8U3gK80zhikP4CMx7GUiMCL65LXQkSH3npRVLzBppl48YpWxUg3LEx57tNwDk
0w+VrVrnj0l+EMpRyi5LzEpLGVCOGszGuI/geIm7Diefn1JBqLAfN1JMmJprtxX05X/hkSIQUod6
jnLWsT6n0Vh1kk2dNMJzlcp51tnMB9Wvfz3UYvU3Xx5rA5eiuouqF00QOC/2pzVPNuD5qVve98NA
er8IN+9xMXadbrdWXMyFkAMsLhUU3SBFonrGviV/Icn4MxiTfPFVYEcP2hwcNv/iAjkB7WfF2vUp
TdjVp40Nu3gdCla4f/f+7O+DEpu48yhMgqtLVuO374hyrR7sfIAMOd99axoSd1bUEMEUft+Qzpyw
4YzVmPTmi7WkO2gwZCJ0wRX5DxNLnSeXHJ+SVCUBLl+zi5tovKh573vmmuSkwpDqjmkj+Eo9oOui
VOMBGWJRqNrNBlrgKBS6n/FKFt9yTiIgCFK2K4pcsfXgFD9xa0om/UO44KOdrGvPXdLfi83zNO9S
TG21DWJ5TjVxsCEWcHhseuHSqhPzMY3I/N4oEmmH4/QBqYm4RJW3wN2fkVPTGOnbWiUjZhNprp+S
aEqdPLzbpjdDPnyDD2JreSnoX/7xuktxSVk7143ER4Ej/J/r7hwjCN/WecTbFniMBWs8ZdMEw4mv
vvfrROKyaOvNN7OyYnuegPd0FlM1hkzRlssMA7+Frf71XkhgoQfGC+DGiYf8jLNUvfHERmeMDgYK
ezggM2GgjJbr00yWkBbGVTiisVFuxN9g2De4GEE0yycWkGuVENUHZ6ys39snN8n9Ql2m4YLCNSem
0QppsP2Fy6LXur5zoLuHguWNutR/cEqB05hLcovektbeciKwpeqnsGBTsLWOYC9Q3D8oaqGzUaQH
oFQluRe0sNX5fdDu0We98qbVaW2x6VX02dndUtCAJ49vP4xrGfcpKq5l13g75/He3XAlIr01MQmm
fOSlyn0hMLlgI0p+LL+68EjSkEMgMteqOuqcKLlU1bRVLq/C1P2JymGMkzAn5/uKdAMMjmFSFwRT
vhjYQMPbafIcMQYUMdCaRd8kZjoD7XyQcXfWrm0vBT5m9fmhSiPm8rV8dPKmffB6Yq9MU5Ui39cY
kitavv6i/YHkUiMS5iHrX93ycnYCRh21KJWinH2oB6/P2vwyVcFZ/WgcJhWX/1OXx9BEquB1NzzH
CdOIAFymyfjxPnX1Ed4Ax6SKWDU50CQ+VeSyv+LUr4i47VEfo/Zuxwag8tuRpD7+6HuYEipGK3AR
lsT7OeXHJrsKBHN+7ZZBNom5EQD1DWYw4j3PTEA2cLt4Xucw7Jg+WD+ig1AIbnS7J7+l5tMkce7F
WkM/nwEBHO30YEFelhxqOpcePoF3niFGbxArFJKW9JFfe+yo8BxsH+JS5yutxXCjx+AwGMnscW8i
35tbubvJXuq6pWFF6LTnCQksDESP2zrpTkAOf5wBVScZkZ40Liy2gS3K6fy4cM/j3XVTswMvsjNG
rPlaZG6RYh+ZizyDNT5a3QMzNolWv8J1d042ioVBmViQXaBtxTn9T5iszuaRDSViRprWy919lmE2
181vCznt00MBCB93s1S2L/XQp9DoaYOpv+XxL/KzfIF5YjcOgpYKFJaHxdlykceqWiluV9r4Dee4
EXHVav7ZpaZba+/dvaQGahFanCFGKqRtdVSrcLT23K1s7YNoZPbb4nGKeCpeExbDzDWpF+sFjvF/
1jQtvafH5MdRXJyxp3oBc+lbd1DaxE+Qx+4Y3SPpDaJzp2N2OWvXm/e3l6sZ3VTVs5TxsqKfuGZ8
abhxdh8ihL4s4f7f8A6L3krCDpdwLAA/hx3J/GJFjWwDSZo+dYlWVoPUlzgHPPP5wyujiVAttz+j
3Uc73EtnskVdKy918Zy6w9S0eXVlWR4rlhPn/p4fHlrlkAUr3UVZlTzf2i9nHUnw/TKKtXl5V04p
8Ap/iziHdxuVQnCcvG38pL6CQqcpW2ny3hK0yo6aL4c6nxsgAUAKaat3LWfCvsOsA8lFgaNEdqzN
NemhsJZ/y4Q5K18IVob1Ua5/sRAOk0jOzF+Hzhm9xDxksZRDIuNF1qd+dEmYxsvbdHmtuy3lagxC
+O80H3tA3vR/y1VgbxENwV+ERAmWvapz7gZsGmwlG6bObbGZ2ISbxLTc63/2kbGpa4dew0YeOz4U
9tLc8khADUBcblxBUsX1TaJcyxn8zHlDqXQbr4aRo78w9lhVUMlIpV8EIUk91yB4tMFs+Rh/ae6V
/A5HXCfAqxtluU0UX2etiPMVAnO1TUcn8WTHkJHmSBKAHCGdO6vq+LcS1TC8UL348yvrSWbHdqwr
5xhh08cTwCMDPGfkQLptwY3CZ3l1C6bNUrqO1KWnO2zehXIyQrtrLBP62bDa3h2f+a9dh0t/DQva
GA6WYm0xCL15ggWFrHmcng08s5slaED1jIbZYvBPtg5+XMF4Al60e+hUCgr4Mqst1K8IC7DMcSW5
Eew8x/7mxfSCj4lpYY+/W85gOVIeM/1bj0wY/1/s4Z9KBNmn64UvXUdaxKFatm2XDglh9F4oNJXS
e8oM60cbj3zoxEvbJGaITcTj3zq/TWNzEj0h00VtbKJvFoauICxjaZIeK7PJjs51UbtJHGOyFR9m
xw+2A5c2mvsf1F5DS18XOKOZqdLTWhiZE2ERZPsZrYZHNGBKVaDif+Q6y2OxM0gcsGfbYKsFH1Df
UCzi/fco9WWBWqfUdMoFpiXKHAiMd++bHxdvCcgF3t9s2WRfAQ6t4tI5ouZ88l9Q4jGANbBgbxZb
ywtCXeROJSfH5JEtAJr5NIH7g+MkBIkZm+xoo9r55aH5dvZ9t10XakMfQPDfTM0abMDNjJ3WpOlh
CheXDo3COs753sK+bKD7TVQj9zKd7Kd3aa7dMwC1Tapt5MTMEd6SV1i0CQ65/shjfntRcRwrDf3M
1QdGU+tiX3r7OaoXqP4ZD1gYc5Xy079a1va3hlIHQW3Se2TQk7fQRLoGqMF5gYmrB/i8fsPtHqIj
znQK9TJCB1w9bBkrpThVLuHyysnyvpwbDXSWbOm4gWmv9o7UK3gNN9Q7tmL+Q/9lQsq2jItu1pLM
wK35pZJivWqrpeHTWAbcvnBkpNGokhuRCRJhKZAek8+Q9HprQkm0DQillLJHi+H3stlaKusipahO
fm+wmUp78Mpkbd9wvF986dNuNNlOn4zMgJ/kY4Ew02YYhl402sHYpszNQG7hncjwTxWGaaRaNm1n
rtM5Ql29dUBIVkvcKdR5m7V8ZKyrIu+Ks/xGIU8hdmFZiGQVYEzGWR1sqYi5pPTruxvCcP0OMSaC
ONZeD7/RM80ddUVC2Vsk6OAauB96rQuWoY/xJBZ9ASQnqXpmGBkXXxsTbK0RgyizLou6PJPB6tdY
HJ4PLZ0u3ruaCLHN/8siocfkCqMt5FPaZq3hN4cX4Y4yh/nktOVDQ6o3f0qxTwKzH+SPMmuzagT4
yWB6Fdk9sFSZf9rEECXbniMP7KUEkxWvOb8tZMDb6p84RcHQVs/Vl3g1JP8uEvl0hLlVh+ThjMUS
K/v1+gMaAEufAa3lNdlTaMHYxjkpoekz2QTyRhhlyBO30hFYtz1cJZxP8k1QvrZuyQv4G/xQKflt
4F6pW2ZquRz9AGLL9P8DR0ySJotfOWry78EYyvLVgWH0+i8yD54T93b5gmNwKkpnR+JctNNnI/+B
eGEhMfMaGoAlbaCTzJLC9khzM3xbCKiFfnh/SkVHvwC0mkQDsuOGZPZAwKn05FpYGRsNcAZJxsDL
AO7JGR0gQyLrlvA5uZCYiR7hQVv/ivvtyxj3KGxfVV19KONVYV/vwx600fGVjjMOZp319cBJ8QV/
wuGoIljc83DTQCVSxwFPYmDlwWnFrG5GPFOtLxuBefEP7kSY3kufEIjhNn6gv7ejxx+KoW7ZXCG1
inHlt7tpBjYDlgIou1/unxA6eooJWfVJUbeFLSoUnG6MGo1MPHPM9E8U8KkR29Y6TZ2JjTDFzde4
ECQtgfAeO3ow1tf8ID0QRN/FWHMIgmqmqLESQNZ1r7T/wXjaMFAIUQ3kTxtCQFU6I0yNi+dX2skU
k3hhlNk5Iw56gRXSWl0DPR9LkSJXT6KAXF2LTcCuuws2+utn51JLKITy7DUdB88bsNzHZuKvTqoR
qIjjDpdNFZAzc1pNVGWrj6/2PU9zqvWBl4v2WFrCAluJ8s0caYtbl3m4hSaHtlI4lWzaONaCDF/U
x02k4+6Awk95zewJ37ryFkLZDwoDqrKKEvzVzKD+BH1dsGirIToi+N0A5p7DX3KRY/PbxIBbxTF9
UXtfFogXriTabwoGc5BGxTDjD6x0gO1a28HZGpBOC/1VWt4pWSWLLcOKH34SJaR6VukAq/v832Ws
S14sbi8RrJw9LscDSGv/fThACq+wecXWna1LL4Hj42yz+D8SXwNoI7dNEoEYCmUtqvzHtvlvv3aD
WTwquwr4VOiwoq3PxAK+v26w5rXsWDQk0+UAOxrAcH6Iid0LXdUa+vtD7K218XI+mNFgapfhLtD7
YXGHhpORNpyj3/IwUnnQFTAOJpojR431nl78Rw/VENRpI+sOSNsmzl8K+InTHZxIY0Ht0WZ2or1i
4fBjmkydnPz+5l+5qwaprkInfe8dj105BBCaRYVYeJe9H85Kt+t3WaMZZ18HuW/cdsPdWZv3SNHH
4LGfW+WOQu7kUz6kTargGQ5zbi12ETNV/6p8lu1CfdUcLqKtwToi0Sfg2hJ6/io7430kC6gPRtBg
bADLOZfMt0giBz3VxDw5fEZbnd6Wk/fuz9LBkTNfJ9Jj/oH7D6wAPMGu1zTLAK8dqEplX7Exkiwm
M42X46UGkb3dUq4DTnhhzw7OhdKx/GkpPtlU2zvzD5hW5G+I5XjO2laOESEZ01qW9TNs8OPBauuz
pQLRZG74SXuiQmiDUpCONlyL6aCc1euht0Ii2TI9yKPH6pft3rUb62LYrbyochU9FHCNRg1JfeDe
jMZhay5P6qttDGsvCK44r1/gKc+PpW31tqYYQOEJttHKPXAapXGp0o17/K72tellAyX1IMoLAJeh
HKwD1pVBgeflG8XWvKbwIO/i3UCl9nO+ooIoaZjhchdPXgVRgrRBEqbNVlhuYeu1jWPb4T/6jfcC
cdELKMirCh01+1w+hs+oA9HltvcDE5thlYNsmNX5Ik9MFpoSVIMgtq1/4JPHzoLOJgDtwmeaGQVY
xOqFK6k919QJQG/uZZOi30Q2BO7iMdHL/0GpUctRt3xTSYO0mUiahlbiAobwNtetjTC4JG8Z3vMm
ACKtLw0mZdB1QwsTtpQZmUxsTsP971v+WkpFYC4FBrfo3vUFZrYrGhuETtQ7/TEXSYDt0AuCS9VT
tucduNLVm4JirjHQNiyjB/EMTezNW3iy0UwcmOpnG6SIZbSz15nLCoY3givJ5+TAlpSQSqPwu52z
BtsswcwFKiu2eA5VU/uiQCZ4ncYujFcTMIohaXU4Cq/eMOQkOy2cbdEK34MafAZqQw2rp1olJI3x
M6wvHIoRtLUa56kO65Qa1Eq5OYMsXiNwlpCrrXWqwhNSngux8b6LBRiHJuxVbbAPL7KDhhE9HAct
AJ1eSbIZtfjYt26k3T0rjQTJNiW7eeLo7zQ9Wna7DUHBMqUqxYhX4upzwdMnbnVU8/fRH/EkdsIN
xFIZyKbdxzPuUPFZx8tQP9+SEi6AjVhCyp5ZBT5crXOf1yMWE1LxQKygT26gZRG1qOgL7tUHaUWf
oeC8ZdHNZXWTFSHhOSe+qrZ3yfJAsoBdfHuKkyeJOj5kE0l7wGaQCEmB5v3CvPKJ7d0azkd29LkO
hSKlw1CiOEPiJ+T7Fawv5JYPsEWQJjOiQgqpX9mrVigQXYJD8DCbG+OisqeLnRhVVki6/Oi+r7/r
bdvl+ghMdp75jM8uuGo463gALGxJWBVkIBUWZNgChMuAop+Q0zACXXH7RjcNKczTul83zWm/u8qT
MfDy6lFkR9cnXFAFU0Aauvl0cTm+eHUUzECNM9HyQj2xxD7Tr41Xzc4Xp7DitLfcKykRHF2uC1Ea
T9OSr1pz4KYbW+J5/Ap3jChUH5Ghsq80hDIDJQhrdG9Q76jVeaYlH3yaEqsKFCKyrK3NYK9QwZgZ
/FpvK5Rnaqie4o5GLOJmFC9oqGat36KVarJqp1jKRXSXPeNTKo/R4KUmFfJWv0GFLuIUSq2+a/Yy
yytyrDa4SSrl4NNMs0gDtZJ89/KCsVZAi6fq+FP4/HcAH1G8jj44pqEps8JI5K4jskvu98Fdr2Ky
UnD+15OiwUbNybfeJ7GPQCPcAELgwOGACkHtpY4+XiuPtfO5Hm7WtWUnIZy/gSrK6hAwqXLeW/5W
iqC3pjM3XRFVxHSFQXW6FvTbhMi9456mZIxRDpqNLlu1L1A33UaEUJT1oUcP2kF0mT8ICrraQv7w
sBf8Rq6wMhr5eoaeqxIWNrDu/0GCAtNjsZu0YIDwHJiOZl680OTV2cCSrHLaZtF3GFSzz/uEIVpi
9YpCGXICCBlWRcX1+plxw6YBUESJkcQAtfGCDB7RaCjMlh4OI7355dACvC8RJW159mqHvWUw23U8
6yDFWH3y43v9jMQEUztxclM6GhL75DyXzKgTSIIb0IiikfkCvdkKM/i7eDOqBT0mIt6x30H3QA6e
FDPnuy0JB1ySWfO2xRC1MYaHRlhh/hec3CtNcb2tVjh28dXyaJtbvH4sBJMmlZHJKDG4FqKhPgts
LR/IEyyucd6NTQe4+v/2c4hoMsklyNH4Kf0nnUFSm4VNYsCMlTrq2Fdp/bf0BG3KcVANWuuRAljq
QbR45j1pKrEHCIQlxBsSSYYZSsZNUpND0B++c2HwgxxsCEPgt9Y/+afzjIx4TMd/PEoydtOYK47l
B6OBRN4UOlzYsDA4BOq7lG9jUNfmHGhF2dFK8UmUoYyqU0Gz669e0yT+w4XUKOPgpGRafL8pDHjx
6nG9291FX8iminINiyvacYkaHt3gfzvpCOrsYP25ghMet5gdDSjpQ7Uj5FtA6uEP3j8QTKWHNHDF
DLrwwI99A1c0JvBtolGQNKtW2Capu6C6ZWewD6ASFRyenxWsDEVKeGPP2kllHMFvxGjlC6+Mi/O/
WYopfGANPYKUDDjiRgnnoPRCx2tKOV6TyC75s9VYA/oHwY2T+cZOaiJttvgMUSXtoLvmeKum5yE1
DEeQ7WFAnjQz0YEy/Pp9eCRhmW6ctvjmm5iwxVHLTzKvE/yRWaOWHHqdV40eiEkD7YPvmAg+HD5w
+VmLY3PIO5PgjRhM1SWGoKLsQNgJwg0vurgqqp6b0m1GyKNTNnsIatrPLwo9/9N7r08lWwDAoNZJ
4VvhYdHvv4DPKffw3cHQ+J0ud2pODSJHgTxpRA0NtEzZez1540VqrjMVhObcEWs647Basuv/Urho
F6kKWwJf4dzmShlvfzHgDxSXNzT8Ni6sVhGKJopqUxE7trIFQQNng0E8AgJdV/tCkNmnS2gIuBQv
CfLosUadDvpp6wojJzaPrdYprMI6NwRUHYqhefaB0aRVIvxtr9icOAB96wpsR3DMn3yaqyLmans8
tE1KRnfTFhng0vQaHLXaBGni/LfvSGZeLt6VNj/dKNteAO5lrfkIKaGPuBBmi1HjnPhojInoMDQd
85QVnRIEeIhlcuVLPBYJkkDwtYFUTih8fkXdb1COK/cJkER99DnlyYOd8l3vh7vavCR1KXoI2tNV
eJuJxehm21zJNDIy2mupc5zMExLuBcWnJqYfTVEys+eIUa2s/X8gXyKg48Uvo0IbjuhA171SI/lJ
mNKIDtA+OQhaABuIWFARq7VzEws4cAXOFrdFSQn1aHC7GYlbiHDEkc3NSksLbSm9q/5Bfqypn+k9
nkkOx4olnYTQyeF0O82JnFKrCAamdp4vz9m744geEn4BTY4MVc8ESrEnq4tH4EjdM+6XRjUMhlaL
r6t9SDBU3GA5zcFfz/eUO60ohI+F38L9+xJt4VBkB69PQUAf/XQgM0ci+4Xv1y8fqPGexvYtVDkS
ah8aThp6ywX8blkcNcs4XJFq/KTfbIgL6Dt43RIqCX6xBjH1T/lAxgroy2BuF0c9zfBUeR9/sE0c
cCGofMaubx7kq2e9nBQgp60UAfysmi87HCBuo6eoQhJkg4UrLPvD2KtZlMVsRo0MwH+ZBAft1UZX
Kx2GUdqrge/LBEvXXiDJr5nkHQIW3wuCBp5kpWZw3h40CNMrlyTFXyWanc19ygRcfvwipm3D2VDp
mhLDYdGXJIhr7GeEmi47I2abK9H8GYR7KRl3/WNcdS8AagoYrprn5MY1ZBuoZW6RrSMXX1YYNcIA
TyNhN1Ade7T97He/577D3gqfJH1LgBFC+mZ5Qtn4KPT6FMq7AltFanihf+bRFVec2Oa6Q6CtXdoI
gTZ5P3T8J9yLrOWIjbU4uHJKOOtXuhBRrcBlkONe3tXziD9OfnNPbnEFm2BFvr5xem+EH5TPsbdz
4CWF9L2VUX9GCZ42xV3HzMP2uM2cC5gLtuUZisaiWUtl80aVDbGExAiH085TIhD1gRqC3CRGU9Ka
U4uvJ84E+Fm8UJOniGkawDmWubCCFCRhaAiHgXvghIukIeBhAnsKGArMQTzvoKpVH+tZ0d6FlYGE
iED39r73IxpKcBg2XX9Wy/RNZiWWocLx9mzyYQT+2pm8K8+Wf210XGLQo/uuD5qwAzC1f3/wSsOn
16FVteWAbUBQhWx+rVHzR/DuLJ82ahsPQZ7J2pgJJB/RDl8gZjtf7ROizLSS/ucLEyJI3Mn3E5YH
kCNDsFFoDgJut6IuQan822dXL5Nca7Dc3vCbwfB6zw51h2MUYqC4jAt4b2Lrynf3XFs/8m8nS2+j
9La93/pB0hia4zS2hBv+Leh+XD4DE6Qy1PpE3FfEAn8rjyQGWitu0+Duz+HslwGhzz+71vNjQEDh
djLJi7W9H9pDDDLmHL/LOpL6oiTrGp36WDnQixiI3nen8oF37QCLHEWj/gf+ZpAaLMW3Iy4L5J6j
ibSSkvIOV/oUh7xHIt7kxtj8cIbH9JzRP2VwY/TvDcEx2cRk6ktU0uEWMW6SjEL2852tmAY2n09E
DJtKSujyyo4fnDsl3HNxych0DQ16sLoRv0Muvemjw89B9HHbfOVlSylU8aRJ8ecKH+Z7KhW1VvTr
MId3leDYW7FLxfT1JhfQmk8aqt5kCnh31PSm6UYHXCPLstG7n2vsmyofnfVlDwomugTGdlWa+aB5
ApboAzX7ZHmqfOUu9mSaQ4OVWvl7stc91z1e5jf0AWIedVZwL3xeMNBJx7nc2mtBoTVk+im0Tmk/
XLf5WBlnepnSsxE0oQqPkSFijNFBdG49sE9vC1DtE0ofJjgfx3D74iXH5/yEg34X0mZGH1wJyTls
e1PJmju+t7gWVvQ/KI6vM2fUfB1ORDoIJGEQvten2eLlTh/12trW4jNK132kia3eozyZVYxiu+r8
ovg4D18lprbOPJBMly92BZBmgw7wTJ/XrJ5Lw0JTmBTjkcHagnAsuxzYLMRBz0PZuewvMWjCJ214
jvWNaZSrAdSe5JY/5RRiq1+NIKTGafO6ezg7n3ToSn09db0ZjEmeKLMEflkqIZ8CVA+SJVwb/WZp
/EINTbAPiYBg8EM3bwvZg1HWS1Ybdy41Ir0qIkSm/8BUuP/3olQW+B/qlEqiVdiYk9LXZF5PlqSX
HoceEANjQ+BfK7hBX9n479yWeaY/9zCnqHPACAtTWX0/TqFb0d0hvgZwkJq3VDJVsk8pqJ42NN4d
A/mdS+2zpgvFExAWNUTMtntYepyEh5PM/kqGGWaxbJ7bxqKmfX8OvrFvSHK8NSLTByDEXD3PfSuj
AR9S0dPGvDET3d4/Qte8QZz9xKxix0P3MrdCzK0ysE21D5YFBjAAhnQgkymnGWGvCu9CbynKO0Lt
c1K/tU2mMg6IVm3OXJmpsv0KCCkd06KxmzDgII6LtoGhNOu7iGRJXHyYYKpYRVj+7JW9uY6C2qZY
SYpJjZHn/cdAhdWjscOon6W5WdoVNaBZbb0bKkO8vJIqJ6CUs95/Q59UBHJevUXsigzDJryNVz5x
lSmljjOt45l0vvYjp69bawMJqcqh+oHi/ht6PZVda8O/vecnKZVcsQwfjsac1VP29CyrFhpBQsSD
uOVTjghfHqCFcWxKtMl16qpbT/tUxcM9bo3PxCTTrymY57AuqOJ/RP7EaRegmGgbafuouV2GEUC7
mazv4dCjctqx9FCY4+4yRHj+nmKFNIpkeJwawIrP15kDr9KoLgM03jbfKnXzH40Ebxbs063jkGo8
+mitBpvStoAblU1IAjJeVkkDRYDD6OTyslNVuK8lKtc/P9RUX7GlPdBFA7kg0itPMks5SU1q2965
7UbIwfwvy/qoVVxoOpW6kQFQwGkuqntvdvKnuh7lv5q0a8NwxiaYGKUPfwMnaxJE6a7425V6fdU8
MGcSRk/QNTRYjFHWWOQmqczwF3QTsFTtwuH9zptfGKRnnh8gfcSJvOh3eojb2hdHoXsb9W/F4e0q
w0YFH5d1Ht0H4gUiVADBG/+bvSpViivu25ZDYQtDOLEKfzVs5yV+tqrG5VQJt75CBGXwvgCLq362
FJSOsb7F19HkBDBBBMC9U3rN07SV4TQ6IToE9Bbjrk+PgKvtLccJIhARilwFyOkJHPT0Ena5rV9R
erhYTYodz7xThAQ8z7pGHJ/bId0AaoypWnjZtI5hmATb3Sk785pMSNmqFoUXEf5YmMNL8vvgdLNz
4+1+b20vEueuhBWgbb6R65nsC6tZP83gKRoP9bBj6rlk+CznV7UCy1cHaEP1Xc6lsMURhh529jP/
pl+SvRBZSoTyKgI7UVoNaMKNeJ3FGc8vTIDzO0UR91LmaKmUGz0wSQhnmMZK7f8eIh2yIJLAExdn
BNpvYOb0mBb5qc36xLOMam4R7TDB0+H8x3eleb4oZaRPRg327CoYaVMirHYWRFp6UmZGXAr3pYTq
bONXuBzQJSfWpawkJsTvJMZjJRcN1TG2roXXd9G95USRzd2H+80CQ2wJwiQLxslqV9nu4gt01LXH
1VmRlMsCe/aWDG8E7ttW6IvMlR5WjKOBSzL+7tPkiE5Cte0sdssK6pZQP2lvJmFa0E/w68htthjp
+EzM2/Dql7jleGm86dQxej1C8pSLWYESgWfqk408pkoxq6hFlsEdJZHNbjZ8tBr6VHvIiHPimFJ1
mpjNc5ApEX6WP1O92rO8E0VDE9kVSer5ILLwBpD4wKe3QVCyEyuRrck9nODbIJPCOkQ0knxqzzSq
OaX01WsPTCvkvQtDkYIIOC0NKVKVIhhaf9MXiUk1qm9A+HWST1OYfOwxGyqY+I5qowNARO4EYXjC
whslLkFahlOWK728jI9ZHJ3mjlhtmy60dQEnUVkrBiqrScu+niLNytMFEngwqTRvP2+O+fUjLuvR
iwEkBtfXAf/RfLp5afrWT8H57Xq84grv3M1TOq62zkSoV+IwujTgSbX4VjA9TNPcvd9hUDa7M2sx
NX2g08N2pqK44C2CbpgqIPB69gosQZF5HFO7oi1zoN+1u6wpWNvCi+s44y0pPiETzZ2meS9pWd7o
dCdgJ71Mco9/gaMYMqde4SKlVP/cGmxoozv/XvQa64ey4zlcWfDul7B8IR3F97cP1XYVK1DteCRM
CmbMBxuuZxTknOY491hn6lcaxRShYq6/zjhqcH/jUe6WuTwsGlwfnzcj8dGvSe/wCm6U+3mvj62N
6xUjDos4ccO2RhMVBAOGCyqpxhBj7rc85DJeIsH81Ct7AgOXLmDqSDihJ1mrpXrA52TAJuJfcllG
4s4f4OQo8dfZ7wyaCckNWJ+bzOfg+TnBLyK3NFikxMAawD+SLModGIGoKZC+fwyW0hVXn9UWF/bI
FCyamMaxLy3+9Jq9uggkceqROIcJ0BbRfIJKc+8YnqV57PpGryIL5ddI8dn1HoVvpVbKB6Ah7ven
VTKW19NeMmdL7S/KzVpGFDhT5pNUKqvq+RG/cxUYexH7grognughqSmwL7vhQgClZRYSa/kipPh3
TYryeKmHseQ3KBXm355YNq5cR5FV5zEMrUDnx6pOlC/rB7RD0EdS9r/U8rsKlJw/84fCGJYxn65w
m+amenLHkTprukYhOlTFx4OrG+BTt6tltDrynGkxoIk7o5xyG7DLJwIn5xrvx/j6cdeGGExyId54
48T7IpCCIzFsO1iStey2Vym5oFROMWeIc/FJWXnH8mrKtHUn3U6a26ddUEaNpbLmag8XYPRkrLJw
o/Zr/nt0yTxxYBXSph53RQ70V8d5PXU4ZTqJOe2Ns//EKnX+lIwLbOvr2r+M2HmYXr7/6xV76sNl
EkWtIQrixtUqES6ZBCvwJlVJd6Cmg4gOw4EtK2WwgKyuRLgPZYo3mLqtdTh7s3+dj0Y3rZeGCBTG
EA0NvaV/quyokSUmFoL/cYA7hvpTL6EVJ8wiacVoAfhiwpgeYY83WHxdKtVaBcns7QBNV6o2a8ux
YuJI5+Zv4lh7V1KeEuwtnLZrN4HqTYmPh+m6/8qjBD1/g252hIEis3ieYmRljhN/WcenO2lA/ldN
js3FDIKd2Sg/YXzM9i190K78nd0LisP0mrTp6zgx6oWT0uKGNYSlN952KDebqc31roHBf7TmfPG+
x/7VnSSWg2NY9rMbIW1KNcs4mMs3rHv2E4hPuYQ2oIPMZ8I2fVS9gdg4UbP+DLX5GiIEJNlvsbZR
khEs2lRqh4WZDkjQOhmY5n9eXnM2+x5cwY0cniOD6OGv7tDVsLYi3wqlnCqB1Y1XbmBNkJ9pvksB
TuAiX83O5D25+H5l7tiVQiyic88ewxAftr5CrkxPHeqBZTXrHFBbeOr14nF50tSHK36IvgMgT7AL
1x0pQlgnvu06yKJOiZvSU5V1BOYI0i8OfPhkrGOT4l/uZU0V42Jc9UxRu5h0Gt2I7VZnsdDeoQaX
RQmZXFYdHeCvJEb2U2UwbCLHqRNwh7g2uVmFbeG+Wrhk0zNQUJwBULLCaTSAi0tfpeeQZg6FkTyM
sWwseUD/9WmmvTdYAfMi78nqrEjOnSsnwvQDqsMjhTAKg+6fOqMn9mgoXSXxb9r4Eq2ZfJMC93bR
IFsq+vmIB49n7WlEb5GDyiCgDzTknOS1OrjgkQnoOHHUH5kQ+chhn3sIEEb9l56amJLz3SXmJkJV
wa3TDYlCT7quv887WqzGbgIYPJdjrVrfvxXX/ZVMJnxznGCuYWB2DlTTIqqb+Jr1TagyH0URk+rJ
l0X0uJN6i8lwyx6I2IHPs/wYaLYpAXJnlbluqFVAEfVlUPyc45hghxNlx2SGtdaW8vPUw4had7x4
yo722lLx4QxbrN+e5qAlUr0TgOR8L/P8dZZbi0dnHTLv4WRUcHYbFNRDJn+bRqwRzq4ZTWF78Z5G
Lp+uywVzn8Jsboz8nuemVMtU7cu6nvZi+dXmg0PANJ5wJdgKwNz1BuHcEP7VTwM0ym+pxRcIy9EL
8ZnkbDCpt800k3yprKUvUgxAwgiVRt0umGwAhW5AafNPZQLrFKe7RcfdTqld5BhWAV9oM87Szl2P
4kuxUok2OCpakKrzNaLCzk87lqrL1eZBNIj80L+CuP/izpdnwxdTzC0AKSMBK3eMoXhFnOURdNn5
Wg3+PkjIbxoMiu2pfNPaubAwchRqqFspWR+9yjNnaOU09jTWbrKw85ne3LPMaAiW08eghv3g/3oH
CTHL05IwBt8B5moj4Y1Zp9ljATvYDjS6N3GI1PSZqu1GUptv7nJ3/c/sIp5svDGGsscATvK+N+R2
T9gMl5rjCg62zUOP3jhjpqMzuZjOmTWvmEAiXmHGzu5Yy2H52nFOt0qVR9eyk8AsZck9VrKI6Qf+
jiCtQvO3XKpRBdI7gVAIhz362fOC0EXfhTFhy4fHHUbhnv1vMFafaI86Y/uPRK+IWGJbebZFD4S5
tabC15G2F0RVXm81K0Fy/CdFzM3dI+UEHiTe1JCfluBc1CUo4dZuVhpW8gitqb9Wuue3ybAZQeS2
wjrTtezqWME1O47G7TOAOk5okwP11s11YMmTmwU4pOVzKGAhvwB28QniQAC/pGGpwdF0XE1bp/XG
dUFKtKmtqgYLyJvAdF6I+JP9QgYiZ8nscVgSEv84ThHGVNV3Gfa/nsO3mKoyVgi6nMvOrGm9zKIa
GYZlo0/8/k/saHJJ2PVbdh+1tss3gpbhBTIMfaCSZGzShRQS6YgJQAze9Jn8S79A2Q+nbV3qdGxz
FoqOEHKnZURIj0J+/e6Ce8E2LNN+uiVGLE5Orcq0mC+Qve/aX27FVT3/XLykllaFiVzO+zkB422M
BOvbJxPvjLfgb0nlvSCuZCaGfOOw3vRvdQj4I9Q2TMVOt/Ffwv95V9Msm231TzIiBt2BbKxfWlhZ
ax27V6ocTOBuUdBLXGQ8o4gZuuPbzSZQipKDjTW14LsPMEotoaPCtDJ77widLHzd3+kYZYqCr9dg
eMU8GjXwVwa1kKbJ7U+yNtydHB1cjbP1RgGGAaY4KTRkaopG0CcjHectW03R24zAXeFHpLqGeW6I
qpjbGNHDY4FPC3Fphi9cLvHdQ2N57990h79PyqiQX1pSDnU+xNiC7wCVbM6xLbsAh6+PCSSuI1Dy
ZA405dLJW3dSgE0+msuu7KSWzWI4cOHqPmn8brcmXb7rIfHPTX+H9T4PE/F1a71FJXPuRiAEYi8A
gCUtGQPVhpL1fYZOdvmOuPgoPlgRFpXrQYRDgEqVgadg2hdvcnsF8gb7QbGN44mGd80C+45tgWro
v+Cj0hUXpR/9Sey2Lt55PXZos9sd6hCWBXnY01/+E514aKEOuoWfniYIMn8qc1yHw9GOn1hM5eWE
65bz5QtxnGrrfnM91Wlt69kEI7y3qyXcyaS8zQV32fTNUVv42WEHISggPMilfKNToUFwmoh6pClX
ggKtQgFD/P0IG2/YWSaQbgBklvOrblcj2+IzmQBVOXfT5DdUNGIKUjTSBEiZgN1O0FUkam4Zj6vO
5eBCwVpc/KKaPqkQyIrSWvgjK8MwoghY1vGJhAYhxKoD29EXtZr9T8vDc5INo9X2dEOQ4L9z7hbs
HWGmok4gX/cQSwPEEuyX/3Q73UaiDgieQQRSkeAzcPsovWqHVrpZh7PzNnG9hU+Wqt8GfyYpE6mK
EPLdyjRZuUUyajP2uOgfpAP88H60GAIkEFus3hLC3hhtvz3tASokzcxOgRkOBefDpFwc8GQqI0x+
6c38iUBCxRenAiizVuE4SchCkjLJ+yhg10HtcyX0fjPpEgylxj/lfEuyUB8B9uafKCbPGR8THw6r
Ki2IiYPAN9JYwqNFozK0O52+a/4yrmExNUQmwWiskTq37YsKCCLPnO9EJWgsapB2pEehxiWeXh0h
7/+D9nzNkUHV7vsiGgk0tmT2UxsnSjGR31HJros7OlCNqtfzGyw9Hm3NfuymWRASK7Ms+37J8aqd
jJwXjvxAnCpGgkMszy1mflBcsicQTviZm/VN9A56pKeUiXcRdyW2lDcv+prv3UZm6W6IOvkLMEn7
54rtqKLEfBwP1yoV6yHbfZz4Y7Plj9lf6P2KCzPYdPxWgFDHqHaujVZtf/udBLuEbNkKHeQm0lTo
uG+QUonmBc5+j2dsqjdCTrOzS760LnS/XBGPEOSPck4+3Eko6nh7kVrbGF7O0hRKXFZKHfSoBlWI
e+BK3BcgqeuqdA/C8FGzJkQS0wfboz/nRMl4rSLxDIvafvUUSCebwyCMOBJTO3NGqcflVqHO7GL3
qZVPqkdsZOCnAwdQU+X23rK1GMiW7kYXAgpeO2fJTbiGKOdSrWw2Svv9fIGZfNIRT9WvljyH6CJj
H2rkZHGKu5R53UYfRkLNTj3xwkipOyWidZkVntxHPwbwASG/AzRs94DJ8l7MZIRkxEkRQWcwUv0U
t+kvGcZ9DB1V+XwCXBDLQ7fB/dopqlFIkkqi8eMz/MfLQ++uW091Ss14q6xn8JKIL3d7o6CJWayc
m3wYuNTDpiOj8aMk8hdiRxHne8mpRGA97TsV1lEU7dDHjinskzNLALhUQ3b2zkUWo8biDTB6OGGe
odP5QodSux/Nl/BXoN9QvwVGVQMsjPOAQ/Exhx4AdkUynMld+AXGvJBKSUjENICKS+PV84IaU6pB
vrB51Dq4tbrUE0sfm057uT4XS3wNzKlnNiAS2YYpIRWgBy5+VvHvvTgqJWYiSNJe5DPydWbMs4mZ
4usFeGep54ATVXdthoDafz3Kszscebq9YrOIeKskuO/j+uGBcX7GHQR3aUXaayBnnZWQ1yZWkorS
9fTMirAMKk3xVnZoI0zhVWEYG1HcbhtK4iEJhR7vF3HkSCLgiRmNoLVOJqXXZJL+ECwjQuISNUi2
kjN5QicpTOTS0GuKd7QdjeIMWU9+D2/34G5wcCkruAAVUDDem/QnEEygi3V58f0kdNkWKV0dlDtH
9bCO56pdSQwXC2yKJUkk2LEe+fxbxAKcFwkI6lx+SwzZ116cDxAtEUtttRmxcltq+w2P+Re0nEIK
tMR6DjDDWTdGDd+Q9OvNsP3EAC/iGYbbCpwQWFL/tjpIhKRWQuy0O3ImiXZ2Ktr5XKjP0v5MCqlw
PHXFomhfrMT0AGxRGDHg8Tr2Bp0vMkv3bB5bl8v1CiqMRpwJDQv4UNr9Z4mP9JniPSHI+H9TyTuK
I1CLfaNBvQDk3iVdsudddqtWdc9AR/LqEu6T83xrlItXT8GsI89MyKP7JVrQdnkjbGLmf6VDFap3
Uoxg3o02MTv/9MypEgUhDwThXem3SQHaSnD5O5nUzTtQcsiQ4RKH/Urbr6jGoxwOU9NsRXJcqPT4
VsoY/lVsTFrfVmFguLfAt3VRURvZ6+HUaQ/3KEOEAdgWA4uXBrTCod674Vlb15j9WrPKfC6c+8HP
UAbVh/z7c98=
`protect end_protected
