--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
g/Bm9xwWL9Qts48W5Iy59pp9TEq5mActhrd9TjhWG+vOpeOZ9xt/YMhhC/t7qozh2ZKhST15PtZb
gAqR0hlOyWXLQVmQQ45eXM7n5Y5/p9HSxg7qhjWYVNjSY/FQ+YInPA9Q96y4KKm8OhhdK01/TxdA
s/QMxLpbbllm+5kS8ndBCyO394r4ALKFgfsV97CeELqzFAU7liM9kTIz+NmQ7tGVrhsEOh2IvHAz
4ULNuxClWUDl72eIp5BiFiLVYlKhbWQtl7whBvUh0A7hdGcNkdgPBn/eMF1XrZs+kOSwNIXHKuOb
d4gbGGYVisnLPPKorYippyQBrLbrm8p637gU3Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="IjvEL4u0rM8BOc9MSqJ300Oc5hFZiubGTIsRZ3Ve/zI="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
KLgMvLm35A2LH4/BYXTJ/42IjUwAnXqoPpd35VKCqOXN2H8+TdEABgnBvvrYOk3pz6qCy0rCPmcr
zAjJ8pRgs/xJd3yjaMFDW7MDcbysF2LCdI2pkUO0vdFtYtTCSzQywfL9zJHwzyvjyFT9IY33zF86
aAGhhYkXNEd9i1fRcaM5fT4Q+tmAMPWDCG7SigU74r9PKR2EPKIopbfE2epVdw2ojb4kcEWBkPmS
SPpRiOBY5cK7z8d4R1jJOPpbg91D2K9fn0LIcqI99WZwzf+p0p341ijynE5SVK8GfLEbXXHx3E7A
yVIJj41S6asGPiXUpkhxGJawcJ2VqKYxHvgisw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Z42W7T+Y1mZUKIOY7U8zErUlZ28aKj3La20ZQlO583M="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2512)
`protect data_block
/XbBUfpQLyBDH+qL2XaRgsnWXFCkX+8qItijjqbwypbFdHAhDVNYiy8TdVhvlmRGVdm1vDHcUeZw
EL/BT+6JJQP1qYbVaKjFfW8mtIoGY2bsJWBcGcwZNkZn/M/UUiXz86lyPDgVfGkpBJS8tIbIlmEo
hIlhoWAbqAVC6RC/XjlYTnQBDmXmDCNh0UfXf+F7U8U1BM2L6377l1yUNjgyvF1+UDwxYmbzFV3H
u5jtsutPxwIQQQya+f0BzzV2XJKfOqzt9kuz8XWeX+lmIZzk9kB7lFgL2CXcwj8LWSnum7sxDtIY
d3+069dxgGhq+P7NUyLtrl1mv+50Mu/qTe8Dx2HIs9jipxDWBDEwphSkw61tnjaR7FINxSQdRRCm
XlhBZhxLTBjKOjiPQZqrIycVOCaaPQ91xAQvN1H4zqs4N+h50iKMNLhYZolgh0xOXmOymKqVDrnu
Tx15E3R0dSAuUxONjYmeFYFyEo5dGo8RoIPaac61Wsbvev/gcDzvm0dKs7g0JDNNyfxVH7Cv+mvY
fwgYFc+EjkKeiyp8hwgW9kEMrJStCAkbd5LIEJlB/trgaqKlAgfH/dMllcd0GQs9vQOY8L8acwU3
dr3EHf2bX1hDLqlSCLnSnekI5CHskMDxXNuLRRjEXSaE0wWUGN5O+VVlVgb3EEStP8BcOBhqJZyF
siyurQMvWjbGyMnyc6qSHaV1h/jWGAmBMm3ykYojI3ks5SHv04Ipk45cyypDXqfmTGzQryLYHK4R
qjV4CfXfphNuFptPYQ7c+kQ82S9I42AXM3vKmKZS4B79N+JsGzur3Qtw48dGszOBTx6ey4wr+z0m
+SY18s9e0Q1VUXm+ZFwRcSTKXqs57n1wVjOn9re1EceGq15duxjK3DwcBdB1EIx/+lzcKbTRxZAQ
7vjAcl8La6dHbTrRqMcWDPJPwTtZI2C8lK3G0h8Lv3z6MrFEDBa3lQlcBkQg0EySZrXWAlcKZIFT
EEjtAaF9RHTJq3bAPTi/8Fl3iYu1Q0djhVm4mAZFPETV++m5E7T6T44EKWUGJP4R1H1ukfg3dQne
K7mPfWSV+e3d1+9d2u6SnvXY7Ud4rtPqVDJpyuAJdEN6Gb0akNX0dCPH1OcfapGixh9t72ovPS4x
8dvFgvQfI9GfsorbLhu+gC55twCiaZxnMyuxVCm3DMqLZK5Wk63m0JdD2l+aI5/XXFqWBNbx1SZ3
6FITxtOaWNgx729J4I+vNvWE6TrjnKCjyUzzRVCe/QDWNMIVsbZE7hQROuO4Lk78Chjen2IPpAKR
8xjhyAIAZsXWcADNWYsYJl19EG6o/QE7Jn/BOHBysQmPrKHdTUsiqhIEPyn1feDodEvUiB/Q37dR
b2j38m9RYNLgmMFKqsWw+vZ+sYQeqxskI28DUZZFgxq/MvjIPuNo047ws8Mz4yJxmRx6TK/OqFJH
+kHP6CTiN0smjS6JZ4cOE4rZdR/oCXCRYY72lCQjs/0bqpcnSvmvfrSC++kQO+nSXSUuhjxRxYwz
cDa5QYXGoILvBWAXVLeiaOzWI3ua7RRMZrMsrQqpZtPyifO2/AHlnKFKLCd/NKnpG+NWvL9Qyyfa
pH2PONwqhePLEK7aETKoSsb3Z4N75bqOxwSWjx9gpbSCUgOBtGrhjrfcmf1kju4lpbA+siDixib0
nILqUT6wjtEXyDnFk85a4bIdv7eQSbrP+y5uKH0SPqufxAD/W9kyVbdeeaL9pA9eGL5CrCoqmAss
8npjj+2iop4Vj9z+YwN8StO/2Q8cU12GjsF0zRZto85PTrbivBU4zvwNx9cHiiHGhz67w9yDTV5k
K11/XiTWtkVZSj3PyGAi9wheCtMRtVvyWz9k/TZhLB16XroWYln8JUAixYbIsUKFRHq0QldJrYmu
hK1rDinzqsyEtp4CC/iEQqyho2BUm9XgIPKOejxdOVaLxFa8oowE2XqaECZXVLTVqtmCuTJiNeDS
P3MMKEM6j/oqTCrlv1KYwqI+oexQNsNiDlYQrYEeY/fLE5yEe8cOCjocIes6zkeg0ojVNgZFfKPu
BJlQsqrCzvvp2ZuGBe6DWqYZQetQf9V84Zl8EQF6YbieaJK0khIcI15krpDgYPEo8LWxqdAUvxUG
rbtA1T3PdWnxDpRbQBzRC0uhR38vnLtcXQLRlBPvoHhn4rDVndzU9tb0ASnZR9XWSDTljjFmboPQ
CVQ2pSpt20EmAjOcw9PW4XrtRt6wFvaNADPHYDXim2uOu2TAqL6OJNOaThg9AjpgEC7aB8Fl3fsD
7vylAevNDU9FCyJuWSeEDKdr9WI4Q958zVdrm91px4a8FGxxKQRJ3ikiqGyb7m4r41QoaJGnzGNr
fmbwkO0KRDIL2W807dTcRybTqTAtFPBVrwJICU0lJ8DHkarCUpbX9hySTEnz3PWMJKCM/bMTAM96
6kT0uXEtsq/Rl7eDfMBWmXW9wX4lAxZpqjBKae3zdTbtUGgoznHYAvY4Mlmputeu9K1cXl+N6Upc
v3y6Xckktk8UFqswg396rFcqu/Fcdnd++5DCw8SF3Fsn6+VTvjms+a5hWqF8vkIzzTC/1NrhblcD
HWZXss3Ao1iABQ/wLqd+hnvNv0AbMahpP+wygfHERXa/pOafK1G8LCVJzTy69+ImZtVNTWKSCSYH
KZ9YVy/V2PoNZ2/IrjyC96yMJ3WletUTSMkbbtEbJ+L+azfMs2o7Fosp6oR/Nfq+fKxBlP+6iSSc
kHNMX+62Mxwg6/5BEgOOCOt8PU3HYQGOJIWd1fQ8hYwZ7miNQbGpoPYu3x5vV8qGxzANCUcjTRmR
PGFdPzdKIHNb7EVObxggqVaX5JjjqIPGRPmSEipxh4uYGUZC6ZvOaID8pYWyl6x0lyY8zWC7ZxzQ
AaJlFiIcx9PUKdfsLYckCGGpAR+4dxMTj4o9WH8I7ZjXLukecyLDsQc5VxYQIDUo84vfSw5uMgOA
cS6ba7+5T+xM6CGziAjyvV8+y7SrLe8u2aJGXTpoSCuaCTt63hEWawiYv2zQsliXlJsa/p90TiVA
RPS209jIsA4gkorF1VKyvJfm5mCWU3lamgC7KKcoV+SIb1MlnFltQRtCPCwVAgw2GEcIsBbE9c0q
vg8APYaiH0qZxOA3bto3VPLc0zQcVQ2T8inV6oAwuOa2UkuvwzaG5sp4CjX2CNbHoSDCIlu+wDdy
Cqi/1b/UgBs3+qbri5Ih1WUMbNf5ULQj2gsU9pZ/AJm8T8ZPORH2xIuog0YhWki8IqWNAke5D8nn
atJFud38h1d8RWwfeYMBj2NO3CrEgfUyeeFR1WMsPHGp/kr6+MR5mgtYudRHd1aAJDB6wa44IoQs
dwY32Q==
`protect end_protected
