--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Ov6Gc1pMi7Ha60jTSswAM6VZbOUZEguh44flpc259YIaPCApWQGcELCebYA3dono+hXRd1qMDvP+
BlcMyPqqJpLZ6TYGP+a2DVFnOHima7SaCAoNGuqEJ1PvUg7gIQxXP5jaPgS3gEbDuBvW9+thWogN
H0N685gD1kKlE49KisvO/Fvo1cojXFCikUoPvjlaetq4d1g0YnTGCP7orhDS1GoujC9R3MnW/ARG
/OEaiiSMGIIbXS+SQLHssBg2OrkmamqaQqxooRdCc144HBuA0RAJ2QKmDljoOcJRLpfEJCv0w8lS
dH5mrxsMHwzhwO01W0oeHc01NpzSL+UbNU99mQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="NHl9BzoVjjMGQNQcgS3w3zVzLeBaNnto9WsCx7tJoQ4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
iIwDGdSEFFa6bD++AJCL7MI7t8td8TNx9m1dtV6KHmpxmcfXiPi/1uGfvTG2RTxhV5MY7JLYR6cv
PrLEj45aKah+avdYZQOViGwpWqwYo8p6vQIZ8blkpSJ1z/5LTFrmulTReyFpPEMm0HrSGObdXGpm
fb0WMLc9Np4sPAfGiSCUpMq02qzQ/1woH3JuqbIz6nyU9K6dD4ydsXIgkUSSIRkthuYyiek7oy8H
LlRdRvKaiCozmgOd7dIsO1IpCBRP+IlI/M096W1Sybwn/5a9DIfXEShsPWZLYDM9C/UZ93tGU5Kq
pb+4WGMcjTENkDkSHJVNUUm+T+ooVUYHBNRO6w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="aKNeIm9pATgYcQp4tRl1IO24fX2NoQN55NZToI6rzaE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2896)
`protect data_block
3uKlkzW6hj8XxU+JuH3vkJOshcIBLzw4EdlciHqDWxzqEZQhYKUaU0D7et6FVwX1yc5B60YtHqma
2pY53WwsjCd62lon5Ca71X2BMKuvz8zWp3Fi13e7GoAOQFkl8nKahj7RfFeatWKkrTEdY3pcAKwZ
6SNDzF3fTvx3YYQMx/55em/NEFASQrKyICW+2J31J6SHre5sg9oBN7pJXMWVcyag2beWabKVsPYW
RyyYlmmLXRHW1VOjrJrqJUfEENeVJ00FRx5iKBqWuwA9DNdq2j18osdTtZeZNq6WUj/GV6h1s9kF
lcyYmr0vWfwxcW8sgfY2KHCqotqddHtkEmz21nZUHVEy/mTlYTsaWRRwr5FIQw86YoWOvbE3O57v
t2XoxBTBl73z5lobdghcYZFtP1IVMxAQsMbWeDU0T+KRtJ+32Im14DOyAFTYJp3xv4Ldp++f17Ew
cDNx15s4PLpcNpz7mQNr2zz0/jYHl2RMelv2/7396UR5716YfJTsnf7+t0urTk9Ba7a+w+k15pcx
MplO412wq3PiwWWTHCOuQbube4RbfnxuE+9euhaITxPZnr2MkxVYrr/dQVkzVZT2m0+FdWoRzcbx
0jJQLYIDfkPF9Yj7iSIDE/+vJNxMRaOmD34Zkr+bkCf1xzijzXsMajypW7eK8ovtAbG6Fl/XlhWz
Nyxst1fa3DHt+COTeJ0QgGdW868ycuhomNRgEwmPWLGleiEka51nsShPpKEqOzchZMRfrKWFEEdL
k3HaKzWI1PMCcA1+C2Vg0S26rLz0w2Jtd6v4Z5hzmqWQZXD53X3bzASR5Jq7rtxjoaTCdX5DdzYz
GLLiwg+C4qHmdfbFQLRDz63Aw43di9lIc3PEWjAzYdG3tR8BbBx7Xwo3soeKEol13qTgMpJGVaGQ
5K13qYLQAtVCJ6i/MLsh0bSwe71JBkZmvRsxe0UTPm+fE4NUN1Oj8jr3s02zhSoxbSKf6Atl3SM5
Aj638DKIsEVxQ50hhJZv4AAONM6mUzAWp/DFfQhJkRGKYmmGqoFk9iGf4QrpCvJOURvYF+xb/odD
vaAHCYhX14ct/dIA6DIirgeiARkE6Eq2lHYpV0bG0v0d7Bnr7YXkUxdCG/LGBVPjEgVRwSM+oWev
OFkCR5OfJo3UVFTSC8BeLe5luzL3K/iu3+NBJ2WNM8b/g52hQlAsMmB2ukIg0bwY+awh4cReWBDl
G0raHOOaCCgyuwlcv+q9cTJhCksXD/IqmDNh/pE27zZLZQTy0tpkWFgYpMJan3HkwhlugBbcyFe/
a3pONVavEpr4Ds3bi/Dc4ga901hoGJVFgXb8CSvO0tNpcBMADdsFmZHg4qYdSuXg3q3Sdzh/PZ+V
wuXMtwc6Egcdy552BQVM78hsTIcTHqUWzV3SsIXBOHVRA+utzTL+3x3j09P3aGj3qVM9TxxVNM25
FrdYxFA/S4/cbf1d75b9i5EwuuInx4mt26OiOidcIfVBEZJaqXgSjSX5aTSxc+aO/lPrCSXlPp2C
qj6GnUPIriLlDCEpfsE3AY/quvB9z4mN7oM1yVNKixyItWE2CmhLgR/PGDhMFQTGdP8cps6M0XLu
WsgiG/Ev3Gy5KETJWfTdD2eQYNXWYqOm1ZWJCHLLVSdYCVdyWIWvVYaHV2r/6vRNVEZIjUaMTddN
LYxZ5e61t1JRIwUhO2FlxfsnAOcbMalC43WqQCryBY1yqXRL1/QYFcd43UX5SWjXfORYiCOZw7fn
YDdV+IX5jL/4N5gM6WvT5MqfuJFVh6f+EsPX0ZEfIiwDDi+bcZT4pCxIuiVw9UT56yykr/1jVK+g
IGV1bGQG6ni+nxRK5uP7+xF3ZHAR1ByoX4XSOU9ob0EZp7tPUTj79dlycqxXXRolLEzqYVjebR0I
6lgSK2v2i2i8lzIoUA263hyDVHPdm1PIe4IoVsgJvL3uWyUbnf0eqzomo0ks5UjJb601bpyBuFhF
1eWogDcZqX/5tn6CPC89tm2qv9if9H8DRwjCoMMyhaoyIwJwSFmSDvbgjgxp1qz3BsldS8CFiuUO
vDMUVbl2ebzy7AE/saIBz1ZfPWR5zvYLCSvOYwmoRtzG2lNEfAxGhhq3Y1Zr+7aq0UHO81MRTlWQ
R/QKPpyPQ3xitIwrEjtO7wfj8bLMdAZO2AvjhjUei4gjz4blSxiIO2euFiHx1ZguOjVTWSechsPM
8AzI05EbSrEWlPvKup293ze9K4u0ziE6iuEubRLUymZOUCyqVp6/5vk574nXDFd6xTCJeUr9hB4N
9Rsk01EbeKOohOdTCnkn+rW7fGRnT/bFrFSEJu/tGTQE9+x+jBAZA8OLLYeW3BQJQCzvuVppGyzK
OOUZnOg47ew+8FfbNgjq2+AlFxr/g7g3bcnDm3Mvco0urawbLAAwvQm6oGywYRzIkHj6foZlfjA2
FK+MOane5GTPlL/c6OBIeyUxinP8VT2/pL+9YBqJUh/upulABv7aZlzStqty4uWTxCGwnhuIk9Sz
ig945ot2cUpyt30sKIFnQEUeiU58vzf3zIloGTN4+d3JSf3uDUuq2Kka0ixtdHfwugZCmNT80wFn
vMYlHMLLhlX1laR2vI9W8qcljp9lz2arSK1xwNmEQZg7sJ7kJ8UgkPcBK/GIjAXBXYOaiNtcrjgE
ZUtMOSVtzsi1A/R7VbLiRJW790z6y+EfviPDsuQm4uxLcZuQkbu6eQl7NT3Fp4VZNae9T7TiuP3c
YIdEMWOkWz3q1xNCKc6nLjGnwu5lkDvIJ8TE7wI6h71kgVbqkbYSOlUIYUY9YYODq7QSQxiw0/TD
5RD+3TQTZ4W5xtp4N97xpiD4qOzTz4LC3+ucQ0t8wnov+H1VtlPU7Y4O/YfngVVSjg2tjoliXe+K
sfTzj95pB08B/MP2ef/RfTFm+tyNnui6Ao1DWD+6zyRdQcgO7YkigPziN4xbiajygV+sVfz+t6Ly
2Qfqg1y/TXSt0wp5LZWQffdz97Q4BTw7DYm3oB64tcY9X1XlFu/akAaRh0WNim6uT21pd7dRRaSl
6HQXYCcrTYL1vBZDABOkOZESVZZDlWNOq2ZyWnLGajTZUuDpe1Rgbo78j7X3ML3h4aXQdi5B81Ok
de2anYUCgwi8U2KPgA07/5Z74Kh07IqgKRLfTDhmNBpqgE2ifL5L3jtBCG5k6lGf0aqzcNscYqzz
bP7tSUOBYJ2EqGSR9B2RgPQm2i1ua5JrmRt2i7ahXFTskdV0UpThaEdFMPkC2YC6psGAkGotMlm8
zeLzxO+itTPJ90i7nOsGGDezmQi/qJyekTWPcvvvizoJKXLxjnu0EW0mVliaNZtOcbB403ji48Wd
71Hapqgbgf5NuKAri/C6qNpsM3WrjRNESarTZ6RyvG/LBSpkBt7+rLNV03uEk5CMHkHmsWcv2t6c
nMI1Yi7q7+401f76Za7ZzcRO3nINLJqIG5CZ99IrCvUbKt8BAPucp3wMNyhB8ABe0p83s5xRLEze
W3Hg7+J8b64oJhE5v+x0FQ+PocKmad8B9vMuSDMxX+uwbG9vOraXOqgHr0fU/QNRzbMNMMFLHOMt
0rR2HkbzbFQ0GdzTHjub+cyewSEAo9wHVqPefLvPt/Sm9+ciVLvpjrohCIA/9ySntcKL6xjal2Gp
oEGRTADR1gWxljzLROk5dtuKjmptDy+hxsB481zRoTe9gZGSCt3qbNOPbGwslXxuwYGwNYYduD6K
QqwPc59mDeIHrZSfp1PfxCwoCWIdmpXFOrEokdqtSUW3LqT248K/oSgiS+ANbdoM0vSKCxHe9ZL2
omS+8JLDDnmIhUj6LR3c22VWctj2li/Yk8BW5MgWy7RQYqoasi3UKLwS8paYWA==
`protect end_protected
