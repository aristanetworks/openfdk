--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
iWToeBlXifjIFnb+mpj2B9RdP/+R2dGbc09sIx9mfBT7UZT28rrqZN3bem4QI/lnOQJykbo3GbLm
z+ljP3EUduD0uiKUb/m9k5dS5QPaFgt+3cifS+ropwS08H5U8zhUlWIQEwsdG2wPAFvfgKmGQ5mP
FtWQ/lFPSUvFgClMA6rFt4g6WmFoCp54CbTyNc4hg4ziaakv9rCt4FtNlG8ylEDJpMUdzN8eSAGn
kQpTokzhvziQVyAW8KJY3977ImfnRzPXR17AqsTVVq557pLldCIRKlmYdYdv6JHIFVLXTE+tqTi/
7jdiKkKOtmdDdYZOQvHe6Yogsj/WX8vrDH3d7Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="X7kd5PyvBnBt6Nkq4cVoE5DCdYkB0gt+XeZh69Ny8/4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
HTwLS1vu0B6O60ogX9M2u1dNkOFNhPMrDzLuhbR3XlCimILV40dzZPPa9/6wpiraIeBKBDITA83w
7EJzat75Spx/8iBg7OxpbM0jjS7iQSChYN6Z1LHDphgWLb+VgMFC13hO1viJmau0pKEs7Nb7YzAb
8OiuHAFlg8g3yr8WJVYP9m+n93wRKLks6P0jNY2vLmaAizBe0LY64cPBLeuW6fczi/CmN7F2Vhw1
cXaV6FhDdrmQn6hmABaU7QgJDvpMg4iNCBDIWKNl8nHTaCNGAaPVkmVybkA+HRvepafVrumzfA7c
6K9HOYu/A6z3aT4yrvJOAMDpyPPGn0X6wweANQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="wTtHmFSjF5vY4dkUCxQLoBWuMf3tzSI/GpbZ/qNzKXU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9440)
`protect data_block
sE78scq176JoOM/H2owdJfg6z/r2+LmMiGpCNtC6iHIDjY1t/JQLfH/MZpu0uvxeLI3JhD/xofQi
y1wte3R5qMwajNlil9WyYsc/6db7rqPevXhQ6EXUuAXnz7U+eVbNYZIhFssVNqjjisxDThR5Kvr9
T3Awm3ZSdvytQYC5vf4DqLNwjdhn9iTnJwXkIthLVe/oUaRw7rT5nPuB8DGaCGirt1ZgmTOi7PKY
NtMtei1psr0vThTsa6iGSWlKzW/WI9Amq1TOfZVDqKuVW8dK9TVMNzFmG0iUBpRoIzbkAHz1Aioe
oMN9srQIeNHSH+2opRcN32vV9VBACAbpqDgohQTE3jUVsg3HeNWaHqSiGbEMFs/EMYFrOyHbRWr/
BuN07/l/Y7ZE8hj8WVQatak2LgYa3+ungNMIQlqWS/tLvKxH3xpMSq7qbexCwtdY6Xi7OQt2dGeT
o1HktkCHCiAPFb+WvB4cCiFeBvKSwjOa55qQLWWnJt7Az6xYcSNEGIvnUoVZPsTWKmVT/EeYZAmv
/sl+6WHI/K35h2caFK4QYbU6fxKXwb/81TlCH0oNaaFaNdRRItqYT77E0Q0JOszJjbCyQ4Y7WbOy
yuP4lSGOkeq5/gQbbjtmc/uwEidoEy/NQmAl2xIYnMH4JKFxhqsxaKFhV6PUI6bgSFvfwxam5tYC
8WdJkNnHZ8Yz943tiu6vD/dvf0tDIvDEKDowqupsTzTq1vrWZ+fEAoKhluA0LibDoORLzw0yl/0S
To91qmVFUOO3dGD8u5ROyLVBSkiDWD5LeO0NlrdJKiFC67N8MuG7e4ZKFLURi08+qNj3KO4JTgR1
dM4qxmONGA79+FGIV+Rpsy9/tCr5IryTTWhKhZD9EW+S0fa74VnftBjEHttUmfOKOd84vwLo6Ihk
VJKGos4W8L7zskF1Z5Qw1c661FlxyCfSRfmirg8rYFAopEbxlymEY+TedXpcXYgVpIKG5OB378OK
173FjrbEOdKSODJtx0hRpAuFAx8qz59Hm/Q3hOCaDDb04bm70aYK68lhe9SltZOiZRBZoFYEACi5
b+vUA/HcsD/xBKmQb7ESTeUdrVzCyOzm8Xrs357I4B8b4aCnW7fm5n6j370UwHgqBRwD8/MGPvMJ
6vdxd0dRqtSb9Xv/RHu+Y0LSxz8q4xajkNVFdkJleyhKPPcfywKqGAh9A00V6vrUKKj9CY+bzHBu
X5UyrFOnXMMA8OlrG4WquEV7pc+5d8EmZKwsano8Lwy6kQiNptGpgJO7CJ8h0j8RyBx9FE8bgyKq
WAZDJqWxHnz3pNnh2xZRTu+9POevffeBn+F9AAon1XLLEdKZA0WMGG3SfYK8+LDamtM2WXLZ2K1Q
/Qz+4aI5iDEeku3VdCwnH0B0HepQC+oGjSN/unM31cb0eovCey35fdIEBQDS/QFwbcvINxH9Wtcz
oq+ktwLUUAygQqHlc7I0B3N059Mj1gikZFyBsWssNO5IURB2pL94vbKYVFjfYtOboEref74RVuhd
1Hcmsed1idZBj8AXqF3r5FqbXObH17YHFFWQoSxXLaXzxKUujStjsRXqg3Rrl5igAjOpixgq+Dt1
z3GxoW70ipapWVgykoPvKLnCRN8urAQ14Dix4X2RhP3iR1Vfm32+IRFRxR7vvlXFPD6tedNVQYp/
jO1QJUBknwTLgycVd6zC0ntHp+un68LETpcuuEl1PgSAa/d7Wh2e28J0PQvTfSTjNU+DphV0y2BR
mZd8+ujweTG/IRBIE1D3sm59RGnkUwK2NR6MPG+q8IYmjsog2G4qokcuXrPRrWxuqHogH4VaeSaU
JDte04IiBiLNZzVKFD61aGjcjlJuU+idLvB6Ql2ZXQXfoDr3u7N6DQhj5qFBMb0sl2qNw4dqNul0
135qIfoApbCnNe+necWG8HMncgQaS19k34N59LLtQjPpxQZ1rqBNH/5pDqnQThgS85R8MOAS9lc6
/AuH7oZ+HG8e+qDYxWRjw8cobGiNdqaXVQ40jDw6+H01LeaPzlrPArOdu3/XR6XcROsX6cxat3HP
GzzVGWR5+PSgqcAvUg6IVuZDUnyjPoMg62MiY5AQpWJbIPPw0j0bRREdpl/O8N8gqS8lOU8aFtF/
KTbTc4LXAiy3WW1Pib0jrLf7Dea1DrKBV6xhiOG/EULL1Bj9TaPIgb+3kGfqageqIEcN1eBXBCjX
6LjYdF5aZ3UwkGDP/vjU3HCeSmcaJCLzkCDnj0RhUqnXmdRlBmll8SShgmEOdwq9ibpVBMb6nAes
MKiXRES3+8QkYLob7xlL0vzqLUG3IizeiOdKMrFX8690gg1dJpAI1ra+jIRSZo0+Y0itWFV+D/UJ
mRwQHt6sCxY3nftmEtCeSAmBAnkwT0GKtUcb/61EFqdW3g87r30Ia3RKLFtCqZ0U0bb6MClQAXKs
R/0JeJpObGMps6DcX0I3x6yOQ5NIOJEUi8Rcm6eCv5Akf3sQ6GYAK0mA7cEgw0eWMOLkrhT69wiK
synbApbmCm6AJW/Gwm7QvoC3WplGM63mICjzIp1vUH/j2A61nG320jGni56mz7w/zf8t5Jf5UcL6
ktDzi9jDVY8YEhFWnB2oacW4s60sPTdYDStCLZIgH2bCerYZ3XArFkvvQ8zSTGNNu7nc7FhZfr8b
p9ZtDhsMpSlxqnfBqV6tyMb2WwmIkHy38DUPEAjvYDFG0eNQdTM+DIvXgXVUMYViLgikFJIIXPNp
EuXITd1V7mx3B8tYjMbDXQrKl2Ez94iTZVV7WTH7smxigtLW8fMPOW6O9S4wKZZ9MA3L0+79tWFv
keWvkcUbnVK35GyAZrMeYj8SurKSc7DrZ+GkPNsk8JiO4gZ1HWXGUIGokLYFyPn97pP072GZB7iQ
ITlUNx7g2wNolB7s8505a8suJ4oqfG+gc/PfY0m493vp2u2FkzispkvZ7SwfszmqoQTQVRj7EbwH
mV1UpwkQSuIfhilPnin154YElzZ56yXVGTIreOn4WcbL/QXj0cyI6sBHq8VuBcFRqgPZSzfWHSEA
Iv6vFaCJCu3hkNYV6qNMeJwe08U3IiGSLOq2wKv4XfErZoSMX6jqJuxiWMCgH0M1Bs87wMVNRwgm
1RtN39mcwNgtupkIxfxwnsBEAvE8ZZnnVrfl00qXruU6bX/mP9otqxrTe1gtaj3Fvww9SeC7fcgz
KPCS/gScuDRSrWXvAZxHIpt57yG0lJlSt4nkMHGMowotmKU12TibQ5zY/d9flj0RHdCe/GiK2zCK
DVs9KzmO2SjvFeB38g6zCtnE6sh2CvhbEywzlGsMAVKfnjoPs64XmUbrNH65w7uTaSFZJXpOQMn6
6IhiPxCGvM1v1Y4VmZ+Cjgbvq+M0R2BKjbgfC89hozeZtq4VxDBTNTuRWkp9Po/YxxwBFefiaQYC
Vqzkel9gKrJmU0yolG8S/33euqy0PyOZ52re5OOW9pZZTJJDVTQPEnirj9zuxuze5BvtaAEs7dfp
P6MyRVbTf7mtBbk1QfJK+Fic+pvSuvwLpShtMyHUn6ED+LKwcgSZBU5A6j/fwts1cEH4RJJ4Hgp8
hiNcmuWSoccx40t1SpCIqfbq0Or02ozTJKWwqyOBGXCHYhGrsbhqPuIZiC8UENLPNGOBvzmzMQD7
vDb8gH7lfJ2cV4cJ67qk8Nwcp7UEDlDg9wqRd6+7oWt+o1nfpAxGiLq5tvo9yQQSsGuRqwe/dKMo
2RkhmzendcH7/QSepMrm0AtNHTMn/L7ztBbbBSD/hD0iQOYgp1jQcrGBB8C+pTs5dCWUWE0AinUR
eHV2w2VWbU4rASU2Jx3rf54tZd7Jfgg2yfiUMPq5WqBiRRyNvcJbpM2KB85W9J33mKqmQFetXV2K
vMOLF5ZLAuafpLlFAq0aT9d9uvb6gdDve8M13/tLdVN1VJsk58ArGTMVb7fTlou+zZWO7nJ1Gup5
WZk9V1VL4sAELIQ38+6qdAER4WlyaW5syjFCysoxWwJCC4fuXPHQ0rZkWsqsph+GN/zIX5Sjqf3/
x3wK7RJ7BFUdO3AKi/Au08d6ACzcjeXTEHO18M9s6Botxa7z54yAZr8H5a7TXFAOJaKUiX1faUEG
bkrh1goP7VNI7zSafKfebo8y2m/tJgeXN89MqSimTPjMVKlKQucymUHcQIBMchAOvJyvLU1ic+1p
ID7hx9yRc5942kLBNb30LIn9rH5M/KMwlCA3ExPgQXHX9rXsLK5kfi0eGPzmUDt0OkZ2c2OtWksX
Lnc/T0peT8HJEf6dqawGl5OGIAkbLqzqXYiHM03dGU9nZ3McbKqGbLr3DheHKRD54klLPYtmFaN9
eIJYveSYfFGrDFEiIw5znWBYZmEaT2dFO9KBnIhHE8jN3wfKL8cN9tNMh5pVn6EkGbqIKa5jMh8W
ug9bOAk3HhmvOw1Q2etPy/82oPdkFp2CSXh3MmoW+HwMzU4NljU+/CtUYzi65t/EFYxX9QCeaOTh
KbWoQ2K3TSrQATlCwWxL6/GL1OY4vhUkOZV0I8jje1LYv9VhThl0TdsPViSx7vdonNBqCAfVxB4W
9dRAUAyPgV1KUzqVnrPXeSGDrOxFdXc1/2IutNhyLJmXMzb3ry+iPfXZOGWHNsJB6LQtxHkQZpDS
AX1695rhKJrgjb2ikAmcpG6itXfP1tJAnMbjDVeBtj06YgNer2iaPmm7Z5NCTJM15jx0lWA8MZaS
o1xn1xPQ3vSdz46k8bdt2YP/z3WKzGvqmy7ja88C0YY2Rev7Bz2KMn62m3C9ZvcN49Wk2/VOJLIP
qg5Vw/tYCtcaQbwbUPH/QS+P15wa7LXXMgA51CZLztKspyqwT5T1xwZwaLZhq8LiYu1RH8zUIjyr
Bg9lmlEQ+QBmxFtjShEt7jQoIbF2oCfPdewfT3oa4KCTWGk/wTkMLFfKNaDxWAPAyu4xTQSepjML
Yhm/KbX7vbmg3dMSxFU1tBYvacMHMaJdBUyw4rFgEZdUpzPfroP4HAZRC7bq4zLjCEuRfBJ1ei67
HlFNj3QZVDmbVSBFVi6XMArpozQEI/Ur0r1zj0Ui02srjcratH5yFKGeOtD0cisOKyjWZ4UFZNfi
ZOFzX7HCrJWTeaH3wDTwsFmDIB+v+eyqNKoF6w7cvVJl2Jyumn9oHoqGR6AjgmRVNeI05edUH3VE
9eXe5+z2WCXV2P4SZ+DW2gNDBIz/Fq5BQTz/WKPopw8MuzHBb/c+XCo7cKorIUcHtgBSGmtDCoA3
PsfjgcXl/UWZkdmhS+N7hS2i6tv7C8Jjw8XxnlJtgb/4LuQFQDkOnqszYW1wAQ2zzwjuvp1a3Fcy
F2LTW9ouAI3HCPRwJM9VsoZkCgCoQIMl6HcdM8rEUHbgNqKX4Km9A/r8cjihGSRrcDfRrv1Vf0YX
7u4Ke0DGAWRNjdZ9EgZ9o/wEIhqFrMwEzXbptEuGc+vjAL/jRivCodrQgHdd8fMln1hdzreofS2c
xG2OFN9n7IXLYsrqL9J/RcnbnAIZLwQgITScTCe8DXUt/kVlzTQqiXqDLLLZaBPoZKwZw7oD8aY4
XCX194G4LnpZgakgBEVMvrl0axJPGbUrTcRfAyyQx0uShg1Q1dAlOorkYQ/fjp64rgF1Sl9LKslp
LhBTDsSZES0PvBb/Hg4n3BWTn9S1gPIyPyN4EZ5FDheOzoanrlcTDCvh1vYDSyDzd1jYQjztj3Iw
Z6x+I3ogOgV9O+QuZzXHfiCsYtECFwp4+UnroAXwnRgxhw0T1qoHAgnvp9qn1EizwPcapy5IM/At
xlKjxW/3OQjZVNjWtLM6e8fpY+167GdGoUiqg2DCjPViP2Io4l0z2MeKkR1Kcxfl5VkU3X10Ct7R
2WPV9rj7fTgrEFSNnWcSWhNQSiCwj5XruUs89AdFlyOZukfRH6C7p87fsLaUZ0vT390kaTB3FhJ9
VOUMUepltPP09TjWmlPutJkYIQZ1+b8SmhqVlNHUtt3cR9uVrnjX3J0H8yMJBW0kNVVqVkmoiM8F
dREH3g+QfMMSfOM1KgSJfdFrIAVYA6ru/GOWePv4UNdytOLgUgc6SzTcdpUWOL8ffydHTSQL9uoQ
YxZ7GNW7oYuzFMbYv7T4I94thJGdZl8tCqUdmU8Xuzq/t5AQ9bcEyfxcSQBkNuGu/WcgeEqcPM9E
9rxWcrwyMf8dA3f2ohTXh08O6xHaT58LIU+iPY91U8W4l1gLiM999JY7aHbdl+fIRGdy/0NesiXC
ONIb1WlqLQdraQkds4gN0ZfOd359CxEcCLVRgMRBX6CaEHOx/Pqh/thejBdJyl+8sqGVar0FJVHf
AttbPtr+DK+TkDe/5bkIvtbx6L6ITM3WhwNbjxsnBcUZkXXthVQm0fbTnvfmyqf6Ml6PRi46jxfc
FF/0b5AJs8de7b5XBJ651ZPAHGDxmUDpVLuCaptJvPLiHiz92VIHf5iJ9Xk+SdbAood48X9AEwcJ
s1ssE6Fmd/14L611jY8BElpFHyHtAsIFpOqAuveuJErEdRGa4X0d1Y+ymVd6VsbkROfzIuqpQNS2
cPCCx6OQgEfJf7H5NdRWiyKgAKbqC8ZwOtuP1O+bmao1xmAmtxQIyXas6/2s6gw4VfaJvknlVtX4
IMbaZOGMN0J25oPV0Onbki3lhZ1T6ASW/UChVOkzhGdkkfNELoeoLkHEz5cruR7fe0DlPGlKt73M
jFmAluf71kudDzQZXtRH1m+KnwRqvwhGXkNcuu0GLD+12Y659P1AAkBpn6YDSW/+JBBneHA0GrjO
tZU8KFFXm0EOeKeIsi3v75vLq5uhPXsLIDJBJpfXIr9kisOHu/zrYbAyJK4VrsahlLUh98yGx8wr
jUBVxE/zeAeWO6nNk6C5bAREYzhkDogfzLGWE1hcXorYLXg5I+Exxlmi8Qpd9EUdo4jui6aAF+9P
LOhCZAszLdm4/KcTLoU18dyZJ05EBkWpxIDDQVUYv0OfQzLe1leky1s5WgR2DfGSestAOEqUT2tu
HB8EAYyYoFoei4FjDIorn4OCZy5jJ5+sR4CvwLJ7RufXaAIeg/z5TCF5L5tuA74vSEQmYqxTzSwP
btzpZjzr8QRqKIpxyU4o6qZxaSbkf22BQMnJ5EumGLO6YGwCHZHzzGNy72W1NJMDs5FI+cNrj0bO
ObtclMHDWC7HHwPdTRIkaYmDrzfkajfwEEE8FPForLULxPT9vIxOYrsMksWVpRD1/QeRQcsWw8Mv
j/rvFffmELrzSEq9QNgXsIR9U1o1pOpGrfwRZYJ4/ZJsyDRtYCF8xxfH+j76YZ5BR00Tzd5fLxMn
u4eqVumzkxjLBORJd+fIOQlvv/4C8dqWondz0Klh8O8QHzfwUFOZ5ZCEdP2mBgAuNF+SpYq48gu9
QXq4K8uIk0KOgmVKAJG2WtduiUK1B/n8Aada4RLvfZC8K64THr1PrIBGnHHcTMT+0k25gMsuaepF
22cpl4JmxsDpIavcYGkzp/+2Xm285Y1fGB/akvDFG2uiHw6Khhwpljs7cL6NSZPJ+FMo93bG4NP4
5yViriatQ5/HCBgwkeScWKT95/gBsA9Txn8E+RFhG8lYgNaXEGxSXOyqgQ1OBBibK8Xg0pUpEKfN
n7H0H4bq2n4RZEHlG4W17DOPJo6Lmif15tzwHspi3TUaEy7M/5UO/KLJMGsw0v8awezAdrsyt0Gj
FsuI23kYKxOSl+qhithtfHwyJi6xdXjwWFk2uHqg1AkVqBuNdLWiJ0m0R2J2wye8/UnT1xD0C4r5
54SK+EuUInm7HsZwgb+rJB5DShjZPU3dJNr3b7fTEFwj9jf6sf4JHU4inNburw90tR6leXpG2wCZ
n+h8LXoj/2hnFZYFagkUWlgShZDEtyUEnfoKyiqeYZPlZybFtpHlMOI5JhhBTy2hVVER8ycrUYE/
xcztgnOlJ0HWSL4P5F+tIJ6GJiaPO1xvJn3faTnqwwoNUrI6gh7k8jpXe6ilJNfCbxtlDfUGeIEZ
0qgpQMeFd1ya/B837ZdAXRoL3w9BOaAQXZnkKs00Sz4A9xgFsGdYcbehcvBo0XvB/og4nlIN7anw
djst+Nga8PeGftDJf/WWJeIinZ0higLwEXeP2zJq1KVEQj2SWpeD8pFdzWlKeeDsShf9KzKtFnKn
TqtInLg1dGWryneXYdqyEyyfzNqvqNSgbv1LOwrTBKeLH5EJzFR0itvZl56qU6TPwmiL0i44k9Z4
oces82ejSSmXnPXKbcVsy343GwFyvlVlTvtPgqyVbGwBn3eO4uYoI2ktSsTfHYrnp/G6SwsM3qx2
9P8V62Dsyz21l4NN/bs7Xlb5ff4NDTyKK/KUNUyI606mfu1XZJQ/Skj6ZmzvzCDzHGsLRlv2Djm3
Xnqeo69QcKBdnoLTF8PQTxGyqgSrpKE2K4oZAmqEZ/KNWzs1wlo3VMqICirDQ53W7yC9/oLG1o8Y
CjTUP++jdY2NwN3zuY/XnRsSi2rPAI5iLVt+fkj/2AEhQZUFihB5ES8iSg6nZByJkmQAN1MXKQwf
TrOcJXv/SVdvFRQAT7uRgiaz3Fg8wpohcpvjFzsi7U102dhsSPdJkG7sGg7pW9HBMB5S1KF5cMiL
b8LjkKGH49jJRBYm81ZeM/dD43SM8reUNRdw/jN1mSxDYdUwAPVx7lW9uivheC4pbl0vtoaCLBcb
IB+sjrXTJbHDI2SNJF6rMF30omUdbObl3pvbv4ZS4HKzo0ATywGE8NB41vyMhCFVIerF3Riizy8X
WKj+xyewMH6RVd9A0FLTEPkgQ7SgznBxHyTMDT4B1vAM+pcw/r/07C23hw5aSgKzngaPbqA45xgA
GAo8UOM4M0HkebnJIslMUqf1ZuZUS1g4uvPkPqxhwMIJlT8SHD+rakLCY2FL53/fLW7W4VCV7oqi
Xq95R0FvaBj+pp1YWaHQ/9/NGaZoLYgWc+vGSlu8wOFl6WIw7aylTZ6BWrdqXL4+XL2sGX6hogfj
m8sgRhSl1DP/trcwxcmhEvYvkjg4JdCtake/yqFSlm7EI7RUnVCL2jGuv6a++MgjCcphOsX+1FBB
hNtjwjJgxV0TFiM50PdXxNujaskTgaCcVdWEnPFtka6iv+41aimcHkLwmx5uXBvLUHJhY0aRjVCm
UEkBVtx3jKUpaRRzTDYEMDxtGtMTUvQ+JR0k0jJJsmAQJ4cfqnAU9OyG8TGJnb0RQFiWIXvZ2/r4
YJj4OZDPmgRm68YF2/pTjAjAGwY8mVBN/+pTTt/Ktmw4jkwtFORtoc9L22kfPHA01hknFRNxbQd6
Ip4Z8HpxOaXK1HTHWsupWoVCNkiIAgQ+NZJ9Hj1mkMLLkd/wnaUotX2jyOSMF5qRgbd7EGPmPlzj
OXwrBCWGGoLav0gcWQTksdYoBylii0J1WrAz0NG/zeBz4Mgyc7WRMJhN6wM7LY6FENxmPw+JpXQE
QLVReYTj9NW39JeN2hf+751J8+I4VBBaEM2GX5qoQ8CAADo5nMltVjqoG4yCcw7n2SUBs9sCyBTF
J8YKPtjgbBARVk8PF1xlmRArbGggT+gO6JAfzxpWsGUf+u+AgW7mRdFBCoDL0f/jhXC845fPxKKr
7CWJVIjKQIfi3tTrV292+yu5Lu99Qff9Ay1YDu0rLvVaY0XOc/Q6eFIx64eEhruNJzix4GZm+fwP
AgWA9dwtcyAZJda53bnpFqSDM7wl5fzY+x/4pC5I2qYBc0Lo8mhzgcdi6Hds6GXzcKkX5q7GWKwW
gN4Og/J6sSCKEceWocPQkMFo8IEz9WGl59T5rAQBmFsDQuxV6J2e0tdJYizYnHOjF17VYWR34Q6Z
Z2KQ+oNOz/VWS25KgEp4ujM1/cEUJDoCg9cY8PIKVulJtG9rMi5Mgf8uowtIvZqQRTyaqtuWg/TL
J95T8TS1BqzKOaK7oC8D86wfrcnylM8HboUzXndz8W7FrDEV7l73YakjMwCEN8hZKeW7xQijlHCe
sdat6drD4tuMpWsRTU0lsYFmn4tQC9ub7BTSZcWoH/BuihqEc+9gXZ/96B7dt0tWO9jd7GHOuUNj
QbAzp8rXMVA1le4LQ16eiS8kjMEeEpFFjNr0JRWPRWaX60VPjFAqhOoRj1UiCJuhpyNR/CqWXGSt
UqJn21TkUrkKy6LqZOhr0DACTrJ77pNWeK0G8lWgJhIwD4By7JKhO9EbbV1txc7ionGVZnspttBj
JlntQrYUT1LnU2OTkpbA6KDvdzwOjq7Ya8EaleQs5mT6BghWTRN2goJjsR0gxjwNvsI63YExjrHC
TbAV1JhnkRDNBXAw3CGDhmJL7ypCdyJWAuC9dPZK0psj2sw0DaHZZt2IUwmPZa5V2sOekTwUfvNJ
runKNTOrKhZPElQ6yzW18AHMdtzyloyJ6zwYirH+F/qronuDlulhvYkGApAENbeZ2ooyRJufxz4A
/xBazB9V/IrTk3c6KlJTrnOF+ZHb5dzYfVERhVRyRV2hxNKd2YZzCyIDAtojdcI0g276qm/xKN9P
wccgz0D5FFB1ljk1gVREqF8Ijkt/57HK2q5Hax80fmI7VjB6ZjOGcmkw9MWuQAVyx13qAiwvmIKM
STQjo8tpPTRuHMOL9CwfdQNMqdoRzAiMDvNxSSvNAaSSgNcQ2fp7UIjHMRpm/tdKUqpqZrPpsAQf
40CEFlwOoIxz3aPgA5Y1fcCaUzn6ae9lDPJ0f+qfVoNxJ7FXHkkdk3FpDcnvGaWcWs4H5yVXHVqf
lT719JnU30kqe0H64xc79wOztZSLUIAJEX8gZ9aEmvt2DIxhEtCtzkzYOeg/sCoPxEi7QF0iest7
LP6JR84sXG3fL8NH/cN/zKEadYURFM012z0gGlSx8cCpM+2KHl0Ne6zRa83b+989vcBrypyQvCtb
O6MmmoBJcy5nUSEmjKK+MiN2JCH/D+WAElFStB5Hn62eX30UBpDNqvrzRBxy1XrY7zJfzd7c8+QF
zEwUq9fI5gnjUrBAXgaBrd1uMiH4/D0gEkdybj+VUX7Lso7AYNpCRAGK4ay8UOratTzWdskmx2mD
zaxrllVyzn8AHswwGaucFTF3PQORozLXYokrZLXJ+yDxC/u+L6eqwy6jDO++DQoUZjfZH6nGXovv
lGZJ8zsHwy9wSIWdRwTThJThnCs3otQDXBvIbXUaB4vYBSaigo9Ad4GvWsgEECGANbXFSzd7D8yK
iVl2lw+7m0x9uUumY8nc/ATh34hSUCUxdHF/uT9vUQwB7cI1y4dvJrAJ3C+GtTGtVr4TKq2VXiP9
+nBa18LjozTRRsw2bLZF/tQo4bj4MVNAVv7uJvULsgO2Ap8EZg2wFeBrGYVCekTUJv604DLTT7P3
/J1NHXvZPcfYPJici5JXug2Vr+S7VDXoQQLBOFq5S68il9GbgzasAGC3zE2UCCoI9LoUOviNEy+p
qbmj/RQTlmBBtjITNNM3s1VOnGO2CV6KDXw4Lrx3KGYWecFMz3e/LyQzEW6lmsPRQT1y1dRv9GTb
QOmFkMH8wcYGORmaL/WCobyY/v3Iv/h1zJ2eTm6Etr0MlbWYsNgh4v4ZdgDWUDGt3gR/objOvE3E
amPTzVHZqNhE96p6hp6RU2DVu/uiH5G8CBogqmNlTKfzd7hU3APH8kruHDfr/Vkb9/CdMgsGJKo6
u9/szfmjUtB4nZ2uxYy6de2T1GC5nE/bq9Xc50A4ez262Wacuw71GVEsI8h+DPs+f8ow0Nl18jKQ
csu0QqTZzEXRdTW4KfxTU7exzBNwdMApIec8yK8WG8l903kx7EJy23zzISDRyxpt2UMMzHRhA1zn
l7PsSHXOCBfGi930F1hKi7+asu7OEFsZd/+LNwRxkw6/Fpn4Me19ds9dr4G6wGWLCxnQCfUdfCYo
ZCFMXsWN4/kgqgx0id+H/ExrR9htiu4QkjEfFUZAoFD3pTzby+MX9BpcJ4j3BYpZYRjpMLDmwQfM
LosXAE4LBDqdu9lTOLwVFEMio68ve6nO3fHjWQTb+AyGHQMVoHq01aK8rqw80bKrVfD7BqQ5IGy9
tuPorl/By06aCN/MH90spFOB1DHpzf63WeFepLxoBbiWLbHpZc0RDJ17P0XcRMWdpk4F5TiedLd8
AyxMDV5QDenb4ce3uH1XTZleqMacz8MW6SdmR6OesoPV2IQyH/ho4QimRgW0vhbyyqDPsvxJCoLj
UhMTBTBVb/GhMhvK6rlUgpmMYMjhqtbZiY3SK7GI2S3irbQt3E/9cD8D8vUlhLfwV/pALOf5B4Po
KKQX8uMWKme/tj3cs7DWBL7er8bX4jor6JlayuIL2RKgF7cULPr0mOZfzApUoFYvG2CacVroN1bs
qwfMIVs59bQwYgytZsuZKgDHE7vkqj1FSJWtBxyati1Zn+n0r6czF0OyVbOKZRiVDpWpv8fCU1hX
hOuv4XJ0uKTTmOjASfKeFyLUTzm4me+Ghtt6aUt2OWcfyB9ipPaCnRLG/gqRMOf0a8ocOMoYGyu9
DasVsjonvW1u2nQStkvfclnQscUNtHc5Il5CCzHyoLpUjb9gym3zEuipceghm9YEKcjiDTpmhVRY
WHRQnc+zu89viZemSsORQAdNbCF928TgnpdbhHwASIuEFJo=
`protect end_protected
