--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
X42R5LIXE7tx407jYzDVCHvc8BFgDqQYc1AYVG9eHk75RJ1AOfTbU78Caoe4jsn1ZdQRmUFkmfD/
S7EtExl3NMMSJ7b1XwWP6xco5MzY187lbkE8wgBKs/oK42c9pdSiBpkr/VwwusUq8KrZDeWs4t4p
TttQWTcpkKDlyqd7uWanZSOwDEVW5sIJn4iS1cZogITpGKZbT9Pi+RyO9j8vyL0G9+oVeVZZFuD7
2OXNktAKE4Wc6FnsW7e8ATVMAo4GpyF+j48RrSOMYiemkLmM5CX2/1EaoG9PdT5ecmslku87G9KI
TiSxsJsUTUnHtPWiCwYjJS5jYU+yYUd6ambAtA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="VFsZcW4vz9u3JRr60IiIco0pGR71ZQc/VwUMlLIeIA8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
i8G4BonJeQwbk9EFEcp8YwX/OzeJJ4F1jUmi1MEnki1dO+wdH/6ifr3qmT2uOo6XG74jtipwwCym
Mq4nvzv2P4G66/2TBasp1Sj6X7eT8qFDFMe7X/BWQyGBfALsiXQXlj5HGOmY2duFR+ukaGGWkRa4
h2bx6S5iftu3GOPrIChBPO29C7TZViKvNYoH5EiE9hju9Ao1ejqb32pVyteMCgs5/tFCLjAUlpb7
Hh1AZSM1awlIFw6w3xnc+cRaD+3aHSLS+8Lt/3X/G34fVJffS8ypPwb1ePv7ObTE+3XEEfzw9Ezz
NvHnkgApwS1c7Pou54BsGtr8u/uXykYZ1RD4Rw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="dSo/H8oMpbU4eMaTEVX6AjuBzhe7YmTFIBGirg3Qoyc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6704)
`protect data_block
wJWkTtvj4kntPZoIoP9TAgtAwX99iwIR7QMboJn81xDWtlKHPiDyujO74dLbsK0KCPkRFS5a1j30
9OgcQggieHVrmsB3h6+YaUpuB9yI8Z2WumCG9B6lGa7ZKTSNaUq62xBq8//3v0GZEf6dTntM1QsK
aJfUhy/EEEJW2tWrsOvTi1N5mrORjMVN14cYKD2UX93rJa+HdHalznu0HVlPAScvq/CEk+AB3/45
gtThDa9+deiLS2W5tL805SoOvVTTk+V4/+WT4H8qD+Q5UdbedOOBZSBxRjVjWt7MtKl9Ez4dQEWk
e7eB+mSnD30IBhosowMVEn3hW/5Az/10e3XdvLoYvmIlXdZVDYWKIgMcz2j6HJ61fLi3UVtGOH0k
us4lCRRC1cAJCPAdNkskWH9P1z5IrJe4p6KaAFiHbbtOBBI5RgHks9/MFtzxLxeUj0OXB8psKZyB
HFEbvVBZvw9mFNSSzAZWrBxicNX9R+8jXdSU8CW5C31FykrSMp/3LHrfmVVCzMpEih27Ihfkhtv8
o3KAY3lUXN6FKlMYEGELGwC3ixXz1nd6ArFXZ5xj79bFfbkPhcmqMbtMLKWceHs5wZ74VKpbB+8H
cGSAd+Zy3h77Uhz3FiaHi+k51mkGXA0QX5+9wbPNKapRFolEPhPiiekEoXK6niVx5w5nFuz33U8e
7PC+YfX2qWachE9B1As7B4VWM06mXZPH+qZyqJ6f+rcJY31nbC+Vj7oHPyvKAjafYM1FI1rrcPDx
wKiBZbc8+E2CBE5vwAp+nJAB16K2kYSO/9LmnJIbowbEc4AbIUxWSepYOW4m5zaFk88oSxjM5Kxw
ru9ruom/e7YFPPnhSUGEgKd5KYDajg1m4KluUFOGP55fYk8TREDomCWL3t1RV6WcLRGbekvxEv5A
NzGM0A83JgDAgQvjkWonK3rk6tCktnBsGmDqqpE3X4FsVeqtDdNbh5tXhb51nXwOldqDWFO7Raa+
sfVEaDK/dD9pvxU+A9OF9r3Jt5fAmAl44hMRdhE38gqTnRulM3l9Ic8q8cfNwAOvqemIXbT5gMQr
roH7t8NG3IVFNukYte5ZhPc32Tp8EHv5irXzbl83uaintsCjKxhy+QUDPNZRTS90I9ME/Uu4JgJv
i2wS7H04pFF89SO+GILMU7F16Y3o5Ym0vKiNTj8MUlSiD5ZvLFzLLxgOLzIRzb/M73vd36DtFi/Q
dlZe+oFnadqRb1yowmpv4JWrhb3r8TUq3OCiG3B/+a69UiyvJG2q4vNbzAZIOxGT9+S5hYgI5nig
VSoxIx4E4CR0Q2m/kKLgl0yyPKNKJGG+sSSg0CDiWv1+9gWGrgPO6oId4kS+jmSdBNUpxdNz+3WC
s1SuQl+g65JsPtku7L9enqLhbLexTOKAqOKCWVsOrt5pKxuVrtLYHOvM7u2geeUv7UO49QXgAJcL
LpNgglLg/YNsb/DZLcxZQCIN5+m+hjPdWI3Y4HitKLq30XmBIlKWZ7hKFWYs7pmjHG/4HNBnrReY
tyoDMJK9/78N1S1GR0Mpqz/eezq5OEvmDyZxyQYnVDymxutIuwrJ7Pmvg22wKXpg5WyDXybuLKs7
qxd25fzpIKyrW9zpqp/SkSkFPtTn1abHrSR73MIc34mkdjxPywF1YS/oVkeAvNQHajzuafu8Cm4H
ZyIo4WsPNIIb5hc6pvu6BQ5UchxJ2ev3C+OQfoQDdL3wkyp5JiM+GdDh685ZsKeI+sI1aDKKkAaW
JZNmVw/LW48DJujFPToMXyuDYdP2GDHKRnQb/lS0IxpO6AYCU2YEBR3AXl1LCN+AhuMv5x4w4+C3
uhrgINnrs9gSapO0E+Z0Up3erf4RwZz7Y5mCN6Tz+RwxjtcFOPbchIKT2VWlgcnFHrUusDYB+51r
VwzGl26yB0bCocXswjpXcN/fNe7sHKMzNspOWpawsGPtEzACJke0KlEptkwlQSaGy8eCq3Cwy+Ht
I3sBZou1/5iXx3fmbf+snEmxLN8C5dbh1AfRsVfGR4K0s9p8akoSlM5ilJ61KRnNv9XeuzSFWPEr
YdYfJo+u2eIqXYcHxzzMemlSzDSnUck0sAFsvJtn7HQXkhVig2/CflVFdoOmrZ4a+Hoxsy0wPIYK
ZwXXM4uzSS7TCaydo0fiCYvByhzCV53/rkfMJ2J1QPrv6jxXE3wRCKMdOxI2+zwLy2TQFIIgpDi8
gKWEr7esRRSHgbr+Fsm22UikygwMIpks7GeMJNtNfiMvXhKdi3hr6UMd4uVAvA9U0O8khpW3sl+d
oNTWgNPoP5S+6Km9J276jIPwkMOxWHUt0dMTwpEvzsCRwP+KH6vO3rzcasApjYjiQPRJen68jlkg
tTg2SYYZQ108k/zE5tnakWiMafoJbpYhQSIYebJXGz9mh4zowqlU4nEEjBihWxwv0/X1k2X2E1ud
fiihkmfUVocHbU+WMdOO5zW82o9jFEb4v/8A2z8vkVqzb4y/SRfZ0pEHM0SIFoKXFhmY/zEEWMql
VddGjXH+1MxXmpq+F6eGpV/hCg5zPAo4Njw8m5dAqM9Znie1B6lM0oPFddK0mk8M+yMadMIlls1b
9yIr7y2W8mea5UnKOfagN+CwPGIkpRaKJ6QyCD1si96SwfqGpWVX+sBWhI/4lRDHQiLwWFijnjnH
XdzNedyHk2hV7mPyQTxP0kwnlWWVADQz25HhJawqXz8cUvR0/w24WVUpfol8xWQfTHSxo5oivYim
geQqRlo+KJ4L1ENJDQpstB7tXJ5nIDCP50JSCkeLiPTq8Q0N4vhymILmmn4aJm2DBHiGBFuk/kCi
LN8XkBZg7aqsEDUnUaZLD1o5ZEZnU36o0xNaGRBCB9fxLUMW/Si3ozfU73dXRtB+UKLIynVayWZQ
FfIIGLICgwBtP5z+1472dLnzSoIrFWUJjp3NIthyuE5wUTv7DBmzsw/ZFPdUWcJ9zQjiwB8hWqz3
XRmNa8EnEIkt8QpNhFThGskU8YdJU7dmDp5XcRSj9RUgeozCbCDF7FI9lmaD+Y2IWKxZyDVOi3Vg
qiQxB5pTJTpGx0GiLZy9+UhIfitcZgFNhjMQidiHgH7aS0gDOwJI/yA1YBABILi2VmJ4s3fJ0aKv
sD9xlibpiuBtW9LUTzlY4e6uhyp7VvDNwgWFUxfpulpU3jvwqKvfdtjGM5Mr0SEwQcaY2V5S1r8k
OyHN09syzwkZ+IuJDAEc4r9HgN35oZW050lgadNkqgkqHThx2Hu+TLgrpGvtMWUXO8oRYIXiCZhV
k+XGNaYQ39kvE1VaKgV/Tu8rVCsdkrdcj06rJIbwTpMEECoxbQdlsHY0VF5Vqs2dinMsiur6D0UP
QA2vzfS38vUJgD8Pk53XKsrrP8fAKVujhJjW1De6yI0hxORd82DQstQ1mJ2+zCWfEPE51nuDqRDo
jnicnwf8FTBOnWmQAxF1v0RTy17YunAoH+4KfGtVW+j4Wv/B6IzOYTOVsClMPlkN9jGje6t8ckkM
q3+5UnPOGNLQ94TRRYC8jkKu7OruzCMULiBgGbcdAF0JPCe4I0M68KiFtCqGevvUbTfWggqVkAqQ
7bbP7AmZGzY831ZF7DpIO47tH/iJa7yV36mYBy8+P0j99EIZAAimNo4BRUhkPjs5nBjAZotxqKxx
d9O8NOT0q1MN3WJS6kCarA80EFPZDccGaK4LMApOxPvOK/vReqg2/+YyVmhDtoe5DSuzYH7HYDOK
vBxSRvYMDnU1amIXftR+86SXtBWWJjvqiDs87wYS5QoHi1lzs25S/pVTMojyZQTGwRg08QE60VtS
EkM9djr1mBmz5V8IwmjHXywglKujSWeLXQHn9tW5VcKs11jw0q1ET/sAVXrdVGuf9T1oTPh7mcRS
+neYf7qOJ7wl+MruoZ3kJkA3Rz6EweDDjYSse6suAkm+Wvo/epQYIaOVivpevC4Ve/RKUsvbEp/X
GJAX+zZRkRfijMzmBB4eim2NTEcKEKL8ZK/Y3f0e/hkj+VL5egdlQLvuhgcWigMshQlaH+0o6w8l
Gf5QZh+LfzxplaTg2c0fgNMuL3rcX7fdzRR22zZDIfD3gboPfps7kOvn031FVSBfkDM6GmjaTFHK
1U3fMtivNDTI4kfhdky9AhahdrXPzJVm92HRlZsQbdguZMLMAiFNZW2lY0RAV4WeYWt9BLpTrj94
J/uF+aM1+Jskcjgyi85wmsG29ntvSQpL/4CsovODyCqcpvTj4W6gxHNZkmnG+LK6+cek/PqXaZGe
W9brKW6D+hTxnFGh7AhBBYj0NOyoxDg89tqKHN52KTr4NVg9yj8CFZfE/p0mQv80N+bwAqOlyRTc
Yym5oH4QU9pjZwMqjh4ed+aU3Ck2uz0fi+r5XTgGBWKrIhkUYGn2HBsMRTm6Fgfl+V+uZnIY4u4b
uJJbedg28kpzVnyrkcvAg22lTpkdmPCrM8iclVW/1n5BUBqfXUNK7TuhCzHnDyV4lbN19dCr+hVS
OsiSjxHpigL1GU1pDsKDmngdRCz4jZpKnx7lm867RPUNQsfAjz7nb+t5LGxmwBt/ogMXi9/2kaBa
JiByhNI9ZuWPv6AJLlhIA4u197qRN5V//ewmRVCGVDtYDS+AX4zw1S6eFEi462GxaKX36ETnx0ey
51S90OPsI79AKvWBjOtrkY+JDBDakwJVPclk/O/D/FCnJHUKrMPkkbWCrj5gELykVD/7mxsFATp6
0aKgiIkYRu4xpAAC6PAerW6rA7GDIXlLVHz0G6rvBeiNwUBt8ef6XqgGEgy53Dz3q7n2us+FKy3B
qd+4ctkBvez5OBsW1Jq2mfdf/iVAW+7RRhzSRvO+8C4VZ7+4vTpUDXm4MgK9Ywup/VKe+BX7bpYf
RT1n6xgLA9gwPoigmjZQFpthEblfob8EcFvgqrhOTofourUXTZNYngl/Mn3MdzKxdGjisSFTRyKZ
YIM74z2x7nDwBxwIvuSoY+6kFTYLSFL6OHLuuoYxeo7HZtmj48TyhzbHzjk4BMRKSbxLt4ihqLQP
ydXndp+U0FEge5NDRR1BgaACb8XhddTGCpSgT5TGq9sAtBffXaqRahj7hHjK/N3f3TMo+iJVLMGb
rkckNmzs5FCes8/d8gu7Ilm7sNhNdRmXbcIsHSS/ROsb4AdaPw8wJ4KYwkp8lvgVKlHbS0iyVCfR
3KbVH3rodJw8O+tkUHIkoiEsrqzHVHW1bNkImiuMimQz8SCCmE6nD8y7SCzL2jEoRV3o3+5TXPcl
qDHhvfWtCcrGlmMresYNq8IDCOIThaWz8itTfuywcoQ3otXtDdabdraqR7OKoBUhY+aIp0NCtDpz
cMbTzUg2ed4gByla54zNFjVxt47EgHCQ0d+3fSBR31DiqlOYqDWWaTvFpj4x3+CUKhN1guT5kFrH
QpVI+3ngKcXukDlyqBEt8D5cDboYpPtXgYva3Gmf6tjTtvAwPlIwxU/or4Mj7LLkqYmwMHHiccZi
JmJIXyCzIwEqSseRR22Rh77GYxCWSiPYGUucTchiRKIi7YtMtDUZ5wtBqgkSJ40hWg1wIJFuGljC
bOQSBHB9Ks2+Ypgm7EEx6fh3fjHr7y1Rnv91Dz8oS2LfGrWQb/lG5L1QJvu7JJFfFx3dc4eZZJka
lHXYQIb8Mj0nKQvx4a0TXAoyLetJRmgpNtR+CL2HfE+scLfVG9Aapow5rBXP8meXv4qy+3hMzH/u
eYP/DiAUvqIzsJ1v3U5ivDuqiLdNnxWSFZXKBqIgXv/CZmz/7KdOJn5WUSgFumSw+EblYbSkn14F
rnTCGopzbkydEv98XLFCuTSjsQMSfLPYTeowCs0Go3GdhRcNA+rOLzws/D7X4rfXXor/x3TkUhas
dZpB19fG/XcSQSBYBdKHsyOyQm9v6dgPn5S7gPKCDB9uN5GRFNCCGlNaoSZ3JAB9C6PUVAUdzdJd
0nMeEdgPx1Je7nP1o3gfZiR4f6cgsQV1K5NO5EpPmLsBcLrCqPbLmmEwDLjdAZiW7LjzTUVjgEft
uX38iIU9DexmixHN9tjMQbJVfFk+DBLoiEyWdM+uFxRfhEEYip73fmzziYnZasbGfmyLjDI8atRJ
2ipYBhecv2cbavHQR3Ze4UP8BA0cfvjp0AL/5+lPLTTqNr+4fs6tuCFQZmX+pHhQvmHA4aOv03sP
Bes4iWs64189jaMXFnNBqvzTQEbK9J5wrkyEVuZMfGhIESSyUUEkyHL40UYSmry0zKwOB48IZwA5
8qh9lG6CzmWEmxOHrX3T6UNbIxZ/u75N56osskLwrzezIhA8Gsl+Ic0vb3FcETEAcLKnKua3VenB
//f7dBOtGRZQnzAK4yYp5Dxpd49PTmunfHK49h9EvJbSMI8lwfrfisCORvLnD7WdIamq8KAfpPsQ
7BC7PQJKSn9xpTXKdi4VEG6RRjj731WlxPXGDMIicSwWSopgVl1U0GCswyAyXDh/AMm5nAayOdwH
bLP53cKvtYXDCDYls+UI2QvkxLtUViBIOfxZXMBgea8XPOnd0s4PluMhsYUHqbAnsDSpET9s5uq/
SRiv9Xbpj+eUa66aJjx7D1XwNs8dsdFJSFUArpek2jmlkrT7hOYAOFHv89PPWtEzJGHZ5EnZTvN2
RRRX4z0gWRYUat9BYRnt1vaIVapcKmmPVgi+ADCJ+Q0cSNcXHClJejJXV6yECusBwygHC65JDpdy
qw052rIRqLzXkhmixkGIUaxqjSCD2ynk2YIIpisSOin3WL3pxmy8EDkPhiQ3uvI7b8A27PSQYoC+
MhekZ3KK7b0k1ZvEKDewe3lfd/KiTV7KAj5z4+XzZNMCnk9EMrmPPFFzqHotz1UKFbK6sSWfz8Kx
bYPcRHoeUmO3RmW4eOwStQckpMIupIvTCNzDUgw/f5jHfI9Es2w5H3oDsRmnvGwJldaaeI8A5qhj
Qo1Ktb4Kb9UdofrvlRj1ih/b++YZzqdexFf/5BLVu0ot5xxx2HtdHNN3JZMGc894P3fDzK3V7gsP
wE4iPUwYg8yWvnHD0925CgAuJ2VciUnHOe9chNhG40h4xB97Ku9ErDSPvuY6kw+YC+mHN2gAICv2
BAHHX3cN2jKT2WEXG0j5Ogpd3vVlwDhu8r8SQ2B05ZZE6qGNoqaF2UWnPrwu3F8RDcJ20Ql9GcTu
t3MkDIfazNCslWgSljlgX+OktfKeIvtD2XKlrTbehLoUwOPQDmrbbR4NrqeuDulBmeiTReiTYIfp
5VjzjV2Cq1lZHXFzSTuiCBcr/a9ccx5fIr/YrpZwceoCG0bX7pVZsdTCMx6/dzMLvPaNqcreTkq+
zBVcw5mBSHkVNJXmGahZOyAvcI1TZH+TISokl4dtQTjHCP+v0/BBI5J/Vy4WosDKvpp7YxAHqAzx
6fiCqOmaGAC7H+TQM1MnFqDxzKgiSpE8jTWjmssi+im3YL+H97JlSq+WewFv7f4+2XToFZdWNEZ8
BvnIDitT5TqkgAMEKfU2H7CdT4xX6Op0CXnzyoUbda+gEx0XPxa4vzbwrYYbtYb/Flx84TCeDfWp
xcklp2xBb9VAmyQszKdCp/rJL9t1FUz0oBLOVuOEGhObjksZ/uwxpNkHS79+9HSpoP+ihabyIhQR
GGAQdRBhmrR9m7MuGCc/RLJ+rPs78NXJI88aXHfCX+i0hCvGMZoeJ8vwSTEMPkMo0l2EaZ19iGVg
A+p4PoqcAO2mbrO1V1D3MZceH1BdGxmboUKuEDKtwOJQ1XBd/aNFgfdsg//JAzrc/dmOLA4L/eHk
7xajkKovzt5i3sUxa4F/pQ+iCeRaza2KYaXnxkzZ6IQ9SmJwq0na+ntS0ZgB7soMbR3qD43ppH15
Q0iWUYsQaUonlNNvqqsryxw7FxQKKcXjgzmWb2mK8+39qUbHc5VdyKroSsvGkdWKQnQIHQ6ea+2+
nRO5Rqr+Daaz97OqRhBpfo37pjUzPIvyoQ0PHowH6HJdyKhgNrWCf6jkONnXmq95pD74KTk4F/4E
WYgaEV3ZrHx4t9fZKFWi4I2xu3Q5kCTRrz7qDxNvJ9kkyUBU6hU8y0J/3TkWBQfW+7F+92qQWwDW
jVeJurNqGBerijkDfK98IpkqC7CFsJk4SWaxs7kNsdTkzHtQ3SyOZZ1DVh056oG/jjms4C7eZrC1
z5IdTBZkkh6sN8ZXDRp3bPg1tl9+dqKNBqVju1xI3SgDruo09ufdIVv2YAVz1Nv7Y7Y/6qVa+cg2
LL43jcI2j8NXdKcTck4ehaL+e8WABkbjY+0Nl7+2svf+k+fiAorLzU98D/ZbTgFjHgworoMAza/V
/jQfpqFyCALrpNmBT3Zs/p4zN1+a3DjL6Qa3kwKe9AURo4rRZ8tKjg1OCEbowjelS/fSmb3czA5H
2WX37h+LxiVX0oqCMlvIcQT+bqUkSRzlntKCYi0akjtwWBMfYHh0DsdBFc1cQi8gtHCMdBfj6h+u
rmZE9Q3MKCcMZiW1L+UGme8Jlep/g8k2Bu/dmIq7lhvtfI+ieyHa4Iq01GKkj96iSiOs8zbQvpG1
yeb7U+AksL5stMao0/IwvAgKDO1mM8n06rbbghKGNKQ6pLTEHEheHkom+NPCglQ269VeMZv3HxAU
cQVr2dgRcGSOxr2UCcDnJf/glkzitpE5SpDJd9jgWO1d6FO35mqRFBhM3bucixPX/C9j/utLeNeK
eAgAqoTLs3gWpNXCx4zGSXROandAPaj+niqarnVG47k/XQ7niycAnNsnHhn5rIrVYOksFsXh+yx3
aCrYw4Vzza247L8HPu8DEMzBIDx481G+HxxAvw5fgqBNoFllSzsmbz50RugyY3Y7lyh9gFwjtZ2N
o594EVKWc2qT/mTtukRqa37MAYtXt9WfVRJD7bJXneja6ckNAReVcVRN0gE4qpj2xh6puS7RZlcZ
X+kBkOqc8QA6DXEvZerH/yGcDtQsJQScOfj/vg9tn5Wvdak=
`protect end_protected
