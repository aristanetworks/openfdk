--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
E1MMT5TD11qbguEsZdGQDUcVKnxETUfxcqTsOrSDl6gIkW+luFKidh8rpvjjsW/YZ3wgBwYgLcR4
LGAn0CyWAu7hkZnupIDVAH4K4ECox2bUaXTb3c2rkAHLLNCZboRAr7vmTHhywB+fVbbHKaMp44/3
QUO6P9o15XncqZl0t8QPY1ggL/mMLVUJAntbxpDQnZ1J0unvEaXxkGY8xFDl5/3xVY6mcU7/KP6v
K9Nhfzyxw+bzkGFFhrlVfuqDPKycaSIPekqpV+6ux+JgjEUjMSX7YSmckkTQjqAlfps4bwzvOmX1
8b3YtgLE6hANQz5a2XcFhBWdtsoqqffxZI3YoA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="mI0IVDaOLn6pjivcY4MixS5S+Qhrvb47tNNe7XArQ7c="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
SMA0T0QGK7bzOn32g2B193fGYopGqi48xdk6Ep5EfjV3sQiACa91Ff8Z04mcklfEV3zjm1lpd29Y
JL0DAsqW2br0lIfy0Y2eYBuv4unGvO5wHQ4vVkNzqrhHxjhdV4wdV74j7WzAgbPpXgDi9vyl2Epb
SDLuv9kIm9yI/tuTeDuccs3931R36r8aJLWbGE9W7yAxLUQdoY7/jpPAUpSxzO5mpTYPuRDq7u+u
76Sup0JwvTFEo6YrmK3Bkd9gjqO9xPYdCqQt4nIltIqfqQbkuaQPoQyz+kE/BR8AMpL4SgroXO47
bMoMHuqfrZGz2XVNo2WvVqaBCt6viuMPDDd/mw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="w+lB95EsUeesEtAmqzSz9YVoChNE4hbbkTmXzz2ORY4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14560)
`protect data_block
c2RudLSSaTlPZQC9zJlh4VSCPbXmXmcR4L5rkWJjowE9d9t+JJ3OXMfzRAh9dgYccsJULM8qg/E4
pQP2lggyZP0HlXd0LK6fLKq6FLLEO1HvIHv0VrdBiAh+1rhekIrVkYlrb8qMV5uIAUYubtSG7rOC
abkpwMxyLscL+czPOAik1AbAnloHlk5R9JlkhiNAEp6KzeiWUGOkvF1YGSj8eOa0ONprlESfgaE0
6+3rKlDlgJoe4cW1hfWByklcmb1lOAdmjLpxQm80rXMnCend0Me/QD7EB3dSzG78DwZIRWEox/1f
NGFTZN65QCeyq9XIPdkVvr+Nb8ay/zQA/0i/tqEvJju+sQ9jVSZ0bNobe6QjuCvOT6HLrER59ttH
80Ey3O6o2c9W0YBhX18nAYV6nuLEO+wrq55idqiPvYK3vjcQm0JMZlp7jerE8zzj3XL0PMPyL97V
+34cyuO+Vt69jqdHtl6OCrxP2v2XYtaX1+8KG49Q4VuHChv4H2uEivonwpf4f2+ICWZNmGBlccfn
7YoFdvDDul2sTIOMrmXj1ndVetWpPgdeT+ItEFMpMZqhunfxxjagPmmNen/K4HGYjiNIhmX1JlB2
p822WORupCq/ih4KEbsVfEpxaN7IXYKO6N2KQWSBM78HIOiD9tcDPEjEVEZPDKev7TMgNQFjoR1m
YFXip8w412aqMilIKry9f7WaOEO9W4jFKEef7ueCMBWZGLSUaV4vC/v7sqBQVfSXvZR6B4rQizAZ
1gNTq/LwnuZdJ5dYtAkQuOHHLMeOdm7ggZBx9o1Y8OVLEyN038l98xHSPZUGz3Uje4byd/CKzlHS
YE9MgbkzkiE9Z1Ju6IWfrC7YZJdvhMXOdrlNTrCXK74m1YkhVHH4GB9zpFjJ75ttjlteMn9hucOq
DcLmFAo7HEOri1HOHNyUXP5ch/Y2AGbrm6G0oJ2Na96/BG2i8ESdbW+6+3g+fdFLm+dI9zRw/lYP
4cjLhFXfinpDQPKIBf+GhdTxf9XghORzOsuVoZhGY9AydzAPsdKkV+4nvaQ3F7pnqdNm96zhb2zr
iCGvu444y2kAstbRQN+MQh4FfJ/FafL1AXC6X1qk4dh5al9KUDywT3GN36N5vAzuG6CcUikRYGyn
cDUSl7ZuQ+U2MMbm8zggnfi1YbmR9MmCrZU2/i9oBO8HV4RprMNZH92sW1BGcPkE8T5//y4j3IQU
35+7vmz5wSoqnneUnsHP6s9unilbisHDIP+Tf7US6U8SJ3W4V2Mp8a2mJngCU7HB3Tu3+qlfO7/3
NPQf3gql9W133It2tFuHZ69GUlflv2mQcWOoUiN0BZitqADx9nZ961kZmbr2Ffoe8YeYNt8soKsS
ed+r4Hn/9aX55hc8Hb4twTDJa4gM5ChQwxg2s4WuFktV4KaU3wsEDORctsXO9cQynP+UaLEj1vrk
TT3SA1oHqqHhhh4FVnZt4Azr+r4iV/rQfgEgRe3Qb8dEoV74m6sbm+3YP2wpMl7I5fHtXe+Q8bJE
W9dRNqgmjKBqSuurtgkEiAv2v8nOxbp5aQbI7dkgI6U0nQi4BZCZNCRIXNjWa8TfcOhzB6HMkREg
U9UfwIyJ0+1+ykulLBEcP0vnEl2TyCPjhRkURd95YcJD0/Z4m9Rjig8NTV/I6KRyZB6NjHJGakrU
AUNPtpQTT4ZcpCPyzSglwtc/1E9ixlUxwEQc/zmngfEVsUn0Tjx2DEl0UaT6+K1s2/uffHuh+2f4
Pode2Zm9Kkc15DEbTS3V7uzKIsLiQ6c44rA4CVW0z3a3f+A/FiuR0sL8vnwuKZ/kmsRdL4aGk3vM
xAxuvznpOPwc8mifSc2a3KUHYnq8oGhvqHtUtHTFHw7rKYxOxt5qZAhkSQ8J2jg2KphfNFSkN7is
g2P6/Hj1v1M1he2ZL18EZq1S66IiaTiDYUp9HxTvXqoGtRXYf/F3lezLB1NyyismHFMafCeKGtj5
fKMnpYb+V3mYDODje4pZTJ32L7Y+SA24fth7su1aM+7oZN8TP8FSe4DYkSCDYgzB/FcqP28B+4Ls
AT6DLuDLdgGCmDXm7WlxtvGIXiFsQtovGSz4N+CbgkBsssfnLtUTCND5FgodHAKIMELZUfa2ejBt
dG7RAc4XFkXKCy0Lv9p7pRRf77at5W+7YpX89NbbXXXiTSGYzUeLIv+cBHlPhMVyfLKHWzHw0rcp
wezxgN5yX5zXKWf54pmzK7PaM2FpoHz+MabE/epj9iw6iyqjRVEUrWSBuKVHerJ6EOCw7HAjC5QE
7IPs6iZydDKi47y4cp30914ijnbfxxHcyesqQ92dOaBmqNGGJLINDV/VJgUM++CPepe1ppkS3rtC
H64XMK10aXS91Tf+rEJRtW2//gVBmiOkGz3/bB4SdaMODehl9EZa7q7HImQVzL3sUB9jtcAA1C8y
InppugtI7NMpjZLvwzGBXrhC58OEVsQugWrgEDIGpUXGk0YasP170Q/hwh6xQDWjEt4R/MvPnya6
6yqQgt+niGWNvIKYmdmAheoJ6/KA3yqrZA2qmVw+jjflcSeyz4gpL1XGhpiEuQl/rwhh9MXN0vla
vEBj1REKcsbRnbVetPYqeNQDWwfKKgKEu9VC54xvCoCTIqi0hpQCAET3TdvJ1ZF/3nqgTfO6AePL
sNIA5ibZSHnBjXqqgj74srnOPigUtXFUupTCwcGRZoCcVENRFJd6oqpaOXEfNny87YpVbVYsgMFa
HwcM9+k2gN4YatdMBiiCAINs0JD2WV3/mUju/exJMXGuE8HsTUGZHKSPxDu3EATrVgrGZ701ocQV
4rSNw6+SacUbm6bfmy7V6YI9iXAd1iASxIaso9PzHHJmQXZAcy7fg/OS89F3z5mrAlo1oVDhpvgx
rUIfpFuueJxw8sVdKvNeqvuIXX/guKRWYxUzZj0QhMNPr78pdHPwkepiKk+T0Wb/kof9EsEQ0RP5
e6UX5H/I0kuJAFfccR7DY54C4YZp99ZFR/WjT30F8f1c5fcDmKowSda5+n4nhUDAZEl+/lp8hdoC
FA35E1Ogje3DzmWcausJmnONnDS82r+vpy2e+FALk1VR3cDxRyTJURSkaS+3g6SNJJFu0UewgEO+
MHt5uSQfwpsTrD/xbxu2xf/MxHRnIVEMnhRb6vjKUDniPlkEvsgaM1iAdU+8/q5jkwj+d56Bnmp0
MOx+uh8NIRH5RxmbDgVWMcSAFCTLles3doiiGkQVH7GR4rv43tOLJhc48Ry9foNL4sMFmtqVSMtR
4JdnF79wJk4p0dZqTuVGdo1YbIrFLn5hBH1hcZCePb8k7oKPvEXr86TdltZc6mVKOa013NmxH6eK
BvTbwHkuUJxsBiR4fbRDfmlWJxNTZfQTIEixYBlak61SIia4zlT/Fzk/wsG62J1i2eGkxvG0HkTe
SwtvWsGgxDyWpVolBACLoQDCqCjRg+dFLfm63FSpjaWhsOP+CCA+g9GVBQiXESuH985aIv6SCone
fFSA7SUaGDB2HttruRvgno++On6mgIrEjOFmMfjDJiKSMlo9JiOxA+1JEWtaFzFSq7bI1RttfZgS
NDaSAIO2mVqLN3Q9SarOAON6asqPX20hN7dlexG3UG9lHchTr9czffnrHSJKCZHqoIZOLflm0ut0
RpRTqyDdH4u2kPmH6ZSWNpVBN5WHrHRCgsyPxBXAkb68UPZBd+eps11SJYEMcg+Z0NV68ERuC6h9
1hN6V2sOd4bNO1cxovwUdgbGWw+YOLzTKmdVdObLouyBi4wbaiLXpqi67qbkmM+rwpcBSE28bTvK
W3xd+G7oQn6Wq9LpDFaMUe0eHSRJsD3qBdGSI/XmuBkwqEqHT1Y3chZtb40qsttuCqFfshPWtKq6
PtNBT0TmC4fpVtnUPvJJe0u3dNom1iyhoouSelE0/qVZ8AFUSJ3GnXmqKkB3srcCyBDdefd80lpm
FV1C5bsX2ku3whN0qnsvvdipxlVEiTwv+G6LePiVdSG7kqROmGPMOyVv+nw7j7clUbYBGW+vTYJ5
CAsY23zyeU203nRwzJadfWW5T2LHL8SUeeZW/5E1TcyAicJg7IdRgfv2VSK37Lf6Su54tYwD/FMv
punhMqHFgMhqJY/QW32dIIvJvhYlEnwk77riglyqhDTj3uDq6mFAlNBCUCoQlkLXqFM7YgnwJ/As
oc/WDpLGvgd8stFsNDV8OU62f/CGnzNi+pmuHHYNq3O1RSYETfYxXRM76rh/hbstLXWwZixWbQun
x94hZuENQO05QfptuIeIiRg1pGGK5t61eRuLa2vGwElQELheI2bBjYI3wC+KSR+OlUjipmcpXFmI
WWzk/ORvKPy21wNGkAVjmQca3j28T1dFDtQA/BAZU3BVbRWEjf/mSEOXVytqXJhZ5emdgok8urux
sC4fWFFPLN19KoyRqjPVfKXJZOBYHrLqvvBiG3giHJheRp1EIHvpM9m8M8Si0KLDGmhkj+5+O6y9
EG4TlnbFWXifSL79J9X9NxJ20A2c8z4EwPsRPAW5ipqsFDVolUyi/CnENTEQYIVyf1wXug5hpk+a
ga/ygJz0gc4i46IQEnFZR0hTjNDbXxNJR9yfIeLJCRDz6+jHEyd+qluIk2y81jfpOSHL43NC1EZX
TcJU14nj2221jyJXAvoykt1tTwHyyibmXuOo0nkDwBO5NLHJClUEFd19D4q2gPsoQzGKX4uMw1Qy
tMdi9W2EzeRiAmduQGxMUyGod/B2jYdV3ms1OLBtaYSgkGBlMtgFjGeVyq8TbOz3VgcgdlT1ErSN
RljIIO4JORyQl+Fv6QATEK4FMIliaDgOyaSXzyI3pJVi2YIKMgRkE/bPw2P7YQ8SyWHPpP9Bw9QT
eeqN/LQDkKDQg0Ej+UsR4YMQ/wxmn/e3wZzjrzbGQ12D6uOisgQ6v4GP8+DmXw9u9H4rrIXJSyE4
6GwDKoYFuKpsFN7GH5KSNT7FFHdvtBHd03i9FqNU9z7bgawZ3/Mmc8lqtBUtp5vR6pCyDIvqBTpL
vRQdUHOC5kVYPzGd6qhVx+36grrKkpT7amx25fKoqr2wGCgOReucBiOHyPF7C38WDflRWPpzkjqW
u2fhjbEWM22mGTUcuV2IpDEmpesAHhyew4/3W63VauDeK2BPxFVc8eN3hL9P0nAmOzaSYU53fQ15
EzQqZJiZwxHq6wTPI4dnzGP2qhenpd9yUCnsjwk4U8bQJ7bXqix/5nXOg4bXP4q1bB5/wZXDYSB2
pHRxAQQoui9MNbm6YiAm93SIiVRODu7BwY97ATpG4XnpH853trTPJJ02/ua9KOyyNMtLPiHloxEL
Wc+t8rsY9sDUqhLDcwelTxT/Qxgym7X5VodC/soA4iFvBhV87R08xgauONnTdSklTEcLDSKzS2ij
ba1bzGwRpDtEndyvSnVi8MLmdx3giS2DCZkjxSxgHvFGdAOfyNUEib5EPvh5vvDJGdzX/XsjK1QR
q+aqKjx++RxlYOq54XRAxJCtPNQCLeNeJZAout8G8Wbm0cLERGtyvaxqiE0y5aG/AV+b5oodu3th
eALWGumWBXu/1FXfJGNOs4vCkuZMDS1RloRtpYr3yoNS/jbNfQKKuCtE9w1b1VzCse0CLGZldBG+
TK0JR5SETarj5ISVibdlKcnuWXRPAaBNoAEv3xrB8h4TEGZ7zFHIWBd1Ww3/tqS/D/Tc+k0eVQkB
bVd+iuLXb6PiXkW1mabHEBiWe6VVJcH9/s7KawbChxFN3+IkDdLcRi0yfAKJFktACCmTp1hs/ekw
yz4HWnqS4PvYM0i3KDndit2aJxhUGAcMwFMuGq6Fep3SmwyGF3Rz3WxYvZiYFO3QvUgEO+X5VC2w
lAMeTzfQiUbKtZRNhBYfuKnAuHrEbHaUleapb7XG0av/dTMC0hxvz0QCkkwtZPIQPu3mMtyf1B1k
fIX3WJFk/+IbeqnsXAkyW921UdIi+dthbEdQ4vc+gbPr73cNBoxM+Txgy5TB9xnGqpEb0Iz5/8Pe
fLP6GNWUmbr5ywSgJOjtcqKvOIGIpF11hH5ZLM8tNzl40Eul24eUuaSbc3ca5puE6b0XQlmqZ4fb
nqik/jfzAxyM+0nQOAIsJCCqmMZrP+N+3XnBYTlbZ/29mRCIITiKyeCV8KDvxhvIvZnrglwmmpJe
Z5juLzMyKu9oxskLgdhrQaC8pTSjFPmGfffSPXDVTiY8lcgXyVsROz2rvJ5s5/UgfFPKquZh/8Ne
x4kfpSOB34H6ET/OLSA4R1Gb3QzBuDrZzvmmoTFpNr+YCAVQno1DGf6iAsFov68SR7PHQxnRcuzu
uiyJFqnzatmXQs3JiJlJ4HCVJNIK1TDLiy9Ar7W3A566MxP57Af92KRlhQKCKk2mNYf3P9Be8haT
H8HkLps9D379vH4HhXbboMgpyWCEeo8s7SMNSIfoA1f/9nuEoyIHVgItI6yO8sLpITSIsOOsDAAl
E4zyyrSjUKV7AhyT7+qX7pCBm5owvrzxkb1ZjcPVkj9t0+nZnjOS8fW9znd6H0rXCFirHPal0HTf
G1Y7ihqLViI3cqc5kBicj+i6WOY6nlLBp1herQaCi+r8oRTwnK26fr57fz3Q2ZlaKGde5lei+Te8
AmxXFZx0P3/rK14uwxJBJMl69gAr4zgTHVr62ImnAJLANwz1RpIClYYFTp1wPeApRYirgfN+iRaX
aL1KX1I114AjWMSD3Lw0P7jtMN0j6NalcJmpct+54Y7kAnanlvHvU65xxk47xA6/+m8Oc/LD064i
668Z3zVQF5eDmy+iDxlCmVv2gQoug0WsimQ6FZI72cP6gn0P3YGDTaDQmhiCtnPwtjZ/bZvAlYFT
zpN0ensCfebC1nhrUerWapYTjHQQZokubAUtRe8R8dPlNYfO1XFWQt+wbFFqtPqkR4Ks3WsM4NMy
UyBcwAvt37OI1p1Ffr+p4nhKUmpUXrSRtzb086Thxs8pFm/nli5LIG2Hpg1VAWqy26EBuYwpM6U9
03E+uz9bhn43XGMBgyQgkvXU9FXvxkZfXRv3Dk+Z8IHj7+AsueEUnaqNoZ4mYcdzgJjCQAfXyAB8
zD5USAbjJsoq7n7hiwuyBZeNkTIjx/aFhoqrIwGLQU3cNsUDvEdTzhbVMf1ApA255BwPaGkpRL/a
PThsVsb0v0cRrc1owjng2ItqlCcMJklA04ORizyU7J5A1Y5pOH7K246D2qRGcOYMDy1F1iYhZgwA
9FVIsaw7yq9IVQ+CAkMNpjP+i2xTZmfMXwgr43gS2OlNkKA/pn5RkVsYPm12VA/eQyrdZd39NUVj
yvcqz5TVXfqKdYrRpEfWEWonwwrFuWIJ0QjDRvzALKlAEylLRGAtgQGLJDGgfNmedwFfg7S6Yzri
GruR3RKjyRjUjIT6fkjZ8KljkBvxgoNgYA/Rb6LikMr27HLZHLKN6lWDsXmNtPDCn/yOU6wtoUVm
v3huEfYhYshg6XJwPFEPzJkCpJ4JKySmdOnNt1IVU9bp5zXqL1CV2RrLJG4m/g0sLXMDQKo/eFCB
Rg9Wo1lE3dCSGwFhU0bqazLveAJ4R63CjI8bR3l7aAI2Bq0BprJlTTcTcNtfwU5caZqabk9XpExe
UDpswWpS9z9LX1toulHvMRvUsvzvhT3gd7zZMZKyXjiFvkZjLWB/AMTpQSQzRDHwIeEUVEnlwRHy
RjEohv2rHCkhP4mYwfkqAHAb4MIgGVoUF4TdKc6tkLZNBP8dtH6A6P3T/36nMjoXmCuOfJq1XUNh
nIeJgFq3kQaFTGiHBkX1b0WFABqv/T8aX342jRwW1s8pXwk0KcbXvpXK3zpyWho1CGVSgjz9bx4L
pjcBtESqT4Vfx54mKHImQ+7CvqBXpKqsmQacZFG6nIZzxzCmGlawkVg9HO32v2tCr0SIy1aU6WHo
QceWS7KTyYVl58kbV9hT1G7lNH+r903ybyCSnJYkwaaFpl2zoe+B8EciiUgdOZ/NT/d71z3KvViI
ObKezlL3iRd7alnoSC8MDLHG0h3LztyOfB8hW9gEhZH5k2BXLARyvhf8W7u/sfmXPwMEdrgXoC0l
4Ie0q1/l9jJONef+MruqoweAja3kpU3d3CFvF10xXsGQVtE/FMuglqKbNCfEi1YoDXasGGW7FqvX
S+dMGwrGHGLbD61l98dWoEbxLTWJo/Gn47cjkOKoDU8NWtRovdwLaK9d5XItitMyY9MEWIyvQwzk
00lTCc1oZLbCJrPI3JW6bIo3cI1vhOgX0ZUrVAK5nnK0CaWQ2XbTg1u6E5auEnsjfXPq4zzEYbOi
qSNZYG0Q37ZfXM3fm2/LMq0zr5QBXw132LaTAv5iC3pHON1O+FZ098gvBRVfDDirgAktvVdDw5Lv
m/2EEDTXEOkw/FU4XYH1NYvKTiQIyoKw9XG64V7YXOdbV1FtYF/giTdZQEhC9w2YdwDNS6zsGEho
+BaJRPfjodl2bGlw+GosHCtVmnfD9eCMGORtNmE1+cMANtDaRRHasJ+leJLCOn8QlPt2L4u8CFxJ
01SYbLgbeFCyl62SPg3A8QrzdR+HVck1+cGe9ZRjg2rN/5+fQVNsinYRlQPHpCznCC83t0aJvEPm
7A+W6jktQ1SgZyo451fyWpyWO8JYLCl4Rd/EnVUpRu5LyVddKnKKbMCI/aeenxzWOaGIOBPcG0y/
0ao6o63bkyNUd7OIOK+cWx5gblfkoNkYeqfS6XhUNTV9lF5t4XblUvoLgbu1IIS7gNZfmGu4JBJX
2MAUFrAg8tiiKOQr+6Icxz6DgHu9CE6U0L1kd5P/+KJHOpLFAEavZuK9rrifGLt4j8lXNxE2uFrp
IAeXPUgliXjbwD/R5XdnaI6dCHZlAmLylVj2T68a5VN3H+1YPIE579KdwnHmVk7kGQct8e/1klzj
l/lWIbm8XNNU1bw0/hBK1gKKoMJ+JeWaM9I55ShLljuwi5YA3YIjJ1R++1sN1SGVDGfJyxrceVaB
t1HYQkCJ+5fe4jvNI6cnFATSlr9ZW5m/1uniH/hxIZIo5QIWd0EbOzeZmK3WSz+2IXvqBUj+Sf2k
0qBeGCILKrEFWpuusIL9RVs80/hDHRMErEYsE9OxrGEg/EB+1Si+FtKStaRTQfhFfcWem9tBUPHy
igShlgBOOIYkUZkEQyKj/j5Ys3JZ2KaL/lwjw+820suIlcSo/kUSkm40lrEIz4J4fi22vRdmcIG8
5W8DeKJ61L4nyrDyKKaUqtIIkGHpchQT0fg2TxZrp31cP7Dh6VYsEsZxgswoTqC1wjWTb62GKXxg
9Y8FFYJ4448Gia0JdjyEIAChFMcCjo3LtgfAmHBoCRmiLsDvhksr/MYc+lGhi2jXqWG6moxjLMOR
Kh7wZADEtdARFPUdfrnvERi7olI35t216J48s5RDW/0SFe4YGEzhPwBAMoX60WikaxxUCFj+Qqn8
UNNo89ecYRMsDsnVcLNTNIqECQXHB4EUI8KVD6AJhHotFRwyhlY8M8HT0f/e6SUg4iTnbt0gBj+P
+gGvSgFJgc3BjABVgpVX94rMQAMfNiQ8Uw6mfHyaCqw8JKgf07AhUgbu8k+t2rXMTg3SiVi62KjF
Nv8LaRO4brNYODiY6XaFCt3CM1wynCZHfbszrKL3gmIaHEHmlHftyamWjQbadblXticlblYgvf+S
j2pZ4Xzdwxye229ux76mHXeU+s7Ub3ST9wIOE32M+5E8y0LVpInNAe6XjCVcfutn+LKd8acFV0dJ
EDgCUMUXOwWXr235uga+yT/YzpekrH498pzqdObhwOGhWX2D6STwV1fSdmWftGt+C3TZCmakTDUA
ZVzMkHJ41jmKHqnPUM4Cj6rVOER5uc6uVNr5PtDYAXn3AJCHhI+BuQhwklGcT/GIqPLXtD2QCZQY
EcYHJVtnr0WnMfgHt2AaSBz4esSHOOFOVOEWF4mQzam+4XjLVHU+0jHlbg9MacTul27MmnUhhPt1
varEENo1fqVCEDGQX94Q328pDdRCQ184BVk9RdRNklHdJ0BvBsSdkccwYXvyugcWBkNe8PiXFLEx
G6zez8+b9dzZH3RNom4Ixb0fUT46GG5Z/ir9Fl+vmbHqnJ5V28cyaiMDy9OXGol8rtnKXzDlDnEZ
YCaWdpmIlK7kJ0ujrOkgPkexrfre+qiWv05u/vBlYqP9c9t2+gK2/RDdb6Pb23EbolT8ssSS3R4r
1iqIqd3Z+dQC1iwHNJDAtfqcBnSVAUcy/Q4E/AbXIBDx1J52Oq3cBjnmY/lMLyvuE5bIFPhEHYop
TtuNRq4sVie9wCvqhrf9fgtro31Zma+3R/N+cy/pcgr8ouK1EonSiwQxtTttjm+FAI4SV4oG3qCK
xvuAzcs11iyqjMc7/St0GXFYOLUy8miG+NO8EZ3I76j1sqdbrPC0a3Bkq/drooso44ZbQzc3ikpw
QKvW6SIxBw67a+6vdRWBi1jFo/jNsZt+I20paUaKOpinN8KkT/QnzwCHBOWoPo3/StXxUUuSFFvM
VGq8izUNi4w61dEQ/M0f74706JHVnoQB8rSboFhO4BHV5pyL0b37VghsE6XJzKxzSlkq/vwcZlN5
6+3np7JiLHtwAHNsSppyM1HlOjAicRu/RXDzVsmchRVXlKA7AoMW4pqImAZXZoAotef+XwS5Zu+/
3bgaeWKzL9CB9XhlmWtQZ403EZs3TrTZDQNgMu3MkJ8A1YOxDH36KFZZnJYSMUx1f/8uKN94Us/l
KiPgqFo1CFeIHLqGMMfQL8pv++Zd4eI4TuaQaiigBctS1ogzFMVvfwc5qAEgp/PUeA0ITRF7/yfF
ZWEIjy3D8mmwKwOZCJezVocsMTCu2X1kkvUuELXeUrwE7RpwnwRHgmj9f9kB2gcvvDjxgB6dxZpR
LAtPAPBm0ybG+5U+vC3q9o4Y/pYR+gq+DM9swYx/hOJvpv5mJvL+6A2J7lX/FnyU6OX5t51D9BEA
sQiK9xdIkWAGUrC+TbJGNHmmF9REo2SQfG+IfABjPZKuRojhdoEPmd5M0xjxqrvNLp2NzIvUtxnT
S4ouhe/mzj4fSfN3PDlB8nfzdv54XAlrVl5My8V4IcwCDLZ+m0EA6IdkFaToGEb7lWWq5qaXxlfV
8l4/x/DB82Ts/+hQyLFe0nSFHCBGzcLHZkn5sCkd3D5YP5HEVfz5DXR8j7C1WeY0Yby4Myqi4mlw
kBCSuAy6F8TqsyNArRReKT0X7etn09oshsIySZP6TuRxaNq8NnSDiJ6qN4237WUSfWvEc5i5sUI2
ck0t8EQ6vRVv+wohizs84J/jwXZ+AOJFZem+p/BSRHpbFdUQ4B7qHL4YJUAt4tyQ1Z/vMw9NgI5x
956YDKxdNhyqEkWqlp7aX7F85hnKbX/DBWKbsZrTlTqYHERwux79D8Rzz4lYpF1q773T3+hEh23C
6Db4HPk/wZUj9kNOOyfsQmU+vy2thNN/NOet5cpeId+40KqJUv1s2se/ZS8vfpAyotUVqdK+JaHu
S1vmjIzYtI0Ka3wHsYtnZZAt1Lqwo5OlDPjfRhLVO2duspBRZXRQziP5SCRKeIXGKZxWYIODaBJQ
+BBizd90SBh+sWQBoKfTZfvi05tLsZzsmqCNw29eqiZCVtytn/hpoXlv25QSbJjXmBE5TxxYaGgg
F38ucKfWStOSrGfXek2Ubgxcs0nz/ZCCURfKvSxQlNP9MvIxfiNLaD0RbDPuVc1gCZ7aRkmdzQUk
K4B2Og3I6gy7eLkXDFRfI+4dFWyDsPfZ8lI2x8jCu9KEw6Ve4xR4Gel/9Byro7cgRixIfLGmErb8
m2egEqvd3jNtenQz/FgIw7OnZDTEOn6KUaYzOXAijDMWzH8aBX3odWMBBk7wTDHEbYFlANcIrUoL
IKlbl642anUYFJIdVP2Rt7kX/kUZfSFb5jp7w1K6npL7p0KwTh3hRHnOyXdcq7mqONah0gHXPCTY
o/lmxNumCPAedBk4M8Z+FhZvBGgF5BM4XT/CO/wa1i1RI1L/kV7yurLawv0qECBjMaTKtWGtqkAl
+WmK6QvwZ2gYFgGz20bwekQGFx9hDk0ZQARTS22/J5VIZdya75fYMeBKI0UjlM92Xy9lC0IJCSmd
sLPC0hIzWQE0X3X+E+fR7uEoboXWRk8tO6Ukjp/ENqtik85V0Ih65AsOx96PVwr5zSGILH6ZvhHc
lYk3NsmpO74KaJYtW1hezAxbLBBPkx+dVd7Z48AprPAdtoYexxh+ct0PjBFHX13ZjZHqmBvz73d4
4B5WqpmLOVKqJ98Ka4MgpdH/IxC7vW6tF67UWYMAM+lk8iVqVvVz0HiLMHBjURa1zdlVN4RwE8FI
c540OT2LbyQo50HVihzo3o7vlBYmXk0uL2g5DkUlpS5JyjBL+HTTR5N5K1kg8RPYHRJHHl84oI7t
71T89ZyEMUp9EHNNMfj5RtEst38ZZVyOqNRWp9MwtgoFLeEic72t1KJVqD16/rCVHK+g7DoeGZxY
ZdNd9JgqzWpFiou/9q7eG8oi5o3QdCWMBHREFf3V+8lFNz7b7tRlVLqD3V9IAXQ96tu3fPY2qT/0
RmY4C+AEi+5O91v74UYLPTS2i/OeuuiDvfbubHzYeF5U7QVIVkYDE0ERhD7ee7zY5MlJzk4MSiCM
Ve6cCH9w10ckAIlSyW6p4G2sFKwsLbua9J+QlI8V+AbxEAEBhaaGouSvRwPYABb6ahMB+t1E93mr
oAdUSbJmaq3mBpEV6fQ+erYGwjyOwb2jdzdOcOg+6XiDzeJoYpkZmsVejP4jPDML2e4giBRed+88
lFGynyC06Pwum8VJVqkfOAh2EsRp19rt7MQIHEVF4epjfxADwcl6dXhknzAtVDbDauCb0sVG2ELK
BFSExJsFclABpKDFXCFLkSdlayUsnciksyEwfqlszjhbONgKSqVCuf4Ige1A6gZPyjvae0zxVMAZ
ASVXHGJTh8NT8AzwMSedh3PbRXJVPFCVJ233CXeH2nDDIzfRgweJO13vmZeP15rgk3Q8TYowSd54
C4kldiyIla/EKsC8A1RUnfLqBlK6L/08Lgcc71wAMYHMtZ0f7yCv7IT89IIGHgJINclJ2SlNVNCe
NoIRFyy1Y2PX8JIYHsfh+yfd/q3yLcxK5ODIfkswHMdhFW8YAydp+xdMo4xx/IwuVEoQCYIe1py3
Iy29EglDO/IQRWW0ZOKFunis4Prfoh2eENaQ9U42HZpmWjCHeIMPjzI6LQ11FJo0v+vU6uFp8Stf
tbX59b/V/Z+fr4EmZ7sjzF1LCNFNqR+Vn8JKERM917QmaIBW0khUxHlWL/vtENXd+XRSJ5AH554W
2qWlDRSdmB0mvjaPOhjYn7iVIsKDCNh852xG6NIpt6+WhN2rLbxRVELqE8Sm+IoMR83GlRajeLnw
jwoAafOQ20HaGX1GfDPEMUhuO1AH6AYKXOTeCx5xzh8CzEAWHXlkuZRwLlNKBHqETwDgutp3pFNc
pldKpVPti7hjOTAZ5WPP/XMZnQaaRj9KbcE1Ta5BQMGXekMCOpAL/recGscPmpeyhr+UXKjtu158
eZdGjbhpCFAb0bPe63iGIbr5Yp3y+bXlW3/6glpIeC3lPPXwc2Alt7TEK+MOtl1TGPa+YSHzOUD0
OlW719tEDths2H/8k1PeYo51vsUaxBqFtEWSEsAfpGap8gzebchxGN0od9Zo5lPMlUxWZWSumEhY
vuZCohgpL3pwSmRpC4uPoOs6ZIgSZvWDuITx0l4030VvZVRO6eJqZ9QCgH092HLS7w5kK9RE4hKe
8XVOcxWTrBul9zZO5wmeRlZrVrpKOZD4CFrPV8OvImXkVtqSgW105os7RTgk3+7Ec7beXaUbQnQM
9fe1mSH2EUx0yfREcgtK86ZuqiydB5TvtWZJsPvMcDmvsiM2S2KWaQ90O+LCIiSeS3eYUpoXAf0O
Ny8VZtyiJ558oBxmIadF6lZv7tMnasanTBkMEYHG7KGOmXl7BdwOX8FD0V8l2GDSpTFkhU3Wk1BR
0fZNMAn0s6097RTN/+oIe95n4gOSZpdj0aopQRTE+KVNyOgsEGwmk8zzHafB3i6KqpJEFb/4Oq9F
RjpSCO2l9Nypyv+ENa/SDpavhn//wIV2iZir997ALdryh7zK3BdHYFbnatWLChv7Zc89DlwluRmG
KL5ZJNJ6UaQFvayfKF8JgTcCnkBXtZfXFFgzUpF1hvQ/IbFQ3XLG3OtxfWscpqSI5lLzT3df4WRK
KvuuLHevGsLkWczXugCcjpdzXaNpu9OTTEyTzUoWrTg6qWz2AnEnFNi6xAV81EhGUq9CoO+k/aO4
Y23QkNaPv3NABhLQIKPhvIskjBbsW8ZDnIuLKG0SwJNaY1k9lUweCSK+CcGrGVFBujiBD0WLqspO
8Yuwyy2bXhw4puT8BYowA/2MwmTihPQvcfcUNCqPcZgTtiJ6mPDQlsZheLD76rzSV1mnrNfcLOwr
+MrwOfj6UofyTqjddHUaCXjoKwL/3NHVzga/O1EahAnBEr/CdWXkfTRJ036KdrnXyszwGRrTKF+N
WQtbKQkPsNymp0wwGTO1bbNw3FC/gJ8XZDLY3CgwgeEjZyOhDhP414x4yWC9NxH6UrNXzAmG5iye
cqt0K63JUNNfAMxIsioD6bqLLMqRtkFmIJda4OR7NBzhxg04N3+ui3SUjVE7k+dVb1GCU3S7SEMX
A6nEPcFW0m3NWomf2wtr9fsJhVHvMHInFBM6z+ge8lbDzE46LUxuddgvw8MRvNGYToJp6+3W02aI
RjIm6PUtsL5bTKHjWMfArbkXIqh9Lx7ARNcWKUBB9MS/PTP8Gd2xGtU9IkitxgR3HodKJVKZln5y
DFwX+6CNO3QbmVnX8Qj/9XOUhEyXUVVIaYSol4F0pNiM7LucgB8Ez3mLvrZGASR8s3CQuFCif+S+
5lylljn/CPG/e8Wwjm4q1pfeZcJ/QfjUVFeSmtXb3RI1JnxhweRSTCqTej5jTSiVyJISAD/aEpDU
8lq+SnoCJLFnbmCCVA1HjQDBJN7ZAV1b828fsMGeVt+hY5lGHOn3Nu7ecA5cqkoxLESpEXZDBilF
e4311970gD1d2uv2f1Lgm7ESjzN5m03qxMZBOP+kKhztCNY54V0ss4Fku08vNb4FLGDP09PubTEk
zZrI/kgZDg+zokrqbTgJttDEIW06Aojv+ox2WJ0TzzN3ANpO00tHYsiDINNecjigD/ToOglphN7e
YuOHrBNOSoFGxPkN9khy7qLX6ldd0f673MbCs4dj9TSH24Me/6Gi8Er9/ANy+E6Wsw3XLasfy9sl
nS0mgcmLKEJfhrik/usZ5bknCi7g2SUXO+4AemWPYm0cufJVR0MHFtyWek5YeZc3F5otqDJWU8Ty
Z01DoyeD6Fst/ezyjUexPoNzfvZnAlW/Lgszd1hKnqMIkLfSfEzljNsGQAtdngvMTwQCERogkyuH
jkxp8ke10NsQJ6BxImgyL6M10DXu+EOb+Ohqd2b5EXqJimnDBL/HNF8CJTtVCMzFCe68wQ94E4//
ARosOsTFSqxeTvpw7QMu/jGAmadWMDxRKCgNzO0qMJzpUljiD8jI/r5qeool8hn4sXwsn1sQKahB
sgMc/2Ej4b1igFt1Nypevbh2p6Dx7X4ICGlULybDMtfOYHWGM/uOAjLN0qNa7SxeAAA3KJ8tRaZO
lfSN8OhTC/lLqNQlNQkD1DWJfkPWlgfU70pf7mNbIfzgZZRHKdTolgx8HKzHfh5IQl0STACzw+sW
/lYUjNFIv41eIs5klGsBh3o6InTB5mKldRBOt4mcntDBL96okkhYM0g9kJnWU/0ke+nH6PL350qS
W20Rt2+xCtwvgRekalxfh2vHCPm4CZmlSpjCe242UI5usAis/NGKCp8wLzZ/1n1j89vsZ3Jo/Pna
Vvwrrfa/7wZR5t2u1GSOP772qCVCej1DeBqIUYWKmAbnAeKUzrY42XcZB4KN+ldtx7HjkBsBQnHf
HaUY95uZALC0/3Mbv6/wwXjKs6RKKFtbAet2XdaxDc1b4AQT2yn7/i1ZMPegrvoTlih61OSlIPv6
BPzOr0fQNtjNkuuoceLzfH6NlRPOMyvsu+PdzbBaNlaouakO1XvHQC53EnHXs2fCEiPgy94/k0gN
Ci+nl9J5NtTLvi7Pys7+Igzn31zFgvIH+uOFlU+aVB5WUuV1FJUEwjO68I9rob42d6p1ea8cKtPH
Yv5leRRC2psCzz3r/3cu55LcrP7PW5piPDVdtSktOj7B57UWIvxLZwRMIHXQ8vf0M/1Cuwswwrp2
LryOt5OSKJcBhMf9x2aQOViGHEereF76SzauzSJiDgpy1bU/ETDwJj7X7rV9sjFBO8q76C9JfUTH
pE3fcHH5k9sP8mV54BwckSAQtxwRA/v9Ub6HY7IWGN8XDSa6dgItr8lGIEx0nP6LgUtmBKMTWhE3
AkZcnstUYX+I9royjEJtijQTtEEApc7evQGHddKLwcKWWOEcdhtdlcfZps33lDiPGx7Cz79WC+gI
SK/quL69MsboyX1tHv7MutR51RijrCjLj2a9szgD/a/bHEOH4iS1F4eWJlDQVB8UhtWuvvHZcxMX
TNvEsqXES/oBRrtfVArLWJtrye9RfI6jG+bnf+TuCe799b3BHliLVSwjyxXPcgJzzACCblqZaHrH
NZHmXjtMNWPsHdxXmnb5mJ1WhmihfjIVjAFpQE9/6PNDAMUzdEGalopC+0+gLBX6XdaMpzqtI6Km
wXtvvinCSq+wPNZe61N8tfbLUgXe6Q4OXhKrQf6Qe6bTc0hLC+KL13EvABra93sA7ymekB5Nrmlq
2NUPNwjhZNCINJFji/y9vVZ82j/if7aJQ7bed4RGzIWzf8n+HRUjqE2rsuoiCmM6QWcCU9UDRQ38
44XNyUM2w42L3RnKbdeJ3GNsLFvpQq6UYxITn0JYW2WiZN3FNocXy1oaXDIRZtIg/621U2Uq4VNu
Rb8oDmyAXtuFYtJ5ss3/qNeMidnRiAXrWt6C7Q1YK9TRdmRQPtpLlyHvjEC4yxnqzqnqvRcjO1Hb
JEN+wh5p97ciiI9Og+xaUis8QfgP74RRwWTqWbjnTyJ9xpjgYukuYcmPOpYM+ZVtHfGuosjNQC2z
eGRDZ+fxcOjmj/8ebEnJByFjRME5W2y999DuqhvWWDT4o24zux8XVmgn84tfvRwtmzAAMnFARJ2L
HYKXQNAH0MW5W0dw4PlONjzM32bcajYz4CdyiyzGbQZE+NP58mIsr/MHGY1ik4/u9aK9axJhU5+L
gv6Ud/jonGo7LTx4KqjFZtqhtqADd5uPOv+ygnQnizwQqnesrErJCsENnCak+E4ttUtSK5zGh2Bw
qq2CdGF8oF9UfSpdkZXHanT6C+jrp+tUwjJEpRVpbH20ypdPUGiP29hmFpv5arOG8vFu3aiJEdnQ
LThfvTV3jFw8RcIv8umQF9fcDLS7jxKiwE/fgQY6SjrI9a1mIeHGKPziOVeoNMCb2kpditZyrhkJ
05PBFvWHp7ECmhYF6nRq11SeMJoz2t2VLeLFy85W1IcdXFDwAYxl8vNdwtUzFXjSpknbQ0OMz5ws
ozoVY6pMZdRkI0dZI11mtsP09CousOqp+ZQu6lu1d6wTU61D/N1ir3WH6c/xSLzx33ckvh1R87ys
jI1eGMYnJCqNEVxnJyYiC3LMh11WWbQXqxoZHMWxA+mDfMuMUUDAXvAbAfi4vTZZFLfsRmYvTHq8
1ACumhnpkIEsDJOluhSZTUum+f349VyfavnyN7B3T4cC/j0M8RAOablM1TjDUMFMW2U5WQdVr/4f
HcCvSwpVqS5ck7PzZr0ymdAvWfekqyZGPqhA5s4i5rVqnOkv+uyKl6xQsPIQ+M+SlNn69PRNVsjh
7aJJDg8bnuYkOuO3u/Diu9CbkAk8hHl8z3UIorouFNYbp0E1HjSkQnjHcRxzKA8z++P5Cy0hZjbk
IfRdF2V4daCf8aS7wePAyq8KPk5lznAHjUY7jDOuZ30bLtSAxrox0bB6zhJT+z3r6iu+Cpk9j+7K
c9rZ8ortMgQlJ2zfIThqD2Z1gCZ/5uJKxMIX+fD+yydWI3m+IzUzBxgq9f784+6PjzvGxS92nqL9
jKJWg6+/EB28H5LsHY0KpACNuNeWMUS/N3zVhQm/E8iAIilyLe795Lmzl/7fi1cgpwMcrHjRkHmc
GT98Cy7lq0xgYjA8wqqgdy2jkKtyDyaIO43USmaoOpnxNVG2DxbuazIPKrTswrhfZ/syGVUzhudt
yh6Z/pKVw1GT7tYrGZK2YmqriIcszoFP2TQ2B5+K++3Uk+h3P2jq6jk77xJb9w4oM9ca1/wb+9tS
J6rQObBRpPn+00uv2b+sbCuciyejzcAEaZSs4EmNmbrvmxGsyTeKky9vluzYSKBOgP0HKiijUtAI
wsgMxmh+t6JAr2grSCTZ8lH8/a6Ap3xDdqvZZzwW0Ug0orFrOBvpHR/rIgUGXt1aMmOYY3S44RUQ
6NDmqkxWjCX4yifTv5nkvFYn1rlvhfReh2Al0ziuhjXLIYGzIMqfOao6cBQjGXJGMFh9mm8jsRR1
ckT7kAo4KndJ4ulHOmiESxP2DV6wAi5j7w4JlUUWorwTNBx8BK2z8CGv80Wmf14MDKk9xf8mV0Yh
ltDEMCkC75YH+lEK4ugABaq8l7HaoFUFjCk/ABqEdZ+N2pZppmFNfJfZOjQ+hF3Fr/GJUC0BsyRV
BiY7swox+hQBEuPDozZXUu4rPtkmOEN10GcP28AaGbwFyqTatFMPLs7sDl3qTt96tqSI0ENu8JOn
gkjXI8h76lEUpXAQNQ9wNL3/Dvo3XZsaae6WN8ki8lDbsT4qx1K2amlt0YFjqjD0OaLWr7rpJeeQ
FtqkaU1Av0i2mLA6KLNDIzriAzAiXauWNgxQJip5NohwchKJoKzcx+UI4pKwIS0mM/U/0Ctz9AUN
eXQjTNVl3ipJJ3ZBmBVTJVuKDGsfTlZjGS1w/oOE1YIy6nEsZU4yMAinzOoDaFTsgXAQbOcfUN1A
KhX3CdYLxZ924ah3t7IQ2Tky/IsuXJxbYxC0lpKsH4nOADbpDXoaBvamZJEnqrTWm9iMETWnYIU3
D71pCeNgV0eugrLThiy9zCgJGBuUQQTTKUmhAQ6g1BfiQfaJKVxkOLnD37EqwY6AupF9bqlHICGv
jlsarwM+SnxxGL46lsoHDgTFAYgw7RyuMmd1YW/ankm3DjZOgvlcG1X6WMcTy410wln10F/F+UqF
VmVy3xpMjMfY04IZcp+kaEzUOcPhH0Azy9cTc9gQIGDVQdkm1Zl9/zeZE6HnJCg1wm4HFyAJrcnM
HhcEgRFBjaqMT55wM+udYXpr4+wHQXAmGqLwHYy4Vmm17uPQ1gVA4B0KjEUGNNgaqREq19vYvIYo
j0BFed6rHMi/GC9f7deJyf+ZHKmPTvOxxA==
`protect end_protected
