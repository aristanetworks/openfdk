--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
RqQrKL+V8si2Fjii4M3iN4qa7TqzTBc7gcRGJaUdLVmLHu6qwZXEjBSI4tO4EPi3ht8h+3vCFR1/
Lh2MRDFvHZcCVqGpaBtSahV6xZVT+ZlplIWvUgfLLBCGyrEQvz57Vh33LEyC4ulnOXikZ9hZ+SrR
GyFja4yE5xuVNzbTvZJHQru9wMTKgeViJuED56BN2KpJqzRfrfVOhpiNlOP97PDkVSarzXm0cxgi
oWC2AxO7hOM/WIxYQXiCokX695oDip1IKtoKrl4K+39+w9YF8lUAvyaEPnt/fwabmaFAKBOqKWQC
ojjakLn3eON/Nz683uN5uG3WSh2kdBBdh9V8BQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="27nIKa6vJNB9tESWLfcjhPxh/YjXV0hSQt45pRJJLKg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
PfL2GukbA4PHAfvQOUozCKb8oSJHgCJewY+8BLhgjRONmUau004wdeYeDyE8f4cvY6TQs/CDt3Mi
BoIj5816qoBvoAAHIaXX60nNVF7IcrK8vhBEp3lQY2iGdU8HwACgmeoL9oQXFHI0nppc+vTwa9o+
8DoZMDCea7qG1Aotfp0WF1ws1whLAqOHVS3ynjjBt6MyeZcVwJqhOHXsqnDOBUNPYdXT7tlUACbv
Cx6Uznz3dFUacqUxS0i1F+MlszvxPf4yXPAO7bf0TrMQQO/LTdcoXn8zfpVgDU51bmwqrGVFZOS3
IbTDBDFMczIdgAdtXJFhzZw+xFb1ORiaGvXCsw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="CS/mjcCpr4FHSJARjNWLmFRReIdQn/Tu1Y8BXXrFGXo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4208)
`protect data_block
Jq7ZcMsqM8zFEe/LRUgnJi/jAgW2qOH+NkT8yDQptoZ6LAExFzF/h8p63swye2XUOneDo5tYvRDc
BLdE3zKotDmxuONFbwy6yR2UY2Vhs4plhmP+yxPKlBdUFt+obMhyVXporTQzJlJ0JBTZoUTZMYR2
rVQ53LuMamaNn37M9A5b4fudU8aaAx3Lnk4fAb7dO8x3UwmmPG/7ya1+BgxTVnCMBMLKHUMxSeZx
T1t7Xl6e9tdMPhmfq/2+2mPKIwJFLww83uLCxBUjmIVfqgAje+wskiwJ5/QaQRMxVRJzy5zBTk1v
jcBaMhKme4m2Ec6cB3rucDjTfgvNzd1QOxNmHzLFb7SQ90DhlIkw8d9tYmdE7hlC+5T1YUByWwr5
OVqpp9XGJ5OB7kwtRfn8uOpVZyLljvqlK9b9LbkSCsMLzoqiH80vFt75X/Jso6jPWCzPj7BWTsU3
yO3Fmrw5dcqWH0m4ZYTZLxTMZNuqHQ/y6mR28+BJmwzBA8Cl0753npBNah/DeuBB7m4FfksB06Z3
pV3QV2mf6EpQXga2GtTFVQkQ6BpNv8EhqWplQR+l27lSwNyHSJf0AUyX4RkvwcU7Czz7y5NoMG+o
Icx8GFIIi6wSlfd3SuEQQqu/XCCfnkCKOSyKqM9mhm8yUjC0RxQtBAa+vGkFLE5t0phZbVjcZeb2
Ggw9kiXjfFakrrVjBOF2ZxUmPcr8afrN9v80ony5eWRJ6ixWW/AjhvpM5rT8sw6Cd77yW/qHEBaH
Ak2USFcJLlt15FbLUwYi+NAXez6rAQoJCuObX8zU+DMYAcxASapnKKFYc7zBEeEw+4NxxHvtGOU0
vQjiauL+un++zWd6u0BdADRoJSUkgG07tvFPGOYoGyUtaGuNdIwhuQ+PNGW8JkL/uQ5/kyMqrtr6
2C+6ERUzmoYqmwmvLsSOwoCqupVdxvak9z4r/IyIoC+wBBpONFOhVHxM0Wryq17HSkMIut6rdBwS
BGmacCsziz/2HHFzHon2AgSdUXcORUmOkM3oD0iyJ8/YKiyJ8v1+rielIw3i5kDv6wMQw6OIwGgE
js0NYEbCF9WNY/HRCpn6hqzcW8JAy08Gi86q6UJ7JnFzPPcKDFS1GKDMCctQM9AIgglwl+Ep9zc5
V+Ogsq0dpzPgjHzM+WK0pc9j4wgvKhzrNdcXWpLMC7iaTf8eBdt002m1wDxrkLYuXlaeNUp/13EU
7i++6wDnYpDl9yAPJUr+vheDtiYy+rO/yf9460AZA1HAAKM8xWTgBW52CXUgXk0XaC01mZNmEMib
RTuEtdVBr9n6RJmhRIDtrM/hgvyo9dQvcbrpPwos2cHugDxjuIyuyA4FrFJQAFwXrrfO7OsWfdTo
zOICmI7+ZLY4Trby4s95MJQiOutP51TsDL7uY6gmWKRV0vCCiQG1Ky+hv2f0d0w/3hEjN1L87AFD
NFv+WkyvIEMYIdqXEJWKLTAhjvFEnweRQBX+/eytF5ln8hTk8KZnGOF4kAwfAY+M9XG56EUYtfHg
qQabNHLabioIjgq8UryVgovoOa6hfBqraT26nTCwW9ZpNKxiTTFqLVl8hQ0hLiwP5HCHpmn76BEd
mvYeXRG76xBwo2akn8IQYeHqHKme9QDj6r9zmpn2pt8wVEXSxGmR8VfYkxXAmMzkWaXvk2DIjwLX
aveNR4GyDGYgPpN2BOQnlNoDGZcfiXYao6yKp01l4oNhqkiYsWLRbG3SMMKLqs2a9OVZvoqGZnf6
LScsdZct1Oox5xGPgl/4gb0UgOlzdqmNDxQgxMs0cUL/+Vncae3NVuTF2FesaCe2qDkw74n+7Lcm
sQa/PQFJiubNeAiSS6a1/+HbTOzn1b767JuOTu8YoAXTYWwlv+jxFMrcTVWCZFrXV3eBpKhSedf7
aVfWCXH2U5DQ5KIhVcCphTO9VVi62xgH7j5am+8e9ioiwL+tLmi8T0qOn3Vyg2dI86FnX8UVTAb3
v0nTidEX2jeAcLz1nv7LmAasACD+G+kRpE40YOYZZWF2yJh1+m5zOZZFeRSdOURbH6rYNY/NUHiR
xHuKlazrMkXG4GURMcCES/apnDSXF37rCWblAPzSiudXfpDTm+U3pv9gaMgesQUddVnwmPAETRii
fbPOWLhVDg19ad7LIz+g2n+saFFeY3P5cQIL9CXjJPtlk9RAzBLcozWJJWM/7o9gMMb89xUoQaA2
ZC1IVZA4OxDekr9QArvfTz4CsUedHZJwLUwTe6RE7Hm/MKpwj3HuBAq/s/GLZLYlPbRUmSvL6+/Z
VccLifUI+0MN81QnslqNIr61NUbZBIAdz3+BafBZG96ctJlDA6bo0OPTJkJMaezcAFCoeYHbnHLw
V3/pq+LfViKOsILI4HtM17R3UKGZEqhQkkbawTIhllSLtSyZKxKMpXdpvfeXBPgxudwkKxBlqhM8
Z+4z+v7i/s0a0lhDDZWal4uq376WveVUkBfZywfdO8UZctPnWZgYIcfTU+vQhCVNF5atmhYxYXSy
QNhokyeBYjWdu9Yug6mwaY5FHDgoXG+i0qadOUB5SKqLo3Eic0C1FhxIPQUWROk6bbX0SxWlhhuH
tyUM89/SjbsNJjgzt/qWFoV6VLMcrSl4PBaphTHvZcLl1MiIYHola3IdyJuSRsNA/eRdmw/lCeFn
n3VGAd8SSye8rKwC+mc7D4RjNHY5YhPU2mJzasSyQgqvwRhZA7R43pt6QN5p+oB/9lWzhNjaRBf7
BRBt5wIduGgUSG4CofVGfEo/BiU/ZkWXwj9WxXmA8cHTiWpN8VUjiUffYSe1Ri3V9hIr7TwZK0eB
HbDQEEPCBHqdKMDHi4/ytnkUeh8Ne7ClrsAISs/W8SFJ/Xqz/I4Qfg92Y5OY7Hqu1jVYrmWXKmEh
ooQ+Y0FyVc5XfrcjJAoHzPmwvgdfZg8n9KBN7zHWSX7ZOFRCwY1BEek5QUC5Vt0QX3dUZEuvT9mu
gblq5iKIymmYZDlh/E6+uoDPHeE6ZFu8p8curNE7ZZ/re+Ic5Kei+sWIlGvqc5okHZCrOggtNthR
aw4oal0CEU9rlASr+N5YxeVyHobMneg9hJn9RfVsCeVzc+Ef6sgdBHoiqnlxwCfzxqyScCtBej5G
J53+Nq/siCYDJ2oNkeH0Cduq+NCQdRgTwoIONLt7t32qZrXs85gFnE/lgzi4zOApZjLRiD51wDTf
pjw6TOJHg+nMs/G5XFi11miD9lNRz0KmIW1k4vPW49b4ZRcTU7KHmHHAvzaeghQDstUwVrpiW4Td
78ZV0gjt68Sk2OYV4GBwsqr+dIpgSvEFV1XKkLSixbFTnPZp/fekw63T+x6caAWwEsNLkBMEOLml
nxO3GvWWoVvCrOfM9o6zEpP+rk1ERV++7uoLDCAr8TDSPrflIFjgT2nE3mAydZASZa+ppdyzPHFm
QqgKf6vqBiCsWn8h+22RPR35JOzCr5ZkxeJ84IcBQUH0bqIvVe9e/v0XYCGMq91swemoFxV1H74o
MT/q7eybKEH301HDVjgYKW45HXYl3iM3wbpDVsTee5F85L5ykiAEm93lF8QS0RvlU3wDwAj1QYpD
11x1A5mQBtTZ9HFNCjnU9gcv5ZVsze2GPvwa783bMhOcRS66xOgvZ4QKkSjFkkbOeE/hGOxYmake
RGUwo028V1tCHpdTb5y+o1z5/LufzwkhubMBDSv6J4oBCtrhx5elwhJrdRJmmoy9IKHN9fE6qTfL
QRb94DxPhB55il+JXM2QS62yUtviHEbWqh0CSyGGCkl/NQPnxYecOTH1bWFQVRRaKd7kbDrU3SqE
sowwktyQZb/6zJXCJQIESabQfrZck5kKsP5TwT3Yy+sJsaxO39WmVqC20mpBZwCcJkP8i0cyEVkl
ySidfJcQl4zx58+UnSfsRXXFURK1i22EWV2/8oBFqFykxMgWfQDKNW9fHwfHwe1n9scMkcWlLDYW
/Il3BnNrUOkqXoBoE7qfRd7IF7dFTheZupni9EGdoMRZky75PdmbxTwbn5PRFMHRADRatz+L7eUc
n1hQc6Y+G/7FSiMD5/cC+cqnhtlvZua8lTUeQp56W4NI1iKJxczXyMjO8T70UVi8ZFahyOtOjtJF
jS+ezdCTzt0QqMFQhoKXTxELQMHoMyOZLOq9gPtpD/mJS10is1yb1DVIBQNjCV/+/4EbyoewOjcZ
IqNuyztNsERkGYGCtSAwcNvM4jovZifXdENRs7kcyT1irXFsfSIdndiDysmChdGjOdHuA1FPwU00
0Ng8ynQ0LCPa7G9VcE1ZltfQ0Ijgm0KMpKEqURr0sS8p+MHYGUeMxZ0EQqFqwS+nhCPp0IOztHOb
Huzm3rqXnYC03iUHQH7PkaB2Wp2MoyfwyXb06Tsz11LzDoDeefvLty8ki/WYwwYSZa22I7Y0x0pO
CCeYqirJ5QsbR2F9AyXFM9bMM9qwxJ/J6YWt13gDpk9Mq3IjdN6F58Tvt3kQHDzmLZE/U4QIzCFw
zuhOD2Z+60vW0aRirOB0RdeEGaBZ4ZGhASrLQ0PA/z5eOA3qDzhJhm0/RheeJ2Npts/ODnVuoj8h
LM7IcqkSTnCacphG4O5oSzmFtz2X+M/fjPYeAX/O6Z5S6JfAbGjW/hUB+594NIKpCtI59Fwi8/KJ
oFYIEIeXqqOwRE2T5pgWAcmjWITDGzP+rBQT1D9d8weOE7exlVCEbMkWIqEC7KQ7uK42yklKEDfm
9m4WlD6Leq79U+B/F5DEfQ4xGewnFaXamqZIvGW7X/a3f7uSPVNF22A4ieiWohP9saUhx1TMUjzz
o12ge2f00Wbri6ZiHK/MED2HZjcwOQ1ojIKWt4MEXiopCRBicJhAxOosjlVXQ30JaCN6uAs2FrBZ
zPGvAG3n7a9NpT8XEugpJbnxn/bxH5dljek3qlVDLwjEgiVivOPCEdGgdt1QpVqCcZGs5xZuG0hw
EAznkfxaUc3Ry6vBJQCE6IEJMo1nqiAQNbK+ahjR3ab4Exdr7aOsaYgymWODICuX+rDP60v2pTPR
6/cX7d2e3QWFJ0kDpbN44PG3T0wcom1B+pNmKbuHjEGY5dRnIjNQmHP8BaDXheicY3hRyckCu5et
5dub84077fjiiTEamfATLzUTXwS6n/nf66KsF4hdP+mIUgcgTcD5iJK2qhF34GDW3f8y1Qcf8sZb
XLKD9McmAIw6vGMDQQev+VlNOaOs6nlv665rJz19Ic8QVyWXFSmSr+vwbcU/UEUVED+n61VmjcKe
nu13UEqnTtgPFDkGxIFFlu+kbMhvEGbgKHRUcJy+Hrk75tWZjqsRzgOMRwMLYENtZWlEus8/1SXi
blIgsE3pKw4/TgjC48kwJfJUR7cwghfaelqPW9qHdHRFfbt+YPNh8oR0rfVjheLSSBiAFOUztU8P
6BnDmlT1vb2f/ojJfYM5s5OuWiYZb7KhesVFmepu+hbpIoNxReOMWRtNMLSozDZ9dG2RIfN53ry9
cFbcBQOwszI2cC/bsf37nRsRTV+K7JUjshIvXtr/7XYbKww0BzZWnRq/qjbLdanxGKMkp1y0Aiax
JHq4aXtjAZH+5GkfVDbN/kQ7yokafB2gIV3DHa7j1jBKGZbOzwRyb4ptU7ICCcs=
`protect end_protected
