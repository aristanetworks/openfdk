--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
XywD57r8jiUYzJAtBr/nmFUWqQuINIc0GqqbqAwspVpCZyWHmxhbyybsJmwo5+4qv5WniQspeIxk
DcKfZ1MIBDN9NAC4WKeAmfbL007WeL3jIZw7N+TBIko7GOVn9k6T1kBgeCxSKBs7YTPRLOTQ7uLJ
4+OL1yN+WE6dfmzu1yHH9yXzwvTExASDRx9epetxuPDMD9J/xI5izUAk20yVZ+9vFmHvkgqq268w
bXtZ/JPc/qwKhgSYsbtAGDkSu8BajEoc7gr70Y+IwIHcwaOEsE+AKspFrTSshjwxhOGbzmLv1yO6
5MyqL6o2/ABg3AHOt/Z5Yik6iDIZjzE/p+0XIA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="bfwIGCWawhKP+zKJ9N2im6X2oBIbxCEd2zDxE/0P5CU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
XblS1N+2npVfqu1DEbkhT2gvs0JqAOqdQBmqcJePP2v5O3ZMkIAFmV1bBt2AJuI8OWZ3NpmuiEZR
cJVNX21jt/pDaTv+kHNK6h8s0KrTUUXWQ14lMRThrSTmv3AJWN41xhXpU1ei3Hy2tY7xXf8EGH23
rJ9xAmMRk6FVdmfnFdV7uflrO+/wI7U/N+Q8Sq4YFCi56CmRcXqwplbhtY+PUmHFN93o4IgXauLu
oT9zwQvt48KC4lwfnKEis7izklJhVCi2caTOBxeqDPFH+/36mhWG685f5lN0CY6A2hNout4kcTXT
uFgFk3/Ul38K3gL2huPv1Ko8O9lmKHjEWdou2g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="59JSQv7itpK/WUoZRCQ3nMgz12eQprZDHITk48/SUiM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 29200)
`protect data_block
yjoe1GqiLM3wV+1t7TrLBnBbyCBur74c0WHYqfM9BZBMF/SJqQBdnVdxyZLX5pYZF7tAMN4M3WNG
1daVb9jFdzU2HuzS0GXuQnQa4OpOGhhl5KFUrXBY2DFMlvQj2DdPYi/5zYcrYhflE4G8nfQXu/gv
IWar+9omhQLwPHFtA9xTT0X00g8IlODDDQHn25oTrW0IU5XpZwTTI1bVDJsosgOOqiB0MK5xtL9j
VwPfhlDwkp7TsbRG3CiGioVpUYionYn6935oiUG+UFumR2oowQXaCRX9Ffa9tAlOA1ELFmXSl3lk
ZIOZMYLQf8v2f6nTqkk37qbzvknjfCCTY5yLJH2mhBHUk3unxsX7uZBuz3Ilx5YOVyf5E0RPe67s
CzFf+ZzEIrUWqO+VbCMFyTQW0ggRH1LimqBWVJ4nLKg8V3G7yvJTqiNxhGO897g9HCPfhtu2c8y4
DKcc8I79Ye+8T32iKLgqzw3P02BWInqOz7qkBcNMnu07+G7j0t0lRXhMLLyiT01s5UUSD2wNqUtI
SsHVRp3+PKQqN/oKroz/PM87zgpMUOp2lVVisxr16tq+KEVIXycUzdZPK4Tg9zx6pDd2lu9ySc1b
VZ3Xe5B1SThe47yUQnDqfLhEhvIebhwhFaehoJ2qWvMM0fziD2gQEnYPIdi8x4RnIJAbLZMXiOs3
Ka7hJjxmYSkQztFwPRsibdSpYqyUi7PwJAWsqCNy6rsBF+Uvqo1hKO7YQNQakzcuqDwFHH3lJcW+
R6xJQuSUfheRMF7/flg4qvR6WlbvlYDgnj6I4ZeqrSGCqVYJH1qJF3A64PMGZ5dsQ6rjU3rbFDM7
XT0KiC+oS4YazbqJ9HqJlLsvYNnaOw0k33B8bdrYNF2a1e7buXhk0TlHIlFmkK6JkOGrRkuBRc19
YzrnwHorQxFY4NUQFWMUUWISfEJVWHwAbHoef1sRq/A5derm81z5PvHFd2cVEZ8YAMZeTzjOjSFS
1ijS3x7bHih9VRU98LWYsoaAXmM7AIFtI8oVQs1p3h6KFsoyCN/eeXCa/orOF7TLIy1MPs8UylXe
GqwvgWHeJtXvTDMAIvrQ1nOdF/P/wJbJ9GN//9Vs9KaJBar2jWhMqt1flqO3jcISuu3S/HCLxzgs
TCEobdSgZopOGVSmxHMP5x+jc3gcqmkIOEAXkiBhA7qZ9+OVJPzWpAV4g3dPifnjfWtoWnvd0oW8
TzyEvwOchk9V/kI4oippXwCHO4fBeOgfWzi85p6k8PHyUYvTfok7SC/zSQwxHM1aOGV/kT+5ysq7
Oqsnk0g6ztncWGIcVNN2pnXGPLHVFHNiE3u2riPg+miJbus3DMruNeH2GOs8QJs6g+/g7M3i79IC
DYvSu5W/AKmN+fP5ZFFMNfVXY1MZw5pXtRM0u05037GW+Hr/utovL1OPSdYuRtx2rMKkZK6cVQ4n
hkeIhlmVQCUxMeVo2ujwGYT26n/gbDCS9h++T9RscD3zKOFBk/eIRKufGraXkpvYevMn9BV3swpw
ON9idYiMUocuhhrrOKqVqOnMTBMxWL8FylzbYlPRSZezfHwbwxSYYuigBYc72vsPcsOKiOQsdcmX
SYBA6wIfi9U7ngN8tpfWkpSiyqYp9zLrBDgIMdlt0GxQJpfB0EE9HBbMx5Wt7mm5RJnERljYvBY2
SVFGGp2Ogizqe35RUNyTvQfRXmIdHoWSATcmdyq1TJk8Q5CKUGELgWTJ7C987aIJ0MbafVUxfyN3
qF7Q+30IVOVA+3czUzxOV7LsEZtb/ksrz9uRrn+6xSxZNlJhdMrORkPJfYvOuPXutL97xEZFSgns
5fcMlTbEKugKzlBww7tEhBRql4p4k/Mdj0EgFpmXZcmpag/r8j28m6jcPfsON3bKbmuPV9+Nq2rY
T38KWCEFH4Jf8iKq9kYP2elGnukyfkv/BdUfenz0xlTr7En6uf9RwrRBtmpxV6cfa2ad5UDAccM7
5Ajl/1r5N+gA1LngMhOA6ua7YOEkZrHB85Jyoo2ZyJ/CPNhjPbCW5Xf0yRXOQ9UA0uHIjBb0Q3xA
M7xpZmzOGsMw4tHEK7rQhyN7CMjcQWJJce7A1VL62U4swujLVhkJWVvnunVlgFjSpPIeSLPHnC+q
Sg3DYYoNGw5DTjLqkQCoDgOxVER07XxiNDXA0H76krEOgedbnQVKvqBxHL2o+psZIV8s40Nx26Os
i/18PN8l3nBY8lgNGjyCRxq4mLoUW6WVHXhPavWwrcof4+i/mpAQDi/+GKVmsdNUe5DTRUNg6amE
EhjWnZoSlcUi1WViNlRuxKZPn//kAxh8Q16eVoHe3AiNWjnZkxCzG/LKNK68kry+8b7A86d4wwYd
hRpVAHAv6lG2BA4Iy7ODI0SlwCyEkwpMZY56hiPe6GrqMWbV6hVfhyTxFf3hbHhbDPRYnJPHl7vs
Be6dopL5UvAlcAV73LkArJ12LklPUy/IQcInhp6qE8MOJudky1y9F3f7T5fQ+g9p3wVoWqwrUDqp
g0Ge2enfk7EOYx2wSunuhxpUFfaXSXo+kJ4MAWujKpjN1NnKNsBiZ/RzAd4Te58YTUAAaZZj/pkK
bN5+zWNhfTT4USsYRQ8P8qw1TBWsG17xWf4o6I5xspVljpowj4oHoUjjxR8eEwFKwX50JklTXiJp
dAoAIUCd0/62Hru65XCpbEltbbHlA4TyDokdREwKTwP2ckpnqIjRrX75btNa1XIS5F6HAquAp2VQ
SVPpQm0wkr6pHO88qd/6mDs9+duIk2/6LruNjYFZF01bdg9qS0NWn7d+dNtAzN85J4CwlkVipTA+
/uV7UXaF7Jwu3xw5fT9LkHxw80NS4WdjCSobhBkSVgbnjQZdbaBgwP6MQjUyiX3BVNM4gcBUaVWn
piJyXUfSW71hJzyb1GDf3+FvB8hpXh+UZcm5j0QDTRKuHGICz681GyDIRuiCDjY3X41uY96yu/n8
oYIhNPxyk4RnoLP1p+33u0jXSNbfaStNBQ8RSiBJrEnxwCOWWmxaWaAn27vXt4YVwWCSLalgyDuw
SfpSjpfIwVanXjZyLEgba1ZTs2Pj3bsoaRjX/sklrI0UQx+XjiV74NviS4TMAmpEecJJDEwC6UTD
00ijtQ+OETb6rW7Pm1fdDLWWMMfMEGWhqLsK/ufEmODyQLblipGaQ0nfolcdYtFK5DNFcXQteapB
S4pVcmwYI8ZGtcsMCPcuH2Es1aB+d8TtLCmu/CGrXeHMKSmikgL56+eVvcuk90m6sPcKQxWYiWjz
LEShb7D/mvumbARfXrgRcJ4pwpybisb9eMpvKUlqra72ckXs+TvMXkN4Fp2IHxBLfMr1PWxLi4Dx
Gj4dajclaJTN03z06pnq4n3BqUu4I39QvVomG6XsVkj2JvhdWKxU7P6rdw0dnYGLNF1r5VHom9et
wNu1GttnXQTjSxU1lrdBfsfkCMZGAGVnew9tfBL97VLTxzK0X7G1pmnFgYOIfqTKY41t1fT2B9Yy
x58xn++7AJV3C4dfcxR5uIlX35qQsz+rbpP832YUWJyRGdOftepEST4RdG09SXsEsuYvDzF8FiAp
Ulr7jwkks5EHFmLhEs+cxh3iIyD4b8+X02xgabQRiNgRdRWFYrpfZuvXvWR38qw3SyMvVEbhMYFr
Dujj9ZwD/8LyhII45wpfUmPDEkvRfBULgqxWu162LeEHAWHh3YSFOOpCQ6vos5NKD3i9Z/+alqTm
oTpKFD4ksPIOaz0csg5P27qiPXvg9sKbTVMOPTugDwF1GrToGFx2QiYk/t6UGlMi8M7z/uOISIo1
cE52MWEj4p2d5QfF+3LvMo1MLMxDUOd857xjIMY/L5EdZCgCy5hS+7qB28/C8W9RAWyOunq44cTn
zu5IMTOYqJl8JwnCuYm+2tAQpSTHNa2PmsOQtBrCkNSd2CKOM+KeJnQrdJ02QxhaQAEzCjRFGl6Y
RGOwC+v4og+6kANym0fLMj82IQN+oExNdVtIwi4CExr/YwFRqStyXWZtQzLYrmCrhcUOzmN9iTNO
AsNZErDxLKdr1rEpABZ90VMbrkOWe1U9zRJ/QgFVYYQLAkvB5RvOdlHKEqA5EqMJMFM65BfrQka0
lJNi9Axwor/jK3Tx6VoX93cfyJBPTR1p8lioy5EV1s0266BX1RDfmRGgLC/pSXfpsrssT6JM3AEl
hSUlzD6pGAxyc4MBTBMbymVNKqe99S9GdsuJmBky66mKCQOS6xL2wTdipct6q4ba3qK5G5pafoOO
DlNk2kxpuJA9nOTVbsSho08qyr7Q1rgOgPyQMmixN/SGE8M7gU2GvYUnQTKGNq/54+MwWmzyGHYb
K0ruQKNaX4eTgIZXSQqAXNroUtnxsiu5mJ97fKZrSkse/xoF3ZQ5O163XpYor0s/e5kXLfR1Xpeu
2UBR9NbRxYySK8RYS88fOK9++yi0hcy59P/3k4udJh6Zi7NgXVwLKKRAhIxPZbV0Jw8fe2kYD8FA
Cc8Jn0oPk+RXfZUlJqvYxCdKkMdlPHyI8RHuX58yzRFI0Pv1lKrjmKuwKYBQ22ujCCmZn2v4hjVi
CrX/TInYul3dsvzV9DJg0vIOhpZCHdrv0f5XSCzRyG5axGqT61ziXVjjJH2mgRt+OrJueJGSoFTJ
XYXL3vDu/55BZAnHboNktlCM2ZpHjyDGOoiezGPvSMFWxsMYeq+ojsiCM4Ay7hOUPvPjQbss+VB1
B3fC4r8zvWbGoNwJDiXThxnv51CwC4m1+7I/KYeCTqNX0apsQrFcjgySMv4pndiy7zeM1KsxTdfr
/md62hjwFi4aAW4CzX+Tp9sAVxMwpX8GU2SJUK4VdDtKVXLDXWQvGOUeGs3hI7+0LeGo4XD0Ql68
jR/9VA77sL5As1zZjToHT0Xn3PN2gA1PmP5NqhZdnmVUaknfN+r+d/4mR1z71aHCQyb3I3dd4kBP
7OBFz/hDe+qH7E10jK9ohhKww0+U0ySDq5L8zBhqwSXRXDFkp3KbjRXiEyCYQ9zo9kO+stXcmjCb
fhizwdJeI0yyzOmZN3vD1aaenqxA8R/x+wr8/TG5WFbkVq8MFuQjNTFtCkcVlANhfQpBIndqrPLr
fVXp06sfqWcLy9zwE+TtgJW4Cut/nfq3myqeA5Zm+AvXVZGRn2MQlKiGWnjblhKm3b8T1GH/uuGU
VAz2UmidGUI4itU7tVopFBeO1HWwFP2LRHcuE0NSnVvOWpzjRR0QLaxjK9j9bIDpwGbJvCtlB1ww
tBRMaq/XmduIRlaTDZSVFuf1E8sAzVmwY4o1K9MhtbU1oMYugPUoAFraB0TmelL0rT28tUGzdhx2
mHz5Cf30bPZxeQDGnzyFoAqKxqSaV2LIqxU/azOjfOIqIl9VQmVG39A2PwQZdKJBcLu6BDKDmuWo
IdYOLWhyJCZ4GVxzA3DMkhD4jZ/Wi/b15r96WQW13zDqxBlCo6CUZ36UCvbvK3HcB84l4KflQKco
1SF31z6Jt0a7Mur5zpXL244CKtuKTKd5kYSfOBqW6g/v1F+0dc4cAPd5upeYgZjVjr9QORcEXIZc
Yyux54ScWugkU42Betu31t+hg+Zi0/Mfcd8Uvybfi15RBA9QD4kJQ6C2hhAjqp+urLQGQyBpjRIB
QMMvcq5N8aiA0yVUyRJkmJgr3CyRtUhby9OPTKLuSoznDJNwMAxDPEpTZ6l+FfjOMfudXFBImwCm
T5+NbiKq4nNK4lBODY17thEDLvHeNh2zoQlV4Mna2ScmVsabsk/b5KF7OmmvOF1jf4yG6UOFHEqB
+kS+T8waVaTqAJjL7niaMVYb9qUVXNgv6xfmEzKNZNNyPPbkcNg5V4Qjb8wFg/yx4oljeGZ8b5rl
QZC+I3kMerz+0gsm30tkCsOQBbrhiq0RVT/R0jjH11fSI64kPc2vEdmE+ZsVkRUvTwjKjqHVE194
D0/oD56Cgd/MEHrNIR87q1+CK0lBXhtbyZsdVnvXCt8vzLme0rzsuEI7XCc44dA501PGUC3xnXoQ
BNqdA0SV58MqOmG4xGhRijqqPKZiE8uS9TyzW09g7ahtHuYx7KQJxN/4G5EBQIbJl7E2djJw8Z1F
mS3LxSzXr5KyKm0zw1tLthixW1eVq/i7jqYQgHY9cIYvehtzUc1PbV63l95/xnoJ05n8eEkoi+1y
SV229/fGxTFWZix7fK7NLcn/OkUxyiLPxY5CH/Fllbv/IIh6y0/h2Uzg0ESOZz+6j6iCm2M8UYT7
LDc27HJZu5VUkLcDuymf9UjogPib7VINy7MJBJVybgEPvFr/0HjLAsuqVsW9fK18TydPdhXmKD/p
GJG4qXRQ2of5D6eX86jxx+4YuK2vFncoCOUwikaw0KrBAzDBqqn11YQaPHju+lbMj9CelCRdhNca
D+CmxTDHyn/vakZ3970oxF1ObIK3R3McneE6YQE7ua4cWQHyOPmgRSRp1EAPrDSzGv+sVW48+NGC
+76FH0siM6rdYWRdu+FXIWQgkVWpnDPOUssI3FIy2WDZnvlD5QO1Zxiv6Vfa7IgEGLB0dJciVLYB
6+yHJbYrjB8nUhMWNjUdIws5ltKef2SBaL48byhIGm+1ifkPazNb6e6sJFOz9NFeYT6nJX6ZL71M
ri3682jAi07ZMI7EHUxCr8NVcCxlnkDDR4M9HVyylsx8UUG7kxNVIUF1G+Y7+iblXqWUYvEVJWOK
/c+r+J8C4ycOyYO8+0YnH8IqbnHHMB1JkRe2sT0dJEa/KdADNNpHPH0OgPQZCtyjaKZLdf7G1SB9
CshOjsDXuiYN8ALfdjFEVFkUPZ+KxIC2DSZBLSGJGwLmGAXA36WjouFYi6KpbY2kCE47mTCnLwFM
zyUc5lXzQE4i8082l0u0YTz0ONNO20PaEOgL/jrREjuhV9SHFLDxscYgpsc2+RgIQ0plujV/34F7
bw0uR39U5tcjQePXi7C124uO1KCzcTFeAOlk7yQdOV6YUN98G4Lkg184FgTeRZDBaqxQ/EkJgTdK
oj6H59BBGNBfLWPaFDuwCvoKEu6k2Q/AMwI1Fij+xbCaJD1Ca+NSnYYfpEZaT2vt1NjHC+fQOKtG
N6adLqYlF28HjrKiAOgBcdYYlRhIfQMAnucDJOF6Urfay0UAHOt7EvUugmYF03l18gR3dYS/LKKl
j9F2YdCyFc26yAtXp/J5OcmlBpLRwEwPGXaWCqiyl6kTdhDjbib+M5sRadyy/z0Y/y764wld1Pzr
7X5iU2BL3r8lzKgAl64aua5tl9pIxrXqN94H/Is02nWp5fM24NVdT7ukLvBSD4+ICkP4sF8a5lFX
nnUPf8kE7potW/ZC0QqVc8gRJwREhMEamhbhLgmdUz5qleZQywUWF2bCzl5kMxvBnz2KT0eX1ISv
Okchpsd/OkuC7pzKYA+4qmJdC3DMq1IEDmpAVOcsJdKNLCsFeaeBWjFxksHnQY5wg5d1E4O2Y3Fz
FgaC0gEGXkrOKIg3tS8eutq1H+g7ciIf3/zqZYGfEwgZDJ0G8Cs8rGafLXUrGlKahFFxaTaY4OkT
43lWGUjkzfHBFw5/dPhbuI0sOVkmGlAkoNRwh+JQgtmq71WdoeYrrzukFD7a5zLTwyCLWymlsdGc
pL0WhD/kVvkgp+YK/GWfp2RDJSeHntf4XgQ5b+TVLiJIi6cHUCDdEnESIAJDpYropS76i+CU0ajq
JeO3Iv/TT1AYcnnLk8B5nFhdDQXqQMfrRCJ8B/enkiEubLUFCtv7j47kAL5zq9LEzjBEMA3ZXNcy
umv4iTlN/hBESBRwqou3S0xNmA1gVporbpciZjSAC3ldg674k8r9TYM9tjwEVK1BnAxLfhIRilf8
lv4m5BjCYXey/AgE2lE9cUkoXyDzS/CnQZsN6lFsQ4nY1hS7rXgWeP3G4arDroyu07vv1Cs9wT3j
qRrzn6K55OD2CttS5iaCeQS2yf/h1kkNReNrLX9SoT8BwXBNEoyrMfAwBwdmpZkuHE1lOGrRbZTw
cs7Klx1Fm3/LnhPdpaRi4Svf+e2bwfJCYlsdW0yLgCXmxcdOe+JuuPETyIbMMXd4Nopv5AgkZieE
vqdRu/27kiZwQn2gVcdlC1SxMaF6BUt+T0OI8PFdzXeo9ITi41jINL7sGaA312DVnxDFrc6uB3t2
SzXZlCQ08IVXFBeLK/gkGD+9dq8qLvwjOyPEnDKQrGztSx03l0sgu2lLib+YZOCEBtJTwi60RulH
AVE3qhj/qh1qbD5qFmSNX0PB475FYbsIOsiNTdEpwFkIPhcG8rj5bF0T2fe+u+WZ3oGukQee/hdm
trgtE5ITB4q3ho064KT6BYcl1fn5oF1/aGhK/y3vgA+QOOP60JVu0tIIMzhcELx3O7dl/qCsAA1w
EdpdHjuput9IBtYBeJfuW2VJm2X/39Nq0WzFzPeaSPirPL9ZQAoO4llJaDK7No5fH+HPwYVt96f6
v6b+NrLHkw2bTr0aOE3kpqjZ1lwo7wVx4zVnI89btCGv9O+5FjDOfX0yBpaIQ/+bH1frvMJDmFKC
PTtsSoIg8iRMr0eWezLhO5On/T1AMQPgY9h0jj4aDVKavSY5goEnNctjOksq9b1pQ+PyoeD7PN6a
fmDFjIy5uXM6r3x1X6Kv4DTt6K2UekWtq4PBMl9ZhKaGtlqeF0hpMbHfiqJvurVyVOYuZYev0u7o
AAdPEnoDpwPRR0CMYwtAMtfAVBblv+MQbtkgvtV/ibm3bEw5nJyrOmFSQ3AewRt1vwYHdr1ndjZr
Z/4CYbpCadQJop4PG5UUUjQf7TKFd1+U8PiOmkwZdt1xojDVjXmQrONQNbk993CX2cpQYppTcyaR
kJtEzZKNAvP/slcpNLHe3FupPOv+Jgaf7kpbBnR3JGvj8giMxs3G+nZ4hdD+SmDhwAElFR+69Erq
kTDTbBT7vtX6rnE4oNK1eJO8lEJZfFClB9s1Rddw+TBb3CSsjxreQY1dL6LSuiuQwv84y3FuHLFp
ljxw9/lEDdO+LKp46AX1NCTbJgOzzhezgn8IIVhdBS23xNJjeAWxasNadEM3XaJ52NkwuQIMjutb
yqxMlXklnR7Jh+kfsi3jluyCCIIusDmUaW1USq4v4bZsp6umdy+OUexODRsJexoCJcUaFqUzojBv
+ZEKdWMWmqK/NclNAjSId79yUzAtkbDgWfw3kAuFaHjgyA0hO7Sqbt73AyO8EBw1EDO1mVx2ypMg
SrF8jRr915ryGo4fdimXHFLC/KKD8Q5XZkFalz2xJKcjqXaOsVA/l1W23ZHCUIeKhlNtKfaCzwoP
CyKITRBbGZNIg0tziWntFt73q6eHLScNUvk0CEyKxbbSg04IEBwfWljxpvM/aYfSydjz8S0AgFQm
hUOvYKv8VxMpHyPacxN/eyOgi4cRbX4zSysfjkWFJdfxBYCpB27VmjGzsgzehQBbjbO09INEqRFp
AyEnsTcnp3Yknf5GO70Vf1PyGm8w5LaCvcUaJg+PwYErKSRn4LgnLx4pSlb/EhECNTET9l8XF9pm
LJN/cpJ43l/xlFsFxis9Q7d7I+KaYSXDsB7JQ/K0ih6H92td1zo7rF/vWV5T/eUlbGu00CV+B+tk
j5b3kOP2ydqcyc1bErmFeQ2MRvTg0grWEmkhYjhBCJG+gfo4mNK8BmGHuHK5MicZ7abTcdzKUd/p
BtxHNK2ShnDnQfP+3Zf21G+36miYU5cKYxcbNOpKJPgdGwOXV5VkteLb8gQuV3C8SuSq7rdHQGCe
80KPA9idf9l20lM69zKD93kM91VajzMKNYsuGuM+y/pXGIVRAiswhaOQ91Ub+bN4yAAdOriMSbxF
4c8TF5eTAfhmIluYfqyN+jHs0WO4Tf1/T8ljRWZur+InxnvNNHREWi68sR/S36TF1sZtu2+s7IT5
ob60Blj2zbgQVLPUoGM9Qx6MztxHOgukmuRHDyAxZXf9ZxqWLcpceIXwJ0CAg1KzWR6iIZgfXfw9
/FGggfIJk0cIxpwMhu6a5Dx1ZrF/O46XQ0ei5hW2udJsFmEUqh3Ah+RszpjNDMQtZ3h5ookEkntx
lV7vXqLbt5hTqntcCmYUQGdKbtBBNf+WRZnbzihjor/nGXmbNAmnvYSY0CRbN+cYqYi3eTmWuoC7
O673CLEm4wuY+I9nr6HVO6/jEm7kkg/VTSogESmZnHeeuE16xtOUXnFEAo5ahPFuISFeWnem59q8
IwbYfFmvGGaC6PKo1SrqOBPgjMs4Nm7opyLwwelxwpxJcPHT8dhSKcEO9VEi39C2j5R1XAIhO9NK
OKlQ/0/0v2QkJ9U4SlKR3PpYgwWab12GZ7JwHu5st7rHOOZdgII/TU9xb2mBqYv5ptfJxZArb29g
Gjc6iGdhKsgyLeNtU7aavDCEGs0we8G2XrCmFfFASG+0CNsy52ar++a1ESZvDQhakQyAxfAuX7y6
P+LN1HHXyXuK9+cJrPTNmXG+zsC1p4nvq9DK6ncJ0wHv83NaNW0QokaxpjHQez1g3nMipsKx8R2p
eDCdy1FSTeHrUR9vwqgxbowZ/WUvcyF6p0/G8rj99UrvrvM5bjmNCEQbkZIRxv664Hf2vXM9nYY8
6e9A8EmB3fpCFceXScevCOnXXdeCr3M14ro9f1CPrkY1bLAc8n+CPtY1uN/WU4RclzPsXDDXKvy8
FSv7IYPDKjJIRiUZjM5sHV9zOkl+N6uXnhG5sw4EppY6S/unqpFXXGnrWNZU9P1ymIOABSbmX5Z5
JNWahhB7HHdz5o4VJo8v0DHqLGLW5WeE7DvEsszg9fTEX0IXajOAVen+urRzHGH9yqVWrFUUCEaO
7Nsv7VnXmOgNsuqZviHkzeNqQgW6T+hSfB8Ox4+zavTLgkwwhCPA4pqbwr4wi62OBAfrlDd73OTr
iGYES1DwThtlEGpoSpdFWVh1opoQDYAVbk7QSesxhDH1RcwioVGfzY6Dhw4h+i+8EHbQUKBFz4to
jm4OYarE8VBf7RGZzZ56lbJ0K72inW2i/1XAzYlZ0dTcUVGqZJkH75wcaSUCVNvzkfglpATsjOOy
ao3MZrH9/jTbjccxImhvhunHy+bjpmncMUWt5smFJ7gRIS5C2quvQOt+sL5F2BrXliMVXDd602/A
PIaU1LTB4nPUwcNZh9i7D/CGXcTswR3UNNC6ydVBufN69gxMLC3XabOTZ9KvOgjNRwWHJMEf3+cJ
XaxbEO/xw0/m1Z/UGEnUEXGWoGR6/8apbunIvBXuut8NbJLRMUuFwZg549h/KYCMQCFZ+05mJGgz
q1qG8FUxo7wcWCWdlalhMuwGQ43I7onMj1lquzZiVUE4UULgGgWgmgciANzr1aWdQSY2ShF+bmyF
59mcmdP/TSxT1UP8Szci0HVDpr7Wdp+O0FKikxxBaiM5/CSIOIZd5olQWQLBfUQmwVowI+/PdbEy
Rz99IbWRE3d+iD28cGn6DcsGtQnB9Dbv+YXdOQXWFYmFzooioNFQRwWFs8qXySGGNMg1ys8TUqST
7CLmh9aVg5lu7qZT3PkRLARANZjrnbfwttdxXC/YNmxestVDKR6bPZzWfJmubBsvtwsLO6/PmKWw
MH8c6uRZu7x+ae+SF6I4IJWPd4LVsRxBbOwk/QGGNx0gVqGAldU2yDmVVJlaMuH53SKNY9fjbA0s
1j/k8arXf+2N4Vrew5GDo1O2BHztJ3NRNAlpU9ZZ6GQYRDDeQd4w3DQSz+Ni2jFvNH5jiPfyMXeq
TvPjCXOiQ6V0hxYd93NnagQSIAcmTUWjPmeShR+wgW3J2F99WPg2cAFdn/v8t+O6RbN5h+fRwM+J
ItOrPrArHV26033owgtCPZ4vZ7+dF1qmXZ8J+su9cutBMCN9vhMk0lwn8ARZRnVSx58au/gkPBn1
QRiL8Y3Y58U0mUXbJao/TVvVJ2y3LnzaN1qVFP1nvQ4gt1HLyGVT2yfncST7bZL9odl+BzB09Rbh
YZkL6L1gg9GHWPwD0KJwz4PbAPC7mwJ+sVPvwTEtoN//FOavPD9BrlUI4TBFygvmFjCw19sl855Q
7kwBCPEpHPDbakirhEENu3biIv9uf2lClVDRTOWtquY9sQYTktF3maNviuPeyPezFWBAePiwhbWi
AzXRUJmWPmWPcogWAdhb4E69xKU/pc2BA7ND/SPEKmh55G56E3FFIP2428/yj7A7o1IlqnT0Pi4S
7iWUrqVwyaPuzJkVygAoO2/n6D5KR9H05i9hK90X41mcfC3jFlwBMZlKkIh5lDhnUDBjsDudiGot
a3wIP3AxGxbDdDeaOVCjuQar2ediw3YkFzDEnKr2BeisPYSeTgpQc72mFGzPGXUxM6rtVRy4Qbw8
PwLrGjucXF8wseVx7AoEKOlkdX1qhlSY6NH74JmzsLZEeWdTjqQyoL86OxF6ez4rBg1ImdkOCkOr
KIms2T56tD1E5Zin+w0LnlOY+X7lHi6IcmUiZ0bMPl0hbYznivd9L3Fp/R/Y8Jt53hw1jgpShQC2
cfWILikZvOs954B9Ot86DflHXhEptz0M2Nuv5HXstfpcnLrlbIZ4P4vi1zWZwkeoPO6sYGx3KIoS
2aJfdScEr5Hpec8xwJMDie1yceZamcsFlnRti8S1w8PCcg/TuD4gPIObehm4COJXAJ8uvaIPQO9o
aDkhIJ7W2KJgS9C7AwMl97RQHoCxPn8FCihFewoQGNRmYMm4ugYbrHKrpVGMgVMw8mGT2DzGK0rE
EE++7XUF6mf3fpKrIm74D6mk/I2LB9cMZy4p7DCZ9hy1q8Y9MjSa7Wj6TA2sElEv4huB4M8GNdmg
A++BmNn865mO29oWUH9RYvoEc19NrktV0F93ywIZgjDtfamjXXVkUQ9WncVEdC7DYqc7pSFksExj
CFlmUF1qvR1kZuKedrUSgtn1xRntmbeBrJdyouKaaVkmAyXBRg0hFtrUFXHO2IzsFRyPkYxz8G1Q
5fShEpNX/J719S7kTRqVcNKui4X/ntMS4ucPliIy0ZbGiFjxcNNd4bm/gRSn0Y0nLEfnS3d1FQzZ
0o2mvoQIKkJH/7JCRHHbUPojikKjS0fOEp7SPOO8Q4KEUKjlSc0Nryq7XsG+yEQR76ihe4FlmUeE
2nU04Pit2BP4bRhgBmfSD2+LO3Ubu5uAPQ7KSTlOCSTvZLtqbkukkznFrLHpRrLU122fBc1Syhb7
NMBtFgdTb2y9XxcdYzZFWM5EHIAqhlprIrdgznGaCWVi0ILIfJRTW0FBKTeiqkwiqY1XCPgLstg+
F0aytNwZXV5N5CRscKm0JoBF0Xf4YAK+e/2pdO0uat99EhYnjWmOPq23sR5+wfKgkiYQIAxY6HN8
vLF6tgSr4e1EVLilN2xa39nxWDIaNUbooC/t7gqQoka2946uAZaligH6PP1a4VwU42E/qvneoK0Q
OJcDqusIXuWdgcYIHZhTiCYO+yvSaqOqfaD6DYnDll/lJUMvg/lR9hiTgkO97ZB/6kFqLlMY5thH
ol1ZWiwylIhZLRe6n/DFqSGv87lmvQe3hLFH6sjL7jsR9MeQuzmdK8r2DO/50y4kr7GQ8ZLnclaH
v1hzgI8p3dzjDSH0MEeOikpAN5iw7IL5S3mXKrXOdg7hB1ApjEFEfFAmJMXyQ0UF1474cnS0NyKr
Uzaf7oPEQji/dkscCUbt0TmaCDU155fvUMmNkPxOX6H4cvVujw83KPM1Mn7R4BqhsebStwWo8hO0
Pf2BYV9L34Kp3zAEXn/QSrsq3bWyZ/gERDSzdgsE4LZxL9O5XBGGGF6Lq5YTeDP68aE/pSASRtjM
h3EOYwaudI578tKhAaRQfdU6am7OcxS1XAKms14dbSDo9qMHDNH8Wmc2jI7MJsQ/6rhGPN7sTQrS
+gztKDUBJWlVd+SFojNKffgXbwHofbkXWxFjOhV961OHsG9xFlFep67N2N4k1r8mKMriktT0Qqud
ZU4Cn2SvS9eEVaDJQ5YlYvlY8yHyAlEfybSCvdT9eXitjGFd2pDbpp3N7klqi1DLBZqG5Es3Aj/m
wqels6WY4NDKQR5GgULrSvK+Tp2xtLwg8e77e5X+fcrm+0qh7hdZ2duwD9y6tcKBhYRcU5cbatNL
UQS8KwczDmLABnb87IJUE0fsbj8Sm3MqgH3pSkvhNu5+laUWOt+yGhokipOmKNTP6Vqy5dwpukje
WNgVigzzH5Inju9tHoRfeVaBlL+ApMrt+HjpGAVKtRDYmxBqFMbSdVWlAYEp+N0AOsJdij2XPeHG
S3Y3WqvlaCGN8Y9nUT3mky0NiewCg+oSq50iI5VZ9JTzClkU2CMdEJm8+F1u61S+Fs4otDi6k0Dh
+JoWyxmZqYwXG8YlTfPakDTKPb+b7CcWK4mXRG5MS49KvCC3FUZY0vcNWQBH++6wTtNT61Oux6A0
x5Bpa9NO1B7fFiI0Bt8/h1JBH9hPhCDhkIaUfxMrcAVtQm8LtK/gzFtSnfl8c6jIpXKXnKyY5loi
naib8wpZwUipjsdx4q1eHDlh6nxgQAy6aMYgtLDQtmdyA24GZx+pFYdy89mPTOwCpfOtazRjmMAn
WP1iFo9mIqlR56nCC+YK5V55uXOlzAQf3DuAht7R+5azntfi8t0TDaO+VEWimijdSAGiIpKHFrqh
mMlasH5Cq8O6xi8/XeRLDNnTGTpTXlGVk8bxuidm06OYlobpmQX954ZMPVY4830tERF8mk7Vux+r
Ro4CXhJYsnbWHHLkNg05dJII3wE38dA7Dat/JZiQyo21y8F9Cxf+CjGOjNrPI7bcWzpIoJJbfc4g
xeWwjeG6pGaACz+DFx6obukAZEwWyTScm+qBMIMBDOW0ZAxB0ncnGNh5/2fG5baPVaqj6IcMw1W5
Dw6MdeuTbDVrFAm9B4F57tJs7mM5UAWMca5ho2LqMgCq+izDZPc7w1PFpE4NJ5V5NnGM3vj1LLkv
QDoj0ruar9cAeyCwIh6L94GEE9sRuHfWFr30QCtWpauirFrHozT7wMQNGYh7dKBw6F2PdvLoc3s3
XXLrlbbwU5BlcmfPYu/7d5pjcej4fRki+sP1OZWI5XextCVX+ZdF0ELqT7blm77juXlIuiRVjxWc
YHpf/H9GrgZ+nrskMnyXAEdzg82PK4OUo53p+9peIvxqEgb1nsqXWwCTcH4qrhSUH7YBZ5f5JIMX
CZ69oS/lJNbldOQhV3IHIQN5PpB2ELyBvLKFm91bKJL89Jn5Y8N1sR9KASciXomfDN+T4ylxeWTd
yiHjJX7u15/10iZ9mB73cuxeDqyYRznEGpWjfXATClASsU5fZYq5UPvjakwL2TtwQvQkTe31wVWG
6/lnzq+90VPS/H6A2tFCGgLiP0zmbipLPFL/JFzoMbCHwqMzuQoT1xd8w0eSEAlwEUf/xgxgARJW
dsA3fRvACOzRLKLGMqD9Z8Xo1XuWglr/UZfgnLoaRSw7oKD9PjEGEuw0LB6md76hLYtKroj47pny
4XFATBiVR/YdhGAgyRaInpbC5I7gyO4rIxICdHOBHFxBDcMw+aj/PoMyKpA8vvbvkEoN8xpSf1Mj
rPpNoMpPdJibJtqeK7UiDzu9hTjTQuujMETR4kWdX+6xBtQeQb8kOFPbBbSm7XRco8QWFi35RLP4
hN78TOridOyFneZYVI0FvCn+BTWkWkMxVEAyqT8ysksXCm+i0bjDanalFPYEEat/DYDvqO0gng7G
age68Mu5TY5n/AUvb7I0GcWeS3rhida7VY59bLsvyVCHtHhR/9LqAp5X+zMU0cmylTSvGHszSmqH
9HZ/yY8tdCmUYQNxPIPm7dTmPa0ZnFA2CyBAgorjMepDtvX0Dgu+xKFbRA81jMDvMzY6t7NcQq4f
EGH+ddI+eGcWD8hHrc9P4MLLYoIGJ+67YHKtOckRlIk3bnmhShFfqPq8wG3lTft4ThpSukgPTFWm
h5D16RFlFpK9qUDBpPEWwtT3UExqrHpJWsxZi1WN9wxMmSlqgnk1dZp1xGbCvNOjbWgU+f4NGoBw
YqUH1FkT7hUV/r0sbjTshj0NDoh+k1E5vRf8rvWmOTo8mwJZhEi4F0WUx0rmD7Gc/OykHsTmhPi/
o9Zg3OeWpBFhU49F0zGrEWiRo5BThCRN10UMhpARTTQ/EniV0kDCKvhgvWhcPnMg6BwbmEcNqG64
MfL4q4nDFYcAYWixsOr7QDnov3i+okbZn+6183Zu0iaI0zBz4qzDOhLnh+qAa1qK3N1aRvLA5z+M
xQC3wNjfM/5Dg7MIzRJ+5dHu7Rl5BKzQfdcolNKB3F0x/ht0/OYsref7UHqVF0HLM7h1pDwKoRr2
nXP6ERrhQKILraisGqefuciK3sMYsdj5p4ghYNmUoDJYqD3hXf6pAk4qTHBjeCCJSVBQ9StF5w5b
HM28dHRIUw4+Yms/GS8dMrPcUOxzHATTHhlNz54ZTeRd9DKINsxN4Iv2qRK/rMRwr5a+3cjcpqCU
VMpSYk/n7G82hjbttcMTmECcZivccHOf7T1n3sk4s0NYAfi8nXV5zvt/Gu5J2zpfqV3rVeLLXaM3
/GP+AIo0VbOs1tXJVAxZNry/yCY+OyTCug7faVL5MvX+we+1GrKCrlcVHNXq5+hlTTNxE4yV7Mwk
BmU4y5U9Kuf6AM1J6UQn9Din8LTkDwSlyRBO7I3hqI7XG1KaGPsKt2r8iqZRZYWvhEG1TSyZsXp9
34pNC667AnR5794sweBjGLTPuPk655ARtx0eQO5F6PfOWYGu515SUtd7uVqebD1BCtsuYFohUDg+
BMxiiKH4N2k2P0Q5s5ammEsMIlpUPe2RjEiwwLT1Or6ePgNUYzOUBN42iL+n4b2o6k+mzaV7+K9+
d9Cxvm49SLch3yvqZbwBLFa2pMqPwbbKubSOuTnpS9yY0RRgyXT8+zc+ZZWI9Q8SBJhajiTARirP
hi/vZ8KOi1rXC9o3QOl590rJCmMDpT7y9dwVAZ8QIBMQUVC5pZkPPmPSUt6XBqUhu2MY5jBh9gSP
gy8uxOy+Xg2YJaApSHWLWV4vAq+OPsExEnVfapraFyjvDzBcbDIuEwpZ+xf4wDiJToJbgNF8GCV+
c979v8zgCp6pzyev50boVQb1Kaby/9WzxfJB0+mUrKofYYh5qpdTXM6n6+7hI4EHcWV4EarWXLE3
Paly6lfhLAH7zOOQjnCPHAquAMUSlOjA8oeQaeiwKD0Z+pUrWWTCIP6o+rabOkDrCxLXAYv+hN/U
6ugFnNLAM1WstWj0APgh/efRf6s1ofdIPIgyGz7YP/Chm7Zzs+k0ZvaaTn3wEAFCUs1sYrpQbzrp
TGwlPUnifOfvLSn/AF3IdUSPpSlLmCLQAzUB1aoptl23BAoz9v9vUMkC1dFftDT7qkHjpB1IwK5c
ugjVB3osM3UAKD+IYC+bIPQOuWMzYnr8t7bK7fIw/bdoBqlnyfJ9tor7N/wvAJROoVpFciW/EClA
iKUmWN92Fg2l//fXHx8eDTrdh/F8m+B8c9v9OU3fD0t+kx/F49d+9R7ghjyYK6N7K9s2ZG9oFFkF
SLrYNDmEWLSdny82rCes36MQi+qFqDjI4EimxFrRnDKMAdLIAQeHOo10NCoCqjQMAGMNti6pbo0X
otMqvqw5o8kPXyeu8vN9jNu3H0RR2tzF9KQTh3XrZgBTafha/4qu46ivCuSQ/COizxHPfC3ZZr2s
GgTkMIwcGZEf+CuNDwzE6uJ3OJBtgirJqEz2zoE50GJh2n74n4uB2cgOITfD8xISG8HUwodq4xjv
4zNj4dc8VuShCaSRHjoTzGl2zmpI/bcK5wONaFcNeTFcecDlNekz95JNkzvcvK+apiv/91KdhQtp
ibIviR8QxT0/97514zbEV6ikGR7MngaP7Tquvx3F0v9sy8FmleAEvs1GAHVmxs+BNoBi/AjiBI75
VMeu9YbMLHfc+JkRHIQU905YPmVFBudW8ye2QP6FYz1StA4Gj2XbTWiyDfUKeiAloWHg0FQ3w6FV
YK+rG1kJMl4KlNGimG2ScIoCJM+tqRBoNvnWtBLIQuL7HTQt7BY3ThkX0bKN4BDGhKVBqP4k+ym+
OiHGeV5A1Bd6h5pagUPWyMxlZKm8GmjbCQ1aIP7H16aqRDLS3AZh+1FETMzoPMajCnxq5HFOvGXV
oANroXeaqoWWiiIsuVtsik8dT15LuE1vhcaYg/pn4FqtLzkYQqDu9HYj5FqN1W9ZzerYnOqTF/nG
BcM1YzXNf/2zg75kFPyvuyv4jU55M8W4l92+k3C2UMD6NNxFPymUGpX/dZLDXOfJ3k/q8QpYjNAC
FggNd1QmP4pOymXOkKUTYm5/ElYkoiAbjwreA+SFd5SfVC4AkQN57nx7kNdPDh7NCC4G1XUQbYmH
MgD5s5fbhDbGGWsLlp96mdIUIKdTRz8B8AjOubF8PTtIpRCJvC4T8/XM5A8Y00OWCvmqL4HOHMzi
glaHxIjMKcc1d/9+sfqYu8Ika1DoUPb/7oVJhDMreHO6wDMvSCTHr++3Ldh3taBSfFkealbQKYO5
9hH2TAiszoJMQsgj0XIsmaMO4u3Tni9MbgW0TwhYChbxrMtAX0LVU5kCMmfNS6qLeexgc99OAopl
LjJastqhntIFlHo6uoNTvCax0WSZSIjvWHYtBDvT4PAwnEa0MchiaTXGpX5xy15+/JgKRDF11BEp
DA0+DIPpGvqrFeoiIkljBHoJKFCWNDBTE/Tp4CHEJOjunXPWZB4kKCjnpfNxMIBKvfq/zHa/uK1v
Z8wVMicYgqGbMo1btTGhHrxwwhNNqgFhqyGaXIQiTlyPr4uF7RgNFchYInzCRtBcTNYGBwyO1P7f
o6AfrZbRuu+Zic58HMvurfJf7Dc4CCvj3UBYHwE+EgAde0l3Z5PJ5Q/YHCsxX8BBgkO+DcSRzCxC
HqwuKf7l9tYgre6atwu2DA6mGZlDf18R2+5LaA3YPRvCdJamA5SO03bR2P2UdXCfaIVs5gLJPfNU
IE4Za6BsXTbosrvSTI2EYlB3HnesGdRGBpkns3KnxoxGdw/fu2P1/MkEJupWXNmi5WD3yiqOB0wN
DIu4ynI4L7QulDU/BnV2bE/sC/BF/hHP4EMd5metUNgqYWImY9JTjjnVroJ9OqNlBDTE2YM95uoF
plfP/xfLkdQAqdLMIiM1Wycz3dBr/9h42Mx3GnjcRWk41+sgp0hAcBG+4aFC1rPf7pv4U34HQX0/
2P2zWb2dr0Y/dR34yfn1J3GfYwHC51UTrVyLv0uB5as3z9HRA5QcBgR3Lr4fDmKSnqFxEDOkPA1Q
dnIa4KuNQG5gZXXLVYeQ+eh6mOvT+c60063Z5iqMOLX44KqpaJjAgDypItrjyTrOJzQuORyS1tta
l2GNEXgigui3L6L6NnuHujqNLsONxvAn2xrnVFCRHy8+wPdW/oYTcE5iOFALJmQoVttT7zN7xkjD
3XHXjikBeRmnZZOahAOtTOSh82a2NgWIeOm6JcMJ310ukXdUIDMtqlzQQRR0bYN3b8Jq9GKAcVJ9
NYh8XvRuW5Yiz3rkx4+eM8hkvoKyOBTcAHbxwl/9xUotB+Ti9mDBLj9+yeYhb39oh9D/btUXz89J
pN43+BuzJGdptXyfmDEpeoJKchh1m8nPpmVbswQlaa0UJJxGBpdCwCSItF0BLxuwUIYi9MRSyNOz
782xVbzTGeB6xXu8oPz1mov6b3rFL5ESXW+dW2iux77uhDbnTNan/IP49XFe59x/mYbvuDiS69EK
dKvE907GmSXMpfGIbDZ2lvsLsEQCcL+99qG1rGp+FANrqN58X04e5HAwdST+pPihx3cgYknTGuei
t4Qu9D01RpDR1TfDvrVN9H9gKO48cjlJtC0bxuLAKpBE6Rjn565MUhekurQTU9YJZkdziqUfhjdi
l/lfDW3lbomreMnYBPYTu9A+m7vKJ6PlX3Zdd9zjrWb9QZAvM9Ic3fTxpsP5NlK0aFXZYuHVKfDN
cX1HigBy1s09AiwTCeN7NKM72UKfqkMoyLvDcN8jwHJXWcqZpvEhzn2trCvYaNw0LI6YkzDBnLlI
YhG9sRI8ylcaQDlB9obvFRcB5jLY1B2jnslBUNTh0ejOqpuTl9gftavEY9/NwlkaLlIvS9ugQvux
kEVmeb8PeWn411cbDD2XkYitdbEjSfliAzZZMPJUxs5NU9Y5w1lqxr0LgIFTM41pUUvw2a0fZ6O/
2eAJ4uYpzvx8dpCuYW4bwAo4LD/SBreSqSoQa6yKh6n6AbPxiRBJX4Lm5bVqxy8ZpG5Yh3AQewJs
YoEbOrJmCGdsTBojeIN18Gdhg6Af3m/qMGGMpV6KyqilNku9lJ9IPMpS7eKJyTTy97Fx6lD38I5e
i/TNFl3oLihAAnpG1xP+/EAZp1RJosUDfffcxpQBFeg9KOLrA20e+W2tA//thgG7ZdnLD14UHNDB
nK5CbSrf9kd6hVH3RGWb8lXLF4Ock/6Q483WG+RiGQ4YuNt+DTh19IURjwmsuUwucfiURsM7KaHR
h1Eg4c9/xB3sZNHVasNobdeiNeG8hUUReP3sZNcl2afQxR2xTmG4KWSHEskPhlEIftdSejteSSGl
c5NV1sGafTlt+Nz2TT+n2lYzAMt85ZgmI1A6oGMhHs4leMup0dCxqwckwqlvJxxPVmRtGgLOYEDK
B9qrtFwVzJ3Aeb92PykL/aJ1I3tcBQ2lZcmDPkPoMcgfFFrzVmTH1hiVUUvh+770zulHIh47jz0s
Tut38g4xg/itiWT1Cn0bjxlKHtg6kWYo/x88xELp9SjYOaAftLusv1zLjoU0qXCxXDjvjGjs5khI
m2AQH1bdIt0IYICsrTR/LEOtCrNn4x5EnZavP463gzxGfnBbVp+5YYIBMPnXnUIb05PsCE65Wd51
GvE71O8y3Co72xqVl+F6NuH3McPCIY+t7TZAHSJol0OfKJlo+0LCsiBst/aIapHQQsG8Mw+qPdgH
MAsERIRwLxbbnwhqvcrmTlXTXTRehOHxnnfmp6c0v3cLRnwTRNTKop8YVeWa1H/8avzL1vZ/A1Ig
wNZLRXVvOoajfVmEeWgLFTWIXwS1gHlLUi6tijCp0MjWE3yjoWJ77GOCPN5S8pghTftAmZp9UDxV
xzu4EvwIVwZjftBFehVADPEFQAIRYuz1VM/OPwCpRq8KB04llJZ9j+XAQD5HjimBiFAk8c2DIuXQ
CPCvmrCpRfUu5mM9MjdLeJwjGhUx+D5hrv3Z0YlRd0CMygrGhjcu0oFP2oVbeKMOlvhka8EGcWeD
Q3czUTlEHFJqgcXEJdzM9vKvC6AdyZQ2MWj0tWCe80n5okCYGTwhPuIbiG/tx/EV0kzu1WpZFFes
Fs+rG/ArcykAZIA4M/7+NICBO6FfvfukoIa0dffxqZajk5wgl5iAsfAWVYm+m4Ou46PVgWM8AL/j
Ozg6lCuRqOwiOezdzP7v5+EuCa4Fzjbs1Cv/Gz8+Od5EwJ7dPDsM937b10U3TK6gwb8RXfKa9qzh
2VNhymV4m4QpqOUxBEtjJh9O42Xwnu8jFdV75eCUpfBC3vnKQMp9h1CUn1uagZz12tZ+6t57Ydus
R0Bl+QmMTZq6iqzn4GAdb0E8DdRMftGiIBwgmJsYR2XaB8MfYiUf0c0yYXHevBAnFj9SscWQpoAB
571m4cq5lsBS07I7MoT6/eQ3SII77i8qD74oMFdGN5sqxk+Q5apBym4QWFkHvnJu6JsR8coTyeA7
4C96iURihsuB0sv9fwfogw5TWpjMYRA0FDTeqfIUJtCnt1wd1onP5JVtQxPslOXJH++jUJzLzKxv
SglZJ+ngommE6LwuYHDdqk/iKG0beBHSgLeQ7hYPQm6V0H/YE1j1iSD2ISuTuvwIDfa+36pAwvsm
ggBEC2rEg6PG8n42b98Bqa+KQazmAEt0ujhdCGjiMsWEkhdX4a9QOPwnGtOkag+S2mLcLbZs8w9F
KpC9n3Uujj4mevn346hMQ14a6pBm+4U6QAHFnVGufQHaBaqTmdB/5zhlgbsxripG3ATl36ln7v7j
lYg7QkModKS5UCwFLjisvkRclD3gF5UahSt9pxjaJYBd+Hd8BjAOfxdcLl0jaVYYYnlIRvjgRR+O
xQdAxrMI4v7WtHCo/yfrdRITvfXx1jI66UosNdMRCUrcmXPrzV2Kc/684oPlfol2cMV1UlofcXVs
UEuWhT7LBI1DRzJbRkCAbb+Biym/cq17zWYJfsxqqFKRcHieWBHaxPmGWIOVRixy/KdfaHR9IxbA
UEaeqjZTuTJUlsapcdO5yxLitCfXufcDLdO/BTitvA9Lc2YSVuGh971LS3mZj43FHDqDsMb5wIjM
p5jfJFWDqA1RXxbuCQ24CCvSg1kq9nN5wx8B6JSQAKHN6y54jLfaXSVmTkN2oyDvflQq22Znk+/1
2o5U+jaAptyccM8tCopjA2OiOj2zKTfZHrCUtGxrr7lvarGEBRMU80KQ2/V/W+mfa29nML1SSV26
n75cgcHYLdDjTi8kHSeajJ38w+7r5LVLZD2hQADUQBFJd4ZTEGEHvzbBkbFIpiN2PzfXGYqPu7Bu
dLgcNKHoRnXCaxuHR3vWQNfesuhqt9pYL88l7WN9aJb4pgUvbTPFKmR/qq31hEXN4CQbIEgZgcBZ
fScvf+NX/ThPAi/Fb9karsdBYI3IeA3gAcYJm7Ha0Q32GeJlYQ6nVi0hg2wkjvGcxvXr16Gn4Zvv
2qBOX8LUL7eu/r9erD8Nj3c7A+DqN6CNFoGJcxaFxt/+Nau2rtD+kLkLM8/v9C/t9U3ZHBRGTyDb
kRBvUQHMMwk2lQRnlU048amygWtgEcmMk/TYMoE033Wsp/sUS3fl27QLxX0ef96sHCcJ4WjizvGS
v3O+f45sMewRC3ztFAmLW71+m5Y7GtmS6Svg8Uyj5+WDe3Ffm/Tqlcsd3A+4xc0btlWuPTA4J5D0
kbGo2EKmhkh7baTi1jxxUtPfPso/JdLijKDUsppVoIhtlJ4ZHyUJ4AH6zqvJaRs0ZASWPxUqiFkC
MtD/Ogtw9Yj5wsayHijGsUD9P+9d4hgkTCJ85E3gNbmywjKl1+dCweeolQ10EaHXlN/ygYtnVe4r
yUl+Ju4vVcgzVUcl9at8i+GnXZXpseVbT4lWhBlQ0zD+Q+2Z1nup62ebNfQrOEUJMwK08ILbOp+5
jKYvYycC8Urk6BKRCmCr26f8EUdnYGTcBJnIUPAgAFIkl9GPhYLO7HPriRZWcAMoo5YkUmIB8RhI
TDB8ErR7EkebXaOyAs9nS6xKneqmHkx0oo8ujuS84YkOhEXz0hlcuLZHWnWJKBw95+BZ6P5KKXDg
W1NW4MOjRf+SPv3r12uaqGZegdprQRIwCoxhaCUqE9RvpkAWaYFaz1B1G6t7VeWSAG1yZriBWdUF
Shf3IInojZJ66VoiHoH/HNvcwD3iPcDG/S5w1BxKygLs7CSMxgJOqwHjKQh5W0VZUCiouWlFCD6t
eSlkQZoMI9H2R3Tzw3ccIGVT2FPLxf6ufTfeIWxd9puCfweMWH/WbukwGflu4ZqBbeTl8whD6m00
DAlGOyh56rFN4K1bgGheMQg7kXyremPHa4LNWBpR/NwG6OYaZJs9bz71ayj+7ku5P2tgYci13gi7
6/4gDjfHdPuCi867RMmNbhqYcCN73ZSoZl2f7Zp16bEdJJE7E4fDfNRrFlKUwDlyXBVHdJEAucKb
s4SDR2rtRacXhSGliuFg3ZByHc29OhTSqHO+cVpuNwcAckUWeIaFDfLeFesuX7fQsoMNgidXiIrh
cShoPn7pkQchbx/UJJrIqbHZwe0murJJ0bMUtnko1Eh2Fl55rFBgZnZ47i/ZfSJYiHqu9D6gBqcu
Zr/olpaQu16hm+H+dHhYp+BOKNsZeFGnxekLFb6vXH+QHKBly4Q+UKAHGBZcWNy0rAH/LfaZKdcF
IJXJG8vk/cmT05JKh8hhs/rs4zm2wh7kPGuAfvocxfQfV+UylDciYAjkVLPv4Hyrlu/2AKX+oRE2
4eyb28KboN0UzyrOD+IUzMsTI9WTITXaGKOcaK+NxXDtYt5r0dHDwvQWZ2sSkB40ZK/arLbijVCm
R2eZVv9yEYMG3Jaut3IS6zOwrhX3zHhltWFPwhvglBKwHD+XJXCPd7PqFItj95osxBMlM9GXvE84
HJAtYtuqOPXP6L3iEp7xd7A18bIXE0ZWmGX89a/FLZYNItJOoVtXgFCSHxoUjeBlg3JyLx+02N4C
Squ39FQM6o7Z4xGemtaRDXFrNsc1LVKpirhfAdnLllXbVHMOpYTK/rHVtu/bzaLf2Ku10Ff+NKT3
HCSfCB1+6nWW5lmaiMMYfIXk3UtR0DoljPQ3LYjgE/2w/cWaRS8lrmmFC8n4/2JJ+6pJaqBktRwc
hmXnDv+iRE/N/UC9X1dv4H2s7TvaXbw7oeQOPqbORphGfcuXxzCWvW4Vqr8SqjFlmSWzE4lOsak4
tEAh6kMBjEI01ziJf8k3sWihUicYavP11gZ16kev29i5RWkAqtZmD2W+nryemdOxCgtNxuEsGs+v
Wm176hiJ1gyv2rOGx6KZnimkzfsJ+mVC7YkIHw6NRNciQ1n+x4a+v4sp3o5Aaand/lSvdoFsfBPX
VKpx9kNPMmAOVyC+mAPtkOa+J9ICsHfJdFrdDezCdi24QWdBUcgBu6RrgMzw2hW7V02OVtFp6Fn+
hEIFQ+8XrkZcgxxbtjsK32Q5iPTEtgcU/JkGRpEcpkg55WBkU53jkinhSGSGid1SkCqIYXWMvMC/
7dVRx/sUDCa6Svl/q7aS3F28jTi6xWxvdQ95i5WnqKrTlBSelHSDkiZZEdvtgLNAOeCrIG0W2qAD
O4vy/PhNuq9H2C4aJx+/6l6GjIBaeqHxjfv+KBRISSQA65NnWxDFhG1htt+lkiMWd0u+QhzpvcMU
6wna3X2ebFmOBrqVWIOWQDsci13MbMJvB86kbtzeXyuDCQ6gY8iH+3CMSzwhKmSkE2LVp3U8X17b
0tB07YcUG+K/sD9mGHu2U8wr54Bnfjt4LKeYIslIFcay2YFUxW2eqXSpKaC95z19dW6LwHHXzDzm
gkevkYTiqXu61dlwQmtwUMuhbD2/VFnH0ZW0OnzMKEIzpNTphAzpr9EWjfa0MIkRJ/XIer+PX6FY
O3lJ/HBw/PUCWfF3SWHNYNqv7tpC6hbp5Uqtz9nZYcnkkPD31tLmJP9ISe90G/bp/fhcRFgeFKJ3
/N0J9PCvy6Vv3K06zx/lYbMq49XjhfbDcxWPIX4HK8NaxkfG7peZ8LSqsLhr14l7Xe4EKUF3OCcR
uvSxfrKV1NM16ICDuAje3fMVldfqpojbuW9ZKgLeJmZ6HRTG33D4kVjoCcKrpHfy16Zbqca2I/kP
Bi0zt5kOfUMYulRE8C6Dp5EpsW1LBBz5rqYmm0FhOEuOyNhOyTVEkukchFmGDwkB98bEXMTPNn3P
RPzEPKNv2/a8TYFEPnLmYwxln4F8kqignx3K4fXmTzYIW2s58+i27cpd6DveL92zKhfkza1K8LD6
qFdeGqxdY6i6iGFIcd/bLto91gujSxI4Jhjs6EwbAo15uXctSRKq0cLsf75APUtOrzW1Zs2h5KNV
zelaFV0/4mXTIvZNl1nGELpK+AvaL6jFyk5+5tK4IWkNWZLtgOXyAum+GjfbZ7yud7IwsLr735li
EUAkQEYSL9O17riJzN+HpxDfInrvfpTcfO3RRr069VifDnYDeBZtkAUuiIj9aLhWyiw78NpZPn4O
0F4gibmqevG8jzkbaK/GjEZxUpCfvujG8M/rMwOuKZX78+UAjmnCjzfeV+ifr1wjExdQpy9QqI+H
qsodl0/2EY2xcF2qyLOyY/C/M5dhxZrmyEH9BQn4bUumSHGTA8l0ZrJiMYOVX/9zGecXPxHcSlIj
J0NaxPosIoUBYI0eDbUx9fUZbyRNi13YzaEKMwMeqyeUBchp3LkNcbhYKF2A+ntoTFNyFQ93bBuH
t/jvy5JxPJChNHKI/eJsASgcBYd78euiNxX3b5P9qpTfUhLYXk1J8HeWMx6A3LkFMvk0pGTHyxdy
CUGsVzU5eId32qaDxib4Q4rKjQMeMYvJ4AVIej0vLFfswOkhwnw3KVrgdnBC1xjIRIQKWQdo/tXY
du2Vxq9U/aNfNwI+0fQWa4Yrn/sTOnBm8fG4sYQ46SgnHq5zvZvOlrra4hVnRTaLlTGRr05eV2Zs
3LeNEW8BdFkpUg3faiQyYclTlWCKQGxVA66bFAuWTKaSs4mZ5EVRr2YFiaHhZ0QYlUaWRWD7RiJZ
tNbJGdhOO2X3dNGKUQOLhRj88hhhOJh/i9OwFfru21F5RLneJSiAa7TQO1fWI0w+pZjyrByIHqo2
tyzLT9LpANm3Fa4a3qYob0aBmv22mTzxlOAUFPY1p7kuA+88hQSeyA4c28cpF0jr+Y4+6U/1HBld
lsgigbf6pKAK7cY/QC/RwRhqRkHbbcMWxcgzF/UlcIkaj/mBtA9udXYy6VtrWiqrmfOjByhiw5fO
9Ynbgx/fxsbTYp5W7+W5tqhVTWW/oQ4l/m7OOl9pX1UOF8m9FxVjqNQT9YVmglFUE05RzpRVn6pk
/erYjshLc6aAm7OBygc59IrXNof5SQAzEMw7HKzQgcfD4MzuLUGEHhyUnPoi2rBCBEPeUSpmdfOQ
R8uyX3bDdEgy+0A27mnRoXIPZMNEUzGL2nELayJ51ePRsY1Myrhs91TRdys08PYiJQD1EqZxPyhh
/YLDUYjHgut36rNQgF75dUqo7+Fm+VSqkE8FSTImY4A8iFf3xEPNbE+hPX5NAhtZ74Hg9zaGYm91
PJJ6o9hJFGSuHKmDtEI4t9rytU+jKZ3TTg8sd31KmKY5WT6WqfCsW3ZNhV4/vymCNLvsdjmqIRMR
nCg/BCzJJBcAm6b4mCXeHxwDh/0obBymxKEm06jcyV/fJSdaOXDxLFAe/l7EgYumOhVa/4kTgbA6
DomLXxRkuyYbv4wyviBhWTkdsH3KJW4dH1HvUPBKNuXH0yVVCXkY+ghVAT3doxhHE/GZ0P2K82Iy
7H0jyTwA8f3Nx+DmULNLzLs7Ri8dDq42pL4Mjfit9gUmI9UoTgaQtFu17yvd+JIqweSu1XUzEDn9
EK+WxL5O11lWM7oTUPA4fV5mIZykTZMJtLi57rzrUA2FvaoI7ccukbNcOFuXnraOULBh5Mk546K6
bOs96hODbyi9ZZHoZocsStopIK95xX8uOD/jc1jtOQTObix+XLLXGyhHLvBLw7jy6o91Obbqv/Yo
+L/PCXNzp7+leXCAiDwHkR63nxQafSDA4S9ygofslqwPEVa8W2/1nvM9qhD+wFUPuwYvO111Ew27
G3iSb37vCf/NOpRxo1S8ARUwG3M1ygFo10mx5mbhNXwJYU7CfWO0FB2XvmuVrjWhrhd7jMn4Vp3T
dJZd5K928wZszJdlXBSpjWvpJ6W1U/+2DxPLcg8GawY6U6VU2KOtpvUsAbSPpGq563AAkVvRqTlD
BcpG2w5520onG4X0dRuDGm3JNG1X/zlAxMNFtzSB/LuhAMJRVsASr2jsigDV61dsGk98lePsBX9H
JwbytR/ojVGem8e5iSp4OXRpdQh29/urs4wfEtvs56snpZoEAQP+rm03K8vh3n0rBVTrqdhD7G/r
JAWTz0qM8WYvCHm6yRwlLdrAhU0ruuWpcsS7BnFUiaTFc+WKkvo0FUc4amiEddV2Zty01mCcDvgI
X6SQMy5kt2TKHeruywvSKUqNuSswqAs3vI1HNa+N/wRhbWT3HTtFnXkROHQfG7P8dO+ohicdjoLh
lQ33yKqtV/lbomL4omA+F6bsLCg9YoyRiaI+GytWMUTOrcVV0G3UZ9hENcccERN/9wr4DzczxMgH
psQfZV62aa0yFA4Bcou/APw2JNxvs7W6tTzk3KqDHdsCbeLp90/oyDUcLj4Mr1zzgQzwbY5GSGog
cWBwRZZ6GKyAKmIW+Ea5oG5C1AzAJnryRc6D1qOpfUNJqZXRABqgztRs5tuSpN566VBiO69asjJ7
UeIDi5zMosASPYAZgJs9Mq5dpPB45tKqEERZeoWbvWRqI1SEhCMlWFx5IhSpeppNpgt9/77keTdk
J2yzKYgXifi0C1nPRge84De9AXv9wBH4SiVBlT8C7iyrbQ9OOVPFfHISjB6UL4wfJp/VF3vVs9bv
H0+6qn2KJyD0cxTQL57QAIOQhY6X02j6kGH7aF8tCY1/yCOarbXeqJszhnAUHOlFpkZvPQ2EAitE
21KrxytLiwc12vd9w+tY4gX2xwR+ytBbdcFTgkat55oX5dx9hGLaDhsD0lLr7EgNiNvoJq7bavQ6
usRFBjcYQ7RRcd3cgKkVJqQgVE0V1545sFqrAnirzZDOAW4RAaH4heg2KAV2lvsjJ6see8Dn3gmj
FZ+XAcbRS3/az9ZsECSv4MQHyP61nsscgi2Y8nVGmpwYO0q0bR2Ip8jAvforDKfWoSHpP8FFTkON
sKrlNckLZXEVfamO4H9ujy6hGRQgF0gAdzQgGDvApEXn1l41KCc2Caz6jXOo4jdEN4OHNmb1Prvx
MurljoS4P9aXXy51/V/sjBvXH5gz4gztB8ZSWjLo9SmcnOhpt9qSRG5gQOequolD4Cf7+z7JJbem
DCirtuRFbQPgli6qOyCNR4Xj4YeyoBwqikd41Qkowy9+YUzEekn5/L1NX1JgCzQNism/Msl6Jp1d
YBzpizUgr9Z5QVro/+FpAUXuL+q6a0ofyYBwqXKlHbPeLKEh6AU2fp4nmVFzlwAAmH/JTJeCA9Y9
UnNqcZAXun8wgtzBOkSibmdOcOSLp0cGbcMdjMm88kdIY0JhTvszZaGE8HTF8GvUXCd6Olsg1QSW
Tn53OHubKsh55TKmr+DY8Kmgzmqj1ghYWcQy2kjbF+OkqGS2XQ9+GVW25m0hkDLlgh4c9HL9Y44i
iQZ0u0HHxLFM/1iQ38MIyPCpqs+4BUEAZrFbgff2LUqsUfWHGiXif82MuCH1QNWlwm31E2WGKttL
pZIXD963rJPkoKHA+js1NBVOjw1Vgtd9eAFzSavcn26ZZtNg7DKu/sVehGvPyp/gkjv0Q09c6FE7
TBmz3MgkczzVfluunkTpuhNn15VD2xLJwnD2XLsVy0RzE29D8h4YAPg5kqvfiMw2E1WJmU36kti/
+vfEnpUIJner7/qJ1uCg9pvxuY+Olt33jUFiBxiwDOahZCyEBA+r1++MWa1nvArXx5WZL2XjJJNA
WFOstWQIPiFFe1I6vGe12flo2mh7e7hG08KSgg3XEAKlO+ZFdAa2QBA/EPqKQPyVNX2OFVoj7XC9
bW6Rma2EkH+YI+95qHfcR2erCvn2BWXM4n51q5PrGZuY8G7Svpd+FPTh276XymP2ykt3/hv0ZqoF
0mfgL+CLtNxELzT2DLYGXdDaaDeNMBa/84yz7WJUeruKgJmb2pjCV4ik+oLGHuac/ub4zwa6KLYt
b6EiopU/LwcKYl3qJeM900Y4CssOB5TLFTpMORPngaXKpbti00rPbZW73ElZiyCe8msIFHXH2jPQ
H084KyE48KHFY02s2tmFatfhuMTSxLr+m6QjWlrK3fX4blVLurryGmQDe9pjEelQt/iS2WO4FKAG
gR+xuTfNlc6EadSRIf9Mwmp/oxhtY8tLeNexyZ4YI88RZsjAUV1ZJI9X/VvyLE41eEvNxgiJAYeA
BzEPP/PpbSuM5yAnKDPUq/PWpKybFcI1o1NJ0t0Cgr/PuBvOJaalm/WtmHky/lLTqsF0K/0AMIBY
NzqjZhRuN0UbPiXPMxr9k0LUwwJzvSB/JkGqRAlhiFIs4P1u9YIy24QHhr3qRcLUr7gGfRGWpQNc
DwnDTGeWxIJ6bkzOC3yHVnZ+qgt9NpI0kPHv5hTA/ZosJHckXzqBHA9UYIJPDyFGsGPcSgeHwpBu
FIdQlh9JKcKfmqYU9fIiWwDo+zSp+4DjyVjybg7nwy8J1f4tE7LC7FFlneNh2Q8D8grJYWMGL2c3
21IsgKHlfhzxDjGZfMql8T1vkr+hnPz1bkHAo3tJwCZICm5TZxUg9agvY19mpIw/WmMxC20Ctxu9
wKZLMgGL8i4hn+IFGBmcPfAZctBmhUfUx/QC+VF0vPDhBm80Md/JxFb3NBF51IgRp9PobGN1KCjp
6XraFHureWjaFil7Ux9n2PKwCC1ZPTryQXs61JRdk4b1TsnhBlj8sb1WZRsZXbtvd3cM1ZC3M95V
qbrordnNDeEhTUNHSlAQcYY9nAKwnC133fW8cB5cug+IHZqcApD2qqTzeTsgFyQrcQBax1N6wDmK
/CZNGbtB+7ABukIvvhzTZ1C52fisEitidjR1dFnvslTAhcKbfbRF5Aqm3YDxMWhIcFtKHUvMBlCG
79FPjtDP7gHoNwCe9LKHMffVIJvfSmU+vyRZEBc6g6p2Lwe7tUkT/PYN6uZ9iyQ4AYJ7V2zucgnW
aPEYksb36YpwPCmjAic0s1LKbNIGIEhv73Imv9ib4g/lbJk2DnW+YYHU2TlB88eRlPbP5F8bha2v
y+fLQql688bKJX0UZQAyzKYKJRKezuUhmkNwwG/1XlFLo4z0+d69fWmsYTxS2yrg3Z5JcvQSWjCo
Z4mKYswFIu3aLDZfMt+ETtgZgVULO0ZOy6Ao9IIa0wVXXDXlXIz99AwPOfb1PcaszgvAgha7tbCQ
ILd0xJ9t0KtAG+0rtwkFVH2dcb7eocgFn6wEu71zFnH15AAKVraPQWKixDpBPRl3KM55UyoPsz4T
p/bWRIkS4KJizVnWqXI59dC5o6AZlri3WWopNHXzEYlkFmmwL5ReJj1y/QImfKuZjS/U9B0ZVEJs
zXSr790gnHB0160MxgDBrMLwbNS4FgE3DHNIw6vSDlsR48FHa6clyCDg4lay0t4j8JX3RiCBlb8S
CKUR77L2V+8Z2TEAszDUb+7JcM+1PfZXJ0gqmsT7jVcWHnMiTHzY/t6wCfQnLs78sLgDB4fVAEjO
+isaboOGC6X8F5YEfq5nNodfi4PcW3FvR+yYYs9poIHw2sxhdGhoOlV9REVQqnRIX6Cu9uVc8WPS
QCr7/Gx7GlDoH6ZLumBqVa6hPdJFyLf/g0bmtmexPAujBCNbLXjjn61uzB2rPi/2bxFMgFPdcFFX
Yobo8/zVYj2UK6lyxebgG8lif2YRkthxwy7YVfmsmu60dTn8UOfGSOwa1tzZ8H5QmbQVZ57UlMjr
+h8RTwLAKfZIu5dqnClCkgg1wTIGdR2Zd/0S6aJLczN010f1Hi9AsORFtCHSRLrgJpHc4BB/AOhX
fSWMQCRB3MJt4z1fyMAFBfvKBsgHKAE2bjULpfWS6mEwS+s99OHKWApGL2Vxm+r+ASpKvfbmWTs5
Xgo2PSn5Mhqv+rZgh7EkZIixz8fpm+uYLwzkSnjxr/kEYCIBnxUBcQo74DBX8SHdG8E3Wpn38CJV
HSJ1SIte31mQykiutmjavGl4n5ER+xSYetI8WyJa+ZcvFuxcniXim89819806W/xLldEIWs9zkRH
9kSRgVlMYHV6VHyOhgg25pSIWxSfELxXsRSZxaNXhfpuyKsudA4Hc/vZR8YtmoYa0WbBKz9ycJIl
ltngiHmLDbghfOgstrrCvN7YdyeRNl99eQiQwG0x84Bk/2Fkj2pgLZEP3cjMc5MqJk95foPQsKRd
dKMfVtpQn7oHJQdAwaBFnZnzvJeYdbZcSuixknhPQgpfu2JiOZdqhkU9uMNvEt4cSxE6vtpbgDYx
R1Gu3ALiXoZbG0OEShJuln40u3k3z0YiqhhcDB3antzvJmkVTljVX59zSf5GiWGub5iJQOxxJSod
4CGGkcVkZn2XLuGMCN2xqUgmCG+rbVmQoGre0GvMpzINTfKFnyPfmtwhDeY9igWipuOc2WWupNrN
lmKmE87gB3A6xwCf87usSf2mu8OVhm/2JRv8M+HA4cxf0yAjpaqj2sYTO3wUgzRcbPcv4waJ+iDK
nsy5291STMbUEUqKBL3o+6oRMzWcSKOO9+tka+ve43eNuSol1lKN54KkqjFWbb01/2u62hwhQxNy
KKAbwBOQpHcpMxR5dp5lGC2MF9HjfJh762X/IO0PUwbXH0IYNEUl/eL7f5TSjim8kc50LiZd4vT3
TRIDKMjnvqVnyZkZ8M+8cL97m9Q3wb8fxWqMPDvE7o6K47OatgrufYtmX5VF+mMLKRCchopj4RVn
wPYuq+Pfoz6cUAimVKOYavflubLikCKOCcvQ3O3En37r6kLupUnfAF8yDDzGVtf8uuCMlzgn1v2J
hortv/FQVKScEK5UwgI5uLfBkMiwKfgXKLlRQ70g4anov5ywVBmnYoYMsARPg6a+UmUWyz6IHd1W
g95KqNvwHYxgm8bess+8rWSxkCdd6IisrX9f/RffGGRxDmuyFywMwtJWgYQg2RVTzuJFX3RpAD5B
VIj9lvYRvvEBxZ6IkqZxM79Vua1090z26ESsfxoQudPexjXCONe4h2Eq93cm4wpZ8Vo+qTnHDOwf
iafTKMW3DxabjD1Bz1T5yIlHGmKuZYX3yYM9zxhIBzFGHAk4+/llcx2FxQYIoCZ03WeT8KqE4wbM
2SswkyxI6T52jNdKzGhdbqDtYIfg4jcx+A7GUfHHxi/OGMYYWGMtjTGyWgzjKU6qqDqdla791xsB
w3nW8DjV0AN8pvIhlyI16+6zwbmTdLIGUSzri22XFgdy44rCaEWganMUaefP/9CICNNBoWOQG8o1
6Hxh+saTHYJR/3D8Lr1sooS7M5BifQkOaPI/FlXxby57HB3QOIbP4RkxO4EXXwyHSBza0AZkZCnj
DP7fogRezYFPry1s98EDo3l/e+KiWNlVi+CF0oHQq+XxIyzTg9Lq07BAF9M5n0bwr5tlapAkuVU4
NQ0H5f/v7Lv374YO2ukb0c1n1QMK/tylAroIt7QU8sqo7KjfO1jUdnDfCensyFPTixOxFHKgZrx1
T+ChjVcWghfETDCCFhiSOhABaWb1YT13pHLOIwIeSBZlffK1bMiGmLLbA6zJ52Hp4WwsTjwN6gZ3
V9Q0vQhRp6rY8IxOwA4JQJ+Ji83QyOYgNRwIB5H7v7lR5bq/uf0tlBElBGI1ezfwJ2tmmji8828w
Jh6yVgQ4XBko96sDjrO66V0ALZSU/KMpHWazXlTZbylzICJYAkqFFJeyTRdBvlfuTQqGoaVIgVN3
CfQMkz9lhyLWPcj0mN2NDEK5Aq7zDXt3CgwHmOKOJ5KWhE2Xf67vnP/B+PsQLdycgdsviW9LbF+q
GNuEzkjGML2dnkuBWpdHm1JEa5d7EH5W/bqSj2o4UIpmU+BSYnUPVqLZkMQ14odEvTpGHHZoQ5CG
WXj0ss432kRi4iRpZCo+epHisdYsp3HQgmPH2ficI+vwcDOTvB5EaCnaE5ycT2gBGBb98GSqTstj
Q+oWx3VmdJ9tAQ2j9HZ2Z+mZOce5d79HYpigxaasJcuyZR8uyHbWMAwCU+oojMRzmJ3pAnxL6rZB
Z2CGgOmwHWDlufMiReI2Zo9U+jiwP9yvH5dN/yZZbfPYk7MpFRVGGNhj+Vj6k4+yIxcsNLA76s3J
41z2EI+U62Mek825XWrEZ/cojwAqd1zywgIfHDRLi5UaWjrWELt9sZe/Un5NelNCXWsKGX7LFzJ0
eU1ettswOLvI0wqaAAlue4JEIFDPpQTr/lvR3mCTRJo1CpmSkGquopuVE8gIc9rsurlcV/F8CU4p
wnHv79btlnkq1m1kOKkg5jClcFUZg/Lk1pF6MVL4dHb5hvLj136OjzPjhIc4VdJNl2gBOYdA7UVM
taLkiR0QZS5InVEm3vZ+7QxohSk2c9qZotubzY8eK6ZSsNCm9zMIANOcsg/CdfSS8YTpZBmepNKD
VXst7WxFEMxGESLMIIdy/0UI0yvbj3s2vpMdF3oaMwIAVSuBjd1q3vq5WwrPS/3Cf44nm1ddbcoe
Sd3faBw4QxfOdAOjzTtgR/y2D/JU8oJY4hJNifJipukk9rxb9CUDUywWkFJz5CzB5FT4NAiGMinl
euU329W+jOcslip5Z0fZ0+skbJQ6+WYin9m4ZTiKP7BtD3798XfMphi2STti1dZZcjeQYOtMnyD+
lUwZdS2oSrnCqUoa/XpKIqsgByMVZ3sP/1I/MM6L02+QYk6+VrTisCLPKcvSb9qD6zth+1LIHWKr
JGj1PUvSe7Hya+d8QIUvFSmCgMC0+MaRd/dT1/tGoToFSbQUpcwJ40yefvdoV3bUaybJ9INo3kj+
TXe4e/mjZUhrf5VTPs01o0aZNIN2ZgDjKfQFP9GRrnTPXvtMMttu4XDBZwa1udRqFlx4yiUMLHTt
SlhJAG89rhqTSa1SadYh6gmx7Uq60FdVZ+INSggP2cHyd1C0mCLGpzOQpeh6DiAgpupkxFf1NmSl
TcRmbmD9nVShKgh17mh9QMnwikTna5PDqdYBGsrg38b1KMSIWExBFRs4qp/Pg3in7K4FkodNrJMs
am5wJzhN/pTE6cq0ra7bwXMr3Lh+5RmbAxsfpn34D7WcHUMd+idWoya4XR9s/yaqOl3qvryqO4vZ
VmJ/NvFQM0BaxHdgWiUH4B9/4mwxm5M07arXlMiJ15F3sKS5g5CUlsDR85JYGAD0nNh4Tuu1ExTF
mh0dYX3/QvpSHhcOllK8ZLfbTquqP5rltTaRvxoysdTyk8sCDXtmrTFaZmGSiCoCnCa4c6OxQhM1
VxAKj+SBDasg7n9eZeX49t26Mw6ULa9TUKK5qmobdBHWaTxZ8/y0Huw/tRifVzGjzIljjqCZVKzi
CXiThiBkFvXoI7nYjpMYOQg1PV881cPZLze8dlScDY9Sf0I0Ov/EKqK9TV4PIg2AglgXAX7Clt4d
RD9N4lzPVrhBdGRCZ61FoBX+hrw4GV2AVj79CJtlOsFiN230s+JNfbLnN7EuBjS3RKD1u7zXVC9v
T/XgurVum+3CCaP98nHJnwFw87RKJoxUooYvHiw6LGtsliWI6/nOblf4Ec2kkGwhP/WdLSsbD8MZ
jhAQ3uuFn+ewmpBo2kzFrf9GojEdAkIsPr2SszgV86d/i+3R3teIrrzX+YeZNCpyBc36QpxvJreF
6tlkC/UurbvBMkC/igicQMG6D57OP1hVl82Ta5j1O9f7So9LTvu824MDgmAZHzNNS8Bl4obnTJ2n
iGu+UBx8SyEgetn5kTJS/h4n2uLGgcw2Y+/FE7ckF4feVtSF7I8jWX/4G/MJxVZLgJQUm30bF1Ou
g62wdAMVaFzNMIJU5Fv0mhmrOX2K7oPGqeNWMvTl7Hfa4LvIsu38XwQ0FLq2nlASk6KEk77Wi2uA
zt1hprOCS/vdXtPeu8d4gkZ8BPqV1/2vCXpoCMCnbzMQVhJuQqPLVzxQaku4rBTBuMURl4f1bNKv
3xy525jQFmiQR7ArPWZk6+SSnEgX6BFgd7gaGw9ijDjMlOwsCLAJVfANeUmipG/eheYnKm3Riu6i
Z/MOl6IMc6i16gGpa63XGXpV8pEb568ZE03UEwiZwIBrjKc0aavfYkAZesQMpZsSkTn+qYTt+y2J
LSnU5iPYCsxEndB1QTDfVxHy18+Ld+Ce9GNBFmK7WWCUv2RAPE1qRwEoMn0O1+CX5UzOHTLg/1CG
+U0wFEAhl3QsDDflu9yRv5o1BSO11Yg0Mt2TWThYjAz6wnSsxoEkWq1e4sgRgHCP9LjZFScumF4I
nXJ2/Jwx3KOXbQ68JieaV41pCqSdHt1M+v23SZxzLCglFcM0D+0Tx9t1uDeHer0hRZUa15oyok3K
Xx7rP8eu6e7VvSOmD8/XIko8Z30muAFTfecINUdmWTCDyeZjNRcMREgCgdRydcLL+AwxpRI4X2uy
iez/7LIIwd/gegXr3WBL732DOkatzz5IchhGd+pjelvIAhTKjF9X3mjIATAlhhFeOZrI02Lgfa++
/NVi5+rM2WjLAL4zk7TBwcuh5/uBSrUpyT4U3ZQPhldeefTiLNQm7pYFMdNqnXgM1rGeSwvHf0Bj
HIgFBJB5XJFRhSU91jSUXF//i1/fx5fJqjVD3O6iDA6Dcr8JGmAlpCR4djMBV+xFcK0vRlq25SS7
Y1HGDOu00Y9JJJKR5vo5IOcx38LweiP7dq9DHhcSrviJFlHIWfaduHvJIIoIBF/zGzOOXJUzPUED
4BB/cIogxExiS0RTvtEf2N5FyF0YbUa/6Anyi0UY9U+f1ZPkp3Mvrl0v13l9uOBn8dyPhEH3SqhI
umKm7RUVt5RAIqZrbwblQQe0oc0l+9vNfuV+KLIPKACVEtLHIjpdawnLMSbFrU+uatxd04TpYCAa
gcUV57lYJBmsZl2/hzLUwXdY3d0wvTFJNeSwRazahmBzlikDLJazuFkc3eW5ax2mJj6CxcYR+DUJ
wkWZZwv65TL2M04WSRsswyDrmV/+Linf9xiS/sgk7xALywntdetLGo5wiqE2aHpN78WswKDv/44w
Tc6AGV/xoi5elp6ZCEUvkZBhSwd0EPOXRtfCe3AlbOFb0ZTJRYX5zEAtlY8zWtkOcLsYtK0Dle+Q
H14lmprzjZGJINzyBLUs/KjaGgp+RAUSqk4wtsy4WsuFG9nL+vZCVmTgsBI1cJ32DHsivdZGHO+J
5sBFEh1zrfRj1lDX5zv+mR3w0CKrEYHmGha5YX/UV7TdGbuNAu8z1P4ACYBEIspZfsmmuydMDiDS
LtT3reM6Kiqy9NF64E3Y8XbXkPQxapAQzHD1EOnDgfR8RUdALBJKk45x6+j8Bs0pUQZ/FjAWIMY6
D3N6cw23wsDy3xt6QKOMxnaVH8f28zHgD6BLeUZ+HOKBwzL39f1yZ/phXxa4+LF44fFGAgS1Mxrm
WaYu6yQFVe/KEY3YtyC9do5k1Y6lcJuVUFF8+A9cZoz++7rvkw/5wrqMI7VBmK0CgTLmd+gLmmRV
RMTkNRtmgYuAXKkm5iB2g89jkh3k64jTK4l86tcT+DiXP0uOxdyEOQEUa0Zpns2vJ6JDSceAM3IZ
taVjQUET5zxlNiHigJ/SHBLZdvNNRzeC7Z0LQUDD2mCVkXrJ6/VypEWLdv+OpMhurBk1ta/ny33u
tCm6ExQrIRtQ1cTe7rmgTppkWP0ynHdTQNREOQwJsMUfF968ZF7+b2suRvCNv3uprdlEYwdrmnSk
a5sUvTfJgDOXUJewXyiiJkhiObKUlQmmzoXzSmhfy3hpP9Kh15+QqJhaM0c6A1bbsmRQsDma7+Ok
IAExU/v++IFl1eNfXajYWXXvXpE76eCYB9UqyKifnwwX3pcIo7ws2A5F7+eEKEGGIprEeeQe9tf0
4yCogsgrQ0QSNItDuHaOJ3U3pr6HfInPj1OhdDWr0oECvatpYAjOB0G399c6Ws/zYEz8CMp6Vb0n
iaK9YDifMzKIkLxDjfdtKdvrQyF08OPr809aW7mOR7745+TErnIV0QtAI9k+GkbTDMBtUqqVM4Qb
rzIfhx2Fp2e8+swBxwx1HC0iKwDAYiAs7uXuC+v1lVV5Oz3f0OyuNMp7eB+PvIH0qQbHEf0IZV0a
shj3eE5mITpMKLkJrATB7sh+19UrvFFfsxWJej1CjlQhAQA4+OAlM5U7Mo4MUEVE0asyp5pCjLdO
41tM+YmmCVD6mJvQuyMLsxiO4jIzs1kj9dKGaafys84eDqYxR8D9fT9gJlcyUP7ECRQ6Vc48znvm
ZNZn46PLla5cuFn3ZRvGmBdN6WYlOpbYwD5Zi7IeSIJyftNQDvIY39WPQFQnhS+cok368lTdjvSU
OhoDzmNGzk8cslLbAq91XgeAdAxHlM5eq4fRPPwZ0pFwSucexZdTagsQzVh6ZosL+0LZ1Rgwsk5w
bwxOq+3grs+vADQvOToh6dOSWOKvIr8lZ6kOV2zFeLptktGkqd3EQBe58B6gX8yHzaSOeP4VJymB
IkOeswm+pRxnv4gtOKqFSE2ppnNB9oNB8gGnD+o70ruK6HbeXgX6pML5lVEmuSlAErG3qmnd2mrF
D13F3RKg8IHbXMyXhHizBQCdJPpqvyxOClA3vmxNeA4Lp4Mnk0OYW8SwCR7IMTI2YmBktncXXc90
lqal6e46LSdRNZcH/JwUizWfcPZRBVK8MmaPh6gntgeFsyW8loaW7W0DeSgOrATq6WlT5kfHQ1pA
HU1d0UJ9kxtuHGpJmLyiXsw5jVPU4WO3xEKS+tDvHVYhT10sRe6BQ88/ZMiTXH+8Otm+DxkcT3lZ
mi5FYRse5qJPmr9ldICZ/lljMpTZjtsZTku2o08+SSLFefNuonVq0bJg3rqBLJBjIc4+DssvJrZF
cqcxq7FcIfdlCvxu0MThwCgLVvH3OpBet065by+1I+d2UmvFDY0p+eqb9t1lSdRrLtbm8XZ+F6YL
u39E3hAabwamPPVfcKo/TysVl+cMGatipBG1iWWaSPPXoUAa7Ybl3OLx2wOMfowcB24B2XxJsK12
Vgjo9gZ8b+vBvGh2KGsIw0lYLE5EweRwICyb6mqbDj+7OwbnVn5q0rjqgzfbu6rx/Buyu0cxsUYy
Na5kl86Td5mTuu75EE5WJxKJAGehmr15sdItEAZ/RS+5fFVmh/fSGU2k73ApXV4vYbILU7+10315
7vd1hcJ6CDCUO8uGuQBvHw5VHHqf/IBZi8gmZcbSWVwOHwgYAupUJLuTkxCRW6WdNaL3ONc3BFx6
cEWwofunjrARC8bal3Cx6RfCYaRqWa1bDDmbbzUoV/LSGbBlAWJqSnDIJm64RIJBnMnTV1FBW2yu
3UekaIi0NFbJwl3xMrSlBMj6QYDwTDWjptl+KehdCy9aHUWMQKkQXh2DpRac3G3VaLK8ecHPXoyV
vc+x8S2OZ6aWg/eORZoZt5Ed/Uu9d5g100Wl3RBD30q2/EuGhCn+ScxaSB0jT17f/fI59/hSGylj
0AnPBvWMSrdu8T112S18OxyVUSXcSI1lUfNdNZyNulaRhzDQDj7KbuKs3C+z3cbQa5J9RZj726Tm
GaF6pMhlIp5icEwrTInT/g==
`protect end_protected
