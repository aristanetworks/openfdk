--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
SVxxmCWH7zXtgJakPvQgoJlyT6g9I0RtZ7vCX5yv/ZIBEZV6dyPgi0oURWMd9ZF7mNuOk7wtKmXb
C/FhnMhG6eiN/xBsJ6Y7329Kt0wQmI9Ab1CgcWkEKs1EFZAY+5tSGDyLicxmNMKo8n9YTEaBgovj
J8O06bcDG2FmfV0RVpaBlBj6uaf+dL6IMNjm65Q+aPLDAw2PnfHVYpIg4eaVyxdbSFV1jgU/SW4V
2Sp05JSXvXs2NZHDxQ8nuN0LyaJF9vt4pWcJDc8TSb+5Viqdf7FpcPKXuKp69G9oEbjOu8/WBBir
NLLrAjFFoEiT09JK1DzDznpDS7DZGkAN1V+Zgw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="BrwufiHD+sePqX8vbAXB1pimXmU4RB5TrUzxVopTI7Q="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
p7uqoWFAGyxDwNgB4GAEW5/M/V1gX5hxiQyGddGL438oyJQ3lWhOD9zd4e+pWvUVYSq4Fwz4Ubqb
h19PliCKHwPGKXcezYxqU7FyXXqAj6yAg/Zy6fC51CpuOi5cNYzyucKj0tJ7JQWOxbYQaonUhZHV
S9ab9ZDc7iuSHxb970QmjzkBEnTWDWfGLw8cQwGl7NxitS0Obxe4stkG17GyrtqswZQfqU451/P4
x6qhUwVN/I+xcxkeL6pLeV2UxIAsYFk61Er18WrbHnoeYmObLQoPS/kUWhitNaUhIXgnkRVIiw1s
JO7b7xlcXuwc/YWs1SXO0T1KNxX5MRg1rIsrEg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Pv+5u3fv4IxTEAKMxDnzFKtaLBqkFxirip9EfF9+Nfo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10912)
`protect data_block
WueOFT43robVdVg1WflkKg+bfjOS12gbRbbpuGqazesBpFjd4Cr6lSTz6AZXMVgBHJhrgpBiMR0R
VNeHsISnCZScBa3bas1RQfNw2H2Rbqyz55nf07gRErA3tahA/HrWC4CTUef24cTHh7NYpyVfFY8Y
r3+03hsKLEh5yWO27TIdEoVlw08OCQPnAUSNTS8IiVaNebmeHCaObrv0Vi7YReJAhHKJat4Rxf6K
3Xx1kvXXkSpi8vdQ5aPeHhCWWMdnW5Z2rKkm0/K3YHxjyJbjfWNehVKBw2sw3uZCMhxFY+anIsyq
kt4B3Y9WP48eb5l/dtddIcATNjo1BiFC62IV20P4XTRrMAEwFOvHRa25mLiMccyUDaE1zfvNQitn
YEAJCUGWREZT7nxNVLdhimjlvVFH9xZ7tyhr446B7/O/lsEUrn9mBISCMFyTv3QNRJqDoWCA++NM
AVKb4Sper6L/9aBSwlaEbHDoMCEt+jXsupm9juaasnWqq3NgKm8ZgM3qvU8ZP24Epg8DOPVcQO7B
6be1zWNF8kbPniqR2BtRosc/fOYWKH6G+4/CorY3HYFG0H1cl7clhgsaKf0ltDBKrjbXGThUrXTw
1rqebZ94K9w9JwsvUccc8USQ6PdxjYykJiQQaRjh9qbaHcg9Ld7NVJGWG28sksNjQwHXBgndT1+W
0EkReeRKT76GvVtWA09bcWFh7uUvzhttbnl/Wr8lPeK6KHFbsjAXia0dbxi7QRaVM0bgjWh93DoI
psvEMWE0ejFXaAfsZOYdNXBipiZ4LeI6UrBE5UJhwHmRlD+ovpUcr7/r+uMmHeUnmbMpQcIqkLIZ
zhr3SaAHp5kHuv47xgFDjMWmxE5cxQnbdDUVCHkqhAV6LqXLeR0CNj86kFjh4gbcTZyAl37kL71C
aEvjxb7Tefv5NbOGvCXO/eN+BmscakUcmUK6zlo2rqhFXQPy/qbsZS3xth/YQfZ2ZLytQGXMvalf
0qQRfpx1XrGNmcmgjMfztHiijJCNv0FR98DLo0cm/yywxgXHH+C21EPbRgkGoCYLkcaQcHx9zC6g
/xWTX2NgHuanXUmLa/qvKkqaIBJcr7ZtGJOkUQiglczFDdI/frng0Z4wIe8jm7XFJ/6TMWddFT1p
RYer6GZPOjt+3yqZiLnyX+qs6aCzrWsawMIBqmsk/5z4pZIqWIV53/XAAOH/5xzMsrZNLHi5TA5P
HaRRtq28GNXVNHky3S42Yrv1JW0n7VHtp81SCzdxzTFEtSiZ5fviCMZYbohjpicBcG2vX98w7iI4
wUaj6epnZ8KPJ0RTzFaRQXBj9tHdfom10SMcctv5VtcjPq/2pLSoTt4HuhFqehK3A/3IX8PSyciv
0jLZaPIw18Qx0+VCuuy6kekhk4crCGE7D06RtRDzdkYFddG3l30hsGmY1BODysFZMmKPgLRkJP5o
Gs3AChJdF1mV0ChVeTwzwrf9AxaMHbNxSyUkXM2Yg9+ERK9Ahk3ir3+5G8g1y3KrqzDkGxbLoU/j
jcvGs742g2LDO83UZUyw+X0miR++cbeoDcv5AykRI7kraDukj3ga58dXKFmZOfGcRNq+nxk+fASP
Odq5QPw4NjAjAN2u7IXBPXYG+eDM+iYshCxjwWAmYhEfPEz0Jl9PKH6aavNKTITurCX0IvB522VP
Y2Znw5u9zBXhE/cKSKcFUXZkw4n5KCeyrL2kVZOoqqaa7IPwS2B0O94jb4/XoiyjeX3sKyYLYCTc
7+KvzDF1DpeSZF7u8Dm2SdU1lhrkxhRZKk9AwDvN6YeRzcxUk5/mya77LVq0jczW87+NjocrIBL9
5y26tvMzrTJTFX/qd/d8vbXnWl4Av89nX+o3QCXerjfBQ1D88dj/0Yitsy/yCN9WTkG3vkquBSmD
IisAZ76NFVtqz74tBblBsDjATzqB546N7Imb7pxeMFzoKqC47FvDCB5Z9RORAuGuhNY+80GII1cZ
WebYGY+51bqWcinSfgpIR/Vm5LwpXzhGa6V6mIg/2NcCnkMFprIBhQQzsYUoUDagAw5tdQArII91
ozxXaVuek76OljCt8jgLxMg/i3PtcDB0f91wIGjJj3xCp0HWXFJ3LZU6d52ZoOGaN78boV0sRKO5
yPfvb6XsNI2phpwh2hRNn+7cuSFjQ0DkA7N8EqGA6bajDBsC03+V419yVxfANtVKgc4cqDs0tUfm
Vcpe6QEc06bUmPB4XZIcPghTcQd5FvQtGM+nLmkx7QlFP53+sD8mg6rb+NITbUNkmVk268WK41mu
aVLzIfb/9G4OTZrcfPwzB9mFWrCKQ+DezGopAA/NQX2yQUAhAv1f/8sSMGuDqlWHLfhYj30QCHVt
yefaUgoj/SBXKKwLrZEQ2cil/GoehXoNCUSYvhUCpUT7P8fp1Go/P6JapY24XMqp4W3c/ux/k8hq
wuMUjEdsGxhtxHrO70BUY4t5mOZp6YtbTtC7YRPD8jInMwjVmFX/1T3ZKrnaGG4dBsy/VUXmxDFj
D32Rc6t3MwLbvukMGfZxvKOEiN4pmnsnzATcMbKS5l+w8pykyS0c3s2BzT8HR23I+LLSW6hVXEQr
u9O5pULXuF5KzkIHZ4tVsKYLg+NUHeO1wsUspu9tBs5CI4/1lKqHtWX/aKKUDMYjmLpaXyqegRr9
u4l50pt66y54xx9s/bYL7TwUSxxT2OjMIQXYDJazIMpWOqzISwb4lZqVAsLiCs6GDFiA9Q9xhmTl
1BnJJWfPyAOpTkXPlTPuKuGpgn5zSI5ifr+dwI5uhPYMkHvn31JXfphcbQ810A9fYcHkAyZA/fMD
g8xf6mpp6acvGr1ZFmYQtQZWD2oBq6TSUvGR0YWNF2asgxDtdFHfU7twKGtHOIFXMdqK5CyKTP7t
h6DSCnVTq5um1H21kvmOaRhPAuYZqN35qQn3Y/2H3YKJ32vSIC5MuPw8UibcFGH9Rs+Pe0SywHml
B3/pIfWmXAFIVYv8isVHDo2MRQG0BeWGYEpHFhbnSGrlPsGTL6HgEFWh9nIkNgVBRFnFZtIyEeOK
OG2NyAbnuijAzuB8TJSB2wRQqXG+zVIVoFqIVep9XsLkqi2r9nm7ZBXt5PQCMS34OKszttocTKEV
ekzw0xr1199EBtkFBbYcqvG8UvLN1dbasEIAnbotD726QJjLpTrzKbJzTcSMI1PrWAWyWRZkAQfm
mdkN+BlVebwiB9w86wU4rIlKRmwZaNVCRerw/1iGw1QSW2BcjRL4b6KE+ABrmwiDEyWvMHVgOZmh
PmnxxBGWl3JkjGfIgIOTKLg/l7xjU/n/M5ZxEyniMdT2ZaOuHE+vDTcT1jfmRTgjWYcKFi7g6VgR
RpTE/dAx4kuhuLde+6Ic+4xltJ1xhJpZ8RqFCLudm/gGN0Cb4bz0FG8bCNXZRXgeSf+aEJ8fTVOs
AxPn2TMFqgeI/KtM86cE+oQ2FyxjI0Er4MEvJYC9+G20cMyh5U78fWj8qi1JM6vLN21LjfKWe6qX
1b/IqkaogmrqqPY+3W48jxBqipIvhR8qrxAhdzOEGJ40VKSUDUj5o8CecP2V1r80xvFPw9kpuSCg
0bIWxUmj00FhQ+CQta6+vNZzh17/4WhA63EL3Lu4xF1bB9lK19dySbmUGGH6LAdnvQXJxQcqnI21
+REDwLAUK5cSWdoAHiCnlX0hgM0aEXMMoaL2D+QpXjrOneZpUZeQ2JdsRxhKl41ta7WhEc7C2Xl8
YJoXAscriL5GwhsRIYe4FvSCv+yH7KBGwJ18zKHfpBE4N7H+BS4xL0YDW21FwNu3s7oKBFyQwmC2
BzY7EfNxx/1vZ60uSHv4kwcOGvtLfnTQSREVKkW91l3SQpxNViRvD4jTB7lcaiR6lo2iSoTvo2sO
/tYJqV7gUIMHYF1Zz0remNvdb1coOnkCaogwcyMXl3HCmnjhbz/MmBMy5ufr8N4Z/MB3mFqT2+Sc
RCflG7BwKpoeYUo+FcT2H1zfZVClxSBEoqfIbtWia1cX0n9NWz06cd1vT5l0yXZrUJMg6dwA+S4u
PJVHtjJiHp73CaLa8ME0XsHXKaGiA9IWMb9B3W+2Ukzeh6FWsNiVh8NC+da0d/NcfmHdEqIisd+3
CE1ktTsEmJo9Xj9QlNwJqM8cixus1g4bTimaerO5o2f07Re2uj+AOk1llGm5hxnztge5KnDJqCiX
4i5oACQmIRMTYWgQ7p2oletDrpZwanN0ICSGfvDmGjRlmKkfQ51NmZHBiDDWRvXGPMJcE7st3dfV
mL59EpLzqBtFIQNqH4naag93xkBlQTjDDb6ET6OgpYis8fKZlWEID90WEVwbWfQDaZE+uKl2rqAR
y4rFOXB2KlEliDak2eOMxmDLsD1+FB6tSGkU+HL5cV6vYj+bF52C3lOa7ADM3NbbXrgAxhs9Lgeu
ZWuVXDtB8WReUKnbcO+68Rj5CKdIv7ZTfEZ5DS2MeZAYb34J3f0hQlZ9rGYY4fLR/JRaA9A6m8gx
7hLe3yVpgOuDM4pIUutmJASAWkaOtWQ1w6g1kyX7eFZQ7hP3rtpB7STe4Sb0hm1wsBHcjehDzSKj
BuxhJmbgz/g+OdT2nNkI5B7nn7Ha9aEiKnmr05e8FkkyhUZsm8v6DgxNtEfPozly/Paua1gqXDfy
Mle7MzbXm6pNi/pNYYZDW7daueiCu84PYgpo6B035bQ3hZKMgSMNPfdNsY1sA/q01MU4d9HnOruO
JzHaoJsuRxtbT7xe6HyhD2uVMEBTiYVrD45wGLQnexzsieDlqxJyVSH+UAeT7wqMFdw2HqkgN0uX
HI+Jt/CWEckY6h2/NUUoGgToVqvxn+L27L1g6SHxmlop6WCs/pa1FTBrtiQnXjrRqgEO61CjqtyV
4L616IjklKAJkcf4mUM9Wu+AiRw8Hckd8Yc4jaAkkPGrxXJJIY7iySvJ87OFZA6zWOTy0DixpKS1
TaIwgcIyBjlvo2LSjzPo/HBSLkwGRiFb6l8hPkkEQ1BTo05tm1sSsK0lUN390XPss+fh3bXoVpkR
UAgeRF5/EJRiYBF8QAfW004ifOI9wrex5RjfEuluO10FVpgZOZFDjn3TZzBMO+PJU3NO7HkX0X7m
Kx6ULN+jWulP5wua9GZ6uNfW9hrRsERAYsTu4aTJr2p+X0rmzM3AspJHmPkK6StXQzf2r/3ivVrM
BrDWu8rpOekWoFtXHxzf0kQqY6dIy/IkWbBhYYifyuheR1IyMktSj8rhEAryXY7DfEyRmfvwdOac
OVpMaO0G1d2bTGy1dJo4S8gl8Mp1iFPyY3IPgO8SIYEPNoFdBmRF/OOLkwCTblrSeCnWVjaUYEb6
AS5RafUkvZvSTJqoMaKrC9ScXVjgOye/rvk87wBqYG3eaIjxpM+LPMt5tmdVnvBTJSQP0LXZ+crh
zUB7pPd0SVoR8KCJm/dbONCPMcB4t6eyOnDKrza/ZDkxk57YC6ihjUL6m5sPeDgBUeS9sWHlZDxw
AqgId10pmJRlt8jbPHCxxAfQcCRL2+paH5G+9OY/xsNgyxRs64syRp71LqI4eRvXwOtCkmagdmxr
TI04UV4pPrc5cGWA/jUGYtTS57VFyaBnOCA6K7QXTxGGbcui6asczQABQ6YHxBuET9+l3HTXUI6C
jfhPwr8dF7+HksqOVZ/JTYrkzqinSnhchmjqQDD/7QCCEU8ynUgDhtMT9gwGLcl2K3x5amhbQk98
Y0bCjNxRydY00SpQXxHOx8YuCdt48cJjk6zwAT8LWo9PoVnXeUFXh1vxc5Ic/cYbeQKGSDNYLVeg
J8z7AIOw46l5JrjTAiC+UGZCCA22dUsSOAvxpPQu4t6+A8FwivcFoiTbxcPYXNXGFSCaMAWkmnzx
ObT+ujY636LvcSVeXiBm8CTaRad566iRyBoUnHBfTSvEWAfrN0I6IyRM1ZYh8dbcVQLXZHxSLMib
wbbF/tyq7/0Dc3c0mEaFBnEHAILzbD8uNiG/TMfEwvukU9SufxS8CgPqinCGlGYYjFiCYenqeUla
dmlwVxW6OmDNSrV8DCvgBe5JUiT24AyDIU/BJBVzHnSOJt5BcH/t8VysfGFXZWHSmRhMkVVx96hU
ZnlmGKjBl8NiR+smaO/sFGxZllkwtIR+PO57cXQ13JsI+Qetl/fQehvwApgm5L5F6PM6+UPASVg9
4fsr2+kVmWn9sq3BrQzZUHs/5Cs7B8/6Lo2+H2oFnI0ZYKJN2IePLREpj6wtCJ7RSk6XWIBthRHk
3Vnx9dnGxpD3f1rMK1JcBeOWufBJqan4r3hREh/5//RYMNiV5Q9e4TD4f9HIKiaAiaRha8lk2YsF
2Oahxyd9QmTYQIj7owkbn1aDe0pESZfSL5ihRs8veXhJDxaazZ0X1YCbTcF6YRKMN2qPg94U2hVF
xf9WtjBBDj1pefR2OGDnT1P9OA1Fr/6m4E3k4krFpZ8MllHg1Ur7aunmhZobORq/L6BA4uzI8Q2o
c7+xYwtDN9bgo+81dENyLsXtt81o4l+EhHsK76shMFlXGyATyoxfgrixxeJ1IYAoVS0xk6Zj62CD
wyOSkMwYv1WwsHRWtJwBHfEriOPcS5zPSm2arl8KRTSoJAnVRDUvii34lSWoaD0AjiA3Os5dB9qa
oLDKv3uD25khq1IVpoUfzxF0jDXPUPNrmyC4I+lx+tIdji7FJwJCamvdN3z1F/MdjMqsE12YHJZs
dL6mfu0jWO7BiUvDvE2HlnyLUDi/S65H6CJJwogQCPBn9zYqT/oZHwZkomltJGOR1c8JRkaJLU4Y
rpWdf4ylfp7rxuzJkZlWSZCEnbQ2PQ0l9PgDhDC72l1bi4kVfog1MSM6DMm2gg31ldFzJbuq9T14
Xx+PUQmW7qyK/Nji99sgCtOo4F5EwTW74G5bncXeMJ3XiTUtdcp5Eb0LL0jhB26b2Orx7pgy32C7
t9gfvAeU/t3Ct89SfiZPfTk2CmNH00teTZeJMb2Cd/+w5k3ALmNzvdEJqKXs5z1WWqtc1mkeQYBJ
KEs8KEd8VP5pRCq+1vLFPb2TfxZ+uKBApYRyZvTMO2VnEazVLmZCbjvkgtMgHP35vw2RyD1Kf3xX
6VcyMEDC7lGVl8b+GM8VbKGkM0JtU0dkWXJyVrKpTBApEDnMflhQd6AvMvQj4kkXRqB1IbUa2S3B
TqGmxUHZVZYxFpoGY9ZEmK67twNpJjrcWFuI//7YjCtX+f5UnKdTE9wK7PhQXAkD6EqJCbn5kaK1
hAf6BvSygl/imN6Mv9y1Lfp2QwE//AZU2zL7nFNF+G9TCD58crKPocr2Pyl++mvqbWT2ssPAXt41
CQqtHMb3w8gZEyJih97WFa1CjfUOT4tyWwV/yvpXgEyVd02BtMKgCBeGy1wlnlc9rLedrYa+2Uhc
h5MEmj0ZTrlOE8iTzisJWneKTLac2Gpo+dWMeo9kqJzxCzccPMiPbljpJhHowkXQw4F3EidiJkT0
AGiXbVvTuEUwjZGWazjeXlBTcgGb6tameuOe6DisBe1th4ZvwjhT/K0l4Nd9XQKWEj5bCmSXswth
C8iJq/lbmpgdlvsOBpfN3AQmEM2PSNAQLWB1CGNaan6CoNoSFbqgl5xesLfKtMNmS07OQBeonYQV
GktiMhBXKoxHPlMicH6P7Pm35WAuWab32Fpj0sFez4cWF2JharwwUcqfqP/mwEBGbhsZmHiIzqSs
kAtJWcW9M5SXpYy4gXXWG1C8TpmGLRVoNQ2BaQofsD/gtQInPWWmULPW+qhfGcOMXSBZF9W4af5T
ysVgf4mtPnwIPN1p1MFLnIwX5XhM5lyvr5CdvdIgUoP3XENVUOkLX12br5bowyJXKjBmSqStvEz+
45uu+AFMWTklYCRIngpH+fdjgJYf/qCVxvtE/5OvK58z865LsUHZgtJkGluguJ0LOOB4MPkzagRH
a+FEt7TdD/ESjnnlpK4M3e1+9hKwmFBAUpogAG2pf9mRElUmf/PRINXIuWgYr9eTD7gkMl6mG7L4
F3kp6WfmIFS+XcYbCFriNxP6FtxmNkSXPEe7qAL3usH8yCn3ilqpWbcKl/wuXB2PfI/X2r/ylkaO
dHpFv5u/wyhyDiZMGungNH1GOI581ZXU7v8j9cqh1O1kitmVtAhDAonrBuDFQmbRk8eQbSYMzq45
D0+zX9QnCCmeh0cu4L3dJ+cmfVGAMEeslUwMOmIEz960x9xheJ6YfC32yWAEAuwelI4GhERqaL/v
/RnSAgRdq2t24GK31UEwa+OWPaaD+FnW7WxmUuevcPc5bEWgdrstzlEWYCqOaFa6D72yfx7KR1rA
caW9YmgkxXFy3QWkELT1zujv/EIqmSiK9DXmO7ri1KHrxHRqTSad+IoSBd3Ivwx93IjW+C0ofIPb
6TjFoM0+Hql1wLHuGM2/fYA1JYS/xuXnDWTMP4FlRTWnLIFIEcWMTbQuhp2hseuft5JwZ5tUlIQO
BIyZWwgqFnCPk8wjonJ8YodGMrR6aZVfitcnKDO7Z6KxNO9h33GJawu3EpYES7wmTbAvSeEKCk3t
zgH+6EyRtAhEpbsqZheSJ6iZYtuyLfqPa3gUI/4nR7E5qescj7Rq19BEGYcwmL0Hi2SdK3nvlcjx
NF3Bb4px24mms7vLP/sw/PC03HYpEWiYa4KWRxyGAFtzyFjUluOm7Xr+RWGwIFtWg/lu77KHMplK
3LtsSc9vV1/ZBl8xR2Vq+CvTyyk7GlxMtf6RgwIzFs4Y5aJAWfikwl/Bp/VK32c1509MWUb8xysI
riUbrIZFNaoF6gArMo0hwaiDI1B57GEDZShHksOdoA5Nx47LlKHah9JQlFthMvzW86LorWfEAWAm
rn9cXCALofHs+SqhH4pXXBjv13vKjvVchBB7HFGVoltDQUBkWwqnWJSU4UzANzYteyyHKCa751db
0VhJzenpWUHCdG/bcqsY31FDIYTZV4MMsRs6tazaLCb+23nL5O/jwMUCm7X/yNxHxNa4/oxioXeu
wZTrQHoaX+/DP0lGbSiKwiaBhQGSuN5PWQ02DWaF2dSG93rUM+ydkuZl/GrwaGzI+SFBEKm76b/e
oi4/hIxJLyVGriC+gvfqoEtpwmmBFBT8BzAHGbSaAdLR4GfE+npYEy6i+7d+U3WqQNCNBN/A71FF
JfBCbSt+Cpe7R6FfbiGljydC03aM+MFpjIhRym49xgK3AuWkPjwbAR/t02+fKJFeR51CNh0ZtdPe
ldebAMpl0GrdqWpeA3ZwsBrSTgRzwwuntIoAsLYihU6GXV75RaGZ/O8S5hlgZRiM5ugHudZp4yDs
d23sgZ/7K0xJ3jOKz++cLFbSHt5prEBuqAAXiBcrKVbqd/bV2ch5mai/aRnW73GTUchCEDl/8hhh
ltblIfZdwm4X44ukB7KXUUk/J9wZirGJR94QkTSsbgsufeJE5ueqzrEajHVNd5HJhcLWxwPIGD81
LndbVXEsNgcvIlqz7veYqY2L35SKJ2Cdq5ASkmJeUNpW+CNi3SCU+OvoS9uaX9UTg1XOlU0IcPJQ
irUqxevJ4Q8XczeSwm3d2eKHWNKXoDEoxaa+yBH40iO2mHaKlqtHul7QKsEl0Jq2IDE0gwVoPFZf
YXWNvGMVNGENe+h440n2VMpyjVbCe/JakJm5FrxFrpdKtw3O22jdAqrKTrbP4JE/14oUlA192GL1
2x3T8VM/zA0wlUFfH0xKqM8DJNH6aGsEi9O3aa/9cQw4GkG9hKRtujCvVsfGuOfG8exeSh783jGr
8IOMCzuYZ6sg0dGf+3vfwoSklRhmjfczWklX0NgSZNdfEjs6Bue1F/4NUQE888w30xm7d+/oD7BF
VjTsBqqKREaouulH/alvK8VO22LJOxFAclw6QBwaTzK7z5+sPBvHEkQc6m3UlxJOevn+xoDCw+x0
SJDoJ4cTdPL9mkIQzZt7l/kX9jbxhf+I/wAyzGm20OtKnS03u7ymgDfT9lvhx9SFOMelDZ/JKt7o
b/KekhomhbubFKGxNZRNm8l+di4AhX0VrJAX3QSy/raGPZFRF3PSJ2RUBQidQhjR7GyjMTSCMybj
0J/rf91IA8mm1mK5ucKtu7yjQ6ngfBhEhp58TaM4mB9KdN7Gx9uWDlPl4CIdcZsu9pb3bz5eE8Qs
jkgemWCgNTYdrK6kAFU8b/pOq9auC6UCZPqes+s8vlR0ww7ltAE2bIvILhIW5+SPpMFy/1+0e6zG
kHzEaHdoURjzMGxApdgw6l0mGAGoKDF5CaEdO0nS3tYDpnrCLZbH6819JtkIuI7cd4BRM2oSjHmI
e2r2K2w+jj7TWEWEhAebWVPGF7UVANbnNS5r6r0YFfYDHdYJOaFcC26rVDhmkFyCFNfgmosMs9H+
J6NTwVt/zKASaVrJBUIeSk+Z4/JdAVnvrbPW4sL9aFHNcqkbaBWRSQ+IHxqULb8ZEaVzAvuVvW6x
oz4MVaOzX0KLCI8F4hQXjxbJAVxNXi2PtrIWyAYiInCrnT0Y70GIPJ1GbxHbrldkgKI3jNA9ShQD
6mGUIKThlUF0uhimZyUz9ty/XKUDLhI1aYNpudtp4R7nZO6fL/pzFs4Ligs+t67xhCi6B7UisgMr
NGNIXG0Lphh6gHUvWSeI/HMtSoKlJrEC89MTt/fptFjpLP/hFqKIQO/GBGEVAA4xnG16i0vEPDg5
LFZkbfCgN7GambZ7ILwc8m6+JktVsSzh6ajANRRKsLZIl4/oT/COt65WB+XlSxnbQhL946zTbM5V
tkzdSJDshwo8v3Ew7WvhmRghM3T24WiYtg+jPzo5YOCZgowIzCgMHCZ5vNtIXAWvhPh2EOftaZdX
E02jxJRIy2dyx3/VVHd7GZ3e2HYxTavMJZ45dUfTje/ZNbBcIgjRZduaIy5NwDxhvIHjMnDqtb/F
4DeM7cpv+16JlQ9SysINONQlFZHIgDgGs1jFVmZD3NhDSmOZxHtNFPuRSrfvDUZXGD9lT8jW389g
dYM8k5U6OwvbIxi+pCzqpoGfvILW4M5J77Dj6wC8oVW7w/GsD3DlQNZmB5o8NsgX4Ny9qVdkjMv4
EMr7L3psr87Ca+Wfs0KiN8bHq5K3NhXOunPjsPl5eSA/B7rJMIUUQ9WmXAao6XRYAsHtfMlYJZFk
sWrjdSs0j9g4lUZDVziUPNRfrP4MnR234z3sqscQnuq+Ketl3NPdP9a1AYLLRpN/tZFLLsW/UzC3
mto9hDcr4GSG1XqHGP1zbZSNqMV1Rn/fclK88aGWuMAqx/qqvsh3BDRXHBFnMrxyDYHprAwXkgUm
xkF1b/mGsnngFmrYFAmqDoF/si+Cl6v8GkZWJuICxxk/qtF4qgfu5wTYR0V/CqhtIcjuHUZqcLmr
3koz9aZ0JRJcmSCJ825FuSKdydV6TuucoZPclvFcRBCP62tl17r2RH8733o6NjwbMMdkMA6T7k0a
QXizitbTi42bkSfBwF4ckUVnfCaTC4g8c/sdHs5Mukm5EpsZ0OJDBYP1Yb8eU9eWPlx6VJ3aQZtT
bReeI65DcGYd5eO8cWIFMLQuueYQappa1FO1hACotgUBssZDKuLdUtrXctoZuyxCNpf5UMQxoEHV
6ehyv5lYModJPGPOu5eo16WW92fFNBbAbHw/0yoRCZ6LRq2kgdPKmp5EEowlL5pcdeJs9E045FCj
byYOWvJC3QMDJCl2g3neThobbhvJg6CT5KwZ95tPimNlISzFcZrRrDK1zfXfFkpQJLn5CzwruVgO
GcRHvgto/DXcM3V1nppCzAn7U6x5GvVKLwitztHNrtAaTn1BpcI13Tit7bQQ6wKAceu/6WqQdTJd
55KxgYgURgLHAdb6HG+Jh5KDCMGjcMCkyqxQxxjGqiEJBB8CaTCW1YtxI+ZpxsaJVayzhIONN2Aa
lw+WOaOi3Qrgi3WOBBBRxz+BIcAgwm3OpVPy9ooelAHkCeJGDDtZGoti7kMmepm1ZsnKcMh8+wEf
hxEs6HBiU30C7OvQzfcKClonGpM+s7t9tr43heuqnfzmUyPisUqgPIpzk06W+qehgSF775rrN+yr
pZAnRqXEficcYGQbBhNagOpzjAgIPJLNYsIK3lrP54S3Pb/bbfhEvxk7VzvxyonsSCtb1y3tvikj
7zTNZzaLffeAYSiITYFwcFzIoCeq8AIl0c1i4Hjky2b2Njg4cdrLVw7xrVtq0eOzOYIvK2yBVi+7
OH3SmaLfCpG+j78zt3hl/Np+Ztz9c2uIwjBmjoZELEwDjPWROgC37rrW1rC/yQS0Ji9pDayJYO0R
GRh9nc+dXcLo5JYCl44tXW63S7rPaQLIth34KwVS55b6SRCZkYD3NoiRu0KgncsBYb2EQfWzh5w7
19uuj4mf9GwbyPW8iLRVE8mGhLwc945piml4GqLzq4nEAApzULUUV4VDbxEksTXkZFlUzOuiu2fo
nqGeTH06soJ3Pqkfe6uQ43aVbwLPBJ6rJWog+qSAkx52+bbiNBRWXh5gMphDNvkk/yq2Ceu0e+zW
WL6p837saPSbHndhIUhX6UNRRNlCWZ/d39LT1lsbc3vNFu76HXWyagd9Cr4hxGTZbPfML4UVpehe
nF5UgZpzNAeDZUtDZlztCzcN9U5BiKeDiDDrtC2hOOUl9YIem3VhnYA/98+HgB9VagAYzcx2OQWE
lWX0y1vcvJdQ8VKO8MFRyxWJ23/r3Wmya6fz8CT4Nd+Wg9xiI78TgIR6QYnnu8QOldAQoEPp2idJ
DW/a19XVcKjr8eV68ggQm9FE/aqz2k0Y4V/6ithiU/rm5K7p0xVc8jlpguJOLYEbBMKoytIr2RJ+
e3TZ/hceLWYORr7p7skZWkeC7XXOQ4rLAiHvGbM1mBS2gsdr6rVPPlsMVqEzWD8xSP8vTc7XlBni
JsXjQYiRXn35muzCZsXPGbHop20f4K52ykhmiNhhB+5ZyynPBVoL06NLF+k64nQnf/iLfpeq8VgM
B5PD7MawISZgtJvk+FXkHlAb8Y12HANp2PiqMjwG1oQuFS4c1PpH+JUzUqTSbMrBIqzfhb8HpdTC
VjZHJuny8xKIvz1ahpyoAiqgOC0ZHRnE9C1L8ZShn8Uzt2zVvSQ0tUvCL3cNrNqMDPDa5Bfl4V0k
MO3lIWoLirfYdGjFwNc3KUBUt1h9tBWARJg12mOLg7FkTY3P+O3N/JNX5FDprWW4VJppaonx9O+0
xRbVTFThMzgUZePhXeJBgyYk1GTlKy+3nxhTrOlJR+hECdegpGGx+uaNr1gfngV4escLIhoZF92V
A7NX1pbpkZssB767RSEaSm6nzGGBbTsV5idzC+aKc9LKdrXkv7P4EwnCUYO8rK8DK0c4Glej5tEG
21xUgeB31acjB1fos6xONh1edHu6WuyTRzmat1r+Hwfwdjx5NtrecdGZu7F04hUeoz/MqSbQkube
ibOKVluYadn29q3TYRYEzRmOR2paNU8ng3VJGncZZxzU75tBM9MtGZLnQh8woxaZYFwqOZgDzpEw
wYtzZsANDslAzV76thaBysNosPiS1pOv+9X5MQ6a/fA0AwVsh9Gqxmo/29/iF8O9UXiPw0fHH2mC
wb1jdqMdXm3/jxlUD4LOmz1oAm2QSgsZFEHdCcOnRKUAvmWeo31/W/+QqJ7dTNHQB7n5HUoqOmRf
1mi4heU2fuyhKOlzpfWewYTNRfL9/Dz7fMC/HcgAaMybfxWOzxTMWG8W0RInvb+vUYISf5bjC1st
hxECkDid4lKjPuicEXiyuYAcHJwfvjG/1HBcsoavFXGC+zP2RHMzhWi3SacTOeitgfxSvOJd7SxA
h8rMlAWWmLWj1lKWWKAqq4nE4buJM0npgyXoQ3Yjo6tQ6dgFpAn5EsuoDxekzwlYn2ZT+aG9bvtC
wcoPtVcPILiBb2LcHRjnM9Vk3Q6k3ncZ5H7pOlFJcCOl3kLsjQ8bdohH7BJiTUk0Oexow+hFKMk9
TUTkyagwF1eiYuyn2Bwa8EEdA+hi/AfqcFr9prEUkjPaOturo89GrUY6ArA9jNMHVN5DH3W2ykuc
VklnEk5ir6aImoN8ix5y1BDHI082MMSeDDFXbzV/Eh8W+QsrSkOaJkPgRapr5schfTUdna79uFVz
qQsAcqIt47C7WdRpu/map7JW+cK5SDHIkXkLA/ENpP1nwbFj+jvOzNHIo5dv11Qbpr4VecI6rNBT
GYztIo1Bjv0DPNDwKoQvaSNr7Y9E9EGgZ7RiKnztDr8dnrNZgJN/YBSoRnGCYhJrvD8nTpCI1S+i
CRUkgN6I6UW1Sc/HM9To/V2iZwpvMlz8/l7EVBzhBDtU5MH8WuEgOH6G2dhL7NtVQ/XuBjpbdPqy
+Yk9xF8k8lWUJezo9JcWVyhrSvl/sjFXYs0OK9bphjyxiB2TZwtvlJH4nheVlAd93V+0z0QkUhKQ
0Rm1VLC+PCLmCezYEraV9eiliSQTkt6C9n51a7L6boe33XdgqVk6tqEn+xtSzuYWQ0EHTFLSOJe6
7KOsc1W3gWfHsoFqyL5T0nIcWkaWW1hEShxbQiT6Nx/C0oztRFcje7QqPIELMzVlwnvTB2rfv/ct
CoSPklPFHo2cBuVbbsKQJYtXKUglciYrVQ==
`protect end_protected
