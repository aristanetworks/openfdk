--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
ABUEhj3lHvwHJ5jOro37ROjPXQpHv7kcQhpNaSz+jZPTmeTfdP7ZX48yuxEGbVPxyiQ7Ndb01dPE
KcNrp29b/DYE5Lo7CnaFwWY+41B11Lxi0R54l2XOhVy6n+sgtuX5d8lTYYv7oYSvU8Rxnvthm5Mo
N0CbFAFFVujwJSO02ZCFXhivTCcuZbnGDxlqqSNhSmZbXKftVJlNqUZMetvUzL5+Csp0STa5MUb+
U3ydYb0q8mFEhC8oTnAKU/c4Mi4eiEDO2qeRwUGJ7R8K4xoAzlom4xAL2wwev2lyrvaugcrfNIcG
d5nWWbht7TsGGzpmlleWG2pYO7kl9wIo/UobsQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="5AZvRmUVk321kzzl8GCshFVylPGLDy2i2J0SKSRGrO8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
mY/50QXj54/tdcxHxTNy5hX7N/CAS1dA6sF4KwEJZ3jiP+VKBsZ4ViKrYxLpYqyGzWQLDV4lPoSo
HnxbSUlKjWrsMmrfhWXn788W3b379RhNH48RCy/7S1L19afQep0U6TUcUZ0vpYEwTgFEFCZ0q98d
zCJY9xYQsc9fcTmom2/6xU/lydl0pyIkT/pfvAdd4rF3MG+20A32Je6GAoFZr4X/soPebZwooxnA
XzCzuABP10OWyZDs4ooMyl+hfWwVG2p6sJIH4D+HgGg0897zFuSwbuOjC7hTCtbG52we5bB5TiZU
JM672NFo3hmFFyACcG99Cr61CPzTNaG+aLbzJw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="sS48wRLaXVGoRY9Kt2d/HRRFNlQcFUT+By8EVrxAtSU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6032)
`protect data_block
EN7HXlNeLYjVRmNK1zEWLxOIjjR3TrZ7S94ppTOFvnvqi/WlQSsuiydG9od5zK1Nne+o5/QoyNLw
QJQMWDFxMfmI4kcn9HzmZHU/eexzHhsvHVO33AAWyskrDtL8cuWrU7gBGrgpO2Y0Vn8vwbixwllP
5ugdilDK2hFqqSEMau3dOKlyTaQIiWC/KRBZRnB1BXQtcB9JhwpSBjJkuDo4hj7/FJINXLwvU9/v
JeVnVNd8ju9UAJwATv4uNv1Mz0LVfxziqlpZr8cUT3zfQ/BFiyvapVbss2qvNRJiI5bZT6dEOo97
EFmIRvP7phW152F2W1OUTBF60pnWcVLDEDfMIIQyQexoPimKXZScxOYXMOi4j+nVAOw0PKiL4Ope
9qhpmZHCcqREDJGlvAdod9Q/nXXeYsq3Jg53gGjH7Sr27IKUA/RRv9CDSjWcx5wL+alyzTtZI0sE
LUk4qOJb6JxnAYD59hAszXqQ6+4A5117lMop/5HjiMhitNrL7tyuqBUXT3yhv8s7ey9tn/qWyw7H
h49QtXagLXurEMx8x/i9lTB5530fceqZp1rYMPsPcNaEc3adTkEe8FUNRZgeyows8aBXoRRVk8Jx
cT+MIkVPgnyqWvWJg+j0O69uohp9DG8KwZlzFKCUZr9kwJT91gmgOgLNnZdnNy3KUrBDZChtdDFZ
PaR8cxDTldwr+ioGBhm9/QUtSCfHB7eHchIkexCALOhfaWfApdv6V91Lvxo1BIb20uBNNm2LSwcZ
254fjATdFuDUOudU+KdF0vLqcGRgwqGABbcygxiKAKCXuSWv+Db1Jdu+qr7ll/xJ2k5vGqTrfzw0
ZMuFe5vEfjAOve9pscBCZWJSBp4UrDqjWldF+OG99vbV6cE8gPlxTso+s8NJqeoVsLk70S+SDhGq
KVppEk+e0gc/lA1+WWT/DMpYO42nE7XL/JXUqJbhl5WNHbcRp0u6AUZbAqymbVJeYlqY7ausvXN0
EVTKRLpN5of5tc3cZVQ39+dnU4KISSt0cInJj981SfoG6g7icLpKk3EWpTmfD2IjZSF4X6yFlPwi
f2RphToaDtT0ZEJwmtsg3wBVqGqGkOZU5qxK8no5gLmwN3sGYV4G0uRXE3ui89A8nI7oMdIlsxqi
ljfGirpv2DEiS0W8WRHbh73r003KhiIB+1nAxiLiA2PUap4irGNv/q36xh2PgZFPMidOD0D7unWx
bUVWfDcgajxDSxDvzviG+XvICXvHzIKaVB7iM1XI8tO4nQzUp7iIv2l4dl7QM8VM8xpqCel3JB15
Oyxsyb477k8BJAicuhUejk9Kdor9lD699XyX6naTonxcSnSM9OYfvY6UpUNDla06kIizHuz8PWgz
+ZhwwtKGlEXr27kNlfrLPrziXcOF9HC0rQ6lQGagsRgCsv7Bz2fV4D0cZlI0/0N16x5QGcY47620
Ttn/VWc8gQ7+fhFc4noWPoV2ZqNtCkT3tWLL17igFP1XLklr4mGvis8VPE3CN2UnvKxKp3GBUqWy
8rjPEK5s59iXhQSi1HULiKrebk0aN9bkcFUF/NM6PTEsnNynUHtTxc1nZwW3ILHktg7Jzm/BQNca
940vzcHgUNonc8BG+7T6TILq9/vn5BT0OrAXcd2/O1FvhSkCz3Vp/54VqeDBLdDnGtP+Zb2QqbMT
/HXSuIQdn4lUcMzF56+FC84VNzC67bPZIX7TowGCqwNWo5b1fVQWC2l/hGiCQfLnug+/y5WNTYZx
iuFpQ+KaMTQWZVOdj8VpXQxrTpXhMYNj+P2+nScpR+T4uFoJfGleiT1rVPVEFn38r2LnaQHAZ1fQ
/vGpBTwQjIG+MUT7emWGy/AyWxQs1sPkwKccLqQa4wA8XwpKEdg+8ai5RodciQ1LrbKKg5asqaDt
ht2XZicMJr2IqwfYAc0jjAGxxPUfWLMTYjXmtHbaD2M0O/PZk7ZhKOlaZC9L49qf7HdZIBFAeOn/
vp1BmzZBDiredZZm4X3Ahxl/P53qtbgaW5cnv37tiB6PyjX1fOCYcBgxlLJKbDLlpq0HBIeZ8XaQ
WlRkgtZX2AudWv97wrMJ0ruCmYkdcoZMVC95p1pEXYA1HLV3PqP8hY9HbOQltFsF0gJvomYfk/FA
Ie+Et9PeEcz+LfCEURB0gIz8oGsEsPl0Hqjrdz6ORfmE15oLOsd5uDhZbITe+xk0qxmdO46JeZ2g
Q3r/bvHVOwIuG2L+/+S1VUL5ShVlRS00FRlvsN5GbKykiXVYxTSqWXTdInTpAy32QegZyaEcZdll
ykpCEabjauaaEtAK6Ko2FOWhPF7ttnUyE9DH5zZm0UpG1zly04rvnfvnqkEhy6Um0T3P8d/omRjq
5TyUAezDFTmY6WwLudfLrEm/ndTzJHChAl1linwKjeTdN9azVu9sB8Dlm5fG37n7gPKHQcwSbIb+
hQl1e2Gc+xMs33V3BWNUu+ivvsy7fgTZch/XGJTsz3ZOvODPCTvUfHU4yCGQ8gAAjipggJUD2D/T
m8F6FQpZpdbfLA/hUSZbFtRmq9MwplnXnFxaVjpLCDyNr+NOMDkvmOIyJnDDNEjHEOVqmV4syxDn
T5tPIlkcbYjhzB+iOhgHKL6rBWdFQKZCBWxtmF07JUQg8YDK0ZTkByPAJQMXxs2oP4TOorFvdbo5
Vw2e6KUC7oKlBnnmM02/oBPL5s5WxTR8pByIwNOoRVviVHjq8bpEKc56rdgAV85djf8bUMhCDzGa
mxCRTX/Maf6YpbyT/d8IC4HYDepOQeP+886FlG6voxiIBz2D9rwQJUya1Frabg9HN8ptDbsb0LJK
J7GSy3rjbkFDTELcb/RTMOrUruFhD1z1bZ0eGKxIRwPqiEzKEuQEixZTSljuWaqvIC2v/cMoXS4r
xvTozKWqJcc6Seg2Hj5gr9P1yrFCksMI41GjNphC35czBNhl58rzGyIK/oa2cxuGGdChBr1HlQjH
2zPUQYRgPRUxL1pE8CecjMUrdXLef7zGEvwAxwHNMoMn0ijsZ6BqJRNPopUzfbxofZAvcJS68O2G
GKZaIZHbZBjxnuLUTpt7K0JwSqUL7/RWRs4GUcAKw5c5hBCE3TxgUzL/xbqvchWpaU10hOfZ64GJ
4A6NmqJgche2KyfVQZdNIim4WSq5yFMk3atZgwIn03JLVVkP9LEd0wMzjwYsqxvRfXcrbiLjqi3r
MvkI5OXrDrHor9MaAHFsCXeGh7iECad+li4KjyYtmCwmrkH/hT6/1TBgckPWxXGbMysW7yWte5kv
GEqSl0UVnADvwIa/nkJ49IRkJn/qUAs45MEXY5DkbctsBHvQGSp2I16Z7/kkeLjOpHcbzxEhVzIz
vfrs8cXKuHE+bdgCPH6uCCL6gNKSn5DOC1sHBhXvyUGpHLC+o4GYpQsjcf/SbRLC5WFudhVaKoCM
dbb0fjQewor9w73P4i4T80aS3iEwFIlRaDioHpIiZzCTUlh0OzMvWWSGljsBFOa7CKP4udCYJS98
w/XrG/Nq+5yhlW3ui0A8aoDqH4WYg/Fx5lYlv5DcTo1fvTRcyGe4Cit1gvs6Yg0Z9VJ1XMNd5i3i
l86t8WcHdCyt+sRVZKNfBvm522WMeqX1XFOiMBfMD5GXzOY2bqO7B9gYR95RUgUld11JgORXPXdf
srdrzjh6HArwuqdMggde4Z0OZ7GfmbUA0dMfcSD7S5CHdNxzdysM4bO8Smi19Ut0o7B8XsAc7jjk
sKO/udToHZVONwiAEV38F2I8iugKYFGX26kE8gc/lxpDKcxAxLKilqPF/d1A+wxBqqwLtqHvPcrV
Z4x2t7sCqpYSJltQGsws7WC6d9Jup8r1eP0PsrY/HtUWcEZn0nG2zWGx/XJtKIadJRLBNpjeUm1n
Iq5vA/F8kmwjkivpN6J5Y2XeSS5dUEkF7dTkZ+Dqgk1IOI3NzxM9wPynXg1OKzBqmA4E0W0ueJ9V
9FzI2T0sPRUp0JUxU3hX1WxxR6OPpDjHt5YZMXeAbzSGQ4jI9MKvlnHJcOW3x1FQZBjuxNrXGmMD
y5iCSORQvh4JpMFPqNIaxh8rs80TQ0NNqQvcAlqZxFhq+Ce0WDEeShDErVWQcRnd4cedawIAbVTZ
U28JyUUuoxS/p0h8vpU9ohDpo/GUbJZTxazBX2v5q+jUF6L3sIdLGhWY8Xx9QT7qEgSeg/MxDgTR
m0beQ9w1SVGtVgKA/LtuMoHZxFRDAML+yrzvFdBeKMN8QhbVzMk67vNCXKTWztR1u+ww1xdvgcla
LYAlH6EOzaUQ+hXdsGCv68GEgJJ7Ht7BPAQ08Iy41SeTgvAilHP9dkGSunbZBNY9LUh2LPno7izx
YcN8CI8qyGytPNc2h0W2ISinvqB9c7Oo5je3z/EnRNLV5DQ81qAsOO8HOoNsMSs6z9fVU9K5c7SG
5huinoW2UAvyeQ8xYNSNrILOS/XY20wm4Odct39zJOBty+4IDqViX5m7iYdJjLowdV2ztt7LqSj0
XDi1MVviVqp49ewPfO6nr29nO/M1hh+pCI5Qh/b1R7uRwOdAzoqDFCUavUivzbRIXp2sXkqFbYBa
ymum5oy/J4VfNb91l//91nj2qiv/00rLNXgNvbLdLfH3B44vYHOMYUKkzUipKDkqdqXZeCQo9HnK
iNUmLcFC8QYqr7yg6RA+a7Rh0Z64m5t5FrymyGhGXs7B2MD7j0bReiWFPZVqCWhN3Fthe7ssHOhv
69q9UGY2jUNN052RYq66S4HV73YY3HMlC4a9qlgg1Y4dVfXldXMijEbZV/0Nj2uW0Zm0Rat+KtYi
Kk96ADLbtc45OHO1AjQOmrMixCNjIc4cumTEaOQrUXuvOcFPJixRM18ko6c48YSw1lOfS/r6+XC+
o9ai0YlkbMo5LdFA1cb/SNJbg5dqHnjTJVYf6eH68wYo7AbWDd4X5E8GCDf/sfHy632CdEQqvwgb
hk7D72dKLaU7qesLaOXdfg5TmI2IZq3OFWpSJF071poSmFglCh4JXZ0WKCOqAERuqmbbQpTePzVC
3BH40DfI7nrKN7TxkMMLn7mXzyoQ8nmK5YZlDkIzcbBrodx+R/Fxozt4PdckrTpygggVN/ClZiAq
bF6/hbqkR/2qVO1DRFbsnfDQpFzSKqXqkcDocIbV2DGljQAPOAI+Fu/FsXOIAfs4WDLKpOeA8vQy
sXZcGLVakSifL63nz1ht90KfWmMY3gU4wVs3XdtOHrugIAEgOVSF+EVgTtfIIeIpTBIjVRF6je3I
7/v/gEcPyNsGwMsOO+kMPdtPTp7rL8lQJuQpjQsSganDA7coim7IOKxzU16U49m4X+UNz6qmsJgB
VGk8/YXA9UmqDcE75MvC4wZy2zJk3ctGA7b8TshU6Ly3uJ3nLlYVrfoKgC3shRnc+FkiV9rKsKCd
OfhcddHDSwmKZkie7ThOPD3KO7ouE/RTAEb8Terxy8+p3J78OAlaA+GutskxY0F82RcJW1cotr1Y
Rj1aGlm435wckT2vRPv/d6KXPwNtELMFiyuyYFMNOJDV8hb2Y8zDjiXc4MaK6DnUymraOmgBoD6E
K0u1PmAUY6eJnztvJJrRhsh6RxhJsBteFAwpumV+ZtyeL8hMiskQsCCAa6HiZQTaZbfodTnOVciC
jxbkEE9bzEe8O8g02YkovD5c0xTdSb0BVX93hVtJRqx6OgCFJwIlMBY7WuP4WEEU1UOFtTpauQXN
zB7DJBKaoL65+WguchnxaC1nMRVB4YmI0PNUgZ2w3II9JMftpycq3vnvIklT5ffIk/Uao5RG07XX
30jyaddgDuQBTPOcGJhN9H5YiaDQA2WuAG4yfgeyc3sEuHQKO9IbRzTSKKn3HHlnwGmkpEiV855c
aaba5sF6MnKL/DdHbFS0qLSeq/UiL8rJAsZUsCOwkvn1DJ02h6W9LlP8BoN/WaltRId7zM03Sjpu
OSB7OstLUxuTqWyI1rLrEkq8+6hndIcbZfFHhWgOWGNk7yMbokTWMMe2DFb+yFylxFpANKh+Sx3m
RtTyloKxxQnSI9trDBHlcGO4/VuaYF4KSfhqNdUcSAPZfeslXjjPJ9jpA3MKMILunlCYctqlk2oT
jUIzYlYUTfF6SfYAH9nVP2MWKobZbICVdIiX5FcH0cnkd7li5GEemtzfOH88KWu63rtkWZeHFItj
kMqUDAhPT/C3XD7iZ+7s8Ci9iURvwRtR2gXHznmmRfZ4zuEu9Bh20RX8vR39gxODo5IKsSi0lRGS
n5oY3/lfxT7Zm6gJuP5Hk2bUNYzsNGL/g8UHjOpSAO0AzZ7TTXyN721yGQjUmXagtin/pP0L03q5
1oTvXIWSuZ+q0A/CnMd7bYMZcJQNwRQtZNlRu6StdxFrfl/pVerA4NLNns1kZjLpXRRNR/1DeB0r
I6ubjlBTAOwYx9cAiB9mFtQh5pN/O8NKidMw6lnj9sPBRHehWXlwB5EXqZicU5tHCPwG6Ojuokce
aSGa4VUqoSXere8CsMMtiv4B/jtbv4lGVhmJTkF8TYLPf1sLIp8V5ZxGH0Ljgfv4LYv9orXwEpqI
qR1xMMa7927ImGtugy5GmKG0lFNyWYau7yxzwWBnqeck56cNU6Fp6t+bUlaW64+C2+TpDpZQAFWp
gNyqCSVpYz16LXOqVOHJgFCJcSYL8v117zxZ4hsehcT0HZq3hSZ1jPboMMm6GLwWFVwYTY3hYFFS
cVYvtF5ssDUnNeKdgwSVMPBry94WQHnTLFayqhwpzQkEgffaQaKaBdH/V17u/ms/nKgZ8ujR5XgI
RcfqfOsnbPO+uBsJ71+fAo5M4MT2cF9TMy5sJ2hx7BFN3TT7otYLUv19482zaCX9iDjYC7qgdPLW
kGWXoLKUVKnXtp1amhiEUtg/xdUkfoDdH301a88dkWUfSnudLNK+I61+EsaGpaiGfLH5/8BizK6C
DI3Jcd+ZfIxK61tG+meU25yE5d2+i43gCgy4qEPahEP6xf700jKn05YCYMNWuk9lNvZZ+hbCqjte
GR9/G42weSQ1C3AfRqcFA8287ni/mFG7XNnsROlZ9rzwYyyPY42La2IJAI41XOV5q/kQTDVb+G0Y
eOk2L0x6uiK7L4zngpjDfT2Qrbq+wSHRNYDCyAoK/2vJmUczCyDBHzmMDBO0C4sV3QSNKTAedV3g
n1ftFcHkOsmmtRp7X0zoz2834DeNIExzMEXBH7JMocGEH9qpDr+YKwen1LZ1aIvnxQANCpgcAhjw
IioBppyCOc79RqG3Y129/Z302UY5qzEiHKzhVIIO2Q9mloqc4Z1Bc1YMrnjV5z+gWgYrMa+GD5+g
duWulA+9Fvsaft/eF8n39/nEq5lXpA/wFIdWDoy59rz8iyy9ez1+tircIPQXkqz04mgWdjq1K+uC
bQUuA7NkrSP4zXDfQC+pw0VOo4MAhbPX16lSOXHsgtttZSn67BQwJEnzhwAoCqNfTyeUZVqcu/Cq
GwaSjb9DosjGHDKKYCQL++IGLWwzsNzghDW7+bNp9GIahQq7nRvrXbmDchcmAoEa7e0TNLQDJkOQ
D38BoSh8hU46jbvGISxOaH+Sri7U6+eCg4YkIRpbFTmOU5xPzVwH/fKMJWIvoFFP/lirLZCB5Wsx
yriDS4hbAFDcM8jAgjlblhZsVtdox3qJHHqrDoDVk4nz5kV2w65U28sNYXbUGkH4xr70qeJ99Jtc
VczA5yZveRyBW6dEy8vPm2DMnlxgL1CQWwXfPt3e2YjzsY90Sr0zoUfqCV/DxjmJwj/Ab/WNx23o
YGzXV1dEK7JZ0eCkRGM26/BUEPEgHZRvSK9uxsNW+AbNsmJ7bS3HDC+ECCAWKS4OpAZKMDiiTw0A
8nOh11ZlhPm14ocho/Hf2Nh/Y1L6Q+7dzcIXrn+67zOi+E9KQ9wjEXSFYPB6UPjrks7uBdcKfk38
I9uqPLJ+K17H9e02fEZHLkcIhmWyPA7vcYh2seV8Wk5TH4rF5+1TMg5jFlscHuxC9dOeuqom6cUb
VcN9Xo9C48/KhDZ75QmtUKYPpF3/Mc5CxgU1BVb1UQ+OnIAp/QFE2Cw5FqGqHzE=
`protect end_protected
