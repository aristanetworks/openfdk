--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
OULLQhqnvXqPBRWDVGVZsH/GkNM3pPCbabAilL1Vmic+ND30IMekd/q53MJi+Yf9TJ9ZWnl369fR
MxnSbka3BAMeP+4oS4eryX5vinzTYbJ6ox+J5eUbanXKGKrIl5ZLQ1GpoYMBSkLZuPgxygkp0vCx
Gz8OKwpFawop4RAUBZ6QV12iLFUfxeSC7XHevjsmkJaHUuO1d89Iuuz71oxHelJLkTZcatAxIT31
wQwRCUJKa6o9IBOVsVK64g4dxJBD5XXs4kSTFdKJbmPzf+6UpcVHbhjSW6jQ+y6S+7Mq3ZJtovMu
aB2Z75ec2cOdhlCYjhzaXJftbyln8RYxIHlGcw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="VcIotSCj7HGGaeGMuw+1U0L3gRx6IRg4Jw32Ak4qTZ0="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
NyCfq8VwO19Sc3VX++zFHKhKI8MwmzUeZ4yBczvP1ZIO6LDo4s/gWtICb+rn+Xj03aokgr3V02C9
GV19OaakOSZl996zTlx00/ke3eCnb4tasxHnHWh2dsWBe09I4u5yClfHeLUgbxSkFkBm9GIlrxmZ
MZvbExxLyIPNBqcNZ1ohUFZoGoPM99cnWCi6NKjhc7hwc2x5iJWqHq+Byts7d34013ybv+cfu2ai
Rxg8g0klnHJvvirxj3JjPCykYiXl1qKwRtczjd7gTg/uBsph4kiVF2Oi/vl8xCYOB61mzflqfJpk
B5HsgDD777dIOs9zDqdTEOISoIFw/Pe2MnxvUQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="MIZ3RGK/BULA5WoCWz4BnmZgn6dGJJ2TyNJ38OwDeSQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2896)
`protect data_block
DIS/FAqv/PPLea0cJiQv8QSZsK1UjWvKlhJlEGanuB0iRpKcMz8pNDpSgOkTkhzVeOX8hBXgbZb2
ncVW52XyMgOw9b0fdoeHo7wmTGyhBjkT8s0h/p1bR9nzllR7D9YHH7exU2O58nelATTDlOXZLLgE
+Vc4OZ6lrTWTDSEKpTvw+sZWEUcbdy9/7aLx8X67IGugr/1aCdWSuHl7alm7ZURroQafkaG7I043
vAD1VbJAD+vLAWrkadU+jNzRAuwrRjfjkD3LssLmBq/1aS00NMx9eqhRoldksKi/iav8imqdqwnO
MRpJY2IjLMhJYToZ/Ar1dNWMaJqxaNfQwp+zbZmJdgvpDBFQZN2udB/7gXiNw41wETC2LoMwv9xD
4e6/H5HDN4leI8kJePHVygnwX3b19ZZ5YbopTDXhNVqiAvvIQfPRzfxhqCpLRUa34Yh5XJqvRku+
n4xeDWPqAHxL9smcpXRdu/lI2kLPZ8sAvA7BlCoyqrhBGcrHW3O6CdDCJKYax5zoT9KkDTFlhA7Z
45hK22Vcv3KjMYYatqLGIpGVaE7tKEcanOuyi9q2m99/O9DJKZKyjw5fTdLSwEPuEt/0EuR/jpJ8
gm4d3+VmGmCez/BeLq4D1yRBq+798Y2ZOYI2rcvO02ysf2fUXI45YmbU7LXL2XID5iXiGMKsz+Ux
03+1eC4azibEJqRQl4VbrzMxRqKQ1PGe4qhcXDh6fyLjx4Jpnj5R0n1+zbuOSV7BF2YO7q2RkrGn
xU1e/N8RcRCa4rYAsLU6SNa9sNKxNkA4aqO+0qY/mdhjv2d/z+BBDfWc85RkYIbwK/dn9WIj0DKF
l75YYhkv7GT6L2HYic5p7/0Csikp4YEK96ltVupzJXNDmLGMNLxkkw0jeERJK6nyisfQtITq7KIk
t/IxworvAuWFzsy3gTt70z23fTOABDdWlrGbonzz8QWY3BgldUBOT+TbIwBd111Xd7wUBhsB4Gmn
/THC/ZCZ+VqGrPkoBTRu5kXUxUrlkLyHSMj/uKLWk0Eqo+i9DzGD8ZsDanS/dfXqfdhoOPMP4YyC
nG62mR1izClB+bOI2dY9LY3LtHERRAOAj8fefOl5jLFuOTMEMy3fKRCFSGANZ+dJoazcXmm1gMNw
QY6Z0EBSqyjgFcBMaIuM41m1bsBShxNxpKptV7lt+bfQIklm7veClTAs7uRuEEuHgbv0DsfJfngQ
7Z2QsygnPsF/VYOMSiBC3Cwv+e57P5bcpQfsAs7kbuadVfjxFDwQ1ZD8PqxPxw8yOXrsgbYMoWlN
1PBaOPBxVsfAloApWyg8mJi608srleVYb7KHZekQBJMHWVWUmnotx/gTW0ZqgA0hOvB71aXA8HVl
Xzzp7jaYWKWNwNdUlrndra4KygdFjzVHQoOWgXgUtZU+gIP9CH838Z3RycauE+zmfujdgYbrxmHp
v0mkRjjd24eSDOmZDo/MhB5ltrwDNeT8dpb2EoWU1vHd14ohg8ohQKKNBSPeyOjHBFcABOG7nSRA
Z3vOwlVQteCkcOsyQW11+lFfeG6XXNY5nJss5g0TyaCtJzVKn7QkijwqDoohik7m8/HtT0j1T7cK
KZM7KwLv3RBQMbeH4SYPmVSqiDXEqpSbeuAfKHEvGP8sy4upDclM6JaDj2WRjI8NtKZS4OiVQnui
x65ORWKiyc6eCEW7C2GlGMa9ubQ0AnC9Z7Lm4GQ9oDSIHqiFk6pv2zOCVw+si8Hj/G4U/kHMGwh2
lgkqQJMb+iTVZnmjmg2Fte1xfNY+/LTIMI7osP6Uw5WA1u0KHuYVFuPmsO710Bh89Rxnu559DISt
xhXjcXoCgUgo4J5ITamBqZOhdCiuV4f+RB/oavGXGIZgDWRYwHfWCsDQ7LcK0ndp4lMYFoJnbfoX
FyXhEKVi3YJBDxmNlcxa5Pbo/PWwT9oJJNafrUV93bnn4XA3VaR4yQf2b+sX2rHz8AWXZoCz7f6z
nIt9o7+VFbZOC92xhzKfpwZYEhhRUOU0xk/m+nPdyQc4JC+doVCbGOs7CdSOFSYxxA2DLvTWT6hC
+jhXWjF53EbL6vzXhA3NjJSsjK2xIXn4sIjopnMk7AZC6TiClckU7TAe7EafC+evms695O+Odfo2
16WKNPRPvvq4wz9sFt5M0JJDjcz96VjkblISRT6yXTdo4IjgEi0EXzgtvFjQw4GTTmtE+VcDVkaQ
aIiyWicXhmZ8ULN73hg8pgZkyQdwV8OURW9gXW1mgfnNPfFh4sIYeCkN9uYfvDqxu9BxjwOKnfNi
bl6W5uAb0X/WM2T1OHyYVRmu/bzF83dP82qISmNy+Ish/WhOwHwskj97Shis5Bj/ThM3xgigl6uv
LxHxzvDztv7+crC2Il6dLu55eL/qPwjl1DbEK3x71k8x9E361EWejcOXWUBxUAIJ2tcYaYcgjIn4
/pa6WNCtdasOFrqXxaxWbG790Nmq3s07d4QODKn0vA/gzR0L2H3grKgqAzpmR6222IMjINGOn7EQ
kDNkHFExy/rCskfuUEzoIcml2RIis2BjwSPwCKisp4OJt5LdEy3BTNgkS4Lj8zYBVhazRhPuUvZU
lp6TYtFEJzEAJvrj7nKbQJZ8kKVwvfD0XYjMJ6iPvebiS/LoIV4leQ0L4yczMZRi7m++TFXH5JQg
eIUzzVSTiYe0hVVSiVz5pNxReUux2W3nN2fx01f1oSMx5M/5SBHgb2TyDR3W3054Qm/6T/hzYaEh
wXsIknl9xngfc/5baT9aSvHdOP95B7tchQaMCT/rZq64bRQVANI1lsOQu94iQqXSWczLFAuKHT6X
MP5t1+uh2uH5BJdf/VAJy6q7FarbJXEu7tXgatjxkfYU2BTBpslGBD9KEseJCucqxcoYr8ut87PW
8US+Zm7jk4z/QDg+eWcZPtrjvsGCqLV5KXm8wwjKi5KZvKILgHGOlfXMItB7bKvudiq2WXtUwocp
Fx1EuGxt1mxdffJ9TBrTCdx/8DKU2UqNaXH+YZ9FxoDMeyahgTdbUOfTOf/8AlwNcilKcqKVc/L5
gybP/9G0aQZrBlKTzgxdrM7Z9ckL/nDBxhPuDMcn8JHoUNBwnIzYP2YRpEvFkYyAK3TXXk/YN6Cl
HPDZ+DHvKB0xNOWG/XNVm2AQ05kGW5OXrtMXP1qEWbS2+ox9BqtiBYlVQFa8YcT1XWAZWqgRYsIO
qsXTfz8o3M29UCR0QEu/wAu+jm2f1/z1+qN5IPS2PsSrV9nA8FMP5DukkGxLQ1c5Ck3WXJN7OWnb
0ypHdY0228IWuj6vtYwaxbQMEKP2a5g8Xlmy8/KDZ1sXlYZp/JYYYBSysOynQRqPJLPDPF+dMgxZ
lFP1M6EC4+3/o9RztnjQYC+MbDPxTHYIkkDb69/vM+uH5yb7jK3cYbvbozlYN2lEUr3eqHq7SYCF
f4hjBgXiI8b+q06xmp63b3jAR6oWcVvId/oLrU4QBUAL0x27fMaaC4VySrRXPfPX4J59V4Qzgtbg
njmCCjV3pVPraK4CrJCJp3PuoLAMyK6puXyz3GEpCIwmA/jGTuRH16/ezxBUi9jdy1evoe1iwl/8
h+sk0SbYd6XNh+Y+t1TA7utGTaSKKEC8X3tb1xcnTvQpRJmPZe1Mh8idyJb/dah7IlO+pSSQZLO5
jFBNbBFyYhGXRJh8gSeRFppMAEo3pBCL0m8VRbJoTrqYFWxOHqMez7m67P5szONGljHMDinJg9PH
9L+zwsYgr3rEPmvkWOzrFm9qi/ktouTrTVBEmhgv48K3G8L2lmgymGQ3ctJkciEhDKruGeXmnC9A
e2A8U9oIga5m+xmf8QybKYinZRr4vJarUNZmibfexwNbF1201YGMyg8Ebpy5zQ==
`protect end_protected
