--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
UcSXWK2JsbyPB0SGr4NAUJLmUnsSyA4r8XezlADU/K+foHbQdzKOmG/dGk3TB1r52QKLV8jmeyf/
YF8hcW0tK4yF3y0HE/g4A43UgAUb5vz1LfP5OpCKTKJBFv/v52gLAKWDFfbvglx3rOXjrL5j7qUq
CSTpkv4YQ528VkFjmpObyIMA/u0Bgb081phf+k5pS0efT2a/WtD3Y6+k1XA6E2dJIEzmjAIdaz89
1oWHyjbOXjlfeYH6eaQWHVSiPbJJffL468VRslxiAfLG2rI5JpRiSgSWnue1f7/ihDEcTPb4cDHn
ijS5wQJieG5qv8NC/zuGGK2i+pVFUfWHMKEJCA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="TJPd7MLMEfm19ff5IpqMknsgwTlpn3wNUInSsywQXg0="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
EBhkB9AgEeVplX4toFNAAeZB1yiBgQLclYDkVX+8/FMEJz7AZR5ca2MjdiuzLITdtSQ4Vp7vKr1z
fXU0OLTFLXwxTQhcp+vavtsd/K1+vBJvlkzXxxgq1WTp9So0n3hKCQfclNL85RCVegh7seSs7m0V
Q2zD9o7EjBzhQV3yXGVRvvjmZv2/ezHjCvnqJ2eT9xqmNXminBHd+//b+DrslTj+/AQiL0B3emKx
LBWZJdVMlhHFAf9GEZA8S2m88pkRX6nqzR3dGyUms9iunFdZL9QQ5jvNA0IMGfwfnutLzp7czwg0
PWoIgNHWFbuLOIRRfMn1NJjHB3jSoK/NQ4hV/w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="MvEqGAZBStLbNq05tfx8cx2F8MckN1vJYZr7OjoeGb8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10448)
`protect data_block
vERwZcDY6uGsYzQjuH0qZ0PTrOAoMVOPghvQECq9Zu4nTw3EBZfvg8/ZYekms9dPY3a7AKe8DE/m
83pAfsXCEAzDlX/iNUSWSzcD7oJxXKQNkbzyyTKZ+Lhmh4o67eOcGnWBDfR38ePojdUemQhL4bUB
b9Hw+Cjcwoo9wiznFicc3fHVT7FFoVTarI9T8K6cvxjOFy0MSzAS+VpebhgAPTfRukrIm2Lf+Gni
De0PeI7vk5dYAd7kowz5x80ANVm7u2VS0hdb4iPCyvj6wS14e7D6JG/TfwrF1q5T7XgZ+T7TuwRh
3ZYQwaDR+CDcxGq16vAF+XnwT3hphJK8ePsp25LEBihePPlv7ahqs/TAfOfjjf70EM2921AMZiwa
cvhB5FVrdcczMVb1SmVxPBMzvfTTTwRuyf3kxCAehU4IwlZG0s8O89Kjot0H4lHLpihInltnvO8u
Lpib6/r3H+cx549v9k6bOnzsV6Lp5jkgXqOj1Pq21cp+uHjh+K5h7dZMmEnWtFE+2whMbh5hZLes
rq/+Q6L018bjUx2/BJYPuT8+QtbmIQQ5XOUTwNtcKqq2+UflG+cJ3LpMefXFS6ytfX1GbnFOuG5i
wVVvu21QnPYzepIMDnWMXefXitbC0vqm2b1LXpHtzNox11/VxfJ9JzNynGt3MJEeVCr3t2AfcXfl
CutGW974WmeYGOD9/H09k36GBaQn1QO+BIifTJngRB5NQbU3aJEq1hW+nLqU4vUOpSBCVm5yRyZZ
1YXEiIZkgoQZ88SyqTqR69WT65XQFJXk/vAf7GB5WtQxtJg95mlH03btbZQmMsaJr7B2Yrenbew6
vNGIITKCj15shXSNHDWZxGj9zjgxZCLfeOOkVkT1qh9o8XlIblvBx8lU8gdv1BmVmjUJYALLcW0G
W5KrOUkG18UJp4aQgpJEXZ4TJUXaLNFNOHvY4Ni3wZiPHBMqTYH8W0Rv2Lsq4AG34QxKiX7rqGSA
rRv+wzO10ggVIhOj1FyQIr05UbbSGOhdqgxq1d2PhcqfK2Xjm1DitQgxdV5I6P/wdhf5VLh0ST7O
Oqo41cJk+uTpW+43Y8jg3UFWhI7Yw0TwL/J6WDMj2Lgq6hE5LHvPR36crod2/tlFutYyELtB4/gN
CpjQGVfk43YM7je2k5t75JcOYOTTPTtgfxGloYb0cZvMHRE86nBlAwkzPARkMksU1BL8HQR9PNWw
jsfhLFW+bU72Ri06ub6LOEHvRqXm7sVC8JxoLDA8/zMj33TjC8p1y4LgFfUZ+G/a140tlUU26loR
q6jF1eoDGI4L7bPWfyffrGQ152aMXbJYn8cPp6QnrJ5z4KxTBOF6M+Kl4wJAkg5yxzZehFY0iQ9B
xTDlFUZkNJgVaHHzU2C+X7rHmHuHz8J1Rk3tm/B9GlpH1q19IfiVsZLis411JWqcWYmKWT+dgNhi
F31ZqGBcx0eFSGzfW2ZYmoseKhxdd8ZnJIon52DPwPfL71MDNPlQJFaGHKjDV4L6ezfXUTyN7WGH
2KTvW27zXd98SAPHF+CXe1Lry9Fur6fiZbnKmxKI9DpoedbQ6C2f9LenjJWBDxP9+3wREVPr0Tnf
B/9MfzBP4w0fU2qwEtcEXzYEV7tUhjemKcOb/K3T3qOqZPjFDBSQlU9m5cDdqKbCrGxOxvD38+Ml
d3KYUHFngTWrudh5+sSdR+EZw2mHugh1c6z3/PbZ7HYeNxMH7DPD03tZ/QNcLHXJss+PE3cqhEeN
/b5TZnLdkAVI21Tas4WAi1qvlyNc4l3yE4DEuuY0iOahK+/0Gj5Qm9Vf8ZLhQ84g7tc6YSEOjPxW
/yVjdwD6d4K7jlGSsaZHEJ8+o1lf6ekmPSLagxZRpJ/4T6aB+bRy+Cdpj2cAQkXsYtc8kHRn+Xjb
w+NCCezEUj6dZdcHIa9saKhcaexDJbqNY/EhGYCb7WwiLwazoN/y6NLp24iq+zrYzg5RPnF732D8
XsuxV/mfLDhs3BZJUr33zMwSEJPtf3F2KUOp3Ce7eUtLC/V8xnmmIDlZ2PmvqwaCqUtD2+MaAyRn
sy6cQKjc+EFVaxmb1DYKgFSt99YdPRsX2YCtDpn6hy/ugmewLUh9M3sD0zoKBRvFsyxKex4BNS21
zGrMJ1BP5wGO0nxPn7Wd6lC7abJnrS99n5ulqXwRW9gy821Xd6WCdzMt7i1a/pyGe1U/s5pfmzsW
RwOxJCMLOIcLkCHMwFElnn/VvAY1nO1Nsa5B6CQoPNmG+EGw7aACUp6vpabLPJAOFp7i2UfErlY6
fTVC5bpm6h4JVTQ25Nzs9Cis/TlRwLrMWp/rr+ivlFPcBZXDesnuorcg80YFt8zFcCYVwvtInO/z
dJxkH+ssLsWDhqXG4LGiPnVEI+XQ2bh/JRy8stsoDFhVWxWMIiTmCpTNz8cfiImtR8bnIptlqirN
XmXkfExhDwmckgDqI68EjRg8Q2+TFcfAUqNHjnUj/cVFW3O9SxYJ7BvxMDzWGlbikmXNbatN8r3K
u4yYI0rLP/kMutX5YZMc3cV9pBtozk7V/NWcUx4tTn6OBhkPffR5aY3f/m5WVK8H5GBQ9Ey/0IPS
TpsiKckkVDuEu2AmZbcviycFpAAJfXm/SSQEdVn3jtau30Pfump2Q0EXXH15ss4TWhGbzsDQD3py
6Lz1hMLEJr1uA03wOLWgG+VOms04XU1AuRMOVwpjQBjfLcy2XymcL5ikO7NFV0SLJTdA/heXt68w
x/93JbGPO47W/VD30Kf7nHCfPsoRoGP8p/yq9MmF82mj3eMzRlUdCQG1wwUifnOo5Vc5HYch15YP
7VJr++CwVR9QGlonP1EDhTidWqFTBPSTzYbxOzFL6KTi8zyEGGb9Zu534pj3xpvIKnzQIrqMS6L+
rXNrg9JClJwkCz5oF824kWByP4bW2AKKURAP0M+eXA2dFjpUOOrSBrmge5XVHohlkz014eORZxzY
qMlA4hU+KS/aFcMIBzAi7P+8eodCGzyalru3JRL7vpKhwpktXcyh56whz389U22Th/msiZPBmWkh
L2KF27bY+C2uujcUI5rNv34ymo3//9X5UIxSHlHvilKyDA0amMoxFyopsTuaxb0EOyWL/dDlBrRH
4UkImcj1VA9yd8X7uu8rXKuHN4hdNwH3CgYr7bfAN9oyp55ZlK5zJszlgWNPhPvPSRq4hkQyLR9c
PEW12hJCZHQO4q2g7KX1YQuMzJiT1a8BgI5Z1aYz3Iuu5arT+nbGVKFTCfOa6RwcZblpZtdL1zJ1
Hrya9PTBpes7P1BMPLi7jO3S9aGjNt6rVZWNHOn7Ya2x19ajWf9EysybZiB6+E1oMT2mbhfAUnmj
p0u95IUqTlcWckgT8Xei1PKvyBcIYiF+ZSXGEyAmQnHd3bMfWJLfWCXzMc7A1IFNKyBqu7jF1Ff2
k1Q5W5GgNEALftvQulTb6CdgdCG6rtkODU+MUXZFWUpLxAZWSYORBtWGNgSAAaFuy4qFArRVz13Y
Lzx5fi+HIj320YfXMwgrJxK8uDP0/OpnceRSGX1j2yv98fvALR0Q31/1G/U8EW4yibSwfqiP96jb
Ti33iXMTFTUd4DMC41vwoz1uzatcCGdNS4j6Wt8xSiag51V8tK0ydEoPvFXCKSzNn6QJQ0gctdxX
Y2F+BaLl/I36jJI4amo6/bFSDQrQA5FyBgVYPBEAlrFvvHr/mdYk6yNBugxrd80KieSJh4fIHazA
S6j7s92YAobBFqKQEL7KLM5picAx9x1Swq8T/0WohZdwBcxS6hXeNwaTTbdsgUgdgphvjvRAysFf
WH68NzYVAOJWhuObZs8B1h8CVbnISo1nEEGpM9sQm8rDYd5hePBiZrEUno9CCDOg0SYYQFvQrKvL
OoX1ZF0H0KAhzQ4QWba1zjggpTslHLFsliVGQhk8RLj/dmyOb0g0fvxoHdLKZ03zCU2DKdl6SO/X
g20lkGxm4ebc4XGmQ30a8KHf+8OsR6VyyntQKHttyWNGxlvdvdUY7vu8w4Pkmrh38ny7L55CuKy1
kuftmrZhTNPNJgvzR5kuKHzJHpGL9EJpIGuIudVwVaW4FFC3QAXdDbXY1rOHtairosLwawHGkbPq
727v7D2SmwtysuSm5rPvdBmVGhf/+wwZA6zycOHqFZq+0La+mWimGaiUA+iM7k2Qz9O5Ob8NFMnT
R4rO/8s4OqoCASnby+oxcsQ8veINHWWP5sd+DDyoXvHH0TivE5w9RRyd+3jCHCqZ0SQeMBU+9tpM
ZmcTUEj/sLBWV9m3zr34ltKeXRBPe1jk0+6E4+mPVs8SiLVs+1KVsgdEl5X8zpUCRKnDPXrfQhMo
vARmkzDQSP2xKjrhEur+lDfddT0kynzjuGO1q0hzgzvcVosogQRJXNZG9gJZggFYv3UejfYMf5jA
W9ukME3zq7sXaRHVlD1upuLxDL4tkyNqHOCKDZNP08UWRJ1831X4NZTfXFq78x/PDa7YyfRVYTPU
OlSvSbZT1C091e8Z2S9y4VHubEJWpwrkn/9mFOtftytPUfh+vy8AtMXkILtCeR8uZ3b9IvO9Jhss
xuyiXojs94K/Nf2GzN8iBfYAyprwymQsWgUIUgvyJsMSzClGcVNp368rghngpXCttZjNsdqi6+AZ
2fRhbps8pJ5ndkmwP4jpTAeJs2SiP/17qpDeCISLGNwD9LNKp0tSG6CPUUn+pGDd5Ais+18wcQXl
/aBHsaaBJQ+tr/nJPTh9r1OgrAK/ws2BqFmz2ftcaViccY6lyfVNW7DRViSGcbb9Vt8zFoEc+17D
eIdweeAHYQuJgiJc68AB14Hv3KzRy0Sgudi7/UeWK0+mNeB8+SOsTLvie6vG/92SUOnjLmAShFgs
X4e7R72QLuPU3BvlS63u87GGUqolsHM97jE74tDmQz5SDGEU+9aSYByBfUnk/xib+LSOrnkQiOJW
18XGwCT82L0y0RnwiiPe3KEAhClnOlQ6WhMgRzb9tqZzP2jbYxDzblGm52F2x+YoN68w3ZqQSkMl
oDQIIUUgCohGov0USmGm3g+o9cPkYeu379wOErdhR0mGkevF/XGA4FD09paHKJ5eIPto2pHektmZ
9TPZmQhaYxtf7dcdzsA4xoAnIaEH30jXvl8nLNPLi4sK18vRvTmgekGaQGtE4H1qFcQMfsKL82Nu
KLiZfVmFCXTrQwalUH2lSnBQBc49a+7pD6q/ibiT9fqwLJLwD1g7ccKYiHcVM2zprQ/WseFxaAXD
QQO5bWfYa6Nf3GczW4t4fUyBsHlMSBzKVCdWGm+dGuxxpNasYMpBZs5KvZbuZv7riOty4Ij3g2WV
zKgdia9XK5kZqvwoo4tahJJpPSpnLOk7RLAHeytuSn64Fsq5nj1m+o6fjRX/TW+G+I6/WlpRrW2R
dYXZidvxpWElqdqgCgwKI/3/VOZTzOPAik7TO4Hf40kYQCsvAYl04t9Ei+ZEYPpsbR6SFxZTJ16x
bu2NA2h2aXwGEEW0tcqHrTIfgP9ssCBtpSgnrqGyEitjDU5uZdg6ripK3kkFI9nevWJenvpO1u9B
Ci4KyWDiDtQz31dV1v0PjZS4ckaNOihXrPFGzGyibisbo9+w2ycLPzZzXzJeQ7fe2mp6nS6x3SzI
DUmoHp5pfBNsjDjFdiYsDKRdnoMP6Za905LKl5vtZDIjSM1i9QoCpsWl5xRtvOtOzPh5oPqnUcBn
zwsvJYd1H2eZbB2arzBgLm4zA8iaEscVfpR3ActiEV1uOdCc8vP9u9bc/Sztjdx9sBVxN4Mot7BL
h4K/dfCWVtNNGd0InLToqsgOOsJQj+HUVSUdtolfi9QQXuye9g5tupIlXAecu1MkGqjTVRta/M7E
Vaor7TVdN68hGJrvrmrXtZ3ibEBnjucwdgKsVIHy0aLjlm4DOLM18GPcxhqCjqOmPf2QTu8IJhZ9
VBZv7znXi/YMHX20A3gH1qSQYiYeEdqHjq28ku1NkcBmFxM1Y3DPSlPkS+f1as3KdJhCzQ0TtENI
TjAEn0d41aiKHjBlzBh8U2h58JZ2B1mH6kI7PY1JluYIFXtdtsKJWNlcvHRWivypOoU0XoZZi8Ql
hKK7JxXeqrcfDEh4HDapi6KGQykDthMDQnBPqpajT9+T08vBVYuS5PPUKdBM4sYaXMWD92tIHLXJ
BDuONvMErjWuoL1zudp4dfKs5JUl5eEUmwdAcmWBsZuu3cG0L2apvFLRvtjCNzn9h2Ufez8PUVyS
eV4/RZ2g1DYPfTiShXPL5O6XUQsLV2x9wb0g1/EXu8+zczZ1G7hOgy1VV/vea7yF3e294DdiAG/x
eHMNx3RHvuPm0D94/6eBKJH5LZdFVdJm1iY9lRsEfypgliOj1dg8kIGthQKOk3k4gjmqakGVjtN3
19b24DHFwGfAwJioI3qHagAJZ3xgXHPiXqj3M3rMHQLNZ+xAZD2wSNlwbMt1hKzLTI6BBq4rTrHn
RO1vNf5PgqTWdWcWTt8z15KekQIN2Ljm9MIXHGCbTc7rkas3xTW2lOid5n6YzEZpUOrRPvlCZn5p
uWkKkqFd/Lz7Ehlc62aNGISODqln8+JmbzDnERYvWUc/M5mrYJz4L682RRMOsN9FSXIah2dakWfn
Gs3fHEyoFn9+xLCovq3zzE7OnOo7lwnZFr828EdtRP6UObxWFHBBcQjK4xtbSLJFtoHTKlq+UlaL
EXpjfzUwln4whgFtZrhB59HNWcCoXpXhlLjUpKMjgWlP8xf2ObSeIg6JhepyTUQQZc/GlOIrWaNP
TyyOX+oJpK7IktB+2syhOKrffDLASlr0+fqVNIjWz1bllPhPV1ias3BfYssNNmIx9PUyNpQNTHVv
i/7M0lMe+IncLgsEhSU2+ou2ISY/H5oUhRdQ7KEu/amcQKK70uXbt+mXBmMCio6fSSnhyGA31L5G
ovB2HH2YvevSOkXRdzlRRk+j7uaSq6t1q4ADvgazLlNsizhcpeKICM/mV/Rr2AjIOY2pp2oaaPAP
3n5SDqRHHb4MgeMivV3nr5FkGYutgtb4vxs6o5h6Y2yOIrIW2a9mi8LcKz661F4cF1eMCYjMRn2c
ocQJOFs2xtDbct7W/9AKsBeMNhCGCYLQfvnjIBhkk5ws6DzDz27ZAZGYheeSVaIa7RqKnIBllqUU
BpCE0fc83ZEdli1AaiVxte7RdrPRnGm2FJvtfVmvIcBpwYIZCs2jvSH4OuP8wuMx48PHbA/escem
zsSVriqOY5pwLE2ijtT+OcpRPpx5OPCC26R4ebuecMbQboq8VJ4vv6pC1E5W1iT/Q0K0Pj0DRBqa
VhOgazTJVHtHlxaK9tfsiiFEcGZOqqefhs2Z4RmnkbMaiLrHHXmYvbeQOkjDkTr4xZvH/mU9iTbr
NqVTQPb+eA4wyfvJATh8Wh5OBtcYH4XGaSyBAschDCMTYHQvJWY8CvxV7nseiv5LDR1BFK5i7e5k
7JE38k+QU8RZzGkcXsGN1y/PzR7PvW9Mz4QPCddD024xcJJ9nMpQ2pOeYt7Dgds48cbBNz4pxqgn
qYnGon7/RrSGWOuEp2l5RHOXAGbG5wgM3NOLqllM4vgJ3fHmxiMNuxRDrlrNpw+iDbj3NeI1pj14
q9GgN5VJkNQhY4aNzliMns6se7GUyYoIFJqOS4um5je21whOSqPOOyYpv9F4mwho1qrkHnJ+I9bl
G0OnbZRCzOX/sOyNaxBIp70+SicwLaa3EtT2CWmUGME6G9LXO78DlKtagfYpPxoRSura+t4I6qGa
PWcgZt06TUQgEnTBVyOtsBL4o3X/jDe3JJZUwQgJkTRJNLe37oSeF9kSSdiAFjHD29lwlqmmMsOJ
rBmduvpCjLN1gC8uuLXVHFU9xXZ7SxmJRfpul3r2MIYkrECzzslLKHlbQsvM53GnEELeyfPg6Q4U
HxmJp4eSMyVomsUEnd6U1/didiAKEshiJKzUEVxH4r18SeFJDyf+3sh4X4KrMrmCZc6pwEJN6PWa
DSu7vjepoSWGp9b03CHaxwwm/8m3J388a4ZN9Eu7Rq7hlSRei7cIX3ohbC6TWw8bXgtLKbNCD84U
/Ffc7cbLEDlH+VuTurdPlsAG9vGqYgafp/GswWRNaEu3LkpICOzLNnDpanIX8rr/wplzTSsHXLFa
Lbdzkl6QzjwZ46x41eeM6F7wGo74MmQy2q+m4HB/I3+P1XRihS8KUtr68Zea7duXV4lgHG7vheCX
gneAtzPQw0ZNj5BZRCfa3AihHHS8rIqeHBcG8SE7rb5+ko/WErKh6MbtDbExixk6DsKVRN1xgKSH
IQwiPgY9HPtN1yY8NmbToZKknV/zrZBV7gPHbexsR1+7lc1h2gwleQo8FuTBvbwxTFeAIVY0XPCv
YK1u2uJ3pm0NI8x/8/vW/9xdimKNGexhqH79qfKLTP7scBP88H6WuzkycJ0iU8AAaC2J+bHpbBTO
RBh2CJzx1mGHiAnT/gH5OuujG+dLy8QWzezN+gClfXNg3OY822sMvhwrs0tRk5HgRw9cUQAbK3HG
BWvRYYGNwTC5cCiT7HxVYXL7KWPYOJPdet8NyM2l5clQX9l+vUcp+poeqtBacOFAL7Ws9Y98vNlR
Xf7uO0TJW9T2OmysJ4ZpV8W7MI8td3ff2ETTJfEELKpJ8hUmkKm1VtiDuQ6hV8vKyHaDHLr65hBa
/y1awIZjR4tFo2KO6hOAGL7cnX/fqVTu97jmXkmdTPL6Cw2CpFe6FWsreSGGx85D5xunSKyAMIrX
Iu/iwQCzyTWF49D0cgM2tXAFjk7zxheh0DShjEaXj1CdrwC+RoPEerQUY1Q+eRzR+3gVgHQ2b5rj
Hq2f/4J2cbQbaXFWdqTgAjmb3vU+EfBKLAk6HulXLoYAdO32v2iHjj069Y3JwS5nCgpvZJouE2vN
cqaftZS4ZO6hsGR+hurAsrkdrWPgBYnrFNM23vyVSO5fAuILnBrO+A5b/PLc3/XEVJNmBssCX8IC
yZEV1dyLnBYkLd1zdJHlOAKi1GhYwY3+AA3tcVWaAxm+JgxKAd45ILWIXERhVOxojgGxNWJWZ60B
q30V5oOt7OlwbgkfCLOzBuZ9hiGt/tcE2S6NIE5TKQkShcwWLnZ/OP9Ooujx0jZt+p2mwbZtFKU1
p68jwa6oPPZAB2EBx/fwgne+OKyTT10Ai6JZAX74v+e91DsfL0c+7A/M9VpbLGY9uDKNqMdf2X4/
zOv9i2IRH5j11r0mxhL3unh6yM1FJNL3O/OEhMkZeCr5X09/2Yf9hoOwtDwU4RFRbCe8ZjVWvNoK
xR4t5BQ8pVFQ+Ooy1mue+FRu91+eaa8oF7z+TYby7W3eKDDX6Phwu7kYQFiOek0xRFc0fTNhaqhy
Kxn+/MYvxq+UIFmF6i9Dfapo1RKjcggAMIAG80kyQWFPt7ko1WMuiDq1Vv2mhlpzAn3OruRIhEYy
zpeMBE/NEIv5h0sg2seePZZwHVgxRIcRU2URNovSWi00ePtvcEHC7Pwb7sDiCERxpX+PCjFwEogG
2Y/5rpmDlNQsd07s2pCizM01SPIsB3HDBeUXdSGDrdY81RJs6UL4Lk7tUavToSJ+Qynyh6yf7P5g
J09OueixoQ9zc2jxRX0Px0QFbyYpMuB7H2t/t6/CGeh7rin/I/8rC7N0GQoWKR92+XGY5ZkthzfN
kolfA49QBTX93MlAgOSZYV+4+AvZHfKxgeOBHoZjJT5JpBhDuh3Ph4YKPN8bKOZ6mJ+sadB+9h1j
/bbTzy6IbF9uMx6SoJh80MeuZXqAgAqpsbAIej8zUOWy7cvbxOZdhFfc5aO63KiWHdWCrjM+b2T9
LJ23o64Ms6YrYUosNo3DKbn/gJCezhQKf3ZBi0EB/5DqvAy5f9SMH55jx/Raq1H8qUgGDn7FaHIf
DQIKG/GmbVWjXBniXIyFOPq0M52+vWc136w71GYeA+/AletU3YSE2V9xJEsBXPp4qafLq21/KFDU
BMTzXH4TvAptUMaGpCSmUjgQQnwIa4wEuQC4J3EKgLqgll2g4//85Rgf7Aav8rppZL6YDQTKg3NZ
nA7utgUKgD+6U39VZma3aVbuO/CeOWujNuVbGL7K2quP+mwvy2ax67tftKDZTyI7ZA6sKf0BIPUM
xnVMJwcL1Arj53Lr8fpNp/A12jPnCF5ZJPHvgItWN6/hUI/ibwq1L8/Oz/ZRbQcZb/Gbq3Do1X9o
iW3To3AElWqAHUfDGhqeazHVw0tEauOnOG0tA8o7CnvLsz5CiRWtC5Rz0Y+zX7nUM4T3ii6cagvd
znAj3BFYi67BRt0+aVjSkM1i5W7D3Lb9Ysum0gxEaDVeXSd8/p7k8O9DFiT3Er88S7k9Dxqp+fPh
aIUuGKUFLvn3Pm3o9IeSZJwtb4cYp12iyvJ37PgYRdI2J4qRsB/HxrcXWKpR4d+O//vw5a0auz6h
fDAqHugrYk8YRqwAg72ceCTuKSRnQOtT3unEu5KD7lGwziJ1RfRr+NkZBNfQTvT3leKTSpzphGGs
I0aGeaj5RR7dNSZWsghwD8dpDoHicePTuBuZ7cxo5ZWBcnfaAfoNoH8BM/yImqhe8VKcOFW0KCw1
tQOJJIHYi9W+UlAYbiLVh8zdmW5dTeHtdVZ4gl4svroYCApb1r8VQIegdQu8jxu6qg125Vlj2IzW
lj3EgUN6yeV1N2hM9+Bllh8N9V1ZQqJ1ZFamZefe9zRvu+5AjMP2tNAhy93Qpqv+cK3ljB7xh87X
WXtdw6e63DtVnkm21nIhNOquYuYiSSgLRG2aZvJ6MjP7sbHOqP6LXliKsnHvFE3eXcPTy2T8iAhy
+KJH+vLaiZKimJQ/50sTidSAHMjGOM0mf4TkxSwheU5UVE2WJZe2HlBUvtn+QQMXfrnCfl8+ZZ7p
PWIqRz7RU+g6zs2y+fKZLjEM6WL/00B68VBlY4Ze1NpEAQoNuUWLFB8rW3M456QV3uEX1E6L3hxm
GKPOBKXDEkMG4M2fBbJnloM9ZeRG+2yKNkPzwefFF1Xm60Y8wElX6eCtKBXXQP0ajHCitWiFy639
8MXQ9YLowI1JMugusBffOJJ/eDuejSzqxyjjbo8eZhoMjYba5qv6V2FQT2nIdmrGgGmAGZtAhk3R
JUqcWw7SHOpyg4itKxo+bhUJNgaHQlDSywIeCnvd3kmNTJdPhV54lGZ+eW+JIl6a63g9tobG2vy1
MypgQdgTTp9m3MLHt7QrkYZEVK+jeLUdspxSi4xfxkeJzHNdG9Z+ehZu6rZBSyFCO82Hkj4D/FFW
y8fcTK4HnYz57oP+s9ovdIeuWUiUGoQR1kEPwC8FLiLp+GCTEpHXtaYd30sqlxA7j6bb30LE9sD5
PB938EGaayBJLUCUEAj7KdnHU2e7e9UwlZy8TZaT9eAHyVrFISiSGSQ1spI9/GmNQQprWojYVgv8
fl7giux/MQPP5UNkzlbnm0D7OVXctj1S/oDlOsko+Q/B8RaPfDfUmn8dUyZq2GJRd9iRauTVuBVq
VMTbaB+2yM+zD0zJM6nsho7nmHppukifP0VOExN5jPDmYuMF+lhDqrkGnJRPLSRBt9mF6np/yIKl
44yIbMMNpucwcEQj7k11Hbc9lCDTjZnSG2uHhB9DRl+E7ognrSTi2UsNCYlNJn9JYKk7Y+JXyKcy
ui/16V7roT7bMl21smwwpckvNmUWszL0Ow48LogS9ec/C9XX904mIgoE8KCQjLRPpAqN7QqtNu6r
JUDZQRYJR1JUzg2Xc53c7Sak525g7La1HII/TbdXiQdroEwGR0Dq9q2TcYi7AXuxy4utI/b9hKHG
Csbjo6omt5j9xCK0U8hKtM9duJEbSpeH10qX86zbag0FZGkcH522YLv43MIUTqXrJXsHa8w18Crx
YrdZWJnt1FxssHLtJ1btl1dwEmfR7+HLNJDSqQHQ7SdfY80QouFwoYy6YhkhFEO+niYrVdCoAtXn
ERjb/T6nTar09r8MV3YUvqOBr1CROCi2s++phnPSpql83KHqlf6to1tjqv3OJE7qJNPAht6A5K9O
SDm0geoeI6LTulkp6VI1yVElLcRzvyvgwJoXLnsM15A7VkrYvE+6Nw6BC5vl5NwNlbPbCchuc6Ap
ebInMQdA8Om757XV4qA8AQHC8NTeM9PAKfZnSSUj1LyPmlFIr8ujE8wOzXh3vt3iy7+UH/pi+N5I
vr3rdFL7I7K1WPolxNAp6OIa8LlVZ4cI6MNwOmjwfnHJtBxdxhDbokfO+LkGOezd1jITW914MW8x
ozYa69CJ0bHbsEMqTJuLxWO5YLAmmfu9JoTCQADJse5lWacxUrBcwCuD7p3CiFuAy5H95QVxa42f
vQDWo8NBJ6a6KcvDlo9CG6IG8rmQ7X9rrCAgTxtX7XFk/2hJb5lJ5UnMH3oOa2yvvoVB3ilKk6Ny
0AhmE6MvAjhhqaHxhHBfKFRzvxjQh1dZU6JuV1o35btbX877d1FbIvlh5N50yeR+CW4JrrtgATyV
s/yLD+hDxd4H4RVAEyRVMg15xMiZ+Rh2c5sdlJYKlPA1pGcr/gjdMzaoePMlYDVtWziM8R0wpWf/
5yA0uOaepSfwDVEVAnhL35V5otBBBTVSq8mtShTs1kUvrX3vJzFmlO8O9VCbmDLBD7R01eOg5pwz
hRIXK2z/0RmZqgWyd3HX3WTrsvFZlw5s7k843GU6hIpRTUhfeOYGnU7It0IvOrx6TMA9/3PQRWOX
02S8ZsKmlxfnwG3QPJ3lK8cYEIdFZMVCOAK6iphu9pztxt+9a9pmz0DLqwtN5VN/glJBpj0oNRbq
HPGaEOO/nmrSSWME5tMWRGVfyn6jwOkwzCRru8ceOtMlEswMSSTYHYeuzAuMuWD6SCTmsyi+Hbc4
zhy2Li1C2DZNPtX0d11MBNfZqMlNKPmlrJz8nEpXT/QsOWvxtdyO5rudN+eFO94UYUNhe2uPCuy/
8EQdSnhVevxV+NbIeQwFTdMsHtkctVPwL3yTCeKX79ii8TjLy/TPiq77tmkgbQtAqq8H7rev8xU9
CgzDupDvdwkBlu39pLvb/vpLwYgyGRxSXwn10lOF6deBx3rQoeoacfA996NseoErmRCF+xIEMHPw
LzcvKBIgdswPsulp2VtFCtPAKN8Rkn0KBsVdCE3eXk5e4cgkbCy+pLbkujrz1rmYiVkoMqKns+aN
HFxz3jdePHScXprmRdX2G0pf+C9eU14kWBcFnbh8+uvwmwhsZ+o82q7gJYWY+oDnJc4CYzmvmWg1
hXUFva63DwS1xr3TJ338wb7ZuHtHLj4GF6rjmGpmleqKYTgGMCQnoH0C4Ib3YzRzzJMJ8eYdO1F1
oy5D2kHijMoPq565VszQBHblTXEcO9eMRRZNmWvB3AulFvYh0uaE24sMpBTXt+mk8sWICVXPixdo
v9IxQfmj4hudcLkjGobgbFQ8AQP+r9jqoHmGHvXChFVqZW0LtujJ3cZatQE6dnec7JAduE9ksi7S
okjuUmQfBbbika4wUF7PfcJJbaoFgQTpWVXG/pthx8ilFARQMM7Nj2dBx4Jr+iGQfFIUIzGlfOnU
FlevsJUgFRV5Fqwd9DuOxGqOhRAnAQEZ3Cju3+lmHnxrSJsKG3Vi95M+vUm4wiNb6oIXIv6OWXvG
GLQ3shmhEzywkg8maSZLEy1wUcJW0fEz6wF8nH76ZvWEIQbpLfO1nRY/6aaRF3DFxfwaERmIhZqN
IAzqJvX+GTT+SW8ipgJeBkTR45BStJOqmJYs7Xt4H2hVRfaAjngqNZd+lSfchjgxQduDaPAFco6g
Hccg9159CTWMMb1+vlv22W/OIrxfla7wXJvpCsN/fQrhBQNoYCunwId3lNMwBelWwo1hxH5/Im+0
rklGKRx/4puWKj8XZlqvhmsGd3QvZPNclpz4KKIfr0N4uj5/zTSge5saowhJ0i2wxLhfJEyyb4My
/BTJ64EFY61blcQsJ+fHyXg=
`protect end_protected
