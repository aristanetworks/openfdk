--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Pa0UGWHrC+++UOakMtqZIvHvczyYHqErbUD1e1D4OGRrDazY8Ret1u3T0W3XoH5CnGxJB3lLC+xx
BneodjoeU0OdY4QIurswjRbdHt4mf0sHDhiCuXeid+Rjn9acDfEsRV/x0jWsz5uxsXUKIhXC3/To
t8P9+XxfSyW7TaY1JTwLAxr3XTXjm/mRa2HHluJ3ysBFT1KEtCn0ugoktV3nISfYaTxvfM4W8cRb
AOllJmuf3KPU6iX7XyIgV1egQaMJR8oGrQ+fc6RX0ycT6eCR5eC9UB97NaCkdAZVmPg19G47oLRE
63ON8IJ80qQ82HfIiC0R6il2aYHvGZsKCzT1Rg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="K7Dtt90FnrLylkVAwNRwQNI+6W1x3WXIjGNCCQ3P4m8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
SKdMJXE4SioAN5dEyLj986P3kwVE8fwQ2j9Lz3zwdOck3Ew9Y3VDuaZ5zFOSQoaazngh1b+4vpKD
exbgjBz2e/TCvPamNija3UHK9fXDGr3l2Vfke7F2BmE688LbbLj3KLR3TUQV5s3gwD8eBcXBSB6l
54euf4uLs9ndcH04n0kQ3ZNXihtHfLoKhDWfAd/XKxYMjxq7NjPaAr/OGca0lcH5jUKfr/i4b7V6
8X5aIo+NyC6vbepGlkYjRsRlURQo/me1OY4nClEm+CMjQggBCan7irQaFyLk78/EPepSNQk0pLdR
EjvM56TlZYrL6GJvFxhfI7P/SsVKZkwhEDRNRw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="TWxfvWNTj3vc3u9o42iK6ZQqp9WL3v7tHVaBFM7U/ao="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17552)
`protect data_block
PJdbFxW3xiWFH9ixN+TfdAMwxrWqBAk0yZM3KxpCkex9XZzbXTj48YutyeeP/7n6BvX/EY57iEWx
wtHxIaBGHThAnSTYC4nNikElU2PvN4KxKgYXtDo0kPDnloT2SxhjKGiz3xf73L4fZbdUnr1zCoS4
1SI819SqmR+6A6atTRWljjOIfRtMEzCLGIJtc3twX4z9bd2by5doBKIHSqnh75gubheopDEWK1JW
qdsQbfFOjXi0MRAqaCOQpJ7LWmd8uOUubi2pQ0uwqVlJpRgLiZKsFq2jvL5dEs06Lqv9hJN1mwEb
CUwB1dUtYcaaEewUD+gxAkoubZkJdY4rJFy2+572LFod5Hlon0lUg9XgHNdyNx6rozndwueoMVY1
IJkAHeNljZfa+xrLtWu5vc555QwU4hO8+OIYNs96vLFg2H9WRqmlWvm9uuz8whbFE+rJPi9Nnhbx
sNMDfXPSyXbuTnTe+JIjScmb+xeZPOZAo4sEsHH3e0wut5jmJ9ZNWORvTCCn+0mO+Af+k1ax8AjV
Mx67pfZuOg2VuOiRZDa/i03SoR8zu+QveETDt+3kldskT+nKg/US4udJZfhYTkRJ5MxU2His4sz3
+WORDpN0tsb9pBsbegN/F7MURk/6t/V0ldyL3JG0JBdxie5tIkZ/VT1A8yHmUTS8ch1oAPZZ0eEB
PFnOdrMG0P2pLZgouFBytgs2IJzy82Y8QlEkta1BjCG3ivUhrg9g7EG543GRrdz2ocXD9Gi8hBqz
DMkurnsA6f4s/3zSOxJnXqeq6xhdd9NZ0ugW3hLBQmnoW2170c00uyTa2KCWA/kTk6HobG96nXBt
ZOnoWo1K1YADVZstN7OzigfpHTIJlHTM+FJuVBbo0LsYoryITy3cNpz5Fs+NvceXFwvh7z7cOEbj
/yO8phiaYbW6IPNJdsXrCpBVXWyfvNB4HCtB76cplasoc7+DSOH6c8iG/D0uzYyX56Oc75f4cEAn
bWFEB35wycP0oRPw01PsNNC4HRzd//1owRjyBqBQoNIOD2ClVDuIsIQ/g2p6W3TG1H+UegkjgKi4
3r8VH/7RjSv2HT1aYOhtxphi0yLV0jxI02z35kLxTMwjn+7nBX8XS/50HfjeWiUiqPt5kpbAlA0/
VflOcImyFx2D3nkFSVukHhpMl17CbdF8I7DlS0/ZUCo8tCLRICapZEkbQInXYxMxrjCAd3AQ++G1
2leXc0nuc69ErwdbsDEacSTw0VMPCI5kYB+KPzwPKfD9mrE0UmxcGH6jjZu94P857XznKUZNJP0D
0hlknRY+2qfNds0f6ooH0/Ciwq5b6GfHpjLLFGNXr9Mux7MU9/jsHXZy8RFdZSeOY2ZXyXN5A1TJ
M2tMI5ZRQAGPBO1JURCJKLrCt0arvIkeioi8SJ75KHjYSUYjjGhTLHkQ0ko95rxZjNtI/IzSeRNW
xRGAovlQBbSh8dzq/HeKxnq+sCg4x4IySK53a9PDoVTOsT83Zvaw/UEQyZmwDRDnrtKZl9GPMBJQ
2UfZ7AGimwsiQzkzx6zWGl4xob1R9/aqJnsLVIZz0hviNlOn5ZRCvFUFdtIiGf9uNYpOGgYQuPUm
fAOugIbBTThgkkaW5sFpF2AlbSGJYvzj5LFB55EChOBL9fEw/IuHP7pTOLkByGEBFZHd63AmRiSl
wayowd2+VcjhCf61L3IGkHLX2OYpT5baqcXmUlyBwShBbmnoY078jx+a4RDADGe7F+2A2bA53DWF
mJv0YnMibkxs44xOhMgjepF1DeTH6b6Cmchf9TYbTLghPVeB5H1UNyyNTtdLgGqRT5kKSzX3/auV
TRTpX8X68NKuA3Dd+7p8lSuDBLIbsWGqFaonZJIfgW9GmGOrUGFyP74qAT69AwkC4KnHUUCN9maf
WxZDCnAv81XJk/x/UKVUe0K83+i0FdE/jJKti+i44XaEjmi3ICPwtkH9PY6cghNnfI81d824Rvks
yHtGkXwtF17MdHu2INNZxHJkAt8oODfyLoIv9dCHgFtboyr02yfYSHvJu/etbYTWM0f6umqkWG2X
5gNhr4JiN8zR2Vyh4lTgRuI5Mwbog+qGDblb3mw4yM5G4J7eemxG/aaGc2OthgvOpKn4TenKhftm
CKiXL2iAA7rE66qsjbyrHF4mzFWFea0C4c7AiIBqdTE4FYonHM8RVcBaOCxyUyAwI95kdR+i3Vf+
LvWTjJ2SpQQLoLURpkPrYSFdY+scuBUjGaFd9/sXj5Ue6agGH1IbmXBNGakAZVh3YmLVvGshQ6A/
qRli50+bKy6qB0Si+vVu2RQxVRr1l/QmG2TOuth2I2oH2JwKoTidfB1UfR/PvlqeV8bVFuOYCDPV
jgEgVkELkBPhAhMqsH+DQ+hAbkGw1/nUhb6TwnSHD28V6CRxy6GHZeEIj4/L4n+aJCkVgI4Ighm4
xANWo29faWkPSes6R8fRCNZR3XjTQMi9fHyJsFlgPLzGZFV/28dmCY5X7TbvO1k5v3qieew11J2e
hBPEX89JkYgR08cJ+x4xuIg5+Sa+WG6teduoJFRLNWtpHg/foR5OhL2Yny3GTs0Xrh0dwK5Fwawa
jpbYMJ9RTP+qtXQJv3csGmiU77q5ptPgDNRqHc+1ChbepkQsF0yDe58CloSx9syGA6mABmdMFogA
34IBP1W365GJkveo/NznrxpcoNhPXEade1/9CXNHhnWAzlVtTLOid782ZN0a5CIoGXDQju9uEs3Z
drLVud9WnwkgX7ssXf63/cAC6TbowMfnBqZ3Js63yRDlB829Aoq3+xks27ohQDzO3TJyzIpfqCpe
pDmPqMDZb5BY3gjeVOJ9eZHephVYPEwlYtIsWxEkkiuEjg7v6stNAKdpfvhgV6er2enzhLhgacjK
XI7nlWXdzFBTKekygHhkZdprL33WcW0JxZvGq5jJaFh2ooVeBZr+usizyT4GrlZH1UHBCv3GgROd
pnSl2xaxXn7xPn8fa09g12R7TMEPOLdWBWi93s6ExIcm1McncPLBXudhykVpE81fXGPSYX0gX1Uy
espW4l2iVc44qZX5UOGIG3nCqV5Z3zx7oexPIhXnwaTkIumRB/vtBvfBfVsbLzCBKYH04ESyjBii
+6EQQlE7d3A0MxJbPiGkhVSehteR60mokg5OAv+LxZ0N8oG0kwj3hZavYoKZwVimAIWmXn71EE2/
xT83EVoKa045U3A9u9nMTlk+SIVsKk43kGmGggJBkcj5NnQdyZRzTMIEzcu/9U30XHv+rd7BsIWj
3UfbHe49/R42cDIfVlUxFUaYWhNhBN+snsjc2tPVEQpnJKVSOi/OoXxq+Tl50U6Uzvg90XIeFlH6
eyCyU2fuNKS9IcSGGz0g7BsNoRNnzv8qLup4+UM+y54kRUNeoQB3b8iuSX6opkJJJqNWiKmf9Dmh
/lyRleNi01gaV7bcTaFWN/RQyW3iL3B/cANtMKqHKkaBUUbcodKNz4sEI+uue2MnG6TQYh/RFWO4
cNYA3pTx2dPv1T0CoHjmm9cMW/TSowTAuJMsyryYonL5DLsYuhMMW4ELyvSY+j06WROhe3MRr925
g04/PqO6+SXluviZS5d9bF6d76dliyOq9NhO5TBpYj+QuWVn9gdBwTgqj0TEru/MJtburvSn8ywX
KDAVkM5RhPFNCWzocOnmVs9g5NEy95Hy3KtXZbuU8spi8VoXRSJhcs0IKZ9U+AC+Iy1fwvRl7s6G
MDXiToV/OXiRwkQsPWWJjV5qZL4os7Ef5PZs8xm3WDta3c7fE/8sWxVcKrFBymTAnGviijJhyHln
sgSS/kXC0+5WBcZChERKpePV9eILfogxOLAL9S424XdcOGa7Hs1mBtvO6n7BX6KBo12v/BxCUCUu
IEWsna5zMGDDri2Z0Qtv6y8GbK/VC+md+L9Z1J5A1HUi8jZOq2BuX7XC0tEMtNkvIw1rMH8BNt6z
SLecZeAri/IU31NvpWISLsLzpRMPSQ1hvIJAGOVFpa5pgk+asPyrb1kwqsKFiZVJEFrIWREmuDWu
V1L/KxQZlJyNs9xe5Y9VsoZ8EqEi3TnjZJ4T9TKy6Qn1fxyBhnGXN8RO1ypkCs2+7sfD21AQNh9t
AN0ovpvU64Go2OcmY0koxRIkkHxf+D/LsBJaiZ6P7Q4GyzxyzV1wUWF2JfKWlDO99G1fmvdjpN2a
nTlOzbR5Kujm/z94aJmubz3SGRpUybw0VA7xHZRNhukI/sHRkGa26+YA5/w89rbeNC52xpKE4bTL
Z+7AHdMV7gXGioSwOfnmdURQVEzsUjrybTqVtMk5fch/6uidpJcLTHKENN1GOF1MbKdg++4YqBYX
QLcFXpFC12aTyTMWrdPiRa43gb9YKipNivPgztJ6yJgWh2FeiBaNK0ZyX2IOo2iWZWLdm9LULajj
8LrlteSPBrYcDMRPDULBsBlECL/I0KJDVX5bM3igT4wRnv+jUyFcbu2vf08vdIuYSr90l3W+MvVo
UT8qrPti6wGRZ/59Xb2L/HqAw/68COZWUzp3cQ/LShoeWRzEjHgyA6XGbWaIEWKf+1xQx7DqoBnZ
eDaH9gODPe31OeFY+TTg4N8YzzRqDE4m3W4tEewkYk+hPntphoEFqrG8i0wlryQI+fN4BgB4qX9M
k0bssVEHoAU26eeTAR/gFeDRqtPq0pw2CCRhhaq8LW1/+oBb6ppDSvcKK1XknoNtgCcZUEvOgffO
xDYmsPoHYxSc/fitb6+4tcjl2MnjfpPaTiMtvYNyWNJk5bx/W1VSO0R7x11lyCeMo+teJRkRHmsb
aaOZ9mOtZ1gbEfgXln8UOIDvR8O1a9/iNm5tMKAUN3/JHodaJlS6wDieTV1MdMZgBCKtDXYY1JlH
GvhpYQfJhyEytP8L6yOHIb389zMrkrr1z/p2/5+E/aTN9V8k5DUqCnrQO8WuU+ZxHmEUebKAs5qY
CJxErX1VPMCS3g6IDko9UurGhsL7E4BO5On4YM5xEe3urJibMcVriIoGNaBeV50ayusWdgz02P4I
XOcxbPpN8/+qyDIGY/xf/kJts8tyvvP9WgRW8hWBli3zhljWukFnh0YBGZav3IHFNKVD1mY1JVNJ
VLKiUjkKKSzEmUx1aCGTvcSe+zMqEYoP8MMKW97svpsHBKS1PYZEwWdCa7fP85Av25JozdZCFs1v
lnhhY/SLIKHQsbB/YqyuWpgwTyisTCisvZqSyySL1dcrBSXrunQ6AHXlN4uVeKPk6wggdwx1JKiy
hIPwxjW7E6xEWhFiTy8vP36WkyAdcGK67heCwQdeWc+AgKhPS7qQjHl2iYqHF0G0qKg0kWzJ6htM
2JE8+Z7k/i9FZuY+XXxZl7vGjPf5kYjNtC8fKA+2gmoAOjLH19WnnGXqZSw3Zhol9FNR2MEBCjhc
QfwwRRtJ4dLVAmfWZGOu9nSLvyC83rpW/tu2dTiJsL+UVAdsHTOOXkIV3YyOueAYshv/BiZVdlm9
e0ki53/1iWkymHjffI7HAsr2FH8aineiAssWCUcMaNDPaGmPWR5oDFonGXmY5JRjSkcp6XkFe95y
usL8j9vWM1hNqLqQsOYUk6fxrCxYv7LyqxE08Yo4UYmpjtsAvNCqvZSVBb9crpo1fuVQ3WcXQFTe
NCqtdDIPhfTQS7T9MbcL3E3C0nIXb1p5pLQRjRKk/1qo0c3dDksnwLD2GoNfTx3v55ndoPqtlotZ
Y/JJBm3AXAXnsfx7UWTIjk1LjtvG5/KxigcWPfo/MHuW/IPq+dfJVGU6bgWk2Sj7rKmJ1mDeOYiy
PI1j/zOhHo2noU4+GR04f3QWulGAYdiXp33R8pVE6DKA+LvdpHPY9UpHvR9WD3EnllxoZbFTPXVK
Ud+UmIs56fRa1u+6oyp36ala+ulYVO5sbsCOXTfQLLno1XhTYRUAsoW0d6S1Ewua7zl/Hgg6t7S2
mc7GOxpU6zrYQG4tYp9uTmeR9z8kNh9LAv6KD0+gLDelJffVUZFANABQ7lZB009/i5Gzv/1WYoz8
Y1aXjRuNFab1CSMZR0tjFJtVKbIX/YsPpWrtH+gb6AJKs8QmDAJb4DJpuOSJhsS3YkitC16tv1Tw
oqaSepGllYBh4mtXix+AwaEI5nRdPmrhv0OtRGuvYYipU2Nd49eHxxvpXwSLKmg021Jmojf9Vyo+
8d99VFzHJdV8pI16kUGgNeFnZ2T6OlV7a7ZoQQg3OZn/vYFcqWqeCwA2BtETIud+dud2vg8MyULi
Irh9tOePeEFWctYG42ZObTzHDWuqTz6XWhAWvTfj0orGMFa20hlwspMgYhjlSxOYkx7pCq+ToFXD
QUNcHmaMEXQV4i9TV7iigltBAi93WEo78yyaZ18f8P0O4ueK4QH4E5yR0JzzwdDTYxAy81RXCanA
2Ik48T+3+PX17PeWZXmxcThp+1fFSiqoe2SMP7X2nFS7tkMA+58PVZfkst8W2yVaib/qhwWamcEI
1ASp8LR87dE+gPidCWOAcc3V0sXH2hgHEm2khKW6PRmy6ZlBcBqzJ/7RusC6aIxcRIjXRUkxEG9x
2nr5dd5xdkBg8X0JUuDDedXd+mR4r+sEvz4qaVR87LUUffD80GTQRDoVBmJnzan2I3j61EEnTLDM
gaRn25QrAK60AFcbsfRaZGETx+b1p7GgcJlRJs106cTvQEURnWpWvgSDluqzaqImRlKebDttDqab
HojpZmQqga7FO7w2ZnwABvYpK6hfoBw5/w2ve6XF0Zx45KWkrPThCFenUu7LzdcvF0O5rkt1LLja
i+TGELxhrlCECxZX9lnc5eoqWO29TwfDsHDRlbocygAKD64ViwPP7fjtFnJA2K9v14VV/m072Bem
ogSsIcT9IeH9UbumqujsTnO/GyVW25A4i0kPEGcYajPDVKvrkjYuUht9r66zy+WfUgWxl6rBfBLo
ciMp1Yad8TGeMIegkqiSavsHnXcYMNwnd7EZmDxJvCRXM4CndzvQcnw3rAK1f7CU60VSNPFSRNx2
2IYm71zMHAE01QC4n4bdQo6igNnLIhvO1MOFZTQzfy4qn5YFTt8civAW3+Oo2RIg/1tM8V1zirGe
Wesi2WnwrpKK57I4QYIr/U51sFNwn53TPTJ0eKR2lkGzcZpw8K2OXuG/+XXRxu4AN67IEJqMuPYP
Sg8X/cWMhag4OJ7fK37rWoYxd2HGGTIcRdU7KuXhie8aLvcnYIWTM1+QpKvhc4ARBhAIFKn5Yt5F
IysLhz/h03ysDWrbaYUezsALzIx++k9wBVpTek2l+MJsc+dokhdJ4WR2Pac73X7S74j2tFB08GLT
3gOiAVeWLUzSlqhvTJXr2mkmIJM/uQOuaMxn9GW3clSW+GxqHVgON11CEZ3rZxN0kWezI2Orrrke
n0I7zgeYJNA106Fxc6f/YM5mmK0//kQW4JNnv2Pomlo3lfQG6jYV+dR3qatVprqmow6T4mRNFZ0L
CcWR8b6HNOH9LFg9qZe1rYJ0cd1eAUUwv4pWOoTRRGcu1AEnxZy8p7df5ng+NzzPm5RKbwVM/ZoB
Jqx8ti7suu8vIip/MNHshP5atGEm8IjOU4TUn9c9YO5hXeQpENjsI3qwbcchACB5PW//YXJPHH9/
gU+JRi4baHCmQquLltBViEPI27sEEeh/YISM5Vpd3Aa3VTD/JoqFHujJNPPIsf0+uBiK5wsAJA2Y
HUN+gfuCGICCEY9cxwz7qXfGTBt9nw/EQQLPCNFsJTJ3Rwzmru9Cbe6puRVMfYwQPAOwCnwiMOvk
agOMX5/MHyMdD/dajv0LH19pU9nl4W0zWfQiqRFkOrHD2bi24Izcs/p64q4xynk0yqaUUxSA4K5y
oMm9/rn2u7fLeDFY4pmzlYmBdMLIDZMXLlCdbD2JJGM+xiVtYWq3SLYbdnJWmt8Lm4QF0VW0WX3V
VhMA0mCltanzZG9AdSsHmXQwBuSC1apzM3eNKgSAPuIbvBPRpgqkvDg7g+FDVnw5IsktAnVNOG3S
pTGY3snvGTS6r7mJcAd02uLrQw+7e+LnX2WtyrvC31jzqem2Bp9p0wjzubGQW039OGnEF2aRB0NT
Ki8ODNocDReS7jWG9lFXJi3kTt+HesPCuBAvvWPbg5nitb6/m0xxYRgv7fv2ezpHX7f9IIOaNofe
wmovWnec2TZa2TE20pTLXPO+0X/OwQ5VnwpQqtaYaAod5boVQo8jMkDrcyM3mXxD9JFkqN4rJGLl
gDN+IcK2JbY+a7yWbYYgp1A5+GEfjKo9vhpjHP65PBa4ygm4yQ5icnENHeLBsrejmHxNq/BGaH+r
Vo7m1O5sfjyGaJ8QCpLsA4dNAJVKIngZFNsC88D8uXbKKzAxOFpgGghevbtVQNdo4PQH3rieBYva
tPymMarfeZrY/4rQpv4ccKwJ8asWMPX9S0k5wwuY/+Y/iUA8fc9VhOzbDIZ6iZko4cdfnKVemDxM
aTYJopaPG0EVfWi2VBL1HtF1xHGyluJPSNZcntmwUUsucwBotyoHD18LuF6RfuCud8kGRoFOpeRr
uA7a8STwaZzqEs8KlvW3CzCzylxVF4tMxRjG6vkNyErK0lCwBURKH7ZkhbqZCZQKLQsgAe7l6Nvg
GlusAFEWgW3fnPOP19nDuYUhqzBl6lzZGY6HSmnmv2/t9cSeMYcEybZQUpOadLmB7PvaX9NdaFCc
c6qnmRxzp3W7eUyFGbjqhR6VO4KNcGMZNWWen0VLfuOftUAWtCP6PhDLmhI6kgPMXYOucZQFRNdH
gev/s2j/v7xhWCckfJqNO9VqpXvtF8Uugw3jBZ+VT/hIM3aqia7yvchn/i5yN0i9WS8ivW1a4aIQ
uhGJgBDUuUFYoF8rZFh1jDo4S4m6lIBdfDXdtgt0ORdBGDqfQYHUjuUAuq4mPRl/atgg43cHEnCw
MxHBTS+3IG4/loCdfS5y8zboQ0w0gVpC9lH4qO7FmdI1c0cCDbvSEX3ZZeycXV1bHkUoOcpPTnV9
tdYaDYcMPCpMYTHZBVKRwV6UXW3cr5qZAfKv1KaCbHy+3zy4lmNN0wn6IEs+P70Q7tChtrbihYjx
dArQ7z7ciJy21DWVcf1eOlhRKjdagnhvqCh89YA9E1gwPwsPKbxgitFLjxvMeWCgK4WbvgwWbivm
ql7PP8ivCK1LrIPOJriClQ8K73QMND/n54SaXE+/yTIz81Gz5m32LpAUZP3wp/yPn5xfl62xwmg5
q09M0RG30X/BSDK96CLRNSoTWxcDoeglnsJeLLd0qL8YsxTPIf1cvb9cThZKgIcoifIDi01nnZIs
Pk/mRx8wWeufj/+wQZaijICdM2FSlly/qvxdWe8ePfWWqdQJe3Tdd5KRBbQSFlAsvmcxJ8oAoCYE
bzSGvLv7TKaeTd4oXXv0go4XnAvLsYUh2HkWNbZ0T4O81D6ertjKOFJsZwqg3cHAOIamvzgeJlpk
1tdlito2QlYIHTBWXLk4ya98SXZG+6m3ACYIOwy1cXSKjhimLspRom+ujO74qJC1uJzGY7uaYB3b
IEZFyRLYOTV9DgLf/CFOsJTVQOWR2C04B10CLydv6pSUXa39rKXaTbRi+bjHo2/Jj94zFQPTeY91
z4KuQ0pTgdfXEO5sYmZWqhmK16Ye19N6uKnXYG20lUpivuGwq56NIi8n181lMTvQdo2hFQhlBJDH
jxkodiHyfUJwaf3fXglPl/CJnpwcen8esBqtDTVxPrjnKM9Z57Aur/Pg1iaUpaD5DmUwAh9svCXU
cAhVsKdOJQm29V6Ezw8b41G7+abY+cmmNNIG/KKG5nKM0Fkr/GQN3c+8+xbh1rmQPVaDR/l6w712
3NHi886JuQP9jzr42zeYKTSN2ZDR1IfljnlXWm6H5dgonxoEIkHKf1yzAiwzTfXd2LAJ2wj1tUjx
qW8TMGxwINfkDr+hQ2vnkGwckqeRVQhcoM+6/vwNfXSRFw1D0VKurobqOa3VYPlXK5ZeV0DKYRpl
u6LpBl/u9sD/uyFjxiNZNgpLQXfsiRQr7lH/oCMDbIh5xZ0wrhS9MSfjqINEwoF80wLXZc4HauN3
2wIJ6uiozxPLx86O0dIUy5Zkjgjo34HCQquFD7Gkppdk71VGbUfH5u0BY3j0IHyxFLbRjd/MIdK7
v2ZxuLDq7K4aC/fNcWP0s9dFiggCgi/KpvPOZf6MowPElQryNPdMyKReDfFyZek6xBI3fhRLMPSG
jc2k/Z/41Uwrptb5RGSvJo1eHYvHMsf/kT3AabTkWrXkdwgeWmuNQyFKyG1JWJlcY5PbaICSBMx9
VLkJci7iuNNViQ0ywB6tzpdPXiY2LBBtMkqyRoWR9phpYfL2NcS4mKo/IruxMtJ93G9t2KQApfoP
rCKEvubjSQj6PyahMWTmaEgvYVkdAy2dl0f5pGRjPuK+xCgyirUfZqmU3GQBDOVUAgEIImFdE4iM
KyB+an3Zy4vzfVn4M+PQUlr2TfnmrZwUqlkJUgFdF/zTfy4NiG9z9Dmy1QBPUCxCzfyQsVFHk+zr
ldRUUxsSTRWMpnWFd2pbgcQbgCfC1YI4gGZjgieKIQT0kQK1LCRpc9wkuwTaxBqWiKadSOb1Tc73
tFNccK40GBWQjfYOetJNlatpTd+tK8HlyAV3rAmcpV13gTj//sKILuS08CEtyczZrPXSqlOXAsuj
EpyvshUMGgNrh4fNHWA29BHaota9AJ5j1fxo87j5xpbJXaGrkIAVRlQb3uwiZ7OdI6z8cG9Q521O
85e5iBKsOKauRU8Laosc2v5V7K+r7H4OAjj7Vt7+aTkj0su4PYIKqp4i63ZLEBHBDkgjvDgI3Jbc
aZ0jxMt1Mfrt92C1s1ZEUVWCQCCsFfRvWimWajGoPW9X59/TvuDP/2NPCQ2tCMDh20hFbg5Npb35
65jhF7eLi/wnPZn4lg9sVA7ybixdkCVSPkWoqt17cFpc7riLTRNeFs5YMUxcXlxVvo0Ug/Qd5bcK
YAaXcBM+l9wsFdtQFrFswg8ssecmBk1ePVyZKMkCXE78Sal0KgwtNSUBmwSMk5XpZIvZxJF9p4sI
dDNGsczdAi5YwwByrdOO5msxcXN/FMBqw1an9uYPxr+D4Fj8VCg//IAHFCnHbDrBtf7SlPZSQcSg
GRXgabEmOdumaBQ+oKQb83nfAshzmGP2yJkeWh9wficLEkjJ3SL7Yh8TkUHCRLZZPsrTvVicjxB2
RmHSBMTS3Titu/8RNz1/fQDk46I7+qyS/yZ1YpplkDSMgt4uLTUM07viAUSSHH1XnGLDzpnZCwEC
Sn0FYUB6XSeXip/a5knG5EKgpVULLvOVuAUym4qq1DcglUF75nptmriIiRFkq7LFgPsaa7hMi4lz
P7HAWjqH6fIZyJaJCqauOk+zrxfgD3Yb/V4B+h1qnfT6I7+rlGuydhPFuUc654ckgB8XPrPUhHbx
MTIKa2IWY9o5OfdnXq70eZ/S9gcNHuseNldXbYT3ZGJqcP2PELx3+96Z4PztGWGXp2wcO0O7Yv8m
7d9Es4jv2miPRzrKfCFn3AeeIp1d2wV7NgybTXUhBIVzFlKULnlqgwboTq/paWT66UV5mrYFv2fm
A9XQ+WVxC/5pE2qGnSO9PF5cwrGo226keksHiOAOnBzwCRBAzCY4wOJ6fkg8n4eol21gkWDzf2Vw
0BNgS8rquc0UIB1gNnsyiEBGO00Dw1QtZs/tf4vkrGXMOfCY5lYjDCfJDZknQTAq4KiSPDoAxfgo
UvOD/dtCisEEK8j00/G0rgRt6k2ut0NaYPpcoWTSsGOq5PbDduXIQqotvodxG6tTatejj4bb4iLG
TCQdOS0LdL94Gz7915nQ913cOAzfszSrHktk2AY0b6WWdNAvo4B+CJ8lJFoplfUrvEsQo8pGCQvk
sLspJIug/eGY4omjDHlRzoKOokNYA9aXolkYIUAzhG0jPR+ItIQx34M3Kj5bYO/frhP/NZdpWJus
nlaRaKR7kWFd/wpMmP4rYH9DvywixRDBQhNFhkTf2RjmDqlfNvjC0+G4r8gorzd0La95S4S311v+
HHQ4z8iPCOW8d3nHfBDoPQnZT4cy3lXgo6Rvi2np/1EBTiYvg+VgulE3QDAu0fvk3ETLSop9qDsi
uyIqmrlr9NW12Zj4P84RraGCRN/yUAzvo7wFTn61P1SIn5yc5OxGYuWFY0FcmJooSElaGFlBAqtQ
D1jZV6GakUzUBpHetl8Y7h5ZvmEwWp5o6g1o9+vSq/fZTxfJ3QR7OMiJVCUBsqQ+H0huqcJF2dx4
bTEr6j+yv6x9pk/gNeusGWtBP5GU630kiXZKGflhmoHmqvvH9obYkQwanFJfIAcK3KKUeCj0XajZ
14oLPEPAAmpUaR8gDDOamxXTzyhtOMDbeQuWyvjOyu/4Rv30Y65sRr5u3OVunVJu15YGwA55hc8m
kNLwQp1h66brxFFT7PEuw1KGnE46EOJAFU252SiKV+Vb697IKEqqojNMOC25tLd/rMRHJQDHL/m3
TBmYYOTTCPZpd9w1n3ZUbJpjVO21VRUby1a5q7+gCi04p7EswMRRJ7WJTpA/lodUzSS4nDc7ioSj
rylzQEWS2HD0fU94HuJTLGcRcgKIh2xfqenoAbSa5xWgX//HALnfV0anJgJRukBwHbmwPd7PN0sR
Oiks9EnlHO4bhrnTUmIAAqYyLlFfbd++vxGkqzZYOJmT2U7vNN3i5rHNon1Eb5swNqqFFdOU5nny
zktS5PCnW1zeajU4mH+G4SbZuHv7i4vCt7pPZisI6Zpw4v10G5WVHlP9XkWNJ2JXYR1PnkdpG5Dl
3Ji788pODYokaHLPQYArRL0bJnGKXuaDWTO0dIV9DB6AU9BSygiayuQUdpzes0E8p1vAIAzMbYYL
MlC2xFqllRFM9/LJ4vNRz7C9QfMmZHr82aMm1TOrXm4mJItZqurte3oQ3zBgtVBdpk1+w3lDEFwu
/+DtmXnjeyu7oS29ARRnReJLU41+gmK022CFHm5u3lcgtqtf9amCoCxvl0MT9DgLi11gV6l9xl5j
26RDTy6itcl3eCymRc/84FxywmL+unnUgwVDnNOliI+4Qs+q2bf2IKRImkkAc7laD9s+J+VQiSrw
lhUBV9Cn1iFGCtdiH/YOs1tCy1qaOAwvg+IcnK/t/q2YDrvSSeX6/XBnSf0B60zd7AtGUy5evJJt
MqzNvjrhBUvC6IZhCJPEZGNSmmH0Fc1eCCs+gMZ6dxJl/SjUYfxjWCFnyqwJlFE4MzHhg59phSoF
napFATkFN3uNyqbpKg1hDWMqtf8YSlzjlW9Tw5CnkzjXl05QxqzYR1LdBXb2qCknUMfQl88uIlSN
DFY9kqEPEHIG6rd/kby+80vffofHE6GqeT/aNEHf9zszKRMIHaUqj+0FYaNol3F1UYgB9MHm/KtM
vqppK4hLi20/YnG9qEl4ctnfX3kehyA1XcI8YzlKjVDeQShtRS3ZuDHxOSoG5FKJpDQi+rWN73U5
fo01+nalAi1uNE9x58V6V60bXa3Ch/hJpFu+MoP6sAtOcGFdLFM2nRTTiMiSW/SYVfDxAbHJ6Wyz
fSBIvdUbHEyNBtFWQLUYUO5FJiApJelyCwQ/elsNa33YmJjikw9TV66GDhm2Eb1d35np4LEFo9dM
2m5wJ1cVpupkLjW6ldtSgWCPg4+IsD6V0AskZAcaA/ldbSP9ee2JQ7eCC46EaMNK/fNw98gx0co4
anU8N5p2oDJQgDK8ko/Oak27+JODW/Nr1iLYD0GmREZIoMPxmwdSepHn37h9Lp1yTHR3St8/R7fy
PDT53AoHSuDMUgMV2oMmbzBi3CsC9R3B3m9Owx6Wok6pSNhTwEuuoG+FbbWfdNojASYiXA68D6V0
nL7gn1/9gGEf/g/p1Jx3dYChkkx5zyQMdJ+IcztQxOMfCDcwYPFWSxplY70dkrm/xRh1Op33d8Gt
r7N80YaHTAYnkrT7g/swI0RvSvUQVLDS0riI3uN2EFOSXoMyLV+HnCDiaylDSRoQlIXY2nsZEz7+
fSPCqTFA5bcNRkKHdo0HZQQSDoOun9mRL+fF1lLWMERv+XuDIRhxfFoHI3jLFe7eAPZD9JFOBztI
YcO3M5MsbFedwPRSOyE1PXjw+n56Zy2pL55/c7JwQfp9hZ9L3DxLZwFIcHysf0d+DDsKvxh4jpU2
etxK395EbcC9WscYzoXVXc7jzELrzKalZQuzq/+MDIFKEk9memkmeIRHXOtyFE4+KJIwFk0hyWIG
oaflvuFdWxaHQF41F2FmNPIR7gIwrrlaNKn52uDx2UNGPqgH9vrXPkpPBijVYXvTUCwePK9BURQX
DJp44j0oWHcQAhM5bv/+NNvA6hkGcCnxiW8wjMpgn6LjLlWRI0lE/cvKtJ9utkSnU2hdKmLCPBch
8ppr9KI6unnLAfKC/GZIpzWibt699S0BzWj8heE776Kdk1GqUDUnF+xqMllxMut+i5cZjxiz6jEV
z0cxystz9hNbKTxCNVUMnqD3jeoNUyh0PMNwIVFg9i2U4W6xX9Zthi/UjZbFUkYivRKOYzX/lC64
nITD3Y6dqRFMpUU24AynWRe6vQhCtzK8lfz/SBn+S2G9EWQmJ93BUqe8tjhWhDbI2CkYGPnQ/zPK
1Yv2FIhbMKCWCCxp897APu/qR5WoLwehjjNE3nEr/W31UeHQWtaTxieC+1klN2NNEI9DhlWWxX7e
GEmcp31teYz6iHG/S2kvdeBt5wvar8S3PkyvHyghBVhh3AZF/x0zUbSQLLrGGMOyNVLhz2IrC2qE
9DqcqiNmIpXks/VK1NuySNHW71jwQE9v5lW7hLgDb9WxACls0QKaFznb+tRY9d8Wyl8QESmmcC2w
g1EgqDRjYgYuJ1R5DpybmDBzG6U5xP1+N27zpTybvCDmvAHnGxNNgFsBs1F/AtcfCZxacgW4f+ww
f3fLWihfl6L5EFmQuGnxHoqRZy0ExEcZsk6ufcWtHe8vpB4AhH1ESny4zXN5Da5yQCzyFuUXFjKS
tV8v3yOw+quwm/k1j2ctWKMLGhSvaBMvWrYg9K8Js7w2JzxH72wbGw4ULdAcmeWiQeN5tulUB1Pd
qXWgBcfoKO0VJFIFOMgS7QuPdcfc5fEAjXmBo1aaEceuoglvIsrQYjOGc6bhSh3zweAD08ATInW4
QRSGNC5iIAXuUHi0nMyqlsOLL+9OjckATsKUVcHJAa09lqVNt1bJLPUvfBQka4Dd/Bi6dfrKfth6
TBN9NfyU3SJQUDtPtywpyaifFY80GZNJLhfWFrq19P4BkkZqbuZjG3t5ht0Zfjfp/u6GCQiF0vKB
BXZD5cJ7ZsOWFAFZdJ2P1VgtBbZHSqvb2aWdBbukrFu99rI5LFcxE0//jr64/l9BgC6DvX2gZSq0
arNOv0hMq20+aQTztDLPhVNPuCG11sIS8RnT2X8D/n9R/lauev29vln9vxkwDxQnVTOFa19CfKLS
12bj4/LuhOSEJ6l2YXN/GuFPBq2sd+PNY5qulSuYFgPUbUS5BMUbtkeZgCfPF25sF033osvQCAel
9NzHbT+TNCYl/Wi9hPF3w/3HJ0+BfsCzQbAAN9Lq7X6T58wtsGQE0bqNUewrDLBlXSrH9gokp7Jo
IHgJh72F6OA7yUF8kbpbTmFrDn/H6tqvGPi1VrbIJ0hW7d2+kLttQDxbeOzigXvXwxwgyrKxcLXX
UQnGGlykiR2hS7W/IRjMEHfuSyTw4cveqE4DD5NpWDeSQkbiu/s1Ebhjdc+umcqT72KvWtfCHGE/
v7MMakE+zUmwQCZq77Ef+dV5mSTQANFl8uloxiyWmZQ7ruvghhufQjficATxkzbXcmkE10iGQofM
Gqi4Oa1lEC9vI4uUWd4mXvX6xcoWDoPU5djZm6ZY7Rspmuehu35lgK0FfLAibonGpYziR1SSsV3r
GsWMy35AE5+EcFnLfKFS+PjiQBve2g2sFLU8hViJBjhvadVC/vnnh+Cz/zSXvf1zhAyB2bWADt8T
P7yeoMnXP/mPjRLtSb4jXiYSCynHGVd0u9IQhmi2ms/L2PXG/YakOUsCneJBNqochmKLuZP2KvVc
smNVgWAvKalvPdoas1PyGNIu4ODeYp/4cPRR6sqgqD8lcSD2LcckgO27sMcZvVKfd5FxuUi/bsie
ILFWP+lybWU+ccKZ1xrRk6DRhH3/5HMwCJ4B2XVWZHcJo5v1/RF3HRA/UdjAIQgpVNTfaF9Tt7u2
zPou148qzirO74zMEVMYhq8SphDVhdSFeij9TQe/aTAnvbY8Zk7NsQ2aFmtM6HcCvhiLZ0wgPPZl
Y3xd77ZyesJzZzdlnp9nsnfEsJXWBxezJ41Gr0ScY3bEjFjyY5Ojfu48S7vt2owg938abSz5zCVk
ryY2kypwCX7wZIwaMLVcITfdFCGNNjr25PvjJwCdg1A6sFTlmnTFBWxEi1J2sPaorNRnVu85CJtY
WfnzV9e9ROd26LARniodNB05ve4ONAywqiQqLP6bf+lft9IXV5rUTBKexFJFtbcviI7ttm2ENHFF
OrE48e3MbNS/EjQJuwq6kBvkp3MRiS2TAXhex1xZQZkPEbfYGOEMSPNCYT3Q4i12gL2In8KNrID2
ueEfSHQtioX+8Q8R4FkIHHErJ4IPOb8CsW239kt67acNTUAgTUKd8MLa0i16m2GCouplYXUlbx7k
phuYzdzCBTJ/YQM4sCVrhRwpExXYkLzl2Cmu2j9lxm8N1W8klF6dRuduoTWe7TWYoOpYi68/PeVj
x4eDf7G988+TSUOKNLHwaRaI4emYJBWHxhcjcBy7Ea9rf/MNYlF0apFOuLTQno3pVam+FvIXphFh
Njfav+c9ljeNndx0fu0PI5MztbvhCWd2aLXF4liLydctCW7yMsgA22sdRsxzWtlOiJ1dKXUmJxQL
XVPPJCHya0zli7wXP+MFpt7pBht/BjXPd0zinNW7vC0PnKQwZTTBy9qUYrP/DDFwXy8KcT9IvohV
Au8uUYpJUCm+tXI9P4z82X16kjU6tt+tKxdreQh/eBUh/4tchyYA3oj4ybLYxXRhDQIg6l9WoahN
PsiTNwZ4B4SOy6vRUx4n1z3TJMfVJbwmyXNEp5dQ9Jbwkx8RNl8GWNCZDJU/qijeXrhd+zuotout
pgXN3yzrgzE+HW6Tq7ZR3s0ND6AjxJGvxTujJQ2JEM5jTPcqTg1DwEWjpBoPQzncg9WueGTSTrAt
aRxdvECw0sFoBcI0z/k10FueuU1BIVbCHgTOn8gv9YC0zNY0E/xZMcah2uYkKLRBqMSY2vngUKQx
rTe113VBVi9axadMEW1MoK7VEyU4nBDOPHfauIUMhkDmstAoJJwPmrcxEq3wGNRWGkfGUDV3KF1a
sYoO8gkDnKiZ5bS5dttCs0iCUq4ecgFlHdfdt2xDdJvnTDJ4otqdm7znDB+NwQacUeBWlz2wTIwX
seaGNjltRp+go6L8Js7QMnYZVYBFo8Yt7BPfn1NOceStD+ZB0FfWDdSBgFckvUKbP4xQ9puPTTaq
Oh7lLU3ksH223DQqE2124HcCR0MYd768CGrSfSRFySEhv+rRPbb/L2HuyS7cZ6jSkM74mVfuhG5h
GoEoG0XDsPBmOr8JEMy16nAgC0JcTAwE6kePm9WZP3zzhePssQLpT46Z+0Zy1TfO/XAxIWm09RP7
TU0BHo00LBjmLLaddraRRffKLRG8v9MKecgRVV2qI7cVrOHtrO2I6bD0IZ/8ditvz7aMPUlSlQ9m
RdACoy5+vCNyDTEw2mkru/mn/RCqorWwwFTpvjoGvubCEgJEoonHsKMe5dDMV9CQAlN1/J9OpeUw
CT/Y/lLrMM36IgN9NQ3G8H444aVWUquD7mrgUxAAGsjiV2yg1HB0nswFgJf/4b2V7M4+lWLyo+lU
KVIYEvDH2tQ/l7UerPvhXX4s9kOuQ8QNa9A4wfGvaPbk8aEff/iGfnOsbQfRIJyIJx2KXROUZhAd
hhBpjBDLfwu6A0dAohzjT3/InrSDxKAhMdqTMZ6VPPVxqfUx476hwYWx3V1vLSvEI1ALRU7oJzbM
MundBp/6qEsztjHZPGUt7Uwjlqen5cTLo2Ke8x2oSGORwOMJ/HCUSpfRtz+dGk0YyjZTNiPuOXkr
eFvNLf3Ln3w/qJP1lIYGn0gLYCLNlKeOHY29f2RJbnmFXpNK+rfKbLOD9gha2NyOETdmZg75H+qf
i40dtiaXGuNkLuRKSC3yAXM7Vt9iW5HAvyengL1JPQaW/ubS33mQ4QL/X0Q2Q2TxTCaX/mxeB0v7
TlvV3WcuChEvpa/OGa00U2CCjKoS6IYokwCURDZQSzUL+CVPprUHvs2UJ/BGoiH5doDEIbXw1SIy
NtSKKeiA+S1KnNPcaQuzHhKyx4av4kgepWDn+CMdIex9UquOHmp2e/4e1td6veXzjy07CRNrSVrf
zVaXrIjz/7/BxIJ9B+GVDHX7iIduLM65P/3rFJWCbWzj6FLFB0BdzUb+Vwk0xc7C+QXcD8Wkr2wb
uYk172rMbZcx2EdOd2cdy7vgiyappqCNRy3Ffo6YMaC9eT3wOHoBkEtmt6AMk7iG8iugN5evnsC3
dNMj1bDvqioIHUIGNMem0Sx4bz55/bl/AoRWzpbkl+zuMRlV2e56dFlYGPBOduK4Yy0Bp8L4b47G
RazBYtwSWONL3zvjcOGjz8BdPNTKAAmzyTuKgeFWqdnCZ3mr+BGBmVPUkuj4j+q9quQxXgO6yz9U
bDA3xkZJiLMce1aydnQaLnJ4/3gIkfh+vfD/e2ZD/zwSk9kuO5dWDtyFnvyxLuNs9T0lh1iSwECG
R4eEhGQIIT8PHO+Uym9mxfWtzE8ZIVcgtzeTAhiH4RXnqmMbgUzkfaENtkb1X6Ip3T0b4qV/OxPH
CFCRjEv3EKsuKfUUeeOwLGKjfqIgW+BVOoAhVvga+MJNZfjWWDHt8O89Ff2ZKRvVDvFkLNu0wsge
FcsgiqT2ks598wyYedrrAUW3+wMorU0HEhoOYRl3lympVZV/Kt7/ujTvgKUBwoaggemU3Dh9mPgJ
dQNsCuK1kqkYY1QgOmNosHbSKv5mU+357tUKORN1tHycSvgC28uFZZzd53d03klRgwhh7kHh4PcE
4psy4oTWf9ORwkNQGc0RgNBxaD99U0Y7TpIshhL9fxVbiaT4EdLugAnHe9XdurmVm+7RJJMjqWiC
kn5aqUXe2HkQudXDGCtG/7NjNJuGI2CRovBRKr2KGFHD5/mdkXpOYcGFLjiwl21D6oek/idI35wX
XOCn2bJ5AUuIE7gndiMTs4r4xlehkmImmv3rrityI1MV/DC9tjVCOw68KuyrMmlzHJOBCKqEZIFy
pXI60LcBxNACKveCeYhKfmKcmDDcU7ObjRURahcGejsfQ0m++t3KCyx4EN12FPFyZYA223oQwqcZ
5UgTPrXm+lyLbyuAVFLCjS2U1Ccvdkj3tdsx9UA1dkoftJ1vTQ8OLtPGczHi9pJqDzrM1rVaMleG
qBbHf2sI+RmioFbQWzKeB1SFwXojze+Mgy7aonX+d54O8K7Ml5/C67p9g7LlanqjG9sqPtKPto4I
2Rc0D2IedSXSZeQGjJJtIM5XO/KOj8XAFZ4zLfhPAhycwZimSnMxxK6bsSvVQYqluyhjYZLOW2me
aJRInMtOZR+GwrDLK4UeVtJ3jg8FBesUieWZYy55tSwmbCH5BdHjEs3U7uC7bcUmXD0Xnl8K+XuD
Zvlz43YAgOn+IAOiPlYSk34B0T/LjtrgjAPudY+yphMcYQDXSlXhBL9hCxUNhmxXQgz/h6D4aCra
KAmSIUjocA5Dwsu+8WQS/0CwHlSxhitV/wtxzdsDbSxEW5Od8FcyYnzLvP7WRtM195ruU6zjxcMm
1krqMF7xyRpWVfjGReJ0wBQXFYIkH1oDzIQileJBrxrYW3pjT60lW7Mc1KXvDNEEfTV3wxsFO1dS
1NJX6eFcFgoulbwxo5Nqxy+85TFWS0xOzOxQL6QXiSAa7ZBcnatSWG9DHu/tHrsl29SYn3bbX3lO
UN+m85rC2mtxBdG31f5I0xPX7vJYRhGJUZNYOth0HnFYgskMjqewdVd3Jc3S2Yr6wbYvxNP5EUcY
JX8cZYzl8KUOtYOVViBs6sQZ9kjjQ8iTjP+7xXknCjaA0r0H6SwQUGLFZEYaPcF6GmelULFhbNKU
DoBfsPa2RZVWVy+BLJ95mfShg81YXj4ejJPyef0/SNTuvYExopwZOgiwfUOylUa6TRER8cItixNM
1suoms67RoJn2xI5qV+Yp73FQZitFDb9WOz9w1veVwSMFc+BXaHoEfzckA8P05k6Yld/8Yhk+jBD
fvrKB5KdiFpb0paTj0mDybvMCQgKYsU9JsQy5UkyiA2BgiM8fl0hAk4Azpj/e2HbMhRXYA3hPmip
fnMuLWgv41FZhkgMrSKmhEUTzemgGkBqx1TcEf5SlTVQIEX6eEdFsfHdqLxA/qlSWjvLZraGE4bM
lsLiKB26tlZPYIkisVjt4allZLs1LA4Vyz13fWE3YZpDd1M7iEfflWw6asREG6GEuGy3cJWMc0t0
U/EeRBD/sdXWiBPm0f4he4Vd4+f1rTppxHoIIs5IWfnke5oj6uWJB9yAYUsySdMyK7dPKWPZmTb+
twyyGotFcQkbuY+Pj+Sofy+YHWQmpzzsaFrUq89wilc21zEq2B59dp7vjJdNQTPGuPAN25WCA0tP
k2nLI2RFYw2dQ7NnP5Q24Aznu43FT0gGWQzqQyIAeDfM5mME0wIkBtC7cXlVEo0E0D9rmxYvVcgt
DrVzjVLn9ZKKyuSqjI4Xr72ig8Zfn9tuW39eJckH5DCgJawZTffcDOWSjbo4r9YHqVCw+hPPk9wK
2C1dLdve+UIkeTx3uLLMHBexaFBGbhp6fy5ETCx2NJS/mRuSo9Mae95d6rOfVtuwgbWQwgf3ZGNR
FsPXRElH+esk+d8NzamekLT0azoteDbYXkhLIJzw70QATmFA+rMLjiFFh+BHh5a5gCIj3ULPg1oX
cDkJr+NmUWIREc5/MpD1MHefptrB2T5P/7M3GxzJ4qAFMxzobpcAFUcWW5AulAKCxjPKWfxU+dsM
HKemcvogkLaMDSQXw5FY740Yn9bDHdsZSUiy0Y/+Na0GsPt+8kDg4+o810Hc3kOkCj+YyRCJb6c1
xTMXswSWcErtIBYYagwbhSdoRmc2CZ6OGtxT0bGkEyt5T4RhVi/PCUXDI6YVSzkYpjPG16eznHyM
tKu9cu1kG3YYUMm3On7+02zZQUDGXqsu98gnXXQA0rQ38mEWocDxPfMdYVahPGG36U+14WIuQGIN
jqGYhrsh2LaroTMRrQpdGIpbkePVevEvLF1/Y3WztwMV7MGKef0la0vYN/jWuAhZ5Xf2/GKJwibx
YjGCaGw30PnoeUYsm1cyvjHq4o8NOEic7YUO2+CEtPx0TxuiFjDzOmgnH5GTjWXndECoGX8S9Aoa
c2R03WfeP3ZNOLyyEuNvbR38tLjiVIbiyc0ElX4CZ57xTrSXglzFFZlGpnO0PfNYand6B01nvsLY
6bfwwYojP++aTkT1/q5Kg+qkkwqj3jJH1gWu9pRQiOZRQcnhnGpMX5Cje7mDBJatGOWV/9b/Rlpn
8EposIj7WBCjajY1vyJTlm+DmGuQmisY3Dbs+sZNr3zzMlSnkmChQZLltBeBZBCkuO4w+iXT9pYH
stckBHwIgcjiKl7RliGLa8xf3PsxM5owBbDYZvmSy7P3EA4Y3dvgS2FHmd4BmRWlU+vPx6a1M99i
ZEA2kzhsDy8QCVZy78G6fgny5ttXSmMMXRG4jdIsYxaQsUNE7b/13HM/bXvbP2UueS+TYjPAXFCx
e1VlENXT9Bvn+W+1TqvodKEiVCYy4+5Xdc+pD8rwVV8xwLW8f08JwUBALdoyYsa4YxrDTtbRsJXi
kTTJOWk8ZJjF6oWPt0AzIsY5Xbn8mR82YR6J9xQmdbMcYWs12O6SKy6a3/BozqLjcbcYI0Z592mk
OMZYNz+iAYXYpvtSCx2dfGx5blAyECPPGO2ZlQnrJXfN/GATvZINcIGShuS60TQtVkfxCt+a6rVR
3TZBGvxN/fOmOLQUSznpvP9T+7KYFimGbXmgLrD2L7LXDiAk52sXwmUwF0R1+7gSnt8ifEHW7LfR
vA9z8gAcbbdz+XZn00Yy+HV0r25eDAjnTlMkQ3y+8lCqa2SyGTASXGoXyI+NiN7X0Gc31YJ52AZz
CbxvnRW8qINEryhZ4M8n+I3Vw6ZJDwkBUlAggvAjVqj1TtxGmRMkiEirRT04NMAZbMp8+Cqdiwjx
ek8nHuym7SZhVFtgHsrhYZhQjT/9R7SPr1DMWRoFmpu9Pp857V0y+TcyyG9ZwCaQeGldvVbF3X9l
zL3ag4pP7D40rvN6WjCnGu8FazJMWFYMMUjyJgri1g0Rmm3zDNWEifY7S0hToEv5wxJUHXL7uyrJ
fjiqZwD2WnkI8r3ONDSX77wRFrfB3ZTzY6BPEF8tjEVRm3n1Z+O/9znIUSHGgHBwQRDspiHNBt11
g94GtuUccF+JHsf39sTQQVvWkVpiq6KEIKwsmCpleHoWwxJHakDVD+WMT6+Rub6IYkbgfiaj2J8A
7bcznbEHLrPOxpl0M0S0TCy9kChXM8W3qsYX3FiHBHQWYfQ74LYiJuQFvklcMlFqDDqJmj+Tr3Yf
qk0yuyLdcBJbpkL9mGVnlR1VvB96IA0y0Qc1WX4pR9AVX1rrZEi7hDSDncZL6l1fSDFoLw/6bEfm
CrN0pbLo/Q/M5qzG9ETOZAgcMAWZhgDBnpkI6d37N+hpaaVM0lPax1sC/3R6xQgiBAxanMLD6oQb
Pnjo+Dj1hOS5rf5me2bJOuTN5FqRi661A9YQrY7kxkROaNuaHvXmIiGendD/21TDx1Y2S730NJUp
kbNOQfhhrt52OC3nt174cHyFK8N+1te5O/A4etydCYOYeieAqzNreWIb6YVUGgBKbVZF9w6mFPf7
L4VoyCcHy/Itr6skM5jp4fKQWkNny2I/L4joIy6Fhn5kcS4N811hTpubux+VIwkHBzV1wlicoDx7
Lknm7oAMlR6HHNisUqDZd2//9ho+1H+tNQlEMO5bQo+F4yVNXh4Wz2OCwpEe+a9/DMq/iGn9+Frp
OSB87G3AmR3caSpabZ6Kti9fPsiaZ+w+xxbA14NW5/Bd1Uo773xfqK2uyGn0Qfi0LYG71D67zLVC
+3m3hTfbCmPKdqO5y0ZTMSTyx4dCCFGU55+gzqP8jgJtv9REkV7fgRmiRFNz/MuuQOr/4Je24YhY
yYw1MUqHYOPDz03JScK0zU/nRyXmePC5480VMpBOYzpk9004TpgDYGziKEkS85g8D6rBgRakTkAJ
0jwn4CPkwfnGbpcqH6Os8GUX4qk6Zd1hJ8oUV+qX5FywtMpFNyNr/vqNnStRX+NnRhTcJSc=
`protect end_protected
