--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
LmuL8z/NukmUvQxcVOkNsWgQNamZBrV4KJfYw1oNmyXybCwNtF+lv0Jtwbg28AomBH46Sz/TxR4K
1A5SwMzzUbmK5PvFhdOIECqqCHG7dRSX3r/81ec1KthxK2z0LhjuOnF/cxkZYFOjHUf8S1K2OVjt
tfHwKdGkxoCshSUq+nwwfuo3hhNzlHWyFTMMCH/Zl3r3LwYNWfDzSC053P2u7VKT7LBuvnUQzctJ
Pl8u36UZ24FcHuiVr3q0kyhATVop0neAw0XMLaci0+DndccOPxgPB8QnCk5Io6D6MF1M+K+Se7F5
X0GOndEkCgyUjOA1co9YGiVHUyRC6P6Uazb6Jg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="DzsXbaGBRbsiaEpNJvvdfR6BoVuBB+d01LIyN3lyupY="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
J9FFJY2P8OLwf1I+LeqMsrreJaBfzZOlPPhnocyaa8PXfEaegilwmev0j6OalLuL+V0C8DyzSpaG
ht21tPqFEQyYF43malJSBi5NxC1ci+zt/YPrAKVKD9cagQfLHGTjfjQusOTJsGOvs0FevRCN3MsL
BNcJDz5FpEmoS2oWTO7NfTv1UyXekTFoVkb7Nt9Smw90/Atsy4Loo2khMKfvt2yLxYDVZTkHgjv5
qvtWFS24xdnmUJQ4IJ98EG0JOG8ozzhxPJ2UQTww3FtrXVtpPPKEOH/xYHN8Jt01GmpYz/eS+0r+
30M4Z2cUa6m9cXfep5Nl7YaN8QiL5mNrJExmvg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="zyuic08uwcclQeGpd7TmL7uPqgUo0JE4mnbY43COKN4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4128)
`protect data_block
J7ZoJ7U5e+9yytjolWRGzzAQlF+uhL1S5bPApzEXM+ybw7cqB0PcxO2n29jJXDbOsZD6Bs/Zx+JD
DBzdj4Pjm5FFdM79ALdTqOkwmeyuBnj3tKMl7HnRYgc64hcPtUERDNHmG1SpgDIdp/rcXsf0nVSp
N0ifuNfFEi3lVmNaGUFa4u7i6H01Rv1yTe6oZ8jFqttcb2fcnBocumOlBm5ENdSyR/hj4KO+BrJC
8Epv5g3r5y9SMVar29ehfhGHCp3Z9/QiJKy7AgpLedqNTYNm7Afr6g3fzz+T8RqnSOLrhLRqDoTv
DWy9cMQG7PbD6XS/9A18dTlsHq6/YzhviamrZ8wID1rtdp1rcEVW8peePz/ygcdPDCa9F74gwQo1
jzqVLHtIGKQMEOX8JQf0gxrM1ixo9CLhnz+3/HUDtlAxRYXoZSVAtSGEqbhbAw3nlkhggazZh61U
a7Yg2Wxm1bDcb+CoiUBOrpr/HMKd4Ll3C3MkHJuUpkayyBebHWx/BSomJK8OEdZJC2+WEulzlvkg
NHBfeRqJfrLTFwmgCO4fEBmY5mvHw1C3ecHuPauPnLqOABvH8TA62kPk4W29kNh0RQwm2ZlsR/Ak
I0tYImD22qNpl18emVUCoyx6CdG++7nOH9P90C5Ag3Tmem3PAUDqVruauUGhe1wXv1UtZtgSfY8w
Gz/bqQlw+yxZ/RglJpK2OJ/oUXE0ZfA2ue9XJ0tSs3lSzaXeJdErZ8/FHR3jcHhdI0j7B8eubP7u
Y4rEWKYAYOxmzlKMLuJTqtX1nrKoUDothy7y/X7SvzbGHByy/yjlQ/gWziP3l1T2hJcqvbOnFDBt
HTy7CyskWvrHf1rrIkwJN7rUs4PjLZL5ds8P1+0vTx4nOmBX+5X2zAqoJe6HAQmsY3d/8YTf5kLj
Rjur2sIG5AJU0Ucoa2NZjvT66W0cjWqBDdRml+Gyp1rU8YoiKqfe7hycChzReIH+HBHK4Ty+jcwh
3me0GzRXADeGw6yMlsXhXnYQThQ5hyoSIWNpneXURa8T0DzhAQVr0TmLkSX4ccled9ETlstfYArs
kuV8MIDlTq9u+rtdlD8+Qi81UGG7R/yah5UYW1EeUyPNi2qZOUWEJ+4Kev5ak9mn5rC87umyZpBP
uUjyzQUyqANAAifuxPFyirvqk+1/GSOh2CSw0PEfJgooJ8pDZuT44U4SGglSK4Kj29m1Vnu2npsn
krbKWZ1kalsuyW2o7wvsNBibX8a0gUJqPEy2LBcMcc++TgnAdsfDd501FBYlQ5Hoap4DOdeyxxFq
tg3E9/MGeo1tOZPxaq1o3qdNKmyS6H8icDlXJKS3DSuiRrfNENSVtNXjw5XRTZ0tIUfGyAGZMEb/
CjNrn81afDz9TaVQTWN0cLFdrHIkBIqgdr2ZckWiTrVBuELacYXxQbr3FqXmEDUGmpHTnDP0SEFv
htKnn1ivWlrH+8I8MBiLee0P3HppUwTzC4tSiTmcLdPBlCTrVhQj1WFjII3QAaZLWC3lZ85Pzj2X
291eNIuus9oNK3EzdsCB6Zyw/UegddRmm7a3DV9akH6T70JHIe/ufrn6sUebxrJep295fKsTdzWk
NnGUmu7YsWsiPAwl+/lzRxXPBrCu4LBoyVvK0SilW4PUzSGtdDeiTof8rBTwolBjEFXG4M0/M1pW
n9lCR4vfzm6BnQyly9XKwiAzd4pgXcWsoRokYYRfkNUKvHJRdO0jXmDMiViKIQJIrwF/9+NISi3l
DtZVEn72Ksr1Humcfl+rKokiAt0tTbnWjOYKDvPkVSheFBLutc8NXN3iFHvavDwlbq2EG+ETE/B/
OtPQQnn1traa97FfUFYujHHY/3BysVXB7gbCl0im7Nz1Qumvu1WRo1IASbYq6wO3cgVO1Yh+tADT
Y1z5tSt16sh4rUwpZcfkDvHkb/skasc1dJVpeOAMGGZkJ0QroSlZKpCzw+ki1F32EajfZ8lyuC5D
tA8MoX6ZJA36l3t8nSv62exZ35/4Pc1eie+pBzLjsybZnyZKxnmAGMKTfGdExD4j2AgmD/dwmoph
NbVr8JsMVAN/gcYDS7aXTrRBi+sWJivqLMQ+fg5UhXCkdhGWd89/JpWsBCdzGQKaFT2f8vOyuGn3
AR4wX1VZBuPp9fIrTBq2Vr7HnJZ0IvIFgL/ya9FVU2ZcYKI2tequv3NQAwj7mxVjqhpMNPSMo+e0
Mfk3ArSpiA3ThL/UI6UwpvyN2InGBORg5Dqv9I8DN4MeFnZM9lc55f7moUl756B1JQ0hYoWYmAvA
N5ql2ARusdnYN3DcKRXt4u1bIicF54wFTVvvhhcCO3RY9WEoY/TujgiK5UFQTGo5ohnoduo2RFIE
/sf9kfebTr5hUjdYtGVVvKHYZ+3bKiwE7zIxLFRShfvNLnD0M31MNkO4Q038BI4IUEaGM8uE5aRO
rwhC8ZQJ+Q6fsIHXOk/KVdfx9Q3I+b8lJsAoUsbuA8KGkPyExMhWoW9zEuSiJWxGhWQSzDxezL2U
kN7i1ZH3t28Z8RF4GI91h07KK6QW8WQUN+3UfNYBr8wdFRkaPZ+EWOu0NGgkwhU0LUxTllisrplX
S3vArw/enVzbMQrUO1UmrakLq3hx7VtpHRLmZ0bmf02pydlRGhd31TTuRHkYbdslQzSlaLFBL7n7
5q9jHyFHM38WDwI19ST8hvlvvZPP19laTcMTGZYJT0Q7KJEul7+GRYQFcqcf9ELp5Zo3y8cnHasU
9TXY7y6VDDRNh82WZRMQHnzmzl5T+V9YyFwyT7MJ8bQ5Kl5Idbl4MYtXBVfMxgN2ZUCp2pqMVS5X
3kYdLMhlWQv3HsRJJ/78rxbSjcpYoioUFQlXC+XoAL6mutItgLgwmwTdVe6UmK3Hpg8mVn7l8sCO
0JrxQINxrROuO3MBSeOgsz0mqRmXZxcEXs2WqspNsf9UxL1YzaKopO4MIw8fL82y7qrsG428Spsv
G7W7Do2fbdiJeqs8XDGUEnHk4WEBX30HHW9bBuvKd0fAT8crIaRaGy9CgKn8bbG0Kvt+4CXGcP0U
S7eEoB7EMW0m4D+OX89Sg7fsrWx0eMWmDCI/VJNuKUd5SfyymbLXh908HK9vFV9ajxqM1jG1+5z0
sDYuB9+umC+SXypms3E8kW+UQWk+6sjsGEoE+RfsDTm9s1e8KZnBnpcc8aoeR1cc5p/DnAJPFEaS
2WnMVM3tyTWRQzBUs+zSBkd9QaDeFjDV489mWEdMUaEV85OFqVyzZMKl/W8Kp5B+8Iy2ZK1m61BP
9qrSxZSwSc8IUqrbtxfIIE9hYiGIWtpr7Ss52Zwd0lDT/kIDg6U3OwI281xfGyBkxedYRhJsROEU
Ycy0mwWbM/ljyYCl/rNkPPiExtiOJO5yVyia6KYeF6fvp9/p/onZVqNyHBGomhAXalpeAnYZkXNj
tFRXnNTQtzy7gj3FOZBq541ImbujDMn9Ei3rUZ71ezgZNc3OWPhRR3C1n7vtA+ktFwSo0VIEYmXg
MKL9jQp6CNinrwyCwnbAaEbH3JsSbcbwaU+864vNQKDKbUNDVzq4ZhBBconOlNbKQ0ReHSrste3n
Fue48A/3NyT+ypa8wVtkCTL+NbEdCBQumqkjrCz+pzhoXwFmFLTwym74GOMmwceZzlXAIaiWhnLC
SotlElNY2TW5tHEzezK9QXX/ka9OXVg4a5029eJ6ygD9tfK6Dca2TTWCvDSXOk9dnJPZYrRg43kV
WXlkBUnH1E6FBwziSREGm+aYnUzkMtUPZ8N9hx5aYmpqruISZjQGQyMOwsgarA0OtWY0ACyJDDyX
iNRSjWDkoDP7SXfhE5sMmWVSKxGju4SyLgpWwlxNylPECxkkP5kmtrIXF7/jZEsFz6dJX7JFOoe7
sd6MgJXxE25BesgkRSB25JaPAN3wc1yTEdZr1yY93U/yeEkVaj0Yy5Xfftu2++EHtyob3LW3Cctj
Y1aisNWM6HRSSwi44Pruqc7XwnabNfh0nyQrVj0EJ5sduO/8EdBWKq43668SPi5r8o0rsBYXmHS6
0RN52cKanu9Yp6vaX/p6OJy2NZJ2SYOI54j+YcC1rz2Upww/bgAVFHYDLfRXw72EkFGkmlxzl3gk
ISguXm+XKV850aAooaz/+nbB9ABmZdiV4z/kytiUem94vmexje3k7BKc934Xv57P5MRXBY9eUIJz
c5yAMiOlH4V2p+iwlkE44pLaMDfnFAkX5Oq/xVrBTd1YHESFLUecVULObYNNP96JSbH5AFGCknsy
mS0JYMqT8anxiri38JBe7wmo5Ni5S6kC4pjmgR3wK2Vn7sorDtvnKh/d2wWkacOaHFemHJSsXQg9
jgPfYLTc37R+zkSoSdm9M8euXjLDvYmH5hyjq6bTOsymJhEV/ycZuPMJ2NTi9S6picW6jVaRIr1a
S5WnjB4RcGhCxphg2CVtW3du+dxGayRogZPf3ayHbGvY8du+8ww+K9pJcrx8LeaWeKkCUs/2F4jb
ShBa6AmQTK+8AiVU+R77HCQV/dk8b+nRrrlQ63j36wXwJtJnV5QqQzW8Q5R+XoMcH5ekEiA8IQ/s
gM1QMx8/HKfB8rygkxpAJZSwApOQjq74hNukgpfGP+wul/VpcqV6q3mJyzd649IiqFyKdSUytRm+
5ryxy9d3DFvKTE17bkXvEsiYufEQRcXZ4+hSa68TaY+A1eQV+84mMP6tGkRhRlfkkbflWAz8HqXB
UeiCcEhSAs3GnYCXIDH2XPJZ7R6VtzxMAedYfcmdEvCm+R1PgNA+Tu7Z3tWwZP/XZXqpU7GM7Wlg
RgL8OhVnvgb8Nnx70nf1TPT5KQnKHxKwX21UkrHpGYvddYTnsEE7mTL05ZzSa2/8FcC/R/oiycr/
gPyq/JAqe4TEIaPkXoYhokjHuY6Rtiqn0nBnMe0XKb/eGdhtLadh4Sjtc4ScKYOHquDjzCcA/4Eo
aeqRbtOpY7Y5bQpI3YnhKn4SiILWgEEsbbVg0BUYq+pDcRr7zIzEtkqiXX/mIq+WxVZfM4IBBCvU
q6VsmrP9kbZLoMXMRz7/L72UrPVGEayYA+bye/OfWfM4JU2aPetwE8geyarV9AQe3Ao78gwOhQAG
ki71Sg6cA0MvllDlg35DE+E9uJGl8pwPP9JZDzgeQNwyS7uziWmj8Aq592GI3gYTGHeuVvqP4FoP
iwLfiMvbpNBVczoy1eUPRdsbg93F7tCREXArgegVEmOvXJNZtkB7wQcpLryOxR+FUoOOW8/lOJ98
ThMh2YrPpmb8L193OeyoVl1TTmTGcS66NrY+9VTpwjvU0uFixi2FhtooLmpnoTrL5RX6GP0IBQd9
BSsLGsy9/sKdDcU7KKwzU3l+V4hqI7zYi9Qi+NqEI2iBxB64aPH5CMl+6g5QoR78RFqbK1WbHRz+
joJksEoX8kUo6tF1vmmwKeRnJ+BrZISb8VAYpwQlgFL5wNSblRwFW2mM8JZ2Krhq7H5VjPZv+sv3
FMfbKdf3RUahblaS9DDQ5y+9DuIjJYO9
`protect end_protected
