--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
IembQ1jVwmN80F3Sy6Ke58N4S4B/jBJHMGVXvOISs19+IDVH5WlH5Yjty4lUgoRCLdpddpvznmfZ
/QUomOf91tP2CQvkUfG3uEw0j9JmpAj1HVWLkdiNUvc9oYbeEOFUUCUtxcTbbvHUrUCtoCg7VgVs
BZj0dvjsV0oShArqwSWhxjtv2rVqPFI9psDqgafzV3MDDuHum1vXzPMWL9++E9a4/8ljmyl/ZXLI
+YO+cKGRjXMCldljT5UH1oQtzCPbYEh4m+jWT6CjH2JVXk05YBi8LeqR/V6CacPo5rPSHEndmBvc
wnnpK2X6FzjazXmDGKewe/uESH4RB5PK1H2LmQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="4sW6N1O/R+RCqmonj0tyRkkSH1SqrXqzYlv5iY+nuh8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
AVZCd7UDwYLhpm47cV9oItBEj4zv8LHkScz0HoAXyFp+wMNeAPTd5X3/cXF+lxE//Z+LiLTaTXOR
LvgVdiwfeLinH5IiXA0qdSeheu/75eSPy0gWo6KRLubwjPNkEIVXJ2mW0rPrVVY5IbXgiTtQUOTz
gC9ZrzcT3oK5RdxuAJu7F8Iw/oQQku2gHrTlraUUlAYAeWTxM5mC2qit/2K/EITq3+khF7R5lwLT
Mnbd5jw+sjX6nNpx4+rKzMKpHZ3f4TkSU7yU5gcKA1N27o6+xpIL1CDezG4Bzl/Uz7pkzqmUAR9Y
8z8M+B9++gql+SI0oIJ3mEdhgiKTbx70UBAqxw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="xPky4C7Ih6gG5RO0USP3cTKolKEzOxLaQXB30a213MY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5024)
`protect data_block
qQ7K8dyYPmb6YiA5p284BcAwXD/8rA42YXlsdejV5vyF/XbKezh8T9VxtjhtkqJPkh26NWlBbMXy
28BDgs59VKy7IoBov6xMNX/uCpUT5hDirRqcE3R/hnYYASB6pL6mMyV8w4I2i/Gz0Y+r4ProWg8M
39xopSqxCqwrR/IgieRCc7FqwE0yEYiT+LsKIGWdiBmE+ybZor/yGkvZdGcSBwHvFFxD0XBkUz7I
fPeqJfFOBpavPNvJCtdgV4unGeSXctNDUdWNHtOp3lNB0Dn/tKflSGagPKgx/qVzHwG2pkRSxoRu
wZnRXbmSXu9qBueNSu23imgW0IR5YFwgrAO1l3tPE/wO4NgKegwUWEz4Dlkgho6UNwcfw9GA1+tC
GW8NaQT1lkRvmGxPFyS+bSe23gzx398V9US3OkHwu4PvefZZ2Pl7uwl+8ue9OEUlhbJjOwHvZoOG
fWt+pdpwnsLtTIAJZpuAJeVL3hjDZjHo/6qVek8NaulLlSjK3PyAeP6g1HWseNqxoPvEuvCV3bif
DIbvvpDE3nYyo8eVHK31qVoFQ+AkQLvnVur4vOhIW/VLWWK9+MpvQkA8G3aS9a/owXjDtHmQ6Yj+
0wHwyoynnGR0ReanwHyVGgUguvLTKzzVZZl+Ww9u3ctyeq4ncZbI9dk/8TwhenMmrKfg0j9q3wcS
jGNE26AlmR/9Aj61viOAh/pyWq+5CzF+xVej69CfvcOG9YHG3OO3BV0Ci5hJA/OkFlrDXaJxU861
JJAQ/JNbxhN4PZnGH47L5vY3GBE4L0Cg3jYWzJPFjaiYpkV/8oEnqzF2JjPpuhVSKYXt1hvf3/cA
oPmOj7IucJz8f7sqJKE5K8aqmycyOQwUIqhGvdGrkk3yessfn5dh4Oy0TTK5FYt7djGgADzTZauX
/qt0zcSohGBatemKN4hEU6Luwf8mbVyga6YD2YRHWotantvtjb8D3XtjIJwSZjnOBozdS/aiZn4D
pMgBdWjCsCjbGETG2p58cn4u2gPShkZidqqeCTTAltRU/AZRlhFoicvy5h19pRpbsG9JK0d+MNm8
Kx3oec9GsGnR/6NuEphRrJFX41vHHaaaXrNVuuINb+N5UIe91n2An5NPX3AdYaaTA3e7B1d6gIjT
Z6QJnrkJx48ANnO/Jr4R83Xi22SQ6CTIzrlPSHL6ntt9lqlWZx/4EZzw7GBWXMfHA2FM74h4nHfw
1lcJSFrjX043wzVyPhqCYqJJiQkZURwP4MSfCgJ+CHUnbrcW9TnB0JFrz62zeqr3aTnKDZ7fI/Gv
K/1WfMkct28GcMOGQ5In+y54AxYORWRUfs/WB8W8FszXAbmqM0jz+dqQ7pkFuEjnGMkixdV63m1y
8J74c7ElTOGVu8OQLK8e0IsG6MHpGLJXpPMu99kkn9jACDHw9bqyBmAUjzysmC6axnajSYzISg6O
D+tR+E2/tMmSs2rB3Z+K6Z4PVb7jo06lT0g+yKF2xOreyXd3VIp8DISUNwdtZElPtUMRMwzsMqPY
9kuQHDoGlfBocjwxLZhNDOL6QEC7J5lhhILt/qmuEYd/G+tOawNv/ZsrbKUjoW/14dqO+P02N73e
bSAevqTQ/FR+X3huuLi9jwHAzqE424XmVnlXuiNlMOMqZSHU18+HgAvj/Xx/powFO9hmgIhphXUj
+tfVf/McBnblKpl845PHPU2W2GHuE74e/JR0GJf79GM8/0QmgCsrkXxCGghcdSiDZMnuBXNLvuWK
osNHQyN43r1hdZWTG4DocMg77J/KPLXjlvyD0iGR2ST0c/DcaHEDbRITeJPFOw6t3LvSh0vinihw
KNx3mZP8oQb8hWoGBc342peKDOvKmTptn4YWflHJuYkYvFrTnWUKCAfm3RbyjAwR9mgXPPKIxteg
ILsSuPdk4m238rA+f95D4/VpBUBGkaVEyUCBa7NqTDkTjazQ+J3rrzuxbybSiKZrjfRhHSeSq3na
xFgLcbWP74zGcrPPSDRwefT2XY2eq58ZwEKx91ayVIuQ3WhMw09zZBObCTXcj4UBXjVBkvVUBzi1
mO0549fKLzpUFvrtn5etroinNWiLVPFHhfObBIfZJutBtBV+MVuwHoOnIkkD0K0w20TvzieRz4K/
zlmZlTCxk0JU5pcDhuhLl2pACF/Hh39r4Gp2SV3PYvygJre5R2Fy0gngEHwdhjVk5OJj2cAeKG8x
Ptj/hRlqi6+ieInc6NjFHUYwrwEAramYw11Z2e5sHc8ELGN2NtuieVBlKmqEpmap/46kQH7bYkup
zGcxK490IYjQCCxV5PU2hX9hYOsxvSvM6ZwK/V1iJ9eBi5VDRkixUaLOE0/rbR9IPI5KYSmtLtNO
NOyF0YoucUak6DJ28+rsqj+CRSs3tLg3JtvV3/vsaH8EmUQEL/8oKJVMrDxL1+OGBYhorwzrcjZn
fE8H+slfHfF+h8N1vfUlx2h/51zBP1OYWffweRQcPL09KlBIwZqEXa2jm/RYR0eEsTeiWydxSXJf
p5z8ZT9i+gWKQquUCxqMOZuoKlmNZkKSJ8DlULl8BK0N9v5FArMKvA3ROJ8DoWUHXIbTEA3T4qv1
eckpA1787z3to+C6YooKVYxdcT/hxqxy0AyrgloDilXbUN2vdmh4bLJgWSJ+EZxFDogbNwG7TX+6
w8NLuSeZR8K5S+/9Psj+VLDuwUygEKf/wm1d4CRilre6bT+4mNEGq8///2a+rtM5f4X7YOGUzsk4
56lRS06FmMvVDhPyssQ3a0jnvyD5BFvop822BVOOCjRYCtEq0BRSR5PTIcUmMgSMLJ1/0R8KzW98
9JQnLItlqgVmw1DxzbshCsUBEwSoJtyFPCcTDueedYHrwsSLqhmP3y4DitK+XvmC1zeRmPh62E6p
IFcFnUo9S1ZjR7IJSUVOzUbz1d9gJ0ZyGy/M9SawDcElBffWgoxTS63bdco2w5VevFfepZM9+X6a
Ogu1/HC2zXtKjh5XjoWu/Fe1VHSuShvSRVJQAdClLZA7nHCh8Wf4Wez3e4FDCNQI9Bgkn5zngxsE
zQaZQ6cF5DvW/Wi88qIsXJbhQo21BHg7IrTavYzK8ssfA2ZEZNVCU6Xo1Mh5T//6HqKtTxmqXc72
f7o6ZzofL3+a9Ms8sSryAjpqmH/caIhyc9m3LY0vN4Tea5oPZ053QKBnjl6crCMGOlkPgeUWFty8
sfY91fZc9MRJ6hLDry2homoZZ189PSXPXn9jjYRucwUr9nr02lvixhN0FlevNxXXRonh44IT7YYN
qvYfrEQ3WxHnA+FwAMYiWfZTq0lqGN8QaBWSf66f8uog/orsjS8+MsapohuKzwQ3RZvMFANin8L5
fslwwvG8TfizPdA526cQawrGWrd0KFx9IxgrdbsqBj6HqyY+6L8mJZpDhxhKLKviDAYFKEYTwasA
4mB1DpS1Yj2K8gy+HBptXaBEwow/Wnylyy7pJ2Xj0QZo5npBU16xnwDd7fSAd2iOVsd3s/skcrzX
N9Urunz3/4r9/kD1ceh8SVArlLfdljdRJ8HR/DpR0PlXzSYZtF/uf7X9InjRp9agLhlKnx0UenHp
fR4z9Swi0VezJKRhY4zyhBs2ANGE//HDXOtpJ45IlN9vWgct3y3pxcvzGcld8DhjSDiyWfd/kLjY
iUcgQXEsL+J9UT26KRHibMUWXcHC+2Od4+MfECXD7+f8fI6sV6TPwk+SmnwRtQWPpjpnS5PF8zIU
9SqyXE6809x+sG4Uk1FS8YWqqZtuHcKSd57r8vB8IDlZijzqur6Dd8f78OOyqLXUtFRfiCUzIn/y
BZmF0Wq9q2AeRAG3Xmqigji1fIVQQnYowcbAZqvZaz1Y5MxlDCq8eAKs9CoxdyBkcVwRQeYxMYFw
EEbCwU23ciDsdlK7RW61uvwsd9A5PXo/NOtamYau21C3QaJF//yx8fY4NkT47wGF5AVtNldRMhP2
4s/KUQ9GlPDYqjFytxWm76/8scYxRbPGtDO7IL+GoxDBMFw3rJ8nZgHBEPAL5uKv00DUC+jiljI5
kICN7o2wUu3rWv3HEipfQlcQh6qntLacS0YGnO3DS5TR7KInteQ+o+RzAgzXQp4V4E/XPJviQ+bF
JqoUvqcNmGNZn/IOCrEL/RFsmAllNTKyyPaoDdHv3BLM6/M7NkUD5HVXhfynIPh0wJkBYBmr2io4
CbeEMMOccfxijSUVHEpidkv/JkDH/j7sgm8rWVoX1iRXy9hrEw+MJjQY0UCtmiRij1FNIRRjNQHV
KTaSuLF0ZxnTUsdgSx0f9HWXcBQGoAjZTM8QyG1hNCCptiqS3fGXhRrAlyZoW9tVutQH5fAXxs8H
aZc6JtgKaztvvNV0/3euIjZcetO5t+NwihpNXQ8/jsjqSCjVrpEW776aRm6aOyFuTgB986QiSFwo
hjt51yRyxQW+f1p8UcIISXh4YI1UjWn6Wfnvr6pVTISZYBOlC2Q+rnUT4cpX2X65uMO06DomERpP
lEOjX1yxSx0xmZHSYeXbpBM6IUziB4e8kkYGdTsdpiHE/XG31G2ZYJXhOZh0fBDp6GXlclRghMlA
+Y0+Cnc3TStNXQ3rdpure3BfZq+Tr4eACHGfW4VDxSubBVPnFFnIGVPgEIHTAv7qZbtT5YMhrEKP
XtCO+MrBrRpWrMBT7zzQqzg115D2SnHF2FT/q9kNfz4UX7/1bQnLCyklAmDMFRXabwi22JLV8Gv6
ZTSQfE8zq3SYPtmA3RE9sjYOqy9cM04RKkeMygMivWc4T/Inah0W3w3TSiBUmDCdxzkUmw3v45aB
/w35cRdZouTnC/VG8H6+AtE01om1XOKWapiU3IRWhLRNDiQQSUQp/zj8AIVrLy0CBpA8gjsA7UzO
Ia/nDuiL/x1NiRKQlb2fSahLBKJe2xJb4/sB3Sone00x2vBwLnuan+4T/JuFP4SmfXkDx5SrsrH3
2NN/7JYG21F5Hva83BalY/75QlB2rGmuYwGRS06ZCGwZegtwpiwy0+dINVtYKm4SVY4nFvecESsj
ppVgEWhf5LzQpW7eOukgsPYnlDzBtw05f/CGpt5Svwdi3GI4zceibJiMsMhSkAm3AxWkxTqR0PnC
dH8kSmX6+LYiKRUim+C7Q/h+m3rXZT5zIghWe6qqPE8PRuvJEWE8zwuvcHrtEZDSkPqh1vr9ERuB
SI0g/whsEfM80gr3OrpZoncXMuMptXwrFXK0UMn6B/+Rcoac5cbPd0z4MHEEc0seFnnvZWVtRfW3
ggPiDxP81e2lnWuxsTmKg2V1sycc/F+4WlCUYWVov/72Ki7RAs2FaV7ks4ssDYfVMHvO+ixS8Ct9
GoDDjIhG3j/wwn/hsBnW+8l1OcH9k7jNO8Btf77vFY0pgkDz9Am3PNRIpxEwajlAdIGfDQKvEpxT
oHK+VaQ1IDVQuhLME0nLtzQk7TZ4dmSgLTz+tPmGbH2vlb7xq6DMmJdENowSCLRFEfZN0efuZyu+
T6PHDpDtrrZ9WdSQDOcWFm6A+UiGbqpe2u6KZiM2ZYkPT8mHyrjjqO1D02e3EdjKpFno0SVAdbXr
AS6vA4cT+HkCC3Hy4x0/ztcg/xcg/4nyVLAsCUh5WLKOug8w95DojbDzn/sdxCza7U9twGY6csZb
1rkXYFPPrZonE2eXQLrkKPsYSXAaskJ5mTBc8XK4M3j81JrB+BWJ8kyui4qxln8eD86KeKQ1XP+5
JqqA35UHLTFbUN0MmNm3bkCUIJLU5tdYGe+cwwmlcqJ77vks9D7XHVL8Ol9bcbYh1UQ3s3nogOHI
opHAQ0YWLvgF4TTPGkZPXHfD4s7eUvBI0WznJ1KragZ8CBlvrREDJNaHnT120mm+l9SDhIKtdE9c
ZQv0gxbg4NWhw1i1IpUhtNWvj0jEufPKENUW69zz7LN+7erXMP+HOFPftvOG/GY7XBa+HahWB2ZQ
gilE4vXHfx2udEsmWWQV1QrM/fMRR6oE1GeWEkqQY58g3wIpPB8hGjmYdf+8GPwWeg7rnuytrJbP
4CCb13IQ+roRbb0i8KxZsSyj9A6BA+kCMq49+NfEy3DcONr0dhB6HK1zRU+68e++xAKmHna3naOZ
b/VinHDUv9rLiNBQwW1fJ2z/+Ajf7u342CsoXJzjnOql4h0TZ5Vn0wEkk1W9BO2zWO8BAdWiR/CF
s7GWOBBNwQ2rOix/AUJmGJbl5afN5l7a+WQteaNsyvFoVqMYKdclAKg/86Q7Bys5koFu3RrSbDVm
xr5ZlreA8uDOUYBXACldb+VaI4qP+ttJ4WcxdW/Wb191UTynqcCAOmVsYhkkaR2KLSOukp1boQ+W
Mw5kbsmGGtBz3EjioPKsHIm9kRmtQ1RnxaiscvVoumcLQFTueAD9FH04h83+fcbnw3YOUNruPKlD
IiJJvITPP4YCNV1ampDT2aDi52mXd/fynHIm0QdVOBMjKjqjRIIlnCKVZYOurJTW+jSEVWa80fG4
kL+v4NHrNYcXkDfauZbioyLQUEnLWukAEDcP7K0VGAzrleRXAingQ3GOENlftD7gBxVFjhrzJYKO
C9Vadg9WUHYinxv1KMHqPr+RFWOwC7yhCiHbhgkAq5DzuePoIPEBCqx7tm15SKn9tGmRGdLl/Gei
8ysRc1si4u9yRfxUxbzrnFMELwvdKctcEpWAGv+eP61+W9dwPMbW3394m5JCxngPlEaGzWemibMa
HGuwv6VCEDE=
`protect end_protected
