--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
K4Bfe8R4IoMm4olXKt2e3zrXULWnjArj3ySYYQFs+NoBSodG9to1lAB2x7QSoW0it46KoiT39b0R
1Qa0Rq3UFF57GoTET+1NqIya0Bve9TunkY2hGOLU6pOLyoRmoljvNTrg9oVrEFdJUVVOHnJA19Yj
Tm/lOzC1Y++XTVxxk5VOFcBGvoDwBEjO8/qQFHXiPQbEzmuDtSV6/bW4F9kAYlVs4OS5ni36j/rI
sEIvnX1Z80wocr4Qy2k/uTQJpvkfgZsO1KQTgyLbZ/bL5cAwxKvGEMWKxFh2IS/7C4NuxitTfO3A
7WSU/5ikmbEZKWZaiYoTwE2l46UUNMguJjAeEw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="gzsVH+p4Hcpd9ZNE7KaqXsG3Nzj4ttwoQ7GWq3R8GJI="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
WRgwclHs6l5c290iT2knYgwZoIJBgxU3Mww3TOEdIJugnLvgAyo20vqj3y3fv5CYEZyXr9iOfw1k
aBSNe8arGdDFZ9VSmIcMhitSQ2H+OBthP3JZYXjhn8MKGQPjQo3RsNBLGU0Gfz5IpvcuJ/54Qtkn
U6VnJSsnCDaHFc4HJBMJ6W1Sk8uCGEdKrBboCNTXEcuPgoliy2ImCEPcxAje31YxsQ0L5l64Xlge
ykFoFGV5g7KTGppCsRfHBY6K/wUEku8OGtEqkFxPqWH0ergmyA+j0z8pCZjGiXWsKsrzJDOi3Hty
W67jShxvup/riRASBUBeQqNT93UFoO6KfcUIxg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="KCUgCmy8sYxkWSu168/QdSsOMNxWKBom/K+DeT1+NAA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14560)
`protect data_block
Ftwh++78R3GL6MMFxiQf8POMRpq6P1ZzzOyDkHVl9+pueZhDA/aW6ng0oAVkyAxOAfFwjZgZcgYW
vOqpMHOyMOchh3Y42Y10EYhqYoHRDuQaPybh2oEoyk00An2ENWQF65vnRW1ZLYBPF01WopJDHXnG
SAAVgj8XueQHfZB8A0SKzX1Ho/GFPLz6f92yrUbt5Zl38PJKbVi5oqugkScirQQHI0xMNIQiM1Np
Wuxdtx10UmDgwzE0Fnw0T/OxecupgfU7xzHT3lylYinjxZ+4+UKgpBOio+BCazLCYXNsBL1AWDSG
P91bEMxqIhXp43hpHNtmEnOMJN0NHMCjQTagfPoEQMmmFjJGOD1RQB9J5LBcSKAbfiscYn5H+AP6
uFG1CKRzN4ygwm8HCoFm3vjziFZ2ziwEgmR6DIW8EHe7Cacut9C87yPBveG2hiUMHmngmDyJkemP
cjd8YOabyjwuoxKfStjg1LPCKEuTOgu2lYhPubZLh/Dou4H1q1nTaVPUIQt4gNwkfjgSg2r8zMXX
qdR85BFLksdfW8eGK/N0URhO6JbikKfurHr/2z7ScGi6xUmwRcy7TyrqA4HyexquqmuJEU9s/4+V
CVJErAdUe649CwMLaoOVlubDJv1zL4Khc9iWR8a2ZUPKqCu7j8I0kwcpyfbfhOc+MB2pVLUscLVh
rXs21YFQ9z5JhQGxAQ5sGUlyrc9mI8QkpuJXurifmI5py+bsRALyhksgvuyHEypjvz3GTWFpcMDK
X5BEIeC0JHfTMGQAnjvWlI/gN21GlKWlgvERZG9ZCobW9wUOBhVR3JNOKvVGW+Bgbjpeq7AwFfDB
68ahLIizbm1noRueqVcXKNrw51ivfxkVP2G+APAAjLRQUm+W/QbfeBVNFFuREcqxm+TxZe03LXtk
cxutWXM3ouFP/dtDyKGWYTL5ZT2FzPIey4mTnep+4JFzLW7OlNmYbI0tzbJgj7nP7+FxV6wRqIJJ
r/lejG6oOLagIthVZAsrbBQKIDoQquTFVbiH33cIiUvOPVYoq0gQ22OSPYgkO+ulZKzVQlfSp1qT
OCHMnFthH0S+AoVC8zHEhv2I6yszq7IZd2jN9BXjZdON9tqZ2naXBtrk4YFdX09zGkD2LQpdEi8t
qRQbM3BkVZN2Oz47abKl1BxW8CMk4QNu46scOudshvuX7q19VZHPZ9bb+bH88zJP9at4t7sflQvd
blO8s1QJa6xl1V1wBUYoNOt9revgu56Qrv1tyE0F1MmeNne1JCFAk3/3XL2GV09fDyf7j0zXqOsY
kN/mjDekdiOnU6QdArQYz9cURib0Afhta+lz9chZsSQT6niqIuqgHQovLgpOheY+1bvrx8XBEa9m
Op1MyvLfGuaNPCD2lvMxAgswFzY1dWwCY1skXzaBcp8C1oQuuhH3zZe/Zgnk2S6xhtwpuLr9FYyp
jY8yauYyg/oF2eDs+Ci6uT9TPk9mgSyKSWCQS0sPz/ATtCSkE8GGD66ph/QDYv/eVgItVHAJR6Ht
aTar1tNz/IMT+Ivgc4L05yflKVOikvxMjwmhyRI6Benzn9b2MyirIuD0QYLpaKAvceDtbfGUl5bH
tDmKGMQgERQImdWs2cWec6gPZHJj4AZD5663Q0a7UGPsYOGuYf0Gqm2bGfoXvCdoNP/itMo0tsn9
Mrwyi4DXDJjAnK3nkaj9hzeB2tv1QMtUxoWjBRKXQtX7mKWResG5DpRKrLeFccRe8g3WE+wPcBcA
NG2PPGu+b5DXci0gUIvZ/wK/s0nZ4o/pgePHrLipfxa3/oZaFWd0Y2kkVXcmtKzrKyLkNVngKgc/
EsPcZt7JsYCJ1piAQStWJNOEKvFkbXAHE82f2TkhNc+zxW6uBihrJb273HkZQBvCBbE7FPNwFIi/
S1SVDS57ZHtJz+AHoTa6cRy3KP9/Ip78pVGiSiynUHyy7UAQ6U79p7BQFQbjpRGoJYLJhuYBngF5
1WWfytQxgOFC3eT8MdhC7AURAWP9osEK/jYG3lmb85uQxLUQPPBHJ4pdlYWT1EpE6rj7HkVlAn/5
cXGw0rS/BE8gSoUSw0SSt5aH7xUWTVzcBp9TxPQaokCNJbW1rs2I4y1tvLJWiGZ0lVFHzJfscQ+5
7nFPHyUaGEAMtW2dSVE2WkXRk7bRfV5AYIoAz3UrJSJOzAO/5JbLL6GZ1b9j79mw7smxdZ8tA3b0
fA5OyqdkyZwrgHr43/4nMq6iisHMpjP00Vj96u+W8zgHtv55rUNHIabrQgU8o3G4CBhqAtqwVmsy
xHquAMNoujOn3SmRdUDarUTCU2u49wXLrAhbE6F+UWm9D9uMLYGxU/xGf5loIncceV5RhrsH0GWO
vu9mb8AGLxY99q140sZibg5Unf3Ge58k/e1aBtjO5oDgc67DaaJtoRxrsCh4Iw1p6S8mvdnz7S0m
rMFzw/d6oKVBZV+uVTyH7gNPICYWaxAz9voKrllAMuDbMFzMGHRT1CrWAjvAnUOPId2JrOFgnkCg
ofEI8n98gvD6N3OdnDuybOXm3IZPaHRL7P12me0FVvUmaIS031Hs5FSJgdUPsC3N4A5rlSPL69ME
njzJ/60W8gQVt3N926+4NTUXjQ2YzIPRIltU9UdVv1KSj7lrj5Rh3IbOlGCCSyMQ9cfGET6XQzOJ
9rVeK60uoHgig++8+wxR1f54eODStZENnjtL8Wbeh+PC0SjCLDUfk51QbAglo7Ib0o+v1MRqWvFH
GeRmMDNIYtUao5jgs0kr2U42WguAlu5oih9B8+kRgj+M1vhAv/5pd8NLMbZN8urNVkAZit/XbXfd
bxNpj7sUSuUEhsIgy43DByiBbrkvfbLjoegeKPSLgr9yLhjLt+UnH/pOZNMEPndTS+pBnYA6iRSI
uMuQTV+JT3sf8NZNmnHi3CeZjVIAjVPP6WDb1FfdJQOx05/zuWF8eguQ25cmCq9IaewESWuyF4US
lunRkBtpYtIvK0aVpUxtn3VRmJPTJa15VlxrcOx5yBaeaXdeBpluaG72fTWLJsgKcf/us38uBOlf
Vo0lF1RsLryo3gvtuE1dI/B/8p/VCgiGA04gMuMENHAMCyk/XdnuBSIhNXOpcfx/ZtZ3KhmwafFE
W5qySO/peq1C/I4ooMqflkqIZ+d2oqO+Dv7Gd8aF99QWF5rlVCyF/rfbFJcuKMqRWLCR1tjHmHdy
zHfyviMlQ5hK1iViZTK9DlpgzLjLrIrOVLfcrrZQbQu7TcrAn1kEDr7551hMLCPyJNNJ3rh8TGsH
yX2I8loXFi3/RCmlrXI5RQ2Ky8iSuAIYoRQcLWzBFfbhQAvTgUvcYSVFSfdv/ajVm/s0Nl2c+vnQ
yux35QKLTriBkcYycPwcpEZoEd2D3+5iSxGEJrHY7yDzs92jfjtgMrN8AokarmXLhe7uezzDcyWt
YqWlqIprr5PR9KdRUE7r0NEA6UV2WeB2WwLV7BtzFZwTNKmTN8C1mf0zAxX6OCV7yo6J4ZwKPQYR
H6N4+tnjAzUHkQjGxM/hYSTQ67rb+VOYIB7yb5V5wYU5DHkhTlbWQjwFIZETGPk/xEiQpWM1KM22
iRDKfz4if9BF4Jmetnrz4e4TIt5/g2p+PEBvZcJHbCSUhbrBvSMSffdZRl6oWXuQQ2RpxEFfT+Ng
sk5UsfU1LD0gavQyLS2rzgw+9WyrFRP7DHOj3Y+GtlC0oY8a2r2djEozcYUAEXsiUIfa2FFWhbBq
D+HYbyn55+TArldfDvDSV99jtmNGLXzvGidlBXEzDmxITDn+LRHUPx4lo/C9WI3Xuw4WF5c4WSFq
xZFKL5S+XicdvFMkX/Au99OrjxvJFPg23ZQTtV66alPvRqYUov9y1bZnELZFeuz8LpSMqp8QPO+M
OTmSlbmW1cE+aM0sJS0p892R6Gt0jjSm5ar97BxfEqV8LOtfuCN2N1vXMeKuVzmQ5N2NggiaAzTc
QH7LqGFE+aYUD5ka71S7tsc4V/I0DaD1gDwt9wjaplADXICO6hToXs7QBk66AvNLrpXX/SEw0oaA
OMTy3LLa1Hj8bjglggNeJHhryWUMfFgmC2sMVP0fg94DSCIJm0RLoBgqfvps2VeXF8Jo1u8OeclE
sjIyzX1cZxFHeEY8nOcSihlz0sOzcb5PrHp0G4vlI24WimDk3XMWRe2bmNC1k8rVR+YILo9m23SJ
KuwKUUx3YGdOx+3TQwGzu5mp3N1W6Eu9SXBFlxKmRB//VpDPowqcX1tVZAWsO9hfIQ+07j9WN7Bg
XAxwNWCzftff2IuaHSwOdMrBN8mUD4ag58UrRp10u3sBwrrdPlPNJTKBNZWTe95uC7QRZXUHx1UQ
EDc17u3iAsTeo3vxfvW6GiNiEM5PtSO6SZ98eMn2FxPJshGtrVV97wGJN4UOS2MkAHpmTV3+/u97
qcojLEoRt3o7Uh6S9qfc0kMhPJeDb7xAHe19p4iPCDdOJO34RtlrulNcl/ZDv4Kdt82aWKmiZetL
NDCOEri/uqhQMWbU73QrnMQr4Kgct3OC0r3mtSv0+Mzuo2bNzLEVFiDVzf0JM5CbBLMuoNe6qx3R
UznTvrcCmBCw1RsifG4ewmCusYTAp4+j3VTm0LvALbub6lfyjO2PXXgCXpfcKjZTx3yIRsRu2Yp3
EmZmrPw99RfJ2tbQEpiWAUWueLjYnI8d1csG/yAENYvizSZDhbyuz2fYM1eh2gpGAvZG2b8HRLL8
GOvxb2APrgpMORGfyljHukPTu6yTcMW/Qz9YpD0P7nRDfuUKNdQceLVQY76lUYLSXqtmhXcMQb5O
Ott/jJQdFE70atbRTG9D21rnVt7VGb6XBhXIRhsMtOU1VO+9+O3M/rUyDyoGp7e8vJU6IwsPv8CJ
4aBbgYwwvjfOcEe5C5Cl4Lw92B9J1HbMfGELeW4m4khKa35QYaSY4ugZUk5yaVO4QzlanJMhYPIT
w5G51nZbsa7egGqiC7OGl3439B2iWVWL94rhEvMrnul2KQrq/vwf39FmoCpvwNcN3hwyxkrnd7Zs
RXYwJpTClQ4/yHXYtpXK0nvmBJ5q9nfLWFHa9KZPFkDpW0MABAYsql80+jH5LXDhznB4jZCZG7oT
UiBTOMb10Y3pjjnTAhLwunP12RSqAYDD69IaiwQXFOb08JJyPRU0kLA3qlhODRCG/oWXU6CMy2vK
PEgAc1wfC+wBo1g+VnWphCCjbHFCi/5LgPUT1LOuZbT+gR3FVh37obx+NG940515i87Apbz2uTHv
SgBcOZgbW2bk6g8cRn6OSAVZZ4D2oJm4sjGWRl+1H/a1HPzbYzTUQqko556VB2fUhB3p5eGVXCNU
WPSBDqQS7GY1DXoxeoaZhO4388VSaLQFhETxDeqV8gEMp3jradgWbV6D1D3gN+vYKErdCebkKfBL
9p/SkhYunQQ3XDO5urwrb3379lhXoRxDI+//NETQMmClBsGycW9nKD6EVhv2tswKkq3nxIjGGeez
0Eqkhb/lPT1ZL0gx0JcDyLvRC/iuK8GZQeDT95Z5XjFXH4p4A5KzK0IideY0e02MKxVdwToXDTYe
Ib5wvLagWJW0WiO4VQHeivnuei9Ghmv3ZDnBHuLqVlcqz7HWXhLLxW90V+PGVy6gZV8rT5BwuNIR
tQ9oJGEDbG+qXa6CaDhHlPuW625Be0Pn826aNEBw82WWORohRGPSrgRRCkd0brWRWGMPhrUW4O3W
mUnyx37DEfeCfHoda6mJuBX6ecTJxT1VK5Min4NpaJa1iBORRd5VlqAHlm0VFdQ3P0GN4ALMRFy8
SsoBiUeJsJTeIaqOdH9hZA/vP4HyE17Ar1BHUtOgD7KoNsaIpBODtFUeLX/uRgdEFoDdCHswHKSd
D3EXPTAyEf1BtYJZR5LtgY2jpb95ht0aLf5HgB0vnhTxfHVN5bXV5tvMcqWffxsbFg/zikwEPoui
FE4PGcvLHaI6xtCyFhECO+mFZfaWBJRiLuE3sDSbcue1knTLDOlVEPq6Fb4EAEFYctblg9B65Csd
y31aXzUxMkDOXILIaJn3ZwVgeFQgVEKF/f7UlZVsU2RYy69+ItFScNDvODPCWePtYl+8gi+OYIR7
upCIb1QgGrHge9fKVM4N+2AjNzoQwTXUYf6IXdeniVDGUJKGFW0lEWN3PARweJnHw7pnnDxlhVjn
lZxraReAqxv2EEItlNog7owI4uT874rgSY3sLeqn5/FR3iqcaPY7eoduEICbdEbB6B2A/C9XeTyB
M7x80GQbdhVKjHU+C2URtdfqYYUykLxLwR7WXuCKWPDHyMTtyW1qUcKX32fBdW1F17RpYJvFNzqB
npjMnkaUz5/D+tW2jaOHdkbpk0nhberBgUQzeFZz8PW0/RazNztX2ZQsE+1+x9MB4g5gRtnbdMha
52QPRK4ZcR8ipRjrzFyFwdlYrqCfqq2zZ/+3QQrrvqbtGcQTOws40dGMl4qpyB+XqjaSLPtWtiGA
2abOQxml0nw2jBjRWsHbhQTkvMMnuO3cPsVagBZVOP7DCVpwDg0DBrucMmTm66pjl7y9K2JfTt4W
6Ztj4QeMs2yRX9b8AjogNkDBpSDMCfUOLNtfghEx6k/rwdP6ivkPPb2ao9lHsR1l0C98AsaPwsHa
+AGxXxAKjLk/bpcDHOm4N+82U4fBhl7kxecuITzEky9U2QoJFaCb7v8c84CeoRZ7mIcIJLCF4NPb
bTmiYtpe7Zy3f/L2SukeV1bLQwpvdbFiuBySgk3dolnv9EWRtvWf6HVltkbb1A3cqD0KK+x9K6YX
roEv5XdnUna6qtelAQgGxAkk8SfNQMDYKCVlq1xfMuNsBArs2hmjbvyFRkz/xM8qygziZdd/1dbZ
KYvy4ftkd/s3LqFGVGTLrYUcyRBJd9PFOcFVeWD1ZWw8H55tFvXQpAQQmRSTSF7WA5X0lB+xUPmq
XSOAOAH6HEAv008QMIId05LtWorel49+GzzVJ+QV6Tq1bIXqAPBsr+3Hy1b2/6BhBT4mamnfdPz6
d3k6afC6pn3Zlfpb0hqE3hcECY8VCkmfOrT6OU18quwHMLmiDy3Rp9l3So5Q0hAR9PNWxW7XnT1N
Xyh3b07RNutNAHLQ2IbhCNsCfDwxbxZWHLCdTpoGyGQhUsetn502rENVpFAwrdt3l28pDZEr2vei
/PeyuQPwh8KK3SORgGRdI2AtXwowZfaXYiT+qaq54Kg5p4bmyKxeKtR0gJqKVuQW7kxzPUc2Jqf2
uz8i1pCn+M1FVjUwgVfC+EtERnDXMHs5Z/bMVteMNxCHMy8sW7XM/TfWEP00sNhSDFyAkSf+zopl
nFKrxQ1s7Jc4Vq8LWbzonMCDNewezlv02CulQrwhW1jdzji40biCvEjAitY8SV/F6od7ymQc91Rn
Zovd7oiYehZ94eMAphmpnXrxUbgD182s22tFNju79vsxJUKUU4tB/vyHb7M//Wam40C+pBCFioCX
rGZ4zxuTaK17TGPZA+knCe71PUmOcouXbL/k37tmO9/CHihxoksyJe25XvE78yzaKwfGFg/Axk7A
zG9sjHqpAbmL6jwFA5KXaTN1XSHwWL5Flw7lhIUrAZ/1XepGQN+IlYAZjsisqPSi4nyJYkK/qu6/
Yc4evhAw5wHJUOdA6451tDgOIz19g2dFCwQL9nKZWQu4VcUpu5Uw7Pmbl9LwT8e64YvCrDdUciik
3JRzT/rEkRK1J/hevo1xYcLJzOvQCdJlUHkGNhX5nvS+W31He2uVaQ8o1lLob9uhPOVi7wTaYLVb
ihEkiGQTH5WJw4h1m9hZQgSgL2IOHwWHMsOjTXakXn+vwpwW+vVSBRaQLF6WhsVLSQH77bylo7Tv
b9KVsWYvQRyFdQ2EKhY59XIqp2HTWHDasY9gDjjyp2QXbDwrYWaMS8FIyH2RU5vsvtSdoYHJcWWg
B5MBoZroqynzk1LXUuUqVWCI5S2CnN2/1tdlHlhoNNKNa2f1A7aLTFWsL2TKgBDmOA6D+2p/zjlA
5b+kSrR2tU42pBbeK0blLMdOB2mlToq+D7IIM8UjtM3u89BIOcw6HTzWu9eLVCR0ngN3aZPr18HQ
7ywsxVsV8MKneMgExFPhdc/918xH0XOxssE5Y9u2kbIDddut7Qw1n3WbhnU42WQEGOqs/Gv26Ynb
SPD7KJUbVEuzLqr/V3g4va82vvltAe9p5XESjZSDDa0WKWob23ojoqadwTGdjc0tc2L3aFaWsVgN
o4IrMqxQkHFJMEoACp/9NNwM23x2xHDri5j/0UCme1CY9S+Qrfep8Sgug7X3q6lOqdjrkATOp5dw
rRxx/sk/1DV/N9Qb8uNIKb5UWnKFBTiBaxU13JgSYbDsyIxAPMnELNbxiRh3anBgq5dfO2AYO+iv
dq30QzeKfcl9fMmKoyzL4kY5kLLc4kTNi1HCmHLK4mmQnXIiCQ64/+pEMffHiZY0DEbwZI8lSila
wBbOqOYzWTJSxXowmMSEn0Vu6hzrtU0D1dVDvrRpZiw1dAMYO4sTM4ZY1ZH1qBcIe0Ejmmf7wPyE
EFhKxqc6zokO1diXzRhTnAMZnt+nGt/5dD4tSNXNblfdgRBCQOfWrukD/yIFrnWy5JAdPh6jNOQc
oUB1RtgKBHt1XEdFgLFg/LXzvPRL9luShoq34ddYGAjt9ADbVavoXZucUOaq+MP8m5FhuUy1EzXw
L7MYINRXW99gG0AOfFByaZXD5n9ueqZeGp+9owHVFxsQjCcmFPQrwbDV+NIFLL8uGaikA7zG71Rm
z00shbfTIPOvmMAdn/DLATmOvix+jVgkyUBl895154gDl82AszVr+rPkkY+J2BqB5Xk1RA7x2Be6
NJeCqmtMU8reJKzE8sEfNPGv3Iy92Sg0IGuAzoH9evyY05G3j3aNJCKmt4gwHlE3sEKlLb+fQs8V
Nnc41zj+UGRh3g+kM2yzWUDCcW8hxsJl7VkIha6Xxr+xQrGQDm8e5IWYQ/48dTJLgfF3MV0vNyvc
xRAxeAnP6dJlOPKzjA03H3ycmGQWtSCSAN3WBYxqdgAgMMGDGso+IIFZYElE5mK1vzztUP4VJkKj
GhC0RJgwJ/fH5zqELnUfI7/7mVqb5O6oHos/H+/foAo+oewA0ACdNB6reu51Ca0bgyA5mzCfaulq
A7oOqZMSfnYWLOS8cBn9za4pOCvbmgxvsNfEtqUOTfYCAxXUFa2zKWTq8GBfZJ+eev9jeZFVcSWW
cO/uMKWUyvU8zlUnWlyGQMRzLQl9PSMGMOEMFZZGehqGHBieVfy+ke0FW0Uwe5sECmhS1vhM1LLl
KTR6yweRK4yLmSjExrujAmCRGE4RpyF7uNqPdM7t4uRTFbT0bJ+uCjh70YiG4MxcjFTc6MChQidm
g2AO+iTAtaOL7LkKsvo9wZT1XdwTfAWLXANrA75LQsJfW4AUxrsUVAohFoTNr2Of8qmiY2Y6yKis
LjEG99zN/aGb3cyR9CdiyU2vN4MkLPiw9TZrDiu6BZamF5/rhVYoowZOd8tTYI0lBbQZ3I7s17PS
BI7VNFFc84XjAzSLjt2QA9aHG8SWbMNcjZbFcE2kcNMv1ME9iLhMNfdWNWs2zQ72kepnKWW+jRki
aJBMdT2ioEGc4EEpUtIahR1MDgsegDXhAWDqh1ztjKjuk1Hy8NkZLz9gzfecLMLZKNwR93WF1BNQ
a2eJWeYU9cObQMMG/p5kuC9oSr5M4vLzNIuEYgU2cLeZD+wjzMePWQX4xxzaazgsHN+u4nr4FEqv
aT3+RfFo2d3++doTGqYBKBTyI/NRTsBbsI7vflmHpbXxLdZxlTRfvASI4hfrAyGZBWuST4h8oNC9
xapuLGpRLTjbs6QxmyUo5fV4RYn7ubpJlwvdgd0w92l1wPCqTnvvmu2NO+89TFf8WA6PyxiQObE4
q+U/AxnI7PAXvp5ygonUl28dpZg9DAJkoVIKOEUmagnpTeIkwAKjRUn52/AvZiUyN0CrRcZ8xB8P
cjnBAXKvWk4+e2/B5URsQfD7Wt9xq82JxxHW1f4U2Qh2XMBxBMQ1g4U3QoinTC3BP2qQVzD8mYmj
3q5fOFUMNL9pROrOR/gXtV7Xtrwwfl4G2J6BBE7tR49M1mSXBdT+jpQHLnSv4Sa0zEcVorSNm3ej
OJ01YsTJ5p+6dyC9HEY7hMlJ8uzR+Bd7DuNxB/NHZoHtEADD62cCSjblZdcqLqeDg0hBUeSlBvEF
oK4W/Y9hvmqB7NO5B9oskC2UZJJ1mKV1x5ekmwH6XMpUUWQfoKwyX/rKZCyi1uLxQF5dHmow95UN
mLbm5WHkP2K3NcPGAufxOdX7geP7w1HY/vq23EXutPWUveeElDS7/ObJ7/lepWifdzTQyAbtKLOt
QYBW3Ozr1sl4BR1HjiLkzAqdvxezhjcp9wzFejAJfCLH9bcXPjVITGQBOT6XRjUpXBecaKY7TWY0
e/nXlnJ3uR9k/94syObOmNU1aH+PfUWxgDQmr34X/g+KdStHiRJfLBVfup6JWXXZpGyh/krRtZiA
MrkqxENyPQyKchSjIYXpK/3Kn9asuWSd32veYWc0NotwNxBH8+e+L4/UEZxy730r9OymIfsaT1Ku
+k/Efr5mjSFoglib63gOuw3+m4sXn9Qa5+uzzbrwyCV5b7HiPP4NhDTwyGihhKJtIYUlnO2ovbnA
sBaQip4Dob3AfkY7zprhcNsh3c1YfOvBVnpBAbpeq4NaFZXwW+pXmiaihZwIUqdX0B8Ac98gL8BQ
2uMdbPrPu1f7h8m74A7KgQdTsxJBYiI/IK6cK+Cb7J7mNoLqzj/6OWXMZeJCVzoJSqmWM+haO+wQ
lLhDvETnT6ZydCRPHyZKJnyisXhL6a65CDIlqcKpQbGDlF1vY+O33msJZuV8V2fdcnH6spUB4r5Q
j+9oH6ufsZ/s5Ty16/p5dywuwNzwEnJqu8wLtxthst8pxwjDTfIzG8aMH7vda/XXzQuibnIPDTTh
ZEdpFALab0pmWiHkCFuc70oGBPmeCxH9WHZKZE1CCFcCLIMxSQlrnbGWDaw8oQEqaRYwV+jkdN3D
j7xUITdr9N/9PsZhSbSNH9xF0FBaTYoPN+L3sUZVct20H/P32IjpUC7Od2A5qFgC5sh2IxtNfCbx
uzCH5+EnCVBF406ikLVOLDnvMzJ6960T1DaS0nvsvuTRy3j4Q9a3+GbGbS2/kZenPCd4yFjJLAT6
qYBGelWYHrfuukEXINWjYuOmypbe+ADtYvhP6rnBJy02Ejlq6viGfLLQCuFmjE+w2Py+8NpBL8EY
570Bra2VabD8cCMn2+jZb/+ZHLWQAFNpYQnKdeBURM5TpFClwkFVQ/b47AN9ZNsaE06ttWaTslDk
0jOvdb9i8f31vaiVzs73Kt58Vx14P+gjz5MSb+1rthQPHqIuYNBNNFVEFpJTgsH/+ZDUj/jkQFiw
lQRfb6YTTlDhKRT48w72liWj11mZf8F8Eu/59u7Dad1uZtkksu6sAMbSzZIs5KlSGWyYDAdD2h8k
NEiW1iUg+SaoGWd4QoN9fUyX1fiVElWT/aqwEhyAM66j+xWAv/R3n9waP1x2tG7RQM29vYF2Trm+
3II409jVzkmwhqXH6Yde2IndIsb4A9NXz7vGxqbWPwFvBFtiehdnDiqb1UWpdIwtxYu78jPRmHoy
yPNFoVN+EiAvZLgu9Pq/lFYyhcAFa4ABbbQhzo77IxIqtl5xVCHuCh9gJbXYvscQaWL5ybMDHwkV
c/5SRfRS2JC/Rx2B7pac/3xinKHRwONkx4jYEjavw5hEJrTQQVoulNhsqDjdPUu2b01u7FxflYLw
B/w47OuWCGV3ZX+hYZ/dm/Cu+3KaE0QP6jy2bwTpMA+dtXWzTiU57+gmv66rEoZ2QppASMeUgity
uMFaWJz0cXPGNTUb+pDYK4eJ/r6LVVO96zvTJih1GpdKIbK0fylm9huEEV5V8cSn6Vmr5mY2G48r
T8givDzgzs79ARoX9XVXjyUFXIfB4eGV7dVv5mj+DCsJBFX+OGRk6ajM50ajtKLgG9mLVRZDR8Wn
tNUo3P9ovsDmg+W8yFoZly4NKQgZ/St+H8jeFbZ2DFMuGMdxM4Ie8pmROBfL/BSqBtu1ss38zHPp
wly8xBq9rmOeHXIT73E1KaZPVCGG65cx0xRyO1dnT4LUc64myDbcAfKBciWdbvWK7wxRhl4d6irn
mu+cN/NW23yKlLgDc0lFlmDtvQChHaOUvoW9dE6X7AHfts6RM1F7qVB7tDy9Q4tF9Bqkps40BQP6
+hzr+i+gUGyN1sSo8aIk5lwqV03S5zNq/fw85hy59rAyXzMh60l1OLRijuh6xQN06WNqH4BTVZeM
Fpr4c07N7mci4BS+qko0pg/mnhTOQTlS1bJcIF7a2d3uhz+xNr0fAhzVN7ppTEWb60feCqCdrOYK
a31eNsCGloCRcjiXZ5p3uVMzAXZLUl+V8IGPVqJnYVJUarpi+rIPtalgwKwhQvE0sI3yeZN/5Wf6
wKQ4MEmZsP1scZZSrXw9qwc0Z72HHcFyr2SrwTgjd8/pXaQ77MZV/ntDQ1BckCG4bvCZzsebUVCY
mzJyM5n4WmzFh1RQsWDSgnTBsGNOc1cnHSRNsgZDo+pv8sagcyRFnyc4UFeWZQTM63fCv+P62YeI
g43j2nHEmrSEw4iGngnwyOrhfcjiU47t8jbHRHJ1NPfLeOXdeQR4HelueeMrSPzqG4Dx5KefMOkH
j/Q7qOyu1jgp/+YKRqQlltAnJCNSGbhQXVxcO5DbDZGa5Amb8rQ3N1GE//f9jzDCHth9RHSqvbfq
/CV+1gl9tUcUT6GtaLTMFeS9QT7te/BcbtI01gAdQdg2x08Pyr5tGGd5Z3Ma7VSjpd8gIUVb+rAR
y0Yd4EoU+3XyVQuoA/6XYEmvwR32X39X6FuCwANEL22NZKMMa/H+MLS8SEl6TSEswlarlFLQp6Sa
nQYKakr7IjPePwJEC4ucHcx3PynHzwHAJLiRvAcpA+xUtolD+prGHS1/+Dym7fdzWTs3H3ppUMib
Lb6tK5gokoWtnyi9qjzfyl5ynOZpfjEj8Qk8KZoabp/3NEYgTNNAzSV2V24n1zk8lQ+IHC8wEqDw
fKF6I7LeTxXhUpBZg0nHGdfDvJHvPtBZbPpYWnhmNQP7Crg2MMTMuR+Hcwyh02H2UfPAdoaj0E8G
6HRoodizmF5P6GTzhmcUHPZ5HfX0YslauwYZQL+N36wmJHHAUni3/CsTaAReVkCUbxXTAj7USI+g
2HTaEgJq323Hl+bxDsmIBwLrhxNy2batNP2a2Z0WhEqKDQKSzjfpZBvta7jusSQvRydrJhV8gixk
au93+DkBeBX7jH8nDlLYzH0/hH3veY8GGxtG0V3MugT283bCLVwy6HLCFwlNj9RG7IJQ9REM6E4x
AlYYNDII+HUoV/PTk6sN0QF+ADKNhI6MOYzHmqpdzWOl434XxeyMrQQi0W3maX3wrtHbRhqWFlqI
fe71/M8iS/GoElTdj2I4YVwxHhny9kIozSQFuWZ/h94Q6zfu/iQhFyDnUOw/JiNFF3QjATSiGdR3
yk64vIHqUrtZXFYmW8DPTbG5xN6UVD++nw53Heyj+ipZylujtChqmUhhc+W9bTQr+/V+revCshHZ
hPBQo6LtqqV3Q5O2JlFjQteH3Yh2Ov8wqR4cNZYMn8+KkiYBOizrEt5s74KxdjEhDYVEBK87u781
TqSIHES0mhjmQQ9F5RGJvVIy11qoMzvNqv+bZTqsQGri0Cz+mHGkaisYzLEksTZOLhZ/YeM2bQJp
hxeItsLHidWVLdHjvLiANKgaomgwS+IeXwNqR5BxIlkQCi/Eco6YtEY49PmRl/cuyrHCI09PJF+m
qqMTfmsaECt8+LI5RYABS42O8htUJWTTA8qRTpidagTYUz4bXCa1hxinRJK30h3ijdh2RGDf+jvg
Ckp8S1nQDF+aZx6y3eMR+1qnq+ah4LkOYQrXhSiIvGKMltl1qtmePree8m15LR8idZMNRVjBEfJ4
bmTqJW9bS6afM/2iZ+zW+7vE2+EWvJ8BasdtRHU0SXX1+jpk9FgaXs0cYZ6VOZ0DbdMNl1OFVwF0
fhEj13OL8HDI9ml79ASPWshVXkFr4bPuBvi1aN+r7tUgFceKqX5M8u+/Cj6R9zwd8YHuE7WTKgQE
jAe1gAV2DbEqI7ShbOAPGude6XSlT7pw2jgpTr5VwHRNERskNqKP0vFQFarAUC+XJuKH0HiOtiSC
DFmtkP+hQFngvHGADejmCsyQDDIk0tTLWw6KPDbmdt4DcXSB9KsaphhvsY+6dhjWfpF2ZpRgJ/g8
cCdHuzfdKOWRl+QyQ/0IpPoIpmJmicAF6Wx1ked4yeMzkd/Wm+pYYjyI7/7ZZazxbuyctjuJInfr
AFg/mns5BKt7ioCliI3BV9Zc02NJWDHDcfnTIomyPoI5mX4bsTtyGyTixSdxmVh3VJj8weD8+vt8
QEOEeE1YGIxDmPA8LMYsJcZcVv8dIfX+Keo7WuAfHojG9SRTqb5P2oE4jtLj8zkVac2SJcaFW3xh
+cvKFaTNDguiNKfFK+S/BMv8eX2hX0BrJ+jgAWB3z7sylsEcDMuYssMufQ2nyoWb45e3c8v0PHz1
QzU7lMdVSxPjoKyGBY4X+tEpsuhgLiYZ2GViBHwViyF/JqOV3/BPtVRk5yuFSm6WJ8WHDRChzAVX
iBPGX2SWZSAQjDnnSDMsyJabH0xKlk4ak8BeFjg39bI4zsbfyvTj9qnl3ckcdSaPTut0iGgNwuGq
MQsc4kicCAKAGqLlVJ88Gj7E/GhBUwBaCKDwcAaNMpZxQq/y66BM8tSJzKF6/aBOYMx2kGVrrJnv
v6HaAssPMgHp5zjOcLMPrFFpAo490W47PCHKnDUJostKGT5lGpBs3bzby/AVhE8xXHHFlWxHaG2T
NjueSjlowKo+9n5J1wMmQP4d4k4S1VOJtvzNUKGyAC5P4QoNHnlAmrNDz+SJWja7yuhIoczBCTY1
DhcgkhyOWpqjmGOzyzbNw7XiETIO4hka4jrRUK5NZnAksQUQjf2Ovc8xfjuIpXQx++JF1Og3ncKT
v+F15fgySv9r+PVJ78wp5qbswb+Dw7//ilOWtZLI4QnhDvGFsDhSUjyTGI1zoyouANSXzUZuIycJ
3Qr+TovBxB7Rh+NTMc3lj3PzThlXgr6z74sdRQl1IxAGJSYQqtqOutsHvx83bKbqDavTsIVrZuYV
SII/XfrYhkNQwLwHlGS7yBrECVmnYipNWNP8Z4xUskyxEvb3LrSrv4u23js3jLn3nQSerCEa1Edh
Suot/Zvr9WKrktPoWjVM3QmEVt8WV9z58XLEtaCXqoEHn25MJEOl72Brccj+DlGMK9rZRBNyo5Wd
uWi/aMx3z0bBQOQ9CWT9XFr1oa+EeK2HwJD6rZSiOkqn9w1Bgyy9nKFu1UYjiWrfpBRh8qejceIB
QTP5I34buWdSI4aF4sAhZhQ5wBjQHR/kfuJtwVkpgr2HCjmIBxOgNEIaSk3GH6+SZXMK49mB33k/
0Ykm8Nzi6+lC9IdGNY7bj1XrAHEkbwkDcqGz5t3iz8+hmAdoLHqye1zMOPa+YXs8BgjuKT+hpqSm
jLozdoL2G7pSBZdYhOLg7wXjOcTYDG93Dy7ZyVPkZ0foiqTJ72hZ+q71KBUNb0e3Wc2k06WIqpIG
QSAbgIPcEbfI25p34U35loEbYMLg12kGliJPvPmqXNcqzURZOkoj4IjKTKagkTImtTFdj1O06zDd
AHVCFU+WSqHgoznBgRHiMaOKqOMa1JwiAkIlDDzTRoUcNroRnfc84KnEUTR2vQrQbPJXt7ggI5MK
cnYllhFcxnV9DKy7S0ITID5ZaR1Iyd1Ep9p587nI+jeKrVFwi1cuxrqdRpRTzm1LHBqfBM9sdNfa
7L/7BUw407MushIOIC9c2imF60k3NaTjQCsF8FRbLIghPTCMhIpikk/9qsXctA1r+H5/aqrADyBA
6BD0fvAUNC9CBWxWsOBNtTdy8mya4hZ57m+FV6aGBloDYLFTi0RJLocIQqBrcFHqopNNnVKiHF2k
osW69F+YqRETkJLCL69YThi01pFZXVSSrrCv/pDTSRg7ynewuOI35hk7siOo0bPGPYIFQ4sxAvQY
C26ibeoW6TU5lOvSiVm0/j6fSCY3g3z0q30hEaoDAmGu1oemBFdT5QCdCHlJNXxewCvI1E6mcSYX
WK+bDejq3Gb0z7Mezpvxz2hEAbc/4KorVLDKEoNcC0W6FnncDoSEeY6F3OjkSyLdKd4jvN4Z+8Do
I5rl9nrs3LpaVLMUyIHdEs2rD4MrpW9aQ4SmjsxatjHRgt1lCH/TRrb9byuaqifqk34xaviMUWbh
aufjKM6qnRUOtw4/jYoG0EUWI0md5/GbQ/wB2XTS/bbIbRtuAWPE9pqvlvZgBcVsPihYd4TfTJF1
AkDeyeP6RxuAVfclHA8wuIK2EWoRpf+ivBFFi1MrpiSGGbbknElatng4uECjGKdVLA6fiUQZ1z5b
HvgihHWqPUEicHpnYUVLj+gqRKQA6tSxsC/JWpAEML91Fhf0QrPp0M7Uiu7dx3IIHzx34T5s3MEm
eHjdLcyt5tRHoCv5v127ZPSIacTpTKieTbVfzMtHkGeatm9R09lrNViz8GjTkxujhMiKSLoTJAED
bNIep0mGcP1dgdzLNPoOCsJINQXb4oCuAWomUf0FUeYTNXxchEsveERXFyI+QICk0x2bZ86R/ZQU
qdw8ZKRhkUcseppE//2xrolGmVtXTmcUA7ZxkJwG7xt8NWSfM2HkamCIIhjNOR9iookKk17UY3p+
TMvEBJleThz3lyfYPHGUtLkO1wuquzNy3X9q+Q2UkhYCXz54RyIEH9tWuqLNrgf7oTW+sdoyscwL
SG454D2bNXxRdWrFw0RTifMFNHw7HEzBReG7YN5s1jh8FI+Ktv6JhImFoXEg8/pApzss8eCwDe7L
bXaH694JEHV9WFyDDEZPLEPkRs4zZ6QApH06dZdytKL4lOVO2FIuNMtzUSV0CUvfJulBhNJd/2Eb
41/Ec5yX3s96pRk+ltD1MnBkW2V8QBaSPedK+cozEjQ/xoyG/ACW1niBJ+SYpxANdjSThvSXrARl
mgItvW15ZJmo8jvbDeiESYJ8QLwb+QczNnrq730Ywci9SznYromu8bk8xDUwaiT9FXyN3Q3CyDYE
Uc41Lx294oaasd3tJDE/7R9D8lh9U+I0eY5vL/HDGpGM3EHinu1QfYcnhtlvPEvK5zPMSnbWU46U
mO2EUsdtafsKJBsVbXY8w8jsS+W1kqe1PYf0s1AAW3VWp+VKao10xuP07TtNC73klag1v4saEgLb
wb6jVuSTF5JpgOBP7MIuSR+DiDkLso24N25oa1zo0ROAD0vTrHw6BL4zL9mIMw9qHegg9mHl7Pxd
YtGNMBbyI5Zg3v8XxUjbk40wmsAEdcTTqZKwl3LmXx3tvQubkm6wP+X8qBow2YzLLMkF9OOe1OKP
KwRlJGA9KsIIpMFKG1dpCYahzFp/2oq1cfVbrRGPahr/8vwDUSb9q7VWa6B7TM6nHXh5x3gCRqiM
hYgNe+iymdfjSCoBqREdgeQpg8jJ4FOKmmmxFTpbii6+1GAzfq8ms4dFASS9so/skvQyJxkffmcj
0DpXsxqsSG8Rt6wuHH8haoUgFmsH8GnOAFGuvau7imdRObqNuviPerd+26lhenPyOSXUigh2PP1u
LTxDhUP7/vzCGpLLj6td9rJ+izNL45elQnWhdcs5wVls0UGOGK7bpQh00tjDJSb//j50hdY6mI7+
8ccIviTEkAlqjL9wVOIm8pNktcsPTNqCb0/r3jumFXolXEc3s1VS+JQWxB9Z2uEp4DyGB1fbMIts
XRJvqZaw/j5u+WnEdNYexSxoV/mUpb64XCsXcWn5IgokYE7HHyg55GeJerz+ngHh2TUKDlkF0ZMs
fKZjH3TbFrlvWAAgYn3cCFzafuNc7CQdUP1Mj3Gm5a9oobaGQUCd7Wt3BTkvf0Xig6Lzi9LW0/WC
HqmC0x7vJFRsAB+OGtoNqO+h+RRNxhxjsKuyuz++/EKjm9zTD08XxV+JVdbKV47Gpw0+lFnIO/wR
hU5TU8QcRuGDW0T2jejh4wK6aUpQZt9a1Cubm01ybwfPR5aDqaYLyOkxtPBNtkFekjCsb1SGtXYc
oLYve5F6mrnYPYegTCRx/dP0X/xDKoyiM8EBHTIbk7KC6EArcMeQxVCilOrnZwkPc2bpHzd2Fw3l
fQG/b//tSY74RJrwI30316Hwn6XSLCv2+9c3zsXVSGyra3JviK+0DWgiH68+fisXuGovpzc/nwqP
xTRi7PGzii+0azwyonGaRFtpeQ91iv23cFrDWeLipBv3aWMgTQOsDqK0IcH5eErTqGj/8Jg/juCn
yC+s21Cf4dxoaUNS3TFlsNrn+AuEFTtTCMiMMLNg0dCBwlsUjGn57cOTIm9RPU7RAX2p5Dqn2sn6
ypcY0cLKBGXAzuLXiBGWY6T3+sFKvn+qPscoToDTa5tUDXK1zshn0E7AZuvfj95vMPVBdCAYTHDc
tq2hpL3BygNyOxkcgnJ+5UkA5ixHxM5InHEPwYelhV0CnDlO7C+4lBJnR9xGBzWVPR52FrQ2hAcZ
ffNsH2zkTVOy26wXsItGxe5MY2Ic88IcYrjdS3r+RY9rUVxpmH0cZMzibzsft2kMrmjWTPKu8Lpr
8mVQI2Z5Y9yTznyQPVhdWfiqG835fT3oZyIRLetx3/ZdHzNIwdZ/peOC9Mzo/SeBW38Sn/iPz/Hw
XPxsTCahstNEtgd6Ah6/XfL3SAXiNiTfMZ1b29M6yzqsicTfyhhRxdB3t1qW4Er0On79Ew4WFILY
v1JQ0H8vbgFlzn8dtZE5ANgjQBNEAlsiauTnkr0vcwyCyVbBW/bN/VTgjK1hPMX5lbb4wzeLJSyW
RA5KD//9HfD+iww3hQwuaSLwqG8RyZB/Ge4U9+yBDYIPYYYGwN8AVEaAknOwtL4vkqfyjT7KA7zB
jnMsSkktK0QVzO2XYAwb3L6qURfasMx5ehFtVWdyehPWkkBq5y30gnHKTECDu2uItaYMO4BS483j
Hw5mVjzZwHlquNjNF5y6KXIw7E0UcwGhHEBfd1YN212gI81QfXO9kRSsVuWpzrNNg9arrcOAbfqX
BhD4SecMdvEXuQFt6NMx5GM4qvLkwBLPMX5xt0rc5x6wWdQYOUU5/OYF2RPWTeCrhiYHaKIjG+Yb
I4qg/bWGIADiyrKzK9jZCIf5GlsGBVH+M4cd4nYCVrXbfcqa9DqM1pWrpW1nd0ueEUR/GCeuqLO4
l5+J2JFrNNpZQ4Sua7aI8QiblwY25fISfNcnLt5Fv7mckoWeX7AuReMbkrnhR6yR+6IF5r4W8jA3
RVWXevWxpuObCpZ5J3G/6C6WI9IPi9l+zQ==
`protect end_protected
