--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
eNEy8hC5RmLXdHKuCW7xgdN2P08BACRQCZjoIgC/+6MnaEroDrpUGjMcaUg2IWyrim5ebfsh1VjG
d/uDZlg1AaR66FlsFtSezdgODQojYr5HZQSfnMGqB+Q6AoQK0uxc1He+a6eF5JTp8G4aFSq2LYyS
ul6g1hm+yw2ychGz/bRp0tmnx6AekW7wiN/7/Rg96KqdizlKQWL+xerghWG9BL4wKfYpy6ROFkYS
cGwUfQkBuP4s+XOjJ7ufXOX+oa4qjYfH2igvbKBoUbneTaa7tFdwT8KU9zSfYK4eo00R1zOrKAkT
EN2v02HO6/SDwn/6u4rcm3L2eOt9JsjN2x90VA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="W9uVFy7Fzq6Plu7/wtgC/bTmUxPp0kVqh2m5/xwicq0="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
CB3VTdI8LB0Xh3P9Wl6lW4TGBv15NO0O7WRm1OJDYjALS1eP0oFwu99SPwjtQk1vKvmsWatAAp4O
XIRoLxngApDZbywDfCVl/rd+gI0rX4DBShy3mYM5i/Fn7PxD6wO1IzjSjH2jj8iuQMEuT6Ikp2as
VJzE1/gkr0D3Qqrlyakq3yJAlItpl45C41Lvjl6anZXrWIextPJdqq8TMwJZXoYcAOhZFpZxmqDV
ZTcYKjCsorERehmx38zPgFLqBFd1Xfyb+Jns2luW+bXgcHlUJ3qjHHxClTTnMGoiSvuQXUgj7tcW
s14MMdrpui3is232Xwn8CGJ/nz6HaWDbh8ORLA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="pxthobHKAJjDw9IDsjn6aIJm0trjr+xwacPI7thHV5Y="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4128)
`protect data_block
k7efbEMoJRK2I1piVCKlU3utKUYaPIDVNigCtXpX739RkpIAWuGtwvgNZ8JNxiSPKpu6qUujuQYN
MISrs6SNJLr0t8tmoZxDQmwS0qW5/yS0mozzcoku3I0MeBvuGnnhVyQut7W97GMh2ex2S92aWt5H
O2/NFxkQGoT4JFjk18xS/w4ugapQfD1X9uT0c3KrdDLmktvB1r4DipMrTdMlOZck6JicMzlBvwNE
KJIhX5YK5OmPDNRMYT6AFUeki2Uu7QBOBI7qPkNrYNtRYfgNG6zvA3z7oaAqN9wh3l+YVZiTW/KP
m/LHX+YhIgadvz3C+bbuwYgx+4wFzYVNjFv4tspMPgGhuIulRxF4wpIkq9CFYWPpMXPblzotCo0e
aNI1DPRMWLJdCm+FjZz1aBGJ4xSv36ZFNRSHveUmZgCoEphuRL/csMqXhk2CsQq5Wigreb/Uwh6n
D+sdRiqjJt0zfvsjXFC+VsZgo6J4aN0xziYOz0BgLeITTbCk/JP4IAahMh253VtxPe3BMWXB3g6J
q0nyYRjteoMMzBA3zMEZiKjKwZAvzAP+YoWH1efhCZ17cCSMtvjNHx7sPLaN1vEaUkeiHrY+zwCE
TsB0O75GTputldzuEDUKJd+h2yJ6syAkUmacedXuTAZFNwL3EsTPSZ8k6LpWGUbjDNdrMWFJKsiv
nwbMtgtjYQP23TuO35e5zhVZrA+cHwHiFOOM7452ZjpTsoeliJ3qvmXV4DQul3LFoFWgC5KhWuRa
7xIH+Q22dm7Uxx8QA51zm9tOGm5T9zXFKxHWG01rbxQu1uDkFcV6iTyxdrBYphvb43LaKl3b/OEF
hZ8POjMbwFnBn5F38Bje+KxK0DEXfXBh3PVOtaUW3jDGYFz9uvSXUZ30U3ZWLbZC8YmQf0wwkilV
HO57DY2xCBmFqpifvyD7VQLuraFO8b1ksWxIiDd7PvElz005vJU7pr1Mpo6NoFEx0C9yY+wimG1r
Yoeqf0GJRfMsbxxzWdDlH6WlPHHDU0IYB0EbNcuBQeJY4jV4gOEkBVzsenxPX2i+Q5tvecDr9LhR
JuaHWTWgJvKcuSbDSHrKOzTjF5SFUGm0PZRDvf9YjA6qIfCzWv0+MNAuPYuCD8TEsFRYs+Oy+JHi
DFXBgxySgAaYt4C6G/Go70QbI3qTZ8cV/5kXEpbVsQv6C0HmSZ6qwhooe1i95r4B2JlG0xQpBM6t
5MbyvpKhUAhq2PMk86vBjRAPuQZt8Uu6gM2VuU5MG2R34JcnVdOALKreokXJ2G413RgzCD++xf6h
0D05fRujwTeRcme8Zl3cwm3/K97KytwvqL0Id8e3UlBh3enUMFdHIf+60BRSukrjFxHVg7SCVHDn
N90fVnrGSfWZHbF2bX4EnbJu2r447Xzs7wGuaFr40M1B9Gn88nIBEqiQod2uO0YR/3Mr+r9fKQ7t
cwjahCk9ztL3Qgl3rcB5ljPNzKBGZVdO5iZ50r5Zwmv4WNJ/pBUoQQYMns0JDwzMHhVgcLzV5cmn
YOOJef1VeAJ5B1zM4GOiISm/U/8UyGMr3nBKYoYtiE1cBvqpMw0iwAg83qhdLeUFg6deQjsY+6rR
bCqxXJwf6hflIlMuv3zod4mtsPusGBANzMi0yDluNthgEef4mwOirumEIub0XUJDmJxItEyYWkIp
1l2lhjjarwsLs2/V/M2Hbet1skF1uGPamfI0TE/usdUIpthMEY34nz9Xoq6PeCShPIDMYcqWOZUF
8/i5Jbjfjmqf7F4NByVuqBuWQOZCr+MsHm4YRTOWAuLspDaoCyBuF0R7t/gWEJ2VFBAhTQ5KWNru
/stEhg3BzrnOvhCKgiOnQBX4F+Dok0F3suM2/gxKtD310HtVSWA0NKK6G9jKYAeUj9Acf5H/jX6d
Z+3FrZj56OUbnq0td9UgT3zOVqFTLMpkHVkVOQTKPxUD0VLzQgAha2nfzErsd8Ybb1sJDfkhG793
ZcDVh3tNDxLuH01SMsisvWvNaFPRnTMjXKbdOnD0ZzAtd4QERuKXqpC9fiCNTEuIUHboSYxngUtX
mcYDc6z8SB0yciUofUzyDBzZQ5mk9t/6n1hO5f2kci4NVCPddP7yQLxXEYPVjYZdV4374QWbLBcg
QX3J27UI4xriBLriBnTUAKe5e3Ztu8NWEv/LO7NQdVsuip2nvXznqKR68c62MYlkFJgip1zaPDQv
LTA03omeT00U6bPF3VobrPKMwtWD79sKJsHiz8upLJ6aI9eoql+4/T/KByxcxqCuUO/gMXFaQ6T3
sOVOHF4u6A8EbVMkuhciz6BG3j44gcUCC0iD8p9PtrV41W8rS+DiCx1nR3bEjFPl+FuQISZhIidX
KEchuH8O0DMPX2/qM600s5Rc94CZUT+fhD7cjHlQ4qy4iJ+u1Vq3FZrIIUvidqz3knxEZA+c1/oB
QxkfNvHxXPLEp9pC5ticzbSAWLorhxFt+ICwsojHxWVuJNCxrbMXV4kZKwlRMqX9PNyTyK7hMqfS
aSUjZGOrfWH0iyfK4r5+KSmgexcYLr50wkkGl6s1I19z4Yzq3dwcGkbtXt1E+EF2MF9l1oshVWSI
nB/NQO9pDGnSTQABxGyWK36Ii5QlZCc0UI8Kx5qTljqJKWghikXfExtveVBUhkScz7zUW1QBjZjX
lvprU0fpvqwje11VRVpSouydYQPfcKamYIb+Ok0fGmfoEfjNio1eAlwa7SChLEZMQmKBzydi/67N
RG2c49AFGQc11SyqkH17dmnGGd3nKRo3CpxpmnfDQApT1s5kbkTqEovj7RaQ9fg1wB5RWm4i4IWj
BUQd+x0f/ZxAYDiQTp3RAKVsBMY8TLTX74RZ6W5L/xkQyxGmpZJfwqAxfz9WnaSXACFVHSsVfQ4F
ImL0Wi/aFFDPCE18eDHkm1jm0qMSYzc3ItGMeaRHzLmc4tww+ec8xS+90F3eop8Ije/gmp+HODr+
V5JnYNttyS/ncgZQ/3TvYCGEoUNXCePSlfL98u8N7YYCH0BUpHlMQ7ix96QTrJdZaBnAtsmOeApr
30DcsYkxaAJGTLTTxYkTmmStNtEUKI9Z+WFNho7bnflHo32r+WS3sIhCS/i/3cVoRI/wdXlOWrog
CRuummNTle/0RZDrMWLlZ26lijZZpE2YpMyLSwDsBF8NrlqjbeG6M20q54YSZmQi4imusu9seJkE
jn2Nq33X7Wj+d7EFQBMTN1ieuSa8PgUDNcyOO8Zp9rAE89USIyxnY1rKCnLcnSfRRQrNHvxPbnZp
oI4Lx/7ZCZ5HLVFfZx04eXp8I5+NuXOxdv3yX2eppPKJWafCsWNNTxkfgfQ6aeKHnGP9Srydh+eb
jrAvhjuWJt6rbxgFlxmNWgqXjixUWyas5xIEIRGSZn7R5mNV3BhRjw98NxN0augAXQw1y/1hhuRJ
MYZWl1wyJUBxsZChQEMNLsEOdWhs6sSqK8lD2AlwdIv5jVjoxE17PPLaM/Qg5VqKDq/4Nxf4Lf97
2sAKwQJXU45M5861JnyoroiG/91x/1J402IQns+bLcvezDQgrO3bD31ZjUlpl78la3B221b+Binc
YXVDyvAsutncrJINqbpT7Lk9yyauk7OVFNNlSq+sORv86uB0dyD+Gpyaup5rmIIYWGpJ63tcOncl
aLA6/2flGSaW0FzMENRDtQrZ2YbHCm+hN6Lb4fUFutwjcmcDERyCBhAxGD0xY0Z3h5TdAlmUHl/G
0l43aKULwJmMYwAZXIs7LPwdngphuTw2AGTzOsacm6d1Y22xGAgwVCJMJI2cSq9bGq/fvE1UMRGR
hRvRPqUFmvTEdc5Mup6Nuw9GorVbtiVp0gIuMmqI2e/DSdGUYMTH8G6KMGaDZKX6eKUKVRNParu5
Eh4nE+tSwa+7aHZz2AJYMRKw+rxN1SKO3QcD1446EsiuLxUDZFswtjDxv8ROO/SfDMLxQ+plfzRw
u6HPwvYYTaGnf9QW9XPavPLfr/YpWYi3J/ZPFLduyhXt9C0g5WeyUMw3LD/zFUVPm/Hr0oFu2Lap
cH4N7qrg5lxbaPJ8cee4pqKYhp0MRFMC2w/ARavqYksWMDmOpTKu/kOEHhmOEz/oWTqv7UJm815h
id8RBxp5aqxEKeOrCvFzEJXi3mt7qy5ulmg9MTC+OiP6GiOlZmzHZ2fJy8sBjWnFL1+xhJH8zBui
koNxS0qeurVX74rpZIp8wyc/pFLDaZ5xsJFeB8wdWsnHbUDdH7VxVttV5yCjgrq//ilFnID39ZEc
RzGFQyn9767FG8Y39Ev87czG848fZzis03XZuHgjCjx2MBvyLUTO/7rP0WAfwJzTZjTySV7LxaP8
zmmxWFoAHAdYYXV7f6FAz8D2kZd/FWKKiL3T3yQEkTQMTYwjyq2Q+/wP6jMhFDOLEVxE2t5lKQw0
661wWmhyMVMIVa/DPBSvOnWTmIr/YsvFZVEd2cXVnZRJtMDHkgA74S5OxlMTDNKjfLLbfaBbkutl
4E14GTxetsNFqf+Gnh3hEHxGYVPfvUuuPJFSbMsFjE4O09517UcID3V44VNUS6riz1TOvHARKz9F
e8dOTnUvIufIXa5YUGa1zQdWjPQanNqRK0blf7pcCK06FOdPP9F5bcU7SBLHNh2aQrswaz8eWrev
4u0bciiaNpqynd+9fSPDVGN2FdDHGWtJUvGY/h/nDnjhtFoohuXgzmmwIYT4SRtSM0t62PzGBMF8
gpcNPujpncgUbG99fH2Ko4UQn1lUOfFc5BajLI+K5BkCq+YvC6Hu/ehFHlpgMwkmgYJENyxe2/Ky
KgrTYI67rReiWSSJd1silYgz+k4s7ZFJLZ1fMoKSQ9mFYrfGtUwXADsrP3T3kvz6VoG5TIeRNa/u
tXeRm1t7xhENmrmgpAh+Bhl00JsRqdlT9c7g68ActqLhho9U51EcCPdQB9IfYKJ0ztgY6tDbPNb1
tQ4OFurYXJF3KVaoY8ujbD9QDa+MZu4Aqz0Bh9eYGs8FPJd029CRJrpm4JH9oS1TNgm0hvRk3yxM
DO4BUFXopeeOaNIb1VAJFOjAOq31xIaq1G4ew+cMTcmfrOydJCeVLG0p8GVWWJ0q/iPAQI54V6/H
ZjziiMxQjob9l5JEnCiqOa/HB2G7A4+IDLifUgNVWAkmcm6nfd5117ZP4u6PpHN+48GDKjYyD34g
yp0rjUKKcVmPkjrheFTpB/CjX9k1Waiht7wHIccE8Um2BnpsNvUofCmRgWbfXxV4aDKgRvEwGZNS
CV7elcsJCKfVctoPxsJ86oG+zYEBvM258j6idm+WWXlfuZ4RDSZpQVXNWiCVQaasFohsH+xw6nux
MPuyY9onuDx29qLnjLvUisdfAUqfegV47Rf1Lugm4TTSNFIfNZW3EbOEwtJ9mEuLvtCwAtO3b4eZ
1brIL6Itii1GzsPDPdouC/h2PAPUu0GhsKlpHGAOUwk89yXvUOymfhn+0c9+w1AXWBZ2Ws4VPJmz
XY9IoR5/mROp5mUoblgkC+aYvc4udUIw
`protect end_protected
