--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
O7pfONldwoB73cPg7iA/b6oSp0goXQ5imtvZUOBX/b8+WOIaAuqq7OxUDCUxdMwNbGWH1PDqy8FJ
l9ADQO1E15j9PlWabhNdjseU/TZQ7rtSnh4WPB7G3eZ+VzMVPx+Sf/3Svj0YROkkLCX3IHaUczO0
1KBiCb1t5GK9dvnn95kA3Uy3bjaa5zPSQ2fInf7OpKYW+7JtbsTz/jwBPKKBHfMqPiecG8F/dA7Y
nOcipPB/4RFuOK+YmnJ+pAUggbVxkE0bM0pcLl4oxMpdoGy+VbncF917G3vX4lcnXCpVFsiZIz+5
o7AnqlH6lfIIj/pRXy/4GrXBcPtEMmAOjdj0Nw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="qv5XQlbYiozPMqYuw3rRrr+gNxgFkTiPT3behMdpgzs="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
cZHmliQoITtE+sK+lB/x4xUGwRx91J+r1zNSby/XMMo6dCAwguee6368XAyZHfhHfoyHEVBNQt8q
RW4fJ/IuI6lAOEFJPOHUQjQtRDYevTv9F9YKff1VvyfnhGz66Zk14PRTCqk5X26lvzim3OH+0ktB
pK4PSreL3EFEN3bTpwCAgG5ofAXe41EiA+ZosKJKKoK3m0J5lLQ+AR6KYiUBU6vcRjcmsblWZjZX
6vBlc8uu7N72X8gMbAbyFV8lARF9ufFhJRqLuOGYz/i4X4fCiAPnmYJpBRbwk/opwVZpjrBTjETQ
uq2xlsVo71Lnf16iJ22n8IlIoUXkmoqqCV8how==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="XJgfbmgR4h8FWcIXKZikL4Yuy0oB+A6uplm0XPd+wLM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 38816)
`protect data_block
mwNkhAYiQXRyN2JALMqB5+reJFb2PPQNY/VAfKu9tq/Vl0JH5S1dJPO0Z0elFU1CwB0EnuZR1gKN
vzV++4Loz8DaSg2YJDSFCNfHvEV0gqGqorzK8qDFizF86m5eDbVqJsIenqMBQ75EcAG8VV46UCTb
+n1Lbkq3slWj2FlG9T305mMt6lj8vrhUw+EkkfvSQUjsVylrHjcQ/dPMKGC3zecTGX/lglRcXN5Q
ZCQYhCrWnLJXLPv3g5ub8opPjadRCIaUgd5uAcsQnFXXotp7/3g/kXMCnyzmDG7xAMKTkkJ3iMQn
D9eBZ+1g9H7Ev7cUBNiY6I4p3aL1TpJKb6jro60cl21LVQ3qTOqqqW+ESo1Umasxep/huizvgldQ
1wZHnco9mMU14ccopQIcocVpZS8jxbAk51jAB/YrM5e/QxlWl0csIltEK9qRQifDC3iMK13XURO3
t9kbOpaUzQa5aR44XU434fGKOXZ2iKW7abX2q+fl0sLxDthKrETe1TOkBU8nl4JNFi6umAVMG1MZ
pVA1/aPhSiqL++NkL55yvd9yIjEafqLn48eVikYlV5Kmz2YsxDokJLw5u/VA+lT/mbxiQBoqQj7x
u+F0A7Jqmh1oDNfxqXug9l3HoGxPgYPe7utgleQBzI4gEFhthqbKq890863aWvzUjwl6zgDZS9dX
5hneT7CTA0GFKhj7xmOe/GFskSmuFFM8WQoCR48VmzcRgtZK59PIvAevjuNiWkmdUHlXNcIYyQtM
kqli6es903i6GpvwrCrRXjX/WlKo37P0SVIaSnbQIdAp8bPI7Na92i+0acZpxlKTJ+h7OYEdBqcf
YtG5EQGCKWcUHKdIM7b4T5uaQ2gTvToEtaIv2p6TAKLcWYaZYGk+VeXzfiJTYaBf91wocbR+gnot
6Oor3NKD47UGqDEMqHzTrHpe6G8fUJ1/JRv8+UZ2AidVj88SjtmH3fE611NJ4ya7B647ALtQYojl
hcVqeF9Wj82RWtyPgOMB1BH8UBGHS/pGk7+x6dJ7ZKq/DuRlPgMSa0+/4oxCG4OjU/TL5jf5HiPi
fXoG1QIY8M3W1hyZu1iFYbEF6HCM6/EH4uqcT+FTZhUMQoTT2uMq9ABPO3WfeW3V3p1F7NHFz1My
qQjH+XULuGYqWB70c/HffLWrEsr7qkUMd1T2yYqU3vYxdMtaxne990ZUr375VSiEC0fWqan88uZU
QNqRiBMykUgXZ6stpKeusN1FcPduytEA2Ffy/7+az8SzKQZFEli9ijSepBgb6OxrAprIdQLFOv9L
/n8T/8zdgx/1lZ1N004382zquQ5I+ekk4pFTETcoxd+R8YHzl6RZsApaUzYCEwE0GROdT6vStc+J
LUAdgx4tFjPJwuk6zYVTdzPOLIWuU8fPweKCVUmPJiqJeYwpC8QWUNQ1lYn3wY5HoYlx6K6aOS8R
fB037WSyve4UNPPcPnw9o0KPsZK77P8E0x/CsOyU0RTUXrYittM18VPNhnsP7FLx/lsA7uMuhEHE
nckiflfHmiB3bIfb/Vc69VNDLPeugrTLC6JrNUSskwc6OZ+6RE1e8kxsb0gF75KCdBNhVr0V07nj
nomZbX6xlhdG8Fl7HpVDMGb4jZqLXaLAEUMbHimUFig1vhmApA5riIOf8i7ewK7u8Jtkntj8Nzx7
+V1Jgj64ROHSSWox6Dq2VH9cI2PrD2tdu6LInU8wAkvlRFukU9h1wWRJEXUUdQSGsueLj98O8PLB
Gbk65rVB6KaJqgm+MJGC+zPg2O5gN9LPnROV0Kq6JLA10N3kG0LHDg+++ug7ihL17z8UfbVlNxDR
YuM88XU3VhSOCavE2Nz5WNWWX2W3ghc3WL6u6jgwSWNQNhBWsXHwBrjBg7b9dsiOs2rTz8PQ4yP9
5NNigndUSVx2aCBb5sQbu4qhsunR0tNYhg+1buStr42FmNiCKxxmCdCk58LB1loMJuEpOQ/+VOAa
7+sR8x6pEqPkAoMtqBgg/m/SEindckzKvx6t6TXkOhs6CZkoV1C3ZYjjvh04aFtmXufzE/22BGuO
DMWQd2PGINWKgC0fhcTHbBaIengaN5/2mp7iIOwwk6hyvvsFd98y77wzqZPWCKxHEpH8HHdWgaKw
0p7jrAZ1o1TVBFotid5xNG7roTyedbbqtuyjp0rlEEvgvtmFldI7DDNmWNrUI+2uU32EuFtOIo/Y
7QIzaK+MSdIreaWe6JlK7wlpJXjxSi7j1uuW7beKcSP5XjEjUI8aCcdH1x56eWm3KR/DLVKlynjO
YV2j1UGxJ+KateKL1WgcWb+Vw+vXV28N9BmZwkcQBYQeyL7PInEUsz/e0xAT37Od+sVw0+vy3gDm
KPW/A3JlNT3IsPcF+n3I0Qx4VORJKUlWs1tsKT2lCescmp7y2q8EblbyFgVeELtaMPhmXdjbiAqT
WgXtW0CydETmnoZ+1PwUvIEWsuF7y7+F2aZ3+KjOjcjIoKeXWYSi3TVgnBgHf6OsituyxHdwIDhQ
qcxPK4eiybUJZ2HkUIZxSepfxGuoltYBVOaT8PywAZYCjCBBW74xKVnNMp6A24EoRCLceu6MbH8s
OwAk18sv1203BBftZrZkwF0iUtqFmZwYVFcOiGDekImkm7LTAIq5vK1BHMWEMTg5192/ufpI5ddQ
q/JAtuSKmJHC8UakEwhDo/yfE6dcWaFcE8Pk8xut+403OVkB0gmOFNCnxBmoSBa5Qo4ZxY/ro4g2
d8+H47knpdQbDNkY/JKNBr9pvbzkKvZoFFPqCZEBEObL3xtH7pd5AbNhMtTX6GOHa539bPTUC1/D
wMiWvlf4PjlqnkM3Dk6Vdn2Fwv+XOHFaQ8+bD8Q0fH8KXIU7/w/HEQSN69vYuI3rPOvWGUOwxkIz
pggRP8B6oQx2DdpI3P2FK2ydCJdyKhlQ5MXwXNktvG2BHjR590yj6CEnrd3REJjQUtBmmY3TbHmO
x36l8Y+kR/4Xo56/L34BOZ/vCvFYoYHnzUvELEpK24xNeNsJleziClv5ukl/5n5Ub/D8aBT/YclU
3P91BlkrCIBgNNLxPac0crae9xMvdWGvqoxSeMQJ8hxJpMb3sYx10sQnMp2ASRV4x+0JqLWqanrt
EIgaNC12UIpNCO50De+cxjEg5CqQW1DkkXlJphkAIXEllpEgfg0sVnwPp7xkz59zTdxaq6NMzoci
Fbf/a3nKkspNNqC7Nq3kmSHVZrkHkfrWmPgvzx+sQ5Jmu9TzKpQy0EmtkrU7XhLFLhEzd2PZw4fz
el0eCnUkUZQc0a6AV0rJxRWzcUKC3QbYsq4L8eSv13Yf5XC0svTHLM9G96HAarWtCUJLwhG1b1y5
aLfVjZ5HD0IVcCyExOxhpplM61NBdhW9Ji+ImMtMBWnKuBNXQS1hqxHgfeQZrFgGXWY7cBE2xDHN
DjhFP1rjoNqWe4s/rK7t5oGKaHWOIRCSRr+UAyC9NNZK0tdY1dOpzVoQQXa6Zfac2T8+rw378Gxe
nkLFjYFKX0n/khm+/Ue5PPc5G4fZA8rh2qGhBiObb6xxYHSbz9tvSEPKXxl0uGEdARlvnQT2rNQx
1GvKCNr3QHD7t9BU8we6DFjEfCvj0R4ssLLPDMsbkpjK0RRFIVG7bVSEOaQIdV/UkMTyWxM+d9Xl
4FH0kjTexUDel2oHIeKlm9F44UBBFxZONbMoxCJQcd8s6YctQ07wGZtv9+cCgVcIxo8D/a/v5efJ
OSMErKAOKSOPqTEvTKHCLgHXnzxllPaYhdVoxgw4erzQCQL6vRvSYTM590x+CNOndigw3cbEy1SC
2Vs0iK7HZS9K3YNeDrW08rcLCUsU4Rh1Rrp9V+KQPi6FrEztQgR0WmMBVJnvmJAyrIWyzoQVCrB2
5yw0uJkXopa/JeDB/aIdWVlsQR0quEXNlsRfNSxl4ghWtVvvs9f4JZ5XnS6fpu6HYc7mF7PgxWyz
WfSMb8hW3ndUV/1PGcpKJzqWYuXkwaNY/oYYp80/Gn7M9V+pVwspIMjRj8P/7QF+XWIpd/8KYrbg
i2T0xmXjqgT121S345t+aVhYZa4QjziSA9v7PPaW/SOwClozsR6+nKEOWb6kw36TP2QoUEZrjYYP
DmdLSt7BNq89XNECAQ3rSSBAEk9ZPGq35Qev/EBex3BuV5o3ivY+MIuD6QQGmGcFxBCiyVx8viv1
aSLVqSwBxSAkAcPf2FU3qtIRP2I4qAxTjzpS20HsrS1xQ+JpSFY9ejvmUPiU0ek5IQ094fI8i0sH
FkH7tHeKf2v76r+AVy5mM2eY5yqm4rFLzMM9en7OgwFuaTAk/Xb67YBIKSou+Uuo0vhTw/UHZ7iA
mKNSHAkMMyKIobTd6aMdY1Vtf/dz23sjwi23Lh6hSHN7S6La3NSroyQEz0X9l+Xqv7DulUfX8z7O
pk4qP9QkQbJtiBA4R3ifv62tMxFexos0IUpGhkINJ6yTH45nKRaazWy345zX94mRqDvhvItn+UEa
Y2eZp2fEMGUnLkb4Y3moHfKs1P5jsnbU2nQu1PqFg6lbrZ0mO/5Saoun8VJmH1n4nIkbHuXONI7q
2YBDydjKmjyr2vIZA/w4Qnragnb1BhkwLC6HwRZAtA2A1ItlxWeZhJZCqAtCBFNUyxOE0XTXokZ6
CvzTCCI1ElZlkErkphMoR4BeDJN7ucctkyQEpqw+/g9spu0ZQuaCuFHEVqROdPqSLOD2eyEqpc1W
v67gpRLLzen/ibFUHpAMRKrTWiGFnJLt0eKo/8eORUPsSZdMCuctZiVlZrhsiA811VOHZR/trJJT
sdiUkqoCBMXna3msnhcE1iE1TP3N1x4v50PhfGhqkSLmdORNU1bUmoT7OJUSGtR31j4NNCHjjcb4
oItuYX5pq0R/Dpb8klHHSLSHv0bkhrJcsGoosvxXv+yPwpT75LorDznrebYxFh0gMovYryw/MMex
FiwzNz8Sgqujat3JJBDdGebJ16FKYVAI4C1jwSg/f/LgPnd8fE1/u+w+7+g+eD9NefK9v1gtMgLR
EMq//pM2TUAz7Jifo1PR1hRe7fTceT2Dc7IbLxaQ5seTzNPMRq/PqOICxZ41qk30vtMhg0/srlzI
N0azK9h3Z5HrDA17S2Tm9gufPbbGHM9NCiRVDoCa4cuyMbChGfN20987NUBfwEHZ1WQz+wM5HPi4
BeXhornDINFlU2F0s97VqVSnOvQ1uyM9yePIYCSQXde459YOyJL74cpWJEO2dueh9pYPzRkSrxvo
a6VldUHuInAUKtwZamUBN2VzrWU95biQkVvz30OgmZeCVWMELBEh3cK416tK5ANSHB5S5gW3XqEy
reP8vnjSEEXxWLVvgM6isTcEmE5wzC6/aefrXnofoRjVdIcmpP5vJYVW6PdRQzDf9CAbvMP4N4Gl
bF+m3JPZHJBxWBaoMdLsvv+LjIwTnn+nIdX+4MLsE6/zfTiSvssnhW6BAbtUS9bcQ1pZf7EflyNC
EoxtLZIdLHuDfw7SCaewT+aI5tEI3AZPuMVxjH2TLTx6s+xHeNmg0Yw9awbGMpP1za3lFfnM2IhM
khnx+vplhwpSimGun4QEojrWnoapJ+ULOeBdruCMEM5mg7xFKvYwLEOfuoCHBkjel1yiH/+PLB3c
vOlWWMxKrgrXv9DD/l1WizoW8jf3M2v+KVia9CvwoFOmkSSOvPALqYR7YLdIKqsCgePj/jHeueL8
/Sg9kP/LVdhk7k57/em1dj5ULnu5AonT3Nkaw3RYYDUmDwHGMEjN8aF0LSpZkX/FsaMBt9qYWpRr
Jot3N3Hkxz8hnk/MaXz8lICabz3wjagaY+dWzUghlSToWayNfy9QfulkyP/YB4hLqWTyQIxVZANf
B0PYk4g9gsXNMdZ6ilOWLW6XBIj1SrZsQ7uzHck0L4T7vzke60QZWfIHs7GRy8Q350sloW+kv9bo
txb3WreEMN2CgXIr+1vFf7sl1O+D+c4CJgs0NUZxLNthtvAiaGEUJmNhOGQdtzwDmguW+cnM9d0D
M80fEkki4JJSV7ArVIPAQ0jS+mHj/2bhklhD+S6uqrN0R5gMkH1wlPZ3yRMpTza79cjyMpDw+hse
R8cmf0anD6pCFERWsEIQiy0eXHuKk8i67Cgo8PJ5Bt38ccrOAY87lssiWH57Fji78Umx2kGLhmNI
R5zEPB2PR5MpOfzYDeDtGQDBzdw1ximu8NW/3/sS8+Zg1SlRKKWhFR/0mxcd9ciTsBy3HqSQJ1Ls
rQ3SnctoI+XwlglmlP8TDqWrszHJDY8lYSA1FEp75fMRQEnfqjMwZ+0ezmBGsEsuR6eNLOFIczh7
YUjlKkUhhiDr+TTrmmDidQl86cUjqV83Tp1Ca//hn09lXvz/v1SVZXg4bS9gDrP5ap37wr9itJMl
jN9Z05DQo9Et1Z66EWWXN37a9k+RCUUtGB5F09/OSoCLhpYJ4TUrdn6HtFLZG4UKOwqvbMuEwPsd
d5rXv+f99vcjaiHFP+5za/i+q81cRdTOWvNW3EJq3ngb+zfLnonNRyDXrsVuwHy1FWkLSpM8188G
7IY2kjVMUgmDEUYAkR2tGiP1LbcGFk7RE+AJyuOLk6q8romB5TcmIjqEt0aK67+c8CsIqJQWg3Hm
Rj16I/PtWh5gllYHi8RtbLhEUHDFSZ/qg+HuW8DLNv9awYgN301TlrgX+4FuqUyINf3x6jCsmLhv
+pSHpQ0Aqh8HtDQjpOmQo+vVbX2+jq0HDvXBK/Qm/k8Z1fDXfNTkolE8dXEWRIrLHT4shOqkPe+x
jsHnLw/C+gf/7Fa/0GVAAs2UA4prcoMFgri4Ki8shzHxu/xyZ69heiVyYe1iNOe/Fq44Q1kXVdro
QRcJWRPviO+0VQeSP9aSSP16M+RwT4wvMm1pIdsXJgI4F8KJzPsPmbk9UL42MrNwUQ8UoMoykfUY
zyOv34+TeMhp2RIqzseX8hlQKEDzv+tBREAjw5L+GtWJjpCcmGRmDiMAf4/O9pue7SFJt4nhHz7I
pU1qBnf/eAsmBKY/It/3zTVSLOhDE6HbREa/5Razoq/FVq8RfNCZ+4QwWcEbWjRWc27d6FCb63Hf
AaFt1s0IuJbsU7kpilQEAQ0CCLG4+VcdwiYy5x7qx/LBd+5FGXU/3D9fahm1T9Dp6gaMBy8yW4H+
Zz093AQPUOvdZzaAhuWxAN+Ilg0SAk36wmOSlkifK+TZbGJWul6Loi8qegOrR6tPwcr6jH0zfMWD
wPCDwQy33cM3PT2t5dGnFQqB3S/JdUyi2ILV5DUE7fk2u7bMjsv1MEHyXEsWGdUPN2s2jVDcbbdL
SYtHTR0LFILDN4iewENPwqgR/lqNfmv1myEbtiMvGcb8/WD7/PpK35Zp9kaoDXQ2USU7HItaG747
sTOVtGNfqs2RvfQZ5crEcKFitZcyDFtkPv6wMwiLMQaaX1giVnedJZ6oVE1QQtvOWwejKOGh4UCQ
SGwOGRojuCwrfkdqTco7usOSxgAUicPB3hf/ETWAHkWedOFzQgzXlj4Imsgtxmog5si4ULw/ZSqH
HwLFQaN+ixY/JVMkcF2SgD+HSyaretNNtuwBvJNVqmbmNZ2yH2Dq10rnTEqILaGdNF7FNVaRvvhS
e8fwXL2L2U1HNGLsrUn2DijDt9OF1BSWAR/VX4b+Kc1T2pAX6I507iy5Pkj1MUki6sh1tUVuEoHX
SK3FU/40ju0eBHAl0LkQbZJ1xJ6lAqGxv+2n2d8v2Fnv0EEZC6lAVh/CEULkVuW/DoqefJwNhl2O
RxjFDVVk4fRl3yPrgEJwnrV46OYSf9uat4BdsYJ95CQYLK17Xvv9M8yNYHB3acBkuDyLrqohtC/u
dFaCc8+JWpDYejRnLZDob9Zah4kUmIwTXmSdVmb99+9410AaeDETWPasbAup6bd6b6+KTGOo2gTR
NVVEBO+iT2xXHQZTgaECF3zu6KgowtIzw+Gv74Ya+YO3gFlFNUPBhD+Q3PnzjV2W/PH/RtE+54T3
B2rkFPXOp0gtw28bcHcW2Lzs3MVdU7m274Ayz+Xt9RaP9xSflUovhlGsTwvl78Jx/FygMv2RnD50
K7wa5W8onPjno1bH/Ee0865VrThzR0Kw5/f8cXH8k2WyRcpwJe6+XGEgZHsm3lGCahKBKp35uMha
eUVyi30MU3Qmvxmv4VFtO5qRsoLy+NnGCl1Gs1Spgyg5SsHrM71joz3gI5caI6KTvP38oQpx763c
JHsCEeYdEdFSiFTKihffZ5ioC2PGhzgOFHe4A4d1IoxoNSXu+DjxjmcLEzLrLbcaCxpJAdkJQYnv
J2tkWqXgFcuoCRNMUBIZF8gkr0hsGd9IEm8Tzx9tSNLAIGV9yZmFzwDRbrh76C9phKPKemau7vow
SPRB3JA0nau0wqt3P809PF1jfY+PdsF41/3QAfqID7R9ju09O9HapTUFhFaQ+BjvpZcpYFrh/8pD
yw8h44+nYzfs6Sx/Nvy+dL90S2Uu35UalGacatH5+KWRs10/NCZeSPYOY40kSYOuuksG7fO5N2dH
jn2e8thr7GJoA8wLJ1s1vT0253gIozUDRqzyrq/iSjaFTWtgmpxnK52A+bexiU8ew5Tue2dwfnID
gEKQD+vbZebufE0uwIZfuM8yw98BanVYnrEjGoptMbRH6BSRK8YyND/pGxdzPluKWXHo3kGb2HpB
V6bJTFJuE8nMLz+HzcfK5FHT8cEzQ31b2vQ/A/eKZQXXWvd7EG2I73KdGUxqHw01AgmolVt7LMao
I5TXOlns9SQBldwcE/5RdBv48dH7RzAArv+2EHpPvkseS8s1yvFlZVih9zWeGs+oduSmzmsnF5cF
Fe2wpmsjYYMTC7fxyePYGCuykxr42oun3vBEANEmpTg40xXbOhRSK+vJq5AypKOBRklvY343bDU0
uhV4mxmdg81RXXeyQHcDowiq43moBlqKWt8OQPEVDu5qMkuFpA41z8uEABRWI3IeQWLrNy1IBten
MeEkAsOVrT32rV9b8Hs82SjXi6RyF7L5B6RarDYVs0WGhOn6F8s48o4WgdLNv7F2hPhdB+lYmYSU
gorQF412K38+epCon3920ZvCUV7RrLYxgLRaKKbvdV8pGK5Kfb58gRG1XcjwyPkp1+2X/DLIWw4n
z3wDd4g7c9Fr72tPEO0jVkWTaR+mAK2iwqyvPpVAADY7x/yn3PqdYkCqny26JUW77Nzug1j6ZN7J
FAlIJHWMwaSb+9o7NCnUdGfF2IVqrj634Y4fKdvMeOd4PZOOqE5L0Qwd6IgXfHeEjCxepq9Ibnb2
Ba/kK32bjy1+S1uoa5Bti6B3RMnXY1iOJVie1g521/cr6oRAWw1VcGv1PN5rLJhrOhuot1Q0uBzh
kgU9El+FMw38WcXH+1vDfABqRietvF35ZpJ4Yi6/ZE3ZukoKR70UlZ/JkINYD5xGTAk85XQVN2HM
NaSVWU4amyqmsKf8g5DoUiV3Eta8GN1IKgZmvzGRmK9GeUKkeZw2e44vjWbRl6bPPdCj6T7gb3wp
bEzDylmsYpFb2TfOuOSFRHIL0VC1EuD4TsNPJ2ZxEpQ6rGxc4HopcUlwn8OFFVX7kssPIy3tsSgp
YRRKi/Wa4DbOuFmbNPZHgy9N+1bwpg9plzMHD07ArOSdKY7YJAG84eoSSLq8Y6i0iP8Uam9pG16g
3M0b3FDrV+y4dSHJm3Oy2P6XQHpqV7v+rSLPTQV76cOcGDRLx0OzmrTH6ctkwX4yjagkyyg2/l2H
miImofzy56fMWegl+q7kmUMPYN/xXbjUAqlXPCPbcYfwwx/uQYLt/MTkPvtdxVzxrLletTAdT6Vl
hx08cJVm9xoi4yq3K90gzDwhrYz4/ZkpAXyuF7PwvF6LwliHAo5F0hFitFdqtnqLXNSkokWIY+7s
PfGmhQU+vYXzoEzbiKR2BliGAAnpBkz4wdUZkTdZMMIxkpdQqQbE9pWw7dc0iJrK3GJqtrDaZDsS
zioaWplEEx2e0MUZu7r7g+SMmjF0wBmeWuNxf3+vGyW1rZEOBMwNlVkNnhC8O1X2crJUuc7fY9iO
lCoTb+Ij0Cgb4XbA16FCuRCvq2T8wusmMQkV95uBWcCFay3Z3xvXrzINIHfSlk+ynk0gVGl4Fmk4
hpiL7XHmyTDqR+VnXm8HsJWfinWqnb1FgpCg6VSsdcksRtvyGA5oi0VskCWTv/CdFydD4nCQ6qsL
jhRJ/fytQ7FmW9AyujE1AWyyiCzwPX0cMn8ZUOW9++LkNUas2JGEGy6elPG6VsuF1VrkPbQidD4T
3x1j6y5gE9KL9OnSrU9U+qK3WUYnfxujMLz9xncN7hFeqa3LpmvoHpPm3Jx1Ck8JKKAE8ssN6zOD
pcAD6MgUnba7h2N+Y7jk1nOeMxfgsHBEOHfkzBtQFUK/fS9yss8nL9VaE+B4Z7ezzFecTq5N3vpj
BotdkdHlYxZXbfFSsIJEUHlauAR8Sq+Bn+pqWjHvzWEW0OlKdZLl2wtY9LemVslUKiekaRksarZp
iF2lrTIvwoWtIlkur1zCNM3kTGro+sb6qHUBO6aIWW5WSSMpCf+GocbyZlM2B3LaS0/eN2z8US2A
zuVeI1IZf6XoVyUmY+35v7ZSBTz8NzHBlajxHHSfZWQUbytvsIrPQD35ZoKCIL/EX5vqUmL06WnC
SzwUiz44/xk7jEpjBEqalwwbJxrnN7xPIWWja4SeE0Sw0QQYVi0ZVr4gfUyP/AWdNm0CDVK71D/j
f+dZobpax1UJbyfu/CvYO+pgi7up/+crfqcqRVWKD0aLvhqNVmY9vdQq+pw+Fjx3iae0Dk1PuIZe
H/dIwos38YjycA4Do9UqbBMxIBR12DuPQMEHC0rEbCehk/7Q2Tmr9Ab868WiCTeubnfdDlNXDOlf
TdNwfqeGtizf2uA3a6T35F9pit0ll2UkgkzKbN+8mQ8gU3kpmwfRjxa0XFAgCQsvEZeUpWjSb6in
UZ68e8Z5cQnnEUOMlZchiZV6SRI7/p079ntkhmYDykhOKUW3W/4ttMLl+JDDhgM8rCiDVVzGxCGO
sehVdXpgT/5wxsBpMoEhvHyrGhv0MGe/GrAtRbbofYaEUs3nzQktf/P66Vze1bV1vV41xgoxn2Da
HS+4KBDFbLQiYA/8w78y7SlLLhZtxY2Pp7bLdOaEn5sdtBF9DnbWmAkNo9IkgEe7y5l9zLvF56g6
kylSwJ3F4MJelQA6fljwm3xVjzePcmfCZhiEuIJcDy7R1RDX/HRPm9GGAqPPwkT8zDh/6gsEKNlh
1BybNtwJUpOXatE5Xlab+QIWI31lyJhEbaUqQZ6qPi/g10MHIjLhJDEWYLUSTEGV+KDMP23pmwwF
xafJ5ziHp3toB/o58dBmYjfR4vqoM0YXfdEI9WG5KPgNb9/ToXNLvlaz8M728ighj48+Xf3vC1Ag
ifbBoSMIak7dB2s+AY/+qSi51upgoFex8QCZa3vr5zRAqb6Gqn9nJpI2+0VfwoXcrXidnsF8LEil
Fzb7OjznJhuH3B2m+UQ1lAYPn1jXiB2mLENKVQknrKD4wxRKAnWyu8ZCd9wHK8g+N7JO6IfFTSiQ
xBwVA8Kyq+/BGhYhpvzGFdKEtVRWsAC31MN+ex/WJKIP0IkfuKsfr7ggQE1hhhCKB/dpVNvXrjMn
bXJpBJgYmWwnTyE6ufrnsA4x5NrEk09z4oukTtzuUNWGb+o6Tuev+GfPphrc+m0fK39fnz/pUPMj
SHJTN81oM6k1sDU7uHM5fSfRZLlSPqPVeRgAO4OdobhBgt0CIiN8X2MeufH7W3udkOWsU566CBp1
J+rh++bJDNP0ZXAP5mHRAL6P5g+yT242vjfn38UC2Z2sIo+lQmqeojzY//T1XwsAE3VnP8v69JuN
wMrdMgUuP+Ev5AseqEOJpdAd4EAXH7WE1wLj3+7+PNqT8dl9qW7mHXOA+l8attzAA6AzTcm4WKqF
PZeBYUSfQOQbeG4Dx8Tvz1gMggSxMTHDd71a+Y+xqQhyDc7afzekzZGhaSbdoFkPHx6VaDkl3bwc
ZSVYQKZY0XMxtK7WVCucez0eWpGgC8R5BWRerggmGVghTg+PUihzccov83bcyVg7GvQzJHyxbUBo
BdkKYZje6HVMttCF9n+py4xgSHExOZ31RlCzTkPMWLm0O1OwUE28kZxvw88mf0uPKoxN3LRosUUF
ufPjxuyHKT4gzCoL/uOtvDTJWLYd2i/aZ50PcRNIKj/mbOwhJBvRGE8QvoSFhY4bC8V000pZ3o+u
4U86482dcV1iZnincePLKmedEp0wVeDzsOr6KQKpWU79lLwBalqQCWLvsS+dXmjnjb0FH4z/Nx7x
FDvCgkjbcwLqgUgmbQSoHOMvbQaUnnQp1r8WZuCTFEPCgMHWczybrOjcDivWd3hjOMkOxRqQydtV
mMa2nKbhkb2/5otZM8Me8PrWUx0Xc3wsphzrpXGt4gPB2+/xrGqsKnd6L3Gq4iKooScRrEEMScfD
6hzrAjXrCnDu+GuWjFP80d3qy6H8UQQq0B334ly9sAWxjyElViuLnXpJPg4SmdmdyfWS34QEVJL4
6nl5zDG28BHQjBeAEzIwbaygMhQE2yoXdmf+vUe1Y4K9eawGKx2ypDM4z6SrjHhTVDz7yC0FmmUZ
igKzZ39s0KlQf0Jmw3kTjctggnT5GAKe69Bg5BUWG8s5EXyRdPX0qibhOac+D3seD2eaiuIjbrI9
KWslVenDxzkBaWwRUSkOfeEjTK77Ve2g/SxNZHAVjcvsOXjWaoOjCLIJsz9EcwWTw/YTqLf4mG+q
mZuUdEr/lj3DNwXpfxp2+opICiQuyofDr4xQt0U5aOGkwYY1BAgoZpH6vJD3zrjVVdXZr6hQstnF
op0ZpMy9nc9Ja7yxD+vWrvDhntaedD9eAVOtLm+O6ojCppJV7MfVHgXPRAGeOiOobigvdJOx+jQF
WFLS28IXHL6v7cMtiTWzxCzzMJsHpC8QZZHf3slB0WxPN3HfpnE7Ovj5Q9Bo6Lp774zpY8uGZ/U4
JNrDv3knQYg+D1Y+v0zvnW2/7l4FPtpBkFdySHumskzF+06ajlh4fVZxU0xTc2QLxSuBqepSPQk5
hArq3UKkMHyd3KsQH4pyTyUk2MZzpdHWTmbqHvs9UMaH2Omgje9R7EuR0Js2ZtCM2Zu/MJYZVWQj
gNWjrV7PW5gLc810u6d6gKnGwBEajlaDgGymJT+QErXhZGPnlCHxcIsNVXDE8vV8KJDCw0jW4CC8
BcuqqNF/jkMv3niiyR7QUtqOO1F1UaXY2E1SjCOsmw0ambcGwl1U/AkUpEA8+L/ZNGwyNuZ6+NAP
jLduDoQLh6HqRXUSk414w1vRLF3fj6AfRnO3xSPiNH28ZHKCxEUHDQ0+YUa1NBDYZUMAh0nL+Ptf
ORWVAQL93MyxHN2haC8j0CALQvoOKONBYArRQtc/TQwiwgEzQQb58Fx7NEINlFUFDCkiZlGuDicK
TVj5lMtwP+ZCmOaHG2SPFCRXQwwx8yB7i1mQA6fLaJdkBgPWu/ty+VQIMQW5IndARFxUAeZydNLf
9E3t5r1VN5HHUWDJtYgnJSndeUJEEJh6eqHmTxQjHwQXb3MRC8zQOPZYo7vYM2jsehe3hzgf9n4Y
Ox50xYqYTuLCI7iiFmsiYBEOKMB8xCAmWTK6xhnKs1ACUQoNeSskoA6qB1psoAUQUzFsX8SMFvWn
D+zNlPEWzX2KK4BAFU4NLQkU/2JWdkojd4pqEecFGMyVeevRWwdo+zOP8rH/EkGafxalj39yJFkr
Yyp9ATIRplRWko2WnE6IlixRLBhb4YVfCq4ZIu6SnIuLvgN+ww3jtnOGF7URlIy4+uGgOME/myqx
6zlEYdxAudLR2uHcBcltz1po+CS/BsR3Ncs/1qfoz6o7yTm3+Lp7CIL/dZV3EvmU12/cbKf7bFVf
690F9aIrovDGGc4CeGYgDADOoqAuLj9T2lcd7jXungwWPIx4HsLMHL+aa3GkA95AyVaI0WRYv4CF
NlSYfa0ZMrJe8wrVVh1wQL/v0czNMwda/SS018RC+Q3/gsdCm5rF0beUU9K/BaWkbaYY0Bg03amo
5Dn6xJnpy9hLxjJuB4PAQqPJDbgIhjqx/RQ8/3nfhjmdoBbDRCnK39dy1WiLLM1g1Osr7DLX4Hv+
qD3aBoplW04SPiZeZ7HGwuWRT8WGbZBN7uiGx33bNfJIKVXugCJYbX9wVyInjP8v3Q245+KyfCJp
U/tsB3gklOC8441ZkrjzK/Z6YnPpU6t24Wm+5TPbZT6WgIXvn4D2/e+WDC6KudO0xoh52RKI8S6R
FZYjFXy32XOue0ncov435NI/n7FEWYlGFJAAD4QWoITMIt4LzGr5MnQ577Q3ZIhqwEONU8hqWRDZ
7pZXIQzNCD+jMnWfpfl2cdpMaG6X9mwSymGKO3kSjCrCaiNKS0RHpSkiXXiOTuVN5FxRWzzTm9RW
4n5Xqp18edsxJ+gzZuXFzqSzPzC5x7G7RG0FE31EwxVsKZ/J1Ybqn179aOe3ls2uT+HkAUNhDGwB
4stroSCki8RactjDbqyrmT6q8KPrj4CB4w+liSM0RlUzWevQBvbMhPfCGn1iEfEmsc6t+u5WswDu
ay6NJURBdRyU0zh/kqWXP4f9zVLF3WbgTVzcVhfgFt3xG0/6vRUZtVNPM6owkPtiAxTXGkSbyC5U
gBn7sKcJy0YivCivoSaTFN5eXH3tgNSKjrE6ZXiRYv2urO5SuROlg5yRwrGxVc68Kq/feI6CUH9l
tmj7lMHilqo1Y8shoQTHyWcXExMZt0CFmcKCXcUEaj/CcVTlpphyWstyEbJtbcOdGkxOd44MyNRK
0kkJUVvdiV1vrUxsAbBRbjbY8AHh7xskhvEZUWyEqtN1+TN5UL+vJsUvZw4AMJihJO7nxdivqkGw
t+x0ZV61HfoD7LeRYqxGt3v1pC92m6KnRjA78Es48S3mfwGCvO2pw4LzmKLwz645bTeSn4KXmMLW
SXy4W0MrKVCEjndRBIp8h6vcb6/Ly1dTo50ONtl4QhwUvjyERncf4HzvfwXHRvQeaXgihiHa0pxn
SAAg8z2A5QszLCHeLQISOerYkAgxvhh5eaBSUZD0xdBUE789FloS30G7ShSosv+/Mld3FZO5G96c
wDxmbYgtNe6UyalgmfFdWtOHKtxsqQJpAWeps8xzh/NAFJ0J8TVuF7L4vnnNlVtgEwl0PDcF7n+N
CjU/R6fCjneoChfL/NziEVFxzZhYBo5bx8kqpv0B39sPOAx27U6nBRY0MvXASBvK+LvIQnRf/9d2
HUohCBnPTsmaX6q3Xavy/Zwqmyn61hxMB/E1sJY6AcZ+v1BJfs9l7V7f+TnT7GJKWrSbO2YDbG11
NFsmo8vRxfI/WAsFXZYw9uIlF7HgBMvSDuX13Q4DFICCDT+SVh3/RL44VIRJdCmD6HnolkFin5YQ
J9MT/N8cRSyIs3SEFm0uV3iTEuxmXw7VZ1bYOLz82CZ5hp79oZHQ2KGAcQbgsbdJ9Oz7Yv4jLO2T
qKvDWFMKj1VpFS7gxHJSICO52v+axbV1vQTUhgY4iCyHU8G6v0FCGMucKZgbQx2d7zvPMdDoQnMR
aR4XOZJzas0kK9MMjOQkPNXyXFu2DYiBKb2T3XMvgVAqQWZrrRztM1/zo8iBJ2h6Axecga11vUFX
goDBSryIo/7C3hb9XqyKfaEMmBvnzpI+jbfN5xuE2IDLt8/PwB2+IcfW75P4cB4rFQ71tjoLmU8Q
LmdPOMPeasfdu9tUmjnQtcuUwcBvWaytZ89F5XcygNVEWkEMfeGPtergAs++L+zQsX9O0gJBzxim
GI9zBU8K7wcHyH5vgCEKWuNAY9Gs3gqLKCVn1F0XBu4gSWEkW3ENHgzZjjhzpoCKNGL9uSbNcWUZ
z3slYsLDXx5zao3FseR5q9qtyAYSP/UPrWyu5NGGgJkS3umA0RNNqD9h9QMANhxMDj98X9O3TXrd
LfNbsoxl9LZwi6rlZ74QHnl3bcwimSYq2+jwTjVqPFpSnRFrChrlh/jLhQptRCGE9Pq2/a4GosKm
nRc0iAGJikhBqg3zEmMSgng2OcLTYnGPSQPx+31suX+RIBXngbm1h119uzaQ43LJ//8j5vs8hFbx
PvUaVVxBqy+ST8OuAwrInv5dT48N4CRHtZIu0GMsM4DKoOZlSwXGjlV3RPJS5N9UUnoOqbvJk8t6
gmYDAIMPi5Y5PF6aMmDPNN+uqeNtgoSZlJCI+H6YI23s/z1KYSVOSedxLq2jVy81WzTx1eBDPCcB
nJ56L6M2gp3C+z92z35odaUA80nIvVIs5xoW4oSaBKt11Muh5RIj2bUFxFTMJMeYrT/g8p39/8yP
9vfOZQoYr0qGOWw9Jxq+M9nWNwerfn7Lh7BEowNWZsa9cSd2nvfUqgzk5bpXFOKZH9xCwutZnEqW
IwMgtGM3djoya0/nPRyjynS6bS4RdMSttCFWiK+aCw5quT0JCS4Ceg5siSpHdEMDTbTT+UZVkqsg
JnU4maGU9RPgQy59F6IpykS3bNmvqM5falv/TLIM90GuY2TVYKRTMWiVGe0jGh0rtyJiMG0GzpP1
p2VYuwf5ugxeHQihaTJH/Q8MOkV9CXwChEUmMXITCyP4EpBBTyeLbQLWM5oHl65JPafXcpO8Zzb7
gKrtr0k7bVGZYtn30nRRGukXLp/t+qgfQoSgkHSZbP3C8mllXQGL0IrtPMOK/PWlVZnJAcFOkqP0
JYvTVrSJZe8SF1GDNKbrp+uqY0GpCF/64knf14tXmvEhcXzDbTjJ7WWRJ/+CBfLGGP08bpE1qcfO
hLQkO1KyBWsR46JEdRv1B/SSOhrM661QEJpxr8LbDOrdoYV5HN65RxyAQb5b29C1o/dTYPrU7JPw
vBZnwBGcmFJ2aJzQ7jSZtZ7Kf99FrdjdaCc7AsO/s9RwSkzA8V5pVtrPYzVl15WX+BaKqT5zCupS
cb7hbibWf5/cvIoozZ3Hzoc2cVjdZjJvag9peNtaL3+9Gok9q0sEi0IHM5MSQe3kl/r/RlwH4dgv
rXaq+aNW6BxcLX/IcwPH8bVClwhzGcUirgjEJ+f9Mb0Qx8w7StBh0ViPu6/+mXEdeHxzk5S+NUQy
I/YY0U3PFXHptHr3BcG+kEDSRhSIrV1aeMd5fYr1GHTtStUEiGSCup1SFj5/XHBzoDT2LM9H7bPS
AtTfOta/dJjYQZ8O4TOw3AmQYq9OJMMymiJHv++2IM9K5TsmPHaVRKbmCSZsVNiI4fFgpnzhl5ju
PeG5ZeB1ANG0Tnzi51gz3+9EiK8AHBFSfIevJqh0rozDW0sruHC56tf15kW8WvKKCZjq8ozGYAE0
FBq1iEae5OMe+MwCrAHGqxIldLmPa6+4aShV685MF6pkvLlfblTNPV5xLtKkFiHBzSvTWfBeCcUU
lURiadqnWGXB72jppwIc4m6BKuGuvp7cIZliQxwQQbebtj60l0QzBZw8S8dXgdLBQ20xjBwQjVUP
aANY7eoCuISViRsBVnCvFqlw5wfukLPsz6FpIQcva1f1qMfam0wQjJ08cTRGd6xeQJkhLtaR1aAl
i/enbnvrrC65rhU5C9bqzEnF2NTllyBONFIPlu3ZNKwS7D/jxWDnpN02gAs4lebZNgUwvBBUUObK
DzcvOA0SHwtHR3nh9AurYVvXmBui3ujN8nSjuWx5zB0PQ5KU3UnbF9VqckrXvnN4//ShgysfaJl5
SM3j3JJ4gZijs61WVVJdXdKrXr7kaZ6Z95urdFjZ6JIVuBoliqubuOfW1KK74fAHaVcnOma3D+mf
EzH5lpDKOePAi449cx8w86smt92n6ZbwgC6WxAkuWxz9cri/bunIC2ca4ejjirRL604pGcSoWAjQ
IgJapL0vmb+X1nLSm4e/AIs+0Yr5Uv43+6vv0VmHYkoYfhYB2j0bTHwKblMaAkpBYaHhukqkDtb+
e8hMH7MNxhEETW9C6IAZHjp8ckpAgSpry2e4hXTntTveagcPFYFBEL5W6ZqXXHPQ7Uk7hkfYZaga
T5VYriul/ymi5w63gsUC8e2Nn/+BXuegQbQAm0IeFHIw1ja9w43mUJNA8bKBiX543bF/jFD92wZc
+CDHDy6xwS0KThg4S6z+YkPeeOLMTwu7oNa8U+Jg5TDK58kK+nLj33lTBTm4bF/8Ss5H3eHoSyq2
VaF6O+JSlDT6HAKT/UpVP505fIxOhiGBFrjwXY1I47rfuSsFbOu4Zdd0yRXZTGhuUapRa63fhGBe
tZez9845BhJq/1I48R8mY1Ys5kANFmasYrt+PfajXNLVxhGpm0v3uiv3AudXkUUiJj+iZCX69FsC
pyvxt2gAVsJWFI3QN8FqBS1C1xA2UJWe1plmz+o0/djXf6wYXJVAFhXLcvZQgBZ4WdnhWZUT4eWN
fWVDNnYEXuoiYkeWzzAYLBrRqK32F84RcttLnuPjwC1jeo/STKdFTzuKV/fP0PZlQ3DXM4myoT2I
nhYTz27x98zl/VlHl5AF5pZYjGkJzjj3ET4NYvNZE4F85vwf+BcNGzXVdx9dNFo4FbP3ckQfO4as
sRYEHJG4hneevoxqmrSiwnoWqAu+9e6YpHfXCbR3d6EBns9Vx/nq6PqZe8hlGTCkVLB6iRD9PvLW
QZ0sEk4t2RABkbXxwYMNuuQmzoK5KG7NA0iY9O1rOHxkZAQtt9N3b8pu2jaSf62WrSG3+Aw41X5Q
Npiw8l46B6sI0Vhj/zLS8woNG7WFjBtUfk9w6TQl6dZsxIiaqSIuX228/cf3+5KkBEPLeRC+F3V1
vFSOKpPxe/dWK/MRYgueolMMvz2h/OdFnV/6x5DfYjIfiUDmQN3I0T9XDzkkBABHy8lBZjpaDtKK
r5GkSYJ70RWL1spWo5AVUt1Jb9vCdZVSQKKWPywzuZqf6G6X5ohu4S0tkdqursmVAHrl0D0rPVim
X6ENtHdbSYy10FL8PiS3MRyJgGhFDR0b5qWBWMpaKrHBxuC9cMN1Xvueui2hbe83HFG6uPD51ARz
/FPZhFuIC1F2U6TdHyuEByW51sXC0osn/0dTvtFjcXZix/9ML8NVkEFaxWkH+ebnQBaxcjcnAu8T
yuvxARCi0p0gjC3RmhuUOxH13LSlnwF6nEyB+WPiMJ34tPJAqwk7g6Bt67mrzF9vRvxsif4m9Zju
T1PC+HeYC7d1ON2SPYEmdUPJer//U4aPN1MM8Plh9vy8Y+RuHHiqmxdSySuPRHMAaIDHv2hpdtJZ
01tdHEZBvd3V8KOxiPB4eOxd1HSxj0dbrnnUHsNSjgfkgIE7vrafdKMKHIutB+YqAbJFnYl3RxIF
feG3Rm+bXHqJxIOK4Z5QH7BprIBv2u5DtK6xfsQIZfCz+Wi07Eb4k/uTF+FBuQzz+luO0lHINEtz
qgyQO5W9yLxebcvkSSguveOwB5pjolK3M0rJIOtuff6FTfuGXLeJkSNQizHZvSvnsY2eMNk3xg6s
uSbYmhaa4nxxXgkd/zxXBuNw0r1EG9qCIQBBnCMj4aXDk+UiVoXGAwRTD74V2AUpzvh9E+bM2oKa
2zXccKIwEOZRqTUFFAnAau/BssxX0StZJ0RpdPhllhpQALtw5Az5v1+dsife2BW/8J2DW3cPPwFu
7JOnpF2cJwasOpVC3ZUTDnC/9LadiGClIfxUbO8x6TSPlWrS/xXKhPpFwfhauoQpHkVgdi7rpcLC
TbJ5et7MCsekxMg2v+RKxTSddG/4hZlrDwWd9fGHzxKZfLuMEmFgu965msj1vxtzLqrqDVS8lhcl
gslrF2p15GP865qMjsjeyOlPaNZ1Pq5T7qEA9hb092Oj9bTAkrk/S/6n6ph3zRqTCU8yUoHM8SPV
zeLSQe0iqomeMuppmSM3BapVhAWKevHuzc8O71c6tcNYfr/GBLCNSgz9EYaWZMYywGGE7P6cg4ae
lYHrJzToX2+DIbS1UMzDCnv6lovcCYWLQ8Fql9sgyNeR2tcWi719pZfWpz90uZt6sPg2kIn/XuLj
B4HhC693U8HIU/yn3hiIvLlPGVISs03RXRuhLC4NIu7sBtG0L3h2IRa66i0ObzNPEDo2jQGZabmh
qjF8V5pwm7ulc4wIc+qA6RYB/IbIL3aHYPzi5BEZg6ed5SwRKf5QSmEBHcR5pB1xtz8ZKKtUmLFi
ug/pd5AEtZJVvuX1kB2FJSwgKhoGgcouEcWB37N4F3zuLibROO4WV+0MqIHVWol2jYHt+urmSgC+
uTCTa3JjPxVIY4H35dNok8DuALgY0UQ973NYSa7faIs9kk+kFpp7RQc+Ua2PJyXpW4BF1nAi6M5b
MZpOjOTRu20US29TtYx3wg7WkiVfySmEl5ttpIXL+V3jhf5aO+oTS2Tu21TgohaotzxhSyLWTpW7
yOLYNV6YbHcrSAfbPUfa7XRQmXKO4hNtIFrVMvVZZZa31b2NvJft3m7uv+yd5uvtKCm/VjEJ7TtK
sKZ83/9/VNma7G3UnlZS9QIQwtUwY4q3UMd9ODXwYLxx64W9KmwMsNv8SIdPcCX+o1fpP5BvLGlw
vO6hrqD42SP2XRQ/wXtrEjefjPzN/mW4Q/FhWWw5UEsU+QK7lZ2NhVkKPOtuIhMuU80FF5+HUMFJ
Bxea9qZYymMoloiLIDB6R7HseIjp2ix2t19VmH6I0o5o93rt3T53t8x084ycocJUf3Z6T065PK8d
Fa5T99IjtTx/wUGjHhmU+vhXMtT0QcGdjhlbCloN8+b9yc3KThBFRY1OxPHzGlRAsvzDbOj2Gee2
JITLZK8Nsv66bIiBCwPTzHb/DYHynszBr86bvPgY653OzEjzSd3anKVzU1hyFnE0FxCvXJ+jdDNe
ym6JZXXQS1AvxVxfFNWfPuPy9/wX2bkILpl84KGW6JsiEWk4Wf31bJjRveNc3s7tcbkq0/XHcsd2
ELeI2GnJfd3XSmyNF/uTqgOTc43C3T+Foj06NjrJJ/St9qEjsF6QFh0d8yCCOQjwdbg/f4mGv26x
zK+/IEBjp020AR5PQRKjGSkAbFA44gqj00TPYK/6m1vS+fWbTMngEpVAhvtuM6TTInxAIe5zgQb1
mYHW4of+Yh+xBsGzRNVFdjBn74q+TqXucRKInLcC3Wz+cdkh26eixFcgV7azyqwkUTNhzWP6at52
GFLCklc86d74f2aglgcrSAMySu2COCslxorDzrINXBh3/1TcniGAVINs8B6JOF0UHPglNftVcreC
fgtW1xgRoaYray0BmqXc6Yb+pwKHhfxFHPMp5wld3TGtcIgNzGHkWBYPj7cYb/q6RjjHZshJcIW/
A+dFL91Uip0lq7zv5FJj4WFIbwiHYLJWtokyVi1FLQfg+NTE7JV3f0pq9/JRlU/f04L9AXT7PU1K
G6Te+zyqpnbpRMFqPs4wtJK6/CPa0LG0iDYWoF/NlFQDxEuRrFiENYwJ/pdWOrtZBVrSRsAKVj7f
QrYe+ml/caK1ejI7VOtL4RUfcNp754fRKYV0FzS31jM3N/sfzsfgM/j8nx3MyiLkcMeBAjlL5KmO
sTN5ZRd5ttuYsm7qqoN561jfMk8DUzDrNtePpREeYt4T3FteoGENTR16GBsd/tcovAus/iBQtW23
MKUIvWdguyHcAO7JCrllaH3KnjjUN4Hkuv8f+wgZAguuYAiGYP708iyK24FpXG6T903R7i4+pxhB
UpEXScN4+qIsLPUS4qfLTDXNtm48gfFlvZNJiouWU4zZx/D52y/hJrdlSbeIMMCCn48C+JfonhLo
GUEuPfcLWeGaz6tnueZK7GllLPxf6xG22079/I6QD8ovCM/c41oGHDj4YIRXa/04ToU745Z5+/sa
oOLUdAJ8jyT782V2+cRj0saPQ3J2v7qiVBtUpDHKtpjdldT+Z6QDEYiIze9gSJR1ONW1UVjZ11Wd
1i117pLj3MY+fOB7E2N7ApNR0S9huWCtFyzTWxazz9bJLxKfT947N3vqVlbI1sTv/tuyg5chKXVc
0VVdhSjBj0AxsHL7mAL0clIs3ZTBSoEUP6Zk72GOY26knLMT4MBYV5VK/Yw4+Ni6gU5w9x5cj2Em
nSZXFDqojG0/5RN2CIkHO7FBpRxDXGsCYU+uo1J3Sz3DBIghxCxCgandoUckjZldiVamjZpNIe0V
wH+REYlCXTAFPHyvSFip867oq8ysGZCbgk1fsOxJP1PmAd0C6hFh+3HWHyiiH9WIu3x0YfFG4ekq
4JOYdSQqgwmtc/uXFrEdG+PHRnEGgY8awFDOCmvLKUePJsADpl1NOHkiY4AJ11kdPscr6tIZyAm1
AIQO3RAQfPfPscWMqDK4UF2GAdejvaNPO19rcuoBa1xi5Lqjx79XNLLV3F/Gc7uFrrtZjSBhaUDJ
AkPVwXm7xxwV+iIRsRZGmZE26snDP6rwU52tuj81AT+HGmy9E0ont+H9J12Jc+DbYJKQVmejD0y8
CpWOLNDqHOTKLPdeZhb8wSET/XZslj2RpWaXVC6PpiQYJ0UgAC1zTw21odPp/RcUUWKRWqMnxugJ
IHNwOPojfRF2sURICN5UQtfAa9Nke3ENDsmdyZaKOGrRljhhS/91MMmARRt1FMBv4PM4Zrt3OabX
BcJani1QjTAa+OYnzcRbTLePzDeoaVUbIBQKQZE/GE989EERfL7N8FehTWm5vSB1KVHEqNefsNaJ
gKub6Vy56F8KtZxOvxzF2DmhuI6TD8axWV4mWmcp89BzLC3bwZDcGycWYoOvVqGwX4Dys9I/oYd7
KYE8ffPF6pkEpQaSgB4t+4JhsJ4jCTUL8TMah2WKDJUu6JHUVPqPGaJdrLBJBqyv2yuiTgs/3kCL
3gzr39EBwHjKNSRsA7XxjfIpT7I4E1tlbcxth2t+rboUye5ZAeli3mcoPUwpdATE6I8zIY67Kexs
7x9A7urWCJv7ry3ULRj6byAXW7S0pYQozdq4Eb5MOF37CN7TJgEjSppNioXdOB3u/3GP5gJkJsG+
3Sd+PimFbbf5jch/bCKB+5A2R3d3RKITvFgMljsn5NdwvKtBIPlon/C9Yh/VuLCVlHdyNv72+WOD
05+vGhE896cyXLE9HXfcEU6fbuo5LCzghm5XYzQ1b/Kt5gTOuJQyafzp5cqLx6h4DshZs7hkPzVw
bbqsyjmZrFE/pyDybJ3FQ3ZlxhwCjpQXaESBZ/s0Ay29gDotZiPtuVLLYsnav2DJm4iRla0KLck8
dV1r0UwqjAZdpqHiZKY9fL8YVq3hlAwTg+OeqG85rUhm9bTzif9vG2EY5+U8WdPslU9D7UKxysG3
ZwhBC3son2x4i8INQo+qwjwjrHr8cTlvaUYsbc/J5c6kOZSZdyGpY8l8QOBn8BZ8522sG96gYO2H
B6IGf2tJbvx/8Kto0Cvl4yuuhBdGk2h1N/feK4Iykq1Vs9O6GSuiRtkhQjMYdsOIu2Iu1higUmB4
2ogyBVTi1aLji2r3U5LDtctwpYlVDFIiXEtj7LKfmYphGs5tTrsT1jY4PZywAX1vPhAAGHaEupNg
fiiaju9CwLBz1kDQnNYeq0Rglt2sKM3+NGZl6s/REpm0w2RSBJV29RsfjwUd+EIu7gQc3Jy0BHZS
Wi2oHdXeKDG5BzGy98nhnEbuQRwgQCeEqYstS2QVRpZwtG4svmeduaODCrIGrDMZZa4xp4avySXq
V/I0b83mnrwRNapCbOLF3h29ERGK90nw5RTdCpH9Qp+FlTqdHeZTVahF/9Cm10HkQWzDX+Jv6cTP
EFJjbQPfzUSChFK1TTcc/mnuUMhtu0rp19JBIU+unW3BNmqFO9CKSQ+06Lby0DihowCe8NuTUGWY
PDHpjUpS2JNjt9QxB5HX4BtJshmK/ga9TCzyCrJtsLgtAa3ksGIv55AyJLblpQRb/fzlDTXP/iNJ
LmK4SqC41z144GYixALZDB+YKxYeHCDhnjB1m96zwdUd2ooWjRj7jmHJ6c1sIhpIlG7OxMgRe3en
yAE3t7bB/dhV2nADgbYGqK6GLG/iJcZ4wKOR27jmmMvUvG8QQvoplJ3YTRhtkhlaWDmsJhCo+uwI
xtOcOU8ITMYHizmihbUscxgPBuWxBYfRRHEVlLDLfNFi0kWu5WCvRthtHgWgAWHd6E64HRMt3SOs
9NB2fKCPnOjAHIdFuJdM3B7SxSbqCc9hAIafNPFkv5K6WreN2uTN4uiDPLskj3EHPeTa8ro+3Z2e
7twdMWuhYdGdJu86i3kY2ZYJvsm1RSgsIiLM1NfjKbkra9nbePHdYP4d/CUlolFYYZGOXirleDGO
md35l01j/qsCnQpSeB/rwJ7ThFnF2RBkVT919mQDnh+7/jE5izZuXALHPMX5DomJ6K+MwIT1JcA1
Ms/QX2whuesnMWL/IVcaHo+LxVoGh+i5SRgSgLs65B7IeKs/nbgSORJgJj3BGGo6Ge8He25VPhaI
/dZNzdYiHqZV7WT5ZjOeDDMrlbYNQkTiBVpYFP1ijQsW6fHetRo8sRktCIA9zfYQ+Gmt2oMSIg4W
PYNOi6RKyxWe82vA8UsnVLpcTEcEogouiDy3IHwDB7n11SnW0wWrD+s2jXrIKXe0EzoScJ/cTfLC
sukE3YgImz8R9miGL884U+xyZrk4sYPMempWg7iz5UT1vNuctafs7OynESkykVmia9XBpDTS9yu0
ibQtpagioe3cE5sc/KBHyCPex/MoaMfN/tCL0qDy7GP8HjYCWHX1G1uzsnhH67WURaTnPd6+SZj1
o7066UP0KgV36wH4B18XtRceFjbaxZyrOz8C+v51SVJoBDs9MrlD3SGGIzjdL8cO4ANp+c65La6r
l8e2lkE7J0VQMTMDRdPJoI5SWqQs3/e0nogpu7nuGsClvJLsmjnJSZdNs/LJjRLioSihKvkjgYkm
wSed2UiX6Q7XDpXc0NmgJjkhRb5gleWhZUAw75OWs36A34CwsfDU5tFGQJVlhLbORfUrEtO12b4O
mP6tNq+AlqC0BrQ88sYLlSQ6SUF/sOfvc6+fcV/smRR9V2K8nSoVtJUZp9EHvf/XSBJcoe4sosGV
gejFP3gfwcz1O7YkWYRoKRkcMCqDR/LYl0Q+aO22tNMXtucbqUmpKBwm3L/Q2QUFboAwD16W0MSH
dr1ZxI+4SMW4xqnnKsZepmiSFiTQfNTpD9OI1NRMSfkjLcmQ8c7gV+8XD++r39zIA/Wok/sKRmyY
ASeQ03PNjW/Dt3ggurN1Sfer5C0ax4EsUnAJJPjpqkycHx/CHFKnqjEXKBjaKhfoR4Hoj0P/9+Z5
isj3ZF6fi0JP5Aks496GVtqUP2Ixu2u4j8l7wY3XDGVAv/ZL7cDAGi25Lb0Gzc+/qds7LwZRY4kI
bQgJCG97DSJp9+7zc6L0CYe3Yu8MlK71b2vhZTtMV7pdMFxvsKyBzfozda22rj7Pvxgful7HfPmY
42rlIJmp+oWKCZ1ARAn0+oC5wZbRXd1oK+0dZMHOJ6QiRL7iHkhdzJ65T9itrUZRyPSTN3rds3z/
3SiNPMWTEA8yvG5Xi01Pr9DPdH/3LX1BYz9b1cXgzn/3kobVHyFhQKqWlHdYplKj42fWLSO9ORmn
4Xe2JUCginX8OqRXJn8tsxpUQm+L6pY1+9zu4RPIkMHiASSElQoOpr5SlgpJ7/8Aahms/E/V1LBG
cb9J5Zb/dJrtZaHgWkk/J7YblqlFxHQrD8T6ff/Uc8eHitZQ+cugvH/h3ekA/pTw2sYuPL3fkBUj
qkyU/AqSP5M6/jFIesETAD6ljFFFCblg72jFr2k4ttyNxQuaVrKv6Of7BJjhyUeQhv7A05IxW9s0
+1RivtCtSBpvwTmnDyMmvy+J12q+WwamsQQa5LkqLb23td3Fh38qWKl7qHGl0AVMSEwtIbggUkr8
jIQprJNw0axg+zLVoPAdLFptU+16kLvbL+RvARCwYyBMWYF0/79FQSwbkFdivSfVdyz5gWGsqAvK
HeRuNo7gYpJVZAjrgsVDNkABjxe3KZF9x3BnYbyLbpbd2x8D2UFYmqfBjFDvv6PhEjVNS5VlEvld
Hu7vP0g2laPSi3fWGTZqZPaQiSH+cZfVYWzZXFfNSvY2WirrCcXywXiUXzuxXzVDp655OAmDUT5Z
tS9LtJrStpYqtIMufxSmJ2YsQzg8ScgMhHEImfnbKZZNyY56pSLNJ69dIRtjZJpPAyRacmj5Ka7o
2MbpyhLigQZN5EzzUunefmVjim6wNF8oGyLSZu2iFWdDBexCYAMRdy1vqJMrMIBV+dbrUNQK7u0O
WWcm/nLkm+qGDu9VXlHbcq9ocOAI5HCL6C6L7Kq6sfAx+dFaWlUZ5LuQHzzmunP4RrjmEtppO92i
iQcRbOkj5YaLDM7UZjZ0BHDmoWyE6wYTH2TA54qUS7KbzbQLVIXcdB/dYvmg2vecv2zuzUsxvtSS
uVciCbmg6rphBHm403lmaPFMPdyY6XDBPcRqZjHCMGGSM5Go1XaSrQC59rZisXcJrz5in0n9+auw
+Q6S81y+0TjeuP+dauUMbzLTqMLjQ9jiFos0ttvQYEv+YTSWgtxvgoKivQCoY29O/47jIPw0Wtpb
dkac5d/MU0p74GBY5hzW8P05xg/+xLm+jvuB1sXa7aFzWdxGF6CtWab5LPgjP7Or7cS3NMbEYNtE
oxlEe0s81z7yoJeGpba1OPW+eFi8FevJy6ZyxqaIIhee3ilxL+cSSOvMJeGjail4N1r9hyVMGfai
H/UETd5jCLfTS590XE6DcEto3H54si+P6Qi6ii7EcYFK0Im/LunBjv1AIxSWEaRtiH/oAEe+ox4L
FkcGfWq+3mMar6/8fpcAMdUJPR1/Of+ezl312XtYe8zUPGHzB64acQ7wyHzdAHbUqQFEAB0nnQNw
/mtz88TOyNwc+R+ItaOKJubtVKvdmdtec8hAtV00rKrmrmRRUwVqZp3z84CN5h53RqtbWpXH3ULU
2na2/bpnw+rkJ87X05KVJOx0mC+zPfXpgvDPaDbfJNxZ5Y8ZyLokaY6fVDd2aqGFVeF8z5miUgmm
6h8t6dGxWn+vn+cKvVbBVlOq7oD93HWIr01Qzjfr/dWCKXFKllSHuhMwpnzycHVRK305QHnZUnUY
/feW28cTM6bg5OsiioGDi9AnKFCcQiI5ECQYvI86eaDSUmbR2d45tR1zcIKWw/xBZk7IIBbiLNCX
7RM33TDpDc5SZAWhtsJXpBtt82GnnUvJVitCH26FojPXKBYcDb9pe9XpFxhmGlx9IZL38R6j/wJx
4g+JE53HcVFfY7bmj91uup9+VVWjpZBxqbGXWfTFxlodVgKxYGxgXb8KrfBQldrqiO2UzeqPXxw5
RpZUUULag1WmOZ7yd9Ko7xjGxLJZ3LcF4ReozKeHWi037HOmrzqaQLne+xuwYexD41EVI/T1C3KC
nRws5rOzD/B6op9jaaif+eV/jAB64piZ22KKFEOa8AV6vQMXAjkOo+cE6yzmbS+deXhXzyRaUZ+c
IfM0Kt3nqn3R7YXYg7waL1gUpxbY+FddUBXJit+NRD0P7CQ41PM1BHlr1BNuR2C0oktCt/Hks/OR
h/TmYq8GfQNlZoFba8LPb1pKy2iI0e9qm4QgJ2XmP1CuElwbKwT25wcg+PlGFE9BPqWieS24dK1s
ac7wDp7tS3UtVc7SAcG8xyiioF98PXxgtHuyQi+7FrEoeptBZCGlxQm8pT3/YX79KTP2MI3w7gG2
ht/2emB8hxdmVipZDFC6Gfit4GtmptuWfB8ohhT44F0Jf2TOwCFIERTwaaYasV1+hGUBSQWiBI03
aumfH1Vq7JdOiwtPgvp3v7y0+nl8OHl4aQY3NfVlKLoRVUZ3f4W7mG2Njpn74kCt+FbP1sP3rhQY
gUy6vZFot4mUt2yyx5BVpgsnK5V951mtECK5EBwe5IXx4Ns4sL6OXQteqjcgIj1laoMsqYuBen+t
P4lP3k80WG94jPJ4d2cLSxtA+PpmI45EZD0NHvgg7Ye6QvRbW1QaPjUOSq3/YbkdjFvDILEy7paB
2Gy9d1cVyCzj9MJTEmsDxJA4iiUNnSwjtMQIbo9PRhRasiWUA67IrkuJJHZDwYpXgEkZDpG5Aqnz
vfMyz53PORE5S4UPcJmaGdrES1IyjBM18B9LNTMcTp5fsI3jDXHlqrQ+SBdNYE2pk+3xpiT+A+4D
TEg1vO6LvHVtqD4RCrz1NX/BQUkT+98TubuNNio4w2QJijxtZzY0YdFISsM6ouJ57jk5qY2Yr44J
TkHb6OyRGehHBJFoJE/uGRzHe7SgJmdD/uPq9QMZCJWsjwaykq/XkqKwbfwt2sQPCnbQZN1vrJ/T
XPUKEIbYXWNrME8v7+Tq93cVIJZFZr3BgA56TrRL8E7/rjuhshshRgXdkamdtYe6ksUff2TE3msq
gW/Jf23uUrzli12mFwMte59kRCzPjARj7c3ZzGSeD23bC6eQhxSS+SRToCqY3mIpBv0TJpEMch3F
sjlkKNb3b70RzgPpJgtFAJx9RzChcjGENkPwVyoGRozx2sq597QDW+CggfJbpzNeLVQLSpjJoXwf
SXwxJAzeoEKB1dqHKetICxbnxzbIFPoukG+Iejfno6KY0dLS4h/luBEoAlucCWgzYUcvu/KYoUQ8
L6SK+L9F4rKSY5a9WYEAeTm7sNdBRXYhkGcLNlT0tU8hV2KMHJNhbfwK6Up1y+9v+hj7Vb3Oo/BD
7IoaxwZh6RG+IGHKDCAdMQpiQwudZEUP1h+zX8M2PfUXg1b/L+G3dCSS5+a0qDvH4CGP2Dt33MMK
q5FcxolTj8qJeL6UjhnWKMCbhdFbKT4wStX0VQhimlCTpSD0fugfL50xwnIY/GwU++4AJZYaammY
OK8bpVWzXh2mtWvUCps4xuqyJ+0tBp1pKWHesGi17WycCfUumkX6sHSQ2N3DIxojJTxubaHVMh6D
FFBt4NFVG8DoVl73aC6kbRFlUkIrDmzgX1z8u+5SvXTOB8lTtApPMLidXWF54LYz2PD25jcnPY17
G+zK870y8WwP8u+f9xFLUeGBk+ZOLE6SEi3uOjojkmdmi4cSLbrVDuiDIqS2DRH3va3KzDVtiWxt
aBIh3Z5LZ4d/2FPJ05nYNzOsP29xJVBFO5tw1v1PgpBm7em9GDK706mF49I0DcuLdGzrr2RLX55P
i8hlgLCWAWX5CwOXSZxJdE62+K69+nFG9yD2RrnfoTdy1Tni0T3FIlkjmG6WXbKb3ONLlFkmh+hB
SBnWmqC7IVanMFNnx/y7fKn9F++HRlyoqDmCV+m4hslcHZA5R2H8HJ3TkQYD+Pgq+qg8uEq8if0z
QBw7EZf5M4G2qKAyIDa0aVYKpiO66YLUt5VuB0IaFm1ar252psHuTf6mqJwxxqIzn9eK/8BgEzWJ
M22/2fYtMljEy6ip+bLxvnbZGc0uht4c7BcLn4qLKivTqB70DmKksir5KW8VlPVfb0aVvU1NEuNv
bZeTp67RP0aT/sNOg1gFm46RRW1HkbPvJey5YbnqU0emvSBbM55kdrnAalT1ZPhlDEoxnLp4+u9I
QNYbreFaz3q5mAlvl+EfncSoGa6Go/XizIYcgzM/Wz20FGxZYhwRVvHiRXHYxp+cmKL+NsVwzV3p
cDa0ddcinO/9v9omWg2n50iRldBQhG7YswzWukYGCoJGzxVuTVBUVohx6HIHcZLe4l435v7g8z+9
SHnKxqmfjCoDHBrn0WFfzl2LDmzWNcuDrrAHEgsVsFilIPX1m3fPFY+22QlBGn7/Q2NYmh22As9m
4gZgABF5XrswzUT8GUw+KQ1aLZTa7sEygSIZ7WnhTHYFeK7HYTcKj1qUvOxnLNYoOsUTa7NeF4QJ
TIIC8MvI29IoaWCiSTJ0Tq/diO4roERZ4yXB6W0qHN0JzeVVe6rVmpifda+i7C4YseIQtQzc1vJl
WPGd0WwuHColzo9QRS8NZ1r8KXv3sXC/9BNJH8nOsd+8OgW8tFz4Gb4Pv97zTplJt/dyHuabRYpH
swL/1smFCphn0r0kQiPWe9pmqIcNZrjOXxu2OwlECgGXLqxmj23xOFYKD2pa52pKD/oU2C7Cke2B
xDCi1Z8bzg31lG5mQJxXlrLqtTI7ZdWIeIFPJ6liUl/ETMO2A/mXJZ8UxsS9MNPJHK7KSpObCoqw
XyTdV3aV437xyHcwF1KU6Z0jlJCq+4NtjCHZfkhX/lSR/WKuTPSQERd9E6FyUobHejruUkvyzfiT
kXgcmAef5PDVZ6NgNQwENj6oby+drmDTbc5zvbncq8jNgXLsr1fbpLw3Rt4IfgTt+3Js9tdKlSuk
0YCgwCju/ZLLny23QnAPJDsPqCj4YZpFHyYPJkZV3Ti3xeNdedzEHUsOTGSH4QTJNigMq9Xc+HkS
lo9mUoHDTA27qok82dbwEAvSHEvNwVJq6U05hjwsJ8iMw+kVjmt7wFesmmEveZ1yNAoSbIevJNNW
zlnvB0NXCXlKSk2GZ1AnmLU0/GehC4hMeILPPn8Wzho9KkmNDA3adhXrMBbeq1qCvC4fX9Td1x9G
LiO5Kus5L6DQ9wBiNe2rsqjBBVO55+t/3FuU5hi2wZCH/isCp9loVplwFc0FdxcGZ1L1xHd8nQU+
STI7Oq+VXhJUZhGldQ9xDWugTMCCF3hZINEy1fCctHc01eg6NKnSkCoylb2lpf58zMBKpM6ixsi3
xLHOdzKKNNuM+Kivk4ivfOm3YY6zthO2TdxKX82aOiISr30ZU4Q8lGP60Fb8YNqkB4Q7Gxh63aJx
/afc9aOD79zmSAK5YWS9BOiGAC3uOHjtIJZbh73/lO158dSzJMMCK6Oaoh1UvA/xFf+VPHsA6zg3
apHu/vgf0vKy1nTHgzNRFV53sUVmUkAKP1zwZ8FKCSwqrGcg+zdeg5iBopXI39UHSbAC7ZR/dYpd
eMrzJY67fXsAtxMZ3f9gvQUKQVOFDh40/ecMY8zVmtJpDlkbZl2H8dli+S65RHGqCMGTCNgYUhaZ
h+wL5tQ6Ua13BDq7xIsvSm7glGhV99jw/78s0+nIDnAZXI85EZ4PODpoBGVNc+rfYFGEoboLKFGY
I/vhEGJFX3Z8MXe7YSPDK//7C3fZdDwztGvBVVljw5Kw1Yh0F3BqPlX+HbEs0oYfmyFxOGq4bN5S
o1LB+/qzKNi8HLBOada4n9Q4WQu+bX57zYQuuOJPyQ2ndd0mFqrj08aW6xDAkHiGRdIUKap8IaBB
I6vlOiiP+2vR6ZCyadEMo6wBjb8c55GXPCxmH+ASK0Jg6AQQ90Pl5BYL1p66iU973ySSl964qA8n
vULSlnl/rRvbQ+vJNBNMq1v8fshLmBilVZX8FC+FxuGNoMKOPN7/+M0IDuENiVKQBMyyzd1WsuyR
RWhUeCMT4mKu7yc7UtylA5OOme1JLaDHL3aolPLGs0CB6z396MGTx+xzt3RyW549wUvbo2JAmLEX
PvIBSSaDfCDykHxM5bS6KVeX+2lcUOX/0FvYMrhyAI9m84godckfBtn0xa/jkV/t9HZ9kGAPRnQA
710r7mx+y52rMFeEA++/hLPqkz6IpGRQMcNhCFzrpGUAQdUXDypUWKsud0qKf/loRJKAQvMm+Wom
MjLRCjLxZKyvp/CXUOLH19EH2P/D7BsbvZDKPuOGBV5g51mVz348zTXYlD+e8yP16VP9dFnAVQmu
dqJR+kGLkINTekA6ajr/H6IuIHijQibtXuxeyoNcunvDXHMCYOSKtn7KW5SH9hDTJdy9NcuFKcTo
WtCJsq5JDDSjAHaSa0d7fNnIciA4I3fCwiUeIM3lsyIc35/HhYWNApeTBR9KBhORuCdrzfRAcm9d
qXBitkEh4BzVGZY3qQlLIJADs6+eAexe6aXyFXO0hzMMnGUL6pdzXoQsXIikUfEObgUO0tImDQ5O
6xi6tftoENHC40Gzu5q+ipaiub+Rtau+tQOnuCmGsHODFn1aPQ7h/hiE8jjuWWzgKl4KU81400wJ
dTE9hDB0uUrOgGiEwKQbwoAYlGXvmeTTWxXSC7wxPqwS1Pa5JVe4zNiQhVNUfhF015e2N+GMaTez
NAt95QozU5G5UB26al1Ldv867RuHAME+9ZLFiNmTqtbTVTxj8yliZvzTRDq6f4NkhvG8U9ACUC0A
nQwbZl9dFQRNvYHUGKeSNrqCa+tkJimjiJgKRUFvsPIHxPev6EXrH8vkd/1pP6e2pNGfxXsLrzZM
XAkJqsMvicTUnO1KoG+hM2OxuRsvjBl8xBpXOAp/jsiRBKkysCosevF64L2FDIzf9t4/e5rCvgPe
KvOb/9/HFN1HWS4w/WJWzwFG6ce4pa1LI497sv0eMZeolYIeAZC+qIQxEvLG5fFPAQLX6ZinThIT
1i579PHMBpFTjQGQv1WFKyhcvobTF+uaC4/gFHrG1Wyac8DKbRxt1D64DEG3qhnhwEnx47GuU7QF
/LuVLZvzHU4Uz+CIgN4QQETHX3BMPlLheMrjlHRYAx2IKpqvJ0PXVHM/XmV6QzoqNQMczBwSR7s7
ZI+04OeK61OMZlT5uWOPz8yLTe4b5AsjPrpHSHMLm5rTkXPTMK/Tut6gWB1IX/68AyP2z3E/bHZR
oLknkVcjZUGLWzOUshuDIUX6cJdFs9oJ2cz6gTrh4DuwkVttp5CVb7T6ye7J9JTQFCQa8j2h4cPB
1nrYnJFdEIseOAbMgAyhXJg++STQWhKI8ohVl8mNMnpzcbjJMicoFmVqtlb6XGD7K9bkfHDqovbE
QmavqwRZEyuq0gXUC4f3mSiHrR5kI6k3yraCEPsWxGBODy86WDDuwRQ7VFupOUH1lbJ/crzCe0IG
iICf3ADZY4Brse46lk1e3iU56MvZR3QB9UQD4UIisHAb8Sl9e9NgZVugD54xF2Pb9M6hePmrZ5IQ
RAj3jPcl1uIR7VAcVPBSSxfisFOv36+hQtrQmgy6K3vC/jpwEvUxEnm4VUr0EToqfA62jGolHLw5
Z/X3na8VJHtczLjaAR9bX5g6Wk1gDoXS/vxpYgNFltgXPbujrn8A9ODviLhwcKpLaNF2tcJHbQbH
pC5SYT0FZnSSuUZRC+iXs6RKLXN3wxN1zglxhS2Ss3sKBS7692anazgRCu05TYrPCKKqx574BfWj
5ix3oV/kZLuH0EnN40gQ7KgsUpjzIi+2urGn9iSOIlph3rzkO7pjEqUPWZVZd4ifekTqcocplJd9
oX9VKNNh1orAM3de5M2j1LBpCQGWeJkNCOUCMtrZKlX3SoxgzL/r+WrFj5ub66UExIs/4dVMZyYh
v+WvzeT/m9CjCnebdyIOsNbn9XdA7CKcwsl4y0/9HsOP8VBF/dsmZaP9XqaBkSRd7+QftBAmdqsv
AlMHzZrHx/LZ/FAxnOYf/oIpHQgbufx5h9nWFzBzQsitOjMiuGmewwcnL5tMSE8V5tmU6TaB46ND
WqnkS1gPAEjZXtAS0TOKLMMaEADo/a7qM7Bq+A0ECM/CCFApJ+VkCCmHqA5PgZtlP0u3TbLJ0/Xn
3LJ2s8eyeugggcskpyUC9oNGJ0+MWSX4k3qlYktpPahLMXZtpbV981CYAOiBJdSiRvf61zFJF9dp
VceiyjuGmZuKq00PXrmSGFXuqRMbgR8ZsJYJ108oF51gAh+eYnXT12kn5uuIugdN0xUXUn5CPR7X
rZU/k1bCA1Wr8J3tcyIE2gJKHl37Tieg15Qc/VYnAVQHqdxFiiLE53V55Bwfzua/dulr6ECVpqzE
EmH7oJVfjhTrHB6/Aq0byqdKQqrZKruw117hp0ukdtSPBdoqZSw8oOD2SJA322eROKN/Fd/4ri+7
zdMM5RTzX3mcxOePVr+0qFVCTTxYNFrbM98NYi0vX5HsuHCH+bIxuIojlIUylUfQqb6QKm3ZRhNh
eNaA9Xh2zr9N12De87QnvtnuXZl1MKmWzA6CnKvuZ90lIgsaO/6Hoz/m4OgwbTV44xVAOYtdEpfR
PPIIj6d2nHmXzhXO0fwi6VBXsE/i7y0coHZkl/51NKFrkU2rWb8SNPlvnbrVw8mswuDRORNXi6Zn
k5SWtAge8w6lGl9Qeabt+AWqI5hIwwthHiMbslx+WTH359/OE00mvW1hWVCRn2XUs9TnvZZkYafH
QSDWmA+HIBC+lV0J8RyhDJJf/kiH39npmrHGEsavW1A7UZ5kqFYbetuRWVzCdmhrqhvIuJYouX3m
tlPPdlcyJQ0WrpbN3pa83bSELXUlZYT8tul3mw9buXOAvW9ksesKaJvy9DIKSkhyWjniKIm/I2LX
0jd6Ylvibk2EMhcOp+rJYXBXQlHvho0EICEiHzVTiLRbYC0XJKXr0DCYspxl09KeqEZMfUYFYOrV
mdZUNN2tVjWyofz5iB5h0drqZWjmnZ7gxIw5g6inYY0g34sla8UH1hsOsbn9OOP9K+DkXBWzvLHJ
BMEz77EqkevSmmqAuFitA3n/kWboZGtG6oDKJXtOKtmkapVpgtH395Q6Ook4Q/UdRCT/dlWPaK1b
DE622Bh9v+Ay9yBaCooiJKvCtW8LnjDlFXGYIuVQ541xzwennSgjeOvdH4ThP28R25SySWZE0VS7
UMmjBvA2gY0DJmSQZTXV7qTopjRG7J4o+F+HrdjDHMMiVR3s0yFUJzaV110EC1prFaIoP5GMGCEz
A41FKa09/mWGIylP8y40x3ZopzNTl9Z2zqMqiv09o9/Ea+OgCNh7uSTChObNqaJ1WwdWB7KDzdEC
2K0dK2i/hds1NzDIu8QApy0sQf1WpTmemUkxskK3LkigARNDE6DYzsIyaFTJsbTQTt1aad1vgkM3
vsxwLPpnbFCZDhuvt8xkpyprEgeV5sRw+TjMEJ1dinCO485XzyK0RULaEUlyo0myJdAPrZBotcQG
M6AlF2/HFPkQs/xXgj5C+T+DoP2NcPVMF16GvP6jrbyYo8mRqeNel9f349r5Fe6Fc5OIRtt4uPDI
euInUM+Y6ZzrWwwZ4kmGVZWLj7Uo6pmnhqfeffKqeba+i7RXWcPzWKg3qFuQMciLhAKYkYsu+yLA
EXjwWGnowR90Kr043wdgCwyIunHRWPnkjFc5nuYV+wExb4Y/X2083ICv8XjUtRE+vvnMZ+j3MaQE
z64Um0sO/M8uWJRNFSRWnQAsz2TAM48A8O7oLfySg8XGO+HTIjb8a2uzLJGZr/V3wzY0ek0Rv/Kl
RLWQiRciu/MJgRrSuJ6ID+z6nckxL3PV5fgKf4tdEIi4F0HqvT7plRhDeQmze5NrQp4+sESH1vCB
2eMwN7VNcl1pQA3Fz8YRoVi22QETR3W4AZTjiHFmfWfJTbc7eLC/5gto5UbPZYyC90XDkfn27n9s
oSbXefxb1vdzqbVaEyGPDRLySWS6DwcDIRKX053xOOZJsjamyVt5n7YDoNbUCp0K6BHGpsAndkgB
RDh8Hzs2XBJvD42BWrpJ8q+9s0lAXqLhruzdWZrGigIytBM2m9olyIKoOMvdf9qIQZ/3irONMRQI
th3WGt1c+nC8nQAuhW1hDOS2anDrXsqFktymt17WXVXNPlgzx+b9t4McQ0EE3Hy+6yyXE2FmiIl/
sM1oVfereXX0RtXBqvnwLRmPgkyD5/90u5MNE4Ygn5klFIFWQR7t29rJnUxiO9PWczDv6UIEDObA
+gKKUDLeC3PEGkGE/s+blvGAPQnlBNGezeUsxwjWMj1vMwddoyxsbTwMc5B275H9mixC7ZZOG9TO
HPzSmGlIli5Zg4JUrpFBNnVEHKSHJfAi4uQ6m5RJ8FquiLCoM/loue8BlVGk6QH/zzIoUZ1Yi1pO
LT0H7L4wSXzikvN6QKAhLaHhIfS9+Z/iXGzrlw7nU4wVgFPZH8KwEz0/PXp5cY8GhyxMs6qgePoX
j64rjvVtGhU7/ZE2nakrVDkwL95oAJ8mdEbbVawvnzbCehIEztz9CsdCsF6AKoMAExmnM5hJQ/PW
bDweESGNNU8/IW3sarh2VbHbgG90ginVea9301M0py/eeTrrAt97WiB+ewD5In9h3AU2KfcX8emj
gYkuchmZSYk+Au92GUrqzT2iR9WwqWIJpLNg0aMUrpO6Qi6l9gtEndhBeixobmeeaDE3e7Gtdz4B
LBd/iKHK8aQkSuJxDyb25TDSgEETPG1+6e/y1G9L1jic5Wl4t+w9pJ6E00K83k57sIn6JI5torUg
S6R1SgCSchET1A5mRRPenx1WVctRzle53flh0iSbLpO3YYYxTXB7cRJivVyOb07XoGDaofFoHVVB
BPPTWlth2DML+RGh84aLq9Ltuc2f1qFkf84CgBI7/o5KAkOgN6rzoJCKJyvsL45IxA0TyQABkE51
3zE4mmlTWAoE5aRCyaYyOTtRiwI7haXdbA6aMTAmSvFZoPMzxVgeVmqIERw/nqw4lcOSScBm0KuU
OM5pdj2/iDO2yeU8ShhAL1M35lDJJijsWH/a2w1tkULuCHipc6uLG7p32oNCEpLYHVi1K6R9DTB2
2MQLm0zaT/8APAFwXeIQKq0lcqUlvBQesQ18BQsxz3ZZ64zmXsMJcfBLBMi3eqLNW8aM9L4gu2CT
CpVUR/v9O3E+p2JG+VUiNDkboixFvUKRRiEU+HxNg6mmGShdctb3q32MyNlauR6Sb+5iZr2nphVM
jML8nXwObYcB1uhuEb2jRoGjEmAedUV1ZYeGwIS7jqBgIHASky2hLm80Zlg0FXuHxzS/ygiTkTY2
SwX+Xn0CVkHC43TyhdT8CXexlQ/Q17sCt/RB1jtLe6GjRB8DsK063kPUsZ1mo1i2xUWd74v7Z2I1
QX97eTboOoNHKWbH6HYdcOzLddWJvXA8qxJX12Hel2SdMfuMEZXB+aqPmrxYJeJMUQfJksmK9ywY
cyM7j6SuOJQXf/eEv6D6Olj2QkPwuiKHpw5zhFesIMNXeQA5+cyFyluBn1+zsBCvL79aoQN2l8lf
bH+mNTF+fFItsETnN6MTuquQnvxvv7TINZQ0ZtfhpoWNvEdchr2vq23fR1bTqVzZ1H1H7revj8PG
Gn8vIZBPdQWydySU9cIFvN13kWUkg0TnINQaRPjruXYIWgVtGAoMB2x5PkZd0zdNcJWnlxzRuBYf
z/MEgQYq1cW4mokF/v2d0o+rNs1y00XMknm417o0XFNX7yC4zwl+W2Wnr7qeUBwhig5oUzRM9ov2
2rieLBMILKXZN9W/rG9cudUVZMRBiI2AnoGN3nnSil2zMw4D+sF7kEtk5jUSkkSVK+mvqqq6EEGT
167sm6dkmTlVl50isYgptEeoOQLZaurMSr8hn0OdeypqdaDM3W7Uhhi5hSa4gkPMLfokqA0JkJdP
2jxTaa0I3BIA7zYrA7ZzVN9xbev+23D0scXjqsOUN0xewiUBIgA8nB3rCfDQBsVv7GXUVa+ZdOo6
iGxNXTvFCtiVxxIP9nsssRYRLcpAcDWKl4GNliC88sa21anU4yrofxjyoWFUs4x+jnN3/q3fbATS
Xd+SmfTzHozBIwEQZ1LEleCkeXDo+iM7klNc+V/z5Zrzty9d/OaXjvOBtsEoipJWwjz0AG+D4EM8
vJEBnmIcURHiRy7M+JQGLUQZs/8JlB/No2MWhbjZa6jm15K/3NZR7u866U2/2EEEDNM1zxySvZiG
e3ZZbGK6tYiFjN40/iReKkGBi4rBTYQ59gSsdcDwF0m+TaL/F8lFPc0y97kjL3B91wcuyv6NoSGF
Z9NbtTxugzbkcPV7PP1SOvkStdKSqFmjhfYmfhzYerVY9VUT2jgMCgEfOxwRyFib9DK61mqZjFbe
pDtDoN4C6QRg8p/dHh3J6qE2RrITvN0R6Y2qttGUWBcx0womdurX99NLIkzNGe8eDigqx07Vcum4
cksskFDfwx85JvqFEKPjxQFy2aBc3xdQSYPd/0oxZM5mA577r49G3s/pXW3qttsY6H1MkAV4o4bV
dBoE68qIvPD7ooR/CB2EK0ROJKiyN2qY+X45gW/aWB5Noe65dgICORhXgVzn0diFLIsQu4VvBn5L
N1y9h/g79B3yAIGLAnGMiFhWs1CSMYYttJyED5rtNxDFuSnv3qCi5TbzY7tbQKBVe65HjH5oB1uS
70WGwgn33D8vE3gJ4fFro1gxl5Ixg2W1gLhaN9Awvsybx3kO2xceNg7IsHq+snkcAckRnXCbuN05
MO/+vPLmWUGwLpCh/GoqPNGKiuLpgNkLG7Z5mckegvn2G61XyiTK9DVYa3nMxlnNtDqi9T5rLlyJ
iVYP7zL+J6tBrh6fXg+7L3DeGfWv8uYaoGMgCVZWE1WcVDVMTD0w1+/An5dMO9cMQh5bgBSXdnMh
qfobA8HmRpDKAs6zgOJMERIeQFXi5s8Z6Pj/VVBw7jGI5CJ3XzhZW2KWLK0Vi9nQKy8WxCwD1Tny
0i9J1AltqTQRKC4aANVfzDMMtOsf8W5q6MqZOvVOO6WnKTnUhbm+DsAIanLBmoiLjV4JkaHm5n0I
hBLOg/YFx209Jyip1NIZS5gajSx9sxWcPoX+phXBasmHzdJkWLasavjDD2E/E4cbWsNeMabIxZsx
l1u8RXYJtJKSfLWAcki/PQM3AsAT1Q7x8ZF0PCtJDmYVmDDtPw47MCmCBRdj3yHuj0JR7aEswPCO
7eOcpkhxgx6sVh4mlRoEi1HNMtRY34unc34FgI2rr2MAOOAJtz0qdCEQt3EJq7TuNQctm9PFeH4r
H9T7UelL3rbQ/hPUuzriKFBVU5Mhxj/Bzsjuc9bkzmblF3tY7bJLhrjcyuaewO9sAEdHVlFlSxsU
/WoK/ytCTzoYlroycHCux+SyFTQHYa4QT3iktyjQw1/bA63fH9M4/2kcqcUj/feJ0gQa1N5COy5p
bwjBSAUUdwPCS6douvHrIyWqioUwMjjAaKyuh0OFcQiX3pAiAqgNQ2vr5tXd233t8RgZ0HgsUNst
xr1X5lhnBNuUdP2B730NbAeHafRoUrQjw+ExAiXiwZHGdhrzpwOgyESYDXU01kpIwGD0OWFMylXr
udq5ZdrEFfBPflWjwhHvF2UAkxapMEfIxbIATEZaXUYQe0O704SePxOUdYr805zqszUgpIydZA63
QN7/jrnj8EDOKaCqIVE8Ge8EI5Wc8caxqCESQgm78bMzGvVwBk+qDB/Sbb4FReLwqV3C5HIJTiL7
LA5AhIBInNdE97H1mRj28MLa2y8VHzyzJpf/825l+QepvTfNgVQ3LEK/v7FWbQdjCZRIgxQyMVrn
cUAahJzGyBFZQ1oC5rCcvrh4jmK50Qy0wzsRRHoL6Oh7MGjVj6Lroxxk6Z469vQim1UR3Mp2s6qk
f99Kxc+f9wMXSRaCWq4Y6ZbJhnraC/kutI7lP73KqVWVJBkrCUj++6dnGLmUckGr5o4NWiDA5YX9
KrTQYMNUZK92VVtypE52R1ykaTOEJwJtmL7/J+Y79ID0uIcSgVXDYPqQmX2SKt/aOTgYwiJRGCuu
TncqZx+FdrGUvq/J7M5qeoMPmjpCkYe6SF4Aojredh91D/lge5aBHsrV6i2952wyqigbCe6kzwvo
12dhdXm6Z1jRHSm+Z7/+DVfSz24P8GXKH6XUVHm7KCVfsAm0kRm8nSdR6T52NIkQJF59vf4wtVrX
ioSQq0n1Mp4PAFFT+AAhedJZunR0ZCGQ23w7p5FtD4pNS8qerkHjw4zMMB9aGcHcmfl2ZlrOEi8v
pcx44v2uvxDYYPooCrIHazM+V5rnh75SLut5qgfz+NmBZMHmwCygVxcKmvk9L5dwrHpatxAjCpNI
+4mC5Hbyre9OFvt0FUIhTJ3vYlQNFCjefh6WK5FlLz/NlE4fxbSIvuK6nTohcfU2vcawMvPlmKRf
tZFxPls3laT6RM5D7L0dNVkWIIZZEzagAcekf8ghByKJWCejg8EDGMmBsdAyoeG+B4G69a7JQZ27
GenwNaBzBWbsnUQdD4/enwh9g4H1m3nz9iYw9tcLycep0FBiqSljnHf+CzPme+LUDydzy11uD1UI
AwV09DKwx23Fr/A3qdKTYSHnAgLWjNbFlK5atxo4ct1SLCarZNUnRNIB0n/VKzkcePLpMSCFnezG
3xZdflJGedRclFLMZy3JBN1B2XJaNlzr2GS3JwhmJmTyNNR9lb3h44OF75nzwXqyruU2Gpa7JK/O
m6c4KszZCO4vwb4RcQGS6dD2+n3TSkBAHc25LeUq0cJ4O1bMeMWTd+slwXpytx4+s6PIBmV/9Ty4
z8O83C2MnPQhvzmV1C7TUmvDEIwu8gGqkXptu6qRwg5VckpacTwzjWXukS3mP/tjrQm8deQu6b7w
muD58+zepzPqdGS8ah1TGzxNnFVxSax/jotSaRAa34XWcHpI2GIGABnCVqueAqrJUxYlXkzFr7V6
Ls2x0iCAQi44ZzXUQMYIRUefrqQPhbPpAIma8ERcQHHp5l9fGcl3as2tj11JXZqMsCUaJIYwo+7Y
hoR5oZF3h1YWNHkAZ7xRjc6XQTHSamar71rodVHiKzd9jHnhTPhHCcjam4uPNTt3bpCAfaT4tBBP
nFH5pSUHLxj7iNUhiWr/dB7DQl8lPFGVEIkNwiN8wrErK0+Yew+RPIyXz+5+fd7u2fMXlZJgLggH
dtve50VKNeMnDmEkcuBeIGxMreC1w3/2n8LmpLjf5SYDWcwVD+nzLARQDGiCcQwQrNcyGgavCuZu
xCLNK62DfCo1adYTNhoTw/Of6aow7R3OTLMmQuVAQTNzj2wFrxh9oMnHk6sYQF49AQcApU8gBF36
vLKLk0X6+y5LNnG2YNhpfry5+Q4IwneHEwZ3OUxxxuT7SpKeYbI5Sx0iKuvNRjkcUiQbyWBSPWB+
qpFjQrLMHVOeCk5mSOFmm94Z+Fl1SZYb92FbGYQjcxdrt4kBb5v82dQB+TW7woGT9V2yufGzb0uj
C9wpW0SH3fe4aaJVikFlLlwvIa4LzYBNoviHBPhos9EVSN8TUf3fygYkUC/F8mhHGXXl8D95t+8B
/0kDhH8aKvdSn4rb09uJQqJLteJlcy+2gf4aSeAG8pKQpIclqEpx7g075R8wuEFZeFtOVknbxbpz
9CmuMo074YLgJD6hPMBks/Pwq/ZYRrWC/SMbrR8DWolTbhZwaah6fPDKODB5nsdRxIfOvnhC0Zau
nP0IzWNHclrAz+FzSWpfc0rZ0bNMcqbBDjednM1lV9w086r60iOuGIACkYowSsZjWZ0jxzCdUARJ
8wPEf34Hv7zLZvjVJvySox+in3i/AE8y6WcbxSygY33YH40hbJmrUJy98S6v0jEghHF4Hn6goKMe
yFdDyKUoKv0ZMrcWpsA0+IHpYCJ4CkVy5CPO+pCJ8D5Xet7pmwGrY8FKhRXajUOpk5dzVbUei2VW
SNPirY7BSZAzdoMLme4bbDksPJm0Nu8Ugw5T24cJ7tqcbTmJh5iUhWFZpMVvgfWx51hTXI5tDtz+
oSSaH02OLeO78FbEQXKRdvc6DPs+N3/MaIs0zPWQH/NtxGzlX3l8M1O7t4L5pwK70OINhUoGNWja
pX3JA4avgH45bE0B3q0F2P0HnrTIOQ/sLTOZ38cKHcRs2y2wGqYeqUkTpULQAoC7tx+EbiWX4KYi
PxbDGq0SRLTu2FFOdu/8vpZbMyM9mxzOSm6y5cLgObiRh7Ioc5LJJjrKBciu1+JAP/kkDaQIjPnl
RL7FDNyYvtBj44+IFlYZ092vBcSlm7z8vVjDwhgUJaTv3gkiR9IGhcupSC7Wo+WMcpI27sxNyCd1
Su+FRbvjBgL9FPHnFJ4sOzwFlrL2d/GcYYlVy//i9oKLzkIz4QgPI/TRKxVHdz+EeBkjPU/37ClM
h9LS+4QrvUJCzsHdLk5oAToXAf15U+P5RN8eP6d/GpwkYqmbEfDVYoaBNw9RuJXh+B56VLwUW7Z2
yz3x0Xu5ztLI5OPD8q5VaA5SzlpGGlmIBIOm7/jOa4WyJngwZuCKqy/A/E7wgBzX2zhht2MTy1sA
oui5L8dI39n6xAwHekZDpE1vVxww1EXa0MQ/JRULYt7W1TszoUUzAcz9XOlYPyklzDgQnjrkOcAK
6p9HhNfLhr7MZdFBmCHXrcXDslzf7Zgq4yaGgNZzG+rWDcSW6ZurH5p8ucH1zjHJZJA4aDyFmHJa
5pKf/Bc1tbvV/4nC852xsfA1DchJRhYqXUzcl/JR38pyNTB8ANGCdhX1obJQ0XXG4aiFwtxGYERV
qRWW5qQkvSSvI8mvaxtdXfPHVnUEinuvQ0hn5K/QdcX7BUzwlXCOKP+gLU+gClKRbHwtrx2HoamF
N2xGE/cA3g7FkHRJbioKB1U+c9ezmTWXDcZxwY62vA5md/JVV3F6qoH2rro6SUWtmVcH74HumF30
NB+cjyovnVDQmJIUcjTZQb+Q7b96KmW7lyCh5zt6M8TghyRqV+2UoPJr4v8Qh1myzQgR0oG5mmK2
WkDdeNPShajZ3VHYvu8OCU79G7QPcLkcz1ROIrp20gacaeeOaJt9xxrPtZLYfJNBB4bRqvaG5zu8
7XFFL1azR26zY9pE+WFXmVf8ySdxWMgCu9cEzcQCtxSu0PPCL/p4x3kVPSlVEK8g+GQqaroND+Ei
KYQlLQAzuXUKzedL+6ITe4ixZMLnDNkwvx1h5vQ+NbpmNnNO+3Y2mX89gqqLdbsZZwtEVPFKHEUD
yzEZMzreMPpIFClDLecyAueOnI+CbYaN2X+zfKxiJIAz0UgCRPDbQTwYkJqSPO2Gi46JRMVpsWK6
kqp4AaEiVh4z1x4USONVx/1B/KOz5NABvtIeV0FD6oiwBmMZKY7TQq5oYxX4BEfJrr+9VaLpLRvE
fN6sPFCTrpOThToLUdAaN1uxtXS1h56io8w7JrBWmp7OaWmp8iLmxug0N3UabfHGrbJ9gIZPp/W2
O63+fUUQu9pVkwgVdumoNbMa3L4ZrLrq+A5jOyRwN0X0XBb5L9tkI1we/sXYbUNxHRVImnJ8njD9
tFtt3JS1w7zLKoJeDCx942yHBmqXmUHwqXWgAbh1lrPTMV4nNErtscrP+7aJakkg0JqspF4famZm
sK3XHsYphY+F6Jncvtbpl4gNDVzuDdAq5AKiHs6EES5iLPkK51i+2EuxMYe/lYHTEDP+ro/aAN9o
pBUI+PhEZbzP5xqeC79vdM0AbOqskzGpOm2rJwaFW/av+yhfJiaAsqiUWfTT5xJEuf8IijgyMEDR
rrzKHUti9Oc9cvxxls7UzAfn8CV5eoJzzKqSSRxBUZBOUex6hlY8hvDDn+CyhyvjER1n8U8zYD0p
GDOU1oeD8PGU6RxpH0jXG1tsMKQS9ezoEUKdSE9yj/lsQ/CgRjrPtX24+RbsN8TaRELJhn5Y72lD
UR7Ek46gg9HhfHor+yhWB4vY2jDqfXFHTpAizDyoBfFiRdUrD7bau4SrHgbLfcLMYZXGghRao099
9NQOrqgsKABt4czEzjAfFJjruGeFC51Je3FJdPQVmzGZNZcvjIADTFcCb1r8hgiZMT8/lxLMd07U
7WS/kStua4Fl7KIIYiNz/lZgiZOVDSE7VmpbG755NlQi4ZMPK5IdjKiIQ/KMFO7MhZf3soegg8L7
zUlHpTogRl7fguWkpmtAfkvdNnvxHQi38lct4AXe+H/zBQ73flxFWu9mbw9EjDcRq7+lNPCxaMvO
qy0I3UYe29TzfTNCjYUaztF5qtIzXiDOVGL+NhIqYZuRMuRgbj1wrHYnssNemlye9CCDFhxRruDD
CXOAxwlaADDF37Es5ChhICsDwM1NPEjjeOD2IGr1/SbSZmXRzHXXJEk2Cp0k8cDAIGGucqX7ZyNq
Vdp8jbrOW0jvgQUx/EO3NuLU8PiWIJ41nPYb56cLxT2G0+iHGCv+fqJ0O+UfV56B+125CbQeIN/H
KLZTcM+qc7wmX9x0Mz8Oo6zDS0Rys0kGSO69S2ILdSeqQEfrK3Yf7bKI+4cAoU9GH4xyOIa5Zd84
mfRqE2AiJ+xfokkefqIil/fhLCFKahQCKdkQIBAVXI8uRwv5WEvIzos7d6C7eohoEQLwI0rwX6PT
zl51GIoHEshOQINzUxxnl/hXxZViLyF4FJncCBkiiWPhTPIR8voJAWzAislx8PDTTeO9A4IpOQjK
iRjLaTUg2FLG5SMtPIl2bTWOpA9ZHLFESkRVbGsmcQjRIMHrzeQYxzJ9ft5jkDyNS3UWn7YB7zyV
WsHyEbwosIITezkUYFEZCZlfPLekx1ISreDPhsRxCKtb6+od5VBEYz8hOmcWJvE6dm62ltpxwTvk
BnTzHO29bW5nolryljQzS4IYRJi9/WVYPsEeoZ/IiczKTA7q4DgMsm+drfOVnybElHIjSrFSXWLf
sf+nKalAzT+Y6UE3wJYVK+Z6/RXOp5OmuC6rOdLbOGSnlTwsQLtcFeO1DKK5MFjuIpF+hnxz2Uh5
AWRQIc8FuUKbUtU8xz00CwCDBaNkvk1BXxlKz3xrq4hoawF4Wu6Nvuk8ssfur0fKxCAHiDZ5o9Y8
QfNZIqFJs5MHzxM684a+3+pJMxfiRQ8/aXYuZEYYjMkxYBiJrAi/cF3NE0soUoAnnvcUURcQ+0dF
VB6UBsk61vxhWvQSM6AWlMDLcCGw8qnEhVFvxdqBxTnzdR0xZ4MKUZHmoGpfkcGqWdo4gu8hodJG
z43s9TgDkdP3oLJCnW6f3kujLmYdfLDLbuOVtb42+XohhgDbtGRYJCrc8h9E/HsKkXqDjLty8KXn
wPhjDk1/NIk1M8cHa5JQpP4eQsq2KTwrYCqZ+YxJzmcqKkwTEb2w4RGjHfA+0Vaic5b2LY/bM1W8
Hsm+WZUIdbiwQiNkKLPjwQi7z7h2tB/LBUjC2wUOCVl0wai9JimO6Ajp5SYp2o7lY0y3nHqqAy8j
PAkKhppLW+JE4jn3ty66t9iAdpAskV7dy8jJy7Tqf7N+XyUahxvuab8+6h+4ReK5FqgdA29T1HnE
APzYmYwMh0OpIoHOQ9gsHhWJop2g1xy9Mjun7C/EuPv/T1EEmaYCKh9WqNvOVWYmIuKQewJUh+ub
CJyMe5+fofTSuV1ZBYsi/zxFPi7P8tuctfYDcMriMGJzLcwO7EvJLUzulp1juRAY3ubL5IrztbPg
RECHLJNBJU+cglgv1w4FYS05dsPiqCW2IBtDKoeaHFJW5wNpgyotwUfeP/PFUFuRSQZPcLLUUFSR
91o4ua3JvDEYmOkvlHKTk6A1DIgHfmaFwPF2Rz6Erb0huVkLBJYksjzOEZH92VhSBxU4Xym2sb5p
cLz3atf22p9+1Iw3U/ecaT9RZ8qQgs9DJWgXDpjTVriDuIfPtyjS3ifuxMmdB2xSqzs0sb3e49b2
CwNkBnySsfLDFnUZv9uT3Th3uJ7/TNI/UrCuD79Rizt07HtejMaWT+q/9tSRygLsfMoHGOnypLKK
yjQlVXAKojWFvkKc/oyj6zT0R0g7WNiNW3B7EaxodYmX2g78iP/5PfPzynmMSbfRmA1nwkh4VfrQ
PEhAXer37MpbBtkL68vjMh+IbviIzmwqRlbmiChq5O/VLG+YLVd+ZmhIPkoYGdr16LtxKuQDlUyz
mbh8VTYM1XhIec61dMVQJdGOSYQZoaHbBvnrzzXWY3SXcl9yeMBscgeAIQ7vyM0ZGq736p+xfE1p
HKGF7fLTWrDAbzbIym4vnvsnPcu41y+IccLSXVR8cZrYuhgOiav8H39sJTuCaDZs9MSYq8EojKfL
U7APeGprkMiFsee2gb6C7E5H4EJ8dGAsx/ONm4OytMpEboNg614GMS5oDMDDW/lUfIq5KzM4hpv8
iizTIkik6yzvSHsogGVd48fSWOoBuC0nkpVFEzUHeq2YhbHzo/njrFhhvrTLCD4U+xNk1OOJOVde
1/kEa767xB+p2z8aaeQLQ6VLI+wXE8hwurWj538JtdC6PxkRlM4yrtfINc+678WrvZg3pQLlIK6S
WzAMYcIPFajyLCoCB4koU0KDWCwmSfG9zL320tZ7pT861j71BdCWjdPucTqsCemqDTJTR3Knqvjj
wSVnAlFDXAyD7qW/q1t2WJE8fDi/awthaI6iZ95Ewt6p2sXgX1TlxdRgV+btyNBJ4f/+S2BSA3Tv
1ITUOLjuj058MEeqyzprgUrHqbFc7hFm2kCaBvy/KYtXd28VqZH786jVKgJ+qLmEioPJFkLEO8BO
UATxLVq4svfsy1FzoGVmyl4MeerOkPf/fI2L5yVYi+M19xwgSH67qzRJKKkMsrqv7jrcgzXrGanI
5ZUBCW1XY5YLKcCFQF1eHRdCyUfYnF2zJgAnYAOptz7urZMgUo4mJL9dw7tSMab92o3ZwoTPnX21
Axcrsw53E0HdsAQ0SXSZAbjw+8g3NkLYaG081NCMeCGXZNKCtq/12B3C6pQB9EjiYe5izQS7E2Pn
rsxJ3KiWUWt+IOswg/izUwJarJzoQu8PHlziuFjtfZEMTSoSzOSWSAJmVvJcytat6NacFl0oKBp/
/M15xCHXiFgiHFGzQgoC989zTp8oL60bEK4FCu1GS9GiKBuzxcML6Ror9ZcRSvj/x0xRDrVEsxXY
nLjUBZQQuVWpHJEPKAvr39wv4Hcw4qHY+OY3fSh0YV4X7b/ufsrXo+n+l2Bgl0i166UCH7nRvUlV
iaoAdURjsGf0QTBOP4gXtbEI9qChW/aMW3cmq7OCthrLvch+mfPxkBS+PsifyCrUE6YFYt1IEQma
qI4GEfAWdTJzA/OZVqoNzQiNI6AHaQ1tQwQy6suxH4HW/WLY/m6jPPxBTZFEP0mZHOnE15RuOF2S
1VSJww7A94v006XhBlkkcRrpE+CflgxCNSMJIz36g1oxPB7VPg4NzelrZfDaKU16hl2ZqMn/z7lC
LhE6GBzVvUNhBWGD13LesbShVSAWKfuO96dsMJiKLZwsMoVJ4JdoHTMXKnRPYsItyb9K00PEcVKQ
r7bVboBMWEIGOHOabSlYXOs+FTU2Ssl2v5Qerdl+VFKZIZ0JpQdOGDhVkBcKR5MjfFqD9FZArtez
uS79F0BQ9eSc9ZXqNrRKTkiSYph0F/WFeExHrf/URig5oNySQIfj1IUNkwEYn/H35X4qJIyime3X
38qd8L0Qe6Ue3luRFR0yIbQM/d4wcQysPLDTNQ/8Lr0S2+p9G2IuH0SyRiXz4RPHCOuIVIf19ek2
YHC4h4KTiJU8j7ERR0GdyNPE/974O59uS9RPPvoUVavkWFvm2/5ickZ5+N8a4pk5mPpq8jPMyxRx
JJVum/RyS4LGUazdoaPd7dg3eepQD8ezhxebrtheAp/R8MIMCqcMlTUMYcNZxuPmjBQYM2XQauNz
lf2wLnmohPe+lM4wB2xp4VcKZZc/NiGqfnakMXNDBz17krSD9PPKoScMZj7wSj8ylqM3QxTT7Et6
zi7CmJvXqqgaCnm06qMYK0a0oejoGd4u1GFB6COcD8jqo3K6jbx+ThjC7XroHRJLNRHZcOFa2g1S
QLGMhlx5pd/V4Jrmcgrf9CHB5DgiwvD32Qpz27Y5FWmT2Z0qweYsa/OAPZOVI/eb7poO4jiuXPO9
0OHJdM/pbHeYoYkLEg1OJ6ieM0dD7JAa8r6wZtqupyWWQjT2Jlw4TZokDD0enHOM0qgbMcie3BZ+
iNwYTtt/RcbcLqn05ZUkwNA5pE5NbOwf8msIGaHaHuE9gsLk5NzTQd2S+thuyyUfS7rmDZAepRfG
NKwzp3bWE7nV3ttXV0FpvKm4/Xbd5CNy5wZx6q/ktNpWcY2bn7PI/W3lpmHoNIL72uMgldPAgIdz
V1uAMY018wwF6qObobLB2lAVYEgSWmaQqR8BZ26GzXgzbY7P8ZDV1u4tISdv8z2SIL8i9/0jrUPF
8s7A8RtCCob9P4PEfP3IRl6sdzSMeHDDN3UdYhRr8GGbpmtoLhMX2VDvviFCDSKwxDJrgOyeKnrh
jPWkgAtG7VwI2mYLoNlMhd4sRKGoFjeD6vqbb+A8s9GVZnI9Itmx1knPvBKi5zNpWUvripF3+nUX
gxyymTBEXyaaocSNuFmvL9GwW1AKAotcJsfeEb76VoBpcQ7CouQ2868bNlrqhUgfh0fhfGbcLETu
HVLLsYiywJg8CLGzqZ3JL3crrb5eH4+EW78aniaSx+TGFjWDMa7bdnegPqybZoIegben1PaUo56C
0Co1Nk6EDjzUxax2hz4qAsMVwlgEmqCqOtHi7HcwacSsEjxAW/4dYOJZw2O0FtqwfuQvW/iPslvK
OYNFAHdsgzIaRnAVIkK7GVW2Uum6AyuAJnBAobm7F0X29+I/U2t0sm362dT0yXCL/UWoQhCjEmDD
ZvYkVJkFuqwI0t1AEo7GZxd6g86fuzMBGOmlvAsRR/Zcf9us7+1mujYkHh+8O80eV+YRB5Uef+C8
mff+NVaVSmFG2KR4dlc5h8eqM0sGQe7z9qjgRQbJx93rbh/rHIAi05ezya2578Nw7K1IfYFPX9Sa
fIdUZhjazjrsW+qPZkuE7eGJ7mbs9xXkkKA3oRUJr64XM08UhpibE7lwnfRTJE2IOGah/XTjIqqC
FRgWdUN36LhTiIlr52yWc4VDyaWe6abozzeteAQkoP6QavMe9DaA8z1sidSEUiUWJK3LEHQ/lWla
0gh0osLbavoVbNeND18Wv+rbn9nTHVOCgI49p9EVRk7+GjVRZh/deA1Fay3oFwfs05Ao5PI1PxSP
Gus/GmHMRGmlu4o7p+i0w66XmkzacqYkKIg0GeFjVl8MICnePhxkMnT6mtgyaauP2TpD26WRW1p9
pISRN+gQyHcVf9APUH1CNtv7LdSjSvg6goV+37axixCnmBOlh+b4zLjQ/VUVOInNlkq8io4AeICb
jRA31k4rbfA5U8ZEBxoYTiK+khl1hZjQArYF95e+ZgcxaBtyNeuWCnKH0iVT3lGMLredCS3smaxX
sTjfMiRFCoZ5K7Uh5XcYLYvqFy1RDGVnIIrGfN88oGWTJrKSd2s3dpFm5hgIYpGnyMVrL08m0n6A
uZuWEPv0W+l8qiPGA23R9mxnQRgrphiVNJ47McaoJ8XoPFmM7Dv9QDl4dw86M0STQA+W/UMk3IkL
I9hgIhVCqSpDSBt29whDXfnKg/NYBeLb9N3iTk/TME5h8ElFulVQRj6gzfguD/E3AzbFXWeaeAow
f0eJD10ZGvnCVTMklFdMK8TCc3NWliDMRNa78Nu9gk1uMVAyO9fkjPd1qn7XGDOHFiw7qfBGE/uU
a75kse+G7x1KDHF6X4ZwEQq6Fu3/E/IEEKFdHQ2/P8sI6q8wGmajc4vf8/JEbXF7YXYWMA867m3K
nmX9B0svE8mSvdQrtIhIESA1li9m6b4j75ARFD+3sKAMtLPmuVoq+cdk7yUVskDTu5WK0WECmDHz
P5HHt8Y51jWSAAb2SjpHKeRc3HQ9lekOHSO+Tg/Jjk/D1pW10GJgoI/HIBpBV4hgrsWbnoy5etnu
VG7OmNUOi8y2bACC6O/YHxABm3iC30+z3ncXSQOmfd9iPDYg0VAh6mCoZlAKX5gDwbFDhiygaeZo
ei2QKV37xJ0xbBu7YbvvgxI4PJ5IjhEoTtyhvnY/Ykjukg2NMITOYplk7tiUomFl8syPtmgHWTiw
lg7x2nKSYxL+bNactQZjjjy/T3xi7sjiMUpp6TXWsKZ57pkIYCC8Cg8T/UgobkY3IYIaAKBLBOfI
RkADGdHakMukpu9P+Zy5ECrxSnTuJMdCZ94QnZkHX1rXiVfOXQtBwQeksWUduAutR3Ji5GiFAmOE
7gnK6xAiSmxXa+NEfAyqyqsafhjAOeNZYZCziI+LNHnv1FbUnlkppkli/+KnWqROHqEEgPfdCMal
Js1a9fXfPAxvvPE9bBITVqFcPHJngxLgEf3QSIRKAQFXe1zC7JbWd5ylJZ4zyZLWrUGVfeuLtJSB
fEzznVzQN1vmDVhg+s+ruFcodmseCRTAU3D/gnTlzGHjZo7F3R5PmqYAALVYsjdLyURpauKC0Bno
4lA7RZCNDoTT2kFd6T2tnXxJlPKpQPa1Ea54cRZEVwSP0ZWz5XQGOutlmUDp7MB4ooyxN51saUnz
uXfhLeMX/NhdeHMDvhF+K7QLwJvVNqEjj83Xp01tMYM0G0z/58GKLnh3DBN4UD5LToovyNyZL4Z7
mo6khhvrLl62dFIjYJfOAeaV62m9VxPRDK3aW7iugU/CNByLSbxWNfbK6Ijm4H/1kYFmaMYBocN3
WWSw9d8F0fKN4P9KKvwmZ3OaSaDEQc4oB7zrcaC8x7GA3iFWo4bIVbGPNTOBXbZwy+RxnMD1XDKW
jDoqh9BW5Nw0hn1M0YlzMumYKvcm5kUBgeLkq5gPC5FcOTe7lLGUgvHi6SXqxZTf7RfrpqtYZZLl
INGzM/VGhPuiFjaeR5o53gwcLmIH44Ynmqo/hAIH8kZt9a7UwrCkz+Hn4eprOvKlRWcSsloN7xnQ
QR4DUC6A7KuailSE7CMJEXlHKwFrW4Hylk8bDK20opr0UDFbug4uElw77AtE7dQISsO/kAe6i0ab
KVCo1pGT1kfeVkgjdlHlVq6rLLI78Hw2O16o7s5cU1ymcKfD/PLq6qs87dCYh/MRICF00D3P+wlU
5ejrwV4wacY33GO+nmHsm6wGQVuPfXh82SC7ZAD2JHX2xQ2MYR3wzp8SazgLQAU+PsnOUoT+e0jU
CKCpDb3oGmirFuTxgB2fFZIKR8aeyp22oes/DIAOh24vjiBzEEBywBg7pUDZ9qbZ1gtVuF3DC3fu
XD0phayoEg1RsLz3bqszAJv/vCDjxFic2p78CBJBJHyzXTsyON0j8pq4GRjQ8RORbnxg3ToiEIXp
V6mxvshwtd07ZThmw73NxjfbH91dLBuYg8xFQcJmwkd+LxO1yNlguVRuZbs+3NvnmN9BbcdQwf5Q
ntcNSmOom2gMLLqKN6qQFtNaEmhuNMMQTfoaAsIiB4oO0+EDb8Rie29723f+LcYI+SFQTzTQw3jj
pAwrGbgaOXcNoW2+TihgzgEwceAQ2/vwf9gU1PLzsKQKJNAeRuPYAdxmidXB5ArdEDvTCfmnt6HD
y1EVSK9il1DoSVEfPM/ci8ZiLEDawS6yFl9HLmtt6j4DT2QsKaUgN6TCnHS+gmhP8nRz7bRXuHgK
WWsSwnl7/XWH8tT6EcFvQ7mzLq7JGdtJCMgqRlrN+BHQSawkiRHVunwiP/hFyoI2MEQfNCe/tATS
qJ/nztxUH2v5vRaJJBmbXBaWy3EbEBPCwdWroUm3GsQkySddw32La/28zUEYuTuULblKNWnckiY6
8JwJRGBnKd4wbrc7HvWnh6QTPQcmKBR2SvTxBMOil0JmJsMxu4Jgx9jOocitpv+/O7WszRegDP9g
5gzXyt4AZzaotGPPYrlcyb3RkQEdqWNL+FDrloPcmiv0Bk5nMsyG1kv388N3lKkjU40JcpYNudXB
5aUbJemB1jNzwnoKPArqFLZeEo7/YYcHkrbNdgovwcSxlZ79lSzXXZz6vmCuI7B66e91Hr9wO7DA
9rV6Ayi28mBSg7P6XqSys/vTHvv77EdtgcxGkoGNkzANi9CNGDNQtKv18tmPhXXzS6niLv/YIsG5
T9RO64g+vdWMwYxEFZsFGb5dTBYQ5yZHlListZq0gijWtneG2w4NCPZqoH8AgGifKltueOSqfXeU
3HFNnA7KeODlS8V3aQPAYHFR2O18/fT+ICdYj+BaKCTOccxboDRQtAcIkjzrLG362S2eBiWLm/iR
qN0FB3cYJZ5HsY6sFyLbmQCNAeVi7MM0cV+ysM80b9zV0hm1b7jr1tQQJxQsPVgHTfXts2dGu8js
woWRfR0+vPEQtDT/RN/LIH5VlL16fTz5W7RCX77Arbtc4ixT0OhV47hI1FZqwEujAZsC+htbCp0=
`protect end_protected
