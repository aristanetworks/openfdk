--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
kCRlG7sZjEbRtlgKSkvvx1AVuo9k4W6A9ZHuNBbWvkWRKe40Nf9ljb9ozuq6SgJ3nycB3dPe8E/w
X7njzkvcKgOb6vmn7FZTHv1NaieptzOkAt5x2LoRcPRmiUC0MtRuBZlYgu3RI2JlU9fKnHZ52ZQr
g7e5fxTEm8CD3lDcjVKx50wpRIa7LBOpxxbBxRpv/UzsPpiYEhor72h0IbHaBEqYJAf44wrsU7U2
wPF7JIOkxUsnoR4XrDHxSATpxGjD0YpEECgxg2mIF0c4ME3P3z2hbIuru+9mj+UsnovU5xVICePe
O8WaDnce48DVCHabalds04BA9cBWMfIfuGPpVA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="jly6Hxch1Yg7HQq2sgiNPX2FzOTez88rJbuBYUOgrwI="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
dNGc92vxKVk174mVl3fOfpKLPbYz7Ssj4HjewiecVpDgZLeFQ1EkQj6zRVay3lIf/Db24/wjRamg
ZeAc+ihjrvY5ojkIM56c5D+4Y3RmrOSRgFN8BdaQjTnV/d7qrd85NeeUFyc1jN/URpZpl651QmYD
PjLuKOnC1PmxhfwFwp3mJQMCoKO1d5Aoo4oLuC8N6qnDKSBRoVTCizFaLRQ/SWwgYTIvlrX0AYeT
2M9MeKVcv8cftvSApDEw6zImMQ7OFbYNihivOLkN3+ZyZ1nNFKF9q5LS/UlbR01hEaBIxxXcBfH8
e42V6gScxMFI02nzNqR8tOcDsYPwiNqBhOWY7Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="d3jBu8Y7mL/itQZ+zCUe75YfGEnCFX6Tns76r80vNVQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14560)
`protect data_block
/HlyZY3ZjD9cpQTle7iHwGoRtQk/TRXZX8bav3aioKhtLLxe7W6st+qaRjVN96rdxod4ouTUYPE0
YfPYOuDei9ALtfd1/O9eESEJIUZXJ1n90Uo93mLl4RURC2RagqWIoTBn8wtjXr/GhjmUoj2Oisly
E4kpK8VqnHJL5h4CQfwEysZiddDHduITrjvX9UJmqhl80s9ta9TApx8E80nx1oWEAXYe0AwzGbBC
+dPU5M1GO7QVcre42A7uJobNPHrsVkx57pGUovKJ/XvBh2lHjPmFmAdF7VDk/pgNdpc4+fphdiy8
tIyK5+b2tkYXnyqhYVAW7sHD8AivxmLGq4b6YGnHK/t4fpGMZOsnN6jtt1e0GfJcDpoqKs8v5f8l
kYs9yB1mkL1uB22swr0puLjuI8KpzlY18vgS5wGJShj1w0luR1dNCsF0XCl8tTiTRoQJmIMNs9TU
XuuWwUUGj7KrUpRnrw+EeKxW3rp6jZosA28PH7o5zpe+6SkRhL+XD8W4s2yfRnlqc8hEdvcjib7b
863TzbIBAq/kwb5ILc9dayFJP66scUOeXossxA5f4zsMUK5DUEHHht2Crcjb/7llF9Ry9HfpheIF
lsrhtQLNgR2wFjaTJqEQ8DNWXMdhH1vA11/3QreKf5E56twQO0oYiKQ6dBPKSvWZM7zMP56yOJ9H
wReqGbVP53HFEgZDxouvsZ8zAQEeULKI/wZyXz62E8Ow62EqmsjB2v5/PgZljGkoN6/iXB91z8ZO
vcj8ZBpq7y9U4GKXVkGbhNaw8M9XdR+KWMyRZ1soKkLCpwUSwz5MLk7EmOEU7UGsLaKc7iUb4zDU
mXCqh5i7HI4ubHCbwMMWLtTo0rgthSoP+TItAj/ElZgHnRjtDaPOmaGrO/jzzFe7pEqnMx0mXNm0
YBTst3dJc+OpkQ4oaPUlM8B1xguCkr1KI50MJ5CbtwRulbiCvkhlNh7pvvl6DsCCZyT4bY0XyDc3
X9CsJYvGPd3zvhJHdAI90j82ubX3OcHtGvBqhjY0Z//Evv1yjhzkMthqqCWB8PAKuKGTHv5+oVbP
i+mWZb1wUm1TeRbl9uzWlnGy59uxHoOz9KzzEY0DXK9RYc9BPwVaY9KU9W5HeeHY9UHfTckBmYgM
x61ct3DMlztdZbfrN0miuApvp2QmdmjpqQynyH/41cKZSCAGw+CAxG+GdEufHc+DSJtRHxY4r5Vo
kgBgopOXwMU3B+zUE9vL1XxraE/VF+xn76epGUM2NXTyXZ5eAow2LMRuXzv5GwHlk6xUjxIVpZcF
rg+kBzJsNIHFHEYpFzFaU1w0rnXnftuO3mWEQNwhFPOeGVl+tjKKFhs7HE+xr8/QEdCYfmQFcccl
/zCyTlJHxOWBtIVxaYxWiZCdhfwYZqqIEqZPTnEftWBwbNl4wUsvsL4xyoRFWKbMgBbQ7k54+Ykp
vDTbHEfV1xDxlEpVoG/IrAjyx7lCYKrEUF7e1rsnj6NicokjVpAgMFUl8p4UsLUIdcrQgzymi2O1
wJA0E030qMY4utYC3Gy2l2CzBtB1Pc27T7L2UJWog7h2LHJhRucqC3te56l0rrfQMPLkQrsf1vSe
C12o/tcC9GxXU9TVVvK8CvKfKwEwlUbQAvvu8Rh3hpyTSyBV1uOkUiyHCvGdEBpZ4MbEiGPLkaLx
dQk72iV5Qylj2BVtmd9CrTWPMrMVy29kxrslVYqdADNpKjH/EdePUhvejblNs/JweEjvVJnU4XGY
KwihLhvaGa3pJ0TX6ac2BNKbKG/sAyuz7fdZm6jGI06rx3UPijk8AuuOPzPG3sdMYAdN41j9ZNcW
S0dbBzIQhSrzSU+8uPmX7N7QefTD1ETYmPDYeJ501J06voKByzYMCc/Vf4LBsFpSyz8yQatwB2m0
CvPBHNY9cOWvnFMU8SlWR17WnrfSd+DTtkzoQx1HZc5zqNcCGMWRP8WxaYMyIuAx1RDHtRVdJRHG
820aM6C0bLSLjoW4VcgsZypu5nFU8Fe0Wr2QUV+bqSSshTJxyiChjVdItcITyq1HkRcmQz2WswKP
QaHA0iMl+pkU+VgAxZ/xVjgms1pK3BhQ84lD1BbqLAWpAe2aDYzXUtziSUqtBVGtQVBiPMIkMWcr
klFZVvBdx2BC1iK/NkPlOkC6wgIjIMT/cPzci8HidrEggalEXE1pOIN+TyVaGqLzatqIbJiNpZzX
R7SX5YQijCiIrbtCq2wVi1En8RLACFczPrRUe5oPuuflQuzzVWWk5wexYBUU8qUEGfnxwZbsev/P
bdoKwHHVnzozGLSitdGbtPp1e83d5jXbxZ40LKTzI5tzDnZE6wQ263oimhraSC70w7AgtEWY5iRD
wX1n4t+HLcNa0ZHXzwfnGY9py+LQ3EGVjSXaMartawRnCGSGuFffVFIJm3aWI2sbD846TidFo3r7
Z1S00xfhVydt2ZVlf5D6I9sgOSUel8oIW9DjUlujxJWvmcMUa6RotDh7AL68h7WA1RhC9dy8gSNR
Kex15G1A01lnzdb4yy0XEKXZjyE71Z2yaWHkIeMxgQMolcSmsY8f8WTExrDFXwH1Neks8+BXKg+9
FcVP3Vp73e3V69pB3Tc+vx/c7Lt03SAbenG6v2Vx6Bl6aEsFrLMLeovQLgAL9z8a4GNlaO7ykBEv
2fqF9ugiURJAi2JLToNjxRf3fGHU6B7l+b4yHKZw3t9HgdvH1rdE+OgYq2AehG2J2b/R1QvnuN5F
6klKiycPmrpZ17cJkBPsxISEnciTeqgmw7nxmJPKxlJjODzQuLdb8VRtw+lxfvIzwEgybE2/nn7i
wLTGgml3/j9JexPwAB7ySk8yhVk1y08CpXIHUiDv+sBXha8b01/+/7b2aXHxpyncz4mNeUiCg/S6
sMaka/evE1RtBFOUebVzJSSwTLDSgwkPDQYUeFfcY/g2MDEEEVyAfi3sRiApfYR67AYvWWWU0Fl5
xk3wmAjWo1eT2jI7b6AxDIlXNCdPMF+Gb2y7+klILHX6zYqFUd9lSeaXKPncvsa8cdo7Rv/j80Yz
Tcv26kb0m/nHB1gq+WxB2nj+4rPhfDQSl7vRBDAMLgfnpmozcauhqEiBL5Wgn3v1hxz8eWBKp88Z
x2HcdgB26VHjkPgE1FYrqk3gB5yeA29zM82BOZ14XfuYDb+81smUbP6kIatr8GxT+rohzpoi2C2e
WCI7mdek39kf/4iq65BUGe140zuAG4fTeMkAY6xGADuvmnQWTEy/e8H3pjwu0M1uBxeuvFG/v63e
BXXs9DKQ22k1v6LT3/r9Ba/Z5a+YQPxQs5b+VPTE6ggW8djj5a3YERnHr+5ctoFPX9hPGQfap5iH
VeREy0EcKArPCYikXnWjMXjqy+oULwIH+GsVzXwgR0ozWjSiyeUuNBl9150X1jLpE/cyKXqKobEd
aWvcBweoIQuycRKcsMUhJZfAp6bhGqvBpgt5i9QSbum2NZWx+EK2oArMhnHxF3lSlgp4imCbSdTS
cYQ2AZd4WxRprNsP5aW7q3UPc6smZPisRn0ABRNmFbe/ZBf6CUUQhrqmUgZXkEOJWrJeJFzGAfmm
e+FdP9LM+VAAxagSYse8cpjDLP3nzJrmqLR2jC3RItdS13qy9ng0hyQM0R5A10klfq8xVCSG6U28
Tl50L9Mab+0FZ+235kE5aGXcZEzPrFb54XAWxQl3WQ9WrtGAosaeSeeueBwfLMomlIagkTeX/5s8
vgBHYCmXmKKpJjpDEhBXFIL+ZXslNlD42I5mXw5D3ihA/MV47aQAW/W8QYu4J4waaZaCP3ELZxB0
znln0IXxPKLUZ2EnnKfDbHnhBz+hogtFT32DX62xNmDHiY2Y+itvsXjsMJusjvNTFlVbSHpEJlpr
udazEteZ+AErw7frbP50rVXkGIb6JHnbztpIpLiRkiNwshketsJPauE0unKJCmLh+Sk8wHltgd3V
KeK7PEes20LGHDIt3DWmHaMyd91GOWCWyRGq5dIxaL+hvn5TITJH2SHXalHteXhybn9NvBl8iOOX
nxkIRstEtMx+kUxT+ZA6Nvz8H04PitdHBM3CmXHH7T4w+G1L67XhZrA8bN5j5oSWSEpZorm2riK8
emQODr2rHffH82rguJMfJiJ5QrVla1LooOMkMvEjD3fbo1y/PLA54YNHD9Dp6112+xG15dmr6DHX
Erb+A+AiRpYDznInY//2kcfAQZAbI6+QCNrK5E/SUmD9nMlZVV7gYPPprm5MBFfMxVPBPxo464Tq
KiNHk4q4d843ZZdAGoUa2557doaPe2FnwwYfJdMq1SqWAFsKadBIoqfU74jZuRzHIaiXlEI7SVs/
nbytT4+25AHQ13o2VMTfV33ayQZPZSvMr3Y+mj+xm+iJwzfkoxX2J7kRocCEluXgODAYAQ7lbx+P
d5tMJKzHf6zV7uMIG6/fX4aUottMW98mHeBVGY4eSedMH0V7E0N6PjIJOhC/RewkOEsDhRnzIjQy
wl2c8yKktKGKdrrUKFir7Gdg1DHPBZnXvAub/jShMWIIZrIGaPVFxTB5qiLs2BbLjA2I8VsbWjVj
/xLz63JtVIFKB3CThB+LVcTb4K8jxpqfXlnCluFWkXExJi9WhuU/ucH/DKjFbrBXWP+y/r2JKT+1
Am1Nu1b8T7/d3EqNXn51Tw+BUyzFtjZFCGG8Cwgic3JQIsO8vXxf6mcnwwCgzRMSys9Ehn9dyY20
gpOyrK5+FV4GmkbsujvF3U0MlrDs9TU/XuDpLIItqPI8WNjTIdNNdVzEdrkMa5TflSHhPEtbwUlk
j67KyNaqnh7nyqv/djgHj8o5diDLSMejhzyMT1sBZZbcNIRCD9choQnfnoFQxbiiAz90DLPm8Lac
RDrYoSfHkBvhWQBq21zIMEft4ISfcZl9KOacF1bEmNx+KSBGNNL8fyXaqP+AE8R/r6nPeUMKvY5L
it1OpAoKoYOtisOtWsYnO8Ip0T8afoS4bJacf51O4Kacrf9Mu7UYUMOAYFjWHnXq3y1dotdq1lPr
iTEsS2SsKtNdA3WGqOENL7RLG9ua3OWtoAWR1gt5bK+8qAWFgt0U2FBMT0vdFo0ReEI/6yLWax/E
9dLk6knrxV9OKZDyEa+M0vi3xOJ1MXCm64pK0h3RU+SbAcyP5pMCsJOh7n66+wUhWVu4P+L8RM5U
QBsGJzw8bSidntBBQWLvI5XnQsM3Jyd/ULWgS99eAUmUv4J2q1YTBpp33Q+RyVnfj/L0xtQ+nYdg
NHf2xu4XC+hDLTsv538zmjzxsrKS4h9towp0nJauLgPHP2Y02xmiotIIH7lPY2jijJfB9FgLw4/X
e0eddKA3a+IpWZSSBCXHyiUSfUYjm5jhD8zwd0XONXgo3VRBr83TY/PKpL/e2S2gsgut4obsJQNF
XbR1qZ9mrok7ZKhNrE8cI10W7puZbv07MWHdU0VRlAx+OzT9rGXsOcH/LnMio0fy2eIv781LCs97
KQ89zsXsBgJ59lSpiwaJQWXvVJ5z3nD4a/yiorzbsNHjhMnLLGcBK0RVRF9CnRkX1iqP+CHj9/Jz
TpJCO7soatJT71ZKvkvXpXSd9NR+8LhLROmg9UCSEZCDcDYHEYxt0merIELfaEAgCsIeyR97bWwO
ewHKqLNpKKO/21Lzzm4mvI1jOs0Rd/uN6ve6VOoAIg+8tClOWnRuv0W4YVmcQkR+7rcE4vxtd049
MzviWYNTV95Ul6BCZKRdQ8BR2cpyCZICaTRHKyuF76wXQ3ggQGNrW9tdDyIo4e5IzvSR9msMCc0e
EIfPmzTb9e9Gtb1wZHCmIn1AgttlwsB7uumDXorlNNvmQ3m+HpnXwz6dbv9DOtXibSpllg8Un7gr
Gmlvg67r7C7ksIF+WBRFBqB3UiXZ1778HcTDX6XcLa36nnBbzn7XTws1TZR729js/qDn0MVSVy/K
Ic+qp2oOiTEOWqnbYktor9cO1VQRHKnhYoNvRtM6PcMxwNgBw33PdxJU37QFmOw7r7DL74/piKF8
ahdTu9wxfLNIUcipNEPAa8EDB78BKpL94WTiQI2JTM1bq4MR7Z4JSn5A+8LhJpxRmH6mFxxKhlq/
mYuYgWWH8HxohSXUZtCw/cZkB1LPJrw12IPW4n7gKH6o43dKBctKRXgF95cLBNLbbs8ayqPrmLcS
t3/vuoexAjAZi33Y1gK1jpmDk4+qhY+DV7q3wMaj87Ae4J4XG09qKuFMXeIcgw2D7hql9KlTgJ6W
Ide1o+/gYFKbS7xjV6jcBZmVvhoePRah1GSEEQZi/Y6a/P6dIWnD5G/OKdbm3AlnH8jtgh9mIKTI
uZx8vjpHkVXdKIjmEbuZbla8BDNl3gqcH9tqO/lEXhAIjVpKn2be+EymrBvcE5gnszIVPpUgbzLm
1v6rQKh1svB7cCbUFMFO2tUU0gYGMBHfbMMvPBjtlruB202ZyS1w2X71frP0Lhwj8wMNtn/eQTZh
Fb2dAxSDQxdO3pEkqE8H+kV6l84gp+eWNkDfFu63zki676F+FosS5G9OIHqzbyL0TAojwFZRjSdi
I4vT7lSek800d+P4URp0kAIp2c9Adm6PMqlQlfvzCxMN9/7gb6NZxBrIoqUm+ZvDYXb2NGreRgxM
OGWSlyecXTIhMZbTiD4XO28uGVrR6+3ekq9JIcc6HEcOCXYIRtqnw8DhNZzYY0B1Oemdtdj5kI/+
KUvu/KT7Udvjf8ChstxShzKgqphbSse+FZgN3FdnN9wJrdGbv5OgcoyKwRbTuPFOeSlYZlfUnb0b
RUV++r6tc9DhJqIRKajlXC9q/UM4R4i7ixs9Eqe6v3MFBmo2Ke5XQhwknltwFAhv+d4azsj1IOas
NkEtuH4LK1wB++ZgbucIsS6d+1Ud0fuk+077NT5xr4nfMUanf/Y27OHNqIY6P3YxTiOl8VfdZHEB
K1LStFdGvwy49AjKVLKz3A32E1BHqpRYd9ll3jJV7A5jgyjmZqORU4DdgcvoIwXThD2sBOfYS6D+
g/Znah5s+ni5/qku0PdsfXmP5Xx4kzLyVM2aOnsPDwgbuC/kM0aOfTkN6h/P6oNl5T0xLtPHoxNj
lwuQfgsOOnQRMZ5Cx9ngCLARB/9wKIV/RAS09PJjM+Pd8iZDeJ0Tohn6vrZ2yszlYH+uWrw6M02j
UYL6saWvT24pRHys6kXsHuaMfwS24gsZBSLeWfx/dfyW+QgCESkuq6mOkzpzt5PIJN6SjsT42tTz
JfVaozleXX1ma7mJtKYSH/CIklGfkPGemI1lC5aiFKe5i3p/m/7P9Drq116xjSUFciXuQ7NE7kfx
P5s6aT1llbw8wwEsrL9mF68wS0OlKtMIfVXvJL7rO2GbpSYUq2TOtEV8hjhV1ptFWhaJ2BpdENBw
6QdO7ANpcNGBOgBMvPu4TB+Pcx45JZiql67j320OI4sDN5IWgID5gJGhnM9sjejHQTZE2QzDMt4d
cZdnwORDxPtnw55gyfpf34NC0y6qJ/jsymGRMbNdyZl8602k5355lX9tnrdUn7Tme0Ncs0s9+bKd
qQd9BiYKPL8yFVj7ykzPnk3NCks6O8RTiAOTUbgrx7d+T4xUttGZL6yrzA4Ew7tOSFbAzUb8lwQI
Pt3PtOzs/ObDaY/MPLHC0EWTZkX/SL6HbLYL7oubzXM30v5g5GoarO5GTO3j+6g4MmyuzOTA0QGl
4y+fDad2UuQHiquIf1lUZ9wdrrDM7XeX+YeXllya7SS6q/0MHJeGS5aTAEg6ikJxbBxJ6DepRYVM
IV22jG+ICBrQVeJNucfrnvN3vjDCLrGrrphrq24U0UG2t0mmZb+xALMrbcT9dI2mdLSdYNbp0mTp
zGgkVW3JB76bfHQ9wvINhqu3mFBrGzoPOKvYKnK0icqmsCcKrlgQzvgmXIR3nbOY2IT5hXKuNkkS
FBWa8ESLYhcYr2E8RIogvPznbLHAf66pGP7HVlCA0BKe8WYwpBRHPMDK23SPjwlLqK+7PDBEmIWv
SIQ8lU16FuO2qspFkiN/J39a9vDP1RsK9eoGUvYjBGxZXrS2BwqVXzwPrE1mGoHhQEr0XzM7VEWq
COeSuzBmpKSNO1st3cbC3jdd+SgQANjE3EauqF0dAjsG5uDH2HGVqPGTlRa4Cz8owODy5cCF6E2j
XdEG//v9fYNowjig3X+W3VDgN/fGgZI0XaKTKy5k2Cqar3LO62zc5O6UfS7QE+bougNoEfRJhMqx
WJeX+Q5v2GGpXj4vlXx8m2fZbbvlktzRfT4V3wYs5w+knh+G3sftlM8wWVuThtHySWE11QH3LBaw
4LwgzBNtmvY4yM+4O4OD/MLLjFvJmq84+n2yb6F+5eNQij9kTXLAMdvOxN9vhINWS3OyyNDNgpl9
imQJ3KVLfD5FH8W4Hbf9mvHkcVyIM98gsmUiUXcDahvv+VAFXi+RYC8c/IQznZmiB9nB2H1ZKr2n
t1m908t85SUgdRoQiONUCdttvrfz40KI7hMI6MbEe7hd99KIjRUCJQYpx9jkpU8qH0MEFoHR48rc
/GljlafBMMF+bfVWy4kF0gWVg2Z3LZoA4eckvfx5rqSrfdByjNI6NAdmaSUv+zwzDYvAs+p+pUnn
gB/ojFbhRqTszuVdN7nIVwW3rExi6cCCp/KItMT/1VWi35x8SQs756p4RSSTyzZSQWPHc4SNXtDy
YygPYzAptskxlehs6860p8dfm3K8roioFuZij+QNiYZhlwxIoo/4AJfmM/P/ylj7nQh/Mei1qV87
sWLcMBh66m9c6YR4W6U2aqDmPzDQ6BjXkHuO7VAe7a25lytiNu5IOACwG2hddWw5POzQVe+DMGfj
GFLV6vYP9rXOaKrnOFDjDEcRy6QLUPZJNPCjDBlwiYQRJEQN8NRsLlOAkojFpuQqnYLUoUeZfEeY
boWpZfPbS37Sel4DrqVcd7nDG9HddrrbrpclCihMDBbHOYS8itzw8EAmlQsDN9apsGjLEPbzvcPh
WdiENPTAiJgjS971pAfm1rv57+7yL0hAu4ZK/ELOpKE4qx1k/MwDO49lEVchTp+nZah6W5FFOUaU
Rjy/Q7nEQmdZAg8f40W7eHomeGO19Aw+pvJcGGJlY3VAexNCfi6XykfjTxXQYR0IZHeP6Jay5pjU
IikUZGPvQn2IKJwtG81Svk4goZFtK4CCxL57nNZ8xMwsWkdaPYus72wKHK5gI3afrgxdlcp+ns9s
4ZY70iS8tJpLmBFo0CJToMbq1XATUCjmZ6YfkGisVH0E7+Bc3Lj57BaoyxzVJW2JZYhpRTf5GG2k
UigyuPzYnXFHtnDROOgL2IzN5Fs6TUqB7tuTcBz5xSv013xnSs8yyscT+2TXDkYKYfUe3dRlRH9X
4WW/eyPo5SL6KBGWXtfujT+4q2u0p/UasER31LM9pQJaAZLu4k9zdSLYlvT1JZ9QstD8NmmsOM+M
aIwchfJxbXdCHbOy1Yt73GIJkN6WRE7+25my6TXg7fQXYATx2sdKnMIa3UmRlN2aaB0pKvlG6w8p
I/OLs1MrckhqCuMTtT1O3bcFVOckxFnowOGwn9aOUlD4ykWryMqGLxTb0Ai4IibICrEChAObP2PU
K2sE5bai+p7Yp5PxaTbxWASVTO55UnUi0NeP3GT/UuThzlIdL7kozWj6dDwN1zkesIsY6N9+Cwvz
InvyZGnUzmOnZGT0oFA5LsWKjQKWp6N9seDfwvfF1McNBR1qDHy4a3nZtsfoa16E6rosp0q3WoND
ekLELOEBvp8aSR1GrTvpxZrrzfk/AzsM4KE+hWmL8N2cAouLp/EpQR2bHY84KzAzJt0iOOk8wbJG
U0i7oNtQCd9sFf17AFk4v4+VLQNTPKB5ae5JaWmJD21OespvvOjsU5YeRDarDIrnKTRUN1gLuciV
UIIfEpflQ9Lf0SS6Ii0ENCctBXFOJph0oBHXsWI4b9xzp+4UlpgRZ9GTZSLaILUj/T3UAR70cFDZ
6reYgDCstcFBQciZla7dqkID9emR5vm8dSlq0qWguLgTlQbiKkMXuzYAb+2D3VJmHwNII8DmXshb
cpRGvhm3tfmq+ffFIhOtuTD5a7kZxLVvDD+nE4U2qgUeqxSe8uU5oJltfaJ0R6LAkhWDUuklycL+
DBhRxUnouF8OM2t1I23VYUZ0JG/Rh6k6hisKNOy8ktNbT4VzviEOYdbewSbTUvTlDvZIAYRfvdVe
l1oGhWpoOVU+EVFEMLBDVCdBqFilWpQQzx/BIpr7KW4Si2T/fwwXej3wykMMXhlRnQerFuvJSBR1
/WXHha+52d1Nqu1lSp/qGZRaIQ/b67UpjpDcPPooehihvyrQvGg8kt9WMaW5jKbCdBtIQ5pkwVUA
BItJMhSzf5lVHVhgGXi2MFEapaq/pR/Ba7h1am6zveZA/VHXzYvWphU6s7/wC/99Q9SWW1JSQ5Y0
Ub7ODVSkCOxXQFFIl815kt60t/lJpUyo5aq4aN8AcBb+6jCQUIredMK9t2BsDM/Zh3xpM4CDQiuQ
Klv3xTPQmXn7g3DSEc3mDCAxKcuQrXiQjt/KDkbkvCx2vD3vTlNEArPQQkHeXwoct1lbffu7IxBp
sLJNWDa9EFXZ+KSCvzcWhPbLeY+kVlDd6N7f2VtDn1WQzIE+At/d46mIfCehAVPxYCE3xJWzWNJ9
sISEtT5uVol5QV27ip8eo47xUZooGDr99s6hyP0isN5wVVOfTBPfSdrfdhMA40XVcCf/c+GItQB9
woWkRrBO44gQ4IvYVE+NR5dDKBJ9+wP5qLtBrDJWuTcKp4GqRPsMXJOQ+Y0kCGdlw+7t8ukF6h2y
gnn04dewW6D8ZePY2gG5JIRo5STlBqGthPj2ONBUCnSq7+ePz+ry5KByYr55W/tW46m9vgDVKJ+X
lp18tI34vjXVvwskwTP8pwWqBheJZfBdv1dlfc09Q72It2fcpdVA2H1b2MxLN1Y3Sdn5YEbnE5ja
A/4AdMcI74NyERlc8sI0w6IMcae8yAWRNsofQitCedn1RKPEENpYzQuxe+78D/dfXF+sN1zmiDq9
LV4W+JqN52qqjurujGKRmP5w4YM5rcp51oOFtZMUA1nca4B3tdya2/1EY5d5OG0HNDvHWGTJqMV6
8M/tDUrrAf73TOUiIm/iGreNETnNobVXWSdUYIsJ23u3hmHAqM2qYH4C65KLCqzjpypf5ZvNBV+B
zHupUgNipn3diOEdmNMqZ7bjkSd4nvRgGZj6NndTMQEGzXlve+9qmtiwfUPXsJ385BkajI9d8yZ0
p7Tg2GT6hKEQr+x3uOAkkNEvEauGxRYTzJxkHRNbZl1Ftgvr9jeEggoBS7W6Vn4Q46KXODsCWwZ3
mUEINjJY/DOGeWo7naY7f7AgXViNq+JQa8mmydQFvAnxaD90C9nXdE/Z46BXjyVGplj0Zv1LsHsD
Zreop/dhbI8VOgwwnZWIPUSyljltdBk3i3RfA7PnINuCCRmNZG4O0lyDK/yuhFgE9a2WvQepT/KF
34zSsswZAUERMJzpKy+kJNIkV0/mbf5YFdLZAbRxKv7SYRNaSAAAXujTcihPTQ+ANbowQruU1mpT
ekouHLghDXRu+qwoQ0rZ7lsIc8HCenSSMF3x40SCUJbQuCQjAliaB5ZvBYOiar7WVN5F1lXYLNyj
5us4UX6/5sjHZFZNEgfSQ+2mgmv8mS4zPg6DvsHSyBZqstlMXZPVH+AYge30yzWIJaNHznYWtrDp
/Q/j0IxZb1vZeJ+2eYDkfWpbIPWME4yGdlmAIn6g6jKcoX6ooV1zLMtGB84TWbdg9HRpoh/kxNlx
1QePF5LnNdO0zpqRugDrvEz6OJCUB45Y9zfB7Jug18NHUSGCKSvuL3EDphtyBdd2ryg38xhicFpL
rXoXAWpAz08w3JwQlKIbh2J/pNsZhU8jmJn+TMsdUOH0Us6igGvxON2ESVXPKkjSjpASYnxptNk7
EIIYn6J4BvL0CyH6tSIGJebgnZyHL/cuVUUE5gz7HveaBgZZdv/gzmk4vNVDLMsfOi3MmnnZxHHe
3F12WPzsmNqytjOzU6X7x4TECrLODVgetZK7IHNVekVcUMkmdI+fAbmMZfGDD5mmD8rBoIWUi4mc
StaovRBB0ME3PzxVuXZla1lMK18PIHrlF7e64fnH+u9/QgHEE1czwCg3Wi1fVpGMRbdapIPSOgVV
8JdhGnnrZNGUSLGe5s9VhgfN9GObNwdZB6SQU4XESRkrEiLMuUlyBPO/OX1uJYXwXACw0VgY+6gD
10ZqmTlueGQ1gPnWI5xPwUa/PXuw8zfQZ4A9gn/wjBvzx1Q/9p4MnfDtXMkunryL+IP/ci47UMOI
jurjY1iAycLSJV7xKA3CUO5BNonsthiXkn9EkrG+0zVMWBgCGRmv0BTB1A5Ei380lhROv+NhUT0/
LI1wEKaH43U3rOOleK2ySKQaGJauM2o+d04CgkiMGKlef+PhyowCcOrb3sj/mC0afatRz9z+TJ+k
V3QwgiUoBd0yaofz8gZhMKkwhjrRwF2k4PdfK51EScSYgZcPtifqRVK/qmNJu0RFCnGvaxej/J5i
wm+XVmAwFRqvp68i95V8yWdbQoQUDHoRKESgx41bXB1tvbjt38VUXopFlRJutxh+MDFHUttkNQqX
56/beCTPNU1Wd2iQLtbGgA7HxZ3JNfdBpq/SIepzEZGcbx0C17pATyYVcM8gbJMT4ooOLY4nYtp7
Yg+ttkToGmV+jgqhSdPRYkNpEBUOtBoLp8xtFEWBZnRtMV6CyFZff1SFKFN3gZ2GYv+LZsSaLrv5
VDdS5XU2Cli5FnyYWeXlLNAmvp8Th/q2isTQud4PSuY7ndsB9vkRHlf5xh/b5EF5p1HT+Iqlo7mj
d4Qxf1HHihz0AYaU81EqaKKg6UpPo7ebUlEm1VN+3qpNS7m+DWnFlU5bVJZa7ukfsfhvdOQRpyBd
mPrK93z+vDOx1LFVJ7qcBmaGrdKp1vHpc1r87ZyYLhfTRCqQ68OUQ3mHxaCBfsYQ+arXdsupfix+
c5nrV4N1CfNxJlgkeOFVDhS22EqfDUcuK8ivKgU/ukphS3o2n7In3JnB2DHx6kotlPCRmrsvl/fK
FPcBzKKaJWawAIpbznlFYgBPIkD789vxkTHExhyCNHlBNLaEqoBxdE0BjXHDtcNfenrL1LGEYZ0i
2ZTtas42KVUhsOIZUBRFL1UHOsyw0NuqkG2dkis0OfpAcnO7lGpQ8lOGjWiHtWNCd9CfaT3fyMXH
EgbEjJRG2ErVhve7bi4ZWr5DaG0WmcgvfIWjlZgAUM0HmquKfJ7phzJFDlG4pTQqru3HO5bKh6o0
wTSiqQgvOVOz05OwEIE8LFYvG/NZKAgxACKyl7c+jwhLzE1mbTAAZQh9hSit3JtPdc5QCdaCaxdV
4VvQjeKQJnXzUj+furBcjDlgibJgZAHzjndHrVLB+GoUt/VmjAObkYv6crVq5xKR0UjNl9nT7pNC
L1fiFC6LpGwjkMG5ube+pqS2x6bjX46Immugx5X3YfiHWkN2m8eE1BVvyiknSjamJ9ppYK8UPct+
o6oWzfL/NRXEvB5L/6ccxNApdOg7TZBcw5SUwt067wjDzZLcdEY0X5GL0qCmzSh44OxgJLZoBcvg
T2RQcwlAUlNoEdP29CpSoYzdXX8w0ted4IEZ9FdV6FkOcLH8x5XjEpGoRcbRYkfNxepgiLoUbMiU
n/MCI+MlUozWSzfA/QegHrCayH2mUL2+CTFtCK8/CVvE+LcAq3cqaaCYQT//25gc/HPQ0ElBkJEm
DSBoS4oJ2FwS1A5iNcd9QZfS9xvA9CvdssVTfcs6nd8xknhF0xr5B1/wZFBjyE41jJbc54NoyxAw
ZFoVjRHNjnTRvYpSW/U648yAYxIbSMdD9MkD2+UNA914fulpNW67xMU33nRgKp0TfeaD0RVLgwN1
HoC+7QlaQ5h0xRkVq/DF5Sa5+b+bN9wlnBFJafrVqyyQZFGBIAenUsFOrCZHF8rkkp26Vo0V3kmt
9nzRGC0aX7L0Mf2Pj+0uGdgmGNtNvpwWLDMKHiQTG0sxQOEOLYCkXCe9AqLOW7+B83zsTDES8zhi
i7zKaBDDN55EYRso8xBGVI7lVGhleKVWD7J3Iq+Ez17SDtBhCbB5VlV8Y9zDIlcrJErGBl9iqXeK
9CfuMPEvGbagSEGRnpvgM8sUO7gJJ/a+Jwo91YVu+QZB89zvAdbCIP+An12pXsPPjxVBfMcJELJa
Hi2HdwKw2lzrEEx8rhio2y8H/9mz2Nbpi87kj2XcUmzRriC2A7pb0ZGMCotqm0msEcPLRln7/q/X
vLB+Ki8DJvk9/uPoowI4bA5mqkWWCsrNNiP8cAwZ898RoRXdkCElPTcQiABiF502AcFRm6nYfRo2
jqAsmu1at15hLI+LaWvsGad+KuYcTpp/pTfR8xboXbdKvKlEjoDf1aq/6SCSzc2jQZpMQE2yKnkG
PfxYp7n7F0+WDCh3gMntOua9bly2lozEbyl83HkUh320FHrYpuq0SaUjGkrBpJK0QDZeedLZLWD5
S15wpOn4LbTtDxLXB4z39n2WOueXBImfWOnzDq4sK839QIHmrm2uY4HaF7xcx8t1Rc/eXhNGcsUr
yTEa5x8CfTiNP4VER/aTY4rwRsfr1Co7H04Jt84GvheFvVF++87vw2rF1+vS/1yRxQvftEG3sODM
M9q47qvU1hpPgDW/HEj5QuwZ+WU6gWdZTT5KOXlqcIOh3tWi6Jt/1C+abh7jfwMqeXWmKRIx7P5W
aK7ysRwc36Z4Q59CtJtdZuO8lw5NCv0Zks2SUVHj6+0TYlr5UMxYAiUnS0GOmzZbH61v/Cu4T2Oc
c2uIh9LHznqq1SD3czeWw8b5keBIzljgo5/09fcwo5Sb8yQGEDynIlprWxxgvoQEKSeQ22dJIAo6
IXD2aTkrIOts1oPQUbR6JWHn0VmzaT9h63972vZM069J+5RfmmdTsFt6h4LopxH9PeXn/ee/AWaN
QDayT6oMx/d4lZkURoUvXkeC+Xu611JxZ2jeyVNPbHWU6R1PRMNRCJXSEfEkOyfPl1KsO766v3Kh
KcPiDwDk+N66uo27MjfxpSi9WAf37k6/LxNl1eLjTPHeUEp5qNccDB+z1E7rC539XEiDqsRuXD+E
kou4KVBdOZ8WeWPKc8ig/HSk10DQIQAmUvyU7ZpsAzr8HRQKYn+jgsDOqVFaS4+/xMzQjPWQyD7a
f855agKERJCtih6McFeD1n9wsDngWpBE0jZxujuF5wo9K/Rn/VyNUBitUMOzK2vtN0+5vipmGGtV
JLTLilTygYavHjLp3AMpMQdXVI7m2D9pOIeETDAWoltdozmjwe84DxL8a3LFbW7guuSYVJed+am2
FoquNtfSUMuKzqSQ+GTS+F6u443QmyIvN9xQCsTL9Gl9vT9R6IdXVwuty8/sJHUHgNOgeS9A7oqO
Xi5GybJKhI0BR8vkqED3H0EOJfE5xwtOS/vIjnoj1QrhOFtZ9MLFhxVvi115aTMg05HYU3tl/Nuv
wI6YXk4nFV7o9OzZ3ikdd3DvT/cyNLm6nvkLMhCOVTyJ87zLTekw4gF5xdAJFiM4PBUbQY8t+6Wt
aiudFroE0o60sR3K9321w686ywAGWcShCh0gsWLoMLQzBn+er1Sq6HqpmgReueTSoDlAw0AcEUIJ
G0bm8516bo205ufQovYFxvdgZ4i3T87/Hly29fRX5stvS0z/64VInsU3bpy65VoVhS+xk6zQQZMy
rpHYmFE3p5w0oRYvrognoiKpVWJeZPrTDCqdPcHUKe0o+ua8kDvv450Rrj5rbI3itrE/3VzX/krT
0VSGeNsT57XzH7ctJt9JjXm5oLcghLeoydmbG/mpKZOTPOmGgJk3gXtLA79llMNV//5s6tKOKWFr
ipVjj8i3MLqgjVcj63TM9qYsk034QLXXvnF1Ct1ZBTHpvLXhTdfw6aInrHIIqKj/FgxAJQv11GZG
h4BtpsJFLpVsbfls541ZTKQ9Ru1EN5gAv/+oyezrLIIf9bt/QGOP+xaMwpyIV9lT9gzLrR7LV6x4
797zUr2fJwFy5izklAaC4iUuH4owinDsDuksvjcpM7Y1joTL6/1cQ6uFohcGRf/T4VAEl9MRY2lA
Jr1WA91lxtGXt+UEcDT8IkgO2EZDfavzLszSQQiB13PB4thEJhwqZgjZF8Ba3RCTz/eSaupzlIh7
/IbvqOvcqmAWyRSevFqExqba8gInGeCx86UNaGmz3T9omVH5UuHkcXWBqNXR2vdAYEixqHgVXrGN
a1e7TD/e58KXPbayv+lNHPJmoWISslVezsAxtMnnq6eQi0wtsvgQgqSy4tr9caQH8HxPmDZ1qix2
/yXBr2iomSIzdEwqU1L8F6EvO75mSmY+eg4iAkNnF4kBYzyXHGsqZBmvkTInErL5BxFb0J6PJ01b
1wS67I7WPe6F+0ZKiebgeFYvmEwQqhJBcfEQuwBxfnzzOm+4TK30qL18J2itgtSn976s4wjoJGkw
OHhUE++05fl5YmOoK9S2PDTG++LOX2MgASDHRysProJH1B8e8S/3eUb34YSU5+09Aj4AtkY7Aa5/
iVOVs04Wkumr7+CUgBw5nlR/kWs3aZ0tDkyCusoukU4Kti5FQzti2mjcyO0yW4fkgBYJVelHmFbS
NAO2HtJpILsobHupAejXwPIIH/YMoECJJDnidKGyAb52lKWERIxslHZscKKOHWPr7NFWv6xWq879
5CCBbMYV8ZZevsn7g50X0sXKhwm99HcTBRSoVGNf+lP6CdIw9SPCxJ4CxzcanRv22acohY7GDye0
wP7vs5GRN/W7D6hQL4L8/ys/sr6m9Ojbb58kufyr/TX5QTVGV0mzRMOnyBp34qlQYAlrtJG4fzII
yttu6m7OKYc/VGFlaYmKL/7GQefsCzDwU2aHhhfXXrkzeZVjVvJqovIyoZ178HICayzHOEhjG+/A
2vkyXDO/Dj3jgduHeHJcIaKYlP6STGPRGkO/O2B0Kfi8lC4S/zYZwWXjJGZ+xniDQuJV8pMcFVk7
yQwjdr6Ruxh8RJAUfG0+VPCrRx6wK+gnKbqNkxAE550ec/c6lv8+SUO+1AOfQwQ2Ggcd9RMTtROF
6m1TjlGN75N5yBskhNq/0JrtV01sQX1YHUKvLmPkw73cob2UDlJYGefgqZPqPDWE3W69o63bNMW4
O9bE9i/VOgSbs50CKmGh/cyiiTsRah/9PG9JmN7iUcajo4OP71DrlteqeE95yVo/nGikOqfANgIt
KJ5mqs+72OFzpOpEqL/o2ZgHllWW4LNZUgqhhyPR+RYJZp5zOuis33/tb594KX/JaH8nN+a4J5Q4
93PiDuXOw29y51pHmoWKI2+ChKw6lor/r+mGJQ7odArQhXrNdqaI53/3SPYrX1Mh8b77ccdiFKSv
2KHPd6VlsgZozVmmCnTmWkVB4dbb2BEkZDMywItiPXOX0NXNF/4DL7hyV6deKfbsngYu3lZ1y0QW
HnglEPUc/N4abP1ABCZFL/AGhtfkQzh6bssIBKtlZVorTg2zx9VXJRYZDWYdf1YqYKOK1OfyQ6gS
XwXHIb46McfTU890hSBxV+UjC1Pzyszpe+yocVZ9tx6H5zAGmDc0RX2BY+iTbnRwwJ48J2dqe+5D
zZUNGIdzjslGSmGGBDuXAeXA8ZIM02IEu8ww7zOK+bMXzInfFUFf7IUoyOY9NxbroyVCqJDxBikJ
KcJH34obsW/NaPJWtJVxakxI0BuIyAzPFmvKfpzlPmPaVCf69U+yqEbPi8hYOURYAxpOn0miIMlL
zZxpukpwy85lQzTECEE7pyakH4JpT/QNoHVVu5oQH/ewLwuF64yI2BhI6Ns3aRtM+tZAvXI0OmVJ
3kJm5wqvfDmVrJcCaMDYkh2lx+tK8sYpLZPAaUTFdOL6HZYT9ZG2Czt7nnRYXdacjXP2/798jGaN
wEPoN50xBVlW4OfxtxNe2auak5ouOD7433Vz9oFhcdrM8XP9t1ujHi1TRbM3MHiQ9GkxWs7XytG6
OH0E0qxaUjV9TsEjnTMCO0uWi4PS/x1JRyFeB6lseI4obWG1Fl+PNKPOYmklfw1fGAUem5PXw+Kp
HWU8URDt5FruU00XJGgJi5v3/Ouj9t/MNaE3XfBeteH2Iehr90yr2XDhLM1fkD8sBsYEA2PqoAzS
iDkWd108VzkJA+05mG6PQbStj5Oav3JPO3Kx6xjN8N676CFopBYQK1rdIFnZbQMW4HCRlzkk5Lwq
2j7IJ/5lp3pGhccmn5BV3S9PF8YRfFElFlZKz3wmhL2jmGWsGULNYBIIenuSstC2udqcG3pDFLyP
xDkWXzdidziLN1JBZg8W5icqiCBURUPpRmwwiAFc2jGCjRNgEX/1BrnHOCJZDGzHw5YmzeGXwwjn
nZx4A0fPiYIsbFU5sUspOL3DXNhqJNUIGZTUycEG1Yw8Xwa/zEWuttzsq6/RE+MDW46g1VTiQqZ3
REHsyzS8YRH7OynBruewhkJ0iNJWPDHW4FuPfYiAroTISoT3N/vQAqG/oGU0qOISY7353A8ecFBJ
Vb0jaPOAtCwTkRjbpUYdqL/Yj1OU0ax3DZY64Bj6LprcasZfu2feReyf4mtxnV1AufSx76OfLG6i
gkarfEXeZme92k3tMl+05aZZMp/93Zfeo4TegSDFlVY/uG+JJ2RcOh+lqwQ9ei3KHfpJUQzxl5N/
2Q2kns1WyBZk4t/k7g7mIBlxk8rKPAqqNrOMmmf4kbXvKjK7bUN4O7dVIN8LGZmIm+o1APoBQEZv
BYKpsEAJu46MX8gqHS55Oz+ZcYKdFllOUoaImkbjNVkOsNugTHu6Rs66zRdbXgzPo22/7im0ok/l
8oymhpDeLvokVdYvwkP0bTBe571X7xx0ATpydvfiKlQs7wS+N0FEPcbaDeg9hNEJAtS/9C6M8au1
d9/NeVN2b3ut5NvbL6L5Vo9Wos5Y12DN/38HJv0dEe5cxnHspiwWkoVGeG0N3R3drxupnoW+0iz/
41gUCza/jjNKgvvsZ7I4Z3xk0zFMEeROWJ3/XauN1De1P9AogExKUQhpuEsx3BspXrnlS47ictpy
BMzeuKH69njhAGKmfKCvz+DoSAnAjAihCgXmq/+ysK78OZBNVrijUdTn1fvN2Q96UbXnVvu+tk1S
/srX0viyrafva1EK3rn3o608UvyxTxClv8AOImGquxOdDWVdjS55b2n4JFvVlQp3VElICvIu4uIK
WORH9UOB0JHPA897lEuaUAmMmcQ5FppH2/v16FtRJGEV+y+j0xeatMbsIMOLLX5CyYlN/4YI1ySX
hArM6VsIdflRA+2l/lDXkYCoJax3ZglmmCHhlkvv1vMunu9fhPFWYvVhN+wjxiRKg4DRtZiZu4sg
/FefWayWWBD6XUc4hWJ1yf+2Jtiah/KbhQ==
`protect end_protected
