--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Cg+R3eoMcTkg7Qlk1kXSOIi+TeFAHVFhkhU/jKtMYV4QyQwmvmySoYqkL0+1QtBDkLUPuBfAmMw6
ZZRWZNss5eepWrgg0RGgIoUiXwMFFpWTY8eHi+F6pnME5QogT1iBJJR88AGfhrhZx1sUubNF9w78
PvTGZi1VqzVHwAGzsGbATFX7FfwJcfoTceloE3v5Z8HxqmOO1MdcAGpimQduC1GPUnyadvTL1+dD
eBjO5vVtcXTVJ+iM6Cfv9oPWanVWYvh+de0r45vU7qb8mWbpSthft9DC/v7JO3+6yeHmm5WCl7yg
0JVFaniYMMRB5LlG4SQWkpfR71BHcyu8wfEGNA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="iORn4fyuPVufiIV//DcwaERLv4YjrS9YmbzUqJ8UXvM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
hxdm9LoyQ90jil6IRiU4DuuuywpZDdaHMrktJ3IZn4/SKGY6SPobDJL55kZjndB1fQ042t1FdM3S
cq92qE0+pmCrZTePiREc5i9RyiHa/BHuE6JIkuJ837bW1gG6oqaLawMi9eRNQadfAKn0oCDfXu4K
G4j2EKgyfKC6c8ecda0PFxF5QY82KbxXaAfBd4AAe6C45XpjRh6IBjHcvpLPMo896MetlT0e2fV1
47917n0Us/vD44I5qkIWNIVjPg3Hxxz2JEhB6e6e9FxvJoZbkJRjXNPqEcx3A/HR1jfY7iqt7Y4w
DYrHz1nnYS7RSbFa2T98u1YIQ58ee6Ysq7LGYQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="jiSnrbm4PNLaUMm4qCqB32pcFQuLpKKiUJZ9tlo1/RA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8688)
`protect data_block
adiT/gyOBAMPwxdqfTTMhRKVfLPa19rde2Odi7/0PPSHwKILNtQ6ur0r51jV8CCcy4ch4Xr8ZBsG
p45lP+MQ4dNHRtXmg4kbFuAL23nSVxPpfDfKzC2bvtTm107ZcJSgC0yaFxKgH1AtO5aoyKMuBcC2
4seE3BH3aEW/OlSTJum85Z9XQ+Iy+LVo6SL0AtPHFaomJC+9m0PowfHqlCWeCiO7bqGVOcWQPIc9
GHsxIx2ONBvNUt8oDYKJ9t31r/fGpLSUDnkb1Iy746orsR8GDkObecz9NbwbK3dxhOGrzexdXehY
w/ZuHuitBfIPrfAEuJq57Z+2hGtuNeRPY1GvTwd1eDtOnyQHjiUBYBxZcCVfaW+/ez8r+GFl6A7D
8SagcqGkFII/08VDjBsbSw+SaN7gTWLrVYG531Y7HqboVmOUxb+vdYqpfh+q6/awfRI3iZGWrPtW
h+pB9bDqHJD+i2dGGzewYW1R6Od6GxIoNmyQFUJ9as9yCd3Sq6Y3qz4Tn11IGMTp2Eo8l/2wo+Io
gLBXn30XVNbvN5JnU8YFR6n2xaEH0FWKMvZy0XeYLsdm5/Nl436n8jxOK8RvTy4DaVSJGeHvmYDl
nDt1zO5wIQnPzBWWa19A/ALeyH/vSKIwKjfawPu1E0wRg1sXOBxFSiuxyhGeoRD3fKVEOZTScVA1
E3MgMdzJU99K3pbp3hBWQ+qVaH40k1v2c+vhVFsbW5/SGYK7mAWR2zU9VTKaIlB/AX1Fs79Nbh1l
hoBXLo7u655C3bV3K1oUaB6ZESPiElKkLXG5rHE+JaWnl/FR9YMg2spgcdsdrgehNL6Cgg7ZFdvq
1bl6eP0gNRpM1lj3oK7KY++xyNoKBikHLEi4n3gqKuv8oPoIib1wryMXdtpTP9AxOVk+hSgzBYoZ
CdQqQOvLJG3801Z1BwaP2qw3IJ+jegOcdRQCVxkEOTQTLNHnU7zrwsT5yY5oV2o4vOg4tqmBRetz
RpolhAbzenyjI9wB6MJu4gxP7eO1QmE4BbOSZYFWjXPKhYKSAngjBQ2k/H9I/bQe+7bOyDA7sFE+
0lTmLCW+FkLQoMEGWV+R+Ymua1FmhMT1i1XOH1pXnUnwlB0le7SAthi52OfjlsJhA+nRpey4oFfo
wOQEJw1fhTYwsGw9aIjFMwbF7RkqV1QL8bxsrKybD4x2LWc/5I9fTREETl/uE5VBO/lJWJ3qmtIC
gVAIbbkvBBIlZyoEbYIY3nc/SIrlorYTZmxV8LJ4JbR+fQca8dHmmyIBbw59SsPSbnsNu/mghKsF
bOhPyGc0ktpSDykIEUqL6fSE1nUvHVMqB1QebTb+4WGREeT7yeMcv/Botm+BMsU5TmWQQTo2rzhP
FjW+ZpbDahCU2MQSDFq3Ep+RfnI8paeVx2upAy7Cx0HnExoLOQeb177umqaO6aTXkNdvD7VUjdOm
kzUmEK8kEycdLgF2+O32M1Jh5ZO4suMsf1dLxK8hYU5qlCkNoAGZ321cZ+JdzP12Uog4JIW4m6q3
0+eiP+3hcikmLMMafQN7VzKddra9lOw+WKSFPhqQtiN1GiZawi0tFFi8gCCj0gSg9hRpdkNVmWvh
aZ5FjrcykqocJzhZ+JJNdmEy/GofZuBC5un9sC36l+tHMptDN2sY0m0AaFtrvKPM6om4c+Vu9b2n
MJ3IbmT/OMap6Y9rhJBzvvv/dO4xdE7YA22ExUeRcRWoypfMXRbmhAh5M0Lbl3q6mpjciSkOCZpr
dvab5ENKg3kgjz8NSwJHOF0dVWYv9DGA75eT2XarH0c0Qfk9gQn1J53zWFlBOADa3ZryLkGquTWO
uQv+oY9+7MF5xR6d+W4V9HBtCT2MekQnkBgILj4un2SPNXnF+ZyXcOQro8ywg4tiHi288IGFOqIS
TN2oQTAOHS3Z9Nrt+2BJOe4Twbz/NDFbLmrpaydgmM+czcq0eTbUX6eCQ11muKQXAooWfMRVWPYP
ckNSgcby+cY5t6vIFfJ2XGmm4lDaP6fU4za1OW6iQCQunp8PUKrt3oKAbcSyl6ZfkCRgwtzvY4PF
jvgwZrnGsiZfUBrnfEJpfungKeAkDToq3kz8XWCQPXqZDjWTnvot5ljXI1J7gIpkULfNIHJXlBWA
9n+d/8s37VcxI+vVt5HvK0TcMtWTyVkSpScqTaElvOZ9HnT2iaj2XrZxlhVLNlVrfPbYazhH7awB
hX8zs9FHmjDzgTqsRJ6Xi6r0Uxor00tDIHBtDR3N+i74JlyCtYyL3XuWeyeIHZgXUvJ1PT4FdN3I
xVfUwT1tArPA8leisimGqQM2WyAGz5qtw5Iw2X8gGMgitGhzA7A/Wj2hxlnFOsSoN+BftKG9HYoH
slYQJ+QwtMF3IUi0efJU4Czm4nOKZ0w1HJr95GajFbjaFosdRdDsjahgKpxiIiU5u2FsrMMP40zO
7Ex5i9WSPIY/sH6iWwudHHbDxpKRU5ocS01PcV6FiCFLjnYRu1QOsEZsn4f3pmDh3r3PskOory3b
njRJnzZfQnoByIv+usQx9httBEIIrBctGBig7MBopOWYPw6JaCKCXW1P0qEnkoL4Z3XqgCHqfu1b
Ct5qFI7j0rQnXDGVY7riJQ1/P4xDoBIXcfZwqUN7SjGwGwRp0wdLe+3wg/M6irg/tVerHWe1/uav
1goJy1U/ypNUpd2AQ2rLe8TWxJmJkejmCBCQhlyhi2PS9Y7LbInRg/2oLIK40EWpXBWgP7/EkXR1
LzyEAh/+PtY5QoNYGY0Qcdk2YoOr9cFnsHHVgaFGxFisyeNMFl8FQ6QDbiaaGxp5DbJhKqWCSCmB
pt07L8EPyXW8j1VEptWK/fAGcGlxpYXxAeU/ReqMCoQGWUZ1IUF9gu4dbp3as54isvO0jwwt9nCf
9+Nvi8DxjZfCrWoD4QCM0BVBxtf351xWHNeBs6u5Ogb2ZngnN3Pz/IozUaJslGQwuhjCcf8NVDsB
e4LAlHoIVykcbgzSu4GibEm4w0Hl/9mhnn0LvG3g1g6KohU1N6Cko+bcK99Q70S5Z2LH8v8zgkQa
VSX9WKKVgZaNzetM0KIucVNSgwtj6yjVIkOoaREBPOga1c27E+AnqG9CXxVUxFYJHfh+EKsUpqvm
nV5Ul/5zQ5pvfvDwDKQACwthK0tSTifx4eUhMlmbjejgx3HqKArFUwTrTkFj+/fhze9Czz/3gW29
u3eGM2Vj4pdHe7vya7brHqST7ekE16TsSITCk27OMWEPBu+GFNFbMwh/0yu7gIxjqs2m6bxSnEd0
V6imScy3f9+OBJUOWdI6WhK8Na3VK2eZQHgt1oUQjZxfK3mWn4ni9H4+9Ov1e+9QsPP5nQfO+ky9
UveOdDWrC35wkivYKgEoPPrvJMOL0y5M8BwqxonhmaKe4o8fQ1/fVBxuy4CkLcwPYO8tFY8Jxfjn
Q+Ef5VC8b5KXbecjueaxvD9WxW5pbat/06H+DkWmWvIoWQpmYogaqHkhgtiWm5hnpEjIrS55TH7M
8iezH4XJ3mhNp2qrFBygZywZHjyw6MqQvMm4nH5BxcDkLscIktwB31glai8aD3hZ0OZGBr/7haj2
4uTZRw9xOsgrmHqpyasalmb+mQ61QZLAwrcJytJEYvbCQKV3cpZqnc8GyZ1uekEOiMnQVj9eUQoJ
ORXvcSyxoEphmd+vzB1ZRf4+J3EwJ/j9TFrwBUykBGhiEbOPOqsqU8SikNyWVmXBrCOIr5h20oyG
pQLfH4tg7NcQ/7O3wiuH82COdEdy5ABoql9pfYylmTE+JfBtxWkFVNZGDDxriVblN00aJsxDKDT5
R3LvT0iegnn3x4dgME5PkS9yAs+hw6NlniHaK5e8SI8bAO2jtdJwoCyIaEok4lm/kOrRblmSrjc2
5U0mopczRwjQJkl4fMuvOq/FsslmK4y7BiJQ+0v8FxgfaEZmdsJL/WcX18TiVsx1IDJ+Ho8iULFu
lQPOFFm7t5XG12C4fWKGrajkkGQkwFQns8eKT+N4DOGdrd/HAw5ifBFBy5AvQyKXUWd72QYW+1Xb
lWl6SVf8kecY2U8yk64RrU649NCm+NBOr+YSVGhrJdo/c0PntE8aqa86F+7ZEKepa6dS47OzWNON
outKHaRfCVYx4XhjzagRlXVu0R2tgKAS3yrJHZ+rTJrW81lRx6ZgEn4cQ5JWjuOuROirl8PP6484
MSq4KvkNgFmWpP1uwXSsXJSsXaxozk605N+3fSm8NatGxOd1DhplgGL88dY90Aq7RYazxplwDrDS
kdxpU9OAZgitzNNQL/vcAfgqKglQMuBD0nj2dF9SlfIFdPE57M9ZDQGcEbsAzEe7U9oUejQToEDh
c/md5jCYHpOFD4buRZSHfByedTiAwOtm+FY/j9AnFFNFwjT2Dd7eLcPSdqnP2rScv0QginN5sE/Y
8iwHD+n6LnkT6Vx7jBVYxeRQpi/pmHXEaWak43rugKE56GU87LoSRkZJXj8ckGB7gQlHjhiwbP8g
cxkAV1+XR+MsGw+vKigcUMhuGkN7P154vUXUqd/qciIss1V7fddp8mqXI0tvY5oCNobk3hEY5CSq
z0jVxfGvCCHJqwbSqjBoJeEhEh3vxiVAqO6OI1MdZxQpaAIbZRQMBipgIf2PHFCMTmNSKC+W/AbH
ihQwY042OxziUq8yLto09daguNtWj8K7BQe2jHZn3X/H8+PY0dykL6bqLRDjaLKroa9s08T/i7An
b6LV9hQcQV9fJHcxDdObdYwerjxOafTeIPyCyV1BsbO8Qu/FVK0a0mRVE87/UL0toDlcMvyZtl3w
3XcZGTFXJnzHPEem/Akt5NFFPzMJo3xHjP/LliZSpxBDL4cGLYolAgnumMHoa1VdmZn+N1WTMKFF
Vb0YAIDJWueUOtKFbXNDBIn3Kt8KE7Ft+nolkC5fmO1W1FFBfYY5CWgeR42xPDX47hG/HILK9QjW
7iUJR1b5ih+F3C0SsUtFiu+f9XuOA39r69FBDdkMS/DqzLjxgsRJhoG5uBohrn+VslxO5vPjff3z
CAq9CVBONR5mQeNWElyHraw5cxoJ1puctWi8G/ou1PGcyVhGDzdScFQNwoEbR3FG1Zeo+dyVeIr4
k6Cm1iCxP0moXvCcieRH8o1kjHvYdMLXJqT2jRGIypMgqquaJEpb2In0TXVvf96MRiKOAwFp8GwM
dJqgeT6l0oXnLLnJR9RELKf2E8Ix9xG/ZEkMAYvHRtldQcpYEO82dPWjniIccgCCalx1veXP78La
Sd8PtK4V4cNOY7AF9QUAnHddAa2W4F37MXNahI+Bbf+W8UHXVXNwvtXi2fkNzhM/HJ8jYn4Tx5My
94dhA0nHkHhIU7aqqqEOzJdULfz+jj5Yk+kRyGLam9engChTrObc2XP0GLaycSNfWrDXrOV0qnkB
q3yYVTxoyV+tWJq3QJSWic+yUbgWnaediuKn8zKRuza+6csNWD0sEPvyhCwmnHYumkov4pO6Ubap
zWpOWdhRqcxkXHWZHzu6qG+2jyxHqnT9V00atZgeBqJwxoDS2xzBeiw88VU1vMYQekv75lls1Clg
6r17j4uy3X2cI1bbL5eVuDK2AnPjIviTVIDFlZIqVLg59ig/qGNtX9qD/zu6WeAoZOSLwLMoQBTe
Ws787B3JW2cboj6AAUh2TsaCYtFzZzbnN52GRwBzskkNvFMHVyxTkst50mmg8RM4jqU9+u2BQZQX
ocgwf+yR626vIaf52yo1mxgSzWOC7P9w3fWOCdmhHOhctQkdxxhpZ8s2KOTQLC3fw5quUNS5UWXO
MIpCbQXvNbYOWH+hZ8MKa1j7rQvkEDfuVd8/JDrcnJ1n6IN1GOdxaxCcT8pU/6o84/DIzFhleKpu
2Ac3y3cnV5Oq62LYfylXMN5UVxbQvT514Xah4evSooct0/z5egrS2eBwCZk/p+ByDPX+QbDLYsQB
6dMIWLGXaELlazpwpjDiRyG4gBgByAbagSBP+rbSvLLBN1JszNAw7MEwtUbEpIZKabdjEmxMSFUs
Q3vVI9M04cQbBaL8jke3yA9enRgIzquuxnLstI8n0QEg/7RbpYo8g1NJZko27KXR6Woa6GC/hJWd
q/S5dZphbDnHOO0Iwc4vM1WyDedrcZuCd9YToGeqc8l3FfRxzwqgJKKTlL0/kKgZ5SQQR4N+6c/9
OP9M0UGeAR5t7Qrk4NQvZ137BD3957aMIjymOAl4PJqgsHBPiQma4OU09ISfKhvzafKthuFRYZoM
jTD+wBwv9HqKtN8JFWsDvseVZ2ujrdW7NyO1ht3/saKg2lwObPatbYhUArNGDQyZomzYgw2AD9Mn
byGpsAd42WFM9ty1HiQ8W/pMffDAZmMHNi6DvsYMyKWtfrLNvEaRBSIE3o4AIjCqhyyBfouICcW1
hdU0GfxIWY8LUp27OODv4QvBY/zCfgyLvgHlWO7Y69mbrIJp3JCxrncFREjKTQW72SxrFEESMWcB
Sv9zFQfITGsGYzxyii1NuIAH68joL4niNXYP37jvvjo5QJfj/OuCvqzXqZxALMwNE03q6SAnqGy5
z2+xD78KvHfrZjxe0GMDpYghstqREwbdYhaoN5celQM49iFiUBCWkysBq/V3hlf74EJWGXkwOK6b
1D+j+MgOGuiEg9h0B9CrGEncZBbNChOzhrP9O6Cu4YRvylyKf6MDmzUP6ywOHNuQ5Zw+5SlvlPzw
q945uKRvhg8LPTuxICDtUwey2eSke8xNuyHIIXHBXW6qjC4aH7p3M6TOX86g5hGOPVZOuuODqD5o
QM4VpRXjX8tK22nrKCy116Su4JMU7TrJXdOru0GyVBPB7ocMF0GaMIwk5lTmYX4nZ1qBufP9TBoV
DGmUwnEq8nyVs/qrxEabf+NDk1RSJr89uE1T4a5gjHFu4AiSfwBq6BQf77TYYaciXHEPfhXyEEIw
SjNVojqYzKkCAO/qMeJtz5/xFrIgq33676mFZDInxlS9GWfR9H2krhd6SfdoPdjsDSuEyQ0LNDPF
nVMCKNx4mqHJCKeNaPzEnpfyBlhnYbHK0ls09vgXJi2EXcib6UBgmmP8HZT+68CH8bIYRYgFZQqz
Jv5KtBkzCluEZz7wsuSu7A0S2cVBjAaGFI9FVbPGB5pAngZzqd2PJbD623CriyXtGBBl/71raB6d
yCqaEjd9nvs7DVrmLQR3M8+FjxJ5AODpNexyHt9NDxoHbZJnyM8QYroMYFkG4bLhzn71v8nkTPu/
l6SEL5Tyhof2vCAjqADMwwVNO4R2x2MVYGBxiAOW+5DjI+PmVXxU1KHtoZaBBzBS+SGv8K8LfPWn
DUZC/lzBUh4p8fKv2PTKEcKYXHBc2yWKdorDO8qxBqPT8y3IZ36YynF0zEOHUWwNSjzfZ3IlgFEG
LiC8pKYdgD1Nyu8bxtxufivW+0Gth01IoK3rDrXxvBOubFVV2+9RUhsoYmqKq8IazWS0r3Qrr9jB
SgmqAiqDIxWPO/+dpIyW3WhqPSDjVHrZwzm7QtOlOaDP7JeuZ5aW+wuHG6RzYgoNqrOkLMBE+o1O
dwBkbotqtD3JliHnh0SyOeM37tslmVVBrnDl8MtusHi4JnHiH5ENapL+6VwGpiLvSvkvCZf2PoqC
DBJzv3c8+zbjO02T7nGf8u5Sfvr/u81ZDiTHnXFehNmcL5Hmctt+ymfBVRNOlgC8K1Ml6nSMwIJM
FoJmzXqkkSrDPs6bARu0VmMhQQtdniEVQrr1Gt0YC7tp8uZUemJnxsNcVyssS139Dq1V4JxeQCXs
1S5YM7cvqd2LD9Tq7dRmW1TZ5soH06p5q7oXKn+PGykzRi+eK8YJbiUB23lmQe10e1vp11ukRF9C
qbUidXD9XZSBSNiF5Va9BxLywmeKYdwPlFtuscJi0yXhheoecfQ/FDnzp1DjmPu6fHSRGIEERS+6
OrzS6TLjFbgQqCxzKzHvmgMjkupxtgSZmr/qBsfuqw12XbbcHq44KmpcFb9VMAUxnNx2oaeQLy1/
J2s6uV4eRerHxfUvjUI77gN5i1le1wcGCwTvVndew45zVVfcuodPb3mzPZHB50+MP0em5eMv8vn/
jguwJ2YLsAxjz2zAMXEikFuq3b89pEI+BAWklqT8Ceh1hqpkxhlheR1z5EnLQFRBavE62uMy8cWO
coSrN43452pGrLyOLjgmjHp3F2C1RJqPAQ04X61JLSs8RyuxmQRnjiCeTtfgUhn+lWLanSZBJ00J
TLWrIKh6k2RTb+pF1T4VrDMc/cKNXXiP69vrbmV4DN9bDcZPSkt4LWXwJJIBBwQjZgjiAoVwI4Rr
OY1E/LFFyCwUZ+izBdzbqikyy4BsUDFd7Az3gvd0SfvAJzQxx98CqT0uUG4O6WuNRQaWo3csCWD8
e02gM+MyAUnX2vyoKmDbCpz7qh3XrfsOGwbDSBabWKYOXgRJQnkLqcbLtQT4B8nHQjypvIly/T9m
qJYt9KEDh5h5XOvgnvOFjx+1yRbsfKS9HsWr9Cbg0wylm9HHkoIY6ybRhX5oA6pQBpFTLHIrfdwQ
UQS2Q5KPGJG5IsOMalXA36nkR/96vAybPt5RnxB6iqZbyHwmPfNS/RqW+Gcpi599WQemmJvwmsla
oOvfT14i9KiKTuKc9KX+hh/jE9IzXWRHahlkLLs0KKorZ77d75LHTEDlSRvJVE6+pT8/7u30vTAl
lIF6AWKW79pW9l7qFHNQBN6x5PrfbjRqhHHVGBUBzTyZX/2cWosma+3a/WJ9woq2exckAHhZ9itX
sKNdrGBjuzCFjSlZuF7zCc0YWIjUEiEyWrZIVDvy+bReNEHXObo7at+mCX1xwTfX4gii1g4uW1h5
hH6eFVCPxScsHBmCGqpaYAXgF49Vet05bF+wD7sH8RtBD7nNlLfjgOVOYJX3KkDN9bwB4lrmj/iN
Q+FlYferHeSka/fSrFfixV0yJNNMEC6y/DWJD82Id3egrgcr6AnI6dF6vWgDC+1BXeTz3jFVc6GR
31oKbfLZPyCf/12jmBA+7n8a5SSJTM2fMgSZ7M2pMbw0ZXLV0hSV6Q/5a8942O3jNqjtkzpRe0We
6Ioybp/72iH94M5KArxjLyXZIa/AyuVsw0ypLBW4k1jbifQ6pH+cCkfkZfPcN0tzOM9Sycnbxi/j
B8tbS6YjJYUVgRz63nvu40ZA58qaAWgr06EWARkCiaxe0yFUswny1trxCCORFn7HcwlGKA3DbNLM
NcH6zxnBYLs2DkNahJv8sRHOZPOtJdJGaERKw2IqYyKGuiljJA6XgrjSTqJgodJM7pvYEQjhLE6h
mhh2pWb8xKZv3BfB6An6Ike2gGfvn5NUMYX474trsCMdJa0YoHlynv9puD6/WtcC2+ZnaJJ4YCaI
BA2Nj2EB6FOuqoE+VM1C6C9WW9zLCuwwiYZ2W6W46Sg/FbX398y6GOGy4IhKYPwtOPBLWRu8fdUd
Uj5c9e2zmalwJsf89Z41Cv4K/yDynOvsUP0AJCLsrQsrp4xS+1Cu1h8FAcqbhUUwneoLaDRFUHtO
5NpMyAeXfL49sdpElRY3cPWHdAZ45GsxQoXPaxZ+/X2lAmLMBZ7J9Jq/+c4GweZVfGsLyG7wBsYD
5Lm2SbkK3NjeLH0q3RqvS29p8BJOY3Xug6MsXEmjdXJajYBAhPPp2qilUfiEdiV0rC1ctK0EqlL4
5t6hb7mgEWT3LfUlBPwNZcbVlZ+YT0BS2ehYdXF+9U+tJqBDd/Bpr4KA1IIkL+gUjJUm+tktfLmY
8mswoPmZnzb+4lZl8MBiTfp7vXgDZSMbM8MH6j6BCFnPy8yaH7RTV44tTPU7CT1hXTPFpWKMHLQW
IJb3aRvyP+NEYPv7z5o1sEVen3HuErtsZlWO5dyQ29jPjQNHeRHQ9YQBaEIYmgzH+UPW1ZawYCx4
y75r7W5QLkdXgDuD3Y8WU83PDMyScyGvl2B3nlyXNkXzBjV8mKCFWIudtEuzwSvGdtZ8Pabz0iiz
ttFaY5irFjdYekW4Q36tjosQ+3Lh4wpiTNLXWed/Sd3TKr7XAkHRdGv3FhQTz2qfgOsA1oiyLQWI
ZCwyjxu0vdFv+Z5YZDaaAUDdpykiGM72o8EEJAmphuDjijZf3FEa1QeQUs6eTB1BjZKy2ly9Ekqf
TNBpfCj5/0B3KuQccUkvLbRDanGPEKxqn0ymAM4m8AmOG0mBq1kMPdVnhopQCa6FAWAS+dfQJzPo
WpJImkUTwgvPKW6SwH2bV1MjKiaCRLw49NbRRrgyCHCAHieKPInbgpiA9hF4erAk/IrlM41Vd9tw
EWFWZd9RSX48Of9voLC4LZVVCAh1VnkM8lb9GRmbqCr9FkS8FWKRakCFvHZAjWeIg8OuZe7u7wNF
BBPSnYBZK0YWw6o1rmsWtiATcnvYK3KRNnujVrsb/4scaSfYPZfhJ1zztTKq5B85MwSknvYW4v/I
ep7AAvgq8MVUrh+AT8XnNhhTMorG8GnTQROO+cbVEpYNYHc42zBjFonqR8gHDQmQuC5TtRUQYu0z
g0jn1OuZZ/as2Qajmc5PFDb28t/UXJnp3i9B0Ql5/IXViAf9XiFnfcVCjMAvJf4teaXJidPKc9Xv
UK2qGCyC2wOe06K94AXKymFJQMWTPKLHTbv+iQaXv8U/b9TD2Yl+wcAmkYakpvsdWU0gjegAfJ6Q
OVSXGlFyeCBiRvWx09Oz1DViTe/GuGxtV4yuUBrJwUQINTFBE22BZ9SAbBuQhyq7qK02RnGhWVvQ
gqWiZfjaGESMf9pAZaGStRkFrxhDJdaFiSfCL0ZklSmiIDx+2tN6793p7eLjj8MMv/uvOyI2NDUB
S24jk9beuZwJy8d5bl21voMbgpPDHvyl7TiUXEfX/Z1+m3Q4WqoFaQt52lXG5JMEVE29s1Mcrtug
ijxeix9e0im+mSAsk/+GjmpsrZmCoYGDoxRmr8SvgxF7I5NEvWM6fFjXGVcGVPnkcQjjwxOO8DUR
shT4UmFKj8qZ/yz+sph1Xl5MnPFXIqFs9Tfo6m3kdZEn2afTIQsVg52prleIVqMK4BMPIBVztv/P
dt7ugPaimo+HUEXDCQG4ejbX/4kyU2CsTbVgzRdhZaEBmAypZRbdipwEpjxhCOZZ7yYaAWD8p8r1
AOKhh7ObvQIYkuO3AsUjm2sMKp0bHxHWzDnAHNOu9t+60eXMMiueIfd1lIQC2LyUk6dMSl4Uu6u5
XdcaU4A4FGzMUkuXXvWtXe1A3GFdb8uQCVmhcyv/l54C1qZ6Q2ckBeyYI3pd31LSDt1DcvbdMaZ9
6dsAJt6toTC/r18pZzBuGBfzJJX4q4MOJ/aGS1pG6Ox91lgCRCMo1iAOATK8lVJdl20iCoedLkSg
xRoz/7Nv2jZFP5zq3GsbCqigjXg9QRRwnpf8LoNpEjfdEoybGUvtR3dGPOuAZv7a2uDHHklxMMir
J+wzqP7zuEi6BUPaO0Jqu/zd+J2r6garAY89BWzNYiGTyTbzkYBkYtE2WWy2dnK43tHAdDVLtw5Y
A8bN1LeqqMZSPMW781z7JmSAp5KAQYjgijDoPED3sbcnkO7nywTIvIdjiprJxizT3+qtu5CZpWUu
l8I69QxNzF7HDgND0aY0Gbv9xnvJYxzL
`protect end_protected
