--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Ors20U6N38izaXeka8Oj+wQfm0e1M8MsAP/u7UEOBIr4QZqOMupHol/RZPZgv746zSe03oK2JpMz
zsQM8Wzk7WvHrIGCRLnIoZ62NoD/Jg4imUJ3AX8Vzh+jAqCDAEjMajbREIFAgIqtHgRHPw8TZKyl
p1YUwHMu4EXjvHnfHlQdrh99Ps2YDf2fQfzzQ5X7pf4mKbEhS8b8VN+h3VYSFqoLHbThH5Kvcoly
gyGSxGaNzb/EAkf7lK9MlyWwhJfE6EM9UwSg0+s1s598G+wc3+/1qUAbopyOQOQV5nbZs1A8BvME
0lMUaKMlNBL3isD6pkx307rmTWMl1kFiMgt1Mg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="MVlzZPj8bHVSvZFzMldN+dkNuz4vwKLzt2rMrRDwmP0="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
K/kQbEZJ7m43CalDwM4V9l2Jb/6n4vydXNmhJoj/K4ViviOaOY4WE3dp/aqH9FXmx96yEVeTeG4G
n68sLrqfvL7zb6nhryiV1JwR/4DcXoq9nWC3vtLHrbnWG7FwOdToi/4BSat8kuSmCF8r/ksIZ+71
jSD4MPZe50n4lhOySJ5OSqKFfJVRHglRr2Vdx4Ev6mf2pvYqATHQeuq2ukD632C+FiGVgiovvnE8
HnfqoCR1euwnCBDGi+Z27cLMU4w79bWEovPsgrO9sfm837VqT7mVEsuzbaaI30kuo8wmLVph2sn7
p3QT499A6kdEeTM/afoEiwyWUpBYKpa/f6xYCA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="WFmZO3uqnk//vbDe3jq5UA+gThJbRXLkWKDk3v/tst8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
RpfXrff1ov0C7FK9f1e66DYLKt8rdIf6rgh9Lpjy0aCOroj6cx0aFY+PKdbk2+HCtO6hn1wOb5aq
FOlkPGxCXETIKdpPd8LRoyVK3tLWDNEvt4hWN/F2B6c6N1kP3NmQM5+FLArrVCWy59tmSjrr71nY
Cw7ZqWUnT9BMKbFk4WGNh2Uf1IKu6BcP85ml9r59iTCbp+Fnthoif+TruFEDiljJeNymBP6zP1q6
GFJReUADP4hG3dJ6wEeJ+iGvKT5yLrjodo3jQKlpgf92krWzccjo3HuVrEPMs1MqUWjzrmi+o52w
4fTg3ucBT7p+cMEIbg+mo0N8kOHeS9UfQ73suxn0xu/B4W6r2UTsvjMSzEsP6Ez1WRQUQH/C6vAa
fnI1QkeKT/s+QLEEKEfeB+eOQtyhjuADh09/poIbPY+wWFFHzgrFFF8IcE88p2+l0UndEy/TDWZ1
Z763o+7CBpWW4MAoZ4GugutgM4W8nSf3yHsm2yUP7CJA5eIzw0rrLTcuQiUj/ISk/Vq7jbQpl5Ql
Vqh+1mRojZMNWOeMfitZHMlU3od2NZp9YAhibHDvLn+QeAzBONongRuVOw+D0OK+5EoU5eMTgyQe
rN7H/lAyBs/pMhcAQIV+U3zUYxeTIorZbVbL6QSG/ZvshcjMyTjZrE1lTTiJo0EEAS8U8Aj1Esf9
I7wpNv1FZ7t1IHrWItmNwoT/+Yx/XMMgM6o5jls8zOUl+XyYNOtwaspclMHbUXTKgxl3Z4+bvwgB
tzsNvdy+WdIJDFInqQfWvZz28UmBwUcI5pyagFZ78qpUM/Az9J9fvtyyWJOOb6wgt9b7Sr61ny39
hRb4TyAFTZ4MzxbPqkk82hJKEF2fT95wK/q6cUDZvMTU92Mn3E525a2rx21llOCWzzzPOmwGanQ3
pI3Jbc7Y5aREYXQIAUSSdo0tEKHRGjz8RLDj9r2V+ynKwf2yu+3DbARKHx/0kmHgtRDJOBu5lr+4
C4eGGGWfkWkvd2x0hba+8tn1dK1H3v9WHeUYCHo8cm3a2JoccKadL+qDeEns4BcMSoucnHieKeQp
LTF5k6RZzz9efaBHuFLwPsetao8qH5tNjtn15gIohej6eTJakAwz7snCPtxccffi+6DV+T5g9BVG
8LKfoHG7uaJZn7ngZKmaHJE8L6r/Sc6pKbQW0y/XW1PUNnXg9D7+4fRt79y6wtMy/le/IQjaBcJP
c1iFjGHgYZpDtiR5/NoErRkOTw2Mje8u3lZvvdJ9jtddBzfZNTeOHFkQGix9ZrUORFV4ioO+axVo
NvQ7NvE2Qzi8VO8uHABNIDgqMYzRzUZzZ9wQGQRzFv8MJN0KdVkuawJtuNsOqPrixHz501brwEd0
BMCtfUuVEIG96rU1MIjp9ClUPo8I87CKdjZCmrRxoypgkDBvesKRn73IeGFEmILhyMNu5TU82P1N
Am2npXZPe5bOfymnGh6XRjIRl7yxLvafgn4ogOaEtcvDPXjU56aYamBPurMzR+4v7FC1Ej+kM2QN
TP6duIMrKTk6keEviiPwFuQAiMdFAbEQFrNh51g8em5wW7l+VhwR9+z4q3eihc6KvPupXErDm+a9
I3SyboCTlSSqw33jg817uN0Myga9XgZYCP8PtKCw6cpKuOSss5+Gt+8mTTe2j7E1wmysYCifJPQ/
cjHp+kzYknAzpPVtUgwKCnzUQJ/Y/85Od3F0go77T92UCRXPtrxPVwgk7aTwvNGhUzQG7iixwhVf
9HH5XmFBXnAKIRrWReBEwSrldH0hQtK2/5GlehwqRxZBsMXfOJ32i95Va9K0QF2B/1aXbvZGEDDe
JCfpWUbby4MwyRomsAOhLVXa4Qvd8sxvLx/QSiPX0S1v9vIOKG5uTQZKlYiVTLb5MSE8qUL+j/zX
E4e7TD7EASZ+h8beat+Mwa/xAb9/pOdysN8oeZfChwolreLFUCx3Q9hy6nGru6DrqREIbYNU8eFj
wc5WRGpYalycLJo4y3YWLyuk4yYak/SI3bBBspwyInq7xVrK3pDjyVub1h4MXJInkIBInLZ3ieWk
HclREoehki4oEE+bkqiyaW9HIDvQzkkt5bGOI0JjU5WMjdGC0zHR+5mkWyAjPcErGTYBsneD254X
Mwz4345W2DXB5lzgrp2haISBBSqpNsAbF/zOyVEoqu4KRXCiHbwXqXI3LaPNHyGQapfN9DRJjFMY
yzc89Xe2/No2FLXNNlfmZG6GtKem2f9WAwvJ2Hde06dqOIirKUh9/EuNpMWNDqh+9oecdXnKIpiZ
rrCas4+Mp5Xj/RmZu9JDUVs9JJB8BVd9SBSZrxgZPNWBrrkdflxyIspu159oxHOthIWXfLpvoX5e
eiB8zqO70GeYaamwRSt9rILgV+PZOoT5Vkf3xCilr5xeYZmaZB2dusBGHF08PfmmVecAwc5WTKDQ
L9+mPCm19HVf4Aeme5h/Gvc6bkTyW87UYp25RAHJE12nhuwOKpSGM8l4I+h4aJWpEaoYQMCE431J
TwlZAnvME4KGwE2MmAgQNKlDwBzYLfIx4hA/qVGOURnxUJoEKGMaEiW4fetxq8o/O5/Lmt86Niqo
pPBNxmZuus/jxpFVsV/ZBWZuwNZv8cUZ4rRAqn8oLeH6iRBNbnsrKv8DG6NH8imX44lJWbcqSe7S
9Wddvd3u/2XrECIpoeJF3b42NR+R9TBlrffKfdAdsqbBXTSXQYsGwuD7BjqP5kGfcSshOKXePQg3
YWvxRaN6aTLJJbqUIaDVxgv8/qlwdLZgdTr3X9D0ZljGcQejuKMf4hd86gEwHxLpssyx1oP8DohE
z0xGDbKjagihw10WewlOJ3OJ0GpqtR1C/qwirC9rbL2iF33YjkkiKrrIkO8Ui4UcSxF6CYD0oVVY
tt+OndPUyvS8HbmS/eeOpdI6mHqtOoJB7gC40N4jZwO3V9oyoXtsOvc1QTi3fX1SbNJXBKN75Hrr
jdl3ppHe6+9fofmn9bdoahbogif0lCY5GSxV81IrdF+crMgGpBEEfRRm59wej6xR+D9GVDBD/bjq
HRDNoUo/rE6iICoCD16yMJI53oATgIi61dYxzr6hlawKyJz3raHcHDkettEbxE1e06lQpBdRXE2e
sgODeQMXl/rRoD4PoPtweWIbNIG0lXQCylYs8t2gZ2zaLjbX2pROWP9Io4CxtysoLUQWMg38opjZ
YpBcLQcOyA2L5yeZDUwMfNpXAjn7daDsTVt+C0tIl9nkketyXzqDPuv4/BCBJPwI+/L8VJ/UmcF2
8AA1oBLv0cAmy8RsY1xbrcSJFPfyO9ClF5JojkepFZ/eF37l/toT6XsRV7lQsXJAPsJNveR48//q
kIBYs/AGEuNyKzQYY7PY09kSeQYGuY6cA0769cLdPIWhZygJE682EQhtSAfihJjqKT75xPZxgYfI
bE1qcTpyreDLYqQa2/Anukw66uCem0OtNxONdafIuZ4HbG0SURSJAWp2lGGC3nJFnTPsA/8H6yWI
S7gcJ/GdGA9qtfSqsVDDLAc/Wes4H9O/eug60ZnL7zIL0XWdcS0vH7QUeukmzaWRMVsqXnZp3Wzg
PuPUw6QfaxVp94Mkt8GgrcmJ5WfKpdWZJfHPgf0Q7+PkD4Fa/Fs7ecpVCGtg9pQpjOdXy7oR6XpR
MtpFOMXr3gvoxugJtja5Tt+IiQUwo7qjpjpluL+mAVm8yS4XEsqpDNWJlcvCK0pJcDVg9w0+kiyw
4lylXNlGGO5s7m+dpCU/Rz5eAyozbE07HbOOKkc/eYvi0XX5KHvzsLIvie6Ka8l+q3pj0TIL4WoC
XR9y4qkdiKdYjPJLSVYcvyJA0CFXPssmXt8eypK+Z5CsRrNHRNJCQYYLU/h4C6yTH1Hgdt9fRYDz
LgN6qs9lqlYlaiwqMUYiYlhes9R3ztuDI/x9ZeRAqWD9f+Vq+9pj1whjFjNyHWaTYDNT4g0FUe79
ASAslymCyT7fWpny9EB/DXaoROy+oQSWN9l7tS93nPU0zhF+S6RWEDHacsJik/34EE6HvFx0W49H
IZb1bKtPcnat+FP+jPOCHTkaGy+hFqd9YAef5lX9wuIWUpGJwA4Kt2c8xmQk4vsei0VbajqXIn3D
ZY5ZQf+PTJuEjEv3CmHwTrEbksy4B2HtwOSF0aCrct9VbI/qHGXcGmW/V3q+ooLQuA8FxElMEW+V
ifHxgzPngltcZ81km0GJJS1s5DhKrtHmJk+uG6yp4sUcci0ZFBU1Dzaz62NRaBDzhN9Ub5lsehLY
JzKD9z5U8CxHpp+YaLihZrvXdotBa8GTnKZJkS40e9ngmLW9Oy3HVyUb0/Lg/MRCqAhoMtLzTItp
F4J2Xmqz3xBA9/1pBOy5DzzB0MmYYeov91jGW+h8EpN7BpmJwMwnBSbzXFFV6AbbmWagYzqkiPv/
MrMNWqX3fo8jqOolXtMX3rst7gW+/YGF4qJYyyePkmgjyseuqjXYKdDClhiCmK8aSxNbXjZWn32E
I0B1PDMTlqvWJlwGZgOW50hGpkBZNj7YJcjQPhTLROMRSCv5VTtRi3ebOJbuRgNpnW7Nf+xJHoRr
o7Dv/zxRDBCOKnGbG/8uddXYxpdI/jvdRVg0lM416WqaCi+/1kD3DLl90sgFmrPrALP5T+bbxuaD
PrUKLvKiuG7/vA5rCmilAXN0ryx1yBrkdpTkDtd7Cg6Hk0D/MAx+f9MSaxFmVHB/2I9Li7NHHTSB
rsfpO0G6SDu4TsNnJ8e/XRWe1SK96qPgiC9y+A4HuRJfjLRIl5yfWbpoaUbLD+cDxHZgve84Rjni
41ogXNKTYjqsC483KWmK2ybMw8dQkIxvG9hEucWQ988syNUO4p+IdBWDR9ACvdUrfEDfXofNEb3u
aYApC6aLhLCELon/d32HJUq5HE+QVDCmuekaA3+avnkzpqEkr1oRmB1K4k4X9CskBzZh2udzkGBR
G/brhE2og3ErjjIc60/RaUnA3XzE8dIaqKuIRVW9Rm2yBkhzEd2xY8IOc49Vcgc3u/t00fE4aHgh
f7Pcmgvj3KUNYb8TO2yOcFjQDkjNvD92tgAyo2rVYAsx61LJrxmjOV5kJ85QOnInoAriHjqopQMi
NbZE+hq9x3Kq8+uuZ6GFdwPY5oHT3av4TuObq5U0v9+Zpb11Qdu/qcFEx1BE9SocNTa2WttYX1ab
zacPSBP+hLj9cntTMnLjmf36BZbEVQc5SnY1OyUbbshuTeWNeW17GzajOkCyc1IaD4Yr7ZyS35RD
VvBknhsOrIwd1Wx7UF1lWlRTIKe2rEsOK/pccy8pi9q85eHZ7zyxYcblu/HgATIdF46lpx8QXtXF
VSDckU9sQyNf5oBwWB2I7sDH57dmfJfWBdTJwmVMUd65TMw2tVQsONSgd9zR+m+TztJAphzwrh3/
klq5KO9S4pEh8fUJHnTVe0i2JBE76ejC7gq6RU03SZShilTAY+6OXwJs+itdl2m77lssfo+DYME/
y4Sj8RyvoXdg993fdBfEHTje7j8P3HoRieqzr+Vp5zFJvVHn9rvDOifmXyGcrukd5hfZaPpeQm1W
JsFscTx7r7WmwLlHbpTnkHAQs8U03BgUsIVSXSHT5KYSRXBDlHHxDuFqmOb3qv2bn1CfaIhX6mo2
XeCMBic4H5z/CVBUwzlou3AitFrmRFmVzfQ5VNUT0ObE4LMH4/bkPr1BR/g39WkxPvZcQikosgic
uDVFYLglebBqLGK8o55j4Yqk3L0IErwccdWuVkzV0mbwjhwoYOr7Ti/rP752jWXdqpmoIa3dwkLm
NC9oFPkBtUW/8MRTOiOpIhvqJA4yStDena6YQbwB+T0Um1bDLTfn0WvLyd7cfQ6PUkeeWJJ0cVWi
UHwrHWwskTXgSADgAcFN3iFJXS+GfK+Cw49Coz4N3PlfSVM33/GhB9N4dRolA1E9tfMN+XTDm4eW
pGVf1EkBmqUXyw/3PZ1jQrupORQmF8eX6NqrV9Fv0MjvMSUpJECFAYNMQY5r9ajMEPbjD6VbeeO/
jW97tg2WEZAiVaB4uKXbKH64xi56RxxQhc9RlnDRuzSvSv7mHuJkWQKvD/8VSeJpHE5J/GF3u5nZ
frTMfRyRx+q/47Qb/TNCKWTDHw4VLlts337csj4aGJP+asFQBOzJ920EawvsHdScycSdwZiYkaQo
sFcP4k14kgEwRHwjqhdV1L2+6qe19hoLtfO7CMuTf0uCm5iBczqR11AtbWVfFTpVqQUll+e6QXZj
76YxSPariYSh7N18CTYC52kCgkSQK6wlOldelCenn9M/dfZTgLejFQ5M/KDPQGBVWp0pZwP3s/Dt
8/q2FLkTI7gGnmlV2BSo2KmlgWR/4gNw6z6Tk4reOALJYS8ugJYIum2iZ3jHqJw+etqlv6EanLAO
l4cTS9UcIaSW5E38K6VPoKbaWlW+9XGQVzs+2Ra5ot/7PGV69Nzb+Pxgld+vTgwajMP69ZslHCZP
rOWpBDOo597KrcKaGVfnAgPAGFXXNLc95XQYAg7Fgt8YiFSzRvhcqy2kxSY+6nyqoQ81L18/mHu/
6+m3/qCqDAi/Ez9GX4aGZFaRzIptKQzFONiZ23mZX1DOziPK0ucCHMANrq6Op67WIjEP/gYqaNqc
zz6561PSZzAnrN5+tLVPBIVdpG5Z28TFzCNHz2aupGXCAB3dwyPEO2ZqpE5DCXaT1xAEqyLxCtjz
FZv108YAQuGm+vfNCC0D2I6QMqkkJu0Qbnm7SuEozmfnwHT8ZrJLI8QBK0skZzCYK/Ix86wb7y9k
McEQhitIhwFmLjuuLGcTohLpUTQpbdIfDxwhqvvJUfa8FsXVJYxR6vlNwEF7Xw9Kv9OWIESBNKth
7kPQzI3DnGvZ6HdyLeWdwTATDTVDgYNstWHzBdaeFbBDr4r/gpy+v/cMLxSWpt3FcKRgJHPICdI/
IAxKMcXuZpQkmf0Yb2Hei+wutbwa9B0JzbN3hB3WphQX4Tm86DBKpQyJ+wNfreUGKqRgWbogy76R
6YfO0ZRcoRiaZlTI1g77lX3RU1JeJhzDOnU84kY/Z56sR2BgmVJEdtlcdLY570HIq4tzlZQhHCT3
J9UdFbwHGthjc1I=
`protect end_protected
