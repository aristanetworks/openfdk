--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
W1zko0f5dbga6ngo3NEcRVhhEv+/Xt5zUvsLUE6WryKw/njvN+C0LWG1cIQ2nrAbz2NbvriNBTi+
8lgAcxTc2s2tQEv4WpyuIe3QsDHIYI+sdkcwe/Txevo3KtX+qHYPm0qgLIvAG3ARb1weWMOscjfN
UNtJOz3rZKC4UvAEoDjkOBe22aOYiEKhdKFsmkhOYgFYWhKBIfNfUAaT+1LaaNjnn464PsC6gIVj
JkuH7VPBeRjt+bG40D3hi5vVMOZ+JA5Jb9DFubfnoGYYa2+/JOyRVLCxouuY6DRbd1KUGuOoeEap
2Gi22Tr9SK9GvikiYyuCW0eIKNSFoNmW3TyAeA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="KxG+Jdv2JiG/nZtNFFyTMZ+XkTL05WQ/1fRZ/IeCVMs="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
FLT3/B/PSSvC5zlYZDetFGxcD1Z5FETc0/eQGnLpTzltp7HUVbCS2uKLnhtvgTBTnYeg8JGjQH9S
/chtxPqhNxg8E1gqm0Z+7wigUse97o3X5yI8u0p4E5W9M6HqtlO7G5ntPAZ3CqLpT5InvX+fswQj
UIt7usjPQ6JwZ5wrRq3h82Xx4IfmqKm+KV2vlj5W6hXS9ueRLw8jronuHt/W9uYLHhTmAulJRkeK
aVsxhER8G3cubtEjI4gbctLHX3BWyzZWtOvb0Irri7pvTs/on/KUTf2aYWdOHW8js/fhIA2fmHL9
XtpnMprT1FAhNkMPSOrqyUEaadUXVpd3IFrvAA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="yc4CUxBQjDmErX3bYubNbqliTuGoh1IOKAWeYaxH+mQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3888)
`protect data_block
ZrIfGigOyWcLl/WPu0RDudasEuxS0tCu53eMIOsplMQ6hEVNyQ40epMswAy+lEALHym4upvT59tY
875Hcf4ZY9kC9Ffx+CDfGA6wvUWSPoOo91CJ6+t7PD/UFI2WDtyjuuZou272Y1L0/lawskfOfhkW
q000tD9LgnTL7lhnrJwCmxxPveSO5vfyERNOCk3bTg2gTXya7fSEB5+XA4Pp4j5XNS6gojBWeFkN
4hSs+BZ6EB6MtNr0mTA7Vw/uKU0UVQL4DIVt0+X297paQlei5YABo2is74g874b1v8v1fcNiR1ei
2nspe5slRvaX67+UC4wgdZkyZDHXuZbfkoKl74QXSQD6opGHf3YDn4siBaR6UYvG0b0Ojw3V4T7B
GtE1s8S6EvmiibPgFcWygs9myRVqc0kylRvM0lJ0mVtKXOPPMTdYrcCw49twBpJoEQHpd80aest8
VzsBDvF8lSJlkjENDuAy5fT7LORscyFukxF0rCOGkbv2+uvqVUlGO6XpIqcKj/YijznTRkrRmsHt
vxM48daJ1yeoDhhEdhI7ZusMRMd+n9SMNF3ERwQ/kRHb9dRIKw64QW7K3yV1OeWQ98v9Yo74qg8b
pzLU+YlgpRqLcJx/J1gDfl2hZ+ZinPCw3czn5D06XrGDR1hrOCePIqFS4mJ+X1IGYLlqRcsi8Njr
FdpNK5BczoR/H8eO4ywrTBXXNVP23ArMS63LmgpvVBpIBCXkUDyhJGEA7khjLG/tPInquHp5rlhl
HG2uvFzMMY1LGSAKN+Hist1AGf1NU+fGQmJks1oV7U4GbKa7i8XFKw2EWs2Foyv44tPY5T03CjdK
DT5Prn3xRVN8hLLRCbIn3Q6xOLZqqTq7/zbIiN13CCHgOHT+fRlPR7sX9DabUI/3g1gFrZvf6g/x
7ElNQKutQ89fMmSR1M/ye4lGBiRLZO+O9oVIfGKD1KfElLEQTA7diY+pEsFPOoLDFoPAKKv+lhBq
28CgOLRWYT1XqQxcLhQ8YX3QpSQJ/DzBZ+NY9CMyEzt8U0B+vd+MPAJOOIiYP+7gn3Bz6CQ1W0of
nUW4HJn9g9TKHG98ClAgO+BoXnH3yXKJC/KwQTl00kLNkzLNBN6+i9zmtv5EpvqxA1dGPFvKeA6U
iGPmKENko1MQw6Nk+3mVQgo9EpER0PhQKy9BVVfeDUK8gWEwBOyMCR4R/85xiBuNrGD0raSFo2ls
Efjo5jppVeHo52PleKHNIO11rsxdfwCA1ZY4Qaats2WuB+zx2+9iabPHJ0uYZs1ohXSVUTov8SPQ
9naztPlHvafOrDOlZJo69uYFQr2wKmizui3JFYgSgGNLJSpHPNyKQLzRaLshXrAw6LGHzS4AKDDv
PTn7Cscxz0iYGboj5FxtSPsF4Xpp77gPutiMuMU05gvix8iI3uiub7iLO15rDmvad4yq/4jJlXiD
tEjovGbv1jVcMqS1yYdu+OKhAMSnREMubPMZbgWYYGYllZvF4C3E/OLU5cuIj7rMKDa+zRmFiKDl
LK20sFIDSrjVoaS5jCYjpj3GqF4tiLzg42VmjUbqmYPlqeBZbHrTo6KXyaRqD1tN6czLOYcQT7Yy
2lzUHqQ65KfittdwJ105HWmBRRv8vcAdoEI2qg+Zv6e5m/Dla29Yd6EN5Nifeif28S75tvwVp+OU
81HR5yDgXucZgfRJK52NAwJ/bJKnSlQ7Vx+CNIpz/iADw8n/SQRUDGXONnedauUzMUSNQbdvwqq3
MOeq1O3b+K2nrhOgI2Bxbr/plNmd20TPg3RPvk/un7G6pgjCBWTX+RNJd8s1kZxnZsWftS7R+kKx
tiSu/+ieCTjgrGNWK/z4P/XL8PrCpl8ute4DjcdkOTiUtYFTJzAIy44y8dHWoIDZzpNelgRHhAQa
ZGFHK0rnIJvbS+MJ7LYvVTDxVjTZjIxa3zNCc9xeRT0q67Mu5FGiKNHW5v6IRNHSirAvP2XgWKT0
YwuaTRh7e+QW3ojX6WbHTHggyUUL4s1YC2VmiJ0KXgqU97/9uiIr/n5+btdzgODKIMqQ8L0W5Acc
N4iD/T8dNzzoxxIRRFYeIR40DqcmDis9bAisD1xQrx3qmIBONZCaTDU30ui2rna4IUkaTgJPuVp0
YX3FrqNebnzbsXuUsVsYn7/koXUSeGYQPEyWBD+AnrqZb0zOudX0o58ksCG0gWXerBqAhe/kLh9w
0RBsHaJiWAwicgFz4Im8QLsIm74KkraRAsjpV41UqIPrpoilC245bpg2EfGzwtZi3kUT5PUKkT7c
ZXv/1+zAPa80jkkRs+Y6gTcdxyOloZR8ndSL349P/HVdfwnoWg3BMcqdKWzeLY18+thgd1fpfKOl
ErwRJOatgeNkbGx+EfMF8oMYxAJbdmGLpCxGJdCpJ8vCTI2jjpQVq9RpChVMCzjTrP/UXrLUvX9Q
Uwt6tZYiaztoOaFxEbiVWaCjCm7cM5htp+3l4i+CIOZADAwAhsz75EuIQ1rmbg2/rDj6A8XEfsZh
y+vf3Wf9W+Q+UIArnMoobS0jsH1b/9Z2aDvOABAhs9uiIMj2aKXX00Q23Uc/l+7sLNWegl7R7OkJ
Hi+k0m0q53RC8z/slbIsJ3PaJCUNF9lC5blnADvi5E+04JW+03syCC/EoTb7QEkJ8roK26eDBz9x
Xb00e3Hud6Fr9iuFeZadYZHkIDvhyezbN/hlO0oCASEdpOMwbt4v7HDrJdMNDhhGN2GjSVCcypXm
oB5NrsjKqKm37V4tU9H0KuoxDYMCcsYftbEPDzICLsZenLy/Iqws+uIfjQbgc89MO/socv+Dwvht
Evmqv4HejMX7U8N2ySQgq4VHL51worRxoWRl5RyxIVNTmldn4H1r9t83u2ZdNDROJS9s+O6rSBsB
y185oGXCXU6X/2xrjMuyzXSNhq2ts+2x+p/5PAns1Nn9XNpLxj54dT5c5+wjSgQEX9UdWPm1ivtg
oKZOYYgEt1IC7SeSvKsHJr0ZIr1GIY3t+doH6GXR4RABTjMYIb0Pf+XFi9htuqP5Lr9qhGMZMHPF
RVo2xXo0z2dNInO6mZY671Skq55YErZhPPEvitWrzxF0h1b4vCcyI1MhP2YQdm6I1bUlij5KRuKf
ADKJyaPsjZbMBpbkofHiBTEnEAmB1x5/E9piJKxsWG35nnDG/mTdV18YuMQJYq7tYTwZ5AVWZI7b
JBsK9fD6bGBkwLAKvhZeTXX9VZXLJPxZ3+MPOljlbcmM68GVCuEzsIR7Lc1IlHvCnU0fa+fZBSoD
s3B0UxwYEa5qaW+0raGEYJGOmg/Wr52mj0WZZ5/Yxiq5uBbVpnV9XYxsADUxuDfTvJ1PakUQcGV1
vn6qpAbYJefhRz/WJOEkIOru7uSLkvmHC4mDHiJNkdyT2sSu25BiNptwV6BrE2NAfM3YEJCM8wJU
Sauhs7zDVJ1Cys6HZ2h5jnzQgmHBPujPcZx8dC0iZWrV/XzUWJW/biaAeA7+sQ2ouCeznpYb3uTJ
qFDA34A2M1dwkbK9fONA9g4727U/ZVzBoufPUqV6RT3URzw43VEGm5ZEFxqG31SVaCdffQugHemi
YtlxPeUiH2ejBpRqJ2DiDr2MajVD3irsPCceGq7wo8uPncntK9C2FNGzC36rzt8oNMNA5fBYegaj
1gMl1gB0SgUQTpA/mjJ+QgmyCLNde62XwYiFPdMoU1B1t+23CSoBXT/kW4Rs1j9IhCiSDUCSWHiT
58LcaI4tJbi0JEDc2gS2wUBCrgXtt8/x2y8ePIaInxHI0VEp5sCGsWVNkhrx8xVVxuHqsOufCXkK
8A4+zmUDxsmrleEgL+uMzQXMw6xPEhOJ3B5T04LlLlsgcZDELZmPp6ZuxcUV7LEKvA8n5yQclVr+
n8zIuSPnB4LzcCPAgnrULK6rn4UsokhakUDVTfakLtoEtm1N94qAwR/Hkovojjo4V+xC7ZV0v442
2pkhuw3Nr/JFGGm3B3N//K+KKoSJq4fgjpFHI/bAO47iMdjwqH4+5WR+jZPzkWAEg/xnjRRehkKv
8QRnw88q6mxaj2JCgV6z0cTe14goUxXILQVh7qxNZSXgCMI7JyTr9J77yVSeP0Ls26gDwJGq6qgp
RYLTaqjU03ayDory65SCNTEXyzttSwJMFrOF9NGnFv/QKf0oLaTRQArvxTGhN4Lko0WdRSU/3h/a
w0suTO0A6ZLc4Cf+4L/yieFP6ZsgFNTHgQhsH7DbwmpAnvM4ndiWwGwU+8TkAdlq0mW/ARbIRePd
HniYBKLxkS1EVpZPOKK0IMPV9fh+LtOX3P7BprrCBHsbP5WIJrDJuxcZB8oYlHWXHspxqoXunlxL
1nND9Jn7GxHEOaOuWwhCcxELWC85AKOJNIH0he50DoO/5DlVh6f8l+0c8nAddMEJGOtyN1mEQwj2
oBbEhqMq/3HSQ+JuqGNEOPSwMcNhSnGZ2YnVILpm2KFEBNb/60MXYWxC/ZXhRL8EiDkXP2kCoVG3
uHlFanp3zuflVHD80DLqe94qT2PwstmN1GLVp0DDygnkm3gIyU2rsV5hbtbDWTc7Ss36AfGsx5R5
KUTZJPf+E4X25AkiK1Oa65/z54N8i8h11d2IxkWBZ9vZvm1V4/eGk20m58gmTem3N4OTM+ojhKtg
Yt4qQlRaqfhBaNxjzCPcnqQv+ZgykvNowZyxnid/+nTTic/kYuRx4GNyfJfGlSjl3DsMYunIpZdi
axwlBpQ1QOk2nbvY4jPPrBp4oQOug4BmnuthPKwbhsdFW7JvRveBILhsBWL5zewwQclyaQcDiXTG
Q8ulN0ghzlABmWhJe2JABNOKF5NAo9Lg0YRbWsTxN2szcnXdmOKcSmMGJ/iJV4j4QQJiWoRk0Xlc
6jZ+PBX2pwphuLoz6nSgS9rFYLQx51C+gIFp7B3VY8+NAncC57DA1VmSy3/mqKGwWkmkXa/99y1t
aFIjfTf8P0x0lGtuUGjSgXCv2JxtXjpZTy1Uqi7xq+S4Njsovf+f5OHIrMkpS7HVJHdaBArW3kLY
/zAIgAHE7zKM14mFY3IipcVQRacalvFybRq/46W/FrETzfcU4r2uf+RHux2gwZXk43IkVO1e3B2q
CsjGnbSMCLdxsCWcbY6N9yFICmXLF9vam8OFNlK6KuBgAxUNqobx9KdikzQtFoi793g6zXB/kP3N
GOmBf8T9QPhaUIvF
`protect end_protected
