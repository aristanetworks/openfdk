--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
CL4h0zr1JQ9XY6045JuUd9orj5Dkm2n8UkyGeNFfJUv5ePsFrTIhf6D2jmjzD5RvZVSVz1TPtqgW
BEcyullIHAK3jO6cMYBm9qJUPhsu3ePmXvD0vu5ErIyeqkJD8nHGWIwgd0UiMWm7cVAuFagwH6e+
rXEivwutSEbQo3bvXaJN4gcG7phbx6qZdnNmaIJlGLMoUGaJFj2QT17v5BQJs5b9LhaX5Unvc7hB
X1x579PDmQg61x+X9ukgqEqg5ki4VDSL0hIoY56yT409roOz343rzPwTEwrIBFv9TLjM6u+eiEbd
PBb6mUw+WQI3uvnVArJ0DuSQN+c2XA4YYWE8TA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="GD5YIFlsbzgY9frIwhctSTp+1osHXIrWdJZwkFzJIdk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
o1fKHyOGHMjP+5HsMVJreFfpi0JYymfim9fOdiCSo2jMbvR5sCYHs6wE5b9knS31UR5I8yVzioRJ
vkc0C51k3zU6zDfpEEVC7sGVW90Un9cJiCQNaWJVMbor/n/PxF3DUqRiQV6yNFHlSss139SWcRg6
fIj00LQx1DFLAanU9jO6gVbaBYNRiucHbnWEBuaawjT0Wjz7EsfQQ78hn7bDplleBbCDlnyWv9X5
PRSAxSruZ8BPVZqJ3vqb9TLKV1s/D3YCpvZ/9DHwQpKogcPyUBQ0mUxUzi5KccwN0ZrlmzjJLHV3
YRpP7U4kyJXtCq7EEkmLq1OJN2eqveR4c73yhQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="KuAwQd/qF0RmdXeyQIhdw7Zm8jrKIfAWlCcQhtUqWVI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 29600)
`protect data_block
sbrSp7t5kee1gW8qBj3mQRdBNEJKZO3vpmNWAHFG29nd/e+WK9j0V8+OSmFwJ+o5n5M2eh2tRsuH
jvNaXs7mg96S4v1YrEAwquaegczRK+WYgkkNhQNRH/avf/XowP21rLz6xus4f3JZpTgcrgQELwVY
CKi39PR3Pn7N2Ln5QvfSvRU2OrL7/bDaPWnpUElaR6qQx9jnq+K37L5r5aXIQWVwdw+i9y63GaFc
+ZEP1osEymTFTFioBa3easuE+b9BayLqNnMLOEArrzEEyV9IG2b2WFXh6Sv2G95bOUsvEN4Zr/45
PVO3D1LVngUKzkd3C7GYnp3zRvzQCSaKFKvsJV30dTOtV2kj7wf0wXAxz2Z08YtX/gojmQwtHwOL
kx83qsqHvaR9vpat2fHgh/NzCOwxwy7RKzawZnFuzdBdJ4j7cs7ym2PquBY9p+FDWZj+7IaqKi9S
grMIVliZFABCMr1GnFVH5aAhEpAgROY8EEQBfzeBAgWRtpsntIMIsnHOsvh9NqiXWzzkph3e4ntL
2VFX6g959pFAz8Q+3v5+HePRvEWaEo169Sxm5p7lMeK+HLR4/sKO4zdm3MwYpQXn7MTN8JSdB5G+
ZxkHpTK8N2jCvrLLCLIb5nemozV/1KhM9c01pPpgP0c53k0HPkVtFmoGtTpk289KQewtDdJgIHGz
Om4aGJBjuwMzBX4ooDV/cb4CvlJfJMSvNNwAapdIL6Zz+q2qqhUjSTo2EJ/SlGtA+0oJ2gLLGgta
yV4QbATeh91HYWDP9bqcCMIyGZ9U+GdrB47ygJQmwpD3qnkvX12cTsm1gpA6ITWiawDy8Xyv+Tm1
OxE0zrCtKvuJcbldFWKWenfJv/3Kaglq4OXVKKO35RTml7+1omV9XCllzchC57hbwnaNiJywrzAO
F4QqznhmLyrJYqRN9/ihs87vYkLc2TwmlAf+nbjNI77KybNBnH0kD00Ie7RAUZ56XX/3uyWvaQnI
C/kRH+UcbA6IO0UqZAqrIt+o1JzdM9IHTMaLFcslinyePH3cPClR19tIUZLusFXmC+cQ+KxtIwyQ
hKVGkX5Ak7IePrQcqY+01GlQps/rtAGowyI1jYWaXnzzZ03RhvIdKUI+sCxCO8V8aDbpb9FppoGR
0jXcG2VlcYbC2YHLA69++anqSNrD0NYIeTNVn4jD8qgCSuc1h7MPNZI37BJxGTNf75zDXRUBpgW0
lFYQ9XpDsTuCm9en0jWlCLucwztpkYr1oqpjWBBaaffnOe7TP2+oPyeKLm0zz1Ch19weAsP+B/CP
0Q47TTRmhdgSsxX+7yJVw60HhXouT/OhmGZ5MxB+0PKauRUw7NLp692Oi2mGh3+5lKoIR16A4Bpb
lzRD7wJrsOYlWdhXBAUEZJIaqBg7z+9sqLVPjPy65j+eY0o1CA262iVqSeK60itIBLsCWT+WZxdF
wRwsEXWXv8lUB0J2K6MC2P3ukJGCaJhZQ3SE6smB3X8HOCqGM0ERjUDMmfCIcuWkS29GDB70xhhl
o5+R6YcdNd1EmQTP84+4jg7hJOqm9BgLa9BnPlaRbrZAOp1HKuK+ttk6oyXwRXCCMGUbHnGGdzzp
9M6CVw59FoeE7FlLno4g1jRGvwcKkzOYNMGYNzyeRYIBOooPALa3Oi7uRkqNNgylxoRDu64u7mF0
yQFcppPRLojzlK32/Ex2SsmRx3EsDlpD/nrEiv35dr1FLHjxiwx6koxqS+NqZwLjwM57gO6KStb7
Srlz13waow/shv+neq2reYS2a48+w8tRcyP40NTSL205+PEa6blupPSktsbkcuFWrv9nYHlXyNYF
ohTJtBRNgX2oXYWoz3r7Ty8dG0drZKo1XIVK46UlsvwaqBCN7Cb4k5cie8BP51eNgJNBCsQxYZqx
F4MfvPSY2MC6IpJxPSMKpJYY4gWIm/PqbM01oe+twZydGLMDLbs7V9K2v/8ULIqc5B+JYfj1wKX2
wVuvw5bMCT6cPEYLMH8GvxhYhm5/mzTahelqIRrq+QYcHJs+M5TEG1MilMPUzZ/+K9e/ghwEmpf6
6SHT+80SevN9L9Z6VI0GLDu+0NoruhQLtuj6veLdHqw77bGEtpJbNCo1Yw+ZeLJ8gaj+tHqkvPoP
acAhWDt6H4E7LVpAdFNnZJJi45tivhKbfeUfQoV6Rdy991wvMJWukLItTy3OJCbk/7SFs5s1gdu/
vyRkuQBkoCzv3EtmwubIcd7k00GQN8VURIsa/2bY7Zdr113IlrfbiKLIZ39ZhzyaTHtrzpNfy/gS
Y6gtrh9hrmxQXJMhU6NllOfMSUhDErh4Qm7zRnEwaKNI3Lgfqi6sAvx+L0rNYZ9m1MP4PeYZzxRu
0KRQuDBALwzMxcQA5bQnmibooS+qtsQbsFS8aPobRWb+zcojPTRGNj2t1gjMt0U6QrBuTtxAP8vY
dU+4KBxZeVUkfQAmlL3k5EaikhNDCvr5jo+uUTAwqw+EfrSHBrGK5DrclxLpOY6tJzS+u8jNrgBc
afshsNRvVXTZaFWvG5CJr0V+TK6FRii4GCP5GD8QsdktSMvJ5+Q6Duw9VPXqBhSVXiHPTEJ85j+k
kpgyMOpRoZ1bTGSxnLAwUzB6a7DEqMjNBIlx0DdI932O+U55H9N248A++u7h9RcInvFvTcFLxyTJ
Zhl6YzUVA8lFddT5t1jShB4W+qPzPQEe0n70DtFIbmCgj/iP+T46gW/yZqksmUVKjQAzlIbr5DNz
c27eoVubHe4gJrGTCRdum3PrLP3wDTtV2RJymIM7uEnffX/qc3UkQ3uy59N8G5Cb9HNfpwRKxYly
9t4Cg8i0eC6Txob1jZbQDmsKCZtox4M4SCkMLiGZSKPZ3Y2iPBeuHYG5hQofDi0tW7kz9Q4B/rV1
1UJquXtknRGZRiJU3UzZvoOX+LZJYodulUbDL0EotFTN480uWM9iMxAbdkN5Qyy7sbve0e7WJ4GF
8Nie/HIRQMqY588rDf8AkUhnhhgZB0GHCSwDRHrWpIZmWSsG6mmqKP1NZAnS4TRsNk+T/1tikELM
rGZKqJfrAWyqpEX95gCGDCMCheNS+bV+qNGwsAzh0wV7223UrCr0O/QyU+zUI3YZvNzVDnUYtxdh
5EqqeZqsbS1/WTs4iT3R2WDqyM8zcy/sWE/y6VttyasLCHzREfCGnhofNlEzfztQrcOpEL4CvI87
hdQMsYm0sXpy5syKziqkebOqkD4pQYHPXZRPCfvmQnzSr8cuKNFfgzaQ8FTTF9mXGI+rGP/ncT8I
NaGHrW9uP/JV1IuvQHkhyeJTSMgHZhJoGGxb8JfMoXnesMpC6oRJ7JiMG3geyDF0peDXQVZ39/1b
/qghrfaYg4xwf74TfH78Dbd3RynJqftWsQ7H3l3CioYDsI5GREPb0GDChBEzc+l4/mpNIodfKGQE
TKTABaBGQe1YAPTfBXU+jaXyw8We6n1kFVmnz+wgqfU7D9ATA3IsfMHmT8esfAmS+SVxyyGvlqkv
qgE6sDaoKIn31MuKwbwTRiLIceqzs3HqQlT/TEpLsuBWdpP4FMsIUFMx0r8i7fXmWwlVBynfATNt
uYduUX0voGWUKe9VlX5gV2/VzxHM+L8VqGPErHo5sVaJFcLfY/fW7wbbvm9HFr3kZ6ByQMt9E28X
7fsmBQQGKwW5GqLUBUUN5vLwYBKlA4elmp9qs5PIHq31w9jcM1FkX6Zb+B+8t6KV+yo5eynZKTeE
VgTRSMupKt+wPo0lK1xd/WkQqz3Yp+eOZb21Gh5YcbCw7c0PF4xLxe/t4JnsT/Ue+JaxopxPbR51
Qi7aTSzE+gHUGDhjOYwe+4mWeqxALPmLvbAQkpQ8lvJQs4muv0Sl+eUQLQDwYL5p+4qboYC5KsRo
nluK4HBA+xo+3blfgHrucNU/xyCHitMHakpRkdKWgdOQic2qfW/6+0g2E0umrO5G2b7BWrBfiVKz
1xqMtUZzWXsXCchS5/MvcVPoG5JXCXuU9Ye0zepiyAxzy1sQd3va8T+9lAZhPiArb59miDi2lyIn
DmugPlQulWhn9GCLIXcmhym3XtTiIbzZb8MImtdm748WYWBZQy2KiDrX6yMb83SYfMnaWE94ChGH
Nm6IjLiKbGHOx53BT4ud48QSzlafO+kIOUud2amSEaM6V6qus2R9zPon7NdtDaUH0Eto52d+6+rD
Vcp1kd+Isr2osjqtk3m5ftkDiBvKy0d6TtzXOYzb51cIfHBW6PoV6sa4KNwxXE71yTogJYu0mc03
IO0+RSu2EFT6fb0/l+6llnFCaZzurBowaq0GSnL9v8pspup/ebTiOasenVIa6E89bXcpI5XmR46r
0YT0t7UtSfYPuOZw41RoNgPgaDWO7Rrcvlxe8KfGeUqquFJF/Ho3Q++EFTzuBGeqbds6ar0VFfJJ
xuMle0ag8jK3qPYjj2ZbjfFRG3FNitqKUzh01N4ohltYSkCa1mEb7mfKHWzORWpQdd41aPzXMoBk
jplUBATgzjIZtnoWh7eEBi+VgZEWjf+YKQsZTIGcOTwAYaBSt4Df8u3l1Wcf7BZJzZ2yomR3EkYn
qH+gplMHkbTE0CCmiU1GADG6RniXLMWFbwLq++fl+/L1NQyf/YWzG9QR6JUa7MH1R4A4TitHGWk1
DHIIx9f3N0BW495l+Bem3AvfGHHyf8qQ2KPnyquxKC2GbCRJwFjwUz5AmePSgKKCWZ9wzAopwd7a
6QzLc+cof11m6AzO8C8npMLJ6OecuUE6rtPfpApcQsttigORIQFqw5snq58OBxirXlMBQCYJlH1H
WAUELNtH4xqoTHrcM0LNKIE0MUkSSJDkWW48x/5Cvkk7nEpvfmx3O/RK5KXVDsszqxsMGK6sS/Wf
949cxOUrOCHZCF5nRypKkOz+WKcnyfjyt2oSBVHrOZSwdk9YaLioiRGvfr9h2bBSYZOdDshtCn1s
bc709q3bI+whzLiGbKA3H4VwfUUri1PBKQal9/nUWMXGH9VcqDSN+o3kGlMLYfK5of5esO3XIryg
NdQyDov4U3AuDI6AnF7yYi9J3uzYjOEIdB5l0J28Wa2ihrS0HhiI7vV0wyZs7It/wkFwXIjVs08L
bCLHX2fww6r3t8VRF49szYOngKp7x9rhVTRDD7h148WedqudbjVM092++1RzgwtRs0XqWj9t5V0q
APWOCX9EoT7BpMbs8AR/RpuVQnCZgiXGv/uYhWkmwXaVpn6BCGBSvSdaO1YsAU+Vo/V20Of2+RMp
SXv09kDTtLTEAk4H8d5IQKpSgjb+NnWkhSMFgR85tC2wCtawn/r2u62LnU5r1YDHvHBN0XONpkzF
fxLzCy1gJpA4QcY0uoisnpFYKW7yjK2N5G/ZoNQsH+dhmk4PylvR0KUiArvyhcQSzdfMY61EvnGJ
ZhBHV2dFGeyFVf4ftQy2cW/TEICnPnOmBGqviUuOV4mb7PrJsR/re5GND1lZMz900BBVUpSE9jZN
NPzmb3j0fkmXaP+VIl8asO7eoTqpDL7Xgtfp6Ma3BVcCGr7uLWMPdLsJG35BT7zr9sfzh1n6cOEi
eNSFDEPNw1F11V6+AijxONzDYCY3pSc5/P2+RcQyI3tXAgRo1QlVi6YqSD+iQ+1dL9jWTMhwn+5g
fmHf1Mj1Y1Wyw001GrVH4v8LqsCueWTXTIr3kSpuXtArEVYnReD9zVJW9wiQsqqqiMVuxp66T3cb
mgIfJfcS7Xu6xExzxVLb29pLGGmPboMjzExqUlFR+SEOxAnc87nmsLStnFSnXGQk61W2CsN8VK53
5wHYDi3sbA+kzWYIhl/fk1t31kYigqUOBvZ+YIKPX7Ynk/PntKPrIW+W7OYY/izgnntdbyXX+lo3
97QAOrUxrPmUdEEOjSngnvufhLkE/kbGiW0HLPbcWC8BkYCq15lS49VD654N/0QyaNUhz9aYy2ih
LxfpY+3ticGimaplK5OMkb74CP0JYz1XIdhsdlS9koAEn13DasmnA0h4CNE3lzMC/Kzq+Xdptsli
wQ24WvwXGvrAs9tlAx0cyWns2xcUsEkGPKdO9QXy9Q07N6SggNvvbMrXdzkkfRu17Cdk/qwY4qne
qdthZhbSHBmiy5g3+1jr1b+ACQULoC+TwcLTRwfzGChOcy6GOhAbR10XdnKzZcyvGq171aJ+Dh8D
mYN7CRxfstdRl6tZhbBvuz4VMRc8ceJqM8RXewg3zZa5bXFGVe39bWPaFiN/V4wJzdRhaee9d0p2
AIVc59spRS4EhugnO0IvQxD6vdM6YTyAgzr725OuPK0peBE4PxmjvOPyvus+UVHyl9InNHKwoyJc
uxawg0JIzdFbXcJ8iHV49hei98juD4NUMfEauRXKVtKPrGXvkjz6lasYABMpcolxhRpend9ZA5k3
VWeG/ABIcu7WGgR3J6SO7I4AseHG0aSNWTMGmKETXOq9iWSh94ruS8ehMDReohksRg/nyYWmYH6I
DF9RQ18On4bFYCiHTOBeMFslxRPIQgVOldLYIwZ4wbFKBws9ydW5t+RnvpTClVlOhuKX2GSOYip4
RWwTW5ijXDJVMIAJQSKN0dVe3a2mtQ8QuEKVISjFlCxBUVUinpAfkGcJxWiCFBGYxMiwwB4nVmZl
M06Kqf+UI4DCgT4u11HLXMRWvIqEQ77TgltK3zxYOdDLyeAzFo4j8PJpp7ToUZ4n6LLWOughauq1
iQg/m2mT0P1WwLQx2Nt9MFSvmMkjGxH8h3l8x/mqpy8r35dSafGhOAYiSLAzyBZ5wNt9/IvYWusm
t3rI4tYGrFibVpufuRplXCBRhuiqKT9vnFkRvtme93XjA1OLZwo0MLygJFlbHu4InSCr8hzNkQWZ
Slexh9WeLdAQfwLtNUe4igXFaTazDdLPeHeoIiXpxMOQkk61usHoTiTwSADn5RGnW0atpvOSa6O9
IHUwcNDV8efcf4aKZUUIZPj3v05c0mfLE0s7WDESszS1DqqKeIMljMdT9Wu9o466iZ9oXwTPxyN+
1hC7FvYo1J33/ZcTcHo9p0nRtwj3gG2SQruvWRaUUnFJKuSmMxASaOVlgKVuVfpqimC9ECRJYXqv
/XL5KjZhsoO2nv5lohdQFQkXK2gSaOZaf6aw9RIuon8CG7HEpcFHhFw4nnf8pWdCQGdsHcb7d1ud
bku48JoPRO0IMOXwLArjAfWMuxzxViN6JCsFuKSVHgQnyeOSQ9dD0567vbrJP1SmQrpqnulIi48u
i29qPoXQLs1w4wAP7mtaqtcjAOBaEzQ9F+6py9xdcMhdtExmCVP9auw8Kzj7mzTBaZRyPJcrSR/d
Y/0+sULoY7zkssjHfNqVJ86MIcuP9Icq3Ojx4yeKdRuMVBgfGub2jhh9WmiuefBG3SBeIvvFra+p
BG7DIZetgRJ8zEr2MwGEnBf6X4tsHRhkkawjGzTqxx2ZTjtXM82K6geDULnL42ylai361+8EoP/l
JCmtMq6FGM0EepcS/+DgZZbo00/z1poVu0mKlcmFSboPDjyLT5BOI16rLfVRLVlr8OhTRW05A+II
0ItGGO2NVUlV2Ikyw4VDaA/i5iauRLQ997HJR9s9XLjS8vief0ANraWo7r8x4HuJGc77ESWb6V0m
cCNJ8iM+QqBfG4DojJGh05cOUGhWPy6b1Vymv+NxfGeRaD12WiMO5NFEr5J7ybnEQ9s/5qHtm+Ei
3HpxzPakdLaFT6QvnMNjFgO/m3V2xPpRAAodhgTU4MoAJk36W+g4xV6H3vUE5qt2F2vAlf6swMhD
2dgHcQ7QXSP04bCZHf3UKCOgIBVtDMqMcdpn9X/y0YAtJ5qndJKaLEwEOen8v6OKYRzjtU047Foz
ttd6HeZVXm0cq2RIsVWtylpd/4z/UHv0+894CEPDz7ViMH3T/o34nKGqniQaSLnWyk13VI71vFII
HuCXZ+STmONAGUpq1E954JWnX3hZarN8Ma8F3bU+1/Rv9/wjBjRWnNqp47pXXLbzquchfmDAUznq
RUarhERkySotP1/nqF2NNCMl7utgJsivLC9LpRV/a0F9JvHHgGHa6ObopfgpgV6iWa1pxLIybsJU
GOrjeo6hZcVnW2WrZmKx7v/xBm9MRUBiGR25kXc+TcLlmsdym7kUUmlNKIurQd3CPsLcuS9Rneg0
AsDfWVrgtR3si9gEd8oSaItH/h7ABGq/YU304/IGZDLkPMlkMD2dfo5hqTictpnGJ2GT2lQqssVf
LP226cml08Rn47U7mms439V85FOoAf173nFBZvpc7vGHGhuV3L3o23mD5eR6971+77Kw22z04Oua
c3tG/r5thp+nMaIAbuFU45PUAmsTIqk4phDYBnR1ZONHumglaG0eEA5QmlS2QEet1gAFVDe/XyCx
HVtRBZKTxG0jG5WabyTiLvxwwXhimvui2uN0kYTGxAUZVJgpHnanskgPNtzcKuHNizUtnYsEWQPN
6ul1QsOmwaKBfMBsVGC2//hUksIsW2BNz+GFDZMqJESguOL29ms4r+GoA9mhjv/07h+Vc7h4X3Yt
GVukG8DO3fGzIbIChE+BZZo4mFJaSot5uWmKcuf78EUoNCG+GsRKMerAh4lTxQzC7HyFX23uzc+6
V/zDETxkAZjXFSyjdUT9buwsZOWdzNy8MF0qvtocJp1MWBEv25OCSqZgzurGN2UlRUm3F4IDgyLR
BE9wZOwJl0R+xhgEtajRpyTAbgfEJTKNPQuP/U+AE+dE93RPUHgHNw8FK7uPg5Odp5N3oR1R9Pck
HfYDaPx/P080q1CBDHu4S/cUZV92Ma3UIxA5PtWOF2u7YXrj9fLTRSN8JbwbgQohoAxozeGIlJ3h
eGQIty4umf1BG0qBhV2wdnxV2CwMmC6mKRtWTHxSDLf35/D3ItKvrFHNoqBDoJn6p/+5Q1qsM5CS
uIiCRcmY0oSqbBN5ENF3z7GE+bwX4Mqg6qpbp10n9S4om817NDwF9DoXNe+YYGdz+qry8hHZtcqQ
L/gHlXQ5V6tLLVgBCDHFaFRe3arwsmBxwc7g4UQM5rKX34N5LUmono0Y/9mdsuEqthKnHb9fSFzE
R15gJ2Hj2rGK0EIrHbbId3z8y8/Bmmxwur/Qe6H/7EomLJJLJTMOwl0A3pKkZSIIpH50FWM1xFZy
evQg5ym6NGCTKGbkYx4cD+lo8LqQM4lalLgCU1PB+UImvQALBpPd4WBFmYs4dNC/6bXjeaRJd1ul
WnDOBlU6hgsLo5r8/BvHOqR8fY2Nk/ANLzU1SVLnRSzLs07gguWqpVzcqtQgD298BXSPjSHVCKb3
BJJSNDRveS83RFDh3N3fDnr3oTiET76EEZsRIhwXqlIoYbOIF1oS516FcmIe6LcacBM3IDJLeVcL
T4f3gsjkkObFVx77MmDdwoBplMiA2KFdZLUuc1rPsJoDMToHp4Ji8Iox3MjNDY0rjoC82WEl8G2j
+SgHK+35TFmheGa2FCm0RZF19qwjCJ/DCo3T7kUdahvOjrGknunbCVbpUbrPbqF7ttjEQj3Dra2A
jEfEwrHiO7PRCxM9FT5UML05OLJhGbr0g9Y0cqLxNXBdq1uifPVquYoxCctmQ0D5+D/h/FgUbRuL
w2mxwfZNYytzI2qdNiwfh47wYmbMb7iNNnqdcO0NFJ2ElwFUZsGY+017+WGwfkWa+EfJELNhVc6C
nZ2cElQkMl9VDVYV5FSIXlyKuPmxFjZ/DCmjZz9ftQspCsYHyGmjGmtMYQ3LXHZeRkDx/dXUrJpA
OrwIloiyAcRhQ0wWUWkQ0uJ0HlN8j1tBof6uMDBHDgNfbSlbXcWoDYvsdmE/SBo5db3Wxqy0B5XU
8tBunlGKkDKJ0cA4sBb4ctOZq6cAPZf1QvJBETGGv2y3mHC4LnrtkmkduKAiNNcXOYjuCn9ziuhY
abjqvfr0OfQmlPR+9B6PWb/JQaXT3wo0x0Cb6lHeiuEbFlwfoWaUiGgkzlM5jrtORdBsy638qn0p
fwL4bUWLmcqRBb7A5fwj8tBjy++C27ww34332IbMXJbFE7iO1HyyLlgl/wkeQlb89voihb6ZHSs3
RjwDyn3fxlPqrVgbyKyCbp8pfN6yJFwQo3IKngkBrtEcgvDPXz9OhRBEvZXTjOnSQDDUywyZOGCC
5lZcIWuH+ImcYnV4PIYuz4YE6LKLTmeuUfkmo9CMXpvFiMyZMN6OLDOhxWhLx3/9rCUCnf59TVHQ
jU+x1UdJ5HjT2SdxZkO+mcFNxyPkmVLd2pTlgQiYd3MpOCioAq+TLVAYXU/bMAFBC+ja7sVlY4fZ
YMla8Mej3PJdkMKaWmiUCQLo3u1rCBAofjP6XZ7MWQuwHNlhDA2h5SAiBqnQ+CdUwdPfeU8EOYpn
yZKLByL9RsXBMGusMNQe9mz+HbgpaL64qH7jILNAthmrI8eFCdfDsQX2bklpizEPZ3YF7i2WVxfn
bOjjsW83pxzfK7UCZ/GVt4/Rnk1ChKyM+sHSExJMsE6iQR5dLzrPFKnPcsMvXBmgNwyBkHGRxQXa
OSkGPH2SkIPy4gvML7C7ME425RE/PWb5mIjtxdCkqeltu11nqjbdG1H35PMkBhYhL0BoOIhVS/cS
0nry6xVNHofHiFBep8L0JcKVq7+OAgz6QRle53N5rUL/W8kZbqubGv+bfPF+QNhNabq9H83e+AmI
/huznVLierUqVHMf+mTKIcfV42RumQwLwG44EgvMojurfemVkmzzhCu44yE0A1shHR8UzCnmDpLU
vFi1VweXx/fTY5Ublj9aePZdyw+6bLPg+PmUbAvUoi077TijDyvlT52LahiRwVHFszub9IClVDHW
ZtNJdV7Vm6SMyGaHdhRtxXQQpzfcHTqSOQp558ROgHRJ9G7f9KDlUwftUbeaVyo3pOaIsM2OcSjK
E1XZ9q4LMjU3WJzgw7ppWOCbmIowfjfuAmaGjJb6hxfuU7VbddSQSvofc3IQx5DoTbVbcE6YO6AR
hvpuB3Rx/3QsDXT5Akp7Dt4hylvvfgPqu5GEaxNfXd4QNU7B3ZfpobuHGdWVk9UlZxgWAfyna23V
hOTd0tItQwZIUJfp1RaSUE+lyVYy6BlxZSVfUE2m6DnpVK58yCjWs6asMciq0CW7AtAKQc1EGeO0
kFARg11jcFqDqAobICLKfK5EV8M/u00xnc59Y57ghkPJY79urEQW0P+IXnrG3/ykBA/aR+/2cPkn
tswpk5IlHPw9NLkWpUktEKGd3aIqrimeriPRENGxFunG8MfZkI70iUC2LrRFYzr901fEWKHHrlcT
WjWyHGUkYb0RwGUjP7bBO9OcTXnw/9NyUO7OV93bvuS48r71yH9K0DeeZAgZZL354U3uPMVWdOQx
qZ9/XHEDSW5NPmK6OueYs/hpdj1A2iYGFwcrhrUdrgxCndZg4lzO2NieDCdEEa0+IDUaGfYvGeIZ
6PoZWsF13k2uoU6WFpWZ+twUsWf4tdrPC3v6gX79y/u25wazYSmQev4/2aXF9bhJIB3d/Di6spYJ
Z4RyhuZEdzvV9DnWMLbgE0Au/bX5XTOy/IN3BN2yOFYDMtxd9kJdqUKc57qGLdGxXqMWfw/holly
R5sZ6DAHI0IDd1a5jBk5Pf6S09tBEw61YZkb0sM+amL8aCSgFtPqwPCUcWjZWlLJ1h9wmuZ3rccK
gto6eeyZ+PylJV1s7prBz0nP4JXf1WDZFsTGZAGBo5ttVoZQPWApxXLPw/UqWyh+g1yjMsn3psqe
TwTtIV6m90b7q18NqDsHxhmoRN4ZdaOxsK+A8LkwwvHXKG4DUfw+tVe14pCTd6onhbgbvJvydsQw
SfyYy6b9sN7iJdgWyKM+ynQjJSHRP4Tyw+0apqyWVi1UpwBLDGmXg55TsLsgyN9heLjlWT8CBQbN
Aslp64C1+QTJiKMRI2kC3H84Lt0fe+ICIQS8w1ma7Su+Fx7chiiXfRQX7Pfw5OtVkHz2vbsKcaov
Oe970qUylSznHM9oRfAUKZrI3hpP9Mnx7uj3l1dlZ4idGtLiSXlbSyR29sCvGIZ04p54uOQ4fEXE
hPgg3Javg/7uw5UnIHclbSocPz+SFPJGVnYtOHRO0UVomvZ/97+yDverPIbz6m/oczYb5jBhUq+A
kjPatmyq6d2I2+d0s1+OLdsxT27Ya9eCWxWGF0jZmL61ggGOJuMi03Pz1wUwVZGyTETRuT0qVav0
eZMOnX/+IuzddQ0cNcFype4euTrwGXeri5Gn3BloWJ4Zpoo0FL+fORpYkAOy4gYUHvLdgm/wRkWX
bXYpIci1hYcv+pxpBXKl+Dm+IVb4RvCRlXYYfzhEoQUAyr6bLZmdpiGDnPyIpzHKq7FKAnOP9++x
nrjI1aneeGD8mccO0H8l0wc7qvHkTsxZn0/nlljuHSngciQuUTPdYwXjmn/QbhP9H+fxhHbhmiKS
wBjin9esjvJqwvAYob/YIDyjkH4r9ysek9Cp78bSJkgUKW+YNhxY0SDrz6UwDPvixxenPdS9XiUo
7+DW4YBHz2HhpykwElVIoX2g6vB2HVD4gpuP8AKuvyvaYEHKdnpPCFTX1IQpXFzlcLbollTHzD+d
FbXor55pz6Qa68rQkl0e5KAHtKbXZsHIKW8FsR/4GxB3+fxAmgmosqCMpEUqyfw8sRdtT7zClWqS
IC20rHZxIt9xS9Of6f6IFuQ0TU/KrtEDp5vlyIHOcYEn6mM2OlmHesMCxv28ZwY8o1yRPzbv/4j7
VZ8Pl5L5wb6g/8T0Yz3dM3VDRZ6edp02imLYt4h8X4AjxxhrCuxY7W9RNYKOYRsFTG1m06Y+tE5w
lUr6fo+N15wEgOhXJ6i4xRrf1LEVI3/RogmFBTOM7pQpU+BA8MOuagd6D6RNnmrlj+OEGvGOzzr6
ejM68jkCviwdnjSLwD+M4ovrybZaJg+3BPy9mvS0gZxiMBuUb5moUyjV66E2e1zyMh8/a5VRiBcW
oyd4KuiPwpqAmn1BbDVZ4qoS3hnaeTrF+bTC7f3gzKQCauN3t0ipDk7YTsdJcZmoEV99lEb22lCg
VcfeLcAPNG/6WIu/qkmEMU3Nr2E+KgwJ6UglDq3wocyEhNwm5rekDxQ3bIabBwL+MMREU7Ce9TUK
l/Vf+2/LS84+72SNwTmDdwzsjtr4aAg7oc5n34D28Xlu69C8DEijVlbxVQ5IqgONs74dbGmQ2ELM
VWgbkN70KrFzQPw9P3Hm8uSNsYV7iF7ZA4dMNgfcXVb7dALj/+56jEbeAYdZZigVNCsVL7zy9wxi
AgJB1OzhyFQ0rVo0FtHIIdUkdapqjr0smsjHOvMchocwPZNpTWuZNhcjxGTb57lD4OuaO5DAFnyD
aK97v/TCbkkuzDF5Q/M+/OcnFRcD2O8SzwEnT+yiCXwMo5XJAJIsaiMZJz1cI8UbGIi244t59/D0
n/snZySocP9LFBdIV1cWG5nEVb6tVglLZuHoqLnArw5rmUOfJpuprgDsgTqygsnFHE7QZI1JEiFb
NUrFCPwAbPGNg8E0BzmKTLVllXx97dFZcm12yxtd5Wggh0vdMP1CJ+d2I/jovJFEu53/GzlhcdVY
D6xeAmWEu1a+YsMGNNJMogxTeJy/B/yClmcmnQlZxLpcTZbL/QIdWNhfr31Kq2U+0Knjgw3vUzGi
fNc5+pLh9kCMxHznk8Um66ieeAA7gSqaMSgIEnogh7w4FjHFIJmgB14gOU8uwqbDsAMgLBasOd89
cscsJvcuiK0xXwtYfQ3xW8FHJXsi4lAKlD++NlGaKlueHbqL4b9RmgjGpzXa/2L7rQMhO5BwI4Mt
00j13BDq8geB2T3VtPxxNA4aakFIF8YJ1lfKx251Nd0oPv6px54ULb+Lf/TnrjZPXhUG6KPdIdtN
bmHLxVMelKjNdf5Lg5/0PzSxqlWYF51k+5PxDOsbwoqB1XqdVgRnV+V5W3oYn5yi2hK8gMIG6cIj
6WkLDdLUFELfYS3cduh+PFhwgum1nV2frgKd8DuDRHlBjK6+hfm3Nr0oFvMfPyPRvHURQcicQPIF
rWoXjmQOcNSyAuA5KpgszofAWiJRfo22K/XLXJF0Kxrg8NlCMzB3UfDHVu/kibrmv08odnqWpl/C
1OPlN3Nh3RHR3I4xFasn18IYZAlppP9UBT8PrxTNUUPkQmxL2Wn7Y39R15osyHTS7NZotdv45Zsx
ojuAAXXRBPZ17Mwv6B0uRO+xXDwPxT8jJK2T1kgCEqXysiK9dyjdXl/+G5giswOybd+b19cPI5Ru
LeJ4+QjpaK4ZqHz643hd42pAutCx6e61B91cmEQqzm3nAWjXHV6YxnZ3i3Q7sXk5za9UCQOqN0Pf
tJb9tFpEuECWnYt17bWdrPYmmhlGhkzSPW1f6YT3wuUg4An36V5djhF6G4Y9IYwFgw/o8k1emhcV
59gQ+tFW34v+tUp+oHEm9+JV0MyY0xrqQsQuxBODbFadKqzTA06e/C7LveuVhHtzvn/Ovx3r37/E
GNIj+pTy5PjS0/BCZRODU1lxLqevmx0kaKVNqUnO8cgENZtX4yzjL3pVcqfhFzQ/nqXwh1hUFp/v
1gS8QSj/OrKSkT65O941P5rQ/4aQ5LxLcs57hpKdwuoXBZ6Zgqq1VuGbDIt0ZZ0voWA781wxUg6B
5MQ4aTZ4jOTR2rm4PHWsVOVZirPg/wak8LMtnFHOLvkFuvqcOSBCOSnpidN0BhNyohoE9bTiTEpL
AvJ2NqomjfX0g0eG9ekFdt+zN0R9mBBVXpGYSXr3icv3W46l3cGN7AOtvenCzWwmQMps+s7RNT3z
oq1QOZ48ndLtOtW9aBouGrrwMTLtC6CVEP65myYoHFaKWDhWyCJXhMmwpcvHHRL0iNCy7FIFslWh
sYLNEbPEHZprEn/fk8hXZVT3K/witWibQR7gqz604ZLv0kwc/kCQbzn7ZKNlmfGj6wKXz2nwdWI2
OUXDMwYNUZXw7Sa4nb8DPebavNbJK6FkYSDCkCzqb7xiazhZRI+2yyWCuDUrKJNABazcRlNEGDad
Zuo69+FGiRygBj3vQspt3EK9i9gYIKBug9U+loAyoX0stg8Z9+KgdtTLnNyBXJw512BZZhq+eHUe
4rcfLYIuhI+I+hBDT60s2QVt+r27W79AERLJj04+zf1GKTb0tM7/CuSQfDUDRkjQSyqOGTKiPJn2
BjlEDtuqEaCZrqUDMYdlpyjYEGzVRasiLZQ6/ntCBwsb4A2CpHZ3G1Dkps4C9q7VTHXfN6wOipfD
rD1RslczXqkaWgsAprHOYri7Z6eWpfGKnG+9+HCvfL9yIfuSp3gmG4yAUGNaNt112Wv+JnEOKNPu
pHtB1GZypMNrALkGeCiY86RofjXnJkG+PY/ZiYOR4TT8tQObcs8eZCaoh5wIXrBxgUbwCnR57Juk
R4r0iwOvCPmSRPzt5aumCLc6F5stkBNZzlxunaQ0Fbf7T0bIA8ukYTLWPgqeasVsJKrgsznxhp7q
l/3q+kVX1NQPf/YoyG0o7RVMgQaPG3OchLj/jXh1EQhjXj6EJD9bZzEaYB9rKB9kvNtHZsUl1I1z
2NZPbHu9naY07ynu6g4Phph831bZo7La9dR9+Sj9Gis+6s4ntM0PEWBHRpvou3XEYxdgYJTK3Odo
nMMhcr9ur80zuc6Mu9gJDgyXD2XY96+/gP+sdGQfwVcQE93m/D0lNt7K7kDh1wQHJPbiFD1lawEf
qvmoTgwJaXU7R3WrhMTbmfawKhpQwGS3pNMQoRY+6rkurSoDPQ2F9g1PMBzGEqMrd0OOX0iye/A6
O4ey0hFyUTgHnZBscRYYtP7qdHxJIKTXbqrMZtSuBE4rjGt1y0Scs844yscsCXsHcQPmSdZs+VSb
dE1sxPx7Hq9Ichb6rNn8SiVJI+IM4XxCYNNxY5ttn8jrOW2yJYTEVySDT+N/3YNbY2Kn9Jp9kOjM
4cpwXOwUFEahgAF790JKZ4xSmd6zVNobMYPlufDRTXaTrllm37RXOG0GstqhGXLCJ0MOVZDQxGbS
fWZ8hwtovT204kLv2M7ICxlOcYVzcGRXq+0JheaLkHafbVhVVfKkvsklAcBKryMfyROau+fGjXQ8
3Vsr9RpYsYdcsrmF0zo6ssmksLVITyDplTU9wVZxkKtcEEPgRJ9avLVks/zwKUDCPmwK83yur14v
/c1uq+DiQfExIzP6+WGS5v0/Po9rw1RXdy1rkoswLF/nSScqAuMtgfqapyBUujKQigf9f2peSIDb
F5j65GBmAgy8eGu/67ic8APwV5jxQkdZQ1qA5AwWn40ZHN6LA1aMdtsKQkAh5RhUvV0GZOlJg/WI
tck366Ehvx4LtMc8kdG4KNgnySKtjnxzO/GZaxVa0WyENxo5JItXmhbOfhEClat6khZaDgokLIhl
49M2C+LXsGeTcSmdPeLg/+5uksdeQN37pMUbrecPyxodv3gdy3lOQ9O+Iq8dgU43StVV9Jzp85hY
GCAIL1l2goUBRIIXqB7E486iXB+JPCVEvZ/PVhaFoZUkZCKxBQsElWwX68eiq7WfZkNqjScpngh9
h0rag07fMYiWU30DWvvkVQ81OZifDIeIwp3Zn9u9NFXO2ZU8FlIOW1yKiltgiye73V35OKhqi10E
5JGWJNjHyE+wnDIbzjvk/5XDDXBe2UT2CD7XPX9Vup6pHSJ2JRBb0a71rkA7KfR5vCsiKyBNx6yY
o70yOKsUoKWtmWhtOtzLkBs2zZa9YLlu2OOLviIyZaIKn9KT8QYWOzIcl+52AzzLJbRXXkdY8zkw
gve8z4Adn7qxE/727cQmlCtaXthGWa2/aHQj+uXpPejY7Q8kAzpP03pEkQdycYqnth91pBcs0VY2
joeApnMIgrGhnGKYsTxTvz9wyBk3z2l7kfqB+fQiVwlKTjswQdYRjFbjwLtvgQCJglUdmZTkJRZ1
deHiLMPYqZ0SPx8innO0nsSkCuOHQfO/AzKDCMRGVEGhPKI943LS1xS0xxsivyNaWFsE/y0DcJ7V
AOwpR25+Sz/yKMhTY/5A6FVZca0dODPPPhGW2aHdodH8zMXwpJRUVGjWaZ1c3138L0zNrSIQq+e3
dAuWt/uMVRXVRnt6Zf+ASBD9aCAt+HspJ+/cOBTKDMcjdqbhdWhCSDFlZ1HdzqIqYtDCm1ScyXwy
GSV0vzKIxUZ0wmhS+pZtfm7t+atEmJrTmEkurPhrDIgQgy10XIlEnu5EkDgA2ZO2FMYwiwnKJhht
pySfAc0AKCPfMCB6GW6qreMWSEtlVeIcHBxAMuzi+IZO199aCPA01fQw8F/E8XcSoaK7syvXQB60
D+c0Y5oy+yvhmT8FJrSCdNpV+8AcRgrT+7mbJ47O0yCLAfOHDcMNSL+O6PNgtBpcHuZuiTXqViAb
NEgb70x2lXAy6YDE5AwANP50+3kKwjXPIy6e36DjP+qMC2eyt5XPlzTnlXrY30/lpDWqzhzZCoAU
7cHOzUmLnGXham42GXKREHWGjacbkGCiY61oe6zt5r6dm7rMwwm2zxlJeQdmLPV/ZAPNdeoj2tq3
mUrZHWekZ+xwe/G5OGIukgu4MBCbQui0NkjELuFm7/XW9zUj7Ahi9peFY65mJQbN1zy8pNS5Cv/w
Qs3Om/2nHibuQi78JzpCN2uxsxEqnBH5RK+jUrjD6QWTmUyrLWOevvtU1Rhwm3gtw0ka187GZ3Sh
AR/WHPSczv+oYZF0KfXh/BYcXZSeqKxFWFDPKI39/eAqywo88t0YmXtLOWULb4LY6zUMuAI6dhHa
+80PofpQnjf45tpH+XbzrvNSde7ax03OfXVCBs1J5/JvlO/BlyvsJ9wTaT7E5YxQb8u1m7WV4tp0
LRZazuqk2QsbXzacTs5fAHUlLn7d8ZxMj8P3ehA9a3wDf3yPkDCQSBlAc/SdAUAbN8AbxNgaOj1E
24N6roufDutWvHr1SinrsDL3VK6rtE2lx9tszxfUSyWJ5S+87D5fFtQx0nzJmL6rKIxE2RsB9bDZ
2ViHaHsTQl7W53Rco6T0yPwaIexjfB+2cDLujst8u5ZPqUCHuv9GtsxkQ/Pqke9aP9RdiCDpynwD
4N94DguzR+qjY64zw0tK7VIkXmfedd83q6lbPMVP/o7sqHu3iWuNqG6iRXhx4EhPZAC5XSelJFwB
x7GhbrrMekLD6eCLCKtNCpXyf1ceNM+MGfu4ag5I5eZuDBIJRgBHJn+G+XSIjTMbJpL4V9BsNV1h
t+kasXcYKBS2j9PbfgKU+hnlXmXmnfxH8gwYleGYLA1wug58OjIwDjOkG7uwDhR6wOnSGa8RRQ8V
D5pGD/3KaT4r/fanFTs+Hu928+Ak7jn8UAMlxbNYc0haHRN0EFggp7ozbMLelmv5mz/DOU/LdKYN
ACvNafivjOXgM/npjrDznBW3GdSiQD6sT2bNnXSM9BYrV0T/AHvdv3J1djx2dwaw6O8ZBl8vh2LO
LO4gdbaoQ3FZjEyDIQ1SaiEpDKC7P5pcFVuDvV7YNYI7S18k0ShwnJP/pJwY8FO2R0y1z/BOfI1j
HEqcPMpkykG7xpe8MTKOJcLfvH/QSLRZcFrDcMDnaPqn7MGs32Pmxg6DwFHoy5VoQwlkuZQDCxmB
fIxbkMyDTrhQpHzRXkSry6xgv3CsuPUASB/4UQ3Bp/tXQhX/RNT21c0cdxHB0Br4gjQmomut18Y3
BbwjI77cQRcUkBVsAqXUrNkd+EH8jxXXO5rw0GYO1Ko48qkRxwVaKB77E/8aWU3+EkZPUbLs6Xyo
pA4Bh94hWSvS8EsfWxg7lhSZ7ZLDBRjmO6G4tjy0n/Z2t7txEQIsOLE6ew9gk6Y17i1oJeU2IZax
Ro6Wt/WyQA6/VjRMOHOxXbsJs1BFJAScHGUdbwi9f/vBbRj5XNviZl9GtgNKl0HnkBw9YyM+reOg
JXg6XYS1fQNlvHza1qnHIO+jHQQPI7Y7SYZPvRJErydpfgZXawgs3WMGjy4Mll7SP9kGpwRynkRN
k+FUbJYIr5wvJh7eXVGhTLkVs9ejIi996sm28HPXxSHYyLfRFpqjJkmtxNQXGEj2AHCjbyCVkGkr
HGnQg4lXtm4lDNAMTSlr/G083JvOZXmOabydZMRQDSHLRFDw1ZcM8eTiGnhIDRn3L4xRJRdhk0et
ltJhklRYQLBznzy3+Gmyt2phJDDg6nJ1MWpN7ijpLYh1X8Ewyr/9sl87w+P0cY1bVcCKoHy2wFW0
mYx9wEyr6BSVI/HNATuF+8O7Kyp64rA5By+v/ivoj+DZhfsrjc+vf1pWF3iI+bBBolTnPU0qVKRv
lbadL2RdS8Oo2gh3cbh0PwgPeOSOuyaqJ3cavC5bzwHUAcjXVhNtdykXZhP/gVkq4NQ9n9QTDTbd
hPAQsQ/7cc0bnOOQilzG30W8y0XhLFXbmqMC7mklSAPZ58yoGHff8Ivx5H716Q2O8cXsX/oFReBn
KkEEbyLdo2PvcjhZ3tveRjzRzlbBERmf/aywgZfr88J+6xMVpoJVr21q9vt2aA7OQqp8Yq3El/B/
W7nnZKvzCQSnzvm798r71kW1Pz9dNE4JbOuPT02EKSMQJkjl9rlvaC9Xe/tSQH0dbWxxK+vuDzkl
ggKOoxiR5PkyGc3z2FwlxGZZOK/83+iRBtkF1IERJY2ndtmV/hotfCy6qYQF1AuCp8Z0fblJaBpU
Etd1GzpIc1t6L04MGnlbfLgzcwAvjhBEwuHNiH8kQqfX97ZE+POCB7FMoETFGDbnvGBKXPJYhVj/
Y7LxCYmbrLh1fYPTe1GrEQAozjmE98gTIID1BCDDC8lDgtpFgcutzlX9zcC8nJkEpM0NIBeC6YVM
3TzJyox7tDos/90b8FpLxSFxWzPOxWiVAUJIMz3MH8hyjy7EyikYxRpeMuYzx1TIkMBrb1EHH7l7
CJVUBWMrTv4/a6MMnCTYxcmKtCyvDLZAFSNC1XAnx52gv9LJjDiThB7nKCzw2PmHy9JaM34gLg4i
2rgwlW+Mmnzv/mky2XZOAdu1/kNDqfwT+eRlC3dDO4E95rt1aU8fAjcniKsnzVKsWTTDUVJifYgU
E5jihhbgU4GsiICf6shyari6882fOFwC+lWVfABeH2+rjLkVFUedHfz/zixAEUQISbcM5GAeRB4Q
y10GbX1o/Uaof+cvQvHcmzh+wTEcYMqXM9PVFlyUKx9VPPAYnfoYtlalD/wx9viB1ew5/c2qTHG4
mCjbccd7PfvWU8pgIjxkrZKtdVddFUh3fvpQfQkhRxGIQKESrmRrPQ2AZmhkzXR0r/i3a4wDG3X9
V2H8zd7cddxG66aSt+r3Jsn25l8WMiIRTTcQUPjUSePVp96FbKsH8cp0lbpkblbSbORsAJ4H0P8p
EdoMWxHHDZqQuYWlb8ksgME3GR9xvUjpoQYCOLegwVS1HrYyejflqMkNC8sb+U0jB8yRy9G33bKv
ZGxwKdxP9e/qAAHujtjt/xCG8uCkkyNzlNSLwSaH1J6Cq4yIv/BcLx1Y0bnmw3+wRT/QA/xkE7Ln
n3J8tyhH//VWan/D3BEZJyqGir7xQVGesPKR2gyO0/uMKB7xu0JigJDd74y8Fw6VvJAzkYyjHA3N
Xqo5r2PyrwwPLYKvhQH7V/TVEp0SUbS6NSqZF2bKRubzBmvCOpr/UXSMAGar1Oy/9YepDh2XWSy1
oPauRVBiRMNfh6poKUheuO9VdTc0eNgQnwAShl9Ejw4fjCD9kGLAfR8YV/pMlverdKRrteVNscdg
/f9AgAgPh5bza7h03Gj/3bYzAf/iPTTeC6AJy3pLwLFXIJ2r6zUy83skkyq7oQ5qAiEKOAvbx5Cf
Cyq6BdjtnOwF6BwTRwHl7qGt5FYhh/aWUqCnUbr00nzibWQY7mkClLO7LYmuI7kTOGF3D/4Iij1P
DmMMWhMEVrgNeFOwu5VJPSm3V5cFj93dvisQLo0zd5EKdSKfRUgPM2JZ4wIXahP6Ub06VAmN2oJO
1eVmx9NMEeMcuimvmptf/+LKd2uqOxUPYs0welfmL9v/juRUL6sqSqpEgzEEVVJGf1LXIFm7w3vv
K+oWhOSvZSNUqWFB+2bbsj/gRZA3D7n/x329e3UrJvc3cUN64InyLDp7iRDtm4o8rkLubZ475kgh
k/BSIuGPQheJNP00u/ShjJK/Hti2Cv3cRtwouzJvQY5krgc/LNpu/QGUNnk5DDQCsMDYikaMhycl
Cn/mofc/Jfs7IKES2rBrch/Nfjh4EJUrMBdaS669wfup/c7YJ8D1nA/HBsxXof0WNEORgCyfTtme
eiWtEpJ3sjDatNKYgpcD5F2914eAiZNCtCQ4F2y6Yl7vEtjrqpJjMMV8nwwFr6/ybkAH3dRXK3Ux
TOWEKeQP3thdfAXDMw0fiQZvjMIYmGetAK28O/r+Zl3BkpGSY5ovVuf9YFGpove9+pG4iwtDU0ZG
rsBXtd0gpwCZyVCelC4dSzupqCVOUi0bVKZpccVPZYoRWH82hGYPcnx6FS+ptgbpjjXS0NNyZeCm
+s/AJOs+JL/f9CTMXYvzwuL3wn5orkPU5tWUOnCQrR2jH1QBaUFdk53lI+AlSLjX5imhFxSRzjYf
O+98ScY22kk/o+DMEOTH1uO46l4PTiGjCZXIAvDF3eAaWeFyijIMfWicAMkgfsNsn9nHF2kn5t5s
2IEavugH7h/WvG0ZfIybLSNSavFOUpyOaP8MWFda5+0sLPc5d6JZyK7jE3lbGaeQGjB0FqFbV+Mh
bMRbjbhmoUiXtDHLm09DQo+dt6IKXoOcfT27i7+FDCR3QJiHoOz4GDIYUXaSxPAQ3Qm6hu24jjpF
9zSfSUlo7S0eqRhEe0zV6vNLlTn5JHyx4wqpColRBLSpt3+dOKkllfbPuAxKGEPPBTBJK216gPK9
jK+3KD9wqUphL2s1+PhnR/OLCpWs75Vwtm81GgIDYlEyCII1b+GHbQkWDpvUb0nEYUtFdAvdjNRn
L3mOZEuKrk2A6WsA/TFU/gtTmtgzpgfjGYAVyFQxuKzc7oWvXvuz0/vnNM44cBAUphG5d1FDFYVq
6lZMNdibD2nVrkBIAhjJ5hqczNiRnDsAIBFydYBO5sfhc68eZ/s3dOKurdIcMOz74EX+MdLKcdF4
qEJK6n1yDhAUN2i/fR5UMXCC+QXN/fKHj0IwQ83UecqQf81nMNPu2Oa1UE1M1cu9lRgfCzU0IqJv
TQJQQum75xkWELW/vdq3NTdnBRKUfekv1G3Tq5iSM+BHJS/MNSz/eLuXPKGNQyvesTM1vgZWk+zw
d5XgApeNwitPfGtnHCt2Yg9doOSjAjDucHhAbZ0/BV0HqPToexF3oRojgbZJglkzQBbL6c9dOs/J
f6jTGoVh7vtMYf0PAuz836A2WER60cEhGQdLdlHgWs7gnmg8/+1W563jNOQwgJcpjPlgnMCX+KEP
KMYZdALkVpaEQ6m5WyVvkdcr9D3HbMS13xYgTWDUvvEnxlZ9Lyg33pQ1k6rP4hrAJcyr8QZ9o+To
YuS/0iSCk7ZLeBmaL0yLacQd3v6a8/U1LMb366q5THhj0nlbCM1aFR5pYnTph1qBuhPfhAQiNBad
jm6Rcz5oiNa2dDwyeMNt67m+0oZ3Bn+ngbH56LL+uUApqXHv0dGIHfRfarLuIsSLjuZHam+9vGDr
IsCBNfFgcPvTlzlcWMb11ZxMiJCevLuaAdjwwc0mZ8CEbyI7OcOkqnCp5WvY29BlrHqVbWXgLejX
RqWr2XlbNuklOTk6jTaypPawvqqyWjTvTip0JQ8jPsl9q1mCd2JQIG+SEoc+BgYRepO7pc+fN31c
kqT+2ALjvtSLc8iGLW3t00K3W2MhP17FUKnV2fBxQ2YX7hz6fHnpsnGGWJuwXNSQRzXJPfBDBOme
FvSpTnM+/MIr54Rw+DNCV9eNLB5stCSUvQ7JvmnpiUkYDn0ak6zV1AYwt7VBctUSAT9p8BEg3dH2
NI5hFj8iiHkj8DuFanYq5zw4e+1Pbxl/sYIg2TYDfEYEJ161zXd5CaKQODNesyr/IAfNOpisLXMC
tWsAxQmBG0X/27Sd6a9hWJliTC/XRrQIhsp2RJ4gEpIpzl4doJ5IcuyG0niXf/uIkhul3CWoqbYB
2Fhu8wJmN5mOTUXM/2EH6Gz/081c1ZfAMcocIFmomEMLXR5M7GWjuR/p+x+4I29Y/WzODjb09kMV
ht2HIbxHUuPvVQWTYu0O4RxsY0sJve5KPO51DUnl1t8VH8bYiOlVt+jarDYnOJrSHtyV9FWA6NcM
qm2fFP336Li30nVpXGxtnSmJqNhKWuS/yuN2wMRaBX4Wat9hmNZCu3Zw3c+F9FN4S7WAT5KfvyTx
4GBpKL30FE0l67P9SoG9/aqMXF3O3CbY4d9H4LWayTCOqlqW2owFjt6wH56QpS+eo2mbkcluydDU
h4GujEY11KFkORYWxgIQeLq4JXleCtIdRWFKJ0//Qghrt/cHNN34Zjant5sshhcA2qTT2ap0/+Kb
+YiH5HsrdU8YmGi4FugPC2hhsLVEAk5AIOpFKZ3+Yv5HqLxcH+EnUjckKt1LzZoSlw6v0DDx4nS3
mY6ZAko2rTBPNDroCyOhbrfMXr1yjcmByWt47BWR+5YFXNgVRejtFbgCvHk+2FLR6KVHLIL1R00l
Bs65+lv3aO8dV5AmiYuFW5/5xaXkKFgl0ntpNzBNwU7boZV7h4M8CizC89Qmn85D9KHq8as9RmEs
1HXiF7HgrSg5QFEQsz4wTerPYb8lh0w7vOwsKDIApB3WSHUZxIOVV368YZis2lpJksNPtTcLeu+d
ZzSpPKInL2KdsxW/1s5XkNXmetAdZH+UXeRz4gifXeZ9bBqCtaS9fH2Er50xRk5t2KwtdlUNoiT5
L7A3EsKb04CWQtGOnPhwkif/SNmXApQ9Up9AyfMiUvOKNluzXaQeuAjLTY+pNQA4BHvxoF+Gi+rt
p30pReDaUFfP1uhqJdLM1IM/V/pyD3nrEWf5NYtq6oFZp8IMb6U0h4DK0kxdhGZ/qJ/ubr3hvZYX
ZUJUsiuG9HtnTY+3QgnEs7Yce2zhPI6lAWBsGnFIRIzZe1k9yZNYtvYXowPJLm+goW5n7dfGAKSB
/4Zy3GKt05xGinboIhtUl5HHbLlaszY+eUUA+audo6Tm0eWrH7hOGvYYQZuQDP+R84FIJWQN2+PS
HuXVy4RxCFUh2Mlp+JLpTpAAZE8vuzpkrG2JAhHfrqCZIohK7VZ5BGA/lfzj/BmR3B2jhJwv0k23
Y1F9IUowT/7zu6kxl3mS8f+/9YM8CHomeA2/sngYsDeroq95iXI6MBiWXISfCxh5HdCJUolOcol1
EQF1+Gs7+Ab2B5YCUQcPA5dTDoyuYMzNcw6MU+KC57HPYIEdbnYBY3LahuFHvoeDgHXmM2UPe6ro
slK7QkaQNVMTcEc3u3jvnPZ4AIeSHu9rZj0z0ST8Z1YJjGiDzuH+r2PFauS/Z9wxUcIbJ4NO11fB
0tfL3a8dXD+IbWYzhl9xIeTBtfgsmay1vKZdRLfHuPZdt3rTqNnqxoxIBrkodH1TQHNxEUpGuKJ0
RcOrmGIi5apjWqfTQ/ElYhq7b93gcbxuKh0Fa5Gxx6mJKEWx96C7vgD/38zyi5mqy8HasMPNfTEU
5dWDRsZIokxAyyQgpOhMNMRUkUZOWr/UzFX5zPQ6hfefqnTvhcz8u13yEvpKigUkR8t/QtJC6ukH
J+TZu0moVzDi2vaaZzWBhPb7dWSaY4fGKKYbakuMNIfJYwvvnVfZf0WpF5cR1rjcSApSelslQ/XW
fSYsRkVIzE5NA8cOeffcogoN4XhYr7Pd4Z4cuHRrdSpEKHAEYMr3V1VRjjxUbH+oogNaq9jrAzBR
QFry2Z1Dlyfuz7zbC2x8Fyy7hLBVSVUnrcTRcPMiBs3nTA55owD9B83fvogtwwPfWDqEt46uz75B
pc2AihEnrQjOgGvyLay1T/Z8i8s23iCtOe3gWx4weaa3yB39j7mvt/DuxBu7qRxM7bwd5/y2W3S1
8Qjp9fCsRcnhG/3jbS90Gb6HW5rhGoXdPP9q3a0YRF3y9KnjXJEEpzifAUeX4+f7okhJHCKprW0h
P8dPYz3ap8Izy5F0qFOgVJoKETFsK7sdhppRko7gf2lFVzkH0tUac7ExjjtFzlI4F7XAC89zZ0Sw
FvgM3Wrm17JelCOzqYohDT5+B1L4PbVNVmtNlCAxTIZyE9r8LJwhKFhXWo6Pfjlo0WkKbjEWl9gm
fNObx0k60CVuGyOBghu8I5W8vya+Iz0K97mXUEs1T16YohI2r5afK6KQMCRnIMoFIxq9myzmB1hz
oz383T0MmSXKQfP6x312bjIKe9YI/qsUXFga5cWM1PFdA8VEhvZ7VulWW5fIyHbaawu2GI6g4BOx
cHQ1JKPC+tB6z0fvnvpyREGb8M5GeTSIOSsaJyzDXa9WDtFpsYCRvR+HYS8eYR8c6F8uc11kZmdT
3G+nG2BwcEzeYYHqVWqj490RJv3jKN8T0s7FMK4wle4OAmZGNFez+EBzOtJLdcbjqlp/YejmHGJb
UWbAjwOqH7tmwKxgdJZXQn582jg40Er1uK/5gPFVTgsA1aAPL60v2WcRYlOZY9dERvyKKCkWsk2I
XcXcLNQDzFvazPP5X2zzwSvoVSNedHDdOe9rxVpfrRBahcAEi1jYMKaKgWgeShqoLF9bfIuCv9RO
sGCameyaX7na3Q+6G9WA0DIqnoRSr0j60+gzF7VVma51gh1FkUEJE628LigxsD2P9zP1Lp9us6Rh
yE1J0Jwwx7EXvLm4H00g+loOE0mXuDRL1MWDX2+UYmcPuVb1w49KTiYYLAQ69YK+W6LFodAzGvGb
gyS8RVLxRFj2pS40Q8I5kezuVABmXRlK4OwmqJQtyXQtA4avIZfMQrhonE8QbntUJpjXR8kbCzuX
P7tz3Fp6YOplRc46AvqaQ1Wc84R+es/gm60XtSImP07qijZffihYjAPVLoviwvgsUsD9aYrPIMD7
dFzfWPKzPzSrKhnCZCMmbIUMdpnBTY/AnmL26skI5ZF92EfqYl5QVUnYJhF/9k1X9ST/8BlQgxuc
xEWfnPC1LmjpvoklkaaUb2yNCJtHL7tq/1g1U8bJaqZ9KDAJLfjTvaD/tOKAOjogbSLdGxcvVMJ3
p1M7mcI/tLL05n64XxPJ9clAQGYEJWpFfGE2zf0KI8J6ESj8AyEej++QTFYkgOThA1baortBzAmt
hxnxcFKJZjMiFPjCkcK5CH5YBEof9zWM3/v8QAornz4gd2fLEXI/+kbYcNbvozLQ0lBflA8Qc4ph
omOCZLluV0YAOZX3/CBJRqKiYTYj0Vmuup3vG3rzqW7LfDrVds3/+GO/r6RBVu+sYP5jpTo9iGsW
bO59immpQk1BPhL88V/CM4cxR5Z9ju9P6FRwH8hlA1IuJDONUecDQGQJL/IEUrIU55mAMYfyElNV
bs7WPnOIUwnVUIDXgSwXpXG/4aMluYj0KwMRdlDXqKVTwS/A0iY+4+11gIyPXA2SoSrBJO1i4qWJ
0KDBgizyja3+eRqUISB+jmIDcYMNcFiDRyMEAaq5Tg2ojh9rz/+Q/GR6q4sr308ZhZ878nXRriZl
huuflRCZadvHZxgUkKPW8RYT6krr5upFRE0zxn78wr0HoSheBrx3q6b4pEgEOfKrS1dbg2CvncOW
E5D/9e4Ql6CAHOxg7cYNh3YuS5V0O+PqwZG4J/N/fu5w49zAhNkeqSXxOwToF7w7SsMWqJGc0QOE
+skNCKC+hL9vqcevwcmbH0PTOD2b/hO7+uM9TLEJhNabtvOoBJlQpGfJfbIm8JelVHbiGobJemYJ
eVMJg8RcMy/iNh9JVfnP16hHDVZqUdpGyf0lEJ10cEDmK8VshB9Nka7paaAJnj1VBXD/d30M1rnr
OB30jeGhWJ+rpiffCvaxwtQjpC9wZrehbcwu8IwXrF5BQHhZjfoPQAg4YBcWfvs1NBGeXc4VVoQr
25z8hQD2tLjqX5WO3NrwT6BzX3AkIjRPLmHQUHofrmcsrCKPnGm2RghXMQeB+kEv7ESPeoj/QaQb
kscTG7hpEC8k7ci8rzPCZAuu/AuTC0unMZv2NCrwMmj8P/tGbW0gvmexowXQwrPVw3i4BCaX6nvM
rjEGOVJZY9jlc+k9UVJ8NlSusVY6Y1dT6Ox743YSN2A4sRQ+H3+O+8c0rVXeSOxf2pLkxZAsbQrX
jxMV8Qnmt3ePswk4GwiiFnCUpvZrYcPVwD36HFWvAnkIrMIgLG3N9frPJoJhHEy/4nJyRxaGUfcb
KCH9NiPVGhesmYcIDkfEkTWCwqfNNMG0rBdI+JU5WehuZScCbmsI2jPkNQqHEMSO3SufopYnSCqs
sCJCMq+Lq20f74KuziYffTIfjKIpP4gddtLCXBU4givmDeuM5QD5ysW0KLQA2qz8FKDGbUFW+uXl
PMsqS4CZgBfvCEMBSlcODiX0pedELldrYtNFvlDK+BXK8pyTXtjwtYgD0RV3ENI2RsA1WnD3fNnn
V5rFRPaWZW1YaJh53YzhZZhRp0DVP6mxwabJivxWUcxzjTJJlV+/HFTcd0aj8lKQXz/4guOjGo/4
uvXLLBar5660Ly41OUkvAaqdqti6aiTyw5BYGUf0C/uWBadhIZzaKUxHmxCa+ngDlPh91GviN5xd
FoWDdGUH8N9lqrI9JlmuP75JMlugpExlxsMlm/vNwlHy3bbSGWxRp+cCi70/OENVtGdbeD4hF6TX
K7I1OB0LFqFH0VU4oPwmAe7O0Po1UJK6gasWjxmAtBZoDPWWioCYsa08zsc+aDAgQFgYOvjo3AnA
XVTXhGqTPG8BRE8XHBrMk+1CPN07cm1ccXm0wM4L7w2/ItRzrqqEbQcE256gVkcTx+QDtgzqgjd+
noC6F2Tf0Q91NR6N5u1TdvCFAFqgVjHi3+CLTyiRcNl41VNgosw70IflPP8kHS7+l5ItSv7F3iIK
S35AvtFwL0AXLziitImzDxauOb1DQjYVB+hSc8TXkaTUlVUmY2PD5o8xqE31Wwy75pKW016ob10E
qcBOVkZbI5pblxJG43s4rh7tV6PviqEwXl5IXjAyBeIJFJYVWuAFp5Okqsfk2AOqPQrKCkkrKRKy
0h5Kamc4cyvnUCd0Y0d8PAefgxJVfTc5B9LrWI6dOiLPafhCQee9S24as8mDSzzhesydJoAzc1x0
E0g3y5N9HSzX+48eI92JLvk7XhvQ30aU0DqUOHu7fQNWJ40UJKUbMpi/T7SrCjw+Fqz/zyQoKvIz
XHnFJ9D11xAU5Rkk807LCZzD3WaEbaaebPQjV0WQ62QTdf2I8SE4Dn0nwkaJLfaYmYjn2+bKVqXI
TxL+W9/b205F45Z2vJEuMbIOEeaI7wEqpZfubOSpUGr1owv0ZIjp7Tgz9hapvCurL12aj08a/8bP
UiH62leqqx6R2X1VuK4phvidaaYA5dlda5JjZytyFgD9/LUbPVtKsdR8bd1IvsyU3u1tr5J3GcN1
qCAmrO0R9pf16y99PlzCnrW+Scxbi1K17iC/eAZO6ZYcO8avLFFi+z3q2Kj5ReuDQ4HgsIKn/JC1
nrJw712lcCx2VwRA9DKjlD36OldzrlYthtz6wfF2nB1+pbiIFlcMGem1uicref1Rw2kOUJ0RpeK3
DevyWa9PGwsCARgF3knaEHrKNribPzLDx/5QsmEqBK/gkkIHAOmxY5CaTyCPsGix4mbpwToH7DYS
a9Re825yRLC1n/JG892MnCNzbRmOyK9gCfnQKXtr7NdttfYDFrJOEhDH5CAfSKB1lh0Du5jOW4vn
WtiDruFfvRVyFv7QZlQi7PwXis/WHr8pPXcvX8jDPWh6Pj0Agi++rz9SEl+DnxOAyEGoeNvu0Soq
AvE2fy3cx56JlKLsbhqAS3/jUbDk4mLJ8JK9ThDV10z/DA9UFF/qXGecY3o4HWdeQzhcTAOkCc/E
/0ipe+lK/uF73hsyxbPPdsgmHcIO3pVIOdI58Ko36H1nErr3N6EpUmU7cPybLzTd3rQ2V5JwC3+1
VsV9hvzBDdMMQx1IqsewLiZDCkjFpK+7S6UqSNpaWXwZVSX2MQiNXfWx6ihp2gr6WjvWr6Q61AeC
cjXWPylRKC/aKM1MVAMH5BY7O/VSc3EC3fArDeghZ9rc5uqSCVie0w5Tf3ClNp/I9lq6zSXIUXhI
rukxTWrAhtPI+16zvWv2QZp1jsYkrGWKyNsCfwFGucog3Ct8Z2lA1PMm7rPzPlMQyDl1gR/8S4wU
urPLMEXvMd0P0fqUcvPHSH7akL2Xl27ycCslGJ1+OpOJrg0D6V8/mTFNBWp0kuh73uDrSprc01L3
dAeeu2T517GfumoZGY3ixM1hzZCbiEeb9+epYh+cY5IkcDSaMiV0BXI/GUW0f3dzxDsiT5j9M2Dt
ws49VElox41ejs5nLwmRuhWF5fRSrA0KoIB8c8tYsCEbMAquX32osWP3mNmYbZEV3va56EH2HJYz
N4l84+wHe/LPvdJZjgHMfRGTy7GTYewhX+mPQmiwYAiy24c8+2zI3LFMDlkYld0KAIheKXZI5kmL
gSLPvHSHD5jfGRfyCza0Gp4IJ4segKmNS0/hxfZtelGLMw/TZLMSTQ7sqvSWLXb32DWSwD1zHzpg
KmnEwQ0S79qxiQimrF8ZVqTwSdCxi9dvLz9tfjJjEr4ENdd/fz58RaKyITzhRxy2/61jtxGQGbu/
T4TXOSxSKBQlwCAWaOveSw8kUzbmTXVz8NCAlIjdlZ91xvL1QJdg6WlIErk8pTNm0Hh2fnM2LGo4
M/W8UwJUG4NKVCDPLFHTP2AA5tbKX/IIlIYs2TGXPR9BX21a5MjqXxYLx12UgCyyudF9RCOuFamS
kTjT5MuGnZ1ok2x9NPaWKOwB8JTlm58QEHM0dYAXkBnMkJ47Z/EHaDeazRE6AGM64+91CnLzthyn
WUEeg4J/uNQmkujw14ph2tXWJMjYyKi1CZKBeylOqzTCGpTr19ZJXSCezeMgUpevudrgyR9kG8F/
8GuBqct9TRibANArPkr+A5RWYOtQKdMZp+2AISFPBagVedRewoVRiyb+4Hw3LMtoGo3WArQSOoNA
vgTWWuGgqBni+8kEYud9M7tQt1nfUHk/ro/FpxonpcTdFkWvz61kZZ4m7ycFGwczgrazt7c06cRI
TWIcVEZF7vco56YT2HJnvzpOuc8I/lYr1vF+HNL0grWrA60PyHdf+3Zs2zXTKzdXdV4zwd7DQRdR
d/Naaw0Sawzc8tcy2kAlpcd92OsEwY6Zd3OEGd0s94QkyQFanik3UeHHcZkfpJZZvNKp9oRe2IcT
EE790T9pgkGJBj/ck3BiNjfeN6Ef0JVLH8icYrfYFobrEIHcFf/khLPfWyFXUN1ixUCeIMCExZPs
i0gaLvGvxjPpFYleEzZxZUAyXTa7YRrtEPbmQIgmfPI3/kRxTk6ugKIcd1ps7Dw+hH6EMn2LPy99
jLzqTOIJsmpz8BmaYVJocCQR1e3Xmjr/tX0Pjf86l3t37KHRny/0VdwE5jXxkOcML3BwAAAmVV8D
7IRBTjUuxbnGejT9pqK22nZV4SQKZX80suJVJEChg1XzhHYZPTMJPCXKWBLpE2F/nwg3YOhEKrnP
GdhDhdVIWlxx/a4ycO4wOZjgL3SGzqJB9cGwBZWh0v5imr03B+7zLCkV8RF+VUond07te4ys/cAm
SGTd4rJoC+Lt22vBkZGGYRS4qOMrUGCrqdbDHuFp2wSAA0b7/YaQSFjDTcsHBUEuHE3Cm2Zq6gNn
yjc8VqS6ukLg5rCvFrlcOmgsVKv/8ZDelj+SBjwiznh+OCr3rlcDejIWC7UWHeVyRCE+ddWP0byC
rPMaZadERD7SLOm7spYX+DYTcWe5KUx16DwsOAKMZQPqYSthyqkqlKCPl5JvYLWt+UVMyRAarBef
TdKI4LBW/SAw3Et2Qgr1FVKqRH5uGSFnSznB0WmvcwL3EVyK8vCPzlNPAllbIvjX9/RpAD5oe3a9
Ta53h00mj2mVZnunHWm+5eLwxBqtaRZKgyZ538pyeO5F3aMNvNbz8cO3+mIwhnYgP//V32ZeTTGu
HvuG+TMBCBb9KxLof6KdgP8XU7b2hBRS2s9rMcH2QJFoAFPhGpjS1tYjRImysUHYv1IZkZevBIj3
5vN6+sXBIpEZxBjAvvFoTOZCqRGv5B0g83raA9EWlBgGxmXw6DD37c6BYuESvGAMi5gYOGImaIrM
GwA+ek+yYfbQvwDEFCiNTBuAwv4tBC3qoaTL9WjwghoReP3XeeFlgZ2X5jzeDltpzOOtRqgXURox
6hNu0xqJezMU8fg7+otcYeYPETDrp92VK8oECFFjlBAMGRfKcP0laE1GsyQbmAACvDi837EKn9HI
955KejGQod8w72UfYVa0gbVtsQawJ55cb3JxOBHvanpsTnTWEBsKGMmMJBX9j6zQdwi5uZTgI1He
Y7fck3SAHZ1TXcCL4V/5sqXtttsx8uSsAHul6vEBrai+fmW5AP+53Xz/LbvnhHWG9PlREGvJsCwi
3/zW27q6lzQmbz4H7Pj0O6mePKCYYX4O/R5MQdSMpgxOV1dt4I/eWQEn0ge+JHGd5r+4D5P5X3TT
8iSDUbPwpOZAPw6wUBmY4gvRFvHieR/jkJ9XHESphw0NEqRGpqW2aY9UZ8PQ5zWLY5CYzKuD3QH8
bW3fW44Gq3X+1RSiivFRcavC2o23062o7HfzORTdYRMUGQi9dYLYDQE9cilgM9C/rWeLmN+/QSHA
hMcQ1OjNBGRys69UgbJeRIfFttQ8megobCR6UfTFBDbA3QDGT9FSvhEc60/bJD4S/6yvtoxhqjir
XoNvM4BLkORe3CsRWKe93I07QSNLlyjbbi7UU9sdba5wmAvBM7+SIdumxEkabigdi/HmYLKxKjlz
ci4JGl2T7DLo8MTQqJ02zoeU8WUQd2pF1eMboo261ZOyZgAYn7Yrtas4mLWHFTvUi29ygAsgwP5n
4azk3VMKTT8fLoaBVETik98ks7CJmKS59ZTJ8oXwOjRudzoKy5cLx775pfcQZPLwQ9G0PIG8Q8wp
WGcMuVFpgzSHpg3xHuk5njwsQVjh6VzUpQAzFx00MM5B/fhVBq2ubOWE227qv9RCtl7rEuFCQ+Bi
aMtz3mFlcbZVWtSw1YkTjt2fsBRWX+29bXqSCcHnXePoaW0qGvIir9BJw83VrHHoQtkjEVNwFdCv
y4EzQpWgOB9Z253ZitvSr8DM9uY9IaSOmuZKsARKFhNFcs+kV3m0vdRQEY5/FbeqZozv7BHvBIOg
fJbelqv9rWvNg5kofzkLpNvvYy9aIT61VO+riy9YGffEP7j3o+4A1Wi+m28EmIhwL47WfZGX+WDa
XJFxceGVt8VW2TP83PP7zufvh2OZb2s7tr2pkq6SgEFxZX0Qnlg8vCsspxJF1WFXJvqrMjFBbUrp
sQyjGKAMhYw7BMVgILyAc6MY0WBHTDXBYM1xp0hy2yjm7CFNzAlyWNJMxi7ZZFhQDB27zl+RciVv
UQAuxTqLQdEfcWzkYh2xnV+OYoadbLo0jNtRndwRmP1z1kkBRTyphX8wZx8ZGovHt6MtL1J5MIzt
AZRVbC4zLjjqUBgWAGAb1JJCQMeTy3gr51EeqmRfhZiSRcUZg50XxEhb8MWloUEbMxP926lxKaxN
akPtgGXSG7FeEBvWj7uANJoq+mjawIZACzRCwDvcqJCOXPZUG2CsdyRDNR7zrBY9Q9do/6EAoWAB
UZkRUlii7tJVCueLMVSZK63lD1IVM4NtFRLXc2Bo6n55UE+92ZUzSqVY6TrlWoK/AN4LPqlUIcCU
2QtJEBjz1XH1THBXDvonw0ymTrmC7LR1RizsF4tgAJY6dQFSYnjZJ9AVTYdNaiQGYLiXRJejKj61
PFSC8RXxSw7MWmk7o3t2FsqUQ9sHU+KqCYfHwsGAR0016LrW5m6clHwocXspeC5iwj+hCOFkxr9o
5gFAhWAXwqlQ9C55YW1Ea2jpsC34Y+aZtuFFBR3wNIZFxN3VQV8OPYB651iZgDuuvqHTu3zMMyAH
0p0uDBjB4t829ipwihrqRfgdtWpoo8Kw4Xp4pDB7MuTN5Bvyg6jgJgge04u2c2I1DOdtlDzSmD6A
K9Pj6XfTKlPODzlqk1TJc3SfztQzo9B7qXPhE6K/fDDNGNb9VPzyk7kOYKGed6x2fAhYI+6Kozan
LbhFBBdnU6hkqx93AMFovl1zeW4iKMhwMy5L4OrlOJ/ZB5gYlTwOR0a2flDD/9H8FpY9ntPxbU6p
SfMOYKrTt9857JI2SkYAenXECArvLW4MHR7ZP32z7LWCreYAl2idXwXiK05cjbfxu/lXc+IRy2kR
3p6/0YYnlTLikAS8wfw8W3/UYu/2CxT7kI3jsbjsHW61o+Ux/3TPE0UsLTA4tqA3ZEbgqFRAG7nx
qjDnmSAgCIbqA9MN7sQxYjYdE9CYWyUHdjmQru20q/4iWhJtYySoThoP1E7UgnVm9UBKV+oSsKUA
4LKrJytGv/m+jkam/dlSLuPQ/5eXR0+mwQNL+ttvgYmEYE7cTfK8cyfq+y7GIjY2Upq4J+g0Xo/P
cA3IkLkG8CO7eHYEtyLFQS7uxqC3sgnM5DanFTCz+N0muelIrKtNN7KzFpQzs2txx+FcrknX2wrG
1OiGXrM9R41yquRzP7gGlJYaGvDenNJX+FaqmJyPGs7whr8QiS7yPBzRIvDbBqUoMVm/222XznNZ
sv/UJKGWHG2nH3hLU+o6p1pRs+81BVSBrlv9ck76KscZAfzx54D5+acb6pSFFILhLmDcICzTaz3a
FwUX9paHpkpFg0Ot6+ErE3I9HTkjRvpoLHhzH13/3HomGx6oGhO9BzUZJzen5yjqjpNcSQlGe/q9
fq/WT9pzW2mNxcB8jf6SJjMW/fWL7V6frlClwVV8jTx0Tm6sn8xc/CtliEny52OqGNAKSt1R8m4M
Mo4UPCOMXgyXnwKnNi9g+Wqa+V5VMFgPhpBTt1dxw3JeHKAuGW0JfcovggIyr5eRuqR9kk+pt5mB
jNOx41wEKy9A1ziO/mNRzzR0D7Yx2W46n92mJFduSMd+iRG3vAlCb+3pdPx22acEn2vFEepeb4na
O/Zd/LmebL4taVwxnb/ftoyhRIzApPswNavxaNNC1cJLwpr7M0yQKCs7Gv/Y0Wr31bNEFbKDZ7f3
BqcCikZu9YKCv/NRuZAWOh0hzw8Y+m6INbYzD9jA8aGaO8He9SuolKTBGeDZ2e3ooqQ4xX1IUlgX
Bh4tQd+uMuoEGPfc0Ogwo9kfqTTzTWI3dqIANC7Uq7CT03um3+np+wynLqebZGyYKbMEQ3JheCYD
H76+0PHi8zkQQY5A7RQmftJduAnkx0cBoN8IMpPkejjfz20xYD5e0+FFpOYXj2uAfcxW8eM0xpwP
gM3/vOpAiF7SLW+WF1icMdEg1pOVI65uotycQ6l9/CRwInoofSfJcWc/jmoJLNKZ5/WPlJFDLIsx
yt3er+lS0wPCw/+/UcbaN/5DDyxa4+k0r65aH7vuaaSiGmq2AdAxArb423JFcmHGx9NFlFupp25/
d/b7UhyuZVuhteCRCacQvl2khtMpv09JT1YXZen0iJLIpGLiwuBsFmJwMw8s/dFzU6xFfV6Rxr+O
WqiY3VSUDe25jxxR2A0Aptxvyh20QfjqDOWqJaIFATW6Q9xA3r7I8xFm9+MdZ+MS6A058BlYYS5O
7iNwdhjpC5EAGug9BFCFK80Q3luDK2OMRKhHEJRC1djB5f2gIHF0Rt9/cGNhGLgTJYuAGDUHnn6X
8/m5OK7O7lc8F/wgPLCLtoOyKEVvZ1UOf9fGM8A2kt4CqHNFIRKK+Z8v9QvDu5IRS3giRTiYSBxk
d0Js3cHJiuxGyZQSIycy3ZybIZ74yMSvrL8UwbTq3ayZ7ipNKRdQAyFMaz1beO4mPvg9lXZ91eaE
lEeOl0FogJXnyEH1r0la+keLmWpjURqCClXdBptSJdHixiCfd8/S5KN/EBlBsL2qsbO/b/xDgD8v
Gv/mUk2mHTF4JOu2fPZu0a08WkpzrGXzbaROeGWoB5SQkKaB4wby4EDlA+gsOUU42r2RPhq79YKh
lMJUHIPlUyVkDx84/wxXfPJg0cn7KU5OU+sBDQsuwRu/TR1jQxkVmT9pMK+aIakzuW7PL/zMkVyG
9cff1XQ+q+eSTSy5h4rYoWfz3gFfwt9yGmFSYcS6c90k+8G5Ic1I5EvzG2CfexjfWG2O5v7Jo/IS
e3bStZfm0h1OGOI9Yc4/CO0KBfJJikX/vQ0f+OjFRr2ZBNXYcvoxeBmXup6wMouwWEjqY82LoBLD
uae3aEIAl42Q0e78CCcL/bsu5uVj31mGidwDggMkm8G/IUIXfDN3DeQ75BxTnjrMiSH4W/acK22o
k/4koSFp/gwQsR2DBObHt1LtnXG/0NyFO7222eiY9lNeNi/n6GmoMd9c7t57CrJpPfJr9nvXol3R
aBXwqkxbHg6GOtC9qoxSZF4i3Eej1UpcAjh5lSspC6t+A+imFCi8ruh+TA2HlHoYUDiO6LabyJUQ
Hcai9bG+KlBDU9OT4AXgO7Ypcpa+7AE7+4bm5eX9YAMecUIGB8SYua7HpR0Zd4aACLHkDiNFdEv6
gXiWpTxxiDbuogAP/5HZ+MRCWG2MQvqnWgxUNb6X2Cbw2w0ft6ge1TQ3LyCAk4loyxDc1mmpde2Q
HLuEQ8FcLPl1cdWQhmhZPEvPxWw2JuFtNj8cX7sWupILqyIUqKYsE+CV6Elh+oxf00cSrqvy/Glt
JDe8VJSntp57Y8wlB8AW1S/pCSTe/7drsCum+EOBMiEfiLAASS+p8VbDDLpflM924v1ZGJSDE6bq
/5Q5qGSGpOKUs19HTdo2K59oB7tJy0tPAEW7LH8TOzC371EloK3hSB1GqUOWqoYh7I8nJaloWmWQ
BXJKt2MXuAfzb/R7C3MCJiK9q3wFnqaSYQXv5er/0D3fyQT3Ng5aOGAPxYwqYNryaXDbiyaA/fzZ
VGzkFAq5HCwbdbkVDe9+ov4FbVaSg1VimTULdHtuyJ4kDVHKe+ef6cRYiJScS6FZIfd6wxhVNkNV
rPm6WHKj7RZXyaY+ht5JkuQj1pMjY8CJwSeEKeyB7d43S0Opg6hD6dsEhsFuUDTuDZ580448hmwH
RZXaI+kgltgkQooIt9zNGP2DlHmj/dJq6Ua8xsW5u8rxrlLbTZsQ5x5foGKcm1aEn0xbNbSHUFxn
wsEtbObLsYLtjZhynnfJ4d5+/zfZgXTyvipAYiUgBg0K0atNRcqAuA/kvTifefoBwDxAsWGyp3Ij
H3kDoIs5qw0klZRY0FTIKOPilUVdgTF8u8sk2lGP1RRzJNV+aaEa7kaa4icdrhQsy61GDk5skcG7
n53NIIghdH++ZPYp6wn8iN9+lQXHxJ5uzvW1npAYL10bfAbDjxR2/6wFvL02Q0xoKZsVh58UUxxr
P4cYdZWVOqb8zUMCUA+B8I3WCt9AuQ9NpT3nmmGkCab2L0rDQtXaDz8sO475av32G68cQNiSYx1m
ksVDzRYo9Cq6Q3mm5KYwCBJ3VxluwMHv6J13VdJxuElhFgSl8s2uSAuXHu5ZLAp4xZVYNdkymgLC
ZMFzEdINFPvp70Yy4y7QthGF1e42z5qBNlOWxNL8Xdwm3PmJfp5gnKm9s4Jshc6b+gS/LBqLZCcx
OQoNforYoFRZ+ijDQVvTbXLP8JjxB2RFUo7dM+cqmRqzJHT2yvudyTpeI8g8c7l86UUijmXS3/au
IXX7nWZg/8c1jkZ6OU6ptS7/rU5P/BJDBB+JhexT0AdttlX0AYV2arGJYG8OpEfiIOLQgC+PX5li
NBMIzhUYA2Fr5fEmvgdNVR5sodBMVlSRs7njLOZ3FD/0ON5dHqm1xaW80s0uGGK6m+na0I+n+YAT
oSryXF4Tkl9jxPYLCxLnH+DJS2Hb/YqhEDTNnCc+49bg1m/RlZ7qWhmRWNenFSs4cRC8IlngagpK
QIh/43vS8oVjiJLlmAgyiaBmgp8YsFnt+C0fh1xAQglPenmaKxO6wf1hFpZScJ1CCtFhUZsbZS2n
6ylfFLluL9LTJce9AeyVTUOHG7SssqrA/wi86sh694Ui77iMS0ZVXiC1oM41R+wvxApETKtSQED+
VrL+u4uxph+8U7g+ROk/XUdXgXpLzqn0PVAjzz+jSZwV2/zzuz2hMbRu3CQ0gMZFb9Aok9F0NaVQ
9VgHQYN0dJzddTPoljqiseiIfzYiFJIL0Px0Ey+5femhThQKZ4CURTgIcuDPu6g8eXQB7YwZpidN
gUcZ5EmSgsWHkdPwGM4UmWELl4vW+VkULaEoP9Qk/H/6p/6Cx6DdQb6khxefOA7cAdSaRVVCJaZ2
2SqttwbOSF03FXOOLoAxDmVwq7lbd7FecQ0dI4/QjysINSh7ykHO9Gh2SKPWJqvE3DyHgTW39YhP
6Yh6yhP3LPMJ+J3FSdCo+KenLR3Utb22ErpDg+kOFM54u68h1vviky96GoHUBSx5EHDEVDs8odK9
jqCZHFU/gKnR0emMYiq/kDkJ4TUmxWdnoo5b9qyzdjOMeMjPUce0bfUAGwY1DcFM3vtaY2U2j075
Nrc5EAicJED3iGjzn9wjLNCoIUREqCe0DFamkYhtMYGmmqCUbE0O/vxbOzUHemxecd6hG+b+1InC
OUTAgAF/KinitajE3Co/TX3kNGgrO6M31iOEXbdtjYiNw6ajmZAgDrOhfXKwvXgICnqVme6TAhOK
4SQcSTgCN/pQhKRsiQmJcBxPL0v7P9SpDPpw++diOmfTyW5iCPnBt0C72Qa6WSU9D5nJzGD8q8z8
Bjye0ngiW/bepRuETyVZS1d+ILeenFYQptiqrwWchpQ7pBMGu6Z79hLfTxZ2dKd+37WnBHUSFiCm
fnFV1CfdH/bq4eTqXKMJ2LyH55aDyJYCY+b3bYV7kHQJ8XuCuswXbo2jnqnUWJCBKKFWdy2RTQKI
cjh+mMscCR1m7jJm7sicS3P5R4pXP6ZS9xvG+RlA6I9ZYnuEm+7n9O0bBl987Yk6ioCA7RhZLias
o1BqIm79E8n3fqBKZCXxRaQ6bOTFWzMkJ2bj18Y7nRWqEGXgyBm8wcugyEDgQto1u/un6DfAwbf2
v2ThqewqQSiAml8uxU2+0v6hZZzkBlF20kgwgGmktjvkUIlRv3k9Rj2eLWBDJeS2K6H7CF2KPI/s
+cIckuPqKTPkWxqjVKU3yiGlAdMK6dZVjtDCHiO7rEZgeBAINQIIN50dR+v6Azv+ZlSPNYGQIL/m
vtOwreG15UaQEmMgBnn6ew1jexYZP2oI21aPhGIbD92w0r5J7SzxT+m1tumeifBaQruirm4xHjQj
XfL9G7ls2kfVkTzlzbt5aGk1s/qIsoH7gWD2Zt1lQAsJ73A31PGRoDoXQSJgzAFgpxR03MyY52jd
D1QqQ0TmcavWQVJj6jkKCg9HPHFjTFhm/oSM2DnhJ6evzXOFRJQBvfTvEYj8ME7IT4UOjJnMz1SD
m2MmPZsVt4nIDRGCBt/QP+YWZiC5ReZrfTys8z9j6v6ghZIAomQbkS4ah8P6qC3EJ3NoEMWQKLkK
m9BdYjDkHEsxmq2B30BOVSUaG0hnvRhpAjwxS4tnaJIWA4OZKZX4zq1/0YtDAgvl1bwFZ4/5Ib16
30+zpgXm6sWElW1QkbEMC3Euf4AUJQXBQf3hoDrXZsfJE+bkBQ55qM84wXL1lLkvpQFnooWqySnk
eD7vcsc7Y88rgvtuZth43kjWmfFHi8tkmRH8kIsSjrZ9vFAn5ICxEcMRtZW5JtrkAt8Uy4Ya9m0/
EaYb4fTlZ1E/C4KjT/jldTNxHF2gspG0n6OC7OK22hjp55KxCkUX74ArdLql1W4Y3F37zvf31fLE
uF0qnvfKDFX2DlMvt58ZtBZnLTAgV3h+x/s7mT6rBOjF/jWzeDZSwEIVoblYSCNzTNSUW4zFLcBL
QG9KfkcqYcXiV+kxR78RDEKGN+fVznsObwKXvQ/RGvZI81l9v/ghPpTvTSlRy4agBJr1GA5mzFFw
mqw0bHx/jYGkH6OZ4MNsyDTA5kojk1fym1fZGSlnnq5CUvLcGr/phCXzgbjrpmf+IaD5I/UMLRO/
dZnTFhztUzPR+ntFyIhBh/iwgTbNFhB3eeyw6YU5Va51kJDzodPtLzkdESvMobHlFrO48/nzLidf
GbOT1m+gqHM/Gjtm+Zv0DzKO0Kl2hV5Phd2U423wiuJ327F9Me8veehVeqhtthC9aNVWY73+GtJh
q7OVjNlbOQj0RJC4C3xHZA8NHGOKXMQljy/j0yfYhLMcDAAlAbX59b3hjr04sO5j4AvnklkFBMMc
410LdLb/qlvb8dQ4vBHW+amBngt2Mh4ihXiO3Twe3fI69Mby5Xk+KsugyI9xgILGdybIrzLW8+Zi
CbMQ78XwPy3t8+eVoTZQOmqaarFgmCG2EDxGFAIszKaeXxbx8YNnn+xuolHl7I2E6hO5KFESYPNO
+xSI3KzZh/eoUqWjrqjxcWg=
`protect end_protected
