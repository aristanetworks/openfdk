--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Wm6YQrWwlgqbG69gLIHjAu52ahdUIlnQ7P7ACNkK2MfpF3t6Gz/jkBTvvGjZ3rAaOU1dNAtS4Bsk
6/IZ9qBXzzCCPnpC1lFj5jojXaLYfMvZhIoT7qsPoyWndMbMmEwg1/o/+Qw4Mj78YaYc1/QES0Le
oe//ywMH15xCRtWrMH0kbFQvu8HCRla2fMYLxhw5YHntH4X8VZcC1IjIQt12v0YIOQ9OJySjfsHp
MIKmO6h9mcobG0sVIu8h8SnB4O7K/9zY5iKFOcEimFo/uuQkI80ce1v/D4WS5FIz4MxXAN/TA2JX
bUXre7Kbui4ySEE6TaEwoeh2RiRT0o5sZzPuJQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="U4OXP51vbeKzpmteQPXW4iwae/TAj1C7/YMWmsyw9Y0="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
avvYZMYa3G/bwkwO2QPUTwJArWOyLI+1tJNJ8L2sdoGtob67pJVZTkzAjikjmfcE0S3ULQplkliW
vjwM5cVNg0WPFLRaOvrJKkjCyDV2ITBP0jaaPzB4IPpfx24MYDxKxemf65FJq1i25AnwnPjTflzm
OTq6VsZrXLkzJfAvjaKWrLX4sDj9B2XhtJp0HvwBplZ0Yu06Do+BlKQz01vSb+AigWJyduNQZC6A
rLp76F69QdGczXM4RU2cdiqpCBzg0SJxidVtZa04EAcSwmqrpH3mRLM3J8tk7A75r6W/B8/RJDqv
92wQ+Yq7AyZPv5XwtF9Zwft1TwKrW6g+JVz3aw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="jhbDQw82PSWWeFi04oIQLmGkMH1O7LZlKki38Zn0oIg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15504)
`protect data_block
oRQkxpN6r9NjdA07eKFD+AHDepb2IjUQcC6mCVDKFgNWWYy/hKLfBf5aUxnR13odwdGcPi0bcJTU
JZ5gE8knxwURM5hAMiuFiMPavi2e5AB4wdrhtw2Fe6q5ugJsW2aI1hnb8HDWbsPcnQyYqTFuKz4w
fDN58js+Eev4WjpT1FWUkVvVbyiMUb9w2+XyEo+2DdFe478Rfs6UfsStawqrbDIj8T49aFkmdH0Y
vvFHWWc8nBItEm0vUfRixzWIGdOdxG5mlQfskQMxMRxE/32e1EIfdQIJ1XiD0rOpEZHLUQ1r8FZG
z1Kx/xvhLX39ofAEM7fZCGYp1qAZH2b9n0IXbebI0ojnRIrZI/t0HlDReZf1Mvq4esbvEUvt0KfM
754bFkJ+ZXILsQ73T1PhcB6XQH39+zR8dopMtzi/JnS3XDDJIHRcKiUBJMB+iTku2fR32pkylvg5
wg1n7aDFSjUuVUOeWx6quW0vXWWxRHZvRPUaDXVEpB4s+0k2MBzeBFtGUrz+eGNLTp9/CZ226aKn
qOLgFgU0b5Q5UB1UCTFx4Jf3rmj9hqh6skibmPoo7LJJENJBJSJEmtHEj3Ump9i7IQwonpMm4Tab
Wl550lg9YWjAk+BJMQzRYmcil2SitcuVXLIQQc9vIMuBnjAOOKlxRBDkoQLD6LfSgMxEOicJ8HUK
9onk3w9wZqeloe1mKBaXeznpVts/kSitFRiE09A+wlnvXuZC1Fy+q5DQhdunNU5+6wEN5ELrySJT
3uP6J1ByioBob0o31vrzr21nfOrq9kHaBWNnCzSqZUIFUB2t60f60R4pRytRj5MdHFjLcrTrBbAQ
bHIlvaKHQ26bGet01ko+V2rzFQF10Zsn8AxHEKx2qWYlQlPTyXOWsOehhNTGs2tlighS6yytayUf
AlHSFlqh8yFqVUAS1nFqLOUCj8VTLMBx32I/NF6aRXqxeTF1DPLuWXe4FS85PDovpoccjM9RKhgR
kbUdvqc0B1R2lWk/Wg9n65faChr2SGj6C+KTgTBTDzgw4jHmeCiNalQnVZdI0TWvl90QixSU5MEz
NEFuVWQFqkiwdgV3hY5iLBQGWfwgQSB59s/uUmzcL8FPULhn1FtRHXirURcsGO5oCv9Lw1h/XoR0
KTdYcKMt8e+SM3jjye5eep4KjdCgUOL+65TBNHS48ngwvV6A1CD2XWybeLLwar1qukC4AqiypXM3
kFqfQeTBtTnHCQoPskO1KheAJxmZ5oI15qgKrSdoNVsKBKqlh+0gPFuONigll+eaK0vrV+yYqfZ9
arOHwAb3zZROVTB3Kttha5rZqWm8ajt6nQ9cFxxmtnD9xU4OtkX35GEtq4dMoWwjN4H/XJVBRrXm
HE3H5KLGVLINARtb6y6aSi5fNxDWlsgHOwowoHH7+RnQW+S9zZXtcKSDKWxZDhxQ6pIU3Y/c9MJ0
1xZhSXP+OuggSIGeELAwbK9Euy7WKX24d3zgHwYFiy7huiqsusGfpi2XKmptkeAYosdzZ62OyiYH
BYKumm0DnFhse9fFspZfue/uRgjjLT83rANo38OvDxh+ERMRcK47E16HKexF6pVyKsVVNmzpepp/
k/2VPVMGwq9U2ssgty6SJam5uPekunDfRM8U3v+J6otSLi5GdKjNrgk2hf74yS1UAPBfm37ISwOV
6YJH56EEvQWY8FBoWzmW5d04uMwdC0uX4QA8kjCfiD6JcykOn0yPJAOr45LQvg0dvCEnqMbrUGzP
paplZdz66X68sY8CCpm5luT06BwriSLr8UkcbWEMI+tyRUiWbOSJaXWTnJVB6A2RyB2UKi60JoYA
1gw9flmUBy+rCjSPFYadg0ZLC871LrrvGvvsD7WKPZmtAbZdMKLXm85DCy6tD1EWfqcPpjBuN7tH
Y15Ms1GqoKPU+BZQ2EzTQxAE/YoOxN6DR6rxwD+OgfaguJuQDQUaAxhgrGmNCJYP+Y+JRAEbiuLG
zT8NJkG3h3UWdT48EOing/4fQJfiGBz8Ufnr90Ob2SwUDxzYJIL4t8YZubh1U1WPX657FWUY0xuZ
JGfk58OxYci4C5cj4CQn6nQIZVzohpfKX9ph9JvUUuPvWUjWyVGaIC0fFLNNv5vsk0Uay+R1M1GG
MXsJBL2eTNsjMXhJtQ/f6QY6acPDICZamxX6FBk8lg23ilWZX6Cap56QptKgo2qUU7YkZ9TZt35u
4C3xAIuKAz1GBBDANNao1jEeoM6o7zsO4yPXlsIyS+QDxOvtLbqm9g3R9Xr4Q3ZCRKlRixqVTK2Y
ykdF+LTBIyjtsS5VpE0dxvBWGgAKAHhTxoI14XhjtqL3YXuTUrWfk6CnFBXN25heTJDa3JimqapF
f2uVIPq6T5kzpnK6kT48UuRMD6bB6WXD/o/6RfcjcqztwQA8DSjt33sH63xTD7vyWs93KTXkx83x
ZthAtEpG1/3C5tY2FigyB5pAgmou0WfLJUx3gXrJFTNxqhucvilyYvsYXydxHkrdOOXh4sTAxBrI
oyj7ThJN/qzhZhU7veCj5a26bOwxV1pw6f4u6jIkFGEzqbb9pPYSaym75DTFoC+A4+l/ztaBGiLz
RNKU+545JxikV7D/g7d1s4BzggC/DWl/ShNv1MOtxVE1s7uGkfbXlvCVnXs0Yk8dQr3cB6TJTfY6
m1vlODq0TDBScsNQtRyO8mOZ8jNv8LWn3VWYTds+2K8SEXqgBP8Et9jLNhVj3+/dIA2RbtDrgPp6
dwFfBNhczbnWnf5YivsUdjTcGtqqvreAI2RvpkM20Dyb6qxW0rWZg8cxCZzjORR2bBnOYekfJ1/M
qztFp/3nzmbrL11BhCBvEON/WBwnOkARUzgPN6QjO6SR9+PkZzzbCYAFzXnhDMzqY7bzzP/iGrlK
B62kn9WQ7AVbQd+7pePhfHgeKirwFDSWCR3faSMgGG1+nHFE80Yd7hAkPtTvZW9IsqbY2qE6knQV
uV0uDuGCHNRJAkQD6ZEEqFeDRmtprhikBCYiCH5ralSxBzZ0hPemAflKRyFiUGN5nPl3bSD/ZP6Y
sEovllLxZ/lKLJraGYBym0+Xq0noHbpUQISUMlZzuCpw+zzfG8AjF5oBA7wDa+6r/0sIVhtnx/li
ePC6Up/9B5qE5DLK0GD6XTBpMBnj9X02G1itoCG54K2GxS4EkzgsojuOsIDwv3QIkutgUoHZ1M/6
lVQ867dNsT8K4v8JyuJhmp4EV7Za9Y/RawJdQ52mz9p2L8mPqhuFbjbfI+j/+mkc5F+fCmzkyfb+
O9x+XGn4tddglCKMS1+W+S3KtetX5T7YabuyMC4eJkjW/H21Tj7pDtrjvbedeCut2BPqnQhgxVBo
ELpjnu6pE531M74rO7iCCE3tDJkxegdGtmlw27mCfLdtNFd5+Tm7gMwrNyWKpEHnwEBBSrUPdHEn
ESFndsH3rsERCFeAHSXM9lAF3sf68vYqG9ZDe6j898C3uO6t58S9jFsXfihjub+72Egptja49TXE
GqQvvpiV6Owr62nnwdY25JDyMxeqzQAcp+DmQu/M6sVAoZBHKhX8UZJt7rpfB9CCg/uEatb5YjoM
iBXZbisZe7Y9/uO6IkapxDIp6zD+e459a3Ne8NqtS39hSSE1S7fDg04wr5NyhxMmdXU+xsgaPzWB
HVMGxMDYIGjhrZ8Xvnr+FwjiolT62d/l1Zl03rOKrRSkMipX/IfTJ5ISoZIsboKS/OkYeVNQc51D
mPR/LuV+2qBSe5AZ7Wb+0VKgL72HBpePDdEDYo5BeSET5ruh6tvEP/5+3kUcV0FdzGdbi4nIxPjd
/AM7qXsfzxddvCf6k0KCGjnHxvyBHW30XIG+BL2dCPwFcs8VuHp42Lwzk4gc/3tb2wFKqS1oLZlK
i9XQHlDf897d2tsAc7/ULDjuvfSH/WX0570hrcXCIqMfcDUN5GNmemtAXDuhiCzEYnHVCeDzDhRN
5/ISfoKgmrEeh9Av5Mj7G6YF8bm9KExzbEeF9qPbMlNYwy8OiiUclzlqvrm8JQphkrOLcXQmEYF0
q581iSKtIjuFW48vb+P759k1enI4uwz1GPwF6bchu9BeMsOR0BJbkXON06Nn82E6O4STjorsxCxz
SLlduz18WsUECwqvymFofRlfp17syhD/v70FiI90eDxDU6ydBAOxMmoYva6q6DtuecFHx8Xmo0/o
XlUhJY1Il4o1y6DWei8Et4cuueH5dJwbZArJr6PTuYAB/BHENoU43d6RRC49L4hLcd0fQrHI8Mv9
yIM5mGEeJbEKQ5b89c3FAiWImyC8c8HmbLVZyRrJXV8C6sCEL/A0FEwM3IkE4xRhgbuJf9VAjEGs
hYRIPul5vqkLUKO6ksaLdujRA/RVFrIJiVhcDwbWiOQltIaLbHLV2vyxDukgZH6dqyiXYNykBOuu
WRvN2iGTVMk5KAjwL4319fqPGuoQr1Q8oIYQal4fKIoDg8/DgCeOqj372ChhStLPehP35Q9vFsmw
QlrGvbbdD2AebAKPJO9JbAAP8SqYtzDc2FZCpR0wh9EII0o74nBL59ELXJ+wD/aAiENYLjbiyeCR
3hWkbo0IOpv2xLuXToU+f6CKqAjM0ek0axLAXK3k+pFvsw7/KdKPAffNnRZEznGG9GAMd3QC9b8G
oZWg6Xx0+BZNeGgZzZ0JhwSlAJnEYonB2HM7+TDsEFtCupbrMduIqxakzBCqSNglRTVguC7IGb6K
k9iMPG7sSls5XsCM8LwwsytsDNswmeL3Eo/RP0XSeuzoDJ22qaQCu3lJ7Mz/bsm7/oC8iGvuhIUy
bcIYnEhlKj0lQFxnrzVuyrcV0KeCz6elSu76KvdjiEwabV7WX9oGjok6tTbUfjOJvDCkO2Kqc2vU
XxxyD4il97Yi6msDl3Ngv842rvcF6pJ1DXX21BavE1wJh+g8oOgV9eCEi42HQV4n359h3hhjGlIE
oG6qGjCA+9vYpNouLIagyD2AXFfjsdimPVN3vSH9cFK5gFJXIw80qmunisf744FmBK5elXzZZtl+
ngnQboMVhEZSE3VsuG2Ppeypeap+hrsgk69WCwEQX8ig+3jD+u+LrEmEzPIKa8NHXXLO2SiLUGS2
QSfefsJzKTSPswDqVKIYEFSiJU8HkNu6gjXlhJsneyTdYz10lUwqsakm8yTjvjQ7JGOkXqtaQIV3
47QAPOUz006XUwNaKAufWGaerfFmH6Xpy/lBrWv3BEI87vufj2RdUL/th7aeo9uki+D9Sb6m4WIM
4gUJ9R0aYy8txtVbF9OvTke8IZyrZ7i9+iHUxx6WpYSh2HFY3ScNS0s+Oae7zV4JtFETlA+F2Vee
vRKu9X6mjIxufdPZoWeXSKtfZSIK4bBXf/r5+Px08AzisKBQglg5BL3dP2N93DFCc6Tjmltp55vb
mrLjZjZMFIKqWFC1zG7kUprZA6JQddg5H9+MMMmegxwZlwmd4QpA8QNtfoq0mDegVD85dNp1yNYb
e7UdzqDcpkYaD7hIz1wh40NKKJU3q8pbTnoPE0mH10Nb+I1oT5ko+E9rXerb9cMz54GFFV9wNKN9
+BH54U81i1oyMiCbX+lLm2N6kJyvU+gmF75hx+9ac6qrN0YMACdq4a99YNkxehgED3oWvw2NIwF4
qUbB0VA3Oh0Z4/KqA8pWviwFIi1jmLB8vtUZCe+9UtDUkSaFgpDTN1lIBckC8M9cKIqBcC/K53cd
Bh8nB4T1pqWXPUunK7b1mkMA4E38hf0cDo8ci6LYYrREGKB3xFzHVAz+znN33L7fA9O57SD2k3Zv
tkHgRFNcawFtxJFwTsXeothBisNAsBW3p9OKh+VaQsqzIROEbmH7SOxlqs9PVQDCPs+EubGW4DSs
/HKgCNkVCJcqGCvU7C/nwFH8lS4Tmft60+Fmc/8zSPENwcuhmt9VtBEXmd6MijTBsn9IpLGl13pK
C+7x3padjX3gHa+bBXNsd/tMGmxXrO2kwpuwtGazlSdXIr7HMd4sjmCSorwSXooyBOMJZicA1tzI
cPb6FsqKPDRxxvQT/TB5k7uXcih86/ek7LoTXlade/SCDmhlsGbvZ+OCNwg5tIOExQ4xdFXbXcs6
n/yTxVd7Z+f431izBvs5NRLeV3UDMWVl1aAtxZ801K+zPLlVq8eHae/F/etA3fNXRQdWUVqsh+E6
HhpNh632qABH7fywg0B2IG0hd+OKXvkErNQcfj0Gk+56Yi8JHwIjjCJquICQXdLMa8yDwJZtjxIs
7XA4Z8XfJiadZJU9wWcVxN/23CtZU2ZqajscQ/t1X5/ERESfIkB7gwmenaqK9FXo7yLo94EFRwDw
V9RWY5lYTcIhS4qcIpOY/i5j7SJCXPC2P6vWiWx6aIT3vvHqpnqUB5VBoPommAD4Bkv7Vw/gZ/cn
PZkjQ8FqA2spNM1h7tamWrjhvd8lw3PLh9CuUiIdCoMa8lDGQC885H3j6RWLNivuO/dx1JCEIPtg
+5HJa9jgwnuDUToZ7v91AheEAbvsjdRkMRDi6lwETYty7DGB644V5aJ/WSmDkZs9CtJbre3v7pvx
Yw8JMW6eUzIivn224LaG4BZrs1Qj2XU8y5DyimHrVKhqVp0SsxkO57f4O3nXzCE0/YIOm0i/nq0C
KeACBE9oHnLkrFbOkfhXfe+Epef6OGSy5ZsUxnecmEK+oNkWwZFB2Uk7RwzPajLvIMzQuNLxCs5w
TEi6IToTwYPDWcy+sJKu9QrsLS6rCJBjMnvcjzjul3L9WuCLyrYzXrROOxIbe1O0RKGArJTKsKpT
TrKuC0ydojRzBKx83oroxi/JrnV3G47JmPYA792hfGCPAE6paiwrb3wLoKCo5ec4bWLgoTzfh9Wp
8kAT9CsG6LMT5wIZKv4xIppJ9XWG+JQ2G3xqWVzyES7/oqxA8aGscQv06Nn5MibNj4dfGPSYO46p
50dOxut2Pea3KBvEGEmQqx+x3uE7IfRrPfGWJu27AmIm3ukr1uDnq5TXLhnlR2vQ7oVcHffm+5yy
to5OVqfb2EhamJHHhCWqJ/2PAiFM5EHVgKCurnjXafSY8Rux/4fZoo0C6+ISiDG3wV0Vd4yh1TYL
OD8D0syOKuoH9i7mS5TXxU3tFZ58ZesN5alIB5rUn4df7AageyhTML1+8GyFHmvIpFbUzUDJZBUL
BNg1SskRVWO+7+yhomSCcJh9fAqH3oGJmmI3UA+yriid6N5ZfVhwfMe4TI8VV4evibGv0Tu+MAMk
oDPPxLhjPot28w6932LideOInyu8YsyjlFXXf8RPXcisHnRoSEaNJ3ttv6Xg9yj5uborKo4cbDcs
wX0sONAfCN1YDLvH+Xvxcij7ztfFIGF+9fJiR1KW9XNAanULz7uelloHrxn9iGaialdkl3TJKzrw
DWwoV86hNFq8lFYvNCfCg8IWpqPUuBHGZ2JuTbC6kajLokpCdWxRWM8HikLO8w8OYZIcH/vIsCzB
8gDvjoc6tbXShnYlybz4/7HIc3MfycwE4TIgF5vS9TSORNncObMa2VjD29JKYt7i1BnN1qfVTtaC
ZOA8oT94ovmVF51MBZfnH9UcolacTJV9UEz+Lmaf/MHRM6ZcYJZdKh+0eiVSSoMY9Gy6uSih9RaC
WTwFb80AuMk+tMXhHJO4jDlq4j8JmhJkL+wGAQqSijUzRkKa8u0nhlatF3S5OhRFVr0mF8Gn3c4g
3GrEqtDTWrtzMWJYo19vorKhZjw3o0K/6HK6rJNdrNT3MKT1kNhFm4QcQuGqXUck1IPSnbcyhJHG
KvqOWAKmGdzdEeZtkI5tdug8uZVyURghE1kpP2zp+RHoJUgjx1ueQJjgr9zoz7X94uYH2phf9uXs
ObF3g02kJ6t5N/eT6I8KwunngSN1Yoh64AwQ/HC64DyTBnr8B68a24uJ25zNxq4S4hEbQcwgm7i2
rsRKlzY+NGn9r+gOGP0ZHW/CvRca9eT3MT4P65Pa43mqaU6uNHrcVbr+YmPJg9CCh7KAyRW8QFpe
AQistK9iUANtKbZKvrve1A9nR9YBRP2oxO7A377y9xmVUVf0JOwb47xzm2cVy87k4jlUk573/7h6
OYrse3b06icyT21kQ4XbZCGb18HGm4icdfPmo/74R2IuVV+fqI0c0rtB1/bPonKZ8l6IMff8Z40C
std++COGBCVcCdTK5/Wr+3DaDXcV5QqRVBlM0sQVNLJRVxS1tKYxck592HO1aCuEVVSBrqSZSEx7
7hesGZbeeTBZUTaidU9abhGeqJjMWfCQ3wabTQsuUDlE3Ee8Pcu8817M24vtvhP1/IQJUulJYt0V
fqwf9kuSC91w4Ui7huXP35Yd4kv1CWlWrPN7eBy/yVxhe8niufHMc/ynCj/C6KkbMrpU+ySS/aKa
icCVoLzxvCvi7gtTfmbI9ha0GBgf4S13Xc4drDTYX3KCIl+GZnHmaD2ZbWHEFRHv9LJy2YuggJJn
RZMtBVPPi3sBWMsiKWpftPxDY51kJ1kLLzwSjnGVkcEkV7DieIcAYK0pmmrImrrsaHvSLbzZM/L8
hvwbtT4I8O8AtRAAPB9T8Hvu9L1/i5El23k0uF9W+bo1ZpK/AM8G9SvPY1maxlVnQzxP2M/ggIq2
kUpDM/AzQL5JyOt5FVm5bIe+WndIEoJkBBDqWF6DS1Pe+/jN0cMqUIV4+HUpYJ4jJHfOKIByo5yP
z8XeglR4BMf02v2sRZFsj5M0jcF9sNRzcFXfmt+nI6KxKi+Ko7p9FxaVU5Gyk3KvMvTDIIFBd0Sk
Z2Pku8wVPp8w0NUcG3ap/FiWKn6tcJYj8+Oj7w6mAqdr6w9VSCzQliNrR+P4G+y5ydI819nz8Gud
4y1yAERYP0IRkkuoaaMMSwj0kLN1D8QsLcIvUKMUl6md6lEznmQjKGsIzkvfKKJPjYZc6hwAEw+v
+PLnbwI/DK2jVkrLHhUj0zwnC6GMY5i9qsUxmABqXYbiRf+gU/uxJNT/2ueoYXFxb8J0kx3F2K8V
/BGzwVQOK6BH89BMRCWiHqXuqV0i3HFzkiFwQlBC+BHLWrsyzVy30aDNqBdusizr1Gkr2v5MlimM
4MRrlMuxvKQcLcoevR3fW+I6bZcqj2g73jSqqOWefDOk2sSv1m5AQnj52VRfmru5bvkoHDV2J2LV
tyJskd2F1dItOAMT+LOVloLhnS18M6ZwrqgibeU3FPG9K2E+mxsxweKMpX+CUub2yADEiv6JH+eS
nO18B3IgeTxoYQa/fM3UqIClvCqEE8Rgs5k8LUqAulVZlpIMLPNnNvsRlHgxyJXk+Fv39lpEUGpB
6xlmwRPJxiC7wg25bYLnNAx5fRwWzWknOBgb8smgByT9jLlNG2BtZZwck/e63o1/7WPQ/9OOnk+K
ot3aJ1bGn/5sFjMHKny7mGlUUzMP2dpeMmQiXBwo8I+tGs9E6gXpR9DA69p1XPkK3nB368UXcbcv
sBKg5Sa5jl3Xcnks/uF1nEo5oUbQxzuaqNco63PLg3osepLpiaV4GsXr1rWrbs+awUqPFbTilhwv
HF0p3/EirHW89FEgtdAs4rqvtbWEGeinXGrz3M4OvxSxbvBVzQR6IuDaqzy7yl/MSOCSPohTXxcM
lYAKiw4kyf14TbcftUJkQbof4WAcugshw12usNcg3vGMmQX+aG0dw5WgxiKijcBGFPkrPWFCvQwa
/H4BioGbSsSYqfMUmhFE0VOHIIrIbsiT7hfp/COWI5WkXxlAvfIOD0+laH1nd8MovL7qku9ozUPS
yFZGBfbxYv8BSIbJvs6uO61nt9inzfwAO7r5EsWU4/jSifhgIzEl6r+IE9ErvdDA111px1czRh+l
G7JIdAKWIYdmlxbw+Z6/hKN2te4V4paYFIVIERSb2ZxTKCXs/FBmGQXpmOxNDHJAxtGXz7WH2LsB
YOnwxeZzkj8gba6xsDIwLo+IILwRG7IMrBVNlFsVd1gaEp+RzM/1yC12bEISJ909qnHR0Lgl38zL
4J2inBzQufCoqTnEWxBpMac09v1ijUY22BDsIuATb68heE2LkaTerQxFfshNOMRJgxNRhS0QfO1+
O3foTV8tiTXjg38mPzga7m4H7YSBl7uNoglWjfSS8C18FpBQwlKNq1Bayg/akgECDSe+Z970nX9B
w4sGPTwtdD6bKR4U2PtyoWwnYKl7jQl4MLuhZRvo1zd6unQAkhbLq0IwaJrCoe8baR5ySPd+80g5
vQv/Fu2pNf7W+4d3H+c5DIFjlPjUiCSv7izhb93yb7NgWMbJ3ZA94V2AcMlr7APdkA3GSJ61rP/j
QHdK0DiqYe27r2BbsW5CT9mzXiDW0IUpynu/63oV+vE7QKfkYOGu4iAJ2jntd7+kVIEiwehPx081
M9BrI4n+4N0bJ6sbr4DXcXk7/5b0tMGirafYKLkuPU/scYBK/Es7wUNwSGFqh7dSS8Ldsb4GmIVc
5gHhtDWWx+nyLYevMVqudkx0H/QOfNn0AfN/eggwc88gJhh/3EYEPeOIyUno6RDoOgpOHvj5v6Om
CCO5mpzJLC26IYSA1lCNL6c9G+K6dxHaW+wYLilbfxlyxJKJ+G8uOuAB6/rsFkbtJGOj751/Ti7Q
3Qtu0Yc0jA19XAcsqcBhvh8G9GagDKGnB15xd4NeYNw4lrXESGItOzbyG/GFav3EB2EHZnWy0f2T
46ztll6Jk6J858keU3UHlZPCIB4jxvxzsZkxmNToHKN2BJxU/DIHJZtWh64A5grbvZs0w31iK1Ap
uizzGZ5q4o6kFpn96oPViTeyFTFzk+qb+4npO4u/dZ5h21vpabUQxEG7fXQ9Zxi7364Xawdwfe69
JqIKD3eiva0Luy8DhvStAqUAQpxD4sqYrXWfKezgDlijOqrB98HyraMyKexhSG5w9AJvKpKffyQq
cf+jWDiYDtFnNqa5Os0lmFvIhtuxP3HZZU4twOvi7MV7Jb1jYVHInEfE/m/8xI3SX5+TAhYcp5vV
RBZoOsTNBZqSmDOR3AYsjudi822ARX2OxXP5lT0RNxxY4sCc+eeppOrtpl++LzWT4U0Cm8tgXhGQ
YBGwn8L64PR9YKzrUaZasjmiDDwBRQOiDWji9JxNTIxLEP9XUxCfxRF/EWkY0efk6mUuyHg2qpFR
yz1iHuWcXZpJFrc4IoY6uopX33lOdf+4UQh7K7bg10IYLzk8v3PTag3byQ4GrLLdqjVKghvyvIBY
kvoXx7I/gtMNrxOsNyYDuCJtNNSHdD0VcHt81+BH5CKq5Rk3udjydXhsDpwcK1fs/TvnvvIZbjcv
njpJnilDsQqaIci6W0jIE+OtNGMwbpczajwXIXiIfoEtzDy6VqfvfhCGWXf4YYQmvxZDmw7qXBqU
UfC4i5+Pun2SdDHbWVg9m/4dn71eQZysNR6DBM68Vlf0r5/L9PHl+ByCdjDkwqLyO/pMna/P2F1x
2XYLlUxcRaIU/alg1hc7FJhgmczYAqmbZCWZNWsmxPSntNkFVE+LU8m2c3TcNuwRyuEZ95/dytkl
eMu7rYzrca0/RdzD0oATmylFhsSXI+B1T9cnuXnEfMcfXNW1scZLPha93BxxILxcJg8HrUK/7YHt
lKBXklesXohF9k7DnGDuanHGdNF1jaMM209ytEA85Xo9JHGyWQbn8WTs6DltbyZDnlHRQA2Uc3dJ
4RcmImGug2w05uRrBCmtieT+Ujv++oZEAiuUnjtluS9oax+ObAFoYr389L0H13e1XLWdbdKX8zJh
2x/WLblOiXyZJtqDlEILiUjjXjQ5BmQssLkWp0J3V8CvS4omj5PmE4IHHnqq5UjT+6DO2gxGdo8h
fH+eR86AFfRKLT2q7wKZBMoF53oKOD22uRhQXQr7UI9OeWpN2DlID1G4R3KEFZv3s9eySHrkLEMd
CsETvSj06J8K/0/Ynz9Zp5rewON6rRUGMc8u+fk0DiY5aKytD0TlXrML1Dv70Y/oTq6XLT/i8IqM
sPt2bgv3A4eu1gxDfyKXcxpxljOvoxy/Fb8uVmZDyFtnOE7Fh8LlVGwLmNFwDjgXYvNQzNvpLNu4
yT3ZV4K6oeB7dxSmrS65K2tKSFC8wrxP88pK8sS86H7AJK0zk1opA3HwBiKaCKogllV1j7q+4PMs
AG/Hsv2X5mmztPQa8P/yXbpAC3jgg4+X9NfJuHQ9c3aQtMMG8qWI4gxI4pWdV0/41QNaRK6WJF2p
2oW0rOML8AlFC/JNOFyVkvDUAEEo1CtvE+W3EXPUbm4FB9QtjRTbLQPDxWk5qZZ/N9R9c2/AJ/hu
oNuwSARP8NnuLSRe17KS6vAc+wIWYIJWLPFokehHxUHANJXuQs95iix2BzBGga33+wqBPMEmCTTv
DJvaLWNUadc1LCqwD0ZGPaHRvi+mlvt55sEJefJ2srPqUdBuXdK4EI3StoL+GyUwqW7RmwcI7J20
yVTTzgNni2OMbkzUC4iO/w4Bxi0869Ts9W+hqx38AtNqMbhT67YLNXWRO5ekNF6BAncdeAPYumbP
YHo/S38V9TbbmezIB4wweKAPpSYUiF2gCwPy98GZ9VZ8Beumiw0PvFpwE0F0M6NP/8mkIdP1CmPu
BnzAYVDjhWncqpYC6Gexp8nVDWAhLvDCivkEA9yz979KwFvG/WWoOkWTd/SiaaFjfD/7XA+0o+RP
QsmjtVASMGwy2sKml69snLlir8WtUEsKW7zQdUYXBZTcFemNUSURhyS8Mrfp7S9VPphzcu2rRbSN
sGX57KJlvQnShI9IUs6wknDZ4X2GKPyPYg2I5f5jo2uTMr/LQhkK2AgTX9kwXDL7nKa/+IE6bZUb
7vkmtLbbLUHnjItAk9FNxOvEzDQNmsUctFBsO5Fm2kNiA1Zj9j3LYXkU2EX6LmEZxKfGuYKWYmGc
zm2f97/VLCmEd8YyTaIVgVWv8WD82lZ57Su83JYIZxokgn+1dWc4ajBHNiD/I5G/OHWMv/qp1q2f
ErHqfELHdHZJxiOLafjuhnqXELErNtS44YEuxbrjER620/lp26KnQMBPqW2oIdaautBhc+gnfncI
jE9gJJ4P1rL7V6b1Kpim4/5J+foYRqmSbGqhBQHDAumnR+ls+xoKp1OWbtZyNrpXf/Cx/654jQFd
9Qs2tp/1TaHv4WB0sZ/LGERys1wkM0O2IxwmUQ4AtbRsAU9PfsP3yIyLnMYbmwF7cMyAjewIJ3Ep
mTi8fQMdhohPDDnHeiitldHRJqWe+a1CaEZfaxDnKroAO7WKBHBc9WlpHltv3X/YNQfLr9DJvRJF
a0N7HfYRTg/n4cphVb/92FqTWxMjjTxJYupR8EzH6/aGizlxt08MBOsLkYFKUi3vb0pPwAThuO97
vBHIBkdCJHN56BAruGskkZ093Tq3rEl8dusJuGoB138E3BgLIeBK9jSdg3mHvHWsJQZBFXFGgZFh
/lZwmO2oedvjetUH4o+dnJpSUY0YV8UA5eZBilyaq0xPtg/Dui92Yv9PzD7VPBsh849/j3r563xB
fl19giK0bf2KwOphujYj4gN08saaaMqIj3jgz1GXpQDZIEGwlve0gnt+gbSwezHmNNKVb4wIj82q
ivBfkDzI/7clxV68/QUdbAoEFZveOIFJWiPhdi8Y9jXtRwaA4vMoAuCAIMs5bvnCO45RzlDTbajH
acif/COynxftevPlIylnu0LcJwis5Fy7uiP3sIztEUcqiiC52rphsZQQpWUCLY3YRe6XHEyoyGZ9
KIfakwKlvMPlPq4r6/UNNuTf0+dMlB3G9K3cYCjvsXjLPYT5eF5iYZBtSfUAsibqaE8dtEREAmLn
RVM0rJ/EGZ0Em2k6O7wVyJBOsfk6xZYeW4b0Is3OTB1iShkvRQ+NpmmGYrl/pyAT9kBREhYp3Ve0
nx2duARu8ImtNtnWtk1gI5dPLBUHKPxYzxeBE/Ep7jCweRmKxPdYzTH7sJnAjSCd0oJ3aTRtIjuu
bMEUxq6b8TUiC92pS2FFL0a1l65HgoYvxGxaBMKiWHvrVLlYZUdUB6PW44YRXeJ+8UOfUESjfpdg
NHpyxLeILt0t9yjmhn9Ji7RTihtc+Lwv1uY+/V/wdItE8SuQvOFLQia+J6B+g0H2SeqEA7lNLQqH
FgtSvPNtY/iN2KkAOkrBXEuLSqCn476J4+pUuqdhkEo+MD+jHWaA1X/wmk6jZpXefE3jHeGSgwB1
KGPtZnOLhKKKZmmCPiTuLDWDwOix1WyEKnSqGkRqs7dyyxaJLmgu8V7kBwH2LA0h1MMpOulIMRLo
Zj9q0WMeO38SCUsRB06PXQK7RHODf+3955iBE/AndnL4nGtHwcT+sLZEhyzQJylFUXsp6eM3r6SB
suG82vb0LtKdAzJTky3TcnsMFmsSUlfVIQGe5QIEfwLENp9qfio2RsFw+3IPp+mQ9xKmp0WrqSK0
ks0k1ZSQ2kOuNANaKGe6THGWb5WKQKgx2FF+cNTmcpRlkFeobiSbyoNnBxc40eDzGGmrsC3iLJAU
NOTb52vuePbDkCRiJKotXKgWHWHffGPDfyX7BhVbxKpiB1C6/41k6e0HYjb9Nzg4DYkDnaQwqOSk
DtOW3Rf/e0HIX3ntNAb6bub9X4BacwZBOFfpKRodRLmCU9HUWAUWASB+98/aKYjrhuB/JHQmJMOZ
HO7efskSjMamZxoLYMqjrmIg6B4L69Hok/+T/j2Wz8E5bxHdJQilXLYujfKwJJqpdZr2hFxrzEEC
DiaYYW/fkn/dqHOxlGRtaC3erD+lE8e8ZHx/5/GbUyoLYzH0wByQHA+MPZ87/I5gagzWa89W06/o
E62NmexZ4+2Mki0QiTAXl86/TAlGW86Ahroki0koHj9TvOF9uTyXLO+mXq9/OHHE/yvv1O5J3Lw3
1Ik+ZMlDHItYrRfIaapaZQU+8ZeiPz0nyu1Xy6/tqAnqpt5aHfBLoDQSrtMG3oKrmPGjWI0xjzDt
50Euuliupgjt/rIdK+LBWGnyzmg75XzuJR3IwgO4CKxYcZcBgCulUbXsHS+cCcORaKaS60fVXZks
+QK3EgiSggWjAHls8XvfSjyY3D3DqOeT3QsfoEZ/MGl5eCJCmFPzwkGPxZqRc+/mSy+nriPqtOBb
OPBhVfWAgD8ShLbviY/c1zeU0WALczFk90TU0p8epM7KHk2zu41QKUxB3sG05nU6YJOEuYuDx9Or
+Xhc54S4bgw+GhOMnOwf2zSD2QGm0MRstaPOfzMizU7MsGD0Sw9fcW9WGFYogLt/gfqK1I7PFsom
H5rs/xVZEo/zi51V9G49IKMCk9gowDV7iP9lFpk4U6BL7FY4arsfncaAZ60TAdfOFxxOWtEZIq6z
urzUUHxJAfsO0r0VdXd5+S6OKDNmFD1f9ZEXcHv22p89AHpd4orQYZPeBtI3incD08cKTn6pb3zM
eX9XERBu2g055bzG8hhm5VDf+n99E19dN6k1hQ+lJlcf3c3pBB20JTC3LDtiFh9gOwexxaXk01Bx
xxoTXTYeHy+BQrTVAgO1MmgR/j+OjemQtm4Nm6nDFoL3wY2MEgEUjqHuTyaZTGIfYynm0WFJIEG3
Nys6Gx+i5jg9a3kpu/ds6sG5Xrxp7cy1sPCqnTIX8MvKfuFsiZaNPCqHlnCMauVFsi/Yao0DGiDX
+bGScBScgkczxMaOyFk7/U5vZa3lstGbOwBlDwbDqFRvcXye/MKH1cyw/8D+k7557NpGuj/YH3sI
L0oKwoLDkLdmlX0kjcbYMRuVawX5b3UdyZCIxR5cFB5Nu2Jb+NbTiOrOtI/ObbNdhLYc45gx89Lz
Um3v7xYvgb2bYdAjitiASfLhmPJWeBtNlYpGq5MulGATz3Uz+BXjn6efzjP1kQa8IUvuKNzcHl48
KJHMANcsKD0JML/E7G768CfpYuv7Kr5SrktwkFb329N4KBdt6UiDS/DaIYC1EXiNYfkcyNemxya0
sJtUJ/wL0AgMrl/u73lGN4CJ4oK67lhwojF0spwNIEeQWwKfimmztII6qgcA82w52Ph2Epeeljro
SVkiwJhbsPibSfx1NyuGKotvmfpeAGT4hSeH7JbUsjjNaQTUX4Nx/gTeozqIqHHr43u2Rne34O4j
smNi836Sdc0qVvqtpXtRQisc1W4VF57PHO/HlOERKWIAcUd1mhkEATfY26rE/35ye7jVRN1jTxw1
e1UcyV4qmruqzINUV77ib856bCD3xZVf/38E+ipqmFvHQ8+g/84W9g7qqZ7ErG5byEmAafIecIRT
xMR/2eho5NT+eUxXh8Fy4S1AXUE4JEW7L/Mcs5iWSSdOMHcYTqzP/lZ1cpRf2zylhy2jgEDQqgO+
UtTG2RgNjN+4BLFqJTuIPhVdtxdolSNfCoTUF4wPJt3ysdSdt8QTBZUXF5snfUIomB0xU3Q7dnd4
7RtKiaawGNTjcYNQctsJv2pvokHYE2tlkEMJHpsK+vVPeJyTlbsJehlWhwJd3twuzbGLoLHvJHP8
GQWiP0a3Inhi1Nv8LuFKD8CJe8SjVOzqLlQ+knzN4skC5qklnyCLkBbnpEjVUeJ7bJv9YIZn5H8R
LI1px6WVd9Asy2v8Y3RYjNGCS2lFH5zjtuWq18Ckx5fVPkJ7LDs7HVN43fZB9+NFgZLtAhLJznxC
HBYHgs6Exol25jXFvM7WpPv3RQLqjtB6pu5Atsxcf0sm6Haxx+w8zxTAiOSVm3um4HMfOCQG/cjo
gHODO1yWl84sE1k5B/Zl6zTtp2kRCzEcmDtvykBTnqWE+8OTjjKBCEJm3Dmf0uNxwUmSKBMhz037
U6P1L8aESTRfvSX/Vj+z7IovIZ4DNTs9JoM0iKNHcUI1v/7/zHu0UJ78DwuVuz34GlzKR6/A0ub6
7U07XJ6p5qrYJiBOmdWOET3qGIHvwjt3gtc3s26FGJIWrk56in4AGedASJ381BF3YABDFdR4XGiE
dOuZ50QRwQoMSH8qnb5OFPYn2eIQoaeAIlNbxxyyP6XeCn1z6AkW6dOiNeiZCqpEOwPZue/866Bm
gwvPMYFIuaQHDqlD3zCKaq9voKvOUW5cgpZ/1EwMM+RFY7SmuCP07MnNChfIbmumdsnZHH8N6Foi
Ph5OKj8RgOguuuYCffJ3gE/pElNkxOXV+4cosJMo2XMW4umwB4zueyL2EqCwL41awjAA1avGQYRO
mCgFLqyraX51scNGQjCvu7YQffVnvqN51ilFrdBlBrXrwZC4T3umamGT0+PwKnXmmDC7r4fST5td
timen+ZfIrSyz4olWHwIbIJ481ckFHNtgz1O/vabXeMP/fzpTMKmTxn7RdoNz5col0zhhyFW8E8E
mYde4FPCSc/1KoiMAJffuJuWyhyPCAFyNC8u6Tafw6otT9tOIb6L0KP0DzbzDtnfQwG72tWBuXsf
MPmQXws8+3Y/rKSiTVxORaDqWDA5pPlRUo6uOhObh+decaHswH6MC0haLcIfDhzOuI1LB2G3VhNO
MKWN7D5BkyRihQrnWDvTq3RYS+aHo1N4E9nrnAt+Zutn7pvxnRZjSlDvnWYJxWkxvYWFuRKXPPo4
X5Xxpnqr7F6Lp0/iy+8gH4VkAX1srlUrs+hIXbpQx5UoFnFQhmTxf1QsBgVzbhcL6OFlVbdO5hhr
8DyoNAmzDpf2WaswIkcMFhTtKKmO5OR2NiSd5767n20PUbw18XSLIwiiSxO3S0Au6z+RBL+8KNXq
/+FS3cNMtjedKllHU3D7rvq6Zok0//UAKJaEAVcCjJipAMyBd8mNC1CKZYcl2GK6ZTzA7RS1bVQ1
KXqVogALQTsNG8kQUu/eMxIw5yfcYQmXh6Xcf/Di71/B8RxZJvQfsXTt7DuZWQ3hOO5ipbBKHMaZ
ehdbRh1gkZQ8R3efc4L1f3Pif7eBR8dj2HEJoitkFB/V1rqCW+wZKNMdQNTe7tmcWcpOl/Cuk8uR
CJ8fVJjQTS0wh0yM3b9ZyacWIPV1TPMqdq2HZyhW8Ooa9wbqbJ6twEFEeQSgX+lBe43BsJPqsylk
a/bperKaJvZOHklzNFPGFPLrf98evWdTxrod7pb6vq6L2lP2Yr+Jw31gvw/rdk34rCb1qyCcUYKi
hqnCfGB50hIaoQJ5qibgwuaZYAV9SCGiHMdN84595PC8a7Ic3WuZVNZE7YKZOX5p/fzVDOnpkD2J
+JZjVcIr4TAwHuPrpzpJmQ0/Vse+DmNCSWvaGiyNZxcSDqMzZ03BKBGfRJID/8hMHUQlsKrLrjy1
DeQEXDOdOq5dO3PuD5jTeRGDy4AOlbYbTDg2ph/dQdzM4nOl8pWnYsc1bprwceEZHnt058z7tCY6
C8vt9zT67RFhyIXylmj6RzLVL9vaFjWdoSE/SC6FKASYSReJrEk24neICBe7CzhoCkJgVDuojyRp
cCm0nfc8yj6TNAwxpGC5KpKQ8T8zS5TZVZWUFgKW05/UDuvbyXSotK/izYj+NmYT79GkohblFti9
XEkYylb8Oymf2loLdjInBzDKtKZUPxfASvL3yVTx4/dn6BBvQ8w7NGoPTGZCObUJdaBYdTbeygQl
vpkT3MmliKJod0I6bZ0nVp0f8vm3gk2XJL0G4QbPkiki+xPBT2Uv4m7DdRZgWQLipiluP79qPPQA
ho/7Ss2AYIBvmDOlhlP+KFzWRusujorSFUxk7QdbDJ9PmrvQRkkyK9zwCEWyQtnfIpIzMR1clpub
dkAXfCVPM4EyOc3WyCU9SxvWOAVrhuUAurAoLIVrdca1bkJMF8tPTvAaFai/vTfqeYRa+IaTlCpK
sbi7412uhbUgX7jxfm8bsELmRbM9O1H9Ttebz0dTHEIr8mKY4x6r13sl37p+Q/r/Hvj7Qj2ZUGqr
l8dPvruCfnjdvSU3NyMOkSbuE5aAECwXHgXTD6/U/TAewIMi9QLtGJntTg4t9XaFRNnSr3bOV79f
7SsomK0W+ztuXYk0Ty+zBtlxkUoaW9D/cPw6XJcUBVfknFBIbw0DmEmG2DtKyiyRlV9CDqXmprOQ
BJmoSr/wf+nH2UpFf2lcTOEh0J7sj+CORrjmIwSn9f2UTYtpKyq8RVt0r1dv3xR7DWQaoGrcBQ+K
Bi5FTZ0zOdXUaVi1xZyx8NQnA0M5rVtICd6Sc6EqnkWZu4/Nv5DaFXE55pfJ1PGoqb10IjZZUYjf
/1WdaFYE7IUjRmKT1+Ab1HIv5/b7352Ozs0ErAxvjWBwOlvUkgyjtBhVPnRFRLcX4UjFKyJ2JmMT
TJ29NrepuPuPSysznsXEnNQj7YvzBw8bDsvwL7IWQMXM62Oy5N2XVzxl03RCHHMQgLKP2ERX3MBQ
FIg5wP2RxLDV2CIgvpDFElFqQ1eNQeKV/lTl/mpX6ezAJpLLaXOFVBSdScMBOvkEF5W/zltJQCw0
UvFwjCvxzj0yNtpP/tPgLdUks76CHBWWiKPVv1txX3AZeq/Ipx0zOhqjeRwBtwP2HPOFCFMFDTxi
FxIRlACnCLzU6NmpxG/hlaDi8od1bN4uPEcoAV4z6erRYsW26Y1PT8NK0jEYNOZhHxOVEvbMvDvH
No5PItL0ExtDCQAQ5xPN+M77caSaMO0LKEJ99JbpDX9EhedQDvvvPdWY+7yxb8RcN7yaT4pCi3dt
QAOQ4mb3tsEl8eV9CadjY8bU9xDw+cVRsJT1baIrAwPCP6cikAuuH5+/PF0rHBL+dbJ4SG61ty+P
fFHcBXDI0x8q19Tcmts9TAVCBlWq5XCjWwxAh0IcyehDcKhp4/sj+fe5ogjNdGOvjyddiq0rjIAQ
QBt8dnMZID/AyDZ+CqqkVa/fbeU4EaaHw1pka8pekxVmUiViDRzhFqXG072z36xRCj0yBm5GfNms
K/pUAhDh699ECQG2uryFvHd7olqvgQ7ysOx3jEiOYbRAQSnoeL+HcsO34Fpw9rYv2yx1FKU3hTpm
p84zK0FvvLO/ZZkFBEiPbh+icv87BZuvmLEVf4beqxhoLLAWjTxRu4LFBXQpj0527A1HLDw01hfz
RHBszg+o8PT+KqHrnoqF8iS0OHLVBnbTZwRJkEBWNRqjd/JjcbxYsmUJnPud9TNo3xTZ7upMDLHa
f/HYsHuV56L+ElpEgBF9H1vcUzddEbGAlZZWJApP1Z0qi15VUbEjDFuU0Q/yQ09QgRt/4gY4tc+/
GpD+7I4vO2+DhR+0u3V7UK2AigCqJke4XefVuvsHdNMl4/LpoJv6VfOhuv7FDyHOib6g7ziTEWX4
P9KjIvR1X1jMT+YBNwnb10tN93VpG2b7j9gE7/985BLgmONWV11aOTLz5p7IKwMjy9cSVeEZOPJj
3y1GnumcocgDjW5qwoylS+ON5RhQ81063I2m8DXrWpCaIDGo+UQY6x/RUs2V547mv0f8HFZ09sFU
kDCxEbSTkObgxgxQJx4LTCrzwzkBp+XVnH7jA8qaPo9eXTCTPE0VqCdP4NcAilkBu8M/yq/rALbs
ezXjI/hGIsrUB0InnZdJTpHJLpyEfEcZIYEhkORaMnLcTPzWqJ0pER2fLlHIVbS6ZftmZq8KYOq3
2qI7061sjHkkz2IgHkaH5FQyHzpWvQvYs8wUTz63BVJerYpymaPZ6/fzq407P5GO+7eYtXB1Q/zv
7EqSWd9uH9sQL6On46AYxKGnTwouBhhJfDiTLvuRPTR1PoBIi0cTnEZDjGcQSHw0oHtzlcS975v1
Vv8arOEwv7gBbM9hrEhehBbOhFJU2N7kIkU3SGPwdLiOs+R/wWdOMcLS4Y/gH38uSUT8URX4u/00
`protect end_protected
