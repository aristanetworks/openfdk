--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
m6Le67aH8JXBws8oCUYDkIjom6Mh8rbo5Ko46bzz33L7jVnAp0isRCU4Fx+sgRoeLHefxrufCrvs
A8+CUK70ZWUrgRUnq112J46PvM7Tsaf5TPvPXciFMfUOoZs+Kjt+WTnD+w418KPCLQZ1+Khh8Bpa
qHWuH6AiW0yPE2SSnhzX/mCVr/ocUmqg5JDEx7iIYW0CdF3CBatu5igZKv0xQ3UeHkRmN+ZxV2B9
nHCNZkBhzFCEWIMg/QcdurfpnB4uNUrKwSQX8xNIpWXU/dOyhVbC3mY4gSJLVoBgZlfNxLF1Wc52
cJdXpI90b0iYI0ASz1VYELSKOO1Pm0YJpvy6WA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="ttimRHztqiHC6hznypMfRpO04phjK+nJqMokwoxjj/k="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
DprYib1QsBUNXQw84qQb8edmL6f+4fyQO6XeFEV1DzZnQKEru9xAvNf9mPsM0ghM5XTDjjwUfkt1
bI2CkoZErGIvWbQ1fNGNYLKT7L3Aajz2bbFQ4nUhkQJ2/j8EyL2EO42S3fN1AvDE/opF/chVtpL8
AyWI5mQLnCp1BY1Mi7/wSdp5XkGzJFOK0F/Jdq/H0ekvz4k3EKJeETiLcUTFuf1mMXqj+VBzIb+9
VhTxtgC/xhqtDK6sft6bHN/20CFn6KmvsLWRgIqx0HoHQOOth1Mcl9Fgaoryy5NLYY2wrSprN8nz
8ckKpyKQbPF1BIRagxrtj9sAeKOZhaK4VnbflQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="chS182LXK0/GGegQWB9VgNd4Q9pV/dbTZKusDU9e85I="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2512)
`protect data_block
ZCZchjrE0cpG29IuV4BKiFapoZ4mAyAclj2yUH3sZJXdxkPesE8A7v5vzSxCsaZx80zYDTLSF0/g
fRgEKZ/vpd2uG6K4/FXUu2HuoCdck+pnZjxUf6n1FhXzmNmu9t09Kx39+l/w/yxDokrLzr2nX0tQ
cN6htQgvBh2tkfA7I451LxMzNhS0KPsOAEM7WlGS9Hl2hk+Gukw3lDt1sDoZCOC1lGV2vZNBsgvw
o/jbnpBeE6Jem5RhGjhmavJuFlwQpcKdEttVwCP0AUOjW3b6OzBik3kWuaNNli3EVPzmdZJSE6yr
9JW+796hgvR51cEXuk3bWyceWpFENUIsMreOSJNfOeq1jG4pecEjQO22bMGSPkdplDcCQ5cw+ElF
GdIjX2LLF4UuAlnFDoaaY54m761tuKFZ4f0X2aUIV7vY0o2hd8fPtEOa3/xcowRj9w0dDE28VD5d
+T/DtO+mFDwmXL4CRfOzxxKm+M34n48ljYjswu608dD0Ran/0zyAeYs2G+z0PRisim5Ad3P/cFBj
PYKIHOtbLpQ6CyYqPAWbkfGOnxbHDEF5JIEiPi8lldxMAeFs/dCd7wSTeH+Twj1T7xJ9Vpg7vUU9
FYjZsDaiEo1OsTp85dOEhG6Qfv+fKdz8Kaw+CSmnbtxbh4t2gzKFQz7FHzRewA1A6+XJCBtQd8fU
MKVieGOyfhCWht8S8ezmFG8ay8zZWzeQlRABWDizvkc49FiB4T5YuTVgrPpxKwsMTXVf0y/5AAcd
qGoTUiHy0EZRY3kx27ZdGJaX188rKKxqp/FZgiqI8mbitn3r3fxNZIuMKk54Ih1sC1nHOamqtoFj
AbfEORjkUIQ63fTNKX8+B/mr0hk/QH5iNcU2gXTJ++1OpzHWLrZ3v4dfZS8op2HrPQ0In63xq/rq
yd26kelWZK654zxAghh8rnTfcpAuBkFXcC8o9qTPZYujItdBD13musm4Rsj2Y5ZuOlo+c38ByTbU
WH4w6pGCrCxp9drZu0FtyXTMdYrR8O0TM/D0DLOVE0sUDi0ZJXRuVx7H0unIuDGPjfuy50cW8+ms
q6ZKrs2xOZJaXUL5DeRNxXtFG6G3Wn/wGtysJKo/Jta1wKrvpbvjaG+I6hW8W8DB2DjFAJb7KPZh
34yz0+ZYIsjAD7ZLSAMJMelBPNs/WO8IPAA4pG/DSmCu7RQjLB3baksbmtLbRq1NT6sdiFPBeZBT
2zeEFpSxCbaRU/gFjUoZyqy22LW9tvFQ/T5T00Mi5P5612p3IEo80f7KPuQpt4J84CfJlx00Rd1a
GFX8yDG+OBFz5GlkH8OEStm711jMDOX0ptkmWlpV4EFZhR9j53R0m5UFwDZ7Gew8TVVhClbL2JNj
B/X3tWWLsIal5oK1sZbrYI9RU+gQGmJarUJHKFZtBGCnjuJ4xxu3xBCHA+ywrsTeb9NT3zC4puat
P3J8Q1NzjZkoGO1lKk+Tk3gnE34zW6rY3HOJnTpHEOuuOJKwaq3ElwUKWdxIigMjyNwGjJh7Q3w0
0223WGgOGDuoTf3MB7oEQ6qdwpT2JZ5nK094r70ZYKzOu2fOj78hkIOEI7WSPOQWlXcfkt4iMNes
67ex8ALnPgCR22gBByRDuK7s1ujRQ8P+5NXWlmjfo74A4IS34Ip4//PioPrpc1+bnSJdCNtSJJh0
l5WbsHx4bhqLOzorVWMRFpkS8no6jg5C5nQQEuZzgbsbwqW2q0iBhxG6yIe2L4hIbBOwkn6XOZng
ZW5oKo08QnomrI9qYsN+cV2uJ2zw6Kwu+QibOXI0CEIuXaTAqKfWZKXeuDwKOLjOeM2KGeH4t7ap
BG/eXxbJdqoTqU7KJK6SeF1F8B9fPE7VbeSAXeTxzvjyMQKoOVGai0D7b1yRY5mR4CT297FxHgUc
qENWMu0UCrehezw87HNY433D7anKVIeyUvZEbJqEYl4EIq+5jdgpvSTJYPeKv8RmbiaGFJuU0wt7
CQmZu2oT8+GhcKiS2yLgLydSYzuCL2w3+a0IYlh7YJn46qQ0zO7S2NmkMfIeewB50SWzVbEaC8bK
u4ZmWB7SjSUL6G3HujXSS2vl9r/GaPNr0DO+/plVip2EqWx+fsnVJjiu3WvCZMDXqoNfTXQZWDbq
awqtaYwu74C3G0fkvWpp1g/e2v6CSlK/qbrG0+JP2wHAOXGONTxNnTGObxKcRJzbQYm46Gw8hfJG
jPra1z14Uthw/6qLYPXYdK5swWyddrVCiEq+TblJjZ9UGO7gFcRyYqxHT11N7jVDeU1kFjhZw9ZM
BBA9KkONZBiRXNBAdAUaFoP8xScmQcvEJ7JZU7f/dXP1+MNOWNZ5vGiIKpW2PlRh1bx832SPub4x
2oMKJZ/xYKbXrulF0V+axZLo9WVDVPAXrgn8cadl+49ekDPzaPjm0zeD6V62wGeTeQDQSlUPPeox
L42xHgCpyghsR4dEJPrTVDME+SvF8cTzOW29OOhRAbBFmjRhF1viwgnd9BfckEduAWbRuoM7G8IB
/n2AzwwpdB/EYhskfyYQP0/ghzPmMPWKmqx9JwmkdhAAcj+B9Y0FpNGPnLARLVhxzU4T8v3rebZG
/NludL0OM4TJ5d5/mXUnrIpvYhH1YD+kCsjlmVzxt5CsayyepnVwYWFDz+7WVpFdO+q4QM4JOBD4
Il6KIuNu96TxA+qGU7zBuwglgx2ynHFm+o9AubSPvc/a5Okd3kl46s5mwKluSa5pLiLtfyotxv8Y
E5+tiiUD4eAnZq5VzSDRFaHA+U3m+BR8s5pckONJUG7+KaRdVv3bAu//cHgpY8/OXjnkRmpd2pVF
W4VEo03ADL4mDKut16HngxX6iF+IL+2njy+aAWcZnT2kSlKQyJweuTIZ6R2YRVJMl7i61Z8uJg1c
k3N5H4kPMeDLklX6BJIrTTyFzHcyL+QyHyisCKCND7Yc7PyJBqK1OSWUboa+q0t9NBvvqh+Djuvz
RB94dcH9YZHYgd+kjnOnzwOjw/u6cZMz4FY6dXTguDaILORGXgEZ1HqAje/hU5KKLWTjL7sTww5i
+0n0AGD7BGvz/VGvY46acq1uPnQRJVDOHQG/f2aqHRYLooI58Vuc5wIqFLJgurqvvi8F1Xv9RwIL
/cEzbOMBP3Z6f3bGuzpHod0UeXlmgvG2q66yYzVCzLLXso66YMUmA5BFErOKbXEKNmaAh4KAeZ6Q
3nuFLwB/zfiKSyIA+PW58B9sFA9sAOvTfYvxLmQWXK2HZN5lBxhNV62YU+Z+gouT0uqfbeLEu9FC
3D40j8BdtE9H1YTS48J0hNn2lIv8bdQoYN2WM+KM/xq/kAKszDiWrYe/BLcCx+evjAYJustD6rFz
+5bSdg==
`protect end_protected
