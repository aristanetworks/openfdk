--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
k9glzVyIyXKYV0pAqyqva8WLgTAm3x8hi+l5laaNf/E4ubl10I3JfhvZSNympbJTr1BwbXhapWV+
oqRGUU2+Ti3Y5cfDMNT5qjXRwTeyTdQ5YEPZYd7u/Q59hYdAemL2IpYIltVjD0s/ECAZsYvmARd3
u0ANyAS0VU/hIq8V7M99PGgqBzob/42es+Oe+su8rk2nPe5RdLx2t73E5JMJmoErDiQpvwNGXo4S
lPLTdHalk/n36gTLU4CEn7KW+E3bWT1rd0+A5pAd9q8GswMihy/deKW1FB6wPP+2Oher/hNyXYJU
MnAqRVjbS+hA6cEYk3f3KvB7lJ6Cf2Wja1kNXg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="vFVypfSI26eqMJphsX7Oaq+YlfGxtWaIHXIRpDBQWYE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
GoeXIpDslCnTPNvBagrtWpO3elgrv6YlFHArdcUDUNXxDScygbD/XodA51i86XdMgJ7cNbTcFyja
bmeqiXI0CBs/gfwbJBrkMXZVDyTd27IeUX5kBAzS+S4MmygqkvMhcFaUa9jcHRWgPvFBTsd9pXHz
AZkOR4a8AGPgnPS1jRcuKyMLv5/9mxjnrFv5k9igwt8ANImO8Eg+e1F7OuT02/F7JXf/1dcX+mwf
WMom3/bFG6BUVtQzzbXHKpoNYOOpo6Eerb+hf68fM1V5c4+e2GcLMk78c97clRGLvuiMeXiLZ3Mx
IsHPtr5x3V07FUz7VFf390Su2uF7XPCz/0NipA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="uNGqyXc+b5yDdJhNNkxFLoS5arbVklL8gztrahoeHg0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12336)
`protect data_block
5GRmFSsg2/cVPdX4M3o5SPOHQHQjXkD8kjGbvchO09Q3ZQIPGiA9qvWCFjxoprj5EZijehI0mwDZ
XWG2J0Zd+ORCO16ft128r9KHk2sN+XDNzIY25h9zLRoJg217dUBpbwWfaYur/u59/xkzFxc+LZKT
D5Ki8hOe/f8KZd9PSghe7rWdc3YqvQXRnj5hKzkgdjh/BeanHiuV4fSUZqUvN+xU+th7G84l5UH3
fRtFar4AxhuLs/j6b05CuAfXANxqjofujx82TnJU0N35S/pcgHMi/CYsLBT13+oSpqPOHzoi4TUm
nfQ4Sj2zULPQpUi1ZWitBukKwGdTHxFICIUVQeVB6UqagX9lUXEwiJvqI9/ctsrT7/NZrDpWdtrc
scvBvpmFBObjidBq6TZdpv5L7VO73TMufNBeals0/igd0sj4fs7JFCj1HeoBYZ0+9I0I/ysekbex
Hs1wC2DJDL2euJcOJ2DDZBzHyP5WnV+ucslBkeXzqGX8O08cvZRZENRajURaf26FYTsuV0cDg49N
70TEb+3ACEdNi2sLcvNMinMq4B3EkVciXTnG14YBiXQmZDzRpf9N0vz27Dt0rmCD6gtv6toNs8V+
m68pn+D9iHq3bkSJRd1ROcyHV/AjzGfasuhtRWeP0BUd8SL9x199W78v2wjMv9m3bvbIqd6lkric
wZgux8igaKQgaOOG41/0qr3gYHmIpEeRcT5k8DtShXMVHxvgQpN+rVANcRVfUkHIkHJYPmtJ5nLj
tBr/cDENUkJsujVa38lcMKFWzraeqw8cRmQHPmN5LSjseyUXrFHjH/sjU3Wfgycdk+jrPlDBOkJB
f4d4M8OIgKDxIaWYsUz0RYtCPnhInxRdr6u2BzMTHvOYeFAI2xrsq2yWsuyiChT90TohiSqEU70H
z5UDKkGf3P6jRG85aAHnqFinX6DEW89hwRhRJRDioC8YQwvx6ZgfhOoCQBaD2T9YZH0PeXi27zCJ
9X00R1TKVgzK0uzqiOfLcr7mB6gAUxzXUAnb/ddoVLtjytuho0g7YNm37QHZZAdvrUkLZQAMbFFp
2KIxq6mL7QuIBYPju1acvSunCL0umbEnpx7U6XYU37H+72N4f6FuTTsw9zEsCJUlF/Lf9nQnNr4a
r8mzwNVTYyRGOVyLcdOEJcxj7xNuMIjz7QFSOo7L1Ysut8/DAN0iq55yAuvAhJY8DPE9AN051K9W
+wn83650pjspQcKEtnedm5BIYImHvflUNAxOlsfIHMShZFaK41QAPJ8z1n/cw7qbYAdOeOs29GB1
ihc6TU2Fxkvk7w6HWAg6mAzyHOV1lRBmALPQzb/5mnsTNJYSfSyJyA2w5Rn0YrYVuymacjRLQrMF
7UztN1ii2b8CTdoEA9H506VEI9vjoH+BB39AX0ziRnc/9PwB0wrFFlx4nYkIg++Wia6pUKI9yeBp
/GePvSk13nYkjGoI6MwrJzKegu8ZQNOcMXa2W/oZEVtdhZvfO7SQTKr0gstekJ/Bx/VnVWv/jN8B
QAq8tUhdox8vZ18bTWz5gkqofA7NZVNWOsPJVKJVpo6FEncjPcdaHPG0c1hmxodMncU6waxkRuHA
qywgh1e+FtJXDoUv5OT+sYLBXMJmrW9RjKGKY356jyxNj78k09L4P2vJ146CkYyQm1KF45I99M7m
r2j1aYOdXyVNrZdch5TdsGzI0UBmUgNXi3RVSzPrtZQcCFD2/RSdA7ZCoiMf02S7LVUWbCHywqNM
w+wpofYT7fuSy2RJfR1mAcI59VWSODg2/sJE4qKzgyuOoFdDA2oG+zffMbLmHkZj0NKO/NhOdenk
KXAxGL9IssB0irumaVB1vD4alvUCgtzL2Z7ba3d+1cAGArP49KxtqGxppHUsZ0zcSGNJDtHFRxGU
rK5UkMP5Hfj33cBvNvtx7CW50wEEqTEI30lphl+L/vN8Wr7iInWsAPkEQmlysMGSJsXN+KGCgHx9
4Ea/3fQXdMAlxDKN2uysdnGbEVVM847VNji+dijMDY0LcJqGR4abUjs2bTWvjDWSZs1BF70b/84U
kKgeMijvZVlL8qXO0ETOFPJHQzfbHkaVJRCxta4tebaKLVclFGbuGiKXFlyOPgqkMMvfT/ZocTdn
Dt9HauM/adAieZZ5+bibKMbvGHgsOgqyUEvwh9vGZYM+qz7V24XCY1GdoP5tVPSChKzLcQzz5Tqq
/j6tFzpoYDCY62xXIxDMikDFoOmGbSVuvYtIbixKe+FMvdw835yZrgdXb5HDsvWqqukrw9FGWy4L
tVMFuuhBYremryhQyGsk1TH96+sA/mUN/ACAypeWJ8YpBBRARubY5pjNW6bk85bxx208jsnWTcTg
0r2ehsvjlXkNt3ADAqCZ+WYmG7FZpiBl6W/R7EGj04q39bYGVul0IQbCA8GPMV95qV07zsDLMTJE
Ew9hvPM+WAmD0Uf0RIr2zTjrE5UH03RIuBg0aY3RKgCcQ/Ib2EcQVu7OHr8foODJ0Dqjz0aUBs4W
kSmDg4p/kJaExpiNyzzcXx6EFd9Ygw/rBTZc3yPEDwmIpibnIe53Q0yVVZBuD14mQ6A0dZDmZlSG
+F7ONc3u/PAkzcaSn6QDj4McfcnpXarZ1/zx50gyloSk76NBockAlZbLCcszaj6Ps1JbKn6Tuyp5
pRrkKwoSVqv5EQ1prTD4AK63RSHn8kSNJE9zhqbr36KlQcgeGioult8FjPwFDkdKaCZKhd94oTgj
gvukes2Wuhw5SiJA88L5LuDUJMaPvwcxyKgEJvFa4Rc2jgjbXGDWKyu9aN2RDoDM4Bu27aVa9kCa
s2OPyazG+URjMVSyLUl3QxNlHWI7i4xFqRdll8BvHGjTAnCQljQvoRDYy6zGjWvBT0RwJybRnedq
izmrMm0fQBRwy4xcsMqgPp8BF994A7dm+/rFKrkk4QYxL27SiO3FzPEJ/KqS26o55AS19aHcJ5B/
WN3/8kizcz4dsZBGtqTtJjedoh8WEDW9IJ2qNExfI20AmqySoAtl5TZtN2QJcNmz7t14r05Zlvrt
r7DxQ2ZAuDBRHCyxw7Zl5fKDknvAv4HEHXISrE1uGmRLVBXJT+UwuDHYEt2QWt2m/RpCFp2rymQ6
hEPuwjYXzSB+6cb7587clROObVSOeM3fUA83edkGskuBvyZcIa/65zjtzwyxGu+8N8eOmuGfIBxk
iBfBiNz7TWqLcYJL/WHMOS0px16k7q1CPB+0Gb0IxzPeCc7TSdH2ZbMh5ip2PUW9zm/Ad4paRtbu
5krLzgSQ3vJfY/o/+knyzsBI/pOhv2uckCb+dHmakdQ6GuGrpNe7zRygKUAtjdWVbGw1sxF8OoCI
aAE0nK3qeN530O42hJpImPEwk4yYVgnKR0/GN9xXkuZ1/imkYu7P2X5Lj92MYtdfkx3A6vWTVs5G
Cd81He5Qy8mjLNzUwgFD+pyiZnbRF5DOHbSQic+nJ1YJe8unPxaMqSYXVx2jy5KhxZK1zKhbdKY+
/ClFIb+PBZlhOTvVGz8ELnDWYyrJKHuOllO0c1af2TBQO7FwBVXJx8x5KOdHnn92pXT5TD3N54Ov
+OBBX+tL4Pk7grf5k2k9CqxNW0fmjZsq2eNbppKsVualonk/dCkbGZVceZWkDg2m0LVcLUMjYghh
6Ux1Z9TgWRoKJufskfxzoqMg+/hyxpBCk2oyu7Z/jXNXnHBGMN+faZg222OqTxcoTJFyChoT8jMi
42pmVTklNK7b1D/GXnuKBETg/BDh7X8pdHMl1LKeUOec77KE0cCJWBKjiEstgcGStlRhCUizfxPw
vjmW6WipdtdarvVVfDXQYl+CaNu50x7Ck/2nCHVy+NW4hUyrEeC6Bm2T/IxBaeiQwY9EsLJuR1Sh
ClZnbu9iOlZOdUFLvzXBfOcAAejfYgU3JJDQN+byJOOp3zHuBiNdvIEfDNhA0mVhWgmIrzfAzlrV
NzZq0CqWUMp/bYEivl3jXnYZ60l5A5oOVytGMF9JEe4P6WXCfu0L2q+dcDssminO1cywmccJg6WU
PlaUa+jTI9puHW6ks1gMNqZqaVcNQ1rKkbC3IECJlDmkEmFuFzZYq3uFCVj4MvfZ+rScSmkSkemk
Jzih0mkQxBh3fD2hUZelVENTTNzSF+MHKU+gJyZZZdJ1L/rBdmbhn0tSQE9Xoj1n4VcJ07SnSVHs
QFs4F3bceWGpuf/hWJas87EexPW3bXjkWl6LwNoyorhU1Dw6ECmmVrZ7msDPMO4O6iVXT4iL/kIU
16Uc6ZmrvNBg7WjzElqEEX0UfEr/17l3slJvhfrx/LYq1IBgHByAudRofuxB6WZAoXi+FVkl3dfK
P6saRsQ539knxaTQxEet2Nd1JGKFb6KVsTn0f3vv++K2KHHoWBAYTs4LOjotjS+pbKnB9uuf5jFX
etOcsYzkCTt4ZWjU5SzrWRoaOnqRYY1NILKgH+UGcuTLa8HRRHzK13EmsIvid6xioxwDp1jW2pPp
RAiu38jMuPCxLKgq7Omca7nzmxuVU8Djtv3ZpFOiApxOWF2zpQTOxCs7RWz+aL+Pk3eWD/EmeNzn
Xtyt9dUCHk+DTUx59z9DPb4ba2hw8WZ/fsfdBv2dXG2luA0unOOLx5wFrFZDKggI5fTWhsM1rPIu
AXJ1HhFMX92VwNfe2fOuKVW0nr2PDssOyyNtguTnzwb1eWA3kyARF0RmUOcOGAqJ6SZJuXY+/LZC
nn0XWqE9k/VXoMxULGEiO1RDATMQrLtw7VuNo+u4K49j8tcQIP9ohMCigY/49ftNzxjOV1B+QpMC
sg0v3B1T5YhZkxdM2hMikRJZYr3NzMnwZXYNV2d/80f/DC4T2I73WJ3c1KdAHc8BfFTTnjHx7ynf
eAVXeS1XtDnlpojpdDrTuQXC9j/U3OVW5FJoYDBbqEDlpn7am59/RdJc6Y7xW2kNpVMJ+ExGkf3U
sqfMLswF/5eXvTDtUNm5O7xpiZSOhgSOYH6thkO9xo/bOaxMVl6KJ0UYfLrPxnUrois1s2ge2YLI
E5goDthL4QOGW96q+RRyAsNgN9WNuNGYbdIkUkOVO+p50pD96gSOfhy6BrkDBDK+tmYt2ldIRpI8
ZChy75uMxLhkf8K00VAFziqjGnKzaxuSI79BgqHcIlpjY2GehbLaXX1mJ7Kq0nDryftYSmzQ3GPM
gXyNZIP0YAOAO+KovmzM7KOntSq/wy9YjwZJR72pknV2VvQAbCfnTBKu4jFCxQEHlqfvh4OKKKBb
TM8qLUboezYIxa8JiscjRY3vlywLY6qBsAfmNgwHTrAGhtS2oJ1oUHxwoHBaXVMh+8pRNozWhLs7
0UPTefGn+IDKUqZubtVMec8WYx2cIfaTpwDyhzf01CYUhWTRtsBTaK0KYJVWpNoe+68TZvnxIp05
+TJTcgzwwwxdeyMPfIeV4iA/b/QaEkvZGmZcMlXtphWjgllSgKquWHGtrCOzWQLqZors8b6VBz1+
IbrSnLlDqd9yBMXxGabY6+7k2M1ZEz9xPL1pxXQNNjo8H/U7XdCETDEd/3RxxpBS8PafLI9833Ng
VhMG2Kf7lknhWuFfTTf7Aj/ABrpfI+wTzWAoGo0zEYgY6q16o72+9CGPDwVdWnKT7ETYDqlXiJzq
30taC12pkc2lg4AOSEOr2A0SxCyPh26agdl5ultyKqjXfP90oiefpp/9gPtblzRMoQOB3mbsWHL/
WdTl71l3uSnDqs7b0vE1zKPBgVj6E4EleEd0cSku4dm1lXYn7xXiBEaPQgjblcMsH2f6ptiqlwgw
WTa96ixppUV6P9QN0GmI2dCJ8IPb3IRvJEbJaLFC4suTmAiJEbnKeuKvUiSu5598QBufEGHYa9br
AkbyVdJI+zt3AvmKIdLuaS7cSntx911Azk3Z4GT1buBqzHl5dWQoTE3RFhwfxHQkJyhXn85Rn4EQ
bDV0AzeqpdKzpwGg2+JMhOB8kHDyXo1adYwDySdPoYjenOJqNmKICn31U28+rYv+cHul6hNAjn/U
dQN4W1nQWgnfJEnFuptjpzGcn2CFCiXxYX/VIbTizw5XMIg6kL3uN7oYwNf2R6ZI/yo6sCOerPGy
IvdKY1KuJsezFl8AfOIBDPPUqbSwl93gkGOx7rBFlQnrrsb5LHCWwivupWKZuIG37KURJybRCyVX
KZvkDjf9KS00P9q7X2OIIhaqQ6u2JCiKezQyo0njdZR2/Zut/wykinqvLUvpNwG3WecjS6he1dUT
8m7hPeLyStx4RsrXIDi8fLdSoQqhYf3GqbTGsDAZVLLLJ6sU2wxR8SOiYfCSNFD94us9P/gOg9qb
WzrWVN3B/Ln0XUo2sxouQZhGzqBzFFAtHvvOzFxjhZzpfaXLRc5xW4FXj8MdCVDbHJVSfEKxi/Gm
LiQPU4vt3MQQKrPY/L4yPqnTJD97QO4MJrOG/s27O1TWuN6bCOnvwuKhIAr3qDavZpPeGhS2hPR4
uTkvYMABJWZBzYc8jPDM6unUGeM5UinZxQ5lyBwueOTXRTA3N9P1wtQMHQP9AaBRgsre4AZ1ws4t
r+N8hc1w/UajT8DCHYv9vgoaWaF3yqmXq2jD3UD/y9M25av+1KYquHiusuhWg7QfPTngZVvj408a
sb2Gym+ftu9KvFLmQ+MsaRWJ1Oh2upu5h7zO7/RgAkgQP74jBWEIwN/zzQHDoAyyQzNlNmZE/u0o
fcTCqL1psi4CzrHY02dJzFrP5uBoQ5+cDKIqxXGdbiBTqQb24lPbJKJ+bc4PWCRqdaZKvrIj/3Cz
h80XdoJgQkz5zjHHLt/Jfj0AovW3tZu2uxh/B6nWWK+5hHkWcMkVzqzKBSB1E/dSBoN0ID/y1hQS
yojxorYnrZOGt59+BJuwAnRRSN7kSaiWUQQ56ytQ8iMMXUVtrrkImVRXhIpVE8Y1kQktgQTY35nL
j1ux9P/VzlJIebhyJcnRJ+20Yq4wIGxvMKMF7h9IOet2CDkH6SwSTOKGonL7jN2jV7ESaeffNUxx
YhWzCpHELnNLh5G6ZlZvAUfw+X92Cx943KaBQ9fxP8AUoM69hXZHQMjgtxujUJQ7IFeD+McNZ8Pn
04OXgdX6zEsptj0SJqpYkcZSymDbdFLNvVSgzQyQwo2A8vl8ZiFGjJwM/oELAuA+i6jke8DfbZ95
dBH/4CFcq8HMyCZMAUhxU6EEW/xcAiCaS1twh3Z1LdvC/GM6dWPbQJ+2epIpwZFh0FDjVOvlMjqU
ORHuqG9VBtJAAknUZbd/Zum6qF2bVNuCdCJGkdo1PaSxj3whHEkzCTnBVs3k7kGsfeOc1KeMP3s2
R4xpsG1cQVVjyfRu4ZdeOSi/21b7eiSWmGM4dE+kv6DmZdPO3E09YLw+S2vBWudJ76HFbK2NAFa5
fczBDLikW46ZCj0u5PaF9RJ06ZosbIif9Mk1uyY29OEsuMNctXQOXrB39uphI+zaRI3EhJgM9aqr
UQcoDjWaRlclYsPu97AxQMFK2j1lJ+1HAqlIlzFIcY3Aa/vR2IUbjLGGv2cBJ6cn/QaRl6xQqdut
ZMFkQxftmfWH0/1X+GJRnCbJh3wjzBJqAdzGnjj4ZSFfi9Olq2tyy3Cvw6nG/8tIbsLAuaLmdlIS
23hc3ywSlK2cnOEHlDyRBXtXBzRqIzPgtEp6zAX+KSGF9e4aJlJwvkM9ufH+ENyp39NTqZVg4wR2
CzQ7sMrjYO69Nj46xx9XJcMjiZB9wDJudcyXwje7UXbACCfDZPA+D2RTZVNLreHjM1JotOhi5OaI
LyqQsb/cF7o0Ll/+sUx9yWJZUZG3tZHUHsVXUWapulNkAnkJDG0YLBE/7Nsl1hrJY9QeDnKnitrj
BfVxSCts9sy28CC0u9ax3fUoqMlNFtcn6cRa0Zt63YjjnpgUwTOqJPYc2vvkPy+MFDu+7+4/08qX
COlE85ghL2EdS23JiD2VgxrXZZHzj40k8KV9dFro1AGD1KqoTkthVxIfoPrdgjCqdBxc6IONMS63
X3mePE0TJjj3CT0moZZAyJgD/Cw81qcFXfodRrGdI36HUZklmaf7Od1+3AzPDi3oAWgy2aWUybNP
072xHp6AIYSUX89JbV8l8d9E3GDS4ZP0b0dGE7/zeOg5ro0AAoQw5RB4+sdBsmZ5Yq93LttV2dLW
c1iV08tMfqPiQoaufQxbmw7FCdwWoKjY31xbHw7ePGOdj+1vR5SEtQgSdlHsfIMDaIWfFhhhhYfy
HaD9KLoLTlyPwYyw/NIUZmhORQLIShvA60evGdOS50zMjcWzWQH4m6I6Q1q1tabzISjq1GC1PDtp
XEdpJKpoCVLPR7IOEvTaYroVJvCiHF8P2IaTNho4gDHvHB/pfuLiejGJxEjwik8QQSx5POvYSQL3
hdrIGkgsRNmEUC+jQ57TXv6qHAtbcw9n+6wg14LsfLl4voYgXmxNfIvDgQouN8tdIx7PUSDN9kDc
0mvNIDH9HpUHMvZr9zG/t9zZY77YqcD0ounfMHQKWs+JvK5A16C5HOqvV3kkC2XEnojXiuUgwDPX
0aqHyapY4RjYeWStPdRtll85C0sdK1cu9AFtOYBGurKjf7koFHAhySj31LUK0R/UX9Gs+2abguW1
x2VqV+XYBrLLJt0xsC0szk0gtrv6Gq5dkhIN+fWyF5emc/mmfLO1cNs8nkg1swLZoGoB74jxSKYk
Yvqz/T+E5hDIcs1Tv8vTQ16OZvakjYe2uqnuPXrwOpO1aImYs598FRhTiLnwe17Tq53YDHwrqJby
6B3vFns3+Tho3JVEDrn49wL4ioUC5M7dxlbzBOXqiJvTswsNIXD8idLglr9UWoBjEenYhfSeW7aq
Psg5xqOy63wWT+cGEAUrK9B5EtW4zMdW/+kTWVXwPf5x0K6NiXDSZHAkusCPjQ6iJs+2hB/o5WGf
XjCGGfklbnTmzq5huZNDXsuBnMoS/i0JfLGK4lpuTNiM2ad9yniSj06hgTr4kiDwQEfRJjDT1OSz
QQzYOd+BHzHoflaH5QLUE+PtPMjm3x/ayiAemPJyJYfQtQsYDf2amLG5QZ1xmEjBTIr3ZjGakctu
d2nMXsevXKiW+K8L61aI2YJTsLVz8Muq5g8v34mnVqW1zTFCskHz4SIeda85/rtCVXXaj3KkTEYX
N3BpvAVd1rPyEvNjDSmz1O/L6kzXEixgIITpdGZJZNyz+BMGfh7IIYbGlylYC6JVrPp1reKbecq7
H/ab3pknFNMn2ypAob+mkOVocCh5jQH+Viq/YUZR0u3/8JxTBkQH92ohdghxAQj+oBStsbYfiBBx
QGjL4D4h3dhdGcaMWsi/VCH2rLxJcJSmlZBL3xkBjoVZi0LY53IAgBRg9a1bSpRWHBg6vPtzReKS
t+ii9aKTPy9mm4DGPCZd3IO9sXDJ9NoXtTG+BFaayVrOziQepnHInfGBU50q7A/LIrcEPaTEQurK
VyJzddC/Nk9ms2KRlo5Z1KPV07mIztoVQVSOi58Q8Rc/OQmWHtipfEwChwcZhajYsLfynTiJVqHc
sk1PY1yPMXB8Idf+xyRLHgxdj87qAFKpShNQcRcbjEAXv0VuxDQHiY1kz2G4Vk2sSckYvwKUgcgA
NM+m0SPxswQqAfDf/3Ikxn40DNcHHsYs7LY4SY17uFlQHLlAo8JlLYCUcbIknWPSpRANgT7cxMAn
5JzlMHPBYkHJJhN0ki3DCDVCXMIiheIjg+dyrl926fpAwq5L/dENNEpXJrtECnVpykZ8f1dztq3d
jX8KqXS+N1YqGBtQsCTPwq19gnYAHyT9S9YRYIHQgl0KD6KCxW4ZCJJnIkTDisiS1rTHLvZv+uVV
7JUy1YQie9c3WIf52H9U2yGCMzSPFzTFtYT8lE5vBUbf/YSXKuBbjYiV/YIDP5+po8oqS9C4PfLE
4s3xWZ1c7v8tFqzWtBc9tUijkpf1ji93MluikJlbUDOLamD3rb6u5Jfky3QCpAjToFLcKfkiwl2s
aI2CFWgiCeojzxgJVF8MskJnzDVN2ywGSslWM3wWoMKDkeDJ0P5xYvSx3GaQlYFnoP853zMRtx2d
VqvCkmxW6UgfM6+OzZrH0K7weRLooAQzqmJYS/V2Krc8dYkZJDFxmsYIkyuLcsVSZnKUxmHMDGJ7
x9MXx4ex0e/QQuFE20JvVNm0/lrbCtSqHYD4BEzJ2dB97KNiMUmS47vK/BTtarYfq4q2Z/BT8f+d
7mu679NEz7fZMkLFgI1yhbKN7rbKl/p7ioE5UllzyzatEaiqOcW115w9VcpK4pCNrlVzDRAFGKIm
4b7AWAhrBNMGAUDEjLYGj0q9ntZBVqynB2MICI8ni6wsMHg9p4qVD1tCtdmkJWcev+q76oHRCUyZ
zQXQBF1Zn7XN4n6CRyf+etMmoCrKlBvATdCRTDHIMToqUXc7ID9whGmgb02u3Td5+A9qSouLR9P7
obzbvMUJA4c+qBZj8OEo6+4P1iMAR9W6fLbFpBqdeeI0XMg6g4ZTWpPVGyCvhmKO1BMM+yEqDS9G
ceppYLheIE/f481/fLOU8FS6hUk4gl2neVM3moI4J0A74s//OasGbLJ9DxYtxRiCQV9cg9+NqD6D
jNlolpJs7T33R2PVDMyXaV4hhJTwJ46gtf0+emPzJ1cMzy+DITCypXWysjcQkUI6mltzkRdeym7L
2DJt4pdIGksIbqddvcIbJubaZ+Zv90Ulk/AH4k3gK62pkiwpMkwCfnJLJLEYKy7hmxMO4vSpA1fL
fru+XLEqQE0Cf1QdvsCiYmBZvkH3ZPthJZWiVwd384/57YpS8efk4TZjo1yKs8/hfv2tujXljgIN
eNoBZRfM6rHpKKEQLWJiOTOBpvW8rBEYmDAMxYmECJJKLaUiw0nLsP9/HeNhp80/Gp01E6l4RN33
cFRwd25Egw0AfyaarKsUST5k+gqizj7Oq30TR2p8pWLsCt0rDrwYVo2HQF6s/MWBR6y7VxD9FnKo
ZXimYBhmWTUwlBGlCNqzoJXTm0h1xwrSUZEOJS7J5RYtnxbkUTlIWEAblxKJWGONAXGpIqstVKbg
hmg1npG/849XjsZar0gjXQNG3yx4mEPqI/QBICJFJLy+D9KuR2Pbvh6p1vEUNc5EmJ+BrQ6XW0sV
toK0RO8Mk8vtXfK+on+6jfR/Mxcly9KHtcfKi4g/V9JnlMX0SCVJK78l3V8Nul/SqE1Qp1y/HAjm
R1yhs5R7pwa+SlmoDIplj0PdUKmiNOhd22vGFqzAqiksTG5abjOAIJD2aKMOPImt5K5xwMuHUto5
o+wx9OozCvvBoE/w5RGdIURnBLP1OHpT7AgFMMJ3JBVXZw82qKq91grHB64dGlPNYs7VD6FFBhoM
GYN5U7BRRV1D+JgUDVElX7uj1RIuRL6fago2HRDKuBTU98IaLKNMvKQ+jF/2xrRC79/LPQlsEqOG
Mu1kn6mB9uqUjK3FbiX9gR5aV9q90wWJaaH+JDbM1xzRiOvST69Iq+uBLdRc6LAbvkhNN7n3cqF/
VPXushFJ0xNdtLZpFrKUm31YxtXij65SEOTha2+Mpl02PPPzh6dy0wSbzBMuWllF1bbEE/j+O5lX
xX9zSOWtkhADJCmbHLfGs0qv0jMX6OitRGXsVM+bpT/r8Dn3Z/dgT4ZBewuf/yjWwJbekyek3Uix
txelIIrCnTKOJZC6p4KtF8+reoXfEotQbHZ3FDPl+XYP5oj3t5gCB/QkLmwoLdAQNvK03ITOG7Ps
Q9+VbIBHNutzLOyM45uX44/aOkMLSSlb1OdJovl5IiNgPiHY3a0dDKo+jwxevk9gVZjtAu1L9+tC
PauzfvuaSlIkslUN0o/u7v47mxq+DgziOcvukPHKj5vN5sZXMGH4wh3pvebOI3uCsjvKp0DgVG1M
WMTkQyE98K/y1B22GcN+ywMtI/TXTXnUAoH1Y6krVWKAY7AcZ7RKcEXQbnXgW+5MojWqTfFKKKkL
qY8HxkcEoMG1MnPHA7MX8U4Er9V/aRKKSNKDYMjs0bWteo5zjqg9QJqRNBSoOwbIrg7eJy8QiF6V
ey1Z1lGk/tTY7zgJZAvPa6rrIv/Ih2M21QGQyKpMSrnq6xQFRKHdnWMR88LKc7pWAFcafzSX3LuO
yALMInktc7dHbBid6dPP7hyK635zLicAkxd3szLeJDWxxQ8StkVYhQFRMRCBHC7bU5/FKW2rgj9y
fY5SgwLzs8oxe5vsZDvFFyO450nMlglx1DcVFIByq8UoOKtLgv/QYXOcHmIXr4uu8EFgy70gal7y
s9vRQ3yZIeIGTKpAsPDcZ1r5p9RIUMM6SxozL2WZGYU0OyrEy8R5Kerz4YtWP0L4qUZwNGqBWogd
fW7CrW47RYhMhMVH8ZVx3QYGDEgNKji1pv41Oaik4FyewXcO3pvf7KlpClLsokOQmOvDcRZrpNLG
xqfJQd8zXvSVF4cNnyEHXMYAfwC00pBCoyFYQLec+Gb7F2rZzdZQokvUoMTN7ShLTdp9HSQvVDhb
cqNgiFpSA7cmUScliS/pUr6tu681BMmlZba/AZFrFbZeThJ9wHWbj/iA7exqhnbKy6bH5yXWEY8T
8MyT7S9VeePnsE0haEWDm/B+YwZlQaDQPk7qvf92vg+TZ4a9mcCSUrHOYKb8pXylw756CX39iVdd
hq3Fe+8wv7y8yX7+6DWuZBYze+BvcFXzhtnEjkvc4v/39mq6sq7hU+9EpVEMAEJgO4CN1gBVuWdA
IJzyeKknMSeanxsmVgo3ygRzAf6+NyiZjSypp1QeSeXHiLPez+QPPl80x/dR5OrRRvFMM5aZqcD+
IIaEuJZaMhps2XjUMOYGYbKZBlEAr9uWeueIFbjwgcutjUAbvt8e63ZbjQkOqIENVxgQugYodxeR
C9eaXUzBD8zJ8SSB8as4yOQELA5l/cV31BFj+Fj9iKBoFJg+Dy+iEd4dhhKeYj89EwOb8XGHTaAk
hJPDYb0NPJfpbNHUAvE6s/E75qfGabPYLfzC8gDHzy8D3OsTGLOmdm1FHTt/21aiSu8/YTyxPkk4
j1P3C3nR1XGPqBbzFvV0BpNzbV/hX5/k35B9hgIzXCtEyZUUcLl5Ox3F9UqUeMxOmHaHwT2sHVpj
l2F2+sb0IIjR0a6Rp8g6n5U5Nd7eCuK/V0EHiO+6J2dhAXH/qm06rqvU/7lGd+2SYD6ytK8+5cHy
QaUf/2MU0rcnyfoTGR0j4bvDx6ykarBcT2jXeSg+5FPq4hKrrfhAIqijtR3IO+pSOMj1NuGbvG3B
iKKZK/zb8qLtdjl3/CV5TqisuEthPewGi1bZIyAj8ntCcZZ/655gHYOdGNJepg9CUHTx45s2JpNP
w1mIEizof8Woy4suzp+LIJkE2ORA6LhHhaOHhINcu0EKS5HST0ryCL/LBT3CC8zY8Oezu4iGG50B
cW5strW4z29IKZJkk2NJnKnp0/08iXQvpTSs3Z2BWOpG/r1g33GEPd5RBRiG+cV3+rmJXQVYRjR4
GV3APex1C8fZe54hCSO3CP1ZB5eUZkE+EX1eHHP/FYLb26IyYOi7z0moutmiaH5Oim/HSIKOzLM3
SyDfuKmtnrd7Uh6cJMmfPX8sf5N6F7iX5fRaZaFcxdt8QAYS+oYGHNWNTTkln1uGYCv/OaGw+XF2
ok3u3lVb/XfQ86gsb8oZlnQ9ZA7fne15ItbkRQBFTcX3UrMcTeZCJmUE4NrKo7k4Uy4FffkM+rtQ
rJ9uXjiHCidn5h4qGTYSJYx5M8MivcGVGTkhkFgO60rFTmjRGL6ytv6EW2ynoyj7rQPMBti0IL2M
ITwFbl4RP8hKmZmEo6SJmhM25/3VLhvS3xX1itOzL9pHlh0NmZz053CoQFDcdFMoWmk6lDPzZUWh
BW+yxNwaL2QmR1UmvxHHjCSUKPEwAQrVaIgdituOIBSBgk2Vk4L+vShMZQZto0XsdbSyik7RamXc
5RjuNODwWr9PZilYJ+KQGrOlZo1QO/eNO/Vv+xymlv+sftdwcfHYsvDuGfpObk+0JgQEiVs5wjTG
xgvAomOTswDjbbiWK1FeG/Epz30X70hFqcWeqXUmEEI3vlhCkrGVtvwLEiiF9PjkmXoZ1JwlDFwv
Oln8mHqnGjJ67V953kaGBe5G/ZD7k30Ns6NFOTVsKt8OwTh+EHQbIAlTKjZLnhHLeIZhjJCzFGAp
gw/CXrsVHzo7VZ0KqXzXhK+Iqm6Blz3kkGcaDqHUvGfJkAP0tFA1m9QHYt9SOe3www8tvMHrkPIJ
aCg9G4SeBqsxTJK8EnoUF+RonwAvxRlMmXdgWUnUHhGz9JftK31JPpQPvvKN9ozhQ7fxB8bzRSP1
evxFA7eKS6aEqgFs+fFGvy8nFtlwkA8GP/ImRMwOmqkSOts97dXFQD4G3k9F+r08Ic7AYSkB1tav
GzIoej7sl1+azKqwT4mbD89bZ4WUfo9abf9Bqd+qlItAwMrugA4COEdINTeoTgvNzGP7PSvDC+yg
ZKc59GaO23QPIWPI/mbAUxQdJXCSPU1jp8RSDG0POlHCg4AK44LHQvf4yNQqyvOhdD3QUWp6KC1t
AIErbXI7vfwE+7eJ6x7iX5fpW/1cM9mPQHsjyoblVOC4TS7nyxbIcHFxMhxVXtgSpNDx+o6//iOQ
vKNS0Xzj8AhSMj3jX5GMdRT9T7C1Zmp+GyRKbxxtl/ZONIsf+nPwS3o4YIjAsdFu2MxEsLng7ltf
rONr4f+pvhzv19pndCiTRiwB7n05eDNJvZ1to+kRa7QEZ3b6dTHWyc+e9chSf4RkwD7bVyCNgYVM
Y82IB3+MHK12Q3vkGIG8vWdKse65srwF5xw4HyLEmLpWBEVaHQP+vpbPMpo00JOZwizWmMLf6Sol
djR/YZaDqYXcoXD/dkOTAAr25XpOdGY61sNuO/zgkteLdGL5vuTgCOiH+cF4/ypNHfnWmPIlikNe
G5GT9oT+WIJndlpBb4xb51fEH734w4OFq0dEVq4h+6OH2f25jCkRk9RfOLxcsus1MgwOwBY9eEYI
cz9pMvz9H0exXEhev2YW5BVbxOHpHdi/DkNd8ai43py/tuYPjiMQbgsYo9CZoohDMCq63r0LZ9Nq
s39UCjNKOStnzc7nDIcfVHiVTxI0n2rmMfRxrNGaJwkCIxH35jkZVrC+AKR49CoL89UU37r2s2IL
Sy8Kytgdg+o2ymCwlEvksqSdB0CwPR9ajSENBC5xGEi/+IMYQasXjHktWr58RBnOK8dTK7SwIBkV
sJzPi7scQ0zRyoQvbE0QLtr+sf5JC0tWARyfxYk5a6ehcNEnN36n4kE/lUrbLGyakNa9dd7U+Xa1
QT2AHdaKdUhff+zd14ES5WUyQ1vsFMcST86fp4UIwW9Bm9bSUvNppk4sXceVpHqN2Hm/RBYqpRFm
yQgAOigw5YL9txonlJBDqt8p2Wlq6IakCeUIJsDIqszjhAmE0t7KOFAWjBrUzrJFs9DX1qSqn/UW
rckLLRTWrnDU+uB35aOZM+N8b7UFISLuYPS7ZSC6Y6/OBlM3EK9qHDISJ7eYmBvIT/1RiYydsOxN
PyniPFlSrgMEFwBLkMkfLjuiV0ePzz13NO+VZqe1IwqYIozdpayy95yJdgTToJzXs7RB7IPrTF72
wAn/TRYysq1OZPLwzLo354v+Ev+7nNTzHw/GqdVJSy6Ayu6546OrsCKV/kEEvwL6fPpNfkosDXfu
ZG7nlYZHKjcmUlX5GG7VpDZYz0vdnQ+cNIpeZzhHZhrIqBjPZPkgCNHLh26YplaPbUZEC/6cCzAw
5aeZEcKBwLKTnpyHR75BDugiu3pUL6yayJLU3MwCuUwQTMYH+kcOq1KEzBFP8F1yYTV9IUIn+C5A
XTvGJTXurh93NnKdPWtMUTnV79n2s8uDyaLd3qwEY4DZB0jAuvL1g4JIBNAlJteQ5P+y/pUBroom
mYYN6/lytaMpiZ92p7dEScQXzCs2mI0a8DZXXIVjnXfZyzaK5BzpmlEzi2VMZSGpNuRUaUv5QKm3
hBvNn35DVnPx3rGFJGXK5Dyxpn5jrciHs5pjH7LoQbnHFGm+rsWPSA7ynNFl+av9Rdh196BjLo0B
l9zDEM7liWQViPrIOOsioG01X8V3E8+kPbJm25qw3NogBrapKWs91e7GGA/qFHAyoKzDFXiGjFeu
ct6wypmM04G648p6yslNuBWXS8j43EF/8nK87dOXPPNKWajFqw9Yg4rrLDzUiJST4foc7kt+yshs
+x001VApJVe2/Jq/JvmD2//BC1eNFaZxkQASbAvxdoF4SNpfyyk2LgpKq52HTW7+Rz6rHWbilAm3
H4xkunvq6A/9dlM7jVyj1ZvPtzwrMM+IZ9lEpLeGqVQPRN65fqpWWW3QN30jFoYN39OHEYEen4ig
VW29xvoTTd4+chHRHOJwD8b9VPRf7/V8YLP/NEfkJAACQ/03LnXvhZ8bRJpA0IsZ5Vv2Y3Zg1yS7
LhRKnYYVNszcPDG3qPgZ0lEkxRSgJeW6
`protect end_protected
