--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
aqDWnzIJAG6/PoKv5RGlHXaxyr6a1G8Vx39HMueJrIxk4pnpexAeMRUcAehOxIcA81ZjufI0LCXT
dv5oZ4QFC45IbFc3GvaZVM0ud144Rf+jwlmvcfEy+9FIxRvG6W2ylDhhJ0xQpPxTwaeCmqA8xdMv
QCFfbxrxO5QIiAdM7fDdKfBgCST+37X9Si5fiESWA7kL1rshnlz+qGnN+fSiE9HzmI82mUtrWsv+
iMuFIQ9cM6S4hkPUoLkrvQjvDCG0JCaL1E5yVvZqFeeCeU5NdvhLPuc4oS6nPvXLpw9RwjFwq0xb
XOozYOg6w/8h1tYq0fH1qw3ZDj0kscaTj/WC8g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="ghtF25yyVgWkURWgLF5WXKGBglp4sJ4WZ/7nn7X+Blc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
ryBYyBA53F4z+dmz7Hn7lMpob6k8zgMmY2LN2hHHEMvIWWgcmw5yhLzk9ujAw16CAQgZAtG2P+JS
FLJOZCAnfeEK+dwd5frG8+SYvBsljRH8OCVxTOE603+PLjy9G7Tj/INjfQW/BUvOm07UUTrMFSoQ
86S6q8JX4pBDb2qEp9uEqAc+s5YohEBuHO2nUbJo9+D38Wedgm9tj5RfZHsH8RmDshFk6GdEQofy
BAsjkyKFplpqGd8PRnNUC1uUFzHJc1KNAao3g0G9/uVra3Hqs10jR6S0JEUuTTUvHAMkkkskzs6j
LXekPKY+kQ2p1nfrwJ5k/XgH9Mrws7J4eYg0pA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="9jm7MujovQTY8cFxwPWbaACf7wEmdqiRzMBsfGmxJ9w="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4496)
`protect data_block
81ijATJKe0OtF4gktnV+Eczv5p2sdYCGi1QP1SYJkY0VQn0c1jIbAVzz28dlmi6dJJKANnb/hxEF
L/Ge+CUopOWAFZYwJYXfFrzJLrc59BxWygyqqj22HSsiGuFDK9+5Z0YJ9/tw6mJr7dpXNFfAQp6e
tlVZdLo/ohUQR6YfUzjjYMX5xwMOt1UiWCKyMaLrwgNiesL4+9rC8tCF4h+660xJEaxnufh711nv
ymDNX8ZGdxbssmw15JJjvxdvya1ostC696Lsdl/0Jb43XZX8sPBjUr7oUWw5PiXrZysrMJWDHbmI
Mg2K5DhYwwhMWsuxygSHY2qwDq0NmSyQAkje+bqs89VOjHrN2af4hUqmnbRp39xdwFyo+gVK7dH+
het6SPGNUD4zVo7onHHoOfL5s/DFis3r7Rfo/UCa47S501xEkewT4UwzEwmmmU5G/TL/xeP3JbvY
lruJJp3RJRUe66qr8pwBiipNXQnHnhg0NNGCCG2J9TAa7JZikLw0LcFs6zTkqsqVycpT8sEc/Vmy
Qa90UROzvXbiKBlFblC3SPDNK2svd0Kd3bIqgkk5uqh3PtEn0o61NjSqHkyImz3j9Gu27bpXKvGI
hCwD+1tywucWL3EJKga5X1m3FnUZ09HA9g6y4bx+HX/kaTjOrhlZxMYBjQD22os0BItT0T/E5uW4
7aNgGV0Es6P5aSZEsPTxz3Xj0T1HUducl6QAsf92nfC8z0cU/ufQT3T8r0NlS29jBAgugodgx+GF
xcW6PdlXapri32LVbVPB5MMBldFMd27sUSjF+dYprLcVGd5alHZfdV09rVIPejDcC98OsPWJd6Yu
Vj5qN1kH5SUI8n4ZJ/x4i4QA3LVcM5VlyWEL7MiYwJd8YMoCNGm3z7YC4jl+U9AMb5p9vm/+E6hX
8KPDOn03u9405abiLri++NQQIaWuBMXaZxqNlNMBwpoKMW5WP49kHom7OFeAMhXDvm0kz4Htr798
eS8VI7CR92cd/XWZ5URmzbPuWMq50qwU7xoVbVVOQ2l6fznN0GKbCDoJ/YgLSXr222/dF5OOYwBl
mC99iq+FTi7ZRAfG87TFu6cJWbhyefEiarOPqSQdSEi37eR7nGTQOjLP4/tpNV0W/UzcH6JvY7bc
OY7RBOniJW0JxxA35bJmo4y2Utfrp+/s1s4CQEMT7/buRMaZVqN8yRmvMEHypZtCsUa6eI+XQPjS
XzI02xfgNhvisuStaf5NsedDhSB9lfnr/nhLTr0WtXQ6KaifyUSa0+4jw2RjP4aIhYoYMtaREC4m
s8l8qqJXjJzOMH6j9aGPKUyqa1rCYdxDuoVjPhOOjgYNxWE3ydywul3+ZQlnhPp5SQa31ZPkpbzX
dAW37I66i/Ng7ss5d7BqXoDaW2qQBHLavQts7UVbRTkzX7DjHg6BEh7usKmFaaXRXbwevOUpp1y5
rKQEZ1MiQZTMACAji489fcnSfaumv1bQ3T/vfnA8al2+apr+7MiChrJdWqokCDKYbCm4beCDmjcx
JAzLlVX2fNaUxuehNiTLh2wWJzEdJZYQMPdk5l88GuGWfeS4vJAB6ftdBl+D4Zh/QQ9oxWCUCb1b
nyGAqoo1HKDo6japDD89hPD0noDFZr1R9y5mSDuaRFFKEU+O+LxAEjOzKfg7RYtzZZQhgP90GHCd
islAY54apVmvdBOB+K5wzOq3cGCV8CAAKHyAuYVkMOVGk9ngQHHzX9J3ErsBSS8iEChw6EGpaZxV
agW/fO5eGI10c782uZSwQo2Vrs6etBj/ZuXis3N76gYroz8uzTzZroKFXiX+jDSesj4NYZudWR/W
B/P9jI4ypr4t2WnSLIaq8pdkuXfMbvgKSIXrbAJ59w0NzpQhEGE5pijgtv9qYP1hciqOIR7Z2583
ioIkRYYQy//i6Gg+LEzHl7+fzReYEVaipvfTpyr29I2EGidvEtY/CclI7Ci5gCCZhXEmyglZ0BIc
LMRe2uMAdNLxHDeeFPNsohY1KdJ91OZMK28tIsfAmkL/BXQOCClR45Sz/kxowdGdRA48M+K3GBf9
fRzZSBcXkMuYfDAiIlhZDhP+IR3QQdSJGhSPPnPdi317v5JZ5IrH5nlIG5Lo9vwl5LT6NlQVuhcB
XTes1Lhl7rtGuZDOAnL5930GskoeXitB0HR8a0FuLI8fnYdGZGrEVPvyPzQzXB7Bv9GMn7eUKXyg
fKfFEexIDQsHXEPNhePul25Am719N4uN3poh4ZxppMkNprG1eNbOppTgZYpEY0V+pxVv1fcQS55U
3CWsRUc5pwF+9LieoGUlb3n36Gj1/oA+ND6CmO8L2zStiicNu1xEMuxBIxMQJ6IMYRqhKrd7uNZF
OCzJ4xU1q3b4L7jRQy9UzXY9uJah3TergdhG/+ljH+og3uJjCFq3yF/BLF+yt+GFQC0QNVjCB6Z2
J7cgoMoXMSkauef73OLEQMbaZyiMTnoSuRb93WZ7b7BDVWhSCFv9NkDIKwWl0u+q4AIiF4n8Z5/c
XxMjBEdUJ84NhvEufI2wIKext2uHzBPz/Y7skKAA/BEPzzuOFZSXB9jT61eVXfpzsxrmCGxd4jtS
FZSMLhrIWmyo2k8HpoRacZ8eIg6iRt6eIpG3y9PB7PsVWwz/hioEJVOPM6n5/unSjkbiISXfTd6P
1NKprS/5BPDuPOCIO6HVUhwG0tVnizkWGrTDeGkZPwnQdSPCivtegG+w5N9uvRbVimc+s0aaMUJu
RIk3ztVinyDLchp25AOKirKXQEXf9KhqhZGXF/SQr2m1upn46yOYM/aWYdjz/RIFqaicJ4KZdFM4
hnOzyGSbCRbJKgnpKFSjlyt8csrIDr+gc7OSwkuhUp4FlYDxGc19w0K5fgZN8WU/wz+HMlZzL1v2
nyV+gDy9aoJ+uKorfkt6vMuCCtAu+UzGHG4Zul6LYhdANQpMfkgpHmLbYJievLOabWIm+AXs2uXz
JuyYSkfGJO5rkW/cIFgoE03twZpqoGpXCAORkOkraEo+tXwtrFbdTu4P+EYSvTw3P1KZpgZm4GWY
jwMXvHuASaYhHS33cXJs1L9s135DklNHEMhOgnKWmCLmPWbfCp6UGO0xcUfnow69V0NZazMYVXVH
iEK0tKz160Y0P6P2+wIMctwx79+bgaeJ9Nxri84CIRTraTtItkzmgqM4MsDpU0lQyHMzKU2gJRcR
VsNFTDp08j1g46IN/vgqQrbBd/9Nt1OW8c6Rul4Dgb+cWo4wVDzfPAjdqHbkpXgeWuJv5MnXR6vd
rscKM69ZogRF240Wyb/23b/i/ozZC6xnywdkOptOlVNA2ZSD6QLDdG1MLEBucujgk2xnPweoz72p
bbSubH+bery4TKzxQp0wsZb1MVmoj/gY1Ej2lwdvY6Xx3oebjAKrrUKeFgzLDTT5vB/sK0MIgOjh
WuGO2CwIi1Wt3Duuqkr/lkEUkfVFaf+GEp1yvSKNcoGUuarsdkOQlFDIt22h96/VJEh33QaqVGO7
14+qeEA/+ouAin9BdNwnQyy/jnxDdE7O5mfErqcmnloubAALFa7yeN6TZ1myBkAslU/7M0BsHkZg
yd+yJU/RFNAqIp170Dzp/+IDdSsRq1jpni9zS59Q2zGn4EAlums+uQW6Ceamo8CL57/txvBfXNqz
UPOJ9s/Q0tm3jJhhAxv6mI5323F9n/QRVjZSpPtN8G3cRI0fjNmRL6+S0+HQbX0/ofWEZ7G9aFrF
yzTB79irU8ymsb7Llf8mMHnk5xQqm2y7q7HeNUyyHlD4azHHCIXS4Vxw+CByM6ZCgrtNgWQ9mwDd
SJ4OqXDIKJ+Sd7zpapfooWYPkgILY65IPHNRcaclLzjLTX2B+ftkjfC+VB7yNrOdvAOATv5BUObp
ciw8k5CR3pO4FUByFp8E0K1P1FijzQKDs1fjBWdd8QWqFzVCmc5IK66ofUyNdzcLmhg5TChlmDHd
OeoC0stMzp0jGyu/1l8BRvSVMxosjgMimb5x2YcZNu6C72Ptc8IE4K7mgV4b8X7JocUH9hQtv8PL
p1E6Do75pC5CyxA3JVKzkyYxPTk8BYCnUhf3e3w5CNARfhHAMJX0681mpcg5LA7CNAaHkm24h90d
uLpGRcGuWZRgaON5JpEv9raMkAq+fIIUH+qE/+BFjeNSEIMMoVl2J/Jb17fUeIXELgPJuu90X0v2
RSsEug8sUX32HS7avIIAy1zE5b6OB8fcBT6+k/v67XB/BvDAomPBV5j2UI0Yq2JqKFbfkCDGiiXf
09WLGrKTpQ1kJwurOb2VMnzjSMIIhGK4ivq2xdTUyfLPCOg4FmqPweDADVk2iwU02S40zgWgt6Vj
wzCjQE6190ip3giRDt3TnklJlcbC77MPs2yShtikWdM8ihAY7Fnobwru+ExjVaT/JveFeHcFks4f
NV+n4FajM2xaDenADL2mPyyseCFFHko71TAAet8ho7dF1wJDa2fl0dg03kyUZ8veIK8AIrwDI6hC
DPpdG9uMGhAKMwJaCCn9SiQEMe6Yq57Z5TKj3d+54nX02duNwlM66YU0iWjOXGhfmZIrXpc0WnGJ
Z2ko1EUdlDlHk82TLdNhd/kGypOiBWaOYAsvTGeglfw99myhFuiJG1HgJg2ZKGGSOFZPjNV3Hq0z
9qkGD8U50HHpIr0INcV8JTvx92+i7qzrz3SuKpOucCbdveb/fnDy20hLQ0JqXYhi6MbLt0chytsm
UaJ6KU0Z2ht4fPM774xy/bPWDnCQUgM/1iFO6l7EJvhfVpQwamH5rFKfMD3Jhsg7xXzuH7DIjhGw
OEtfI4mdX84J9qkPWbmBOMn1gEjt+jynRbEhh5snAVFTtDSn9F0xXDTIILC11KxMj2Y4qymQuusw
d5FI+VonOyRwZ3u2XYHoMHjL4m5sz289dxC21qKuWGVii7HQ80DmAN97/wYFOlltbFczhcBt+GYS
a+XIe5Bvv+2epFF7I8/C1N52nARf2tMLNJjgjHYwGjBGdYr007BKEFqIFs03IeYOtndD7W8xnykE
Jklwd4+LmzoyjN4QwFb8QupLge1evoZgpFYDjpuydql4cnBMs75DlOpu3holXAnNRaIsdQz7eBT1
LkhBK3+DRnyzpP4TZWswd609fV7S/GxkFoOafOJBY/2/Lgfe4ddRPeWUuewpo8DTUvkneTccXCyH
h6BxxF93uV/y/BOBwj5iAucU4Uc1JgHqdFieSJ7Wc6mp3w/ETg9u8/8k6+67Qp+ZIQWKbHI+jgwQ
A3x17hU55Sbe/MQXZCICBv98TxDJI2X9ehFQ8MT5mcvQDnwKOCgUGNMSZ31t1LoFKigMzv9NcG6Y
e7iaTWvM7OEMHWQPlAZIVKsVKOvZBKU6W4QHUr6nsFhUFRJW3vTOCXYnc14AZRjl1yTxJkZDRbPP
mTjHOo4D0J2JX8Z6s16TGG2jYDIlyqEr7ovXxJh4uxZc+18jL4L+wXkuwmxVTQ8mbyZjlzXhCCR8
lXLuC3xcfASWkCwtwTaG3ahDdvA2BZ7/lA5J2p2BgrPxquftnoG0R/2ZeSD5cZB1x6tErnbyWU0y
tF8WPWX2n0mFgqQfBzZ9ZQX+fyxKtRuNmeBRZMXR+Hb4n23pUuPHJzbF0eHlEx/oLOdyNmZ4Kgaq
I9cyIUppOhf0cjyimCr2VCu2ZYAJ+0lRzjAssEXev4D1MWJmyR7qdczyM7L5707YyCW6huVTggCx
OzLRjt7sP4MWnyYtpCZqoA53PusCTQqSfXCzFbNp8/BGd5haBCF45lTs8VoOcfm2zOQ2m7n98kJi
WOyQzDNm4ijZC66e/dNoodcaztr8DRgMmQasyygAkZPRRDnR/PyNCqQP0oMZXBEAsetzZAmLcXaB
H7yu1vMR/dvQI0WyM9W1/zfIxTlFxZpIGa/addAWvB0sx4SPlRHPFY0Cd+7Ll5gzmgp5eTgy0cYW
ZF+WtXk1rApMxOl8SS097wT2mpSwPPqU9NrSySYrYDjrooI50UUFFOIZDE/u/b+HTN4=
`protect end_protected
