--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
K169iCFTr/K4on3tcV9fA4gcyn+I6DFJzAKxmt0l7M+VUAN79auMOIk7nhIpkD7TlMOpDBSUlvL9
6vTlMfDuKpoh7rjZngC91Hyc2sVYWS1ylnhrLiIMxontP1Y68DSmQ4+PydGQZs1NCVpK6DIaOXlE
e6ZsKKGtMwcjtSA3YOxS7c/ZvQPJ1bmLxTZUZ3JbjxZ1u951C4kixXscVY8afHPkJH4uVbBHTqnG
qIUi5p7YXWrFHaMax9flIlD8tg+XIOEFJOSQUvj793dDwCkZdf+f4tV3ONbi7TYcwojBF4jTU6Sk
bgCdS0OJpAHfRFzVwGysPheJ23s9eczY11fpUw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="roFDEGetbfcosqBUTdzneSz90+225ObRbGh/77UpFp8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
XbQ6cITZr05BX+6uMCGOD4YZJdbU91754UtxErUr+d2QZcwgyb6L7SPFuXPy6gGWKjz+W2mb8Zwc
oJNs9jsLLvAcU8cK41mz4SLIMmy4ZF3rujTPM7LcmGquwP3WOZ9ZETck7TNp6HXUtydJmrfsMJK6
Kc8+e4PTD/tTVtqZKsSkXRAikeDlBj1aBPdbtdAGhOvRoz0rArfF6N9IcQhfFWWlrnwmvKkxLrRy
h0oBhicuoIRDAU1mTsvn9UYROUUG4riXw+muCjohaITLZEckV+crSbL2O3HYuoVuCan0Dckhc8Cp
MbXE0gEA6WcxvPU/HGPqKO5VFUM8Ea1cysBwZQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="kanW/4ddSPsPL2+QP8pHJ02LRMwt2BTV+r7qx+lCmFM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10048)
`protect data_block
vLc+06OJ9NYt7MZor8Zdg52VPRQEMFKh+dghTpicQsTPfiHzF1lPRwjk2a/0bOsjMkSHXc/JEHcM
Mphc3Pv+Gbox4B9iK/ldG6tvPyDsZPh4mp6lTZBcJ2lAop5sPedtJsndqM9YwkFivdqY9wmcEzUX
pwSoaPY5H3e4aLM3iS5qXubF8JWiP35qU4Lqdhf+WJyJE/u/ekf8nD/Y0vQpRYM4H5Z8v/rA8J+y
qD08a72Yy+/7jjKRewOgMa6flCo1X2yl7xmyUdZOYoW2rVp+fUX4VFlVS2Ou29OG5f+vcaB0mY46
DKHt+YzH5vxXcV4xH9BHdsgTQ6APgfw2amf4ZPmDhz0qia7tHZW9zAWZsupG3uUYB8xOn02uT3AG
aWjx7EiRpG26bnaMrXxMiFJPGt2ckHYvEqN7t+Q2niHnQvELQ6nGoeJxW8AugE4JNLr2S9hv5Xph
MqU1WW9q7/7mvyP0a7jPqcb2nf5M/ko+GwVgEgsdNg0gLgQDrdpp7p2KF9S7Si1DnCw+s5QUkTD2
IFheaa5RQfnZ8wIn54RG6TEGg80x/UXbx/qCx91wsMyuGdtnTIBXyfywa2yLRznLja2Blov5PHim
AmNtPgJbphJtCaiSM9gi9unHRuqrl5ZUNPualoGO+Q9EGz1r9WcpYM3xNpXxrycvl3svUAj5kSKT
gbrAY54XO//jDnAYtc64s2ROo2jO6YiMVV6YomI7aexhm2UrGMAcFacEgCyzzHilDF3jU9joGPlu
K7i1cHzHh/qyjJlUnhjSrGIdSqdfbtjeGmP4SQr0uJSisYLnaglzUtVe1LMX4SmSaJ7xWcRxMddz
jI0C8rW23sfikGYnV+q7pZdsr72zVKukA67ntKeG5vACQR5+6tO8qLGlLCywm/96IK7T2CLRFysj
Ej4FYG5GyN+NT9/Uv/LeGQVSu1yiwGxQSGC3PpS0jbkkqMS5ouIc6FjZlGDjDEqWKAXk9V2slFLQ
6BoRPYRHkFBmIbn0WaA8NXb3El9PvpRgLbnyB7uM6vgcYj/fM81blgWoU6EveZeex3x1wz17hOSE
JJzmN63MoLTCbTQle+AcdBo6kcB2OQuTuTpsgXuzhON95o07gb6pby76Wk3RkB2iwQ83oqyt5B5M
v+O8VpOIUJI06S13N50ZCwfbGQSf/1bWCX0dJIFMtsFmOu/Lmfo2AVX398Onebn19sNRAazqECQF
48e03AcojqlryWIrPLcz8A3HUqrPavmdeI2eZujoh69nXl7nHLei+9ogPIqc8JPSvFHjO9svA7NP
uOOy/0yda+xBGBQdjzzERB0PSRGzjH9aC3BACT8HtBIoVs9Mnry8LEW+/SdMpRa4zAyl+srn+ZUM
01EbI5ixXWSg1mGdbRcu1rd/fwIyZGcADoKnbWfhHZL1c9ww5VNQtXGApXEDkkIrVWBEKaB5abEt
YYS6SnHXkV4JLkEnOUgAZDQhE2XWg3rqHeDHlFZFue9PnKLS+RoV9UK7Vb0duLMuLZBRVGGyuwcI
9Uc5COmecP7K7adlAtF9RtgFjS28YTB5zDy3BZvrQr7JmJ1hNCXaAGp5Bk2qnfJCU1A3SFr+X3kR
TXszs2gg8SqYSJu+mODQbGXCerLcAJBlmvEoblTDen3mSavXY1GMsCxsfr3ZnPsXbxftrrkPyNbL
U7SFqEAeZkiy7scsxCbUskRDd5HqZnStpYHQvqTpd6D8WvRISBJVZfcw83gV1Vur7Deqnv8wTqqT
RnDPzY4YbyoTk28OHLZTev2BZ4yRuSv97GAwBvGyDFPjpr3hwMhIqvXGF6lg8ngdCf4owAObBKsR
bHkIQ8dMBHO3EahehElRu/qLYZcnKGdX76Z82RolFO5pfi1zQZH4tZIEtSUrO/s2ZBimC520mAXi
lKgOFRRbPzXpf10pA0PEX/UroXSVQU2pwlgQaH1o8hlCNv8KaIChGYE+GKaliXGIEdZ6f0y+otoj
6q8W85jq2Xf/TfHZDbmepnqqnj8WdlTz2+QPG0EDvY67Mal2ZScXI0K+KVXViVP7gFiL3M/m2qtu
z/5GF8QBBAfEgzOtd2dvyVCRshXiMK8eD7N4Zt1hmQlUHbG6c17OHZaztjtfyiXAuTkNTKbSGfQ7
pf0tJLCUoZGpFrS+XflKJMOI1f1oaGUmnwivPyrOTc3L/vx3LscxylK0makRjxHuLgknE4J3Ttzd
M6cuXnekvqMN+vWrC2OmwagYVTRvf6X1u1N3FOzsE4hODiwZbAnD3CrbfYUEkyqSBG23HMevOiJJ
f/XDFUoRoBrz5ijysuFIlSIuKR6VLh0WGUFJhjrL9mCIMDXrmIwmLLOqXzhA7DMPRnza1Ypiw3Zp
o44rtVrwgw0OgNuH/jsOHfTsIX4Rv0eKHtDA0K4QOtdWPWwU8KlndGx2KuoDT0EqX2nVMSXnQx2R
wjZkkZelIz9IJ5esGzZSdq5lITHWtzUqHd7wKw+c0rr/OOHM+uYpb7YFpkWjxZHzwrWARprvrvse
7ywG7xm2tPzOjM/FIys/0x3AIpMwWPXVlXVByZwf3RcbXr4OvwyzouC0iCXWp1uoOLi0gsib9bWN
UdPuu6GGiZzq0ssiiYyU87BRWQwq3a4FByFE8NS5cqJLnCk4dnpJrb/uddAVDNR8p9MEo71ORscI
ZfNZq28wymzr3YS91Xjma30oDOLEgQEUfjydJCCWb6NkJLbnJrff51WPJWX70prFbh5wsoNkeeFG
CGB9ke1WSXjOzUxU9z3VvyVtLXOr+cHNBJc9uiMCLma30dsOcdr8X7gquCfQe8AMGKx8wI9HK1Xw
5Q48XM/Os0iW8xT1vE2ntj+yXjtQHnvU3UBr4a9oLR+uy07QLOmQAGhvctZ1TplIzML+BUGbSwy2
wXVbUsOWzvel+CvuUd692Vvlq7IjKhDESIQatbL0S3Sq777TNnrt/+5T0BzULWVJiLKCW4kyXnp5
JjGSrSBhG1ecc+qGzYHy0Kxcy2m71Xp/N/42vQo3pSU/zsz8EITmp12X6AU2FE/tPx46+feMZ0gV
tH5rgx1Khl+f3yZR1Mz+ZrxF3VLBta5Ql3m+ep9ENjPkFQMRN77G+Z2EnTK8TcGh6e9PP1onIF/d
E4x0Mq0O/H8X5z4CK3GFKoMhrgsb7O2FDO0jMcZa2IobEa9V4Sffybafo/K6z43uVWLnXtuTuTPN
RZVG0vmYv/XM9z3IFBPEHU9nqHpvgoe9pyu6sp3JzjXW2SJ6lcmz93wOXg/n41lTXekUOpMgyPir
DAw7q0I9wbIWdmddAqvncBiJ3H5yJ0QkcHPdZtPq6PnyrX5nDrvfSKSSMJ0YxgofE3TlRFzVIQQU
Rhi5CzhxHTSC4YGvkExUkgBcpc6bpIo+lfnby3/FhN4c767+m0Zp1oWEHyuN2yvwvh2B2hbFuV9X
BH79H1gzNJ6rRwzdypStgN24MpQR7Yxunn2td3EVis2AQQIKIiRkfw0zNhiNn6DZYYJJQVFPX+p1
RTehVuuLONhsvNj2fo75D/wAH//1cvBB6sy0JF55szp7JQUMJb+Kdn7STyhJj+qy+x+qQbOksPj7
hFZR0lctnbNKW0eib/EK/9a3ETu6X51TV49qwghV0t7zl60MhSKCkgVqOEq6wPuxKyFh7dwmMrmI
kDKoDR9Qhg3g/u/MyuO6suK0laUZcXcn05kaIrII4BT9rkEH6WFPXjWO9qfj7EjE4VxoRG4rtAAw
Z8DaDO+mTbC+l71ypVqqjRJJRKEFqSsnaASQsRocCwZ3usQD7vVnd4QOEFAhRXTHb6e9deXq+mha
o/D7rMPX3cL1OAF2kt8FH5OeDVNxIb3GvSzhrelva7IvQe2dH0tigzdDGMvaXADwXMLtSpgtjPn/
B/SwQo6W9tgCz2wL7v4VaV4IuVTdVrgEn0XSbAON6mQwtPAQqz/WiiO9ip06c64FzFeFkshPMH3L
HKreF1fmYAtUkvNqL+TIkpJhxa1V9fNUqxqXoDWSMg/9tnTnNOjfkrOYYd816L8ysEWXX+rnsVB6
UbcRPg/eLAUPQMinBJ9RVTUUSsDOPK+gP9nGZoTGmTxbxYhFGfesay5jrDenXBonnn/EUmyIoJk8
EcKKve7yw3/rE9KEseKB0WLjimZFLK86us9azagUeTabm7jv6hHP+BJU7qQZC8fnmYO7z+WgGhv2
lXu7uJVg1dDR+pZwhriatelkYE5M+vK6g+y8b7XkquBG+t8oFGYtXFRD8FMooGvJ2H56zYaIj9Z0
Uhr7eL7lP3ZKGrZaQKajH670gV1WVmk6niIzY7B5kKa/sV9ujoiJDeoARXn2aHegzd7cP1/Dbbc7
zqLFQXOFPjsOuEufXi46UqyLHyDHfk/zpMFtXHXTVRhjXblG/Sle3abtm+saChSN89X5RVRCfegJ
HVWCgD5qiuLLta6BlOqJge/0yTM1YP6JnDwstrJCpnNO1lXRanMLNxO/igaLQiR4huUtbqs8aXM0
iNjOSl4uEl0uwq9qYETFpZ6nwE5fVpXaTG2wTzmkUkHnPPOACLoydb9d5wTp5Dp7lZ284jMPPiQe
+aiepDljczOjcrJo6UCnECJaYK0mA+9nCBuGMLTj/EkxndTm30i7UfSRtb7Ty1hCWA0aYERANZHR
h6lPOzwG+sq1rcOkMkrGsj/I6AOjqGD9AR/5BqFXZN3yaY2gjeoXCq7fy50Yt45VATKSKVhgfv1f
Fv2BVvErm0D4XMHSgz+hPuU71XO4OqyVs7owMcdU+7Qop8rLLtS7BAxNimRasfTYz20L6Xp9kiZB
GpU1ahjBI5qa/Jlvuaf2aTS2EZi+/Cxr+WAbs+yUGjIiatARZgM45mFhy8/AX95p4xxbsUZ5pJPC
lM0oxgK607j0Mox+K3oBlJiDyYQjjKDrMEHVbca9h2MBvAmZ02d706EmngIJTgG9UvicG16SyfN3
0kfbn/yCTmz84gLUO0fU2m4kcChmpy3x/O9hMUwAGsUzAh5QE9nhL5B2sfoWcWCwSz22mtFLqxDm
mq4/04crmhLpvPGF5O0uWbiMRHTDFUxCYzAXuyYO8Un1W+KWDwrkNj8L2cBAeUbohdUr3fEnHME7
nb3ee/rPWuc/BY7OEUhBRk8RoSYH+OHKROPjNgYRNKjghk6azyFF8W70wBK94tiob5FkqTHKMKkG
CXzjFYuhLueqKZNH4A40pg+ECSrkl8YAehB7vUJyZM1MsH629rV9If4D2cyDICNH8uvayGCRZIWE
s7pYGcNnBhW8AgXfAR4IJWWIXsJJHQqHVC8oeui88FpuVTdpj186qJxvYrwHSfTbTs51AKUKDwc5
orTZFTJ+o2LWZVoCNHKAfJXdxYMf7ReAcu0oKwUd1hxXroxzkyKydSgN130CAmGE4o+gEapKZQbd
lS+ifF6/lN85iZhzDQlDx1u97s6yXVmbl6NrlV0gzHO188UY+tNDYZx+rhJtkMyo99Sn2v2Kk0os
KIgpNyozdZPmZtZmHk5bA6Wffov3TYi+EF3pyjswxg/xP3yWfdVD9nFQ1uQlh8ecIsMeEaF2YniU
nqD74KOzdX4NfCaw785tQuhn+GFSsGDbl4yBFS5ucjLyg96gQ7EQSu6JUYZXw7BQlvu3b4aY8i9e
TOrfv5FFvhkO80sOoSrgRJi3mlEZVN73dEfjVrwK/+JQ5wfC3wjh4467lmQEJA/UiPxAQkHYEPYN
A3YBAUpX0iz5YuRoR29YEx5K8NxT6MzEvGZr12XFmEb7w10hfgn28slbREvFSYun/ewgm34NkBdm
azTGZFr7Q40VJ5iLMLqbe3uw6+Z4OlQvCPirzHE/dMgUVnYOKNlx/T+WsxLWs9PiL5RXe2epOosk
LZj8gigIpOoZW2O2x0EX0Rm88bZTkhOXPG76wsAfZIWIdH0R4U7ZZMxh1OComQOt5XU5vA5MHFt0
AsjvACSZ221g9LVISyKW8owGhciepLBg7DXN//WamBAFZY7iLInlh3dnvGFra11wXRz+RnV6Oqgo
xU0/yexERcKEApLgdWeR1TU4w8zht7rAZDLhvxr3dv/PEwIyi23+IKoMi5lxtjfplnpmL/YDJntN
euoclYzL76yPXEeSa2I2I/B5X5DiH5zmuT38cFPBJbxXG/c7t1ixZu70TjzXov8uSSBe8hWtnHlW
uCy80Oor69n8kX0cTV8VcgXw3yya1ZbvE4U+5thR2/nFUv61QuBtNnkFxHhKX2fUDmhOmXK25ny0
sS7ycnYOv1Pcx2n9j5JYFvjUULQMi8DT46jC1CkZxfsoIZ2Y+nnVBXnwZDqv9bVIPZkcZyRBhr7D
0oMZ8JV3H1sFjFxL68WVg8bWcN1Ee38H9gQaVhJm2cPGozQazUXZ+VsGJPs2wmOtpXlgIvQvCdiJ
UjordUIiVE9y3FOEO2xRpBdCmKvmfgTrI3GKdP/wopq50TGjtB3ESxgig0q5rG99dgdRYG/OmVvJ
TuUx3M80oRBIcLg21/8dX9NO1U8vSihW5VEBfcglOiWa1KD7jxc4m3Dbq7kDqa5nopG/Esx9shMQ
jSaFm8baqEaXnRlBJqhdTZv2Pp2MZuVLcQAdu6G+7qC1ysrDpVL6brR67pv0PSX83GhKmxhvYYm/
1DV/VAdpRPuGIY94lJTgC6QeeyZLAhONzWFfoDIqI/l70z4Ut+nKv2J1YOOumxBRs9L/EsZUCcNC
VV9YU/aOxvvo8qG4ziQ6rUzSuu8bnlF+yDHKM+TnhtcBZJFKTFv3QtU1gXkN5DfalXQOChtWBeXW
1M+GG9/tMz+brXnNB2CJ3ObXfG/IluCSOVC5ah/WwfITHJN55PmIJatKEKJrpzKbtwkTrRIkCvga
EOpg7OWAWfElfJ9FsTzNdUF3AZp9q4a3qoWbZt4qZpz4de+a6vaCwSgysT9N8Hk3KCWQpb102wiC
NB4Nnn+8qumpM8Wvl96mbmnOWVSWqrBpfeE14VvL8vmvrUQFtAn6AdkLpqG7Qqrr7j3WSxbrmu5V
3ifW6FhPPj2ULPm2dapRHUydlOQ+TrVqR5IOi30siUaeqdKC8ed0RT60Wtzpj7dLBqmtIX47c4uE
2jtkVw9GqosNHT1dnvK4Rs7rdXvUaFYtDCZu2xb7U6lNYFyDrjsnjvulbA4gEtagaToimyDyX/Yf
Pd85KD0KnONLUSBPPlu7aBJsfJ1g9FsiK9LIkpeWfaRQjAXW37oOHPiDyV76eZzpuBN6f4yLfMwy
Hd4ilNvzs7qOjSlDiGcIo8Niwh5HwAuekWs18v4t2VO3FCyPtJruWPE4bn0tUctsSDsF8c8iND97
7FhEUGolpLcTPMKY3wj5zbD4GkfJE2nz+ZU3eiNqXsuayNl9r1qIwu49iCqqf+40xPuhzY2O2fwD
ioaJcQcfWn2iCvBcGxSuaKNGaUfaULFUnr+q7Z+mny8t4pdIg6BHXD+QQWTgA7MS9x3QYJt2JExD
wrs2YlLnFEoxxp+r1E0Zj8rAatXUUpDfDQq//v4C97PUU+y3jlpBLBhPpN4OhF5DZa8EySxoLyCH
KcU2yyavGGeLFS+g565fY8iAmNpy/m4OcEIku8A4TwKnymIs9Nv4qy0UCyyUor49HpfhkSRv/qRR
XnmuQyHQrcUGNLtHeXUMT7o6EBUCCCz79sGB9XNbsJfEsPkXbMjyBqsXqO2pgJnSmoucuN9pAeJP
c7Q/KZalhY+vqGOSkSbR9lmVvmBTfq2UP3ZNTEb0z8wCD9glzVKLdfeiFyR7erJ4HE4YnV77a1yG
wNytDG/fY4Yo/ihn3qSl0+NMa/FBksCVExNhyhJX7syGMGn6InyvtdBoyqJVabs6j3Nt+dJDgi4h
fkkIE/Key2LiFjRYmStMR3WzLidx3h9DL7Mls5Cm5JxrQEoX7PErDxoIxApW8DiSVTGIzX7TVfb1
0GC3EdhsSwqopEgqovOKClDqp8RagT3AsV3EizkF04bGjHMripGnLjTgLBU4wsAEXGgencVXUGzW
t5np/oPPLR1dYs26cG1xTFiMpz3MpU8SUChJMakq2640zu4lX8EeZ+80sUlXaBXf0mBM29Br6i4y
rP8tKzOAzeF9tw9Dhn3ax5vHuxOEH2L91xEdBgAcPXY3c7dxjvjSYP2ym0NDfsPiV0+jBeVBqIPC
AlLdJVfKd3zFFvtvF8shLPD8tMHk7N54zr+Nsf6XlrwwpLxa3UQxEQxBcDrciuOcaPKNPhun6MKo
h7Kjci7bxguxNvd38D+oWBxQpMW0GoIVI/xItSyNxeABYIOlJiivHKDjj5OAU55kmIaWgXRdZFMx
SvKx4VnxFZz/gS18Nw3ZFH72ub42XON3X3MwkG6k3gtDaKNJgCOvJOPyF+q2DA1OIy0pzSZlxNhn
aOmMAhfkLo5jcjPz41m7mMmDPc++f9f7xscQQxbzZynPP0aCwyNaVR96bC3TE4tFF7AwzzxsBgDj
WNKtwAg3h7t003zBeIjRrBJk/T6VUZLqVX1iZk+/Baz1M04tX08hqdotkoxoT1UcnaG5bsRWbi82
VAjGEAEbSIwOdfXVmKw6jAUou4zpkvDnhVbESKWJydV02knRFn3D+3NnwP148uHudspxsfMUNKge
tp8dagvdikhrA/Fo08O9CQfAj4d11N2HXIf9Eb3z4Uze2bXVoeBF+Dzw2g26F6nhnpFSyk/lsTF0
PqyVkDnlgPLPJt/od9CHqjSqaLfdmKWMYGQbDnJfjSi4fSy87pW2ELAgrC06Wjrl9YO4y6rC+8lM
sZkSZWURyWwhNx8qpyNTIZHZaPxr0A9Ly+NIkgSnXOgQARTO9vaFIzh6VZyiVWP8bSyNpAvYLFNs
srXYz0jwH6n0YgwA/9a8DD9zDpZRdS0ABIuxVKQMAFOX+3/AQsXk7wdE4mqCnQo/Cefuxx1GANiZ
knmwigKPqnjxHK04Dt45FGW1TL9ZwOIHjQlBKjgvc69GYWDft66sKpDwFXOZazbVzT6t9xnXeB+z
3wuIrYit/woYP0ieaL3J/SRWg/dX2bI+NIhlpDW1XwR0JvBM1h/ZWn7ks2RSheRZ+gAFg+Go0tnx
GbTLqhDcfx5+63Ip4B9t6ni5JS/PNG+kyOx//9wAE2oGxcWnE8YnvIAuYIXDQnlgoJOAi6JX+BRZ
cxO4gtCe9OXa4Y5yYsWmhYO98zM3BWEzg4XPk3bR3BoMgM7kRuhgDE2NNIVz02+fQfewiedcxz4b
ihPRnd7I44LMI24RKOhVhSFuYFy5QnGNrH4MkIQ3j+2HnPwRf6xCNfFgLh/uFQq2N9ayJJ4Kys+N
DMN514hNIRPUoulMDrwRQ2OhLDViy/LY/Ul3Z2XISbGUfXhiYymVx2Lu3J6X1hMCwxHkv5v8gy/t
tnkz+qO+12QfYc6injze1QyaXgV1tawBEZOVaibuM2kdTa9lE7UZ/ZX+bnNApeL38CIZHOyjdOmL
rNwP4tDRZ4jjY4MuchyXgbTbHZ4Jf1xxsBsbiEzK/0grvhTUdZSGxAfYdb45c8fqHFLoFSGD6zfl
Y6na3PBs6zpX5mL+Mz1zJZAAMkdSmoCJ45W9icYRoj1hnOdpYNgwKXsfaw4nzB7T0B7M7M92lNby
xm9HUXgj9yUjR2mGpdd54Xkz1J7or4M7mOjblibYrj4DsN+GitYEb4JlWSev2YpyTC8mNIqfasQp
ehP/EF3qosHdri0fXZJKHbh4M4ARZ29eDnvDVpuzJASCAAbm3rFrLFFbeT5lrB94TZRBBCYyDfux
Rq7cfRGaCxRu/eTj88r2gEbpF20iyp9qqn0ewj+ZjxQJeXuPZ/ADyjF0sFYzWfUraMDyZdjyBK6T
FSilC0c7ZdKbWBxpPT15xeMujetq34Dt9ik/Hv6IWZkymD1oXnoQlh0dM4BQNqExBF7vkqYZ+4Cj
hf0D/UUMn6yfO/7KNLySSs0xzR5M0KFAqwhQ20O198knysEX0A/J6j5v8ydYv5lzY3BZ2IYkf4tC
DzQjNjhsauhWrsv4kGf0Lot9bfHMaeSyJJ19yFnWtEt3C5RxCv3AKWmHZxEmLTyZmCssEkslt2Pw
BCbRw+oPt2oG73hS46NWWk51xfcH5rkSNbRF5dV876KAHxAU2zU3ZG0xJ0xUXqLF9FLVlM3Oc/Lm
qaMT04r7mvDGNVJXut84zjOMHaKt7nWN8Z1IjnnUARQfCFdOp0l1wgED8w/UZvoLXLiJaHX04Yk/
F/S+4dJBGObUvM7VDhswnFgCDniAsz7/VYZXr7LRQ+Iju8ZYdE+FDbitcTs5xnDfG4iIpxLjkA3K
iOhio2M37ugjR841x5S2aO2Foy0NzP9sdw0EfL5bsrodeL87jl1K4X3rJNAnhKt4PicjWsLzq+9t
fc5M/HNtB3TdzvyGTApzRHNNlmeJSMcg5+jEeiHCf1LaWg3HBH9PTOLzbGJKlDohlfm7ZpaTQMSs
9jojfKNJ+51AYR9Q32gG4pGnCKJU/LDTT2jkkeoa02wwYsGSnus9vkuQrtzRPnncQsJAkvCVnHlT
b3SfC+ul3V+wGdN0q1hkbz1v355jpJXVrJmFKXlPuDrCx8eeHmTEwg7W7a4zZ1qWeWdnfq7pYlhl
crpOiS+t4enbC7xVrjBB4VP3s1taWzNGqIPE47Y4NdHU2p/2jn+Rtlvsx8JBPOSk4mqAAETaaEze
YGUAcDCgVpGJ7yG4ZH93tXp9j0krKZ56lWxnssrsCX2ofg7fOuaNEr9dL8QeXCMptcos/wRmtFCs
7iUxED2wmgTh1k/B1iHtrC82kuAH2eaKdptxnoc+jF+U91gweZLZwIebHEyMmv2tn4bwJA8EI4sn
EdwRZCKDKEGVeuwIBMiMf3yvKqJ5C/z+HnKZRTIyGPyJuGtudj1b4vPaJsNpgu4Rv17saPJsDvqY
TLFqPPdN5hD6Za2pOu0wXtvQIiHsUJ26WC9EPm9Y+ARLIOc7XQblA6k8DNInHA5aav5t8Kngggsc
emOqPl7EK3j4tJl5a8/+6Ohi7RkN+mcRDlCQ0pM+i7s9xF9QSfECeVl3fMjnxIn99DFmGgYmxqrj
qOfBW9vOsmiol2fYtp3bLBnkPhD8XjTSdMpxcT1KVaZ693g+enTO/RZx5EZVQpTY69Q0qkVXeEfO
WkNPnP5WnScNC5qlEg+J3+Z/ChZfSw4r8XML26AAwZW1jblaggBMfEWl194cYvKe6nqVnX6Vrl4s
hrtFI82ClFh/R7y1yU586ANTKWn6WF/y7xYRhlGpD713s7vUDCYMzdnSwjsOLD0evz2kjMRN0JMp
6I9DPTwOa5f6Z0WXDoyVWcVi86w2chIsaqX/QIwvp82pPxjsQJEdY6Hdzx7Lk0bUF+LOyZOuRc1b
HDg2barzQy+pb1zk8EmNVIID2MR9YvFy2dMf0C3OxaxcvofIun1zXlspnWUCIBMtUG/diHthZERo
ReILYUxPB4TUreRhxxt0CfxBbWQy3RaiZzZpWJkjHVgKzCnfhJVyMC+qdNnDFBbhQFspSo/vvWwz
TwGOCi9gPwrwiHT7zujg7qJ3oqItt5RUwEtsOT4p9M14NouvRUzn6RH1WvBPPVSro/sDZCWFj9fg
fZwtLPqZatgLGv3EcxiNMWTneQ0x53g8ZMcgftBGoJg1nYxs7xY9NK9vtD25H/bCartbQ6JIRlo3
jzxVWqCpHC17Abe3xSOnGV91e9PBXCz2hVedf6NXSnQDX8k+HHAnaJHmrXSEqfhFgkPEA6DdDuOe
BvDUiQES6t9zpCkQwNgQxnQzQM783et++dPjjTd5lYCXf3F72FlFcbchEwYHMcSepqeYK15NmHh0
rwpZW//tyOuljSFAPahG5HmMwchWN8I+0fFg7DLg6xzGWdlLtbI+lbbAW0tHFWj2EPfenGbZ/FRA
Ilg+bRoUCrLF32AKiulqPx98AFEBXiN+L530yf6XHG77bTO1o+6CZ/cmIOv1YXZSi4MmrHpkQ0ok
duP09EZTJ7JznWdsdGP4GlOgoc6DVum4pEmA6rSEKeEdIjUSDEnvq/5s5xzWuAFXI3n8eRES7Bry
W3dq/E2+mwfJu22bkjSgTUkMzmp25d6+0gE/LZdI1tu3VgVm0+nRmQjTVoCw7kGEuQTzJhHSOSC3
kSI9TEIyYqvD/1ihOmcjhAHVTOmo87ipO/jRw/RoRwMJJPQapTVEhkQcfi6zI+WLPpS8IsKLCBRm
E/mBopX5yE8kKGVFJ3xIHiG2iUCSJeX6b+csq/ZqLnBqflKr58kaJxydb8wI+YGIz8T0efFlyixs
PPQf92O7iqjz3Msd7TY5L4lWe51XIOMcJCaRbI5lJMhltSPOWYIVmHx70xsj/sqQatfgamllMImj
JoltYGB5YDBwqt7wWn7iO3Fegj9m9jEFKPwwywqSm85kHvMtVbHh0Rab3jYfUN+oyS0P3YeHNuZb
YFYvvm+UmhirZ3bQFscq0O9O9mN2TD6O9ZZt1ZL6/o2lG180eINK0Z7A6DWla43YTfpBgOuE3mWc
q/VKpSVotdLL+z7A5TDTKVIxEMkTm6JaqaMbNU9VWCdLtyPJ44/LYI4j7eqT/jorvmfyfD0EXqc7
b5RHrdLqTqjN99PIgQfaDwbKU/3i7drFPZrOpIKwk1vO+ZSctFFfhcxOERV/gDx6+YTGajOTd2La
EmxKzgEBUJafDFBdU6pcJP+Ml3Spt9Q2ETvodw8ZAPO1cD22vsqwjjrqQbEoSZfCFMCUUqzmLWgH
lskabp8wssxW0h/9iN3BhtkB5DB9Me32BUU317JGVLzoT5r9hu4ekTkYsdAilfPg9TUXT8fz15r3
tOOXgpRJgj871EyxqqOk2guKJJbSZhf8ZHIqxQWYhpxCpy9Lpye5ct0rECXAdg0ugsTz/SN49KjO
o01um+YkiTAYdmWPTRECj1vw+Wcb5WcPyGDuTUyMLeRaPywR5BY3oX+7/Gqh9O38iukw2LLHRKcT
WIbEwuNWB0jq3vOTP9e6qqDxPwQSDr4aHjqF1tBa4IFXGGRha0IEHSJMojKDXHeIlH6gTMN0YWAm
i70aK0VvTJtOyd2cJJH7RK9adj7smxrbQxs5tmgYVjk70zuCMiE9+mJUUy0W9osR4wy4VzAlOsnP
laABVK+5R3474K3l7UESY/6iA25qP7rI3zP/FpX3Toxcq/79cc8HLyygHvJFm/Fzw3D+rWXYywlk
MgQwYxAh9OKBc66MTKvtiBuT/Ri+XnGFlDWvgcDOisyk7rSquCSKw/yufy8uFpwiknDTmgmKkD6A
AUj7nDUktIbcyULlF/qGkPK9+1LoKbFP8VK3lrIH21w7YzTGQMJ/oItZPWxhs+7pPjNGwApY/LyF
BWP21T8SYdfaMlYmmUEW0s9+auXSZm3BKg4NY5wkMmSpNAGj5CfSQlsjamRDYY39nqoWAs/tAXel
+kKjNFzaGY5RzYiD6x4pow==
`protect end_protected
