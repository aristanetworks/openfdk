--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
HulN912qd/N4BoH5CH43Vq2zgGYJfB4Mue3O9WpygYNgtZwNQqQxHxti/vibGbur36Ckb9Wp8XXy
bdnAnBe1QeWDliAcWVWana8IDMyoY3gh5XxfRKex7t4ubj0r2laKeljCW612QYBQWeWiXva7NQzM
haQsXQ5zU//uzl92hnaR8wdyESOIV57NLluI6RZLvASxby9D+yaKSev7x9YCtuH06Vhtzs0xae8o
mdLIBKTYhWJQTcSjy9S8jQFOe9CW8xgW3VblRJmwgFUkFW4mUxhMWKZwY7E0sYFFsjBSWuLgqUGk
RKXU4ucjpEHJuAdJ8T3fbO56Akbfn3NJ/m1KfA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="17Ql6okz6CC8/C6GImltfKRudUM46JDasOZkW1nwtWQ="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
f50CKeDdu4/ap6Uurmc5QNcgUhZlk9SaKxinNcGCoWL0kEctKEZKpcnOJYKMwQEcHufr6sqB1Q8Q
P5P5ir9Fyx2AH+3sgWReoDfXyeo+6yO1I0F/jcTnF1VWtgSQwkbGQ+Vh01OR0DKevi0cPFKFYwTa
4Z7mphUvoyMfkVkvMelqtDyxQj3XXiFUb7Le4oz38k0EOjSdXX5y9e6GAtFTQr75QpGgYk8TaKxw
RkkfEUVkZCmnNp3GJDRc6aVSBEyzL+Al9tCzY0LxVz7ASSVifzeBLh64lQCtrtuWlF/GJfcRPxM3
Jy0jy/c6yqk6mmH5VGsmkOuaJxsNwOoJL/Mpiw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Fpt0ttWz9NYKDKIEEqq08gqYjIsNn6baL/vE2ApLB7I="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13888)
`protect data_block
mVhhyk5NC1CIw3O07NW+wCJb86XEPn9PxS0FAUPHqieZtsalzkpWZPGw+v5ojcE0RG38TgBVtkDj
p+t9ocTzgcuanhZG/Z2cztAyS2IlTwHSgHYUXTi9sKkWOe4lfwA2cfVCPWfKSjlMi31Kdw89yBEm
0f5fKM4NwedlBlOit+ffkTsJfh1gsPVCyK4ixJYTw1FxNGak1VrJMlhPBsOFGssgasy17yzvmdcR
3TxAjRseW5GW76RJZCTAhAVkpomhdSWd8bs7SH86FbUHrAhG3E+cwr1OqdDhliEA/U/Wz4GbT1pU
UOL4XOYSB3sqfgVf+809woT0HFKdNZ41iRlJODjveBmcPgwrxVj3KBAL/S113MkR1gGxalsQWiFz
PSYffj3EEkfdUFC16Q3EKhXiU5YMmjXbmkW/z82YLw4Um9HJkfp004G214Ul6Cf8LlgZfimstY0m
IFEeU6mPgzloXffdBiYSWKDSrQpriAlR7Q39DMX8Fh0ShIVzvuzWfN79Qak/pJvEjOUhcyOsEcV7
D5JV1RaAeiJ6BOdLeyr5AvhoV2JwiCoQ1oBIgVkL3XAVF0c3islbyOwPuwCioNO/u0+vtqTb8Qs8
sBLDxnj9Q8KEao44r7YN1DhkMvEfJeTxiVgRzepOhuk5g2yxbyjpw1gp0Mut+m40DiHAL5rgMhUp
NQu4NWTiNC6MX3lRW5S+GqtazbDceZ/xvkr/i/9TznUZcpevgLwEG654uz4BK5AlPYi6etX4GMeh
pxFptGBhUZladiOhCV5OppxAzXsm+4DCUtj0jdYEuR1AmAAvZGUWonX0eLGRgZ8GMPS8f1jpLTL3
C0iGzXg9vdYOQQ47QAoaghoTvqNe0+WoVjsjare9yP1ngNhOWzdyfX06kIVeehGDvTD7xwEfaH8K
8JTUe3dYFJU659zBAopNLUAA8mJtXMDh9/TBGHnMHAE47c2T+o0ap64OCPoKkN4wFKNubX7R2nzc
BXzx+aJT49UiHJ6z3huXXE7TOijlRQloMqrblLyMlUJe52HjeQl7TNt32f1ZyKjWAA1AoU4lCKK0
fHK0FsKz2lxLyQ5L9DFtnvDc3oii/DN0G402aSlWNUu63fMYa9kkznq8+uxpGIhDOOOIHFvr3HPj
xagdjfcaMETOJSfEoZOHNlokmvOR6j34bWYtDRUhq9Kw4DY9BqSKX/txcbXSLopaVvsdZl+pzmAG
Mxt60PBz/BgUjrWAo9YMPY7YWyy5N2cLaRj58tyNBn4X2XDaUQIe5S/ujLTDC/YJg4yV3896Jgu0
6oi2lKhTD9tS2NtWdJmq4H4GjTFB0SJ+MqfKz5IHHtQiupisSRT6xxtZdWEHtyTrO1arQSS5kCKk
K/yNUQCgje62I+rUklCfYouAmZupPs+dAy0zhRvyxCc6V3MOwivWBZQY8SMFVv00nrzP3sSoIKeI
eUEq2y7E4PgvmHo60yFSIsmnVjB5/dUqkUf2Gt3Lt9zyU7gWiM8ivXXz65TedMw4uTBREX2siEcx
qXf58k8TIf0NQF2Duk8VjvyYhSE0nMSXuGrF6mim9q3JiR2JSz1xOZ/HmZX8Z7IU7D1ME06WQ018
u+nH/idxYmlWCIkL8Jh0NvYrhnZRlqakWkLEglnMfdajzGSlU3MjGSSeUAaGOR4zdgv8oNVWxKqO
X6+dCm/mavpj6eLcSaAOxfZx2CY0jEM+9pmbr5SJSLzZuhcWmOsb99sywzmjvgegFD9omS0n6Icg
ABM5eIGodnW3a98t7ZscfQ19k7RHwKtjN6oHUyVynIhg/F825sQbIQu8h8isFHEfjZcIpA9YYYSb
26id45/SmIBp6D1pmsESMzUTWHygIeWV0JTOWh6wTQwcfFgLGvkeVUS3lyb4qTaekROATZNog7zG
zl/QSSxsp0E0A2pg+aMUrJLps1GXeeK4OpGDJ65LSg6z2y3nSqGjKio7T6BTEabytZtTZNK50CxG
TkMeYq1VIeH+aCabb26Tv06pl3dMJu4kwRuntZMK55VkycSfNvEwV8jNwXHSFLT62X41zooyKt9l
bf6I6mbymeQnnPSljYqzpSKFlQVEz8pCqE4MqP2Np5pgRDVpqchWkgF9Gtzxe/7tyXVolhd+kJag
CQieOjQWFJrSX4avIN3gOJ1g5sTqdMfICIEvp/U7wNXLSSb9Jat0IuhbrdSYgzTjtcnlI2rrpWfo
bBKwWieH7BCQR79y8hih0Zhv34vbT2II35tlMISGAr6MGzdKyAb9Ii4b5QZ0ohOffks1dWD1cVEM
iC14TGnDKrqcy7ddBl+o7sdIicbvAnjVPcX/lxKWxmvoLLBY8hr63R9gQ6gPAmPK2yZus+FlKps+
eYhJ3TC9RzE9k5MR77ERLjtS9bp+TDvt0eEQJ1ts5IgW+tqJja/sxiFrEjykUwAtCc4B8UbEZESN
hHoObtsZdG/dlYLDMVaFMEwrPNXv0GM8+0ZnkU6m9pXlDo7xWgY3pnniF5d3F7GAVpTqfKYBM3hB
5D8e97aTC+UcvvYaSxEZ0qYcAUXcNukk156q/uN5XIvZST53kA1Pq15r28yPp01uGFMk+AEA8179
5qZQLT2AUClnsX6MEbNJQKo9Kam0//vEIUCdlsTEgn79/k81vDGVjyv9RtLj/X0P/C2eJssu5rgl
XYSFbzlpoofAUjg/yPqeNSFm1w6gmRJ+KR0r59DE0TD0fXKhYc8jP387e/x6aAZ2J2ckCjsmDZzI
UjIk35MAAuuSP1KzgQooONvvTYS+s4b8H3J2KgUSufAxxoFQqbZlhr9qUxgfPN7hZ0/pfMN6RVDa
RpsOAbli63qsOdR3Wmpwea+H1fc/zR5vvIBT+363ckyEXGoJWZPh9bmsk5F/dy7KnC5cVDiseAdo
RGebQjrEY859KDrpBhhBwFaqf0MHMO7xfrRAi5u+5eUEL++kdlnHxlwq4arSfv38NvIiJVZuHhSN
epWFQ/+d19MzFuAIXXBfYfnT554B9YF99CXNJjAhGjQtu5JRNizN4PHzm1dn0C1kdOIU7EDstxo2
YwuNtgLH5Anrr4D3IfX7eU0DrV+QMJ5gsknwfQ32mKGQvehYEK1RXj56J/EJXJoRxG1HP8h4b77j
eAaFOYMK4vjn0Tardxz2vwTD8blzkV6tWIu9j8JAxbpr9R8f7OamV63qp3tp65q5ZUSdcR9C+AJX
lFVfFwefjD6rowjQem6bDv98LDhzgpLln0ld/npDtfqD1A/u4yOx0SovfN1bAJ01xe7IWrMQTtad
26gnq0Rvoe1HrfjUIVV7fj3wpcJJYi57EMAdppT3Ivf1ihg/oUufOh0w13DFC4OtZ97t0UdY+qgE
FKhZxUk9gVjyPJaGVrE9GdsM3Qp0DZtQPQzo+kpEF0PcZ/9gkdJZNMfhy4KU3d4DuuFwP9c7kpTO
9gkXZ0TMCKh/foHucnvfZzKr1trncaWozhC3gDbttAKE6PrhXptd2TskZyMNQvZtSB8D3rSTvQLM
HzJ3s9Xy7Wg0ycP+DjAJSc01+f8saa4XGUdKl27+jtARD0pToAM5iKmVvLDnVBKryK4oLRMseBJA
eUFK0f4S1lN4LdPU7lTo1YVwTRChcEFyzLAQyRWvFlGRDKlQqrgssMr07pavwJ0kafRCooZfJ7R8
LQfw0makmB7luKB5kxgxfD4o0s7R2DOYNgPb5i3TblnQPxWwAzfGlRAYnkKDyctnQPbIrvKf0Q+2
3ObVmblXGxNnmttwGNwkG013cffBYdGE+VWiDPJJRAXa+UYeajzH3Ni6Mzn5hpwFOThQQKBQ+PzP
YhMvh8Owi5gUq6zhB+RNjCzm2Vk3aVYrS3ydfbxrxUdaQgsM3hAsIn6l9bhR7bZuFAkilR14PcmE
Cwtks/VokXU4InHt3RE9qiOUqFuNgjcVGbkmY3jLZ8dFlWiixm7zegu91RSPRc7J4h+bGaK9wIqk
HJ8VU/xecbhTjSuzZMu8pB05M5guSmkIPdn5b6PN9DaDLkGx3GoZIzXcxFTrT2A1qzPgDUlbunmF
Qg5WkPA3wsPKZxKmonPwrC0qRfc4+G/IJ12zFFfEzOLpsSfSuMlvJWEpwT1znFeg94Fn83FibeMI
ZP1tro2tzYBi31wQFbYmfGHGCg9rzTNplhbobV6DRTTWkw1SMdBk/RUlPux/Rrxk/+s1nWhgr6yI
cda7+5Mq6E0EIi2Gw/LaPi++VPTJ+9AL4NKp+75E0acqZnoFE8vWQXNJrV1006YeoBlIxeen7GhZ
ybDLe+mJz4MaFKobk7kFqW1pwmnE+gUDj/JFh0KhKZCMsJ62V11dOVwPqtFbZe+oT+a76034Vux3
Y4Hy+0tqwLHAm0rptdaH60zXmcyR5chypc3XvRvYsyAwNvRcr3MEhYcFYfA2c9/ey8WZRckSKJaa
XzjzU3T0oWZ3TK2g5SsUAkUQU9btMgHItTHUzGIyPiLoFQb+5sgni+MN8zbAHS/GylIhO5Gcljxu
qFiH31YibGOwg6CyVs4+omx46O3A4Av/njPa8Gk8FV+OJBxtaYgcpbEWHAnkhJKN/zWW9PdvUaz2
voNSFjbES52FPdOJ2s16Sw1Og7gS5LYqSp/UHkhG2zy9qMd15JtdYfjCuGMKry6H4XZu2QSpn4Gy
NQXGLRpHrDC1muoGndZOaJwH0D0wIXUYbthZxyk2vvK9z5GJN786kw3bzx1bsq+6eIAIwAtUcpk2
ScNZz9UVTFlMjzVZSZo2xasyR+XEhPReTWahoBm+Tz7bvE5AdTXgZOZlaUyFx+LE/XDH5ScQz6Kp
yrXKd25bEYcY2SLDBF7GMYhpxbFMmSq5Cgg8uX21VlNbDlsUJsbJjg1AtNzf3YeCI7ubJj0qNsU6
eKq21YEGoBZ6OlnA8Q2rm5xPRjxJibdFX2lI2PxB+ajFMtE4fCyrG0gPYcPl9BHAyqQNX8ktRhUu
qi1OuyWNU9R/8dLx5HBQmEkOH8q2q8k2DY3DCDoberAceJsi6GVGFquNAbYGNZ3Op5PpNW6Ve1Fa
TTBLL2ciPQPXnXm8ODUh7whKN/8bcaEWYhcPjTqV/n8jgSotBMN68kKL4uOnBD6pKnznr4+mlOXb
WjZn9DaBQGZX4ygc9990NYNPdzM9agYEhYVCJs9wTRgHTZICiKC3mhzSg14Fjvfdak1KCsRSMZc1
0Z5ssXKTgeZJViig0r7ljcty8ksiaMMXSsmEdaAMg/zDzU/gScl1+Dz4R6Wsqr2k2UDq7DpUzAQY
rewRQxJMsvQs7HSx3DQ9wW04cdlBL/ISBJ6IWlIv+8lzcOg7LLu6ATicMuEZETngeyLLVTN2z+y4
kcgwKZOqvhAcOIrQTppA98AjqN+EWjE31jhML4ds0zojjZUGWeNKjaTtiaAo3gwf9XPsZBaQG28G
A0/P/xHPy2b/I9GmZSQ4tQReHLf+kfnxleTGHWIxD8ugTIyXalHyHLVELbIDBofGVPHVWdwytD/K
OrFYO6EpZUo9gh+UDNOGc2bEnPjYkKMAFZfNfyf1yirkeJ9W77+5Q2UN5LPB+as8Grbx0klBa5Yi
MkNF9h75LnzaCeMguRMnU8pB/PGV7SCV0QSw9Q9HTAMxwDNxqm/soJDTPMv2lQlH4BbBO135dhT4
6OT26G3/cC9bAtPr4NT6ehz6CI24GdfjaCfS1nKEk2T7Mfa++IQyT6P7Z6WdTZxKnJ7vpbgWEIqh
cHt8D7zbffLCYfi0DiVXqAuhI/Ko3fm0oi4Pai4focqaVjncPUQglBuBvtq68WdAzrO6HNoywRrz
knVcxRWZYNFAAzWEbaG+Ud43RvKjzTmYgBFD9Jug2UYGQz/AdbMiuWTsL2EjPOxjsrc4C9QQf8J9
T53AahMigXIeepZbcM/Ak31JJfSjZ9fDJpOHf460p+eIb9N2x9OQLgzPB25qN0BX9HXpGovGdKm3
VL/O3tjbZb5ghjp64BAQ6xTvruCgXMm2JOgSrKvfhEHzjg86SYfwqbGTfHn5qpRH3O0Y346UP6Nq
4Mfegrfl0I9FIRbB/rpIRpPFFIfP1n6w3AYjG5IQZ9VelXWjk//2onjeQgb9ssp4uDSe2bxZPbtf
CfLyIp9QeQNWOSEpUlljgwNGLk+8j5DmN9dQG5DM5/da2oy/RJ6fU21ctQEuljq0ymiPjESHGnKf
UMv2SOl3vghGEDslBzHHrViDfIN6whXbALVpixK1gaEIngLi7nyer2Iu8FfDL5Cb3Ka2K47Q0zKk
bWNbw1z312ZWz5NkDGiq951IbjYY+WwStlSIZkwaKE4F1v4T0tOHG2Q7wHT1OCDXQMMWm0y7mr0c
0U+IOqD0FApx7i4GCFEI/9nq4jQHVyYzcxJ4ElvuWpO3qCPtC0Nv31ptWerOQXidWNMBJP+M5vsu
WyI30XMzenp7ERELHy0tO3msPJMamKpHf6K+auBVxFt3V5DyvwiE9q3JBNtKW35RMMZkh/u4l7lI
kUqmyqLCPRztzXoK8aUjia92DNjsEwtCSy/WIZHD8wlhdW247NTJ/9ycl1b/GoMKhhVaCCbEAgvU
mBgkfnQ5LQ0jZr68LiQHNi30zCnUL2aOebJqaeZyA3zpNxUqhz0ms2+XneSY7oMRhy2/Pl98c9Hc
HNmr6PXgO+3pRYadVc3TTUj0Vt7Nb2QFAp9DQAXj+YO5mR7V/QZdYS+DuCWjiJlEKv4ecc9mqAqY
uXktXhiNC5cK2zLMnvbnXLhg2CuzaKldxBlkMXG/nZcmnyi463/k7l8Ior8rqBxOE+NrkaahzOC3
c+g3VOxKbnqlqSdwJ9EBv/BWcyhsK8tiDD9LXAqLcgk6C41YRTI4RXbupFvKPbpUs0k2461t79w9
WytSEMYIKfAwZgMxhT8fug4j/6qa6ksEX8yH0NpFWfgoEfj/OHpNeUr9OBn6hn0aq6DVMfmDOD/g
vcbnGxXHPnRszHWQe96U2yRJjUzh8I579wXQy1gTHcRT2M0c094A3436usQiLRozP7s2hJRaGKLf
sBasFSaP9NQlW+hKuCPmV9otbay09z2i8Hi2VnzULwnzaAolJnCGjSDFTmjwqSu8xkn78nGlz/44
1mgYFqnj59GtGUKZb3mYaYTtE7UVvA3RDFqDI8Z7xZwQUWVI1LUcMej0QKr4OCpNv2k+7dp5y4nk
ebXtuoxpOwApZG7mrkv4wFOkxLNCQJAMxkoEEIM6A6ljME0ou1JB0lF49FjlozthSseiHnT3Nrp6
/KZKr8p9ssKsBgOQptTccY5HaS/b9+VLQi80Y16Kyfah8b03foXlzl2PBeuW7u/4AOjgjVfIJ/kI
2IWe/DZP/uxvrLMyXlJ9T/u4NMdxl76gEwM1mPSrs8fxNYI+n0j/LaWEUf6IpYGp4iNQ+zSZYOG2
yyGxgTuI42LLIVb45eXCyMH94W7OasPIGoP5INaDiZv0hgJJmJsov0oyWnYRjvO1EsxTsz1uHHUy
3Q2HyHuuSoRNzjFPzZCg5sxvm37FsBRk0q/UfEzzSRYUf+mOd0DyKf9EA75oLXRryQB6E2b6t7mx
D0auPh4OUF7pt6sTMAHQZprjZs4YSC5Iqxg9tRnPXtvxCRhl+Wu5tmnHhCJ/f1mNZaauDx+VHJyR
6BtetW9ZnGfF/oSd65cdBd+rDCuxGd+oBbHzmgtYVxHRLuoZa4yMzJLvIe17JpoNfoVYv3X3ofnN
RDeC3PcBPm2zwwtyOi6AnJJn5dFh+IyOsewhjY2DhWDYUO23Yg4wXXEGQatr+vAGCFq24j0kAT5+
kqU/vstrD6djiszP+0ARL4YSDvnWd6bLjM5dnsHhFdcmWmdfrD9VXpQYGEObkxgQtQ/a3GE67DXh
ur1K3fPbwAg+92Q6gvRB6TTkiK8sqS+h5Zaj5R3dMGLZnWvsS+ITHLPzs7jA86kOH1uF9p09wn0a
Dnsi4TWkbz4RxtdBdXtkpupQ4CR8DFNIgNfJaGvzKeWE7groZAHbSj/u4Ml0DC+o+wNUsq6dtvdi
klqIOmLcdC81p6/UmCix7ccEzfGqwykb5T7WXmHUu/HKcmKJyn58E7DQcvM6sFL4vud95dTGs6eH
HbJEormr7VxJqn+1sb8ArX2evPrlNa7hgB4JgCZvrNfWFGmJO0j/cxRwHBsKxQldKqaEnRzxv1jm
7q+hpJ37pRsxNJXg1ArKO63NaT4FEuzkIeIRYPDW44l4ZWpV9pxMJvhF0rqiPhF15DKOaQgOlVEh
Q6jBUrqIyjMm95hLDZ1mDKV1/MIbklH1LJ+JNFlAc85WyBJr/gpeOpQqsGXbFZanh3tq3UuLBOle
23rbrb4KbPxoK8AMD7IKVC6FxdRPhh6eCzN4PbCZh8P3rYvr0fYzG0lXzy9HbyBsBKrzHqmqpiK7
s34EcjRCAsCHPFKmkP+FwarBbYKwnH/K/jqZx/FnT+1QoF7wCLSrFFJ498tydOIXXA9kwyNbIGDw
mi33zfG0oqJnhXFSEir3XZZ0eVU7og0IxzSNwh2UIV3foXRruZnQ9ZKP0sjaVotoo9wv/FS9DmP9
jSnNvFB3NvqBbQzjc5dxDseHctEYYHp/uTozyEcpzT+E0wMslR3MiSL9QR/+4LmoOHhtBpDLystd
cyptlyVc8PwPgeR5UhiqG3Q5pjGtosM+7rQ0wzIASI+72NjDoePkJrwomAgtz269yIVSYHrKmEMu
EuJZYgzHKgeFHGI9WP4Y3iQhus2p0XVuTMFkN2193jn6YcC5BTIXsR3P1Y0rIjwgqTCS1F06iE+k
JuOb19YxmuGfxhTVMn5vyQdS+wO0MqgCWATgjPAiOR++7OAKNna9DSXrLAliZCYpwJebPyYqKsep
x/aq4UnIRRTParCuFJ3SMJzO095V571k/JQkMmrGZrTGBxIPa3cJMAPNjFvemjOpBMxbcFpwaple
3HJU/UXH5Ft/c0pNezSwEZaEdnyT6/oNvnMlKY05DE9UQHxoy+Qs6XCu2ZvIqxp9u+358PgsJLJV
6jE0IC3ZRDOOBi/feXsGyP1qnKRkxKBAcdQnDGOnDim6qAfn/tWOvyqKeAu9yc3w3n7x9+PYoaNz
TD4NDXLL69udWYy9nq6HAvmzoFn1WFBNKUfvXMXIx8HRvLGXd3Nj+t3QyidPDR0rm1D5iX+Kejye
rYZ7v1P1o4yWC4skux8uYBCu+/x3G2jylaqcQGQD4ZaE79VhFV33KLcIiyD0wk+siZ4HBJe83Kal
EULDhCU3A7bezlH259BrP1aMsV+my16UUfCIqXi326MLKWPL4nImAwVN6stCgH6WDNbXJ9XUTrnE
6uxaSAEQN+UemTtUKhrQGsO1iMNNNtuQ658jqMnFtEe7S+D4BWfrabS4/fnxBJnblDCHo3DpqNyv
o8C96y3oEg5bcEUpGz/npAX1kU4GCuJhRMh4wsjRHvZIg9CByfqIGldA6nYlcscB3jHSXL3zxlwx
/T0K6/Od47MvaCqmo0HN8N0QoH64TgBZ2JuNIccONwP1+X6jdwciUSRCzZjmf1YBXNqWzMtmyhv4
ngby/cx3wAVhOgDbi20B/+totm5wwm610cB2nUc7uKV3wrUcW0BgsJSjrnSdVCVmPUW/y7uHlwCA
8MvJIuT/7IG/iyWPsbphepj6OyPeuritlAukB1oz9IBGbEbz2t7G8ZIlnJ/ly/I+AX9MYRWC0sg7
S+iCurB9MjwzeinMxfo3q9r+5XGHYuFCqA+3VKa+Rl+9HwAZZo686sHqmpQ3dv0ootcF+N7ZMWBV
55ytoZjqx04SzzIqnmwEvXGD5W91ds3WL0F5Wk/zvcqQtwvx+FWZ+aEfGXrIhqDSwKW/ybuuMArj
wSfvJhbs38IpmZZgsfxN/i2OyDSWZKMGgKnGGkwrsYh+8OH4yZZjYLzXoe8QHfa9kxN08ueEOy2w
JYa9mhL6vv/tP6uWFZv5eSAluRB6lQdhdLlQG6rEOt/jnKxv3Qt2f9HsP/CFIIR3SEV5/aNkBwq8
Czf59RfexJ4OKR1xMDzvkI/q4JjoIKHm43gXMbERXP10mIVM6hX4dQe+LYTg49iM0L+lgZj1lWHu
iK/fMjzVvyKKN+WFXm3f0Zhr7DUuRzhH6PQ9YpMZsCWJdTmN01Hk7MEeAok7zr7OcnoZgmWj43bU
btLl7fhsXq8ZUm2b/SaygSUVdLIBv3z31/wKQnFT/8oevaludO1sPy0fpnE57Czdy2R/q7Kw1PZw
70iaTuNwjwhw0h56keO4HkSNJzGeWOW7y4oRePJfI8OagGlPMF4DOUH5yqmZXBINVDxW6z1Jvrvr
2zer50URzFyvbBjivBhSqorIVRCcuFY49FR5jnNzuZUl7CyGzUjsVNk79NrzofhgKXxAe1ehi9qE
5axWcLD/1Cna2XEwP4zveROivu9RbwEvpCJJaOb+u4ZI7eXZQy3XXTdIOE22nBMQdeEOLtlMbIey
BuwU/7MAHqbln7DjYP+O/Revg2SZrT0fJQogvvC+YWfFLx3yc9BDtBIaEsvuEGN5uTuEIkF6vO52
NJlNdvoaviHqkKaSzmvJSab4EQ9hqtJW9h1LuCeRrUJA7SVThuMkfhzLa9rNNQp78j9I3etpi2Sz
fKv1CkOGz9/HaxyMwVf/vTvdvv1v5qVzjGRxtv8CNjsjq90239cKJGuy+hdLMa1E79Z5NCxnyZSX
8pVYxW+4K5qrncLkfp7Yvsd7T4B89C/uFD/WJJeW6X4hiWvrxvNwp4fhCgMpgMprhisJjryN0FDl
K9HYumhG54Kox38YjEuMlkmowsV63+/Pg7VGwbHFNOwg/sDuFIBM0nUkyRBgK/kKhozayGnAj2s9
7xlQLnaIjkMYmzj2qrsa4R3x0hOQZXHZ3Kg6jB/hixi3XaMvKHEc3v4u43y9JQGZHO3aT/4wemle
q3Tt/8OKbRQPsVmS8U9ov1TJthS8BsiTr3bt2LKfQ9rI/UA/fQrGm/NLtJAf0y4P1lPdRyIqyTXG
n3Qn/eWCCAQD+KxSxnWngNGCQrIG7RJAZj5e7pB6ApYIo0BCgCtib70fpAsXpFWdo7tcbzL+XFNg
qbwcxikgRkFO5SV0i+yOsQpmbRkEJ86YpBX2twJgP9b1pl1ZFhvsZgnL+uwDun+dV+BsvJU9c6fL
3+QzRXNiOjljlo0swl8YtvxDLK4azX0d3DU9SjW8YDZ70HYGWIqjE0zxbJFBX77wzcdlbcPf409X
4vxunXrpCpKQPBQ5ygLKhmF0f2pjj6FTPT0REGuuARcvLGlimCYCnG3ZwuyGqECXq4ElCpCEG+C8
S9qFwX5JtD+9zem6mkUgQzNldV7f2fqumdXl6jCvVZthtBfiDIweA/kIeDR13MnH19kvP69vPLs8
ZQxbH76pJyZZYZ0VRlqihZGiCFcknIr97cW6FavzdiwGkYY/gRBN6LV+pAaJzTlFkNjK8b/NtY67
3gYunmFJuWcDVjL2dYA6ncDg9mAUs3ykwrvA7dEhh1WF70DhIn5ZbRF/FxpRYtxBWflHa2XZD1R0
PifgZq0dot5yDH30OzJsBl7IsLioB7mG1GKh6LrXsTuV2ueE6oyrMZNSB3/uTGvPTsdNAC38Nb46
rzdagrkaIx16O7dynE59gH9K64o1EEzK3RSeT9BZgmtovdEL3rmMWImQoWmmmd/q+vYI3FcvLKvG
O9O/wjV0AjJ9DsD/HrBdHBiCyTtGNUXBG65gesfw4AdjEIFjvbbGhFV1si7RX94MbW6rz10yPeFc
NE69OcxVF72eREESUwN5wcrE30Ac5h1l9NqMbG//2O9IWzAYjQ1+QNUb67tbIUlPKConq/6zJb18
qJ9gA6iXadXsdAD8Q5GvpMdgc4iLuuWTWy+WXHCqd8NxDbehybyaMQsqRiDph1C194E1wjHYEn30
PSjXE2lEhCIFxzJ+A2SgURS3x+4cS0lYzIvDSvJfGI8/njTVTGFavaPoj5RafjmwlWNztc7Fa29n
1Yu1cYn+koQ4ZFZb6E63EVulcMnaj+KqzrUV4Sn+JzFFWs9sDEnox1VRBZLpo3HrU8mI6MMpdMd6
bMSIZaR3pd9DxNeZd1T/6t/sHJE4xnLgQEVtrK/2oWVBtn27AftnDrvRvUT4G+QycM2Hix1gGis7
ufnuQSzHPl+g0Y0QbxxFNFOQVQM7ROR3h1u61Jq+WiQZl7IVBNk06pWogc3b8kc8e1o2ab5KlTPe
e4TmHX+0V0SICeutVf3SGJ6EhntfAw+zK/OiXYtjewi29SmO1ik+UEW2gWDXZPIfUCqYUefbUgoP
/ZGcPKIpW/1ZVBEJPjHUe00prv7dRLTx4uxe60WTemM3KspQk/eY4Qb8tzehN6/rPLHvjpYxHA0U
CUvHomc65FmDvdIhgCANceClg/4TDinc5khOEdnsrhcnYbDgNv7ICFiP2QsyWBsiYnuz+ohTK7AO
XMbv9JCGtXDMie83RsL0coBnqwQrWShg6E7IZ6irQnv7FQFVYmnQqd8n6HVOITHneBfujNu0ZGVP
0d1Slpgk5ixJwHQi2Bzm8G63uwoQy1DMJMbwhdkICBLU2bFBjKTMNo0Tuoq0V7zfzKQqkx1oGgwX
HO9OWQYaxG9cHOwdzfGm+bOybJefnIvebrVWfTOVemoYU7rux1J32W+rmgFUJFVkoC0sgPqkvI31
Nbdk9VeiG9L6SIjJ6ICdhAFp6Jpz1gCKfvpeg8zJ7vETVQ40swxEWoXchWBK45oRJ8JwAoMX3wiT
TE9A1AIa4/fgMv2REcDLUFlanWJZf+iGbiEEqyeBa+YvB9ErrdL73wyYJnjCrXMY/GvyvuznpUDG
2EtfAmi0y0MVNLi61ms13X9NN9QZHceFjf2z9BXDJtnjPTaeHGqG5LiuQGrN4nDHRuwMIepikaPR
rhxzUCyqMxQp1JWJWMZfiswSJSSbdA0bW7rHuPbNqdQLLM9e124+zz+212CX5r4j60ZWIpZwS322
TkXYUxFobJzQCsh4bdJm0FiRVpV3hL/i0ILk9Ut5pLfzNeQqgrd9AsKcnVaBb0d9fO/eBPLDaHsC
ZBPZouQzdNIC3GXLprUqIJOZT3VOGBf3ptuqsPs5MIN2349aSejr2XcqaS+ljISa/idtzNEBRm2L
LA2DOcAj8TKFZGyWE9dKnm6JdcZ+mJiJt6FbC8aplptmjFrL12g80ZdjK3zOvSmGsKz2IBBdclce
4ACB8qhvSLsYy5W4qC82q/fhaftFkGAJBEfChyJjmPKN/bhbbFuuUCLP2u5pUnyCJK9QhFgmsyBE
/Gl1hGdOdN0GUPFK3NfYaKH/DfAv/wLhyQMw8a3CUFjbG0AXmvON/BTZYAaWAJ7eTeiXZ3rznamI
6NPyKNCFqA4MGs74CuYWBC3oWm+cRYh5N7eoQfCiB5nuSZay2SsxmaoEjBaW22nzAhycR6qfhPGc
GHqD6FcqAdMCiFZgG8BIW/ZABEtReXoFuWQNAiUSPXiqcYuWwDk9w8Guxj5rE+OJjzW7EiYOlawk
bnTuc+l/Y4S0G9fMPH5cAvlZ4bKePUWBP4MyiJvgUNl8g1EYpfYdHx+R+kbUyfaksefuN/LAYY76
e+YEdQYlnp11LHMvMtZX+h5+Ij0uU38StgQxnugiJMs8N+7DSaJgCmyFjI3+LFCARJde9Vv3sH6o
Vm66MV9xDTktD2jbtR5CwIVLwpjwprFlOKC0i6VgEt8EEt5IHgUZxTRbhXijiAsVdxssv15AMUEp
/1nfG22EsahLA7s7UbwRPkvt9iaHRteXJFqpkDoxMYSUuSPrwNMpHR/K3VskDFpg0PR96UtcEN1S
KbO60efLkXxwQvbhE+8bjoXP/vAAVjjYot1bnvpljUQ21ku3AtQ+fKCWbBpKJVN8McbFcS/HXrxV
JLA4DQQ93gvGVnqvR0ISylZ3aj7L8kSfYWsunykeezGn9XLIGwc9wPOuENBbwI/67mlj9Bgr5lqH
G89tzedFwkm3xkiSQFGaKORIdE89PsdaETxVH2pSlOmRRsEbbAXQZ6/vEmkFhXeAih+9gN8iI+8o
6mMXMtPS5gNuphOVW6/sL8yQEVW77ogNQUQizMj/iZ3mUd7z8UZwjuNB3jFlWFe/rb+JKyKfF3Bb
6VvIstj2Kw1c0zpkBzQhq1xdrUM+qvk0V8tX44r/lCePwRibQ13O4dkoFgkxase0X70GUWaZiAOh
rp/4BNVBVsvZQLPGyrSvpkUyvxCbFxUbNSklDEmeWxLWbXO7NU79iHKEOTwUbHG7F6AZKw+/qSmv
WG7tuiFt7pCsKqNIFYHeVp55+O4pNXEtY4DhT7hAXgHqQrkB2rUv+AUnT/cJ43XVo0X56L9g+r2t
CDZf+q7aW10pFq3NAbSLPQcAjFQy2oJqRG5r/bVqsj5mpiMCgmwMdX154FeaJeTOpW1M5p+CDLFL
2qWcN1yco5mUTi8d8aMXcXJKGNhxj1brBT0aY7NmVuC/B8ZCE9aCtPb5fRE52WcsBerqrP8RV3lQ
qxTWH/Xozo/5QlWatRCJUHxTZWe4UAf8iCfRFUjmBEJEZOhPoJxV+MpMO3Z8PU7uK2QTFFhRjSpN
HB7SwrdB8EIqI4o9VebaCFDGcRRxuxPHb85NKQ6L6+TE8yN3lw9xdW1yOeMWQV2c9d1BR5EZBtyO
6Pl0EB+gUm6jr/WhF2j12PgCBFyFcYS5bQxLX2RtLymPLwdDlNCH/WKVQHsHKYj6AR6otsMCbUTH
dUhJa8mPfJlcfSLABtpyCgiw8mIqKZ2z+J75Gtg9A6VOWYCJ564vV/JKyBMzX3Dm68X5aFqklYgJ
9JZ8v9qtiwxoCkQJlzuX8+k1ChbCsni6KNBxPTFPS0pAzTPV/tDrKQXKt6OoeUNGcjrihZ7NGdJ2
wcSwUN43MborKmq14zjNCqJq2QxGbOglDNwp1Rng6JlSdaB1lBOR/UUQ3ZCmHFWhTT62r8x1EwM9
rRklK0e4l9U/o8QRnLLzYBvGS1+sMCDCaA0VceOAoWYOZD5tO1cZFxq8sOONF0ALbc22rxhmQTiq
O55Z55whf2a3GFqu7GGb2vlo/Nl4ka+Pi+JHxSsd0EqRLP/cC/aOYQufoHjOrimaEpxV/gan6Bar
Nj6eVgGbkgRaau4jpreZCif9EScOfreFKRrQCqjV60Xd2eiRMYWnPy/0i0bFbOtG9xrO8iyCEYzB
zaYP/8WoL1aOOvSpxNMOQ2rPizE80zAWitVThFSt6ly9pWGMEuZjuo4ikYE3hFiTkIa1T9aGSrsX
9k2o6Lg3zpJU3uc6trSJowZ0OHXzijm6Bld4pvhHdA/G5qlasaJ6gWGC59tYAxpK7F6+A0ge/bbS
Ce2NngY/8NTvCHeikUD9rF1RaEmoiTIQfQCuZG7LmqI3oV3tu6CdrlayZYBIfwTJTQEcX5l3HSCz
2J13s85xVoHDvMk75CrWRbp5knnD79O32zqOP4nwaqW9boxcecMxbdP1k12T+I3z/jmqkN4b7ivx
upNsDUTBv/jGVofux0gbgp3ucJf/UaEi/s6k5q/zHuWVoS/hmxA3/Sv9QrDOiJ82LqHZyjSwFtp6
UyhZeN2vdj6SDfmJ/7CXZWv+s+22/727Dor6D94rUygWswtI0JjVKTu/ZPnjeuTnJV7hS5hc2tzp
4vPj2446QIGdu0Gw1wV2G0GMNUmnuu98HA3XWHpT4GruKclZIVfSygNkopEvPRYs1nNdjfxJ7YbF
siu8PP1nEhbDUWq8ATGACyHyEg8SYzjO6OBL/idZ+X6CFkBayqyz7gxOhMHiDtT0XPpjTQ8sOLHU
aaIAmP8jAb9Qz7HY1V+aeCVX4LdnXnI7zaU+SXfUaIyDGPMIXgPqwzrQliWLHkGBclcZF9ZB9OBe
J8qOhtMh7EZm4/Am2FLWxDHkMW3DnrD0LOy+3FPdYqUL6vS769dTn9hsHwfZDVdNR9Phy2Xudphw
X39s+51Z1+lor3OIKmwDrRwLpGahCvbiYysOIF5/LU1rp9vgxDcq5wIkmbELGqCsWoLJ9YVrt+2f
aEXhWihuUi/3iGkJo5NhhcW8u3/LP30O9vogv64Pe/ocmC0ESW1F/ZQxgeODsm3R5Fnd/Ac36WKr
fceKd3z4gJHcs2Hqobob8hpdj61TPo6ogFPf6UHhRTuvoC8FpjEDd7C07cJJWnIWN25lPWJxla1N
N0bXdwsSaUmM+E/bT0bsB+LIEbDFjX6Lfr1+Ox96JdI/x8DJIj7CKbPSB+nWYnarB1KRh/xYdhGq
SyUh6zLkVS3OWMDuHdm8B1mvrQK3QPMEFHnpbhp0Ze0AixZpsZvEPtM4oIXnRIFI7l/ar/cHDQ7Y
GosxttfRNNh5Mrb95Ns/KtRkZCg0ieC1+eBtvqa6zSMMh1bXPBtk+Qmv+1EROAu2zEt58t9WdfUq
pTlha0Er+w4X9puiIKvH4FckskirIiQK1nJfUrfVTbbr+1EXBdlWbalotWHypIdFWpACwOG72Ure
2zvx6x1mef2wLaa6hu6nXHbFSAHJyLczFs3dt9SjWifMX9M9Z/Aoss0kuyZ2BmPNWqUVyOaZsuBU
rUSvksAm4yip+9lF/snjKjQ/3xSWIlTLhWpZMj6gj4vR1EgrlLGkaeXgfYwgfW1xqoX52/zCGJuA
Bc/m8QOBksKZTcot1bsW7Yqok+/j7GzWW48Wqcq+Iiz1UeiHhj70RshH4ld6zxjrU1GaZh/xl6/a
+Phyc81GpD+PnxYjry4F7Wk5VMQwOkS/s2Si/7wMX57ZIMwT4ATI29luS5+nzPOZGi2WzMwWSdZa
mH3Gy5qLuYVisO6A13G9Pk8ug5/FFsJYR7i/iY8xmIeK9E0cLiZtEdi+s3WWvKM2pJRYFOiSR5Oe
icUoiLq3NqhQtzKsDrc6TM0t/pSoImvdp2cSBdRM3SxBUxt1hiS/340NrCdWn8rZ+FbaEDhlv8Ki
XuA8qViU/Cxrthuy6rzIvdmHHJLLMqHymeCtqMsIjmVGPP5fFxSBQL4ClCcWw/B+I81oMdPVMFTF
PWZXaOPNdbP4dFVkm6y7i2d05nSbZk7+4xQWvlah3jKnjBIm5BWElAPitj7/RTdKQX+VRiTqADp3
q1zLNY3/0UgkkovZkDLo3/q/6KWGsx9fjREIL2Nv4cBxaS9oNlMO78lqdw4V4SdbVOggXor3A9H/
yO2zLhSRDo+gjloxlgwbue5HZLbfg0OxY+XCSXd0DGkR45Mw9+pNmqnw1hvhs2lxa0tM8wPm+LAf
eJCQez0h9ATN9L+RoqHqnmb99xB/3weN2MUewW+3/zI4BndZ8Ra3m2+QYDIKkNsHpXSZwabGpQmN
hShMN1hC/0XeFRywuF4B6G1MntAkKiXI3jug0I80kOZjUJ+uq+QECs5l18X/xGTxP7UZ4pgE9IPp
K8wRhXunavJ5el6TRi9/XxMhuQnQZkPm+kXnnVsqA228WNw6G/OvpIKtUAxcHaV1aXuZ+VGFYmCH
RIZcsa9oRlr0ATmLXVpkmAfI8m5xqfSrxiVUmsBCFr/S+d4S4iuBN7QJPBlssrtaqBT7wnpAAzDw
QlIhRnRozRYv/X3VISUUZrqZ/GO4sAr1AFvPnNap4v3oddg1/jkdxNvvRZYu99uO4eIZqop18KLC
HxrrtVh+6KicZf7lhxvdMphLMbWMtih5mOYFtxRJy6O7ANLkjUubHecISXNYs4xpz59wtF30Q9tY
cbvc6wbI29wnHZr167GcwcrRqyPDj0GDO+3WyaJmsDCIZb1wHYe1KOmmmWEybPlkxd5S60FdVVLc
wUgrohNmxWRGU4heS8thFxAz0qcjDPIJ78MMJEqXKFE7aUypNOrqNCe7ubuyGERLqdxUxdf18T8d
BBHJ/ckAo2Ekdz7bk5IESjum0SDZNG/IFopUWpbNEuuckqDUEyAxI/gDWTTLzV+94e9/8pm8v61I
XAR+hFhSdLe81teJjcJPGIH6bqEc3lhOj0e9DhrZGQ3PHGZm+fOTUFTf1vv8sVkd08G9wdnCdkWK
rwR+3aFc0t+vThWlT+vGZDYFagfc03/yQME3xkwO4KnvlfxL2v5uGAydGQy5TpQ4jeKn9TAHzBDM
o2MDb5JsbN5RMSCsLipvzF9jqGFjO+uPyVlFiVd3AhPXd1RawmMrETHsIXldsKoTH7ifYndMa2Bn
+Tpm+FUJ62ehWNKcK/dC4QY/w7+v/lo6DFsVt0jpYYUs61PZo7QPqYtRV4ak/lNP6BA9JmDCYZcX
v3xlGYJvQrAXtZvjyh93WVhbjl2Ln3ZDUFTotGzmIIyjCwXuxIeU6qDRDWA/hiMc7DdZ0XP7/Hmw
9tqibtcwfae37KguCCsN2q4Z/TudkDx7g2GkCvoEdfo78bxN2vCdCciuWJsdmxkRTGBrU5KNWkHk
176dkE+VGorMgTZpJ7Z20EtaRnGYDpmAScFCDAhPB0weSsXuOXksDmCMoxi+CCOebjMZIAOdIocI
iMuVCGuwmxnTMX8feRo2YYCdMrPG6HEmNISUOIWz+4ehbvHbPvy4GTxrURQb+aYhM10nUXiximTh
FxdQTEB6TAcF9+5XP1NEF4oRIZ2SoMJLmYGZPpXYzd9G0vAGwQ==
`protect end_protected
