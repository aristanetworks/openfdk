--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
YtslHZ5NBLRXg+P5QcxolVADCR0rQx1lmXMwFEivtNO+geLdS3e0nzqGEmZLYc4hb+YiUCG2QRBD
/u7eVoc18QSpL3TCCbAx4qk4medwyepn3bRJ/8KqNMS02hamqDMS2UoiiAuEkEfErXxLdHVlhGKK
WWrF7s8jpjZgx0N68RKa9eM2CdBpiMhA+hkB8+Eb31f/a7wwPviJgQo6QNPkY5JyjWsCMZR6UrWa
2H4/old+B8vHuo+SYtAdfM+fwUALxdEcX8oSK5+CotY+uKGUDJCrELNrXc+c5x9BoZDP8kz6ZYAh
himEcboSprn6T/Kod9ZYJM45uS77ABCJnPrasg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="qy72LnnR5zFICADflWeuUTPd3kMzD4jPmuSTad875g8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
bIhB5YxlVw5NVcqjrAEaCCWro1Hhhc2A6cvMREieqrj/AzT8v59821CvgdU74cMQdJlGOyAAD/EM
ehlt9VvnzZGnBpznNnTIDIxQj8KyHweAFwxxr1yXwnlJemxhibg5lynzIgymNlzQUy6nSD9ZVl9X
LH8IIcv60FUyouQSIOM7a4uaF316CeiaNpGADQn98ApFX+E5faeCplzbYtiiqzlY37WupR1XV8qx
fc1GPFSAKKP1xZdIUbqejUo1W4jqg5bJdEWJcfCgx4uH0fIFqZdeqPOjUW9lsae4xlv7b9k+NkLO
A+uoH5YphbQY2tAcF5juuAezHdw2YS6iwIncYw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="3a8n4WWrR0s3eyaHgDYam96kBwN/m+GOD3/6GlVE87c="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6560)
`protect data_block
G/V6+hWVpWISaM0K2Pv22WNYFwDxgmZD37jhEuhnKgDw6Zie+y5m/QpUWMKlkTu9KBq5kSt97txj
RndfKWsAJvzPbRyZRhxqpq9nJONOI3oHLmNOKrxmNfF8JymAj8s/tfwXkKNevZRHdcQ9zJO0OkJF
MR9GGMn4yFmeaiGm9dyJGK6R3/nkODCOUVekxwgY+IkINUVHdkObheU+wdYztPy2e3UDyLlBB0Le
8hXlacsQ5VmarIwVNlVClubfQGRTA/LpMFkh6PDtXdVCrl34B2tSaTmGnyu/ABlgBk1+wq2SVMS2
ZU7/pYrNfE9atEaxEdYpNwZH6xvF7MiYVE8BqfUeXDj8ynqrnmPAbaSGKxc3nM9TI8bFG4pnwg6P
bZ3SXfMz8WJMe0jL8buOGiC/l5mxnYkBH8IUSl8qL7DPZcgoiD1M70jxYJyA8bddIxQ2JxcOC4hv
R3xrx+njQRZ6aFnwrXpyKaSysBFvLycrKBj2eDa1jqzZ0w7vgPiUwhf+9x5P9pzKUPY6du6cVAs1
B0GxbhYFeyGDELmCZS1PMMS64TlFPvCA/Z/niXldIBPoh3ulJdeMEU8Aa9RcU0VGukhfTv3pDj9V
xzMuqGj4OuefzkZFTjPVkfN9jSh9VQ+ilUA+jbBDY/sbWd7I8C1ENEq9igoFNXoO7Xp7m6oL8oM3
C9SOD2bkGVUgOI9lD6ClyUPSf3hSSOVRV7BzTpQaj9aij2hESKScV875tgLO6XHAJtAV+TcBKqLt
fjEdLv9ah78tdt7P4ZozbCM8TfZ8G9s+yLC0o/w4R12eKZxO/zPiCGBAIj8ahfs/nFAKloGkvg+t
19Q+3lyltU7cE121t+YwlHzVs6rLrIE1eEu+3AYn2z7mkLIy9tBeqdje1DOqOy/vxSpEws9FHvrS
TFVbiCxmOnmg+MbV8p1snABUE61xBJPBrKHBP2bVvScATY9ZPvd487sBWisq2ujNIlNsJr5CQN90
kdEjR7x/C0nlKfTqgJyLKu04gP7e6XV9P707gAn6fDZW/WgFm9gAiPciTcnMomCpxcaXhH0Eid6i
vNfT/n6gWLhc8XMwscNnwCXa3339rSYQKrXV77b0c7jOogkZwjWDXBT+ZGAjU3SzWtWVqaiUm6um
bGm56JBqD97YmmU2Z4ztrS/j2rcm8vT/PSS9WAdzAq/P21G+3ImlWw1gKyYO+xt6wCv4PioMtJzr
CZrGjGVP26Yz1X2oBrqFuSO5I2k/UlFdjOzrRkoDLspGF/ginQ8tQ0NYVA6EpkrLmsWT0HNw0R9p
W2gJc91KURMvLnbC8+/SjH6hLg8Vc8MagiF2sUWmr9+MP3SrCRaxk0FJLnrkTURKU/n6s6tpSZyi
wIwvNSNTl3MVUxhhz3RYz4X7jNfmqBAIF/bGbO8lE+otGOmaDMAZ2fQ1KNUJiivRgXqMtoRqeadt
slTfBAxi2ItY4U3/GJFefAKVPuwCtI+eM7LeNQLSb3/h3bXYww2QW9BJzOrqdcahIPt/SFZ7CDvg
yBruJh9NoK7obZaYe7AG32qM84SUBbTNFpn4vtaYeXunnAwJwih8RiU9eZ9+vftWMFi8wVyE6lin
v3x05ivFIFyzSVawNYr1g1HnHaECbpJm8THdXewqIi5l1YBGzk3fA2SGt0UISU1v87VgXoyrl9fG
ogTeuNucLosRUW0QShU7XINJd8hFJDPncce/fUS+E9QwfhtD/xKZcRYgOHy9EsOxSzoaYktDa9Xw
1CmqIwC3LSZsdrpoXZqAcutVcatQIptNZq9hzvfLy4jz9p3+Xeiev2uCf3p5p0g6OaOaMJp424aE
crZGoPh9ojTJbyc3NIXz7hdkeNx2QyuTYvmODFn37ZP21irNkyzn56JqvuswKIjUKF/wfLgAUkvX
y/eH/ho3rAJVOwLylRE2nZdGXRVCOMrLpE2Ugi+XYY1b07sIi/qE6CSDdLKCoGNj9dTpdnXIjHPZ
4yf00BOJMA8eNdFH6AtMVlEw32o/1bVDn3uhvm7OWFgGIF4Dc8DCr+2jXaNzIxQwKGGACKNILx3W
lSPP1mf0lnZhZQPW9bMz6q9aaBnuSWlZEcoRqNr6dv564kS5KnUK+rysUm5VAFNEWN/6MLdwAbDn
Cctu6lP2QqPatbSZpTQrAWAa7CMD/JX6PcC2OxcvHgBbtPEnG5iOYJ5OWt6ENivc7gkxC6NUo51K
Yxni3xGrBO+Nqe4/zu3ivzdzD/JlTFxn6wpkEW86IBtQFL6C99hgBG6r0jOpUm0fhMvip999ugZm
FPLFh9BoZXApWkI6zsbn8R8urrHYUVLabAyYBQ8OApYOLM5w4QuXgagpkp1XBRIoTR1RuJaG/aqw
MSMiRz5TAd02nfWt6qcFqaE0kLPAgCMLN/IfSciVWKQFPTSGpP7Mhin81GNadnouUYCrPZaH+XWF
wHQkgK1EhZSkXevRMFxL6maAF+1AdH8QKKpcplmpbc/WoIt2qhvPZWqy/OEIHRw52Z8A9S9dMqkt
t/Uc/eIpgv/ojWL0sB2N4Y8UQKz/KYKhqVz+v+rvaz6tXTqNCmvCn+Ua3TeYyvR+olI3LBgQLqz8
uHUlB/RFZVpd/2LTdTxSYGrOExysakX+e1A/A6ubanCTkIHx8riobx0SdtCfoqXhrAJ6cwZfkngI
IgdyZSw2QcIr4pWjqMUeJMWRQSSBbib9wLhjJ5J66t2WeaSaJ77A9kiPI3j9at7n3uET6Lck6jmZ
Tq03uSGSXySKrmaLj4rdR4h6tC+naSAziaQMVaDs8lIEqRYk1K1UsOb6VFTKaNE3JPjt+So/Ocrd
yoeyd1aKKz6akDldRXYusQSCqy0Z0mWtmVNVCYK+6d2o3lyBIGh6QgazwZsG5Tv5FhEyfrea8XQO
N6ID0AVpEr9mMGFzD/+edP0qw9C2j37Gc/CZ5t9xzRWwD844lvqFE8v8PG7DSAfkpV3QBsqq9LsO
Rrof8VWdIpn8u0YtzLiT/URE6CdrlrAnb0ZvPyfO6sMbga93Dsi8xZu00wwC31KEx4Y9FKfwFlOK
S/LsNqMZvSnJ4aMhvaaJSvrhW0bY+v/bcpG6nlNYLddv3ix7+6ltP2cqhsqzmKGmfsU/0MShFJEh
pOHkZMr2ya42vWkuHDd1ssg7GN6Iq32P7NXIp0T2suKnnXLZC68i5pMPJKsfsWTAaUQx+SG9I7FW
IYoc8foJ/YcWMgmy68lP5Kl2woabgzw8vUgDAc8+b8suAkinimpoCcVfl3D+AQspkSQot5b0/4Pl
4djuDZkBoA48EO6WK7G8cC22/tZRAk99RwvtG6PM4QtdGEfAB5fBLBt2KY+3CX86DnNA8LZkbvs3
XvJQNW8i4rBn6KaA2YE+BhjM9oB47jWYx+GEMUheBGVVB7y1ljt5gWTUFQmnuTQQucDDeLxNwRce
JX8yDrwkHPNloyZvAjYGssllVW2f0QNX5uuCu8j3xmK+l0N0bkjQ7/2YqWraHOQMk/E0ofEokfpr
SpLcqrFpUVsWmQO7O7szGQftKRBcBSnsugSpNeTBylBWdWU2zNGz5G78ERouJZvO09G4T9brbhed
NPSAv4IyJWVYdX2UhFggRPksmjee8Tf2c+Z+gV9A47oC3fI3bB72g7w2EHx6HCqvmX/L8SuFSOhv
FR3col/a4DcQdc0E5zGYdfXcK9xeM9GW3sK0rQ+yrV9J1UiWEpVbHqo4zHbweB0Z3RAAuvvihjw/
Q/qv/mF63N8He/uSAcez2nj6tDyics9qa8FaeZDqyj0fhv/NQI/LFlPrJBbjWuVJIdTBKEW16STB
8qVgiLpjGqluVRFWEBlxCNrnUiBE1YGKQBRZ8tVbqXZh8CvvlSZyTCRHTE1Zo621rRWQiZ0OO+OS
IABCjQUzDps3XD7WI06TAkaePQHtb7S69xJwusEXV6vvHM4554+AmPetCooOrj4HBVAxbOFLmyoP
zwVlN7D6HAH+lWiTo1CJgtUO+Wwly50/IOYopR0s/aG9aMWg6U6EIkqmUwpp+2jhbjqRGelkQaEj
TUGkg/YVAQLP2ll4AOOqAq+aFCvB+R7tmUYG0fwHpAglWCdUKuXkFmSslUi3V3OwzLHzXc7VB7oj
L0JEJFkVMeDq4fqMaQkUkmbmWasPAKvxsIFRMTNWg7/Mf42dy5c5+ceeMOY4onsqOQvnO4XqDXu8
28avPfIweQI24DCn/kfnXqJHunxyNAOpyPYoDBzXDormiPvw1oZEjlDiTcB5KuJR14AiTI/7rm1U
bgnkZcQzwGRWlBXjH0L4Bb46tcc3KbFNo7LuAr/LESkzsRq2GaoOnf+ALPK8qVXqQaUq936iLW3C
s4kdu+5Ej19W/Cfkx5bDc3HoTd/zhK4WFjjmAU75VB0DXZRWI+qsupzBe2KFWb5D9T8gAsPa5j5i
Wfm/LkKwhFU6nxtdNcWwqV8S/Oump+mGqIWj395NiiaRKql+GWjb/A+vE2irVoqk69r3H4iWnmVF
CqtnI6tib/rkwsAWBcWeF9nWzRmSH+4QiPPQe1VCFYng2PHH/xAPRUusuFYMOi4Ks6AYOAza5N9J
hNRkdPmFy9EbFtWpp1WlBHK3D19KfQyQPs/REkoYTf68Nkp/rIb0qRchhIwm0/J0K/LLsHyz5MiJ
xVDFyZta6AIP5q2avYyQLg2BDvzgg/pfJxjED8XzJZvgvyDlu1exXyPX50EYjinoX8K6XwWZW32O
QWOmXCVTDd9Cvu990ueEQTKejw0Y5lSgF2pKsbF5n6ntL1iVhExCNBWsPclCk5emTv2nHQya5QIb
DWBGBLPEuVEzSkbINEaa6C6HtePlq9hG/+wsrq0eFWUGxr58mJfqbUCmP4/SIh9xBPR5yoK66orj
nBr3yPKemfUzJwYQmJxowR8H5ecDY56p4l6s1PcNWGuvNA8U+Tku2wrwSESqfd0PmdQM80eWxsF2
LzM+ke/RCNJ0fEMD1NIG2TdBCJV5hfcRlptXx5jFs3ZQldeFiIue9JnaGJdeImJJWFLddluXgZ22
HeLKiqnyr8pClRxXA66KQUMejzxrCTpC0PPpGbpIxG9y5rRL6FWpKBhZk5FWarbywlZghTno4pkP
YQQHOtuchNwc3k9oV1acO0r5UzSGK/j4Zc3imPF/bDDYXVIFZHSxzwEI9+HagH2hZZTYOeQb8A08
q5xookwJ4OXkqvUrTsQbZzv0iIu8Pyk9FeuXixp8eEP6DzQKgVQ5+TITkJFYOL49fiEJ/tpGZd/8
QqE56kABvmwGMVmM3r8yl5Nw/D866duWih2E7jb8cGs++TgtQpO5AryDH/YytQXCRS5CS/A1tU6k
Wz5O9uczF/LgTw7J7SUUqZnuZ65oGJ6tHYHaYRGGyBr1Hy8s+Y+xDnvVDRfKxwbjqIeoCA6mUaJ4
27qoUw/CvFTz4m1iJypbb1M42nQkDOeC5fjI51SnZW87aMNWFcB4K8IkThfEJZizspc3p3vRmABr
S9Lox2GDRaNb8CHh0nfi2tCK4YU+0+x+xTNnNzpc141IzLci9dxt9uWc0lefAnfgvdccNuK1OfXx
3OGgeYP5wdQ0VQ5XwHrxW4F89NHWERE3y5HRQDJcCLA7AuIkfiBwQgLhf12jA+VYeqUfyLMsagaq
lYWGhxIYsl13Z4gQbj3t27xS7TvkZ2W3phYtAR5Gzlb5UtigxQIzsE2G0RMrahWT5BGZeKHbf/9i
kxJwNVcvd2jGm6MCcainP4WDuIiiyIahF9E87v78x0x5O4t6xVV8hV4z2KFfGNJKJWoDLKJDBAp+
Yu/x+tdnDc2prQFzYHxgChfnXUG98Ty5oP3MSZlepnAoeExorpmOLuLGZONSWNqqGO2bfIN6akzU
Axfrbw2OrLuWOX8neI30Sc/kwXFspasrAw7t3e3O7JNy6gnWtX6A6mlVEVfpCW5BB05fTmtO991l
7w1LbblVkqcK9RZ2af6MSJzAQVWTQifthRBV8f27+q6YxVsVC3GpLqpitGzLngVSfn3Meb6jx4Ut
Fdnfrk0v9bdoCj381qjkV+vWuaCXbiW1PrIvHEz4oDUE6dcNLf3HrerPwBNe15VRnx8S4t3prpCu
aFCdwyRU0p3lP5kSHRScvVnIVcDrz7nXub0gwZrt3ByLA/Gy3MKdQKWCqGyDa7jRvcRegKRn8LNu
kK/U46mRSo1+x9jSuc37Xv1D06JFWEsrjnQ1CiGZ5tMn6vi6TLYv+iTLuxxW4x5vX5iuEbW8RALv
1iiObYBJTHSxBHP5Z8Jdodnd2hpe24AxN1lVR6cXbOOwjWSYIYXa4Upx78El5mzKCdtNqafJQfO1
TbzAjSg3r4F48+l2PgoCDh+EL1IR8J87QTmGkD46dTAxGDoLo26Ez1+sAt+ylj6UE7AALh8Lt5XQ
AzZ5sycVzEbO1IdlpxsidRpmNazYFRksaHbcyfgb4DmCS8AMdVYmHtZGYDXMi1ZPD4CGubxWWH/k
cRyxK5mkFZ0gr/dQx+B/RbmlMZFU/Z0doWhNQlTXxeGWboF7fzeR3kA3RPQ/JEVemauDni3PwNDL
KD0Ek6WJpk0MGVZARz9SZSQ+66ORZe3nZxHaiojXGBufYgUPiUUCjTe8R9PLALV31yeDWsaUcwU4
nM0eLKOu+VgSglX86VI+ah99wE32MW0HW2DCq7qHA9Dh0cLC/ouqA/rqFGZcMpFMUhBvOC7B/ZWG
7OHwGHKKt73Z2B/AMqZfnNQRUrYRS5fB53by7gTocP331Op3Nj0aClAU7ELS6kByaTNFQLg/VV5k
bSkUULUK0SdbLK8dfsaXuqG0GFNwuCcjfaqlefLjQW4loSUfIliUcF+NxqcJ7mCZfq0/97bE32ZO
u1PsherZRxoPr2yTJQV8TKrBBy8/oasncEjfxi89VaoiQt/TUr11iXBuqnfEQS91B73yWG1OD6zZ
zswX+oj4e71+cvcBxJ9dwSlWUr4IdxiQUgO7FA3kKQNPW/k51gQVUWXETgVdZEQePUoMFG9qoCqr
DTm/w5rpsxKnGI6RXSbO7nNgXrT+oi628S/V7zJa2QNFvcGg+BhwrGIuUrwXL8MdLpGVkI6aKOsu
UKicb4ZmeJJTYqUVXCi4V3TrYJs78oMPVyuvEPEnECtDTnKgk8wknJWwMquFSO9cALxYHwjpNBHc
oxEZX3zgQVa4gJWj2BYzNjw80WegZ5tuNGDSpdhUWhmlT4Cq9w2AmaFBI6Vv8ax/uuBL7ZIbNlCM
B9oYfNXXZMWEpV1ei9El/dmN3NzFZLGrs0Vol3loKhY7NtFmd6viQk/X4y8sVytgVtIxZatLk8WX
lZ58ZxOWamoPvDi5X/pU5jN7fMPbK5AjipUXgN3Y+e/Djv0Jf7MvueD0yzmb7zyiTvAfHBqXIpXU
VKjjplo2K/X+1DhHj////d5SYJnYIYOQo1ONiSN/6F7Ym3XDRQMZaTBQkwsJJKw6VeyY1yZ1kyfG
piaMGNF105EJ6V4h5aKgct2XeUY0dqPzMEuc37sdo8RxQYKM7IF0Z7iSge8wPAs2/PkBavjGTIqS
GPBIa2LyAmiNHSWeXTENL5td7pa4DJqXybySanws9yaTIgQqPSbqZR+DK21zI4LymI1f8uIoZJ9Z
by6QiLr3UXG1blf1rikL7dv/AP0DdkWVy4d6zX2/7TDze3v9qO8a+PfFrMDw3D1y+BNKJgO7axv3
G/bkMxncym7NcjrJwbAdunutM+f2AMNMKyNx3vIYEnEmKtDUSWjuU2896lD+IiH+Pq6cjWmte2dD
4NJ2jizJ9JtIWst8+d3V+MWI8ppm9Fl0pNPZrI8+LgLv4yRiP3mwi+txUTbl9ouft6zg02Ej+x/b
m0rfBNiGJGqKe+21acQRHcPA70jj0SEoX6FaM4OQKsibq2TNTYrGcI34S7BMCa773W4LYrjv8ayk
4GkRb54KSAS/0w5RqNtZveO2z+OrVQHfaiFWTcVWsv7KB9QRe9xKgW8o34ZFzrUVXa21WiYcIpTh
Qg0e5oHlV+JU0sE/xdkHdHwLLeWRq2bQNYK4IEP1sOLmPRNlMuYhV+a15AX6AY1AB9ElHJuB6LcF
u6XG877+8Lolbbc3KPQ3eZURDj52QFNO30xJL2bwqSMDciCx8ClTqezdeYiarr9gDKW0scAZ5i6n
4S40cr4tLhX9MGkZqxwTt2Y+9GRUm9RItdMarfq7CrVPzJuxACAXatefZ7e/V7FB8YhHBooU23EZ
Azo37dteDMiACT4xUuF2+QDq/duojJ4CQo+R94/gLP1goHiwHR7fKUCOSwG1694sWlEP5ghAzXn4
CL+pJb9/sEGVxwpUzBsJp+xGSCbDhWNNqfnXJGIdLu1lL2GUzPR0UdPHLlqQd06jiFrjDie4jRax
D7MJQhW81TwtaRaqcoqszVKyipz0nzeZSp0QTXWABzpCaO+S3SOfwmtZYmphxBtLw8Tovg80JTO+
TVjYXZZcnSwB/vKg7uI5+OIQqZysIyZ81/ogc25oXXu9PzeB+xPVYz7Gl9VgH5uKcB4HESshrBi8
X83fruclVlbMdSoA1yiKMKw2BRsafpc7f05czBHVDCi5tWAHDBQgeQrcyOf1eMzwCpK4UbVJJZnG
Rk/t3DN8yTPar/i7RiXg9DHcsLWauTuMwOIcwLXhPIX6Fc1VYWLxJjoyB+yufOOtb7qWqBVjF9af
3nN5bFTTAVpanq6MSyQFm2apNVkBoYJ7eGfIr54RITXDNHoYfDKnOP3nxwShVs6+ymvxtBwWuKDp
Lzkr/EQ=
`protect end_protected
