--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
IzCx5QbxEp1QVailOI5RzwLX89/LOVxLgbxsTsICgAOQqcQgRHDAErrhq9pi42GEfbdcfP2adwHh
3ZS0B9FOrqgPZBbS6Et8xJtsyBwOponsMWZdKiK2KGptKocVezlrWRkfGdKqP5PW9BxWEoDRIfc3
GMqrZ5ky9A/iKLnpY+HB3Efoea2HPCAYTdbNVfdyt3ivA6oDRE2tsIyusL652viQAEdlTF+fto2D
tjhgoInzRSDzV+5cAqfz2FRX3T1VEjBVrQEDmn510QSpXiJdE8lF83BvLsKDyj3VeLo97qCSuGv2
WBWm5g9i7Eioq4j3PGf37bPVMI42diypn6Fr/Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="qh8DPQvmGtk4ThJc6D9/ZxQ+mHO4O9sSEztKn6h0uM8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
bfsfuFrjRzbuv8IcA4v4zoBUzhHAUNfVK/bgU7a0s9ynRBzSkntxBnyN3gD8VXEwc/HE3X4/lQcn
5s4fwpjxPUzVV2/1fc4G7EBPqRrOVzYy7WWHTEVQKQMPQWzX2JQMbhd2yTBnsj8jIsqOWvR/c9qm
bO1OXFiCnbKuSoZUVCRhKt0jSuUGmCthG1ufvQLVZIMuni5Pr9hXyeD+FQl1LgK5ddj98wP2ASTa
O6Op4Ieorl6MNZg5Wpa2RPuD4cwJKMWf+cx5CAj0xsj2hEbMkovltxWOtYe9aaSgQA816aaXFYWn
Jr9yk3/gPfgVUfUBwZTTzwp+C5LPfnZuZoJ3ag==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="RDqi0G47wvYYWTo04XeCB3+CUGScS3o0FhN5IeM6VFA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 38816)
`protect data_block
WdXkybrLH1CUXS+ThYDtsDjm9Oi10AYl6B8oXmAYUcdxRQHX6x5LxP795s6pTVZwLtL2QX2BzEh6
LZHwpZDwkJOnGIbCDG+tQyaHn+AhCt5u3tokPb6V7h3nRJaCE/9fk/530S/Tl6MX7w4QwR2YT8VK
22Mmwfckf7BkEpUNu+cU2uWtMknT2g20R6g+nRHiJraaWq/hP0E6s8bgw816lybTgPWvArG76OOT
W04p7x8i1bFKIGqqwwFBDMsHvayBscuqec6TWasaz0RPB+c0BPBgVV5/uPx+0WKaUXcecEdMynCE
1UJxCDqlfupARj5AdU1GQNic3gYaBu+iRDe+WsyJEEXoh4I7B2HwAn7ezRDFSuePL5Fj5v/1vPYO
DvFPM/J5bRHqbviJgVt5PhSuUDc1unJSq3vHOq3VO1CbAe/S8A0UUDE2vRrqu7JmRwe/cKW95bJi
hmdX1ggnbfdYsYDP6GhUOkw6+jmnp/BwW0i43JK2UwTylZdFQYE/JezsozEuiJoQJ6kOl3P6yWaB
/CqhwrGyou3ORM54r3F0dpJ31Ayoko4n2MtRRowOuDl3qdjyBqL6MCltqQQ2N+DOu2UfB5x4I/sS
K7WMUMPFq6wXY9YfTwrBODBhOp3Yxw+hoNzQpGwLroHK+Z1n7OsHmoMID1jfRotuDB5CdnkcYJLy
vgnHpkB2RYnG5OHthL4E+ftsGS2OCp06vtSq1YVc1Qd+jPSaDJcEcGlaioEbQrOLkrF+hXJgQc/B
qJ7eKBo5SN9kj16uxAJxDVB0h8X7VdOs0EsYJVdflNLF3LGflX03XUDwDWCe0ii/ZTPX8LgXEukF
GLe2PRE6nnQGElWB2ocvBTFnWGhALfHN+qHP0HoBR9MPqKcyWdZdIY1SAppqBfEwqTqnVrkewaHV
xKilOmUhBeVtVipYEmQ6iQEgWvLshg2RbTmnmoJdMoPlJXud/hI6Bnf/Ftn5UG9HpSizLyfK5M7x
rnwnA4UFIsLq4TvrldHu6rpGkPOtHt7T6jV3iJYkZrTrs1jBAnQiBnLCkD0csoXcOZYJMNu/ASSE
8xjCVqSNu/nJY09Pqj+MRX8BJk5Hqavv9UtEKnFgosIP/L3WGWv6z03DVSMc/My5hpn5FmpjVJXX
gCuIE6rpNaQBINRJZSwwJil6QZyYIwZwLqtOBsuk0EYEMv+MMNz62VLNDrRAR6ZpoJ+2ECLeVF/U
LdGxNFUmQUMYWF3J2V6P8t2kNbwqyhrWmrgogXx/hR0a+KIhd7g5F/nxPjh5L7vMbpRM3gYmY4D2
d5z+Al9SPq1BlIW14wc5w6Vyg+RiT2fpe/RKTMFtPszwhZc1FPPXHTvnjtSHpL83een6//EGWSNg
614eQgbW1OZ4BFgkx46nwFcy10rldPQvEfzpS0xX3yA0ijGHOWRw9KG07m6u+ZU9kBywa1FkeO9A
f23u3jIhYOjMqgD1oh+sWff2pvFPpVVvs0O/Om7BDCJUEEEhBI2ZD6388x7kGYCJfyTAf3fi9Ku+
LCtPjXobYwIFru3QeuoulfIQ21ivdWgOWadB/Yth12YntYJACGd7aIulOZtPPGjugjlWxgXD1xM1
efo5aU8o9OsMo9K3X3gh7ZBHEN/NCqqiXEHKNbHuMOQcQpTLFPs5L23Nd4Xj8PrMnK1ng5CnzAlI
x8EdumWlRsn9q/vQM0VJiW/RZzN4cmJ/BmznBWeDrZnk/a8y68U8DgnMYfVGXkXoT2b9cF6JHfnN
k3sNe89AbOq2tAK0uurXk2ua9SdwN43J4VqTk/bZYaF5rK+qwQnx+fdQQaMLy2JJrzFiX/WtiriG
V0LWSo2iluhfiMYfP6AlZWXPRQaPF/cXs9r+JzFq4JVo8kvl0KKTtSf8A7vuIPKQoKUerBD0xFqP
YAPeT2NGFlDoYA1dhftYMbdryJKT2HfZD7IDiAZyYf9BaJmY3OJ2Nxu6N1BGNglyDF82OjdK1/5e
5C7/HFSD/YXZGtPpz3qKnotVZEL0kk5aL27PHxZxcN807LPA1MOkztgnY1fscU7l61eU7R0SLp9r
r4A3zoYc3aQPGCBDI1/ldfUljiIRwtNnaw+gQ8WRiUqQYMtn/OjStR4ViDk//agetx2dY4k34cWW
26+SJTQ/y6LHSq6o+CgNP3QIw4u1/cgaPwJF+lhgk9Xe6nQmv/mEDQT7nGH73uWU/pP5PoxgNR59
r9keqkZfrAyTozzAt1SuwWTsrNmk4ysG/PxFmsgjKUT198u/vnyU9h3/EuQDlyStP2Da5oogUeEf
R1ai6qUF5veCgrSyOUQxlOdpvf8xmWU06pjVVJ6oAhz74ZFpwRwwFIkYhEw0YTWINHh9cBO8CgH6
EMk9OXkM0sbJijGMx9prqIA5CpEmKERxxMdMDChynEyCmK8fMIdeJAtqAfzfue6lBF3BHIgG643e
Hln4FMeMVlfXyIxgVlpau+Z7rZIThnngULb33RPM6keZXU7HEOOQ96zosx7EcgultON2TK4eOImL
J0kmKGzJSXd4i3399lor//r9Y/tf9ZBmxzQf9zaKjx0jN79LEjeBVx+i2Gc13n1ZArtnHOERk0A7
T6Hkcaa8hkYbNJ77tXkFYxzb4crpX0DCoFqYgLd8oVRUlYU31poK37IsaMQsvHpq/3PvqvFgmQ63
ClI/ESFhIJNRZaG8Q/y/GfIumeW0BwB3+zfsYVOUZW6xq1bhZvy620Ngi0QJllGxxg42MOPn8nLD
3JhqUhPEAHp7fiX2zXKz5bfpe859/IYldmv/Nn/hjebcqfr0r13W7wIOxpoev4DARDzICt1PezSW
bqP70EXp97NGqLE61FMiAOr9BQt/qgTE7ZFVxlS0DSFq5xrMEtBLRwwfjKVAOaq2SN/0FGjxwJDL
PMU1GjVG72ndwCAYqI0NMNh8ccvhaPV4GD4VpnjKq/uZf/UQ/UenNAynK7EsjQe3aqYxM+TxxxNl
sMzB7+ApnOqE4uDesPFFUrmh+2jb+WMSO79nLtYAMQ5vn+ajUl3NsITJSZygrKZKA1VVVMmNklia
+S1A3ZwBabyp3eGAshUrJ19GK/SGVIEWtDlWsgm67lx6XJJAJ3/8synGhk5i+f9R8CkiTQXTS1jL
B9NcTkQMlq3Uylj/BiQbcmh4GkhBATSZxntzCtwARKKH9X3PHL/Zwp0E/83fqxEuX2lJEYVFk1a6
7TOCJgMTDVw3rAU0kYXFVzI0eWkPM2CNV2JdS4tYmlVhKLzM7Fw1Y8mfqPQoCX9XTPsDOBr/vaNU
3tw2nliFmpgKU73GMvylL0+lUmbUuU9rm0/L1lEAdUR1mTGIvKg96nPNkPKVqWibxRS+F7li10sh
urR5UpCP3ozshMAewFjO3O3/qWNMNw7YItcQxiYGjjQVf3BqQtxC+negUmHPAC588HoFj40OZK8t
IlAs0aTmwOdtfpWtWKOeTnnsJGQXW41qkpIrk0rNLxrnKjK3+AFOpO3oMV1Rw/dKX1wSEChRyEnT
h05chd1C3Sq7nFlDNC0p/XXupS8eFsukZY4ivmKPYs0FTUsN3c3iabE8XLBBanYgWsdUAlY9j2m7
de9hz/ggjdrs0Dc4dVNZh1IENanyI5qesi5v7JoajAGKsJEVOgAtUok2zXqMIp18HRQ7nCb8BKlt
Fr2IEpd7bqz0/mndJenNbmffJ73HYeQj5syiI/xmv5isnO6XIrP14Fkae7rcvw5bXJ8O671ydNiO
vwtahk7wOuoXxmPsmT/KIpB9A1pEpzSjoBVq9LCht/hfCEzx0mIZvHUS9EgUI2sm2BdSEeutT7JV
d69N4ytf6qiM2QUn8jZtt/RKqjF/FMoZ4HWsv38YT4iEiKmpKujgQrNKo5Hc9qvjcwiq02AVuGGL
3SepMcb7EeTgFiiZYnZoe3zXLbN2n017aJltUvY0eTqWUNoOOf41h69B4lcQHNZAujz2SIbxZ/oM
RItlPDc3QRJQLy0P71TodUJebYuBx1FPJWLBi0YN6lUBJYV5xIYgK5EVMiQVj7AMESSjGLY4WZQG
yf0WidPZFPVKj9BjWjy5Uljf3cBltUqyoeVnkxn/yb0W4ntsYCFA8aymICat1wwn6AZpYFzq1Ogj
Th2YkNThtEuEfQ3x6LDUrui+0I9QUkSW0C4TTSQSU9WMnrLkUsfn6VbaHxRln4nH+WxxbPh1zEi/
yD+sZOUXnLqh4UO7B8EEqu+h8JhzLJmdRQXahPoNmcteNnacz6fvtBRvHUCatDgLsflwkozZR9YX
CwxByjHGaIUJRaZQZwBNZfqAf08YbG0y8xbXrBfIfAkuvC5ehYvTkXcabJy+Gi5M52YxQ+/a/DMt
WdHUkthsWOlIWJTJ1m6C+/RJ2g2b34P3rqVqXUe2FuMNaTSxGQiv3LgCbY/yOfRf283zYi5iYjum
O9/yvXpXGaPwJBW3v9S/PkDwdcFsTWuCvZ7/yq50xi/Ym51amXUiAVLAYarfngL0aAD+MZpeek62
h92Ab2R+wJrTxTN1sVCBSvpLrKobj1zT02upj6/TIyhkonxXld60hzlgdsNk6uM154dlpxbNzSZS
5qrwsYD8hRmiTzFexUC3n6SpLBIL/uuKoyNGmDxg1SGj/rERzmRhLF44f0Xx8xiLuMKMP69nocsn
q21ELqktT96a24+D6md0WPEKwsluF/IJmE/uMmf9s/DV+y8CUm8bf16UDnXrAyku3FHU3BQMk7PV
bMj167nIsrnBEFZFNapXpauP1qXXfeEvJx6/ao3mw1vI5XhC0Bp4yjgrpGP1PMaS+INWNrB4BQkX
9H8LCfk+NWHGbtTKsqI3etAH8a7Yhu69ggjjpcWXmCUdjZSI1bvyLo+HDvFEWfLtREX4fYa+6H/I
9/6cRofLPlgvFyz7oEaCHeFvrdO1VF2buFzfqnWbq6ijveKioU6Dac3HD64yBWldNwBju/Bvf41u
HyOwqtuTVtFW9OfHxlL9Qku4oq1QP+RbTp+twV25dP+2z3H6bZZL82u4tGFDlpS1+zjmCyO3kz2O
nExAt2UVCe/YIJYJMdXkEHdp+HxGk8XTWGjT59MIEA1u3HznPiFBM0Lvkq/TwoVyZwUCsiAhsaNU
fnoqDmzEYBCDUihO63b70/OUwFguJGIr2kxPBQIGm4+d4blIWm/ru0/rSHs8xtz75mOKQzpPjTt8
CwXO7AcwfEde/sWPtLvqhPTgxTR9TWTWBAOpVWSz1HNEnsIvfCv3y4XEH5u3LpaLw8V/fZo1Y3GI
A29/SCngZ+DRln3BL9Th90fitkvYGaK9tHDxax2KlMPgkv+GF+JWEHj0K8t5YuPCB3uB1KMiqOc9
sapdHXVBmR90O/QYA6wg5aZqkgwoGxvDAJLd/w1tnJYbCVnExONg+/2zHSyRjTVnK+eIDF+Fk0w/
44RxScBzseu0n9Ta205rXqi/HgGsGrIRjEsvq5eBBy44nrw5MY8K9UqwuQix6550wwUA0DbG9+AE
cZrYxJFp46sYtBUuG6vrkS64JCi/DL0b1/DDmF2PouySlaCUvafKMqMHit9PpYfctJTjR2kKX3a3
Ml2/KRCU7+dAHG4s4ogX3NsIh6kLiSffDBuQx10iqgVglQv0b2+4PH5D7CB/5Pza7pDv0XJRRMtV
r7A2nHGvir0WcL8q4uBY0i+Huhe2fQcPFdTTUTjAOfAEnrO+lTDCNnPZnmgR2KLk1/x4CXmPDKU0
03eaacN1dgP2URwobEkFlt6X7EZB47EO3CC6KpO66QGLB2QyWsJ4N06evWiZoX9h/6G72Ll29oDm
/XmW4mHtJY22dZxjnYEUUcp+eT/GD3+taPgMA8uamQ7jU3BerOy1NIDdRnKHyE3ecj158lIK8FGN
mr3f3KiIODlpKG2Aw6BrcKOjS2s3F95r3QScn3ViXd2qEIuLrtWrA2Ag9Vd5LogEZZ9AAB966gV4
iCCXoetdlj+uiC9GG9pLZvnuxRSCFMgsN+H8/huA6ZYEZLHku5z+lxKETyDoAYQweJOJc8ESLTrQ
2FOMzZXaQdEMbFVU4pHx7bRUj8nbPoh4e4DL60KM51VxSuAO8NGlTAkyU2daHdup9Iqhq8TYxTOv
fRcH4t1Zo2WVa18tWBOmSJ45Awf6CQDfubUkXOkoj3UlniELfhetoJy7mc4mpGbuYUj86Hh2uURe
pXKYTFDUvYRQkrVZjWmldT1Wor63xpMQXZDuCS7SVSmX59k6hoxfOXuxBKrTh6/TDtN5Y/UKvye/
OXk8O7BZqHwED6e9jpREOATx3IpbwcCiHk2uTA+mf3YZEmtYB9oqFokMQU5irKsaoHL+Bwv1ILS8
96kqMuCibQkM5B0Nktsn6YmLJIgAuOs9k487+O0pX+7Yrtv/A2XLTiwa+gl6P1KDuSO/QRT+gyxa
0WEflCCf1E02QlLHwJ5wjo+22MTC9tCqxvdNbDPydPGa6bBrm1g5E39I9pcNC01NB3/2zvpRMnBO
cyCDplEImgeMFp/e7LU+/hz9bYhc4J0rrY7dOQUQ60Tw/AH2ZSQsnc4Qmd4amKY7ErYOJ74M94Ox
QvCOf9xW3owxCF/sT0y20lXsn/kFhpoySsxpETLo6mwiWGSOXHZ+6Q0XUY6/vIgcbcDT5mOnqSa1
5c51a6nGpnpkSzIp3Q64hN/8icitoxO5BBWyhR4bACUHO7JxP4Xq6KohC1JJqwEH1CPZA4GZQUeK
ixjZ/XdGKFW2CZl4/hq5i33HfA2uIlkhgVKDfJbWYrR2ntsUSn9L5KSbUCVRXeEUCw18X9ZMWgnK
/eOgv+GYwYvAed9KK1whbFpg6CX5qONDL4PYulV4MSmjMVl7pYNtwZM0JTNK0/LfhB5FahZ9cdmj
uqay2AR6NX544nG/+Phr3NLl1iUnwG8jKt8+3IPbJRy3fdLrqp66SYq+8lKt+Dx2eyJMP/9fhpbS
QLsb0A8YF/OnnhiZShHjk8DHYW1Fm+nEHbdhhVJy+CrSZSuRh26KVMLCz/gaZLzkI9Bp2Iq5tYjt
LNpnIxI/v1KF6XgqdhelBXkUxRQDkQspXtia/xOXBqO0nujr60I7JUx4GwwH1Cb+xntzYYwC8n2R
aCtIRZ+wtYgFjC/zOCNVDBjU3zkHDe4GYxSu1xq6oS9quyPk8tz7ddx8WRVOHN9HCagxxmdX182V
FghLrLuu0+rYA9ECHZpN0JZZzz7JVwrZ6/sv/yLbcThqJZPxgj96qDYUpEBT/pyEBhsRoUwzlR5c
b8YueKiTl63TmDCGSaC4Nt9Z++9icqq+UHqzLBLPGksps0nGRISZVQShmBltVxrWpBGjnu03Z8+X
939LQfZgxR5ehIEn9zZ0tMvuhd9JOPXwYANpmBkjELhmy40/n4JFpKK2njvPmADqleQqY+cOpHuQ
D5SwSxplo2mLkIVEPb+Qaj8uJhK3g2cOcEJeoIuBCxxXkeyexN31NTtQfrp3t3zP8YKDr9SNfOiW
qkArOY/PsFuNaa0ewKddb7zggdCmuNfb16ViP1hP1rM9phcE2a/4rA/lKtSdzquWw0Dwb/X0ErG2
OQghajxkkCGKWmdrZdW/h6QxGqK85WTUnJZzQhj7XnnJemC2BD2UdQFSAx+NN2BJu7sG8VrR7VdB
SeTzgobINYrL6Ei/ofF7cat6zFKtsSg2/sSsMlqnkFvNirv0qRUjac6I0sansUGIT/A+vBvTQWcA
oeUeRianyfCe8hx/D5fEUdaUl+qXlb2SvQZNvMRdZuxsG9h4FHUrXyXNWmajgFoUwvGXr7K1ZiWH
/oea1csKS3k9dXHvrsJ7eveRnJIm8rTD+KJDXnajCnqjHf71ss+61SkGT4UG+gIugTyNwFM3/XOs
AfBgptv5Tzf7z3sKzhoMF29rJflQYFIbK/H76Mcyuvr1HEO0vZAl8x4G3FtPTnSR8DRuFANBohhj
koVAdLNHXpoG4MzIw+7I6FQv9VOUrdhAnHml1WZmgQtYICMhZ+9JFuwE970X3MZ4TcuKqK5TSWl0
WEwfzetfGPRb1yIoU10ilF2uOa0bzW8Dxvb5hbbRXxMKK1szNzrvJieFY+oov90GE5URf3ErulsX
pfWHPuShjU7jF62k4mIplZGDiUIlVuCfDswYST8KHkyDVveJ0RW/q2v/Sv5vtUtWupkaaF59OxRD
b5J1KOQP8GWbD34CL2UHoKgZwU/ABdCcLPgMi6vIL3hQ8cuwGIGcWODe4l8MmgpkB724mTpXsTeD
n9rb8jWlFIV85m0qkfTHX7NEDXoqzF6MT1EDGj+R9OZ/2Bno3t6WjIqyU8OR/d5TGkycWZISKnHG
FPO8ufZEtvXUVo2d1zmTXKsbdu90d3l9hhB/g6Q+G6ShC1754nU6T0KQb8nMNVIZwKOJ0D+ZnYdD
6Wql6DDshce86Z/QxFhvkPeI+cnCFnF0c2tU6sShZ6ubVldClGWPy/+l2jImJYj5eKivUtqh+xIj
KNSv2zfOEVRE75GPu71QLLh3UmGmYlDLusPBFG4z4Y3mWtGES0vA79qFoC8Mi5qOUBchRzS8l0Kf
yWwzMhMJbFWOklYw9Mb05wHmqfubh+Tmlste9DxgAuXOClawlq7exInfVezYiB5X85N1fe8NDL48
VtOwLZQtTmFOdOmcHu/xe17foacaH3ts5XXRR0uHedOgZjjqS+OfuH6qFgYHMnzdl9C7URaSfOWG
ueE5sOjapFBF6CHK0KKGnd8WTfm6Ew2oVR3r7Br1zbJolkIEBmzgngFV/wSsW/uB6aSHvTJIuloY
kZDxSwNwZKU2Dz1IQPV0/ty8QcBv0FvpWWdb3JLMXEDwB16Fog6gpwBElZK+Evd2hhgEIV4+cQhH
nDVBxNEwPqxUjdJ4lfoddQfNuWSxJPB+yHn43BKEReKdKhNFRphl+XHxl1D2MGO3oiNLLAO9lMSl
lyKNTaY4wjDvAuqFO1RekVP3Pu+wcsb7YYr9IGB6QYOh1APD+KIflClEjwPDDkP8PBLINGOKrqv+
9QC9JpzShUTLYp1fbIZMsTNNVSExXHE3uJ9q2RJpDDB/aAjhkCA6+ifLlovlufgt+om8oABnURFA
2S6Dyei5JH/B4mDHK4p+nHXjK98oKHl53gE8cRoQfEYaQRkIo1U8ns8HH4HHrnjWq5B/xFYIhYFE
pzPz5Yk93WNAZYhlwM6Lujp3yfnyQ181O2cdT2CEV2O2R7Yhw27slRT65rVoXiAfUetXyhyT1Xpr
25EDH/ZQlAk+C0FCGpH6/+DnvRVCbL8HhcPGefx+PUq8oRBVg4NA1oTz74IoEwzpAPoKFDYUcTzC
OpuuZDvvAAEK2CcGFCzVhomWCOy2U9i2X0eVQpCIOHLFRo9df+sEwnZSlrYEjxDCwsBB9BYHX9JT
uN8P91g58gNQhANCVgUrsu4pa6aNgY5qMMKZCRgZtyZqdm0DwwL5tPem4zx19WCVKv1GK9O3fUO3
7qjhkpGO92wBMXOFEUQsOZ6aqHd+Ki6AKebKaH4WO8DjYyQMcURt10T9t7yO/ugfh+CBmRbb4IGY
TQJ569yoYePgqpSaHNSeU56vmywEZGcygNTPxpYSO5kRYqO5P1e0U38w0htFuJq6E6P4UkhwO5U6
zoRRSsyiiqA6H84aOcdIZBir0ECX96SN4YLlgamAKbpeMpQfum4r2ZWQbQNVpMLyiFQQljqppcp+
6Umma2m9qr05gJeQHOazlPeljazG2tpoTREGPFRqEo9T06WEJU0aQFSJyycdcrtzjdvWQSO5otKo
V3aEvNk/H4u+6LTdB26n781ggu2rCcOJe8bznoKFyCp4vgSM1jxnyEeNswcEJLlfZg3LuA+DO+Iy
TitzznJ0P54tBF6Le9V9ITiGg/Kh9vE8bpQo9wG8a3YO3WvhkIvwVecnq/lciuhvPYC/MnYa/2XS
am2S05I37qaWgsXXCepegFejabYEQSFGNiDWyMJdQNS3uDTRTONKYkv8t7UzTB9lnfHdf31FaAAR
50z5pVrN8wBV+TgTuMaiYTUIhICTM2eySfIgI6qGEJ1gFrWhWFYrau0wa8lzT0h1vLSK4y2WVPXt
79n9JfNMfY700/4elk2tXWQbHPQnSiv00jJHmui9cJc3e8Zlpqp05hOl7v4ABrJG4euGizu3puci
7mfkkVuc0Fn04yYDHRnJsLRI8R4ssXZW/4QAbYvSFqaVSLlYIvJxlakHc1URAsy/e4mfPFwsPKs3
p0zsVwdQjN0BdF7n1YJI7U6h1fmBAUSRpDiQQOnKkJFxU+FRf5Ajikv+BJtLKFM95eJ3kpfkEmAX
50dZbyvyozqqHPZCOw+1hYnQ3M9GJymiVnSni6n3sfmqQ+2Ddj0eGLWTJxANyqzCqRuQB5PH2L4b
JWkbXN6ctNrxYGrtB7h35Snr3ndmNAk4cQy17X0LnNf6V2+pgIPKVS7G7ygIWWW7k1aqky9CIwty
MXk2DMBoyvcsmOuDt0qu1OecpX7RlPoGUhnnnGOsmO3R696ZDhkV5hLrkCi2wxQNM4Z8Mc94nsO1
egFMGMyONKQYrHowT1ajtNH00vI+kkhXWfOKM94Gkf7KmQTgeJIADwP9Omfm7WyF6vg3erVlEqXm
UoXLqc4hvB4TqEFk3qozkV6CSE1OxISmrFdOU+mmwAOz4Zp9XAr8wWIqA91bXGUnrIlHnxECsiJg
L8wcfbRJlxavCoBmbxVAzPmF4LcdTypg2lrfxLKjOqR1pNoxMaKOl5sFOKOIIkFi3kO+ND7Ktw6j
4x1OFVHhT+pqrm6EA+isvS8Lovr5NBbHu0eBMiCDRSkSnYR0qaCORXL6zgnrtMXndUHOAJ4be1Vr
SYyoXq/+YC5+4p+PE30tqsKnXshNC25IgCzjnKIq9dhLVROh+xYMwcZjXz1WM3Nxzp+ANRLITt0w
A5jajOh3Yfmie4YsC50bdVeZHRii89QHRV3yVgUONNJUhQDzqrkwxyJMLT6SETYKsY6gUal5rHcB
hzgLoH/RNJJ2ERY7U/uj8UzHNvseiqnxjCsxHt8lu6JQKsSxE4+OV7F5hojrRqAulz4g2poGTai9
TY3XPV1bV/1LERyt+OHu//6/Tc4DGvbFCID3sQpQmx1Tw12dIznvaYiFSIlJkHN/P8Qtw36J/Y6+
EAwc5gqEIlcIeqF5eyUi8391/RoSYluYGn37y/g/+FjZtRTjWgppgAroDycB+83rEXLroKHOKmBG
nIRwsmvWpOyuwFn5kH5LhJZbVUrhqw5qE896fsWLrM/lK2T3vVH805jzDFszCRlnu6zjXjBCzg8F
qts9iWu3vZH7/+ufOlDnKJ265xaVLc89api4D6REJfo6YGqJB1w8WCi1eKSr58NXFfD2gvJyVPug
fKDjX4NSyWvMhfAir2Qv+1XsMVXXPRAEM5VMQ4H3kdMgKnj7Xz9Q4H0HDsTXeJjLMNfbuV0PV6h5
r3Gt+Qoi+nz5zvLdmTG7aQUeeUzq390I825exD4m+JcygkZ5XeMbE1aAdcV9KHNB+TYiIs7m5Xdz
+BkhHMdEILuvczUBWThWHiDg3r1NxNQBil0SR11Kj/YQJBWGyiiqpfN0bXNv91wUGTbeKFMv4wmg
PdJ2iLls/p+dzyAA1cLl7jSVF1Ca8nK25DvXv3c4a9qVjvfuumgXRgWkANS/v+KzRzkeAPYN+0Z4
EN17zZHRNbV3wnKbb8Kkveq/cTplbFeFdeZglpoVuiJ3mQl2GV7CbfsEUNtVqPl1dCtLYpzNJ2kz
/fI4kYoXUmRbk8YjuUAq5dme2a4APuLzjJtP9bQUajmJsKT8xhhjmLpoFzJ3E1rcoF2tkTriw2cO
UeC+LBOWk7MEAm5ZB2LNlhnvMa17jNGphFDaDhNkwjx6L7bxK+zsUn6BZ6S13fRsu768+9m/INlM
mp9jTUDQIdlToJ1r+ioj37OESMNTYt21PeeQgc8Qo8eHyXrzZH4NU5pZO5OJV2vPjnzmHTzh3a0k
RP725AU4LEWD0kmu0ie2gd4Lufuc8MBhf19Zz/pAJUxc2PO9l+O83P0WWeMP6hFpTFzSfABK2/F0
atgdZY52+bDbvjkHnkvtndb0THrQt8oVaCcUSzTpkhfyXopBurLGXVodrJKHwftQCsxaOUMLdVlX
IjZRU3Qfoa29KGNqEfSFuNwuC3bjrhgmaw4ht8w+oxR4iWYW0Ge8MWvXOqqPmwx/SRe73+CtxOgs
EgRkQXdByZPp5bWZl+0ZlpR8xyccAWxMic9ovEEkXxZGZXhwk1RgkzqzkgKFcNBXodhVjanb5j/Q
Txrkm9K0hbQPfL/5prrkWuPOIgqiAecK/nkNmeg53bpmsODJAgAjDJ0y7iKtk8MwsJA0S4Jx5iQy
py7L2Bm+FIxg5lWdRnv3rVonYmo3i6bTcXQOCxUm+Z9GdcsCRh5c825I+mqyfdF/3JJmHbUvayER
b5u0rZJPPvcHx/MVbdUbekZGSjlRudR/09gC96fjmWSH3H3w9bIWAZbxzgCSCXveUfJIXkUAURm3
A0aqtu/UAChDc+zLckTROU8GSe6E08+tINkFjd2cm0hOzlh1qyeGDFt+CBGAXgS7U/TfdjCAfudE
7Qw9yvicASLWOU8tyUfbhHsVAIh6YchJmJzOiQ7qgo44umIhXLoS3MHbTv406Q+AlidxlAk3y0am
nZ049Mxq/Kquj2bye8l94Vxt/XlPbjsFKIv60hMAqJJd9jDpL0O2dJi/KlUESrfFfdch88HI27Yf
O6ar/vY4q9Qn4dy3JS6LraRYDMfqbYHnS2/8UdKO7oqfGF/nbCnMPyJB6E8bMwXsqTqO9j28OmVq
X+aJL7gTRZSdhTP5XU0Kna2vzC0itMqj9lBON9XdUV3rCa0wduvXMxKsTnn8Dx39JRoDwSwsA/mw
sGUJ90WFUFf2LEAj72qbOjLHpO9qD4ivKgy88Jx95OEpbuhzZwUOaSFi+ox5k7D8JlySpAdIBbAl
U/lXLoO8NPoQW2ssqoH7er80BrSRG/Wwn8xHqyttW7UYPv7bMVoqAO+Yuiv3TGlxWSkh4q4BUlkR
KTHmpKs+COYCvwDWfwk/9DF5qaSEB77jlzBuJArAKYhBLNuEOcRJruU8RrhcuBsU0J8k4ZLk/bGb
M0kYp0lw0C5g0olRdKIl4RRuIsnu4hQgi0PoxVkPTNMXGTIq/5uno+Se6a/8J/XhH6s17LV2D0FF
eOKj05pSzkH+WKMNRR14rSDHQZDtpa+B45GkwfsiL4n8bmli1cOWGj32I/mjJlDs9Smp8gn2kC2i
Betc9mkVEtgXk2YR/faSLtzH/3UBT69pqCgVj5fB7Blw9Lz9hz/rizNSQUfWiz4+dJkDhQNsnN3R
k8J2krN3Tle4J43sZJFATGRUleXhx+gYRUpQKu6p5eiWlPievIc9yIg6TtEKhB0gqJ/bI+KjlfRG
ajHRlwSs1V46ZaDzfRtyOCNehO60Q2UkZ98zLsJenHyOBTRWb1idHzDlpJjkVyoqv9KxThOj/OvT
Ae4YUNdlgrF6ZpWcEXNkP9aLuALg9rrkvGoVOCP7c6FMLBQdgce2kHW9DZ55q1zeMP2WU2rTTbVF
M/a9bZPL8QvCvNfME9CCGPtB8AbONgxZOZFuMylT9NxgbNFXvJK9ISdnB7a+oVDWuHXb2hbcX8AF
7CXXKvLfWfggP9Vl8KUnyWvGDGSRrYdX+NXeB92KW2iTxmsqZssZUADbJASAyMfLMQypUje1/4QJ
CC+p3Vv+spZvJ+MaZOmpnyMrnMaYDwsx7/q1ZxpFi1P2SOBzYFIBiiL3bMM2GRASqiKoJzvFOrOk
x7W9FARP+L4Y+9sASvUIrTIZDhs5TEmWrNSYHv5mLxZsCZGJjRRoZLmuZb9izyWkHWwJP+9kDd6F
p+QLPk054NjeGYYd/7EzYoQ2khLSXKgG7EvPhgzRT0rDI1Rq/3MBAGtKlT65jMZzUGpM6Vn7vkrL
J4OHXZp/mJGeiPSeAt8JAa3WLZ1xlwmUVzf9QchM2MwAGlF5mEk+qv+0emZJ+OThe0hLcqZh2vN7
y8otlAs5AtAzgnlIQGola45LJtbVE+9REH5j4Cs8KbDPsDsKmavWkbtu61qcyfa1TocDyDwjIpKe
0WGRJB4bBM5KnLNCfFQ2iSob8X9embJWHHvE2J79VFRnW2gbCnnWX2IP8XnjNHKeOVKqra1dA8V4
VJwvqyXpBQdJMdvFK9sX+G0NpLfUOn5OeswTQCgQdOUnmKS+SbYc0+R6CH1HxbV48EAincsqWlEX
mp5DFT/dPQa+WH/u8IcPaA5D+4dGEzeFLfdbPq9KBayvxftKp/PCITyhE5XsH4cMPCa86BR9LRKJ
U64w/MoINlYlig6AUNkGnwZllcvWCyGr5ZsIIvRNjbIQ2qb6zcz6Xzmv3/B+QIeaATvJF8qvWD7h
DsaNFtHB7/cbRMymbqqMZ+t7JXWQC4lYyvjdnF0VyD5FfmgqmwzDu5tEFdMuUYfNQUluPXrDGfzW
DjgKzpYErDxRpgffh9QZCiySs3B4JtDWHgg44X3XMXvVOoCZt2ujZH2A9gjBSIq5UexDgjYzH3c9
fCBXf6SkeSvu7G5C7ZDAr16y+o2tTYKBs3VrV79LoKgGeAXGk9JeF0wNadjkSes0n9gcZhtVYLmj
nrh5SN6ZLVMAXtKRvwrbjrX7A4ovOId5gcaVrMxHpJEOBJqBX/AKEPXuz6ezmiIU2yr2/+1jbkI/
LCooRkL3YcYlvQmTVZpMNl7pf3MGoqRLjpOef8NBjtpKjuVOX16GvKHIBAXiSohPSl5iml1mevd4
AarQlSQ+MUIBg2DzOVj06HbU2AAQ1FNsrXy4vdzYGPzvX+VkMGD/qvlmmuitDbUsOyL5Xh8zUpGi
/VEERPORqs8nEmoamvoOhC3lHOkt7gCpqm7p0tva5UcsnB4CzOdyH6CJXrw+xnMf0Vire6Ei2j9u
bPwdzukVFIYJJk2QW6NAWm70gHooK1PrFfBrVqOQljYP7ULTxrzZe+aE0h9Fwbjs/BMQY3dXQxpu
pp9UE65qqhlgOazECqPwizE5x02aW8sRISUhzrvsg2vay38qqSD3Ndx3BL8wG+FEqy2BLRGinyRh
bzCJ04V/NZKeSZDF1qo2qG+41JDEyXknQbVqq2Env1YOe5HbhV76uaY8IHeMjdg11bl15qI/H0ps
CnVtUb0uY7PG49nI4PTt6lAJkXGfHOd5Yl6WRx9VxmwogsZBqHklj2mV3nmyw4hD/UmFElzUBZ3z
V0mU4LTYF2qjwPWT/IRsk3DPT3Imrs93ewJW4E5I4wWQSKOQkzwuO3+WowBRK9S3/7VwYcurF0z3
W7vbG/Z/Rh35G85Je9o+OOpE+qzQnmIGRskb8XURhXs4XkGtvNzjjTncebzyCrTZ9ceQxJ5IFcrA
h0H38EitO8Bp2YYZ1naOn44XoXezFSyQzm/j/FYiMViHvz77rp0oi2tUIRaYcJyy9m3+XSUxqgSZ
56dmv51EaFXbffZl3xSPMe+MyNwOTh0aIzuOddwuKf0RbcOyUYj4V34UYa31HekXg4hd2xVQQatq
RPtdd00/rn2Y/nb4dvqubUSIddiXdGc8yte4w4nSede1i7Os57fU2ug5vRnCwKp6y+426zyMbFcE
BY0LnnOo+N1yHziJfbIKLzTsJ2Q+B1WJRmCtUj7JbBMWTm058qnFQDFFqO4ECi0uocjQruq0smDM
O6gceuTOxqB2C6x5IbN3a4eazWn2el6xoHtjBgTWlApN/MKMimxxhzx6KxPEGgxu8lxwbHMbNWLa
yyyGFJ6ntHvpb8+rrUovugfu2X8Av+23Z8Mq3lSi4y4/KYxiIOLxbxvvb7uKJVvmABsyiQTKuQqv
PC/R9Jl2MVxI6/D16tpFhNnrOzN3gV+BwObkj1aO+ypya/C20O48ZrwNj2PkNHPTdgEae2+lz5Gq
+Xb5UDQ8OQ3K3w2UMBYebQpi0wm8WpQ2l34tLEk6OZVvF9oyGdm7dJzCB5U0iAeWZ8b2Lei8F9Xz
1uGPDlkyAs/deG4Pu7eagGqAb2ViN2uKbP6nM3bLStoyxgmnkuGmTk3NpvaZ1Qy62xzkALYWJQVh
EPNZQFDCk1uXWzXsFx720ImdzaXz413ZOGZlLupxCBJIJ+dwH5bs9kRzI2BKR01z1gr8zHXAMg3F
F4M+bY1fuSTQVRw2ZtPcmzs4kbbcN5M1HYYeVv4zx+UsQMuveIKO2biFuPh6iu9TJK20TFJ5rykC
lSlFl9Mr/6TWWkOAu0WDW5FiJ7qL/lrIypV9jfna6DeQNV3oGVnvlX7Ijlw27QqDRUKHnXHDMOE8
wo3xXfbVDa2KrA3pegyfoQSs2v4cSR8z5Utqr9AexqHY8agBZOAYNeUIKC7k4t86JI+4Zbv/wzt7
zWSxjXhsiAiz+0fVvKhdzM/+JPZ6JFxb7Y4xTz1a5ynwx/aeyI7xrdoZFK4Lplvt6tr/DV1Lx4h1
IDQIh4b7E/hE7ZYJar5C+pUoaPWTFnkPZUsHlHLsQUsiZQavmdXcuv3BgqztbC+2WRsebNKNoSKH
+Iej+kP381UMGfqzwvIRzmXyR8z36ZidNgNY5Ng5kSGl9BN+FeVczpoIhGJWnXPbtcwDX36dY5zS
quuk/TIo+1gyC2smFm34aRohOheSmaR4tQPNsNrQU6DUomwscm4AyMouLk3G60oCldRZSACb1kVa
Ckt+XnG6knJtk5h/2lhOed/sZbtlbzXwjtgbx0Af8mpqEJmFTQJF3pHkvxVBaeOpMgYnQCwWvDjZ
DRMp1CGA58kSU4Ro7XTj3wLMhCU87eDbL6ljFxKsjS1I18tLgTuuaudFgjgAk/4/QfPBuBw7+for
lnqT/R/2s85/acZqE6rjWVMja9lrIhe6JRAbnF+DBdWTYqC12Tp+4kkDjOlfMssvhNfmdDzPeBij
EKOzfMIDSDK9t8+xMJ/cLaIM3HXxEQ/yoaV1Y0fsSR7KDXgHCpiETwHicTRpvlc4KOe588ZYTJH6
kObWvc0LpFIvDIW1vr2fvUT86fnIWsG0CTaX4C1XcxjCl5S4JRNMli9qtg/6Lnu25hroPkYWzNiI
lFi4kfr58z74u0x/OVErC0/F0SGENAoOa42Re9jt581PC8658Bx+/TOOBCMN9v7sLF78UL6ZM2NZ
ac8h586Us+G2ri6y5MAGHz6L+BBdE0uO0w1Sy+21a5xZIXI5geJFoZazQWiFXKlK6G+59dtiP3dj
8i7h5WB3q6EVhE2LP2fLzUYduoPdazXa+wFqu/MRyP/qwWw5a4TNyuGT5cJak3VTkNFtHe3eJUkY
JctRhmkE72p7QWpJjrqGinD6w5/tyqnZA4GfiFn0MaLeX1wYTwFMOGq8MJIApH2rP2ETNZ2TdVDu
MPJQ9qRb5Bzj3tYr7WIWmh/sijVGB7qGmHOxdlI8R0Og6yiFbkXd4zmR8WycLX2mY/BKN9bbS1xP
4jIHA1tLGNQYJ1LzqGTZVAi/NSEY2ECTCO+A3U2LcaFpOz90EhOrWscrXc+glKisQAeqQ3YP1oWG
vv/gI/zsnsQltheisN0NPlw9vViF+ddbUIiVo8cke6Hqtk+MtEQeAIDeU9tB5EJeYiQsP3AIPX7Y
/pbV8lLw7O2gb/pEK2CgKcChF7+LMMnjv1Zz7p22KVwLMFAglOlSO2yLD3524ZNv6glLqU8Egqwc
1g7nixV4N85uCLv1stvjMknRl3h3Jw2pGFkpd7087Rg+9BW6Mj2Cs68YtpuQsYJPtCiyU1U5cwV0
jIVLLcSO9o3IuT5ohtMJcMWo+hOKeXhVPs3l0zmfKt0SxlP8D4H5PTSE7V8IDrgklM0J9mekgrr6
nYX7VT48ZK4xo/wQ6EeTs3gYd/Pm/orbB5hbzDTnqULkCrIrkqVEXvLryZj11Ra/V9PSMUClTfl6
g1shxKDKHVpfgetVH8mo1Eg/7AEfr2hJRDveb3vQeJ6ToCmvnSmR7J+s9yOshQErm2OUsLlF0v3B
PNWMIuEPcQHYJ0KPTvUH1JLGsIy7x+AnrzBnmBQlB43mwdWBv5p7RW760iiRouwYHMor/uavH7ep
CIfFlm9Pi8XWjMIXe365tMSG9x0TwuwVxDiabAWBWNgBHiWjSZPzsHHlaRAYuVW3nKnAAJfOQlom
YMxQSsypCh78qrLjIN7L8FeEPEK9iQm75bAz7Cn6JuZ3icr0Hq6E2U2RywOsULYqZ9RPTIVkjUFN
sCoi4NjFMWnyAYLOX5/LfNmmq5rG+1Y68T38uBLycvilOnhyLDY0JKC4nhWXK2J0OJaqq5HVkQgP
p7NSOhZaSNCQ6rlgoJ8xpoBmehQeDJOxmlbONJ1LgiVqGAxeZa59dnS+CzQmODgH8XV11Lz8VKqM
Ntb17mgz1sliTOiD6dGPT1jRnmc/MCJ8Ho7QHrMGSJ+Oc1sK0His4hSSlcMW5byM00hsJ1qVrkI5
O2M+HSxW9u9F4PsHD9UXQIGUVlMk2vE/ppK21UDWhLqqXTNSNNJX05TSQynvvHbD5qTVY7T7Y5uP
JuxQOrVZEOOR0fORowb5rVxUY81l1ewofDLF5sBo9XWpEWpWbj4kuYLPfLmYlONd7OIpZizyVqQr
YD25YBqDthsurKnh2UBXqsMXoxwvLR6YKq+HeQycpRb+FDuaO6jXYmCXLqb11k80osToo4AkQlQC
JEXvIGq0rIZjYMDvhCXf9TEgNi6AXb40H3ZTnxqpp/p4VKoZsgoYD8nrY5dP4hN/PvlhoNhfKQ74
ca0b+ww806zZaglY2S9Zjl4lsvc8ikIDS/AYj2eCHnBfUYctc1BeQsKwgzH5eyPJIuchtd0FgmyQ
8YqImPbcsQ56vE0FKlqvMUQfYF4f45VUyWR+EpPqbuXxSj4hkGaYbIvLa0HA4P/XPcSGWrCNJ0yT
xSsVdylpqfJTwHMvuG1PAwf08fPmuHqs/a++LqbY8OParYvXNhOShnWo/P2hhm5U7LRqxr7dABAc
+RhNQFsl+MRh6v4TvrAQ6wTHML5VHIz4ARaSoFpD/ir4djF2qevKqF4aTKMZL14Dtzj0A/DX0epU
9hTaEAOS8B1/dNjrirtYyySG+KS3BUS2XqDmaWPBYFeMNQFsTBiT+oq6F/L6KeQ3DR4ctIFk3k1o
o0GUqN2NIF+GvF4qQjARbQ/t3E0NXgMCYFpjLSobVsC68vIsVEuxkQa5l0CJ2FosG4dOe03dEhal
VJ/XjgEJB59vPl0V2z1r6fKfGB+uNuK7S9pNvWHqzZWuU24n47Bly/TgTPlKEZfFDIiNZo6Pb2U1
L3mZ/tvFe0nTbt+EIPG8PZXKgjK7PVBXofyqubmNsn7djeCc7PBTKL++xosn1dl/z9DxbVMITUU5
T9lACM2yN0vLA9QX0TMp29gD3BpXpiCooOLGrhkUG0L0CGO99fG37k/P7W51DOQY3XhZNSdYftuz
Wt5pB97dnuaedMjnXndOfQGLDnNsCC8AiGDktvsrRg2ZwtelUetqhUAkeycJuvYF6rjek/hexcZg
BzKiG4lh9LWp3sy7pqAIiWMcgRP+EyvITApMWQIN9sIZjkwPA/xj9LXa84BzgUdNEdJVftOU82Oc
92oJuPOVriumCTV01sPq/Hp1lNgkJZ5B64t7Xh7pbIoh/IgBhlWWbdd71S/4ibjecXRTgcx165uZ
bXy9y0/zXOLVXorMn13WJxWF8qDsiZAACiQ71amtzNEJV8LyD1XnxyBShmTdXX+YLea4Cy27inLC
KC9DuIXDv0r0eiJuErex+U2tK6HE6Cg0/AOSWZXHtuuUPDzCxlFITcAIK/UAvV9EqX6gxZTzAN6r
8xCJkfOwqKRsvxADPzC6KJ8RkbCApg8E6AiskLAU6t6RnlG2reAbRYi09QDlJhPG15SIG6zhjLWn
2kKwAe+XAUh+fwzytFefhJbT5hpnTJL1Xlc4xU3j98T/8PJ/elkw2gwfJNr1zVTmHEIISwWkRI+z
9qhRim35hpHmh/womDxLFK49wAZ9YynkwGHrWqFioVOOb4oHH18S88y9uEIPIOA0Fl2RDOq3ABdf
siz6FhFZ2Shj7dR+K/zaaDS4nVDL694wf0+ItXLLIEqmMnCcGXNKcDv+FoR9dY8jSpxZ4FSDNaQT
m9z8fo5RnD/VRystYsTB6WNJbsInmFW0dY6EYPxg2ccPrE+sVd0c6869keaktNPcSriiu+nNpZC1
G8Mclskltih4TFVzR3UBopFpd6qjjEq0DwRjpPzgWrecAoVZLM6/Qb2byL4KFYBMTsJ49qMH/Ajk
LaqaP7ADTaZNR+IrpQqrO0Mb+jBis8RUa4n5zz0ZWg75VT+pc6iEirfyMS2GCGzt2WQgZN0Z3d2D
o7UvVm9feE3rI7DelQRWxI4ZpYkmZ+2c74D7tosFgKNmQNdxyFPOIIWosICwg7S5hg7aQ04Jai5V
iLmct/EiZD5jmS4Q1UxSlCVQtCquyu7La9Yj9PZWUzwv6Gwff6DdjRTmV25eXwBG/iqjUpo013bo
wJYEBLdYNCQGu3jjK4w1jriTvrzSNTRRhYapNYWkqqwkpFSch5myqfVTn/MEFeo+4Zw2NGfrw62q
U4HOZAc+Vn51imSAFfc4tK4hvJp/KEv8uN1+xEP+TW1k/7ahqisd+nFpn+CWkgCcr5BirojOAn6G
S5XcyttBSK4/lkOivHkB1wD+vuJKBFtx4hvJhAVYVZgJSpbgTGrjQ8nyocc43CIT+qZYDLPWwEKq
IKOvNp2SvG0cBbSNEp+w/UmuRkVmaF//pNBzjD9dYZ8px2VhPrHQcM0Bh5qacuTV0dGTd7N8EjSs
4qxJoKqnOHwrqgy+F1/qZsUJUHVlT+vZ0OEwto8GjCZl9DfS0FbshkK0LEDWLThP+N6P+uRxHc8o
COKgDSuoQLM/Mqj90st5SsFh9Ja1KuH/otczycZkUgYSPgsVSMvRkZJmZUb7+mtj8WTYYYPPzZjH
NIdP2pR/8GkQsvVphM81JaJx2mc1Y7qxVOj640ulhHC/+o8786dPgy/aM7nLHFJ1QLTWGr/qZjzx
D3zJH2gx4x1BGnJU7v7SpiXwYJ0O5X4Ddxc80JaKxlJ5oJN4HXss2rMaF+a5gHrrQOvwQsgKZ8ev
1uf3Bf81aH/ZSPGPAcgbSfoSA1KHebqBkCkLM+46mMYDMxApAtjXRXmWymVstL+BwoiMdccp/CW/
HzFN2/XpRV6oDlrr9c6oGmXqAZzlJFW8hP5mZjigW60j388Mgzd/C8k9YXeMvyLBZgqbGasC6W7+
Uih0b+aQZIIns7a7P9r478PcJwTOvmDKKrx00psePnWztkhWuzKVojXZxI6S6ybNpSCmM/UjqVrR
W0dEQqRa4QT6vAg3/eSQxsPnI+COT5O+RAXNGkY5VufTgrJe1LxNazpUSu0nXzocLhUnJv0AniSB
b4iYXWoabjIcg+JiVBuTxAA2TIYZVXNoI4gegu5F7bEbZikNRGwQTzS56Rr94poQ6z3JpnC9Jaas
REeQczEDofbj/gl+hmog9v+8bJm4ML+LoIh8e4Cxs7Yi0ntnvgDYSNe5R5X14D1MkwX9YaneRNWw
xXJQU5FA3ya7Iy2ji/iDlxzTDQ+97Lx6cUkJbh47jXNIxzrJNc/VLiGUDs5HRAvNyNjb5uDzJSLz
IjJjK3Qb+1/FoOTQMzC4gbsobkJOnUeMnraX8sJvTWO7xGpJpmTudLbaCCvm5v3ftnKYUIeN3MAN
2RyzbNn03sUZe7AtzcGMCRZYlKHTKPZzUOI2UTNxmGjVFul7kDAJ2rXUSHYFYOp1edpZUfkHybfB
2HpmiJ3XKF6H8QazKE6ZVGb5OQMw2SVPnPONQ1lcGX3simO5DTxaSm9RII0iAQM8G9oWsp1cTxT3
gJ8F5ZUx9ej6+i8nmYo1nYaSt/JTsfhsMyMFM+LQkR52cic3tUuKqfzOWvJmZQlA/Vra0d8nuYvW
EOq7xuHRPGbTwDqgn57XjSjM3bBV5Y7T76zzlrGSvO+4eJtloJZjgGrkVqSSfb5TpKpYD9FOboSz
fsKOR5cKNksxh88EeUpoADXo/l6UwugSI6IP/xmpoF2MJamMV5rQksEAUOJ3QDztRPzNS5pvxx21
bS+pVCK1ZQHK8NwTzUSqq1+M58dZYHg8RVvoBMCV2YlZ4mHbRlQFKKta1ubhMy0jKgj8B1jV4LGn
iLlwGP6ooIq9tppX4YGZNjU2SBkNSaTUPUHXn2MvFaDBN+M8rXgLQT3yrq5vU83f7bFP5p7bkuuf
/asX3MMX500u6n/qfWI5/bMxYEmzwEsOlVEtb/zAOd34xCvNz6/KhnAMGKLM6+qZwSRvEqJ+yNW0
wWY1rfap/h1so40OdoqDWX47L90XZDjWRnjkZ+BcpHy9963RCGUVg0nwFgJSr6u+Ju6N+d9aAQvf
M5bNBE771v8pLu0rh5hZ2v3nVDyY87cAoGt6QBkvvKOwi75gjdj6uKSe5JZfqZnY5XnYAF7ZQ5sD
rMsny3KS6gG8SSkTUPfFWOtwXYu3ZBNlkXVEv9uL2XDRIl1n4aijNG0dkEfzEz+1jLlNB0NPi8Sq
1e8dim8K43qwxPdASKPiCzPNI5Atvg59DBQuZYM5QxAPok0oLyorzUDnWmSvnppTkTl15xQIV4F+
m91HnDGFttwGJ7pggsPvZ4rAG0x22XSZRaAEHyeidguDDIlqtXsr5IaDQmN7QBJ2ej6Wv0R7Wr6q
WNi72Hg3Wi8e36S5C6Tfovo0cGWFQc1Co3/vptS+FG+yN5Id1I4a9BSKan/Qlc1ei9CbhTJUlyTs
puyuH/2PhuaoF7aaVXDOzmOyqI8fgGw4FeVRwvlGF9OVUAx7MN7ytdtwo7A/PnIx8jJvmow7RuNc
kM5K7HxccJD9jCry1+Xgvc6P5IFgVgAuvBVDEWL9AH7XE3I9ezQOsxfVGJGAHrH4AkN9as4cAaNz
205mf4id5U9bunU4ykpnnesMzoREl7rl/Nc0BqSCthTp8LuvZul10pirTXLs0IfYDKeMKe1PBIwG
/EZojSJ7cyWKnALFvkmtjvldQZLuBWhHtFuMEh2/KPdT5R8oGbA8aGeUwjM2XdVRpKCylinM7zYS
VCHr2osT49qI7f+656D6JCSeoll8QwadKUaqTm7KHZJUFuYf60NSutHg1HJRnQWNF2rC5D12deEb
tDDiwbbokGXb92b+U1bgTNHBN06X0Q/M6ErRHeoFex53V6BiMawOG8d3kUBeEp+YGXH/540XXbiu
vFj+nDI61gY7gYMazzu0uYYeMhgV1Va3HLLYHGhHrYOFuOuxHwMRGnMUoVJ/42fN5wFm2wHWunIG
6E/S7klIfsTPxNRyjK6iQ99fJw1okkWZxySOO/A+FeeaSFupM2zm8Q7AwVaOk9klNn5q07F/SJR6
jJLRapQQpHXcnLoPdHGD3iNilPzxPf8zHjLq/Tbkn0TMo9Hq6PBCnzuSOTouyFSOB7YPd9x4EPCF
ITpvONEP+4SR/lNqu2KsYDNi8qI8yHX4BDzRpisM7Rap+ivzKbt0Kpr99iaBkKsPDdn3V1ekhld1
M2wbmUxLcT6ISWH7IBn/Px2t4m5+S4ljRkFUQ2l4krgCaFst2ndtsbYlsZmOCGvt567CWxyZNBc5
RuP46PLgGQ8ur+OhG8xq3VNz254klPrWEKGnUhMX1JbdGD61cmS62LTZVVPITx1ppQfTn3luZukN
DC1JyxZiuSvyra+3VSsMP0ZscGrBthpB2h9qxagVywzM9yVuqIZRyUdEsGDtWuUCn4OciVHUBDpy
IT33DI5hhdQ1jMQURcnAmrBBVAgKdReo1R99wYd4RKXfUUpRSt1FDbEfi2smOyvSq0NtaM9WK4pA
1azuiC+PSP3uTrc/jajoLYIjHDtytH8nWvLn1Z7RlBeBYcJkz4n8/HftA1BwOuo8zd6CJQHs/Ldr
2XBXOIhQ+pU6u3QAYuVIzl+NIroWohdTlYLM3GDAaZwmhu8OA+o2eKbaIEhUw45joau9NvWdWzVI
uu7X0+4UVhfoIloHgFrfvJZZ0PYF5PZHKfWRMxgbTvyRhblbzKrtAPc4GJXWIkZXaNC+/Do9mZEI
sp5dwI6EdfAEdT7xugewtw0ammV9SeUBHEStDAXbDLhiqt1oY3hYpLvMr1mCW2hLlsRzAHg7gBOx
/RaLugiO2KKIsU7oXMI90Yue/Qimd1yeDQYkLchqnCPlysBQvWS4va2q1GDCcMc3m6gQoSiEuWEl
3FTcW43mq7W7HNOdodikU6tfn4QhxhMObTzmCrDk4WbzAfWHEfvTU2sLhedbuZ3VAdX7ZxnJEKy2
N6aFKolF/+GrW3b0n8PlkylQu+yihPOBTTQC+unHCwHRU5G3OeRS+v3wtc2mj+p/PCFriRfJtCuY
R/KpcTmi+afxB7tWjXf+rhc6gU0DGo+G9EtwzQTWhV+pH0Ao89G942Tu5nj7rOliYChp4ltOMHhQ
ry/tIBntOD67pwK6U32wO3xznUxKP+pelr7O4qKDpm4rLZr2R8mmp5gmkp8zA5Th59kGZThGf+74
edVw8PRF7icd079dM9HahovYm2juOxfWPtBOPKvbs1wdqDwGYJctPiUDiXTncuG62xYV9S7ETMwx
fUxPnflyja27NAO0is2bsmTAbUZgtM7cxKlHfMA/Xq1izKEmvsXSQWEvaj0JlwTCUKdXNmOz2CVU
OJTlC38HhC2yA/IX3GnguctcgFWpxPDQHB6tuH9B3QY65Hm7TgOCMXGcoRcZwc/c8pOyETcvSZZl
Uyp7LUss9p0CU8MzAQwhESfqN+uYv3RBTVIktLP0HkwgROg3Z/dmQihUymiOdrA9oyikOMlMcALD
BaFym4eul9Yu3gSo63H0cX250bWDRtJOTwUMP0ntg06DafnvlGBWr3oIyMExQafW2Y0Lx2dJNDb9
lILqJLGTwPpFdDrUTwk6Wz0szuo+B+8L6DYt4dYypgGgpruWAV2K4HBDgbYYB7n3svw9L8B7mgmO
olbKBeIfi8tDtt2gNprXAeUMYRUSFvdLcJbjnqU2cnZOG5sJxLLzJetlCSj5g//rM4AjbewfJ9om
PQU8OFF6m28+WMDoIXRIeLump5CWoBomzU0XpopbYu1hqa90lJSqVxID7pniQ4Yp4Kdx0GA0HMCE
nT7EoZ/DirEWxwXQgqvRUw8uIqklR7cosKMACMeoDFRUHGAv7cjieejBgJnxSdCFPiFRI671EnvT
Iyf8EzKUOWulB+M2cOyoRPpm+mjDbD/ah0UZmjEJhsQk+WYeiukK0YkaM0w1aZklbma58hcpbIVd
9oZ7C+d4Va6kL8wa/IOzo8QQK9A1q9qjeiEZnwL5lwoZKtTQEuNCF8sjA8fGWf1zlhBLhWyO0hqk
JuGNwpaVFQo8IzVNeph1TtEdi1R1lwo1+a2KIIxWM38pLiGa1zOR/9tAGkhUNSdd4qFETJ+Yf/CT
HUIyRgztJhns8qC0ngkpClSJR1Oasu8/vusMCFyA2Qq/O2d7flEpK4tUm14sad0uKLxv0eShiavT
b9+e6GVfBdOdACteG76Vn7qxrgW9+N9GVTy9hfqQcTxGkXaWzWcIr1F6f3rvmqTuRyy2Z6HGdkGd
JovcHulcrUmFB+BxBxp/ZwuOSyt43xAM5ZLKqd1NXdyyXOuJotdx5QmLsNA5Z0lytvD9DN0esTRj
JfLrOPrilIx6rigN9xa1NEAkjgVxKqgdsm9pR68DfCuTW8PDLYhQVdSV5vz9Q3aRzmaAuylEeg7e
pyudT05sROc5QbA/VGi2dljXUaQARsT+egWyFxvJBrXlEtH+wRmyvx8G+lQ7NLaJvfeIjQZDV1TQ
Z4PZjNreu5Xi//EUm/RbHf5rfYqA9z9m7HoCSoxx0WU2sfpMkZAoWEcGAMWstfGG6L51UH2kFywk
dvjwbk901ifD97db/1wHLp/4hUMEtRWbxpgiGyYao80wVi4M4hTHT+hET+pWewGifmc4F0ItDl1Z
fERf/c5U6Y1PdsJsre26OMnxuJKdYZzpGCwVcRfvSFUurDDcAbANemBlfjOts46WuPbrNy/EDteU
qG2vH4Zc/G4pTI0Gm5xOA8Xb1KnVyZlSLh1YO8feMyc6jvHf992ysO7CCO6AbERJWzLGF42EqhgA
Y9Y/QzURSwHk9qAacCGY/CACMetcoXa2C83hUIH6jxMx/oQ3xImdQ8c/v8noiU0/ywxZrf7Sb2l4
dngfsPluhpiBouSpHfGYgIjlWIIO0ucasb9/M4GymcVBCZHDA6y+WRzkKKxQ3EMSZhPrkqrmKU7c
5J9IS+J8gyCtlytoPIIxZDsaDxdUg8MTcZdc38DwxsiLwxcP3S5hlw5TU3NZzOKlf9swNjB2XhgL
Qz+9J/5+0fuuUEtDoQiICVj/6U/ETD4JWHZRCcE3+ouZxdKQVyQjXjjSHQ3bDf/EhdMzkYiv6gRK
w2kJAS2mC8COY7oiQO8eSJBEVWj3+ilpiHMyrPOYofxTyl7x8Q5f28XXKnyXWTJGlbkz9puGopvn
s7LmtmlCuaAYJHRMEd9UUN3w+Ib2e0qtpgk6OkixOxbGBuNd5aBRE2CnBlIvHmQtUzEt7G8dviQ8
MJfyGYnKZF+1v8CWJICFI0Nco6Xs8rQX0luw5D09d0d6E08gDwHEdNSCqrheqbNoYFsE8fh8GCkH
L+QAScHxJdckmvq0hFxIwhKUcFGcTbEVFTEU8LJupfACnJ75EEGs5mLElfSzVrb6E/NkwBYbX0rs
Ua5g2uugh+T099S/OYuzdU+FIZ4Wv4DwvhxM2uXMrl+YpPvWgqbnl/mAxB0rU4rK0iH6EucT8Xjp
EJNdwxMhU5/8EQKPlyGY0+Zj3rYEVcV35QiqKUoVVf8DDKwmppZuvoBdU64b1SNO48x7ShVSC60m
BbzlWGMRbFyfc7TU6ZdLlY19uW7R/Tsgc2Rh2jHxYjMaRVF9Kx739+wHbw8ouJ7I6u770ayt/Sch
3FopBYI/oJ8rV23HzxFHgNlu8B8kkMvlljW+wuFc+X+DQkHjQjPTb3DmSPU/wDbdO3s8mu+4KZ/S
Qw1oSgffxYnKiisol6G8aIw1gf0Yhgm2AmOzWeKGtJ8s8/uUwWpiW/Z++owvGcTxZ4cF8m0gqGrT
/FUmlWOtPjJvRQK/9l58EJPjN08Bd68vTf66cygmYaDokcz2MflLmHR9AQ7sQ1p3CFGbFuGelK5O
BAcAAY2vBr+bCotmLwZJpJW9Qh9BM2NJGXK8pZhmwHmuGpb+4ZFNuSAT/8pdJECZhEgWroCPTtEn
7eN9/h7m7CSlW/rKLw6zbI4K3uQRCwjW5QF3b4g+TEU+lmG62qvGNV/ksDJSyJ1+Av0YgoBrhAD1
xoBBvwSDgQ+CvV0wDYwm5lhb3eZjAic3zN1lhCXAyfbXrVEYF6etKFXfyM2CFl9zNTnHKM+CceJT
joLQfWiDuZmeA4iALJaq47ZKJpftO49e95OGSEy7bSTAwx5+oP4kfz+PmYLYBLUMZTPUDWVV2LT/
lMJ5pNKz+1JwX6cIUkqlMuU8PVTQCwwzgxvneCgnGKsvfk8sYtlk/2aFUVyRAx9cqhXSIS/5FMZO
jK76uSwU+XPsWaMYpqinz6PhTlghSmL9eeP2Q4cbtmuVA3wtdbHiroBM95/57O+vSgBlNZhavBtz
i/mN852z+nwxYb1RqdU01Z1WvM2Euvw6v/h8j9CKta0inB/Bf7YvH6tjtfwvgw6AznTgpFn9e0Ge
S5sWCmw0NIAlBqjvzlEUgOREXCiQuv3z+Lrr8uOn0IUhBPAR+yf0lnAC0HBlLe/6IdF4+JSug7uI
W8RCw/PkC4toReJL2UOLjEQkAo19oRzCGwlTT6+Ie1qy4yf6sOMZ1f8pZ3C66ptsCll0yRfGWsts
JY+XmNCSLvANAgsHEn6nnDah6dzm4C7WfCglRZtQjyjAom0Gin8LBQnzJcmKgf7lpZkUUdYkqtaP
T3NRHRvRKrQJOCXOja7Lnka85f0tdeeHSky3vGQTUVRh5dvG0gjtZPA+Atmf5icBun8kSYNVw2Do
GiythvYVn0EM02vj0A97kdz+gp7qRi4rHrhrw2LXvn5cSMIjfycaGnGf1rbAO8C32PJ2/ZBxcdC+
ZLTPNItXCohfJxZcCwowVfqjdHtHQNBfKo2CKnUJyth9LBWholtedFt9+My4S045DNVr0zHz4mfb
tn2N0Ct9L2XXC+0nSIWDw0QEFuor6pRw48dBV3n4Z28QDcDfLW1sjlqNQ56KjLDRjUy6lFHqK6Jb
3yfOD1gcZM7+TSLdsQsbI9PD3UL0j6Ew8YmaEcwWNcukcxDzSWDh8Ym7vP1yvjj4b8IuPi2WS2T8
veibYpmiJde1u1vw8sLZYcFvRf6L5zCFu+k0Ar43B8U1ET0deo+QHchJHIQR2fRoL3B1kVPdX1aR
hogfTf2mMouB77zm32CiM5jurbr3H29/6ggCraNLGO0PQa3t5dySj5bnAB+V2KeBDXyQ6zfT9esl
xOPxakpYNWZDMDYy9pPyjsnnDoA0H335d/F7gBqDjhUbtWSDA+dWCHUEseK2xlc0BKM6Oocx+mUQ
Lzfbh8BDX8UjK3TELNlzceCXXo0LoxxiXDEQ0nZW06xtA+SyUJznTOL/IBUzLv7UX5h089Zggxef
zb1sMV0FkRJxssj/OIePpcTFRqE/w0SGzVQF9adnYd6o95/Y8oQD4h5SLwy6URywijYfyB8q2T6P
ecogtmdc4WuJJ08F51V2ShAi4zNY311ETGDyi4qSXUQPbuhO13efMsdgGqvvW5gU6OeAZtL5v84b
ICaCLYif2qsFYRaU2FCFIvmzTqzErK2cF1+5fhdCZWTAghCAPmcWZURpI+Hy6vJm2ylUD2ssjdcI
n/R4qkFbPGCbvHmCs0k0d9w2ULa0aZapGv9CPSGuP6we6LcWOGYV9p/uDE+n0u5qRGuA1uaOh6vJ
azXWe+dNsB6uvxpXRzelvIILh/46Xvm4zy2n+SPRCijEhKk/Y8lQWTAvsXr7yjP/cidSend3L2aG
zbVY0jwSojoIO75fP8l3QHz+gBYSyU9wbXdDlc7v3IfW0GJqQIqe9ghW/DdK8wcHn+zYljjuFLlM
8pjhrrbGKSQGqC92gnIXuJHLeUe1/8t/XSTLX4CUezZlOKafmX0hCuaCnu/BFot2vWKAiFHrdJDc
6MRVZxOEKzYokUHDmoPIEOMFS4BCoMrP+TCUYjNsHO7NCMH/XhuIKkmRnQFT1R80+5xt9IK70CZt
SlDpsIQU0Jw3QxAKx52Ftl7iYASwxzTCFKL3RA7aWwufLd1ATGaQMFje6E+3tZtbb2mOgDQSVuWq
NsUCKtbez832KN5t7J41Q1uNHni2xtix0UFaC89ebPqGt2thXT7Z6w1MfRPikII1are3WkXvsBX1
X7CUrA3UHn/PLtnjz1JTDBvvbwaygKsICbekdYrXJBp8ZaCH7I45HYVpIqFseCvYckoaT1jzjRmH
Zip4ZFyNhig4D2yYOJjPs8Fj1wuHCBxuLn+eBNuUFIweu3zFPLa1Kxux0kp9Kseae7OzMzn+wTUH
l/YkeBcKLCi9q59dIs7J1p+GeloZ2yI9wzbI1iSBv+2Pq+1P1TZzBfCmxlz3t2BunYMZmEc65jKG
aBER3VTI1Gg/iJQ3e1jCqFvyr+iqjA8xlu9G/8m3tXJAXZuA8Kqw9LpRig/ylTDZJBluDdGWAplD
l5Of5qswd9ETlvTCEzZCMxpC1vWaqUACYXWgERcqolV7c8uoVKysw/Zc5/3fjy0dE2PUZbrLKLX1
ZMynJpxi1t67W90pVHg0utUa/zkyi7V2ofU8tAJjgi9/MDG/w4UM/y2D9KYKtpLDD8PSdVSRt0Az
WJfPywrB5MrYGehvJuaUR0MUL0QF+X5x8FMOe6+DPpuzzF8ev++TZYtUVi1vQlvqUVb0g7OdUF6V
DJDdBRhqrPWFpyKh4pEtI64cKKeYAMWnqCNrwIFPZyliTYMZZAfSBgfVo4F852sY+0O1MJjbJxRK
Xsmpwmyg92cE6+ZNU/VbQrjSqXN5BjF2B+bB3E0Y3wN9R/lQezIAXSfxrH+Uj5CleAITnnaOsqd3
+9VW1PFfJMZoo+co6PzCWSz1UGv3RZEOTo+hsOcrb2wWuuLqVhAQ+SszK4Q1PcoT5GIUL0qfBzQP
03LX3my1SbIy6drSoUHtflqTxI1wneBuThtUG+N7oNhUyc8bHRDtX/IPUS+xNQ0vexs32o5jPBlU
lGhF59/C7ykmLCUhfhGFcwTlxbziIaPNFjmvE+bbQgQFxw8yrWPt8fT52xWtkRXPu4kU5r4bHU4T
LhW2sQUtZQGtvIBykTJPobCwxZAfdg8tYgqas39jH8P60s8oDs46sIEWVsWWet0DkopQVNVIONX4
a1EAAdzufHzKjW29AbxGDKkqrD5BzCbcbZeeL4C1lr4r6WNmSsIoOTgm022yZb1wWu7CrJV+GyyV
wNB7e/NaVxfX3rT+gcWWnc7cx5od1+RfxLPNvJ6gBiLLGv/g7Sbhg7tzB8pH28zjlwXTGzvA/XfM
jUgrIx3Q37Po3rrRXciRKFSUsB9EulezlzdLLq95ifC4MbE1CgTca4Ok5E3beZm7VWQvITapE1H4
5Z3P9Qb4pvrmq+HEviHPnwPnznUcd0fxiIlhRxmExVA9c9fYL5CTb3OwPLbOgNgt8WDI8CCROanA
J6NY2NC7F6m7ntJIPTfkZZpqiF3R3SnVB69BsyN//3J2N17RLRe+Y8N+F+ZylCw24Xlgkq80OdAl
fEU/dXtTHeC+VS+k8bYg2aQRDJBcpA6f+0Emyyt1IdpqMExX2uJ7Rp/QELM6NjNnxvbY2gQ3d7pJ
ZhzElwGKk/eiX8k43SQ5qvLEKMtLCc+xDrk0I/uds2u4ZxsthbMWx3wyhaU6JKWsmyCzE2gJRsR5
ENS+6p6AjwZgC+gyTalR8P1QCID5E9T/FzLW+SieyYYGW++FNCfAU5wxp5iL8ifeZNcwYB/YrCP9
AEpLj79tbjnxdsaZ/bsP0QigAewlI8Rowh/Z8849rPiAV4n4I09lef84rZVbIr8rkYlRE+gdUIJv
sP8ppDsmf2X1sn4THBWYgSTxJeabqQ4evMf4zben97HcMyNq9j0BssznnjVlVLw0QPMmJHGTavxT
u31+eLqO/y0umSJxT5mjloOeYZXZjcPJ4/PoGmuzeTL5ZYlUnlHYGp9lVAWuOZg224UsFNe9+dWS
X0j3k+7fEHDqpEtPelA+BKMOI+FlaxZ3irMrJ/G4C89yJ/HK9eG2lcZujdvo7Zqd6bF2uCsA2AUR
XuOouNaxfkgn4QV4LtA9KA2oqyu42gyJDgFSybAymxI0r2LiMWrYbzkh1i9qmHbSrNNHvdYniIKP
wsLkJehQOMudaF82xPDHhtwajwOEimsV8zTxjzpuv+lzoYgdXISFZIGI0WBQDownbpMXAsck/OVz
7f/KcPZ5mwIqQmAGLpXMgXPIehkLA/QEtEtQhELh9mYU60KTxUXa9U6rC5qZRzRDKGn+dHiFciHb
DxLLYgtTJ/1W5Tq6c7cvLFiDpixyRa/Yt2SNi02LFc160GbvTXcjllwwRT1fS7rF2F/qK2YsDpUT
jFGshbQDR/tWz1t7nGfONR/gkXU4d4IX3ThDA5RzKEpGTywYcuq1OephkwPDo+Y7RUpxWQe9XmPz
l/6nu3H6d+O7HomaAuG5okdqB+gQEEFYe4dSoS31YTPKHTUCXWuR7bBtcsF9Tj3+oA1iK89QktUQ
x8TWf4fgHvrGL/xREjMXA23TNhyPwTC9QDcRlnfigv+0XVA0q/OoBMN9UN7lNe5/6pop1OEPBnOv
v8FrPph1ZX2yrq0bZr8UwQYkBQQ967lqHGOt2fbV6t4krxHPx4rJ/mTb4DGWCcc5dGA/MOL6xBNB
gatr5BV53HAssfq6wVzuM/FLu6rmNDAhgs12MpDEF35LuJUKSPeFJS97/urJ3umXG9F8CWybiUEa
zjDQcwCZNlDOsWb6eHXcEpwHhyX9yxQKo04KZ4xKbJHHqeZhahPuP8CnXVpFyzpFgPLtDj9otpLR
WQgLIGNb65j1DE/iZw98rZrTlmzI7tEmg/ZeZRsxa0oY4J//X5+QqQodUCIi9q0MRwPAUP2vsZbC
3GOCpdpsu7h79zQodwOA8Wf6cExbiA/0hH+UFZaMn7pgJTJtP/lAUQK5cL4+tHJaiczNNzXbnKu9
2fLZN0lxK8Wz9vqxx/YO1G463VYuYdUzRNHxlv46YBNotkwmNwoz2b9XlQKHdoiJ0fPr9F9ZHLzT
PzmSwZIZX11/XE/pzcvorZ38Tt7m42EmgzLGr+zF8qhbWkS8loDv6CJlqSTm0+mR93BGJRxjLNt+
7C9aapg1znU/h44n+9X1OZSWxCaHCsLMJFwwObisMAe+VQh4KP1rnY0KQYDovS3fdm8x9j3B9Vz3
Kv+YsNZnPtU6eBVJuM7CYuEAoT0ufqrCcc0byEmMhT3id/BhJbyRX3h6dh1LjarhoR5CIUCvrje4
MzIHmFCMagzrzsBEg/XtKQcGph++2pmcTbAFXVobmkpcYYKYCE5HKhEt9ouBgf6xW6VVFxWRqKpb
qrEzuFrUhin6ZUZrbkrV3/sE91OvvDnliKG/nQm+cHtneb1y/NOO6TfbpY+2kq0ykdHiGVm5Adl6
/dWOjjrfb/hAdHJw1uMWXNxRiFfIiF1xwVbgDq/MFUJMYdsScAdjZq27PEBRxoZ1l8wHdHtc8k4r
zY7obgop1BNo5RGJwYsfnHBmC1j5tzBx/IJMqsisZe5I8FOlRHxeJidkOMaUmC5WPITtzka0qalr
urOwIVWrHGKYTAaOO7nZtOuGGCu8UTtpK+ttoQ2cYfDlfRZ6Vt0RT2XFRxxQT52BZYpXrsL/ybq/
+owyAKQd8Av7g3Jj657UdRa87PWAWkSyWvk3sO7Jpz/KOS1O4CiuDT0sHhO3ZcEBJyjiZubUod+1
5g6yRWeS/IEe608T8tbbKxpXfMvn8EXYsp5h+lLPtnoY0F7Rs0TBxtbrdiyYabvvqW9Fn1U4VFoA
EDHnQXtvBj/F9l+RHPKRZu7YUHCWkd6MJKQtDxCuR/vKeeNSQvtmQesNXlQ0Kb677gzQ8uUd/Uyv
i7qNpSNQ7eFMgHw84a4UKsyQvDD989PZwNHnvxnMNSJE/00R4EeDGe3sP/EmD1rJMF9xBFzH9vM7
qPDMuMT0BO4SiRQld2YcO9K84PkaWLpAAw5gO+SlghuuBf4tPWVvzyC8vMdVBOkgayoSjiPaW7ek
WfhmfpLSArwQQdss9/2KMqS6y99qT6mpfZEmqgj6irIZ+mwiOfHdB72z0fkXnNTjjI2EqblkFbuw
rrzthTbu9dNMYIcq4PwJb/Gw/iVLqUfYf98lzGQif73BUezqy9XzFqb+nZ822P9cDCTTGxxUsXK2
bdt7NhQsL5IWupiDnyVAi44XW1nSMmHLOgMRo8iozWgMbj2lW4RyKS1MTzisGscAyM4JomeSPu+v
aYo9lRXQC8IF9adKDdJqtvMQv7wHnRYPpx4QlCObxfyQ+W0c1/d05r6s1yEaVZZUgBeV6Zf5ZLZb
Hje/CBTXqSWQzXynG92PV9jPTvXr/MLg8YMvWuPUVY9MgO7Ixny+Yuz5oIuy863KzvfaOUHmMBgg
zS9O8hlJKSRfoZrArlbUvrPe2IG9dRVPfmlRwt7UR9mNGtp0dFMTo3AZ0i+u+0plhikV+9mpWBvg
5Ndx1X7iT9OkqcP3xs2DTRq+PssnzcHFEcAKlygpoZAfSHgYmHmycwnwMLEMLADVeYDM9MPUh3mn
99Dg11A17MSAFiWig1vvWs0lP6A6NC9Hi+r8O9oNSrtZT2KbPU7Rj8gWMApXvqwgN17l34+g1Qgk
MD9FXZti6e5C6fbCgJNCWeAYu0VItSRyl0cp1pS3KHXtZkulkoezWkYVp3KyjvI34jTpDgbHTmIA
UAUcZHE15qQD1I3+XIlvHdBcNg+5uT06L26wcudN1+swYGiAm1OrjFCAm5LV3E0JpEFGv0KziFWt
SqPWmbUCMWPtNnFYmGEhjvDsPIPGbIifipnt2nAR8J+OAqfIzDcTzVlaNonIa2R7UqPVSkW9jJ61
r5TPpQIiea6ARJF42SmNiQpYuz2ZX+B7Pmhzvl+3Mg/PjASQZvov9EG/B5kdrbqL6UDqLFTzz2ad
2XdnWiYLhCroy71VTjfu12H1DjO2k+BGUwM4pyTAMhpSnpKYOrcC6pD8HYtrWKrW/hFBwkpsX8J9
YR7g/hzQn4OQ7VNGFKR2Z0TVFtuvhoJ/jkxrRAnrVD7s22ZsMxwCPu75PFkSXpbhatpBFKWXSWhM
+oAUDfm/WenzlUlrUePSWXEUj/a6kLHW10eBtLK5bUF75R5i1qSwV1LrlgQ2+GWyOKJGx3GFVeTb
+aNxNE5LurusgO8LMoKCKPdMG3QFddipagRLc5I1UAuh7Dlj8d2XLWjkWdmM1e2ktP0+UapHYT0Q
DT68mT+5/xbpoJa1MiTjWyOgJy9VHcq/lqfZw3N6HTEBMG/4kauHQX3OwwBJl++rX/WFQSGBZkfJ
HjxYyc0GbcTBGo4e8KwfPoIEKXXCopV68QAat8R3tifcUcYRa956ZQF6WMWmqjDY1+IYppx5DET9
QZFKFmWZyzueeNhelHkL5x6OPqPPy0cEkgBO4L9ttRpSfHOJ65OFVUIWmsmodRXdAnqq6KDF+WK4
eco1jfbawA2Lh+wV1dvKx/VhRZT0Tpp0f4+xQhFUTpvtxGnmyaMlWSC83SzlJaqZBBMB8PAR6U8I
ZXESOLk8U2oJHeXVBY1npjeI9fMGwTnjlboWH1EcV5P/UAut3kp3coQ74zdEfRTRX79RGZ810Z0x
eZLK6n8qCMFrV3AE3OBi1R3cyZX99VJ6DOkAOTa5XGGrvoKmkVquDZHVxtMXvZNMb972ZRDdGmi/
z2vZSOsMI9IojQ3lZTAYyF8K9vdFCSwSPNAAueWFcGZZi6MS+iuhKAnharMGXGXRrqpAReqaGTjo
tHtcMUHvyKtnI7Rhv83a8cxDeTamLyRIFad3WmfzKFgmSOMhLyAjJGRboB+6CpQfYW+MJLgaL6jt
Jb9kaEds3WpPkeQ0QKr2lZ3GLdeuHipfYYQdm4kkK3LVqFKb3D2yem+RAMigY0ZtllR0lxOE78PC
c1bAJF7K//Ie2qCU6pFYUnpQf5vFtoi67sImecQLNULOyIF3bbvMzhj9RHP0bH+w1lv+WONRHS1X
OJ6hIB5NKQA9HMuMPJ9MC5SDKwJ9kIkpmnylFYXbjqO3KjIAJRQIrcTVl+v/Rtlk8Y1QPb0Nh75D
usGKoxkCkz3ttlgYUbRje2czaRFTfCPPh6mmtkUhfLH9IRBAw00pNCO3oyUM5ygQ6sxG0XHbln9+
xhDr3vgRpAg79WIOPCLkXOt7379SCi4F3rWoIuhkNFkaM0CFaaAPpKk3yV8EOLxEg94LwbtRpcBY
GN6Dz+yTx489bZAEqnd9vBzL+WtocAwXTT05pEY8RpxC/f8au/sUd9Ve/aj1+kqNGPNG7galSt4o
wmVPAArEEDG9aGVQQsI1g4tZ+wl8PRDLwGG7UBJjxz1NBz5smOoQ4SKdLRGiypaoMnnDoA9PLFYd
AYz7sz2wrWsFp7vcBbJMtcLdQG2ISJ4zbcsrN3iAcQ3qX0EsCbYTVn+Tf4nFm1bb770aO8CJNmCf
DpVKCmL1evgG6R9dtDEWXa+HFg9CBPKyr3lYVZeOELJfPQEqC6Gb2kXqlgvmgl4QPUnCUVQpQfAy
DTryxLvh8H0iqfTTF0taypawXMpinrIGEHTB4C6iqGvyDYc6KW1Cd5JX1JEbvIygR5CQLxB9jd+8
8qhN3JMmeolpx9Q6skxRaj41/KrxhJFvHJQnJ8ogqFh21ud/kdOPeKj+TGHip9AybIEKST5AW5kj
Xy7M/OvkxsdKayzVU/SDT/WAVjkN3XnnScesRwCdJWoHoufildUrFGTXz+xP07dPfFcJYvPHs7hs
6eHmir3HGTCbDSHiMA+h2o2R2QfnA70PML6RE6OPPePPeB0GPtdteN8OJrFyQZQunANteC9aJ66H
th6by4K8M65c9LpOxi9XJSWKGK+LYeqkkDYho5SpFUXsk9rU8nQzANp1PFkabNyd4qtdT0a0+xkz
gmnQgVRNIDccci3TTj3krAuAHMvuQzJI+hbd+yncKJzr8ZKzeF3/21xztlBug621QwUaRD03AMAY
QaIcg7BnVKpfxQRapCfZoW6iGQDw3AG6hbDEE6UN2LkI32nuRu+r929Ix8t5KxeR1r8Tn+rXFAoM
iFFb5t+aj3+t+co0h6wBWJbBumHcyUONI4dF4qY7Tk6cbC5LZDH1iQsiud8nRFJgDtRzxnGQ0wX2
nRjeiHEB0EGMOLupkQ0Q2r0DF05mKZf8vaKF0+8jABZPmK5Uv9cPHfhjeb5xcaN+D3bOqYC56iaL
GNVXtHSttyL8HzL2y+fSybXxwZsYnvJqvTmkJWyS0hMtfVGYdTgY5MQQEswoZ8c0FPv7cYYvDyT/
WrCMGeYrfGIprVRAlSGXK6jKWWXFtmRrrE9k4i87tbPFK0S/Tfbx9gW0fSLwwJ/sb8TPeoE13lP0
p0v13Jxa8u8ikPMy8EHCD1vzaZKF55gYxekTIcRZ5bZ1dyzys8JXqCwMaWtpwnM068EBYDa0dxMb
n9hk0nD2Fd2Xpz3Mt5TS9yAR/YhPNfZUFRhW7FqmpP8zOK+9yd28FjwwH99xWuE53cytUWu2J3z7
sBeRaje0Xl5TK7aQTDBUKsqk7X2czRwn/NtW44MtCaFl40XPYQejU2Mpyo1UMMpgEwmjdnyzxe7y
zY3zwzHncGvAqO3ZzJb/mu3djD+LzJiVtCPcsLVbL33MuyVsD+c7krY/2AARfrkZvOjOdMrjkPr/
9+SDWapgE5WsWkVSHjsslT8lOoMPIxX9aafQUS3lRL9EEHmWE/RC1xpYrZPqe6LzmMzx1p2w1SQ9
e6MEFfOEshkpUQMdFULogKQd436i1xVKyB9DgB7J/WkUraTk9hxNPYaMF1fVihTWBr8eOWrkdG1E
0Ko9B72vgpCzfksIsY0MzoWdkApL2kgUVI0Fog29AV3Wy6SA7+YMHzvRjz1XlinbLUIKoH/8GCge
E+twrOi3frdERNcFFsKO3mg25S/U1daGDpOyAo8AuUokCuAoNI+JOoEXxmJf4j27c3ujcwm125Fo
Z65gu8RbaUZsT0zbWsbH4Ss8xy+ZF0nmtN5iOO5YANmQINNmTU3VmWtUZc/jeQU1p29eF8v8jcE1
k3J8h2MDBW4TbHD6k7S4BAk6w5995jXljLUANGOy8FIo5RDIe0t2oXeRf5llInTRyVxJ7v/F3IwI
cLJyyFlrQHvsJV2sIGuuovAlX7HQWJdub2QV+FwglcUD6ho7M/kYTbE835VHaYITtO+Y3uNj6zFi
gNSff/S72/JnCSAm9BL5c3CUctsx+c6QsIAE8yq5pg+IqV4W4iIhYZFAh/J1CsRaj/cDwEZ2qFTu
U9dvUHi2gT7MXB2TOrDTK6fe6vBx1WYTuhA2ZEytRnTRDujrYQJv+4K8sGzYJ6VbZr9rAF4exXsI
R51hYf90UJU5llwF+uqcFwWmcSd0T1ayyZMNU2x8bAHZjLtvBBCwK1wFAwtFdpRqXjyZ1YnX4R7g
7Zp7T38dE8kJ94nQrM1LY/gbGMvDf4JHzTZ+tQRDHlu98ixAiQNn3u8dA7TzgDI5ucHdNxI4vYBH
rXSElGDkv7/b9zIEZdxCtOKV+5/U7RNWvZnfTLPYj5MJT2Fx9VAMRPjRhjVrAy5ZPd4qRoBuAuzB
IZSzuY/FE2XEfL+rCxGhfCfp0lRxqfrk/bkpgIfg1dFHc/JnNgkJobPzoCBl2uBwUcxzosDORRRH
N6ChPh4EBX+Km/PdAG60WcpvTOIKlskk0bHUsyrP1YUQeERJdW+7ZpJosVH6xmAXoNNs4qoR/hvB
gF6vDb5kcxHHpGRQkwlQb1UXsLQ0qr9Yjfa6FZr+zkzwlhnL7BGATrDN6Nb4WDTE0qyLI5iK7e9e
Opaj8iMEm9DXhAqZUztZAkdgxzkExi/N7vbeR12TqdLsCx/+nZEVDRHOVF6j+/IDUEWR1Nln331Q
+dmkrYzUsDE4vM9DG4oxoTuK/LgSaWvDqrEu6Wtq0fVM21XBwF6L323r/a/Y6cKw3wzQ6sp7nCat
uTNl5ovhIeZx8RDwOptS2u7hsyUnjB05lUoLEfsDH64UaMlQPa7W/03qFJmo7GX0Jiub3okTc4/v
ytQbp/FgQin3JEeLl0XAzQh+eX4pcCjA1xfU/wxpHiapiRVwWPDVkn554QbWHIcTqidOQwY0I9Ip
w2dFQyHZRhEH8TMX0qj8K/FPonoxBARDjtD52FMiwk9kkIeP29ORfqFqyO5eiupT7XpYCnoTDqfc
REv7+a28qmvO98wHvAQrVedGy8AOB9/j4VgDcj3bCRZsyGzKJ48drHzdJVHMBQcM63Tg5mI1k/AD
f7SJgGg3Uw+azMsuzIlgkMKsh5ThonH9dqPUQTf34tDTYVpkR8MrCx+1K5km9WqqEe5flEE96Q4v
bhDJwYpsCfe3SsN8tnYOrhBSyE1Ljn/rwjC+I+s+xmRp0CIn+1trWd6c8HdQrDGI4OcTYTVDx+Pd
ACI1vVQASUN+fwwsqMeAQ1phX58z13vn68Wm9EDllFwvjUcDZ6BwEa+8ePFvAQuGZzuOwToc/86u
SRmqMVtRZDIrCWUrru4hbGrJlZsV1R927YIiu0tX33iSdW8VUVnSpbqpbPhztN7FU8p4vz2afh1j
D+KNflTLstnCj4QVEV/6AeggSI/HNn/weKbfcCHmY88YsnB8/ItTczGamz1TLJbWrv8Ub8CNVmRR
OLikpHVPmahrdsVXPCf04qfuwYwYthjHpP4Xbct8/BkkNGLt0xwiJRSXq25i4QZMYtDTXWP1V2H0
2Oq01yCNq2vJb/VliNMtpPjyk8P6nYMqsxTJEOGfEetiqIDVyOEYTB7Y6wkH3wqWEcJ2JLgJPCfL
f+BnYV+a1Z/Khu+UYJkBrHiISFTSNdBwqfDbhLABtcq894aRJ9Na0qUNEu1MCUEWE9uMpVZKUasF
aE1UkDPGj+MHB01PgmZnaX7Qe62qF1cIN92H7STJ44XG7HHwM4xP6VW5apIAopLfnJFGuIpdmDkf
3Fw5LC0xEVjQVQHFwS+zyI/vvaEWck7z/3mCrNU+XCigIUkXjQUB+IGsf0DaXjZwq9slHcMaz3Yn
rG7dUiuEB+nx13k67yZoaRCyW1SahB5KwhYQsh6zZH5irNHBij0o+KCpT056PVjUgjY+eM2Y7EOh
bQkYqKAXSsaunr7t/nheeV7sCmE1CHr/swtuYvphwajbPi8CDKtlQ9ugbsYZzJmmJ59BVrv1MkOw
R2Y/o9FuUxVRF6v1n92DooAqeKzw/FU21g5O0AwkeL8nbyp3trtr3ru7NP9y1Z8i1QFUz6Uy85ha
rV1T3ZDC2KaLv8XdqQseKU18FtKRD3BZlFt05YcEA/UbbmTS8IJEnyTZJJ7xAAL+1l78g+BHdfU+
fp4JJwa1Fj3Ng5HXrrsRPNRjgcTxOJ3unOfjiGqKFRMT1N/+cReebN99T6ZXCCq4jRGekZ3QySO+
CtdKtbozlWxBs5Wm5qw0BTqafSOQMGviAYCsrE9YAAnvI/QA8n7m1EFO9e3UXgKyvIh2yCdJJwOX
nazbZ+S+Kh8rYtohQoYThhYoHE8O7RIzh9floUKPl+p5ivMuGOgC8fsGaw3MfErHOLXzvoovDeaP
7Ysg9L4/D89Jgp3QrWryMAZ5wXi2+9dl22aYPJhDC0jrl18NSKBX1fiT8oZymwwMl3kcP3BAG/V+
08tZi4gMGc4sRhtVO7wPUy3wkYorWh6flVa7ytYgmWw1lRO6bK8W1Ovj9WJM5A0RGoPOi7y+jZDm
bllcqJhy8j3iXpAs3CxK/IZ191LG3H31x06KhTHwNUPT6B4mln8wKJJJ2OfsAoJwbxA/dXgv4tZy
xCJEQ8N9nTp9pVhzyZi8jq+QSPTj5ywbKPOUc/y+bnln832RfCp6OXj90acryMEKamNleqjarcFJ
8MN+vRiY/dvEhtg6muVSPPgjqF61G1zYuZmbq+q2PdQh3qkKDDVAzQEegsh//eLDOcPEnTsv+543
kyJ9htDcsqWGIHjhNRHvlMKYIg5tt2+5JEQB0eOgDSnNnbYm7/m756Py/0k+xv62ciOOH6VTNoKR
dp2jQR99H3vGyBUzfDN2ijKtxGlpHEZ6+aRH+G+qv7femGN2UyEBIKMOubxR/WuxrMkHOe4u1QKV
ZQEPXfcKIIx9raQKxaNXVYmJ0yzUtZGdQg6UPyhnXmSjRPY5KEB3mp7f5RIk/WAzNGhAYHD+xCGg
DeKQfNfPaqKRCI2jA3xVRoI34cgYAKy/LsnrRQD2dElSO/heKI7E+o+PJL9VMO7fEqossTPrW5xZ
1i57dtcsTvq0UoFwtkK7gnNCB4f3SetcbRTtJossjjug0sk0dWMw9HglTH0warYkinQpu8DPSL0U
/RmsdhZeT+q4T+PrSE1KbZBaqT5zp4ctX9imPEGIU2cp/pgmB5eekGoij0k/Xbgy2XgHKumNSPjK
pHzFGQcswZ4KWlFiPoXVrr4gpkh/j75NsPyUU+KTu59qPIOWppk40gM0WLD2x7u3rUzkmhFr+/0t
a+v6ORsR0fDa4iYJUCYnxN7otKHEv3/OCDUzUdHBjs0a7eNCSb7Ig8e/zI7QNyT75MEi3yNTj9Dh
KvkAMnaZ9UytcD/4Ybz46YH0H3PVKjHXxhjUKEWDWzlAus01H5TvUFam9twLzNsljJ0VU/O5ziMG
EhG6NX8OjSK/uGE0A5ZrZ6GNn6Qx9ICDF95+TW7zYn7YTJzQd8BiEOd++AeqXxKLaIxuk8TdEG12
3Yos6BUtkVyGkCkIVurtuWoOAZpSDh+XIRYW1V0yRPOTvu2Jxn0+VT739vRq1xK7SVil8SPQketK
nIZpDqyUFiYtA5KGmhZTIHnC15mfF328xP1JA7ZCd8m/rZsRDdu3/J7v5gxXKbDiVHcfi7TGpVVn
jAOu24DapUWbfGIvlh6zDWBLP0jpubUjOSDuUbwIDZ367zKlIWOR0rDWN/7oI12xyTBp85QpXIEb
7ZOGGJtslIbyusTItcsV1eAFyV4puPOb0XmKVeHR7u82fXadc8SqKTWiqEyqAOyybHHyYiHM+Ha5
uEK3yejb1N9AAcIs7biJjCoQkf4HqH4m+UfdGs8Aov879HGXRt+HoO13VSHALbiyKwo+VO4leOrB
MVnE9NKOq+kGBQF5ZzXdurH0ODb+jnBYcTVXW2qp72xULr0fVb2PkdJ+/LOTPoDShPwD+r0PVwvG
TURHzhM2Zxguipc9qNiDuecNanZBHbWVoWakArdHYvIMaZd9fWh200KYcEHYL2V6H63MtVa13kAa
/PhSyKl8K3uwETarj3sjqX3b5Bg53fxlBT3hxTs3JDsl3PawpUlKzk+kwXkk/U3Ptnlj68VV3kK6
1luMCmoFn+4J142ZkOqWsc2h7/pZgb/FLdblwLN92z8JIH4l5IXZq6uiw/SZ6YnwPTF+R1IMBBTp
4K70+Qapj36WnK/+iyraqo8iW2rsR2EonwxPo/6jyoGsZ/JMKsRE2pnz9wkUrohwHq9XHeCR57gR
HWy8RWYMphE8TMuDF26SpSGa2EKAwgtcmAoiyJayj5Z0kmU4RVeQ7/v1Z2qXlvJWg16/GEvFzJ+E
zqJZ2GxdXcFyxrOgXChJQW7YqYLMvwd6TTvQM0Ymu3+O1Mc+Kdmw2CVfYP8+OsDkXd3mLMgf/Uqn
MjbQUTltgQwLLyDgr2+ihtEbf9MfeSy3UpRnjRiA33QWyUpppPFVdnsBvb2kJd4cSIIESb1Fk4Ed
hrGQRL/4XMyCQXrem7ajAf5V+/V5U7DXOS4KcJcaUz7PEjGPOOFfTQ1SRepV2Di5GMkgy/W9CO5h
WlbQGop4IbJc833FYaWa/9C+bjJMC1QZofmvZkYkU/fC7eOg68jR2xoQH/3k05pmZhXfg9mUIN3h
18BiJbLGLSJyNXAUki1iYRuG2XMsvBnKq8tbttqOmwLlwZSB3wrJzRKrYwK/FhkL2rckqneQtX0f
g/P8AjhWYOTGOXxmB72pefHyees9fYdYayptI2R3PHfVg87JdYvfHJhN9rasvJy/b7okTu3xHR2B
12L0oJt6zlLhPERFvh6FgYlfs5qO8T9nsRK4NZnqg7ny71nV25tm4uy1cWVFVM6IKUPC//k5pDx4
aF2K8/aU3DVINh7qELaiOddOwOCr/j9MKYRAuHWNA8rODWEflQHj9Dcwtd+exXurGyGTLK/29mOe
5gSpzTUAnl2NoXFDXrMcdrcFLl5BW0zogS0Hn0CtPaZ8+esYd6CZDNMj5WRgAt9rnjIgrhMkdV9r
7sRdGpfgq5txjkUQ2ztYPLFy7ibPC/3XC57wxps15xktHkN8BMnM9mwVdCy6z+Kqs6396QVI89WR
qC7mDFsloUMsXgChYkYHR+xUVISn58DLh62VFArzmz/NVU5psIQ8cDEhpHIlbCtsO7bZv68Sr7hW
O86sXP5I3PvESFufdFhoRfvUhWYRbSVGrS0Dziwz688FIQzwBlnbDvvHhyB1D6Lr24h31M54p315
suI4ltUubvGLxRBmyPS/EEDgWkk0M4PYU1roIiMC95VybLwxht8Ejlgx7G/xOU2C5NbKNgiKWkem
etrsAhMuz/KdU2JTsS3My7wPpyT12jjFCgEAntW2Tqe5JN4SJIs+k4ausXIkyVjS37DXH+T09Sv8
43sM+dozFGY/20gCvMTUrR54I2hAbWrJgBcIf0cJKtCgbMfFaAk13cx3BmtlA2yXkxrjTjlbQ8Nb
u21ko3iuluCqh/iHShdOXLPYi432Z1uvrVJhMK+TjDOTEFHGmnkafr67bFklVIAlxpNg6lU5Ghnd
wj+PsCnDTCzvmmiI8nKSRQy6UiAjPIdfS7gsPU3FBsKRzYgInTzZ9bdZwz4xs2DtdYi0zty22a04
4nTiRTDvXAR4uf5NKvUG26ORp5RgXGTUNJ+dirPt5zkLiWTLdDpD8U1uZkQ6WvdrfxJ42jn4Vesi
AxqICWCqhlT+vQieLWZUiLM6RLatpg+YFShtirwKRAO8N7BJ9fxVaLr+qUlIOsh3f1qBQFgY8dAq
rccMCi1dXKo3vpXkX0SKLkPhXtu+nWFciff5Hq85VS1uQCJhuYG7d12nk6cjAflOa4blELTdJ+l5
ea6MSKa4jBfKBAs1JGwLNIw5LqJ0cmZtTiOe3Ei1xqt9lZBLG+Kz/saq3WIbK7TzhHuum5bPL902
L/bjbFvpuJIUgpRY9MxoUMxW+W437huIB562zA7CZiiecYuGvoLELfwhLcOby6pG7xCeuZHSedoc
06Qh2gs/WkGH9ZS2EzbWnTqjDPG9GjI3TkioscTZ4kf4D7ZBSxcA5BFnk+wn/kbanxpKc36rU1ub
5tpmZFLIzZ7ja6c5S5dxj9Y+gzs6f4UTKJAiwRkWWKV4teBNhmBB6Zv8i5MIrOLmPWhOj3EZPgee
ltomZVH27wS5L7vXXnPKCxyhUfZhp13CyJjHK0hBaiIM8PK1SXMudJfugyhC1LRergtlR0LZtExJ
RNRTEjHWlWCHC9jTQDoWxBMXh022eo4I75EzthlTNLugNEKd1EFKo92VpwQe3dSS+kiyR/LDIc81
efx4Z4oG+IK+3usnKnHob+N2Yk0WPJ24c6opVeF5qHBaSXJoQOKYB4d+AnKG44e7XjILYLb+MLD5
XdbNNTDF05jJCShxp2NawgEkaPDXQm/UC0QqtntMeoFjmKajfSJusNkQQb3fQYIfZYba02OLd7tM
suSXY+7Q8RWqxIvAJJulGAA+ee1XGHICCAC1gCidmiFYvM00oK2njp0orvNMAxs8yOudcuci3F7R
SwpuSr44C6jhYenXgSBPicJ3r+wlOS+AdZYrwNtbe5HbvkydaUTruqEHEkFgK28UZgR3hrKXw9wi
4OGlrc6HRhiqdQIc4jFRQQonRakQushDz19RA2CS80gCBobfgUQnkvxjsR92iKPR+cbMNBCKVhYO
XrSqj8psuXFVTUM39ql3cSwGHuwD9VMGSuVwDDmdfVqvUBFhySQZCpObXqM/xWyEcI9gQQsRFp6I
26ouDs05t8PsjpWZPouWyse8yUCFIaXsQ/HM69hpfsApILpBngwqJ0iZ4Sd7QVwqb9eVaduIZKwP
ec57i0EUIMRGXjojcqsr/NlRKSeywMWI8YpHCspknyperJ3PzUVpLxRMObmEXA1UMtpicGq2uEyD
1dD5kM5IMcfjN9eyRvHSZlwnjTVvjew/x3F+X1rumvCSpK81aIFzpRUOKTpoWrwd52aylhqRG2ah
DawIY5km3mjAJ/RYnn5Z/tJaX2vKiTy5xZoBzwb9+p9hDN1NV8be0FtG9077Ua8d9ISCVe+7Gx5q
8cp29xPoe4TVJ5fwU0WSqaVffIdFGxEOim7e7DWDyW+YTCIVoOmHC1T0lo7CVyiAih6/xeS4yYEt
oQ+d4sY3FruO++NhkKAcWN87FwWcuzu0tsxddBudZkqtCsoMb5WQTENdHMZn+kZXQkcmNT03id00
BVMpNGO9dC4Pbw3RM+0oCTJpos5B50M1nfOxVyV6SJbDj9CmeOtbczm7AeYSQPYLy9fo7r8UBmun
vB6usWsAg3yiL8UUMtTRDt6gmGHwRXel+TNzHgGYm20xpjlyAwFm92iLgz/Dwq/qPnHykSODdYGc
Q2SVFe6L9TWMreGq+ERwRUMhd8QR0LG9XZ/jydvem2E4/dvCz63AcqRdxqHUTBh2rGv+ZWSCCABf
p53h8+w2TQS5x/9CKEyEJHcnD+jyouScCimEP2plLx1vzzpzvDDvE7Vcwid5a5Mt7UohAYkYWEqi
yCHIlqSbEl5LSlH4o16StZK49ZVESQZrXUAE73GFMnEGRmgw+lsSen7zwixbpzeWXnvF9UCu5vcw
zf/59T/eELDWlx0muBNNXke2EPH2iAtcfE+kKJW0rqNe4UbI5NVyd7eLgVoRxmJSrlBW/BPxhB/v
3PBfoGJxW9usst1swlhAbI936AMhPri0VXynWJMPx6hJonC9nKM8IHhbyeWV6Yuy3AY2OJxLxMU3
OGu/plSPawHfY0TGBoZ2PGaH+psZbnOi7bNWEDghiVTYNP02a6djdSpOzD4x5CgBnDyfvX8kzOY1
E2c2DmBhGj0wkBH0cI9XElgwdL5B9KhxwDYfv1of+r7A0HSuZtk6TgLXyEWF9NT/jfpIqBejaIy/
eDgleIMRhvJCUjwQY1cda3ybMaCur45Bddg+EftakZeKfzYsYw4w5Qea99fUUp6YqAqShvvIwy3P
WvcDac43iZf/5Gf9sXLF1rDGPZD89T9W3hFb5+02K0t9ap588xTkiVG4MaM12JPPX3ly9+uodUsF
yLDhqGrJTJJIYZf8kL1D/e53HcT9CAeXgglMYPtiNv+UE3yZFKoxBlAMjVjuk4v2Azi0hQXDFxAo
Pgp6pzv6d+CQ5aRt6sYfnb+IRmHYQexeBf3mwYp6i9CZyhby9zI8r+DVrPGw2cq4ONHrX8cBdZvN
wBifBVOKX2CIbkpFB/hOvMDhiYaqQlLJxhb05MyvSM+5kcJKJDrPlp0ECJQlLwk2G0fj4ANW+1Nv
fKtF/wKUHWWBLoOHIJ2RJsqO5WOdek+rkrrMkbOuoWeQEyKKoXSkojCSnbOatM27/BBC3UBjcluY
CaBxPKun0hRwAvG1ZZT5DnMGQsTU/Hl1BjCocM/qAcVHPL8gDiV2slgcblu103bWFr0sMunvzl9J
LBgO6O+WUugIQ6jZ3wSLxFeBE1p7Dk3eywIodVEB45N4lx0Y9m48pJ5ASCyyuTSdMcURzGnjyVaZ
YCRFMxmQsJIOvp4iNB829k90hoJ7CVL7VU0y0gG8IdOY3QyJqUO/4Lr8ni8oVQOeDAkPXI+8f/wx
GJNwIU6bIG4UOorjZ65EOj7rCd4nxYDaKiYVr6bToFg0mtC4CCoI/9LUG6Z+D+n9DFOZ9MfmuCmo
F37ZT8bkw7D/agPCCo6t+i2dW3MjLD+IqnZanbIYLdcPtmr2FfeG3fpI8PusmLZY1sGqmNWQF3c+
Jd+nMuk2wJCnISPvWmGPh0CnQH5P3ykjtRlO987XXq6LX/HNhJhQok6qQPEVminhKroJm/9F3dei
tNljBCWNqVT4BvLhKv9muldwl1S3e+gIBNxOylVtAtM508YvMX8HBv3Y52hq2H0IbWqjwmGtZYnW
4qTGeLCeApil6tnCdSCQjL1qdeU23IoJ3bCpaz5NSGax2pkzlwRAJfXyFtYOT79XZ9ChIBDB7v0r
aChwGS5IFXXwyFhEjzGUSUpayLHZJQNIyGdncMS0jxQRL4yXJJhAYPZSSDZSX36l4SEl8wzUwOdJ
vc8Vc3ZofhyFWnT1KMZeIGhkBBs30pBNXnNxeUeDRffdp8RP97giqyNGrd4ZDA/ybxVHpiaqSePR
Z80m5LpOoqsuORaSfMhwcQoixf+gI/RuorEUxtv3QdlQVU7lqnDn19MmqG26m6mWigI2ExGSAWEb
l51mLSjw5lQvTfpnC5KE7mX9orhZY8JEeqif2yR2RKdci2YjlkweZLiBAWNlkwBFtg+iKahC3zCF
eUoCK/zl8YPBxAw5bywrbBhOqD+fm97rkH+CX2dU2c+lM0P7k7rW62AEmf0bdSPp4omkLFrIMQm3
izJwi5HdO4oNv5sY61p658sLgU4JKEqWKkaItNIlE5I7AcGeqPIJoAQvuM50aOdIPXOTyHE95MOK
wuBvjhgCJEnYhKDBVR82A6AbfiO6fBu0o6rkdE7bX8I7s/pjK7M6Mr5joZuMgjKNwH2xbtH1YP7x
bndacTEBiwsO7iv2I+BsjpT9DQ7Hmip0UvPzcwASdKNWi9ODxtZrdhiNGWAI4kDfCNpYdNm/jsLW
kGD9Lb9nXTGWtP0vd11TsQ4SKyjVJdAekanPq+bPPIp49ArVfWhuPnfgfZRN8Eet6HuJtWiHUVeN
9Yh0f1UG5zhGH9jj+F+CIPtzM3QveuLHvd5c9MYAucGhVzR7nbENiS8tTTtV6FiNIzCh+zyrl+n/
OWxyrn8RjgD0cPSZFVRYYsgedRsSNypeJcjLMcoRKR9axDizq+ogmL1+WJU6wCCvclhEzGojXS1V
ffoR5Gbeqi2EN5W0xMVzkObWQ3me+Qpm9rohaCxcEA7pYYrtfft+3OIJcjxxjHQJBdsQ2iH+bUmq
ImhEVodQl58qM/YRuIWgRvUc8unnX+xrmJN9WV3kjmewAMzBuAjGpKBqsblomYtUUIlYi4W4rmwo
DwrpPH7CZc5i4xSpxVFFD5POu/IOUywVz6QCsyZ4Bsvnspq+6sGyMfBYtbHptw3f7USxt6sKKpR1
bqXYlXmNj4MzvkmfhJCLIzW5Z8oR88AVMzr83upRIUnmbf50ipyjTEHhHzn4P3s8P/xK60ezUXZR
fBk6uQQb4cZQz7BkpLNVACXkyRC76k0vRTSi/FZBL4JhSYvoTKBbfvPM4zyHNodIPETvtmpcFqd4
ufzcqIVoFjdzZpW5g0Bd840NRTklQ4V6xFcrMk0M77okKFjSwDGN+EKmuRmJKg5w+uCLRlkZwFce
BB6k08Qp6pm3AVKSw90blkVp0zc7gMxpokFXlmMk8KvhHipWb4NNSGFb3RqiOj/jnN0jywjEBfG0
SkK5xbGjrQK+vVqfMCrum/Xz2oeUkJvrVkcni8XOxefDUQF7UdwjWnD4qeClrSN0hvHnuIb/GYZ2
TlPtYLMYLXE0lbQO6L1ulb+3P9TlzyqJUm3/ufLnhUIUWHoO1b+bxAtTYc4Ix/mFkVdQy/eMWi8O
VJcSCVCx1396QJtkXdMumoXu1ZLe4yBOAaATQPW97Bj8PFNfRLH6RbkXDqqHF+uTLGSbqbjmbRc5
YDMJzCRMqN0Vs87Hx8FqoP6xmwuXg9oBQ44dW7vzGKkyDZ3+UYLPfS1XlKX4JBQYL6q/J/J01CmY
28Q4FqMPSFbbXMiiKY9aUS6766lzEez6g9PQXtUPnPXvRpEDXKzSSEQyqd1foI+0mt39M+rlvgac
BbaWkMMD5TVs5kddsWm5ZIjiTvMCYGc2HKKGqTYOCNQAtRh8dIEzCcHNwUWewLPAQHoFLuVqXllE
3gz5uRSh0wE3y+PoLTudXcNvYEYIm5FNNDbxRR/j+x6aoT2Mu7UMx7Oghbp2OvGM8Sw1jGYo+59R
w+BbE4vmK6XbUxhO9CQCVmf3XEoQT3SgevvNKlRb5s8n9oqzweYXRggvkrh80Ab29X9jgbnc0wp4
diN/DgdOmtotCK1xGznBHeSsiU6cVI+TtFhaq4x9wQ58zL3kU9S7RIFKEvoaWiN7vgcKCC5a+LG8
hEtBZU7kCphy7jKiXruItlqq0PXw/foFzrB37LaBM4oQ9IISiwfgd7UOYn0LOhbcN41Nac5tZEc1
Zpwc35znNmoSvxtedWNhCSh5hu3Qat5O/oc4iRStrCBdm5oaJ7EE4/5rk1phcp5m1YYCZlaDErn8
vBB9mfS1WjbGGm7YIP+tPKQ17PPwtccHnpLsltVnovqG4XZN2sFShnuVz+WFUqvO7pNGP82olVHn
2+epB+ZNC7Amysadf5IhOvhWT61UHJf1wdwYc49NBxS5AQxxyzSE92WgRs/qBwZORIOSDC48+5vG
B/gzvZd305YD/pT7DwgWD2MWLMN8VDid7avHFQZuzMkXM+4IRLxDWdGt/mr9qtbTvk1xe2XAJRlU
6CesgbM4EFs3hp4flRupXc+ATnOnyKYa7skOOlx0jCSOIqhradrqVcpNgf1EDPUXLnTjZ4bXp2ZZ
r+iFoW7zKRF/jNULjaycPf1q1Xha1BsOitftnxtfd2R52Rl1I94Fxw7BBHZcSSjFutXze4ppRX6s
XeGsbUJS7NvhmIYoHhox19SNNFQIqsrcHEcz6wTHJhquKGTzxY2ckpP7LXRihj3145SNeDisAQU+
QNd+ocp/8s45j1KofC9zbSUybrcmRgu0GXbkxmQrQnyV1MNmAceRRqH/KQDoXBnBduHbdyls21Bx
dIpLjCpv8+B0ofB7Iqlpaw+2+cqIqY6VcDxuOE5FBtaVHfeR15UYGcKAve2pHQI2tC/BxkFKuYYA
v7xr0fC+cduVJfgcw1bpevFnp/AF/aiOd9hr+gerdfE4fES77QwVnEWpswTOUBfrz/X9M7JP/PA4
ZLITUnB9PeUFvwQ6o8g76k51iyUIUZlFBWs7YCyuYSaVXDyWhsx29Q0Y+xOUGyWLIsZRF25HahSV
8JKI86u76+WfoJ+lNxhRUx7ORTuP+kI591DoYpzd4ZZ3iwB9lddPlXhrhoqfaFYk9yIycdLlq8WO
B7lZpGDo7hpQuTOsHhom4/p+ZBVsaSjwHingDt0p/8QmBCMPUyCcrhUMzAq5a/Qi3dz63LPzOiZW
91zCJDkMh/w1dTlg8wgnCF9olQxedmmekOHzZ9JR5maVq1LM9IlL1qyUmjtjjn7nsVYrC2etW+Mx
WgtosqsTEsWBPAjkAHdy8LRrph3G2kzxsYm3x8T3wyLPFOKG7N7Zrb0lTOYlP3IiW9240XtrI6PO
w9IBi2PxbXiec0HjD+7DKrEQbQhM9k+HYRv6dAFNwQKtTnEPdLIMIlhCSNmaNhxNWjLtUrbsjXsl
evHMlLdCjsHlfdUXD+coawGSfya6HBCCxlO7YVl8XJvCSR1P96DIbaJSFzmXSZMuWeV0CQN0m6hi
ENTXJYnMO/a4/ZiYel2KF9aupPn47Ya/dgBNQUL3WFop/v7FwTeoTIEF6SFbWQR51h9Nx5reAZ5q
aF8rMbRIw/IpBZmEbEDqNTd3t6bJEdkhv9txx2LAo1FRtom9zttEYU7JrExeKK//m0gkU9LSPcVU
48VShOM/XgGq3uLj7sqZzJsOP6HFTGWtRm2fuArAnM6cj6+5c9zfWfkUBgYjq6y7wiWvMR/VrXLf
ix8Iwbb0VANJOZTcVWVAxVsZsO5MKtbkQF6S6IGSMawOki84hmuMhwpz4r60Udqib8a0nN98URpI
JW1eCvL8FSBHP4CLPDT24GDcKjAG2cYeWAMhBe4zgzICjOMqDgopBKAK7GnYlQep64HBg3fRpj3+
i3B4fGgwPSl4cV7FHIdmvgY7lX1I4NjyPuJ0lB99an4fJQdH9dQhLcKMPjTXIfbYHMy9NE93nePU
bg6tqvhNLUoHnGEDbU9JB1pqWUIWfsSnkTtmztKp8BPiDh8vstFJt4D/ys6GaugnNPJAuPC8Clh2
s5vCCfeifIt1vMpyYRvKbEXZprOcjLnu+gitrbEsiw3EXevqaE66u5de+9v6DF+IGD8g281drZRC
ruDCqAn8XVfMI9Zt9N7LNMsNeE69WuQxCW67+kj3G2QOSlGSrcy8QXDZEES8PkMKjNsDCnuXsE/R
EYSf7wI77CZqZf4z95I1O1tPKNds7rV5dZ9f5Bwdm9GbQgFPRAQ1+YQR1pLWJ+1VnSX4QXS+a5SM
1CABlN31f04Sal7//KGW2/UWrffyuV2o6MosAeochlheZUSNZttjmZy6Wvjb6ahzJSi0qRiumcZ/
DXuUazPTgx8t6udL2eknYDZOMPnOCDXIbHWiGp4hSJVYiqGDQiRxfJuVyIR/b/kea7y0gMzGPMSW
suRi1nfF+/Rvl0yDnT+mA1TpHPizUAgrIP+2cscUMsTFhyWKvOe5ZMmdAuMZIyZawyfCR1Hm2PBK
0D3LP88ihQ9H0pwS8srDJPIAxGwntF681caW/k1uWulm3PFQUX3HwIcYaLzBrQf/JswE2HQjkzvj
oCzul4I5UU+0BzIUR74GhxUAdF/IwUHbIkHLrtOqPZobMTvKX4jtP2ITEB33cMCa1Q5XLGeUesa1
Z5J7n1qWKGS2RnNWTmDx+kokgzdd2fohO8+zsPOPTvYrblePsqjyzkW4km6WdmU5TwIZwOXDZVhZ
cqYz/VGvs05GAymcpqb8rAgCBChBxfB5LvYRw2B0p2V93z2ZfrB6IuYFiKuvk+70rWE7ZWy4iPWb
kwtogZ6FnejZmx8ZrYRepkyOfzT8a3618M2KFNLbTvKdBXnn8Y37Izl8a2HXdekf2RBKjO8IJNzO
Qjedt5yUBVlYnt4xzL3hepRWzm25DYGz03kBMo0Of7faEt3gHoyNGIGXlOHYD0rh0NMhAxqIA/2k
/uzI2GvJkATa86jsgiqbBQUa10rLBad4fsZ9FfXwlpqBnngH0f6DTkpBLY8lJLQ0dRwfrUDaxTcR
OnJfNqpiC27gJXpKtQyifIf1lTBOB5PhdiSrlh0rGoK1rlPnl/apPfUL5Pkm3xRuK5JdYazvscnJ
SYgXy0wr2lDeNiqPb8G3oAKBgO7eX1LWkMP+OS1LojzmwmHH9PSlNcQ/1kTFxB5RgRG361L9GPrA
rwOZO9zgjG8/KTGKvGLBaA5YlBaT+A4i5Fl2DbHypv5XJjBnQoTssRDXXVZzdxEd9ZmjS319pF4U
6uM5vty+zR03VNDNMM0TpWBOfw+yiqYuHyZkalMaoievNEB+M45IedzdGWz+dQsFkUhiemHfFYXZ
iPx8U7iKnYbclA/0ML3Vx3vFDZWuL04mmj/C3FS2IfxQPbWzoTHUz4u1M732lcR4FyLM+NTxSr7+
fflB393V0DMCtsn+hKJ341kG52HuF5TLUNFi63Xk3/qJCMHEeIl9N8Ik+nO19uIV2xJzRzTtMJE=
`protect end_protected
