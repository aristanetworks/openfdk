--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
euHb/s8r2MEK89yHSk0pCIibjjbHRie4F56oByziNr+wogL3ir9pmTGBAojjuNn5wFztcuqWjfbr
GsgZaz59916A2FBU/A1GgG8gffF1vOW96BHcZWzpu7DWXWlSoSQsxqC3Qso2wx9wmpdUI7YEuHDV
LOKafc+r85R6jmjaYWXj9oFOOzhHEJXh0aYytEwMb1HFi69s8fUTnrhEGs9S9kAZwYP1m19MTTNf
EbSFivMlJUvBWhSrkTvrd00X63yMZ59LhQ+CThZSxdpsPuVOpIG3s16g0X0EYNTncAxBQO8H2p3f
DhF4MmYMhYhaj4RRIKbmA5NhcUszvR5VQQYfCQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="W0C/DvJHyZk2WZ5okNjvd5or7Ql+CLm90CohTxbsfec="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
bRGdR6nLedMmCHfCr+UNHk3MS2j63LlADimQlFF5oZGkzk2SoBpXFH/xJof3qXEOvjTmsV05W5SB
Ze0z+Fud0J1le+TDsx/zzTpIwBaYBXK+SGfElL7p/Uv42sPkAj7hPTyz9nIz7tzzuW3sZnqxAAY+
LHu6dMBXWyYnyFfVR71WYZACcF4V2AKJ/yuU5MCD6wLs6Y2o8EAhqs/xi7QOmZ3nJ05+QW9wCGG4
+cnF3vR7Rb2K+5R6JYnu6j5MfRFxBWd2dijWCyNPPSj03OCTguyazwQE6dCstt8UcJ2g2veOR4CJ
y50yoG8dO4eEt0M9VnytuU8HPy33TOlyyofnyg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="WfAjOBvD6mf6Dddk8lfF7sgN0+Iv/8DIzK6JoUDmEQg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6624)
`protect data_block
Fc7uZPAy53Ro/OaH1p8kCxc4HPx8r7mffmWE1gashGAk8OecR8miyq5yTHjBwfhFj98Z8zxWtX0x
kI26PNAVy5HFQMbmf4d9eJdZujEQpYxeZeACw/PdPwCRtYc/CccI4Ui+429A9Sron9zmmHhIpgn+
ejGMe8pNrI9Q52xObW8+AzsR85shcZ4r8b/LyLuGQqQXBgL5zGA+pFoCsv02cIR2OQjYrNkblavM
IIL7b0XdloCqn5QoxD/zxr2Z7VZ5JHQQsQC1dwftObfni2rGjbbLcKT0XFdkGiUqct4KjSx7bh84
tZlO83Cr2Fbv/s8ibaKWIG2BCEDAi+lb4BGQZuM1mY6V1y80nWrD692nOQO7y2y5uOPKVRsgHVAY
dBvE/MYz0FM90C9Q86XorvSyphesWYgEEHtYrUk8lN+dS5LMc1IWrQ5uZtlHKiHDAhjksx0ZT304
1NgZMQXyuVe7+YdIlnKMP/RWFawLMCsHZxBaoZ20FAEXyNE6RuxZnCKa6rMNTNlfWrWsdoCZvwZQ
p8CYF1g88cgOynyLbRjONzYtNwW8Bq79hCCacnC2vd9n53vrSUzQVhncewc1x892BR0UVe1zFRzj
MNnRS68y5KoSghzgZHaMK7ZgnJT4ebm51zmTaieQf91gCNEuAn7ersRu6MR0OmQk4iXfARvf++K8
SgVx3sqZAO7ch3G/gqdSkjS+zOeRnCDNnROJQnhHT7gs6CZppsu/GFRJGIsslNNH3IzMHCa640cl
1IudKdMtoapiHtiWMO73h5jR5hu5KtOHXrCIhlSsLbxz/KGpOEq1YCm6ssUEQCRE+Dj/0zZ1ZjnZ
oyyWtV2p04JzpvHst4Q5/oGTQiqY7M7cJczZ7muKEamDAAXZT8VjfjNGX8zFfFFs1JyhlLoxdk2R
sDehlj7C2hKHDmZY3jgMp0pHUq0yZq0BGZPgZZKwUPCfe6Ua3VYFb3Qh+C5M7LZBAmm0O8iMVsss
UM+PVZuDVIT0aVq6LrFEiaMf4xuvfrZiuZ0YKXXOM1Cz9UG/a0LId9TSONeBY5TcYhnS+G/8404s
TruoXZmhiULPriQyyl3TTsK4eYx4dbvie83EGCILZkHfjzWyJnATxHG0jmMEjpALE9wclVEcYPfu
wSR9PnNzjurOBsA6rvvKuP3/+72E6O0LB4fJ/+3tDszGD+P0KQxrI931N+6+nRxrkTkRo6YpG4HU
oWD3Xw9OyvnabSfzNagBv22xD5Jx8PYQjA3lDuKqxP7Mppa5Tc0O/P1tHl/+9DmQPm4E5QndiL1g
CeMafhu1DgWGykQlj5IA93a/O5N34DSiKQAK5zCjZdqSdEEXunXZSvt0SCRHI5eNhjK+glT1+OJs
K4zpyfeU+12RbTOjNAQeQr+cWd02h2DmEITSbumJF+FXHW4OnYMXDORXZ2vyiM5+0jr+59wgbbPd
ypp/RqpW6om+COIvuRSU2Ml6D67uW3fZDi+L4+Ra6P3K+CjtJAnTfmYnILO8574SbRWn8GgkkGgq
DVLgCOvCpPwdWrhW2Bhj5uCUk/3ExRYjX5udcD21hgVExZI/SjPLnF7H/LgXe913CRne7bF5PwWZ
uVoqGt/DA8Fb4P4HFIfO4keSOpUMdJXYmij85QbtLqMuK0pFg9gIObF7TveSHX3ASrJFWS4GQm9S
DB36eyFBKOYaAN+blGSf6nE+mG58UHsv4JP9SQmOe/e8mApGxTmkwgdruosABr7a1XcwDAp9h/+3
hmM/6/jqXrGCNDyz2Gu05maehsGLzJY2pQKOQ3fgsSNThHkZUJ/mYeHc5NFkoedFLb1PuzZlUtzc
+Hbq03xCvgKZA09vGCdkUlcidBqVFweisLu+4+ACRVUX0Xbjc6Pfi8L49pYTRowrrpm+++JVGB0d
Rzt8ErD0wEnhsrOA3KeESiH5U1KsQi2butS5yYw152FE8fqC26r1bjTLWhykNZDN92S46bS0K1TP
gN59rIOjzRvf2sHu3v21aYOhu8C6TK23UIIqbeR5I1H5bhgM3iKIrgCBd6h+Neei4TsKCGpniXSA
omJVUgLHntwRD0S6gVYwOfEjwHoNluJkzDP6P01dBLz0lVAkbnhgJR71MUQ2fKLaeFaJb1CMmEMM
/mVHJUxY+Y03jPbgHK23IXhQuf9I7RDoyqK73FeZKMTNz+M8aHs/hQWhUGERihRDcqyxdelmLaH2
vHGg3rXEAA31CdU+olf2HFMpbTDXSA4CRDBhAeLIetQlb3dJfxOOpji3BhkBdmThGbeLCFqXG1Nq
uuhnStTJsRvr/y3fskg7LN0PtLuViPKpXMjwj6/y+kfRFR6rsJEju/66wBeuOdwSxnemjiSw4kUb
itqPRFTivt/fM0dEdtK7unJkizbv76Y6qPXD/Qz6UnDiVPuWYJn8+PNOK4Ju10dh15rpCiI9QIIk
IQ4Xpv2huuysQLKdSyfRzHha6k2SvyU+BUnp6G7lLNlBT5mqxDWckl/n0DXwToblnjL8rYhInPsQ
c4kF/rca4ULIGrGMQCglFYYT7mQhbyFlKhxazDRDB/i8Yt0LZgAI4mtFAKiccUWVKlNiRUMr+nke
mlfGIXdOb2BBkL2dxDEnew93CLEYxgH5JNitWd1RID1B0CvCU8BNoNWvP50nNJLAj5hSW6UTWf1d
Aoy5FwGkgyI1nHEfPYJKE29NpYa13dnPbGd8Zh5kfmgrVxhK9xRQ3r+fN2WpPlVP0jPjXiBgIOkj
fJSJqWQLIURe09FQyx6Vj387z1aQgP/oWatmvI9D/AJ9AfQ2P+zEJ/nKB9rr7rOEnfWM5oAPdcIW
q1chW0HtyYBUes/ZswJQBnLB6OZLTcC8Sb5NcqmxIjAMD1vJSh7BrJHZjdawkMHgESZTHs3e5V2p
dBVjsPZnyuth4x/2iOOvh7P60nkfu+k43vENxLmoaHEyu6lknO92AL2cWINh2xD0xzAniwVXMM1w
6ni075E97qbiTBYuu59ISIXW6JuDB/CsJSDQie7YZ0uFOhMQriinF2kd4R6z/sU1Ob8gLKExJ0Vc
C15BwviQlzXxd2a9aluty591ndSW/dcAu8Xy3C3gygOvvRh04JUq0o3NdIKm3iiBMFGfDIxT4XCV
m6N2pLFkuuTbv7z18/sdd6jNgSVLx4cZ9JbvntWBdIM7GiP8Zs0flznvmHrqrjQShgeHBaWfy+zy
Kt9ZLxsimgAXqcM8580fg9SbO8gyqo2bpqFf1cxbqFwwNHB4/tlWthZGenq0TxfEhKEx4EWD82Y/
yYCq5cVI9AYfFD1imnJdqqnodHxUfyTWHZ4In0o1Gy1Lok0A/8qlwATRIN+1rISkTlYH+uAG9Ndt
5Rtqf2qHedhXdVPaUdthXKkdY0TRnKZT6s9u0qdd+bBCTQA+GYsEcOOhJRCcMY/W8a9gYxn4O2hn
h+LwxDktFazvhaDUYPyDPOjuXn2qyVAJpIvJnOtVBePGiXnW5yrDzG9n0whluviUT65/oh13/rgn
GDseisLjZDZ6lWM6/srHwhgamFk6Awcr1OAh4yyq3kifD2RBrf4ox0kWshMUh9MG9SQ7cBOyW4tB
3cmgqR8Ll/xOjnbYO5TQrk3WawU3AvcjcP3UdSQiKbpn7eUtov+OecY4r5K//TN9AVbWQ6K5bWYi
1E/5jUTjtqMsPADmGNRChMa5nCc8Xffh0X2STpF0MbAgA2I/pCSIE0nKoWmY+QC5SttdvRcU8RBB
xl/82ZgseaTJea0fmcYzkqTCrv2A6CStXpuTKU9otNw1dtJZHjn6iVTxCdemZeBjGfm7NhlH5jcc
zKnD2l51T5JhThQzVOvduo6yHTPD0s1ySoBIVCtl9AYTlSaWgb4vix6LGShZnD8aX2nk5ZvNrPmf
aTrNt00zpJHbRsXrL6/nH1UqflYVmgrW1FsFN7ngiVwvw2oNTDj3QCwzx4Z1blfxdu8j+HvS4JMo
6FKlI89kmuaMZsst8JFQDPh/EtG8AgIKmILPRT1syh6qvehj9ZsQOzXYjvTU0rUwbVSr1YlKQk59
rn43jEM+bp+B6GdT0BVQX8L58rFmmv+vYHUmj9uxi1yviXwYeerCn+rDlO9FSZ1qf5vPrihEInZX
MwDqCUWhQzNnSOcz8HL1DgvcM1b5eUY5iznBRdwLjJTCLtBZWr5UWC/jZjMy0NtVKllhVtCABhVh
jXPZkVsNeDX1+xcbnguE/uVUROx2MMQq8auKBlKrVG2kym+y0uN9HbvWstG7mlWy+Ac9R1C6WC5o
q/4L+KvyrYa80glW0XP7xsTqxYSqnTdAu2iwOpmen8QlzVphWqvFVB5kyM320nzSd+nxsdURLidm
loP8rQ9Gcim4KoFlQcwp1zu7E7rW9uMG8Z5V3sbmdqsIJ2PoF/Sf+zqyCr/rUOrwvKfoLS3FyGS/
bci7ZduUEp9ETM1c2DowldIqeWzdntjSb8r95ZFOBK4ZzRB33suOuY9fDRG1wNgF6c+zxy3q/uSt
9uzy5ni9rXb1r0LiexsoLPb9VaLDyg8ys6Kyptl/6o7yeghQaAm0WTxW36feXPtjyOYx4XYRRoOY
uf0d6Xdmer4kMst6AhydhL+VuR96nRBJ1zFdPq0yF1jFuNzIOjq1dPo9pfbVCryIL6g1tBjrSvPM
og2jMzgY6G+28Gqszb9RScekIUzeNbB1ph4T66x9s9w6bWdUUKlZOBu8Q43p86VlaqqEtgTLbcqs
GinTCxkhP6om9zTA2SVVecA5JnuwGNajfB8JETRQmjnmSKncp7iMavXPGs29BjdCwCcI3zBmLVH+
0Lzc4PIlaVL2pIhWPkxeWaCGqimAzF2HeTM3O2ELzXxdfwpqaGXhd3BFHBnMmzJKU5pHGOIukqXB
Tqjwdqi9L/srSmBEFdf4P0Klj4IkFjsPA6JDjuRJckMr9yPjTOCXG5ZQVqNHncDneZlnGd3A6+Lm
SnXKjPXyqrNGIKUIbYLqmxVznqTDch6BaQ4y44AMQD+yXke75lRop42z3xdI6Eo66+k4zWT6l4+P
5SggzYYmTBx8pHbQ7pxAkByHrEikF2aYhUN4y9xXErOQakgPX1gFmgEaTyeEZh9B6OhhHxKBB/Y6
zXXS/1AudTKZRp2OW12rqi1pA6weXLlBUSyimvvxePDaGkmlf+IBy5mquPVD6/f2w7WfuwbZ3C7G
Pmdj0b5yuOFpO/fRYXske8Bl9Z3mRTk1nDGNGWpE//rdvYJyStWGO/wxcy+SYVes3zurhkqTFEAU
h4PtiohelhpNflw6pXr+9eL3ARvWAJKgC0rne35MrZbuwUu01kNR6zA5E6Znfp/X8fCYecuZrX7v
U8SEvuoxrPvi/tU+COlMWb0fXSGrSu27w12Frtf/qJiUmuXRctdxmZtfHh+mzda100qs61TAKIyG
yC2olbKGkZPq8qd66fbHRVlr0tb0/c04EGBr5m+ikLD0plMEMRuJBpgt8Wj0UGImDtvMJQpXQaio
ne74WfHMaHCi6omm+QZmUo4oLiwghb4ZWz90epridH8X3+AeYjmebhshcTYi2r58wOitmI6TtlqQ
NGMpT+orGkIL7CCDL/Gfdk6rBJCUt+Tt7TRwYbz9IjdDPmTQu5uCUMcvDF0FEhi74wDIuXmkYeHc
fWpaEjwOvSEf4KP29JfXtYmEvVUpTvbXpjeRryZfSRSG1K21ibFrwRFnM6W40o7ARaFJS+u2b4NN
yD5atVstx13WhQFFCSagdz2EEs1b0JcpSioqhwobsUOr2bdj7DRdWk1TmwhogyfVrTfDPMSLiGYz
zDPPBx7H2OhZRky9rojGGCMtXQWGpzMPTnuKjtbiJWZ4L94NvPre4ny28RzVYbOFgpCQ4leszPlM
J1RcUgqO3MhTBI9HSAkgWB+mQIi7yfyFQk5lGXZyfFwgGizUE28RS4xj7SeKIeV45eeD7OARynPz
Z9mnNCBCFQRnyVVqfXHIX3hHSIILcplSehGXWbg3QjbHBrPjzQWVyPStRBorrplILbm/vojw5KR8
P0wVVYwQvS4JSHXAF2XJ/+N+xJyvmj6UKoVXsgMgTO7aepGnuO/1MI5sI6o/XWoBYFRJ64fVgqzt
KGhhqd71n3O5cmO50hGJ180x/fU4DUXiUMNCxdatP43yqA3Zn72SfqDxpx/T5KE8dxQxhSAbax2P
+layM+U+j5hpsWgt8cnRtAmzDlEPIN8xEr4klsxMOPaYIQ03QUrbucDcszQudwd/Xbt3ezbjxt8u
l8Hm+HcnjhnuoHX7hToNTENbLt22J63Sm3OUiu8MBgamaAYpjCkS3K3WZmblaM7cpB02dom4IL7m
spjudZRjBEZnyCHQdHhn/drAibXMTy9O+qF664IReb4RAb+IQKBVHTBxj44rX8uO5uGzHSqei0he
Pa0ogJrHE4OHE4SobxMmtz6YoZNWgcH/s8iCWURwAoygK4UzJKu8Y8nFB84nlbTkkJcnaHcKckd6
KomXbMiKt7NqLRT1FiKtFFArDb30hdyt37ctyxoJt+V4yLjjMR/Vpd44zwEAVQtMU4vGyubam55M
OEYGl/VJoJVvVcC5eCyvthH4FD1Et2bOOiYHM7pRE1es8PY8IAsjXgk5UIlTRAq1+zjUJp7AY9jH
JTB52xEL32ZUgI8LBTgpgCwY6ZprUDnTnWe2tF5PdJzMmOXOZH28pjKK/3dagaqw7DHGA/vgrurd
mW05r0/nvxInDWQ7l4mxbdStqnQCsM/1eECLbCnn1AdDfD5ep3OepMXVGaIQwzhBpKTlAItCvaZA
oegnkkOB3OQp6n3ko/m8aqdjbToSxMZQ3wJi0Mru0+XyYj0dkh8yz12xfOuPc74vihGp+BDLOpIu
4FqwvcQHpZqxnfTTIlDr0MpbteH2UvBeietE/WgdFl4IGQkHgKX6KsIrxJqRBczYJDohz6EiNbgH
t6Vx+w82hYVRWhCIbDp8MRylAx/GSPQDZSSuS/Gu7eeIqE1X9373PE2r24tX/tLFqIc3WadODu8Z
zjY4ZZ6BDzYu2NYoYs0z1rKbKq7/7CzKm5fIoN7ZcYWzgEl4bq0b+nuoS71MaawhSl+tqr8NZ53C
wTOh74j1U5Pd6gXoT5vxyHYCjUiD6oO1kp5mWy6MhUklEymlm+JfN5d1clwIdLygp584CMfGeyOu
waFozJuFxqyHZAYEyJ1ejUyfAXK0Z4359jCnKcJSXD9KE9yOJpWGJMFbLeGa55JhsoUb2uyX5eSn
Gw6XfW60wSwRhHbn1Gca7hIUJ88U65012/dkofSQe0UK0qbJJCKkLX/H4ji/sWagxJysGVift7zY
MqiNda3+LrZCiLNpqBtVFGu20wPf3SrQOk2gcGjZ9A8CarA1Rm9SLKNw5KjovKpA5an5W8LPSrbI
iHOzNogmTrlqaH0M1rYC39ccbjJ2mWKJxp5srjXrERuHhjeUYxuZZp/Hdoto51nXS9Gm47Gb3ziy
1lWGV7Ct4KXqIEUPqpbf+jkXIC3qmKN671DLyDjk/jQAMi8WSWL4bNkWAKUA2SM3ky1a+wAw5z0W
CRn1msixJPsyiVXR+dvqfpcGOwxJYWimKFQeoeaGVVKdNiniY+eGgyYYIn1rOJq1FZ7AfgTFplTc
13QAaUQ00NOSTBAi6dTZmO7FHYDfnXkUCZqSoUbnv+Y73Xyty0Gh90Ff1/d8OXeBnat0jjmFgC1l
d/23JMakiNUDKQhFX9ISYFOo+MErxZGAnsl6l8DCRL4M/KnrXM58Jhmu+Gv8XXCVQn1x1zSQ9HNL
KKzMvXgV/fNHI1sD5YwgTl8P7baXWbqwzWdMxhnZiJLH7hrV5ClPlkPa3123Xqv0OY/Ll9qfH3lj
5kEbGDzzhK0YMrVwSp8QPopp6x88m4UWCLb3wfOgfaCdNruBlfSM48CQkcRjGTVgBepUFNa76ZGx
eQK+rzBE7df+aYwIN92uRAv2S4unhtTcDw6w3B6eXeGT0H62T7CR8WZTfKUmsjMK0Es9/bHYLSqR
rjJG4chgIO5sXXEgPVGmYb/Qn3/QHBVtRfUwxr01MXJY7693vCA4W5ZZ8BviZMB+oI3vQmqYDX9M
RNLUv3mCGA0PvDLDvH4b+L7oIZxvltjnnz8O6dFefEjqnNNU47ad9b262qBQSC4e249M3vFzll/f
slaNe70jHWL1phH0oeiSqytroOW7IKB40lm+F3DbzLjYUPEZV+ehDX587Sqdt2hMEbUMyPOVxvov
RdydVYehdK2prEgi2EFXFlZFshNjL/lSapuV7GcALd5BTuFkWJtvEFgY6RQDpMS28KUB3wCZrE2T
DDNMgLiKTSNduzljQTb5zc8XSfc68TI/q5kC6B3csmshNc1reE0yMeM7Kz2Y+/Vk+Dyn53djjYg3
sL4Z6my9eBgiEFJKsZxi+q4vxER0Hn4lFT2nsM0uQ5MsbwTC//ikGwCsotDXKaZP/0VpgbPWDeVl
wwjDyHiO8EB9IyCUtfYnYNTcpMIyVRTc2Bnw9/sdMUwBiE8TTSC3DwLX3SRXfBYTab11iEMMWg2q
ZzHilB1GL7f01NEi92lw1FEAYxhEx7ivnkcn+NYOutK+Z2EvAu+hanStHBOvxSjoy+fXew6sRAa+
zSv0g4KQs6eY21ea0OvUX+K4m2hbyz0N1EZ3XT6yyAxLiTQ8HA070K9hFpeUDAGZm38WgtbP+39x
bssn8WceNgcy4z53GpRYDTFIlQcgHQHSjlsNKPBBcrAzGl9mQDHMaNcO76McBMIdu8WxanR5GAVp
MIS3c/jSi9M8q+7pb+bd5TvPlUjHaj3CCJN5ZO51H1JCQmdQpwfUld03rV1Cb2qztvG/baOgfs7p
S3Bc1QdnVRZGWKy5
`protect end_protected
