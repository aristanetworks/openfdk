--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
oIOFQ3kERl8U+fLErG97UqI3YIxvVEdh257dqnhoXam3iRAwpaWh5v4LvkvfF4msCznSwNC8U+c3
AJRlAlJ/NR0uPPJteUt0qNgPdz/SYlUprTppnN+XaRtPq6OOCdP6ngYaumo9xnCtXXgepc1dzaA6
2EdWeSHN/mZSmX1mhDQSbNVRkGrGVDiFw18Ae0g17H/7tadnD/NIMqxS/JvfrOIVkhfC5Zx11Lcl
26bqBTUIFi2JCNdHhVQqOQLTQbetIXYRlcJoYXywtcvV+Otl3Y4BDJ9PdBcVUt4JsGTWYas3D6HF
GlpsvpqN+H3u3Mt2MRNP+Nx37UeAzZx6NgeR7g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="4q8b6LK7PFmMpl/WvmQPTuO65QWmK7BEbR1LhfYPrF4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
UZj+lCP5TvYHnVAY/I4inLgApsynFqnNSglP2bnV/IEb0WXBXSCIYjqqUMoq0DfJiRDe2sXZF9Sb
1dNUXajSJMvVkUAmbBARUa50XgtE99B13SCT4cVdpmUBBrynu/GK329pXea7MCA1R1hcONB8heKl
ssa2en5/DCvHdJXke6oEEDrALPxLyu9zZcA+uWdJZflkga4zUga59cLUR9vXxjhsxeIijUOlbQG2
F7HcwrUvGKiW2/CycMsZB+iOXi/2+AhQeoUZTbqnhezIn2dCDi/muf4IxVjZyhPcO2OMufI7l2Mg
cknPpNDvAKeXgfZS8I8swEJJy3NpzLlYXlllbQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="2VeMFFbRNOIzVMO6EIQwqTXabK1PvRSgNg1fdsdRVeA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6624)
`protect data_block
xyJ4hS+iK03DrhCGqh+C0X8sdwFuUhc04BN/uD5Ys5LJXIqs0+lcLwvjyB7Yx+irmYTlJEXrebMS
BY9xfBGae0gHIvIgBl/9+L/7+3KeqEGVNvcEG9DfZKvybK63PcnUv3XDSLclZ6Oqlznb+oDwSpvA
6xTNTzZE+SdnxFvgBvckDKJaNz2pNhsC3c/Q2r2r+lckAnzyciDs4kufr8R0bpRDM2RFh2/dcECB
R75gQCT6TyRzp/licVa6zriObh6tTpO0LWga0A8paTz86PZODDKwEYqrQ31tZ9YZG8shba2YGAjX
NxZd1StxuO/i51K2pgeKO7MlG95wTBJNZj++a9YQPtgwY4NquBnDuuthW1uXrVxJvSUea8bCv6UQ
iefnMShtJUPyMwQhxNS2JX1QcKSJg+VdfuI7HXhar5DpXgM9oPWatjkL8JknEpCLcBWj6CxUv5fE
vGrEveBaSMWQMGekgsxenJRO7yyZWSCJgOZ+N//Umk39J1wFDm0VKl/bO5Ey50h0F+owtpUv85bK
nxTsa088p7ju0OJGLrA3QkaDUNL/KJjB6NG+2cXX+m0riGfEJtWXPV2P5xQMsoIVh4H0t0cmxjUb
/NOyA3rt13y47doaiQp+MnGRIhEBHMQ6UYbTKI6RrUR9SoqpQtnNWSEJtnRQV4UGIUBbZQvuKEHK
EZ8EPAVmvEx6zZpesv4CiAOWPTif5C29TwXmzea81rInol1eNjkFuLZIwzr9iHdisxjNiT3P5Mee
dAs1u3Vde6oYKjIcwWY3CKbz3OscM9KbvMlumXFu+/Hnh3OQXO57RJrbUWXhGolw2zadrwftcPuV
o6ah4VD95ub+BJcpPJ4oImEcsRrKPIPxTtKtZr+HURIDsFzmbH1+QK/JrBsydHsk3RyfiUWMsWxZ
VzxtZ4/3ZybMv+gyuq10QJW9uVMz6lgNL1wKmUK3GgDEfKYEn2qTMgP9LtrurdIbs7YzNn9RtQLF
3rNZlInNWS7C4NAQcfZdkv2Nl21WHgPQBwkusS6p1IFD60D8pNvP7wnQbQAZmlBmuOAO47vd7nhZ
Mj/fLKyuUYGHEw+s5JOyBkjZh31MX6Qf0Uv1WePTsTOn/GL8f9hsQNl4JD13KFNu9XomR3QQDfNA
ABUfhXve/S0KpHyEUPtlZyarcs3KAMuPiz6Lsjp5ggZzi2Bf9HA0PS1Gv+QRhmDaS7VyQeIfYjKv
5h7rpUA3kvRzeKx0MGBL2Yx0PJaj37wbdvqrNYiWDyKxfFfS+RSbS1LISz+aW5QWU4rGRn0ikoEU
8RFbqbHegeLCr22LodmL5xxv+yi+AgGJY0htKQvi9tn8CXQrn0m2Wqw+nTCtzM37FciRvhotX78d
KbIx9vNSDhb37R7nmQs/fscrRutbPLXy7uIJMbPK2KmSwhIjSPRy6qFG4wY4NnDUdeCXVVnqFtee
58CBwu0kSi0Me2AYowH788xOhh4+tBNG/tWSJ0ovg3wo0pAe4A6R9GFQXBFJ5uHetoSZeTibBGLy
KfSF2T4Th/OFLaj6qb1GFQTqVkz4SkytEmY4yaxEE6MSL8QLl07logVqzQhxuyilXsa2NTd1N+jc
XKvrFu9umrHKw+Fo3KjCcbFcTxlbp9qz+Yd1aaAXVANpn+loJPdPzxfWHo617YURXMwtJgWHshQk
XSRVCUPGfilt1nUgSbmC+a7C6tAR4nB5GZFRZchPfA92g5ll4C84dtUpj7mEKF9jKG86ww1i7g0A
tnP0vTflEOlfqAms28JODCOu2AT81LuBvs+zrL63lXVYXHeLzRA0IX6cvLmzdN91V8xxi7lrShWF
LQxDvFBgElJW7xK4YzAALMG0OuMr7PCAprOG7QOr4owSQt8B5T7frhN0QD4bAcmw0pMsBoDpzX1r
fCjuvQC4rHYh2ADTee0IpZLtI5DoEjVzfmICPZKG1FgYzRhzzWa3s5gA2Q3gyLqyDrLYggWEvV/R
avRITMgaK+2QvGdtylsxaq26ZnchukarFeBMqiceIcNZ8JzT371SEWPiGDWVbOT/AQQK1q1Ybc5A
KrzG9XyhH+d+3tGQEa7Df6zQuNMFy1RBrfvkTc+TtHZW9yx4XhVGmdKxidLylJa42jE3k5ck/08a
FEji87YisJc8wtAPclLAFyTMYYJo+9tPt4dsnnpcptnL2Hjl7rwf58K6APSlLF80MLhb4shi34AC
LeUmmld+3GVAUZKYSv6NlIYedaOk8rdlRVMlQSTeJlhk1WCMwlqY6YbNzCZ6rubrKdO0AaWj78TQ
8EAW4kGUoO67Mg4rgF4znOFsqOBBs22Q8FUIZ9bLLQWlcDGgb/mmzqCafCAwCaDihmf8iywM1A+2
FBj8nSjcfG/XworyFwxfIxRLphXj3cFNYmeObNmXO8Kd9fcXYN790tXJ6OAloH2mSVkhyclqP93+
cRFz1gSsPDgktLRNImGpsG8JIaZOK6DPaXTDRlVyVAZjnbASThbg6mZVVDJA3fsrc0W+Tle9psY9
7sPCu7+VTu+ycP3ga/t8wr2X7WKQ7qFUpx+SZ2XGlytJoRx6ETG5DoU+pOwAKgn3ppAmAyIk2+t+
cpwr1TSFAz1LQ9ohq9TpxKzApTX7DwBOL7zG5PxPNuXTCB36BuS85V2BA3iNoyYqeDnrabQZTLIH
iQuOmjdvUk3fwSQn/2EXpG1YrcSlcpjWmVuv+9SF20sr5dma9Wi72r//50bflKYUCDI0SSD9IhWm
XTXRvpy32leCrl8Z5uSLiee4XBUOSpFvbFI9sitYpqm/TCCGDyXJHbS4p8Xg8yOq4beBAjfgId7b
+0BRH5MY2dKOxp02j2KSPoAboG75RxifMPvhDbwpilxGyFDBNcHe4c8MUb1jjb/ADehsYc1k+IXG
POtfGMDLgKpcQJ3/Q+3lXdjFvmnTvQd7UqnBmtVHNkL6Jj0nNvgmmLcyY75C2EsIwR8u3Fs7eE1l
N1mBGfOVQuUaec2kpKBYWx/wXXSY7wmpg1AiYO4spfWskBbFQwz8fTj3S9gLLxxDgAmyGVezMQtc
QA9d27g8Yyi4O6N0XfvR2EjCu8p+we1nTLALvlKDJpwuoIVoYKnkcxjKgICRFosiC2C373QxIriT
6KcZtBxzLkzbCNsfgo7C3eEnKIqpzeWZWquq3p1QC0OXym4vXLL3CzL01hiJngfx0KNXwNm0W+Eg
De27+vrElTuivezWAiOpuwd9kP5CmzO2gFPsy4e+IbhXS51FuKV0u50XT2Kav62PpcY8WulhCgjI
bOjk6rAyeNVynW76wDEutpvvfEwamtnfzpoCkI/2U2D5wJPRlVRg6ckh8MpeRNkj1ip9ZFrvm8J/
+o9cQIsVGORj4U2kxag4eIzQV5npjvRjEIp1TzwDsrYA4hko4dK2VXjQtQJahwudIYA3nZ7w0tMU
BDiw7UgBEG3+q5YYae43AFWIR1fXkWBW43q0vVEL8+dd89RjgB2ZUie7GZSESgVXvEGV0JnhpVsV
18z1M14lAfQzE03wEgLgLiGkFFTK4Guop23mWzRRoOY32UU9KOe9BNfcAfsfiR0RmHYSYFJt/LQG
wQNi645ayItedyh2NbwJ4uUoRD71LD6WeP1U1JEAIbvhHMUwslzVvkcRajLFpyUVkeIj8/T90nc/
GAGFB8Rfyk1+E5Oj71V8qmgAZG7Yia7gA2VdOiIozsOwfsHKMhxVIykqT0C5s0x9o4mEJlh94Pmw
F6AuDEEL03eq81OZEAfSgixbQd8xn2k84vfpTs4Vznz0xls+/oWQiSIrmn5EypCCdTBb8VNk5o76
5v7TU1zQDizD2W/O14TJ1gbPnKPqwDJqd8zRMqUv3UTAJihYYA7WLqZlzhCwQzd/gFghi2RSvI2p
y5nnUZ/vEJnfAldSpQ4xXD2VMYNei8hgUPRgOS6T1QVFLMkdFtuS+qKbaQ5nmEEs0XjPhVt0y6rL
Bz56/P6Q25cJCs79bisuHamrCVBD4UuqaNpd4XQC5p/xQ7mRDtViLelNBuJg2Z19r9al1igvTmIP
TVY1WK8Wmf9fWQkEsUYKxLdoet4ykXq7E5C9mOKgmG5aGnmXDT55Qut/tbWq3WyGpwZZgOnDry4R
OyqxEGDbPrM35scATa1bBjLPn6JFe/eUdgjsMkavl/cdRtUghfxRJrgttmPSXBb5x9V/71M04+bC
zjsHQLre8BWUT7apKLjg4CyAUturpK1rIOgeWwOBumyVN9afncOqxNRe7lfY1RrRhwOnLnTEyMux
NhRsENtNHaGo7GZn9WQnHolfEKb2MDR3D4+xGlKrnoYnWYSidoZbfm4GJCay6WPhqL7sRPM8OqHR
b+gwHRNrWHQPHN411zpmFC8JjFepbd31IQK0MkEmM3fIlt1lUPYcN+6NcIgM0Lb1VbLw9bmbV4+r
Wq281ICacLz2zjYT3IBiGE4nH2LlINj+x4lSXABqISVZynqihL7yaRnKl7roxlURIDn6XoMTUmpR
MHIjk8KcSplTtcNl+DWN+/8d/J8u/J6B9Iefg+xNS8h7izQBoF7GH++Bc/FZ1qfMj33rqilZp51b
G7oJgQNM7f8AUMKCq+R+/QzqX4jXWTsMu7bcoU6wEi5jb1B2WLl3eWo7QMkDS3O1Bba53/oVbhYO
ULi6IlwdyREki/IS8/UBi9KhRRT009QwJ4cWwkdY0mcqLYsVMU+dMQAlH9NzYkwqvEhftaVGek0p
MUd26cAFx2XaFCzwqW+8G8uj7oC0EtMLx8UOFGAldF5R/gCeh+0vDhjexaZxQxVXXbtyvV4lDyic
fagvTbsBi+xYP2qCYlDn4HO4RISt8zRJdhedylEgWA2idaeetFjP1l7mp5N2noxhhTwgyr7ZSI7L
dapaDoK8fFECheY4ica3PwDh6I4xqdz0Uq5CFpB0f/hPDBOvuetlZKxAmb/IScGFa8PiI+OcUgII
4aHDqpRs1nZtev9N1ZMlMWM2vn2YOpSYER1bUkO07eXQthsR8mjfUL+9FzKowxAgNgM2C4jpsjnC
UJIvucK9J7CDfO6gsS2UPU3s9dgXsw40nahI1QFsIrkg202oArf2zckAJ8xVqxhdVYn0Jj5+Q+Zc
AnZTHAwO9X5wRmhO2nsXZekkFJnEwVLKn0xTBBDLmxbYMQPWGaV+b3SobDwPr2OxvqFhNRdOiPj9
gsdZOZIWI16pfmaQOQ5VJpiVHn4lny4MHTryp46IjIK4mf6/zZsfjrJ5R4XM85pvK/+bWrgdDXnq
3JgT0l3jlMS8e/ljvZQBzWINwcVunbMaGTNTkNmdV/vXRmkeeAYDkdO3yLkfNnL8X+qnabWOI9sW
qZhObNG/MwQ3xZWJlx7uF38RdR1l+94OvAZNEwBSNYHpjIiaCr74/wMrs0bkfOMlGurMzxvPcw4O
mqMww37X0vzMgCWODXoMSYSAKfRIyg8wlF3aaECutfRYn4UGpMh+wKk18xf3BChWUvlaa8jJsTPX
sH4lgWaC1Lt6TJ/XXDhgRDMvzqaTFTrz2/ywXJCLcHIYyXLHI5ocNXAtCV3LzKk/gleDPpucYy/a
757D7jnkrTys14wpqrsjQXA5moqVOPNIrC1/TJzwVOfsxYQBDXt0kbeoJp5STNm/C3KFf9C+fosT
9GYdxUBGgOnsgU94mp2jFjcMstflGEBI2wAvtp4TZKrTDz2DRTP5aWqvVh0J15N8bR0pwORcgtDY
5ixODCeYIuRG/MC45JJQwF3IBVkzy8iib4bW76g4nBXJdkvqq0eB2qC/5pOpQqSS0thm2QvmInXT
RoNlWdK+9L4L5+IkIUI5wtpogjX3RPAkc23yaIwyZP8CWRR3+D/ltOIpvIArw7+c6ZAom6zm1OAJ
Ov4KsEhamxqHrYtx+3drclk7DgRH7w99+G/CnNoXdMOnurl+5wGTcoh3s01e99F/1GXz4vZfqYfz
qpqraH96ibBI0mRkCmh7FBAhQZpVxdlAuHuYCp/Fp23sSIWkUh72SG/cQ5LDSt4PpIjfCmZiu1KR
PHMf1TxKjrxmLTQrF3pbF8qU0dqMsUtolXu9RztCmco7KaCF4JTu55gAOpRtPf1DOuKfc8btVQEn
DM2WKf7fAuWDPDSpABsU0Ti+406XaFbi0d594r/GC9gYcKtI478ndFDTvafgG3Rt3LQVRW117fkN
DTfm9KizeX6NAS/9XWZl+6Wz5ncBP2RrhGUCLuP6kItUl+yd58e+DVJV7XeV+tppQMWr7apThYV2
q5+EZvVQ1lSqfqdcK4KUdsCzJPET/NV45gKun+AkAbymmk6R1KvKi7aqU96HoZvP8WAKdd5bl8HC
99IJKW0lg/CFODyFDHOhcgIgdPi2Gv5pbTJPdogEzej1eulwSDxveG+zr4L5jJHDDMkeC3/i3/RO
uwerFT1k/qF7KgCuQiBzhTQEnHfWCkapnJ0hY9psdDy9csFWskrONPFCsUuYWVqtwz++dKHURSb5
zJP8KgNfTpA9OfsS7Gqk8V6tVS2NerEOVBNHBqUfjerypkYWmYaH57Ptin54LQYcAyVIAhxtsdng
YvaqXYJzazkCnRW1TsjI8gdrDw9uNuIB45JjwnzfB6bFoXfQv8pnoHAqxZGCFiGTNyHDO1JAyHVE
J70YpsXuadXpQaKWx3xNqCpdtlmW8yVqjT0I5MFDK7Yj8vmW0KBuu5tYeR7TxhVnUnvkSLz8dj3U
LDmIWW8a3Qib/qr8CVsMgGukQB1isVc2ZDWUPJIkR4X+pTR2eq9TiW1ZRWqNdArL1oxe0FWMtmIE
v0OWzHMB4F8uSeJ83ZMPo9tsqYp21eiWvUJU7+uDn+7YI6XNFf5qceD+uAJMgLnqczeThNLiEZi5
PFtFkriqYNfzsgZDWpThCUKwqpZnkCTSXNL9eDqCR8D4XtBggUsTCwDDhw0SZqBAA0QCN+1GRPUn
pi26LS5ee0YfvixnBn0lWhsGKP/tzuXBt6TzKbELK5vNiqAiCa6jABELxV07QO+FBNxRwNJ4Q3VN
Kvuu7bHKL1Va8luSj6++sG4JrUCoElBIt9+4+o26OQ4ncLzBp0YXfcIaRKZkSkh83LkNkX60OJoH
3mjGKI5jVAdkc7FWNQpT+kWvrpYWYBPYW3x397vYr5Wz8vlPeTrIMC1KFbgE+zNHomUCcMD/Ptk8
Maiyqmj1/6oQMRCanlJbWLOD3W9dA/2LZqW6HGPBj5KxOonl0C2J1BbPkfYij6JJ5aCzi0vK1sjp
KUsDnQI9BqUXBswNSJ22Ws9CpDY4y3cpbwOrvWHR0YzwXTpve5EfbNJW7Dauk9GZpCf4ALtRAyNh
Upa23hHDBontZiFd39qSpKbbzyg78t4O5wDFTHBJuFVrRLEvjS8vraAOUx78ISKbqTw1Ja0Ta13p
ReeIbxGCDIlWQhAWpWcsE7SdhA3BGxJtdLkVBIkFLaWKjKx9xmjbhwjPUd15bZUzMCbTsmEVGVku
R7SL1nLND1vwnGwqZEA3nPXrCL+REquPrJB7rhbrKij/4bDUJ96Z3EKFoaOwU7UCg/FEKSid4GlC
2FKziq8VD4k6PXeU0RBn7VqwvsM3+Wiu8DBnTZBWmZvX4ky5r/v0QTqSgrS9jY5PjsXwy7Sp44Kv
5vFEaAx1M563HpbCkUl20ZycH9bKID9lDF/mNLzp9qvJC7RBoopNZdeflkXs1438vt9SsI7hiyDn
UKdU3i3BVRhxdsRM2Ck1zUHtfz5m9qkGygRQSTJBC33ebhG4rjD/1RpHmmqsIyiHQM0PxJGQFj/O
ie+/z2mpO/AHmRVI/U7g4fkn0vRaT4tRWw0nbebA6zZy/klsKKMq/x3iqC4Fv5UGPEFg3oCnKZu1
m298LQ/tWvwTiUix0MfNjnBbK6huqcRr8MSKSccXWnMf0OVfvIdqoQz7iWpAbS3iD4Jx/x2t4CbO
Y04lAJM//EPpxqGaJNbt7KdiH1TUIlwRR1GeqGRu0Ln+QotEpi+lDMj5xgCiUPchXxA3Aim59L3H
hNx0KmzaHGBzaHJE5jew92ML0VlvP4/Up0/dZ2aFra056/uULBWt8UUmZGMP53lzfWguYI+BLXuL
lnhgEE7h2KROTadYbQzNBuae4VjfNXBBv0YvAu/ZEdGu4ICQg6vZHbwTquN4GYgNFhZR9jbHmINl
H13mRV7vQw56zXg5Mq+/IZj0Ueh5g1hTn6SO2HktK2JBVb+nneDJ3uLCwinz+S55IVXhmucIRyn/
XdD75IYY0cLIfY9Yx4bmDcM8s6+kqwNP5R46IC6LdeFUa2+nDTYDy5JVE5N4E4V+0y+onyge/Wm+
5q+cdLTC3+OfXeafQ5ZcIrUKyBlziXPpbH2y6aV75qkoF2JeGgU9KT6u/lIz2y93Ex5UuTmQn9zu
mQOOU8ucV2bjLObwA9FEpwMDg8MgvhppnAukHVfLblEE+88QzbD6GIm+b60fRizPoiu1X8Xe+qkb
cefsa+0WPmIN9wySL2n3sSzWWq/Iyp007AtB6mcWmHLo3ygUtQ7MWBIHTCZKdBI3BmJMs/0KVh9y
HPAvyJspJlYI/FokKMIzIK9rNBs0tq/2TbWsPlPvGVwvKb5n20hIfoS/24fdcp5ppGYPiYE9bQ65
aW18Yi8GInay0eIwTXZr7eZ1r9QZq93gUHfDwCA/qUPvZ1D2K5UQC9BBwHDDzqgqmfeu50zd+IOv
Fczl4VcEj7+ZB3XoGDcA8BryVSPUpCsVIJiwDVIchjGeh8LjWNfAM+ND2XFTajQsjaydBcbKLp2h
3RHJSlje8bCpGPctusFJSMYSUlAQZ3V/Dlc0gB+Sg1sOaotkldoOEUKMREuS+CjgM7D1xFIbzs1u
4TXRe5yYlZTX0zxs
`protect end_protected
