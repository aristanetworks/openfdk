--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
OcODJUzEt0MDXk5EnPw98x4AqF+VNbUNRtbbN45bzY+0JuNLOWmF2ZxIe0Fu0bhyCaZ9JMeQD4Lc
i/1R94UJJHdZuBEsy6NP/fmQ8obQwYM30fq3NkK3g5naOuHhKNlDqNPYJOFFNw0E63cAZLDIvPOI
+5Ls47OBhtufF/JRONQp/1n2odTCY5wnNE38EzqhfCiq86q+k17yVPX66yQESwt+v2tnde+3nJ8E
g/8aSOCf92W0OGzVvJMqCIpzwh9MdWgGJNbndzwXgHBcaHHA4GWxuAiA8aDxARe6cF+1ftM3sMY8
glOltyFghqVL5aUV4rgrhX84dagz3vBfUHUyTA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="+cnnD5gOatx67wl04vxuLQxgS2r/b0PcB7Q+W4BCuvg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
SXfiFTS3dLqv+7R586/KVYntVLDPbyCR8AL0T0XkPvvyYENr0uQVl5mTLOdcXCHPzav+sGGdD8qj
ldB/lh6gP3Mt06nlw+t+wEHQvARFPVbPbxcgAE1SVj38LuEKKXjH9wP6/sA/JiXYdsj/hTXJf8Us
S9wqMU1CNYZHwGQg7omp8CGcqnFdXEZ8tKrb9Uf9YpxREQ7yEY/og0mwFLVydftBZC/vnK5O0ru4
TSlrRAcx+P7jLL1kan8ShSaamtt5s7GIfqDRhzX3AFUxa0eD5pk4+e9YqbCf2DKj/0SkfUae7u7q
lRiVOynLGlPuLDbZwIOg+iuWat8lwV6+GHrVEw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="tYSoFR3KlbD8A9T6fwRNVKSaRvt3pFQlZb4N8nidclM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7632)
`protect data_block
/IZgobB4jA3N600Xv7sJ2Jj5uTSooNRSmTBgov9sPuJ9JUWHIMnjh/+GNS1d1f2O2j7GcgAgrNDA
R4Q4ypifK0CvpHIVBpfZyy/AXY4JStI/e1omcyvZ1eVL6h3s9PZy83czRnjfpB5UDg2CBLPYvW+Q
y9l0rGzI3Tce2oBZUibPZlckDIPQtzVaK817H1ogKGk/pHbN7A7hKJ4Kr8kggGvK5yj94GOkKTQt
1lxsJD3VtXut+gJmObNJV1cewy7TgWqmH1960Kbwx914UNDfy1sNWyNrif+iHYBfTIvR3LbaCEat
pdEq5wVNg3VzHd9wJ6pH2phPp4EQP1FU+RTn9Z7bCVZUOFsPz5vsl8+cZtj1YvVZfZXd4+gsS1bo
P5gpAJ1cJ35bfIq6I+F5J5TLYG/sPJ0stCwsD8FuKv2+o+MAtsmSgoVzBZxkFiWkUTry4R5mauxk
XZmtoUwoac8eNkCIZCtfEo+6+VgXtdlxJ3lJuhL2INiUAujURiR1OvEnxVK1o+jGwMXP1u0FM6Gw
lcAiX6vJiZfO14E0iqtvsXrXIFnsHfIat5lQtotvw5AScQpmTpXj07BZCUfRvki4uDPJ9eJdhK50
JyXlEsvWHVntF1P0lUAUmyjYeEfkderygXvDPkLNfp6lN3XTS+B0kFgWU9MMFkrvlpsp7Vkj1+Xo
RXoqyZFTwE1+JXdJmyuxG7BXZIFAZYXsXaviafWAqk46EuP/Z7V31mlO57FdrnSG9pDyCEhcoFo5
fiAsKci5+FG3x/CmH9Qcvjfq32bN90JIWRwhcGqeTqXC5VUrgWrxT0wQMQ6Sk28JSpcxEb/4EfEa
tw04AedtDeEpyIggqhqFr2AE0U1wRH8q2jrhOXx5kOB2yTRnrPEbcdlalI2tGartwPXbE+LWu3tl
bmu2UbfbxQtSrOwEUAdsRQWZQfoQ8U1Vo0R7faqqmQfSe36sWfDTtKz2byuQIG5fX1fJa77naUdX
iupYaR8o4D0/o5dWFqLbcsUuEQwdsRQp2Dj7IrMKI2zNHDxMmPaylifUQ3v33Pw2KGX851hHYpMi
qIrM1T/EM8NyDmuaAS8PumplNLk8OAskCX3TT1vWgW047BECIbPgjKhLBlucOr2ziG34BTWiofSI
aDz+NMAIAThFhahCS3nEIoVb2cjI7FAbTSGx0rM4v2PN1Dr007FGEi57MJ2Bn8p7aVfRGbVjjZjD
dtopiQl7O7zUA90E+WwjYq/5ucXXxssIoxlbDmieWrmpSHQSfiDF6cByclOySjPQUk0hSeUzGh0w
8uWJMizO86K+NqShwcsLMbjm4UoVufVfIX0ojxKO+/mLprElJ82S0vsxClLA8JFZMOKdasgvxfEf
gfyr36VcIj5M5zBX/3k9DVLvtqq3DlKLsTrl7NE6efcREW7f4V65gB7e3B4MoEadlmQRUvguTpSG
JLflvKbjCpL3jBBWv1+z+i3HK9t+/hsa1w5IJ/B76egLkcZcZtLjw2wOf/g1KQ0ouPEbKNnOV3J4
bjA3+7T9YMy741hLkZP+yEVUEmctlSw/dMCrP1e8POOA6S+qV1CG9CrzsJchr4kjszyu7PsEdMJ2
doUegnAK/xRg2sATnbjjhGpjedJ/ZEsRRlO0BORWWxHGr+BNUFbwPa87oaru/su+l6FJqZOiS3p1
bNA3XeLwfpSMpO2EK3gphtMPnTICSKoHzOc2r+9/pjx+tRB9VaaUI+9h1cto9477zVjUTRe0eMUB
dmUhV6jZYkvWChgsuvzpNVTgSqhdMsPgVnsZpLzp73csBNPmza59jIM6b0u3yDyxiSM9mBdWJT/q
JyFnk3KNtxFpLHt27Q6/4QGAS4TeTAmpSdSv/piOhwQQ9rExeVTwjaIgnODnvpbohoFJcWHqUths
r1dL7amjM+WKFxuROm4tdcOgjUOm9ZkmTb9ksyxtOc6fPNP6I5Q3zT+RdNkloqUQGW9a6UlRq1s6
Q7mypR62S0XCArltatFvWvz1ZB4bIS1peumU5qFVQ0+Z37i+gDh32R5df7vl5gnN8Q7V9U3J4mhs
4YYB3BKYIrl7F3JxlYRSVufqdbmbAI1NOi0AvCs6NjR4H4k/CIwmcMG0RqwjZuggwnweSfHEOvig
bsd0YO+0GMLVJoio6vvzTqch7Ls/YS+jNOZCQqSRPe6fX0QyeMCn4ozz0a8rEWdcAgzKJqDYp8IU
OEir1hG4urmWV4P5CmS93brr0aMhWpXKrcqvCmBFILJ7wQ5dXvEids+xrOiPrwheWFnWnvBzwh2S
T7GGpJaN7fkQ9jtFAZRTBjeapRBI3wl6IP0A8noZcolyobVtdiNVT/GQkoycQ1bzcnMxRILgtGeN
GMUlHslzoFW24YoP+n+8T9jFjJxTTG4tiYuyCsxpr2PdhLCj2oF1Yn58Cg2rNAl05tXOTeLd+QZk
HDepgxEXAd9/ncxi6MYV1HHkCIRY3IqEvVAWcudfh5nmCUKbWuHBYsv/rgnaFEZUX2e79c7+LO+i
jF6zUrMXMmHisdw079ltG1842ejhmI90myxwtcteW/Hi4Koot7STzKHbeSLe+nk4Ed2Nn+7MV5P4
loV6OVV4UVYAsK5ILEypGYy8oo/V5g4zpjdiNkzdYjXDePWDA0ywHchYawjlDhvBy+zqg9FZKm2k
jz3rKI0+JYS7aEYfCilY3o15RA0eVBKb2PDIrgQs6NTzwGtS/Z2VVWlpDHY6ugJWSj9oNIcvhR7z
xkOhd/pJJEyMpitNEtPlTyTh69msctX+2/9e1MyOxbLRgg7u2/bDrZacJwVfM+xYtFBB26Qxfv88
hzy+uBZHAgcrf3+wNgnW7emxnEgTo/N6rZm479d+AuG6HHr9s9Aamske0hY2TwtVRjCG5crssyW4
Zki+WY2NOoGqWSx66nwCwNywoA3KcyaTG8KHE0UYQB/9rkm4pfznj+/xHYbfCBDQ7RX9D4+tw+j3
2cCCbm35/v+5tJ6FdBJUae89HyVDMNwr01hQB2nczHc8SMPkulHRU3rqhmh23sFoAYyahoB+WnWy
fFctOzZpI60jYfj/+dgg6rSB0YGwb9xvHQWAwPZfXZezX0eJ0m8RYKlvFNH2f8esw3KkcCwanY2R
b2vH3qSqZqy05jzV99vS7k09MoasFBJpP2UwJHdd2R2K+j4goBDV+bzrAuwyChZFB9FKHIdIfnY9
VdlTCJfTDeap2xxyLuYbmJzeRqcqAWcCNMnzwROSLn/RB6WzjWD6Gu1/1LnZc/mncOym1FdGaEy4
hmKPE911HlZHR957HlFMEJ/B6BwB9sCX7mSfFDCpxGsSIRJZOtMICzmUGsZi711MuTJxvRG03D/b
jDqh0N/eDNJliNDSQSzL8zTujcdgS0wYaDZvlkSAxqDvu2uqn7as3gjIDCtS24+G/iYDdapaczRT
pLfr3eLNZ0gNyCphG2bof7AMbhYpIW4P1hhbTwwweLv/xq+as5eOwhlJDE8D1vkJo921E/pZbylN
DUfuyIOt6xt0kCyDUYVGMoJwAVliw+PsRjOeDB8XyLmDy+YuxiGDzIM6ibFnwUsGJvHHfB/1+aJm
IYuWEoWR0eRSuL12COpHBKNNxD102JRMyMdY7N8sQ/IMKbce0i9LArpbbybGWlC5x4degwS37Qp0
wK2z/arHRdqyHecbdZukyYgveAsusdL7nXjUUEn5iYLuZRoFoeVASwRp/F7erg5qRO4Sw2P9s9/j
F+sfQ3Hl4zH+ykBbkJfa5To6S8cM9xrFwpyWAMM9FDXSjAj1HdiX9WDLnFaa6AFXcHcr+BpTJZNo
FDbPPK1ohuBIF6atYWV5o683OaqNdKb93ZfJgwL95SG5F47tXIKIFiS4+kUDg9GpIzyZFUfqVwTk
Aozfs9XTnC99Walfrukihk6Jmk8VbQqAZa+3bNtJnp2bjvW0JHrmekdCExIciaFy1NMpG8moBwS6
t0bCqN9SSvfJCfv4p1ij0mGdnFtpaxrQk3zh3dCPvExx+3VUPYi78UnZtOfr1QfHEq62+RX1m6GO
vVeqcw/4N5L7HA8JpZyH1NtzVmMDzr6uoTnW5KQKKKuGxqXOkOl6dg99wu/uNIv45GhMS/nwpLkU
xnHya03boGeQqygQ/yEol2r6bmr/25jb29PCohKwNJzZZUVMcYre33Je3bqFPRQTg3iwEEfuEfJF
OV11cOxwb/VqAC5OQ7z67jorZ6mkZSMvhGsRdx6/CrkT5q3bHwTZFSn3mNTLbWPtc+cNhoTGqXkL
jpbL1JkjQAMfiu8/Ftpe1tZJ/bZxz+gEQgZWBnzK1eWZV+cxIysmMXaQL63gKM+g9EN2qwBSuSKW
ae1Mz7qnYEkPU+E0bQTKXaLDWwr8UcjXk7b83DIVviH1sQ/11Mc7BWboVtVyv07R8BTMk+0IU3sY
v85YlCgUZ3dv6yZ4wnaQyYMrS9PXU3CPioceVF6SZisrXgZWVkYW6GNB0LSOHcdPRdSZ5y6bqpXD
OGcYCrnVNppmOtdRgqY8lBbXXcax2//hSLpMWFrbqJ5CMAOSpmblb5YQy8ncY6SvE5zIUVhAvFcV
l7Mn6Sy70EwlCzVjqFV9KUAxGXLGsMp5RI+P5xBalvqs6Yzr6lyuBJxtBvOu/bDF9pwuyOXzDpWJ
Eg3demcFoXqo+AY+nVVPN/5imX9n+Qx+iqUD9kdB2ocGLFn9nJ6gBuxjJIsMnVGox53y/Dyq2fvU
uoQ7HjbbRcfGDLp3a3/cmxMqC8RMGZd5vWaugD/z9XUeowUA+jfhO7Yrzqym9J+gH870PzK/UZyF
hIW1BlFEf/21KCPKaeGF976cOJ4EqnzCpWTrD1KKXKgYLbWcJcYpByMVtHp//ZP6lVgnllWDHo94
ptcjLPgeWbj4ZtnQ3JehbbVho3jKxfURYRhXpEmti4fS1YiB1bvT8qYx6ZwQoP8oTObzDA9rmsoe
9sLiiOUMQ/wP3j1Uf/5bXiG0oeA395oessb5C3jVB4hANCCGYYm/QAv+q13yQko4vcReQiWvS1uC
Vyunh+htznNLGucBKYWAvIU5X6OWDLWpc3uSFEZHv7vSDhZq7boEJWAM6ZySIWfcUwtnjbDvirlV
wS+2pSHFHYac61QLpdJVtspPdPMsP3jzS15ItW0m74XntrmftpH9liAYysggQrzhg4OXA9c+A1r9
jXuZvcq6ftAydlNNcPqBZaTognUylBSZryZDXU9WdMpgUDv1bMDrNO57VQKx1GHiDTuuRGzQzK/1
s/t3yeegKOgfLm6dIwb3nn+8XaHSxAox34OI/D+rAibL9U1TeaDKpqNcScuaVVFClgEz8yIHvaPX
VKseRFSRoKgUNWtzNGint1KqYeImwToF9CQXmP6Je9C1vZKe2sc7cphdgPkOdgNbJMg5EDuFN4aN
y2I4ln9BNnifPjngVCsodxah1oVehXoSd/akmQ/iGy59+r5rtnx/uiOLwldTzs4BgWbv8nn1MSXG
sa791gwq46CcOTKASoFHfuFam2LaKC5Hr03J+V4UlMKF0bSV1JuFJbfFp1sh9JLnNYeKCm9Y4IS6
dE28K3Y+fkm/6VcibsXGzsV61kdYt60HgAs4cjqGryzP7M48G8135dp+xlVsHQCTkO6rjnuYsyvp
sXxMxlMVL4aFNkh0EPIVv+9FAyu174CLUB60uqlOZZaXq6xB9VfsJ37rj19daAeQSziGQvShnmdZ
KqPE5vcfvUCOZIZT1tD8lRuMksoq3mKALHlDsW0z0bL5K7Vk7wYF6xuQSGyLhqfoQtAD37xM5lIQ
iB+PNg16jecZm4GT68VKeLpW80lYlcJLLcXI+uCyZqXmm8Am8Fk+kp5aOzH79LvvUl/TxgUTyxL8
5bh5I4q6kTb2Lu1wL8ISeGHCx8FqYX7HmFnmEb+4Utn1N6SxkF53LSpcRDyM+ykjOPkQujfN0Vut
nkjdM56VYYBv+VN8x6JwADATjpmG4gr4tJaMslKgACSb0JdjEJfhRFNrwCbSnidlzyNAzpKRyXac
DhsStMl4/F/L/ff4JFOtvo0G0ao5k4XRWKevXLO7HY6vjTaHZDADbaIZXfWlWKzV28btx9KT8ZBu
EKZe+Pra5RSPis5u6Jls89TzYPF4fVO/wN03VMeUQsD++cJAeYbZYhmuQ/g/czqLmG14PP91T4C3
FDXeCNd2Alp9Vug0HOx1ElubzAuDOXr/vFJq9VkBLW0pZlsJ+X5TDnpiLd0EDaHUEucjbQPTLZ3v
3dtPrZJJIBod5pR8zsgo94QVT/SVn9nbuC5NtUDpLKFkfr/8pPALWlWEqcoLzN97ezi1aifeqU5D
jjOpoS/LCpawbePnGmWP68QZD4jUJPGWMGwSkKtr40cuj/UP0O0OY/UH9PjxImzC/8da3S0mwIRl
oH/10PsFlJtK91tIH7Mhmvm4VipPuarRCSMfv5XYG2/OE2fbjN3u/CoxteOSwT7bZLnww/B49bnp
yV5Ghp6qZQNtDSjJpirsfaPMW685JPtVerFKHCowKQ9j+91gtf9mYiBOynZ0O8ocSnBxpEUJjFdT
VFf0jgpUOi+FcpeQxmph0SvEwd8bgcBExJZTJKrDw0jWF/mb5fQDpV4Xn8TRRvfqRK2xw5jX3NT3
YBB32E2xtbwpnMUIvnMejA/4b5RtSgj8bcMbTsSSsTtoku/bTitSN+WdKG3JCA7nFx3iip5Uvf+B
fKkKW1lyiHWikId3d32pU/IQbFUEuiL1rK6hh6L2piQUOH/gh57S5AJD4x8zU3MSEU57PETHGDuP
r4YBUuavfpsJgimnpdwZ+7Mr27Pla5mrI3bkJFznAVH2IBCKbEZC0TQ9FSCY0G6HG4vSvVhn2YYk
Qlz2vfMSHSCqM+u+Zw/8+8/5g9kBqE3WGlPDrgEKHNBDz9mhLHG802NDWZQQUgKCR+t31NnVrTBg
3KZ0FpWJl9Cv5v3DQ0vQf6l3Pin4R+8RrskRHkwTn1iHQaHe5XgTKMOiVEEaN1Zla7idLPwKEt/H
2svNZd3hx+XH4f/8fmF4nYlO0+gQbGVFAZdplGtAnbn6FcvFNckiJfhnL2ZbBhdISHwt0/j9gwCL
98982JdeHkCS3RfhVK+Z56LYpPtQc94ui4P/lw+E5GuMk8RC7HyCn+4r0WEhRasYtxHlCTf2JQde
wyUf/XQJzbHPwAkSJMWzDPcDfoSThfozyMbdIUMu2rREALeBQO4WZQyquJUdqAKcIZBVz3MHB17g
1OQnlJqkcAC5ROXZlLs/58A6HnBINa57o7RH9oNABQSxdl+REJzQZGOuOlaFXEyeE/KxrwTYW8ta
brz67850pfzNPPjnBYWcAs01SeODzPAqZi/4GzPxVVqsEA2jjO9apJYsnIHSgJ9hk/720MJK2bUa
1HDKEuU1e5QcO8uy1a32EDUjpv740jRZD+q7jDKbVBOo+93SAQ3pitHAzFvlPoxL8cqsBhu+dmZR
9UsIsF2+Kg2ni0AMJB5JAIv52ILOAt0fGmf7Z8DQJbtnIVpHDVDB1VbN0PJTqFE1t1+keBvClFBo
+FOG9igjlA5mHsbpgj7+IOB3vVNf9Oo6bkohKPjd0GwEFwsF86sQLbS2wacYQevFkre+P6ITTDDN
2vraGAz9nMmzC3rGGmDJ4VFjZHXlDA8+4Eagf2rPFwgjkUhlx7vN+gD1GcSiqfL4wfmXGoMwyelz
7LR8fpXAsIpFsMCSAlrxK7vLnpT89JndD/+poTvuYqlKjBBHpTTaRNqkbyuTyyaFPXkasF/lkW30
cfY0MG7FkW8domioEP/NRD3eW/S8Wh3VfJbTfbBjR4tTNd9X+uAf5yPkSecGt6ScE0PAw5JfGnSY
smTiFkmrrPy4prCUV0PzsFMIxdvX5F9sLW+aXU8DZqxPRcyVc4QQNrFcePqWsjrz+5cISJ2dp5Dh
Ve7cl8ysw2O7WSmzFVTkgSTnWGkK03roiMWFnCIJBkTglOa5e9Jc4jcyj1FB22oXRLKuq9NhluK3
06sSceHwo3O5ivIt8/TErBbRjJNj7k60yCG6MIQ6rhJKlwu+0MQNkkt9YLsQczeIUosrkty15yfh
hDT4xH/XJEVx/1HeyNjI+WCx15KopVI/Cbp9e6NgKi3vRqt2CIb02HvUfjO0X2uEwj2mUgtQhWbe
VW2NUrC+R4TSfGOMFYWK4lsWA1E0GpoCjaX7QWlqVVZ5gh/HAki38qv6I+oTkVg07AuD2L6lzFA0
/BhoPiMBsr4z8y4BjQrrtgBvU5RFiyi+/TZlfr5MVTuxaCoQSGDx2xuExyU63sfSZ8ryOTVvsYoi
P+RW5uAiXvyDcQarViAftpbBRv/ddpq3DVR+jp+jTHNplnz5dOBNG8ePgsL6/ssIOc9pd9UAgMgi
JREOB1fCsLF01CBHNG0Qq+sA7N2GPG80h8mSRORpvriFCpXyBrizZdrtEyz7Bg6gLjcIffPlg6E6
62wdhrJJTwc93dEUoagqns9aee1XzWFqvts7VvMJF4TSEiPqFmx+eEb6uUnZbF4C93mIU3v0VmxF
1zSljX+rG4ssHlaANIBYTsdW47U/JzAgizfNd2kPIPSyg8QeTxfa2l9kR2wDVicolj0tHsNUr7iN
ECf8IBEozO77XzorOLfnjJLO5tTZrvDhznOv2BMPDMEXGeKGIkFslHLTkDqNtCXvEI0c8xwbp1Pr
ODb4xFpy2vYAX/HFR+I6G/xCIgsYZSMyJX+AFg2QX4BDsUy2lo9ipS7YRR2VLspYLMvHpIN4cP93
aK6N9BP9rEVnOoe5DWuS5VshamVLfKHH8OBdCNuCKk7Xp4UdFA3sNdupwd5lGw+egOE48B7PQKVF
xe/ivdUTSqTRdQmBfOuqfQn28+7oonH4/dvrHxyybZumEYWE3RQ3A1ucOyYTn0CnIZS0rauruAGs
k6BuMx99uDUl4/lrVxk/GOsIiFAdMvWN6cEuW6SEMwn0ckFZICBFKq9QbI2Lxt0um0kHn9oZfXaV
BjgJ0NVJJ8VncvqjdAOOtqs7Jg7Ra1+cIAWJEOJgleyUA0WYW2qm5RLMs7aMgscyurt2s/ROVrGp
v8vVx+jK/PG4egoJryN5mw4C5Gg8fzHM92UHRk/0Y4iS0joE8Bg6GC4+FjWCNZPxWm2M1DK8yYB5
1rqqVh3CHnJbPRp3sftfGJDC38NV0RDFUw8wTHC+Aby3pZu4G0bvAwI9u/6c3uI4IvCPNr3uh2g4
1NQr4Fv2wXqtv0zUw3R9GSDrDiraKo2mZNwjkfvwcX0hZh7VbIxZVjHT/aNeJf2aIlBTatU6zDkB
ftX60lyc1fHB1FI4aNBgKtY0o1i58+grDuWii/TnCQ4kaHYz0/xXIvROy7SNtSpZ2395NEljNf1R
tnvpcWNGn+p3lCOh8DK4HKLZDYSluhMbkfZuosBDqU+rYjsrzMSE0Cdn2KcB9XCGb49SQyZZCOxG
I7LbXy+qpOYpy1SYyN2qLOqcuA0mKGnvnZBFvKm8rCKH8iskz4n84VW+Qb1dJ+1SCFpWecyXyZbu
hIh/7S9zBFDcDAo1WP8VY49S+AO+8s16EXSjFs1SSQ7jFOO4YEdWKTjt9umvC+UwXZSKUtjbM9Ed
bo7rxlDEaq0f6JMmr9s+9uji+8lumJNesVeH4o4SD3wkfB5fbR5YkuoBG2nZPf1uJlXWSjmg2yUF
VrLFX+57DjRz94a9fCJtl6xgCC2IBhWRQGBE7GEzRv6+lmobVOiRtfBpkwyr1We07uaIqN0TCHng
s0EGtv//PicGunJXfvuvJZ1rrMlIjD9iorwsK2OjVD4y4w516pZyDHBXQI4ByqFuwSmI8mpAFsSf
2rsRAbWCrVRDYF5P+t6u2vgsDnuEY+gikaK0ndjJvv8Svq9jqlYGwSZWfYl4YlAUCeLM3uLEVBMy
ydjDkAN98vOyhUSZ+7Bktf5nF0TF5ZL0CdZjQe5Tv0qCWTgf5LH8/9IZNbIFzLz4AhbHHYDa3Y42
SvnKH+3HGwW/BSa786hfAF0HMYbck8CnQ/+q24BvaSxJDh3LbAYLkbgbMGgu0krLumz3E74kuTvA
ElCDzznZMq0zU9DUCIUv+BbJ62/yqqYHKZpgbzCBvakES6iBi07ejmm27yDQTVyfk0M01Y7CMmrX
GL4dO3m4/L33++1/oMs32y6itF/YQ9Ur/9WSv6Kgm5EByqZtMNJ7xMRG17JFHhrI0aRD
`protect end_protected
