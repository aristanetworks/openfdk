--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
LnuPVH+aF/MDKi+fBye/hdP0ZDEJi8OhwobByNioTmLHoDxHf8dojCHJi/zCXNAndeQZZBaGXVRs
TTqqnclU89+s3To2S1zPG6A8H086XU8LWY1p3fUzS6uS15gRqfVu+o79fSI+ofj1WvZIjML8hb8L
Ua+y3yyPNiXmMuetYBTPn1ahb1IydpIWdbSRRdG6qswuzNT/HT0dD4wCvLtwkLTtPcM4DDZHe3Ft
T5wcFbdT1KIDrBacHUOSOCkGhOdSHDEjxT33sbKb8bBSnwU9xjTbG8tOD9Xqu0uZB5GwudkesOPi
eC/MRNg9kTLh9d6eAMi5+MrcOep4fVI6z2TLYQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="85nT9Pqo9OosbDRo0woV9zuFI+N+S8mxy/JFft7Y3lk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
nyO5HY0A1L+642ThUoz0hCQPz86mz7yGRDMzhJFuMezgr++lZvTU8394WQAEY3Q4MmKKyd1vYOPI
wRYBRrwcCQlgrhpcmhJwUPmkeco4zV9TiL42aE1DcSEFl0s+jEV2TuZzpcWzZXdiZd68tbT53hfN
O/71Y9ixjPriVIYcya3gbrQQS1nVoLrjHaUzpY2XljWT+JIquYENERMfL0Bnu97K0dQEHjy6By1l
VXKGZEr3TwwVwTxV3UYm9j4syd1EPyVVobuEC3rxF/6mgVoGLyxgJqwAHv7wKo64OhjwhjkckASK
wJ3RDEHEULQOwvY94rxZ+Uo9zivUKlNJXDke/A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="t8yu7f18v3V4K12da4bcxHq9296IHIiJLdB2TFypUfw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13888)
`protect data_block
q5ab7fmRGeVrkiT6O2OotRX47pTY0jMWcC87nKDps14iDVImNBoaWKWk3HUoskJWvP0iZ7Zc1xAv
wRLgFaeNJQR0F9GcxsjMSgI4ZrVgqRoEybX4txNXkcV8ZjnkujrRXRBiMXZ632+DYAXsl+CJX3/m
EcdEmG4Xw6pJM70d91Y59Lu9ixXCsM//xWNaZMI+ehKyA3Y5RaLlTcJe2RGAS+up1jsGdmPEtNz1
0G63T3+/bSitGAJUv/sKE6Tv7rQRi3VUmD/PnPRK+ZF0ygXE7CK86YVs17EToTwHRcdh+Nn7Kk6z
xoITE6iYSxXYKBFxN780pKkl2HOsw9ltDk1AjEwCziGEg94ZWWDUGy+sz86zMYuVjHoVrNt15HMd
30lRf99P+3hXoLKtNEDJPYEqU6R4/INzmU9Y4hFC+FyV5nzU/rXPosere+Y5gOyvbuuhkoAVuEN8
3pRO9cTYT/bhfTncBZyJdkRm4i4lr1+DWKd4yk5uko5R32YpDelho0ST8ByMb3As706J8pgUBEPa
98DcctuKjKHIcvQOCvaHjDMdtfxSSg+aSXME4zHFjXxB5UX3/Vu5pps3IEkMIu/CAtEjiEjJFLhQ
M4i9JAJKzBq8n9lKDPwlSCQ3aPb9KL6jj8+/wyW/CkwzuVT3d7b44ukAHhbbBt+k0lEKuSABHryR
iLqWxGiUUvcrBLkUjTempiwm2D+NV/zvWkXQtGxZ1A29lVEq2PFZom8yEty9vHEcYqOKwcAS8Vrh
ZvOL8Bu7PcQUvmpkPh3dKH0QOXwGipCt4sOkKGUx1/YAwrO6cK9Bbsgen1faxb71WYvJmi9Bcoug
WMteuYljkQTNj9RBzwQYRjrERZNdiZYfAoA/yC9inoiJUcJfaPSUjYVlsPUz+E5pao+e9kEo3Dku
NiKpzJDfFLVWaYBQ28p2P27Z3o4lLwzTgb/AqOvE/LT3r7GzCeDxUaJtGfGPSrMlVBOoKXJ+FYX+
2WcX2BTfuUDrCy++/jzSaZDFyUuHnkvBT67Nn7d9yaDBZMVM7iZbbj8JFhrcAG0xEHsM3RIVJJQS
ja23nLu+fUFPVpm/4ir3+POFCo1SOArIEBnbnmtCoQp8t2uGdWgoylefQCSBf6GX7NC6CLOnUzdP
tt0/seWjGMfkshyhEkw3RiyGj0CG2UMtAkl3YdCLHMlMxelbGZsA9K1uBkkkGi/kYSgFWGAffRpd
B96HIecRqetePXDWAU+3gM1wMJf64KDS6SOWqnTPOF0zjG4+a9vYMKc84pyUX1ipA4ruD6XbH3kC
94lZzA3GwUVcZRv20bVBKk+TH5agziUATs3sLSeZofBWv+Kbz3yHFZvk/RffPO4Ic3BJgcUswHRL
Itjqbqcn1KMsdhCnTI4FrWdrgAEOtJPL4thb1QnVa+xvOAaiD0Xr4uTNyfOYGtCwWKW6GbHP/Wo5
fB6U7iPmlQEeTvY2hKscQmCOZfLA9aZ5O9DxtZ+3Wte6P0KICRzfLtfiSHy6YadGt2huYTIP8Xiw
nrVFWCEi/ToC6uljHK7ll5Lqg6NZ2AJdEC4kVOTkrZ/7+at04RVMl5CTsFYKycmFfNtzZCYL+ge9
gxG5UzpIXRwC6nmxcQZy/kW57nC7YGy0ELcavJ6tv5kom1W2VdbV+tAOVThF1fDToA5PTc9l5xV/
RMz165bjAjnxc4i7DuXb0hHMBedp7N1Q3uEFZiATZ3KYChM256w59WpACuEg0u/Pp0aaBAccpekT
novhtNudVTdDZ/CZbFtAtHBNx2/xYT16bKFHrUuqjruJ6hB95MFTwxjT7qP1Jr5mx4J/YAJOXL48
arn+Kqi7etuo2n/mCiQfmZ+hiMvuMavhm27Sc+Fbc4g9t7ORYkB684ayErV6zdB7dCMbAFMYY5gk
UcU3rMJHqOAEDHWH4vWqdPcEPv/vzgQGiH66QG1x29u6nq8zVsbSSrDtDBbaIAbWffmvRUBk5G4o
O/tEu5CgmC4mWiAt8D40//lTNbIhMOzb/pG9MtzY5GYe9Rybk3bRiQhlXIYK4x8ZoyGM6l7TLtGq
GixjBOxIv+hMJmHzKZTRNZEG3fZhc7v3h09ZZ0+ehRF/CG/QAJi8zMkEraLvuz9IDupmG31sLQq+
PlV+I26PLYVYtc62Wek3PI99Z97bJC0oue7OlY86s19DIf6evRbsvIqt7P9Jbb04bjaXd7U/MJcs
ngfmtdjzfS6RVmricB1tC+Weo1LuddcIjeQJ+Gq4esjUTc2V4fb2yDxkgIpcqG1LL6p2WN3gQXE1
Qt45XghxEwvQcIWI5ltDjMbP32t2KrGp6zYmfLF/Tc3IERiv1oQn96KuAz2rz3sy9mL0smZQmZHS
F3o3KHlGYAcCELP0TGZEIY/lK4wG8J7dkc6yFczHTitcyZUE9sVrLTHCEHU7cN1DRTFowrRjTJcq
IqgCjunVJORaBeeX+hA0AyOk5nPOSjXwDBuq/GsOX0VgkqtnXFcKYMdqEtZwJWWLQUDjIDq0onlx
s5HGuXmjrcgtawQO8oxd2eGoG6XuMYQj/1SUfbAJx8v+cxi+KItJC6dU8Nquw82jtbfmYaqPPnL1
Bv3fRL36/varAGQM3ODpvUxAKJsm2dT9jS6j67XKProBWKT6oG4C0bX9ZnurmI2O44Kwei2uSm94
FRunv0pvVyO146UlxyLo+R1X4QGjc3nl9RuYzGsRBLBTI02jfWqFcrx346ISh9sIRzo3hMO2B6Wc
XOzhW8rJ+6RXz62NTqscG+tuENiClKq9pz1BMmaBX+DlC0iLbPK0Sujz/8tooGgXwHJ5m5R3YWZI
HR/lveA2HEuNMHl+H5xGBPOwTnC4nxbkpeUKvHWhs+ylWbKkGBAY0L+It8XjXarr3TLMNRFBtiIu
lgDKMEmciB1yWJVT27x31Cz7R0SvFi7ZNcJQAP35Ej5eh7U89PgeJKbPLiJWC+c4oRsy/zCTYOta
P+plUBMPPvphY6rpN3b78eYwrpFoGx2cWKkZ8szzUREtsH7S+z0jVbpdpCzwqGfPp3E45Q2b1Qzd
GJsdJb1ZrtpFmFdk+FQJanNN4rgd9OwGoINdpPCBBWlAJtE5Ycm4PzvgG3DGWUBC6TGVQd4WoZ/P
Tj3FEqWLt+BU5Wlgw4JNdg2c7jOY7VcBgJJZfpZpDRPh4LtsOl6uSkRH8HaEldt4bflv03XLBVgZ
/pulYYi03pVOBuGiWwPQp8rxRGZZS1HJVZmaZYZNdAvNUmnZ3j9sZTIt4QpZav3hKJafnr1G3Rmd
Jhj/BkD2k5UQW3FaRwald8dY2fBzVh42rlYIpE3Q0C7N+53arN5p/nedmWfgzWlrltH4eic8yi0T
35TxZ7qARdrnsFhFxY3stFGcWdPlSAfm/iLkmVZtqrn9g5kXI90ePwagwa5vofLKMEYr9yJQx36W
TTOsDttHLWAvPXPd6N3HvZ3T5HDBVPtgcRuwMTkPW3DuHnVdCAhiLh9Iub8Jll5luikEjbGz/yuU
LuWywjSgQJaKaFu/o8pbKfmH3yB4B+Y56KS5UaCOsBRZz1sbk1dpbysvXKSkpeGekGU+YxGwJVgo
SUtfWOaczZn4xOnbWCN1KzZLkoaPcWMNmLa0oo3dEcVmhkbtzOr3Y0f+hVMaRG8IEUxAuoZFd5tY
whMCvfTKVuq+uGdgUU8M+GrWN7LJo+FZ+OfWPLOwcjyTovtFouI5qMzgImTwPMB9lXl2pjPqMG4N
PA32PuuBz/JscoIon+TiKYzYmcTWJ0QJIMPhUCnkHAVCKLmyV3/X4oifCC6lk25+bk8APy8AH09C
67BYvBkdJOpIeXdyHXC9txVZjiLSUereBHatVJLdxv0L9ZMLqwwG2TxHIkmqB8WZ/nDonBI4Hlkx
3PcA3JYOXBfOlh17i//TxzW8qorNND3T9zBZifFaQ5K4rWB0UdYTx/xK9kVnm9k8sATomS1KUVdZ
LU/ANZC0TrrKQoZBd477MuBSRjtI14G2BY+PoiEnCcfN4+sYfMQ92kRlxaDeRrMy9TcynbWDX0XC
QgpFxnNYgamJKQa3W9ygkGoGOyTPwuCvFa/D25kLUo3OhkafoeX5CGSh0oKtq/MhYydorbG4jFNQ
S/vlOJMVE2fqcemnjoJDTMYzjZweagjGH6bHzFfAEK/kLRyRnu0B8633U+j0pI2Yk0oRe6VEGZaW
rEnY2hK7GlycSq4etdLpG8SFUzoWabOdteJp+uM4SkTtIh36vNMXycLb7QfrrjYv8li+PVxi1HGY
yY6+jtA9Uv5TreJ8h9B9Yx7JabhCaEbcM8ja73yK1Ie+ZPmhuIfeP4ikF15ul4qdvPfxBfG5L7N2
im2CFuIbtcjMoreYr0Fcc1n6iC9PipJNggXqAl7m0rKXqrzb/jh5DOvBjpftvtZIpnnZ0hw5D+mW
xmYATG9dFTchSzURMBWWzGTbBNj2y73UtN1zcpsiqLkrff0DdLiJ9iY/C7ShspVW9g6DGfgmuYWa
WVef1Ze6y3Px+xGFdOwIS1XbjIMCTOKhvOdn0sjynvP2p4+1+TdsaBoLBl7Y/LCn/HyBhPEgjbOP
sAoyoPkGC7SOvdWynOs96EhuN15gSqljaUSsIZQi/UhMkDgMXs3tmX4h676GSm3XId0XnNB6T/o+
jNwLnFmkQzsh+H0FKGP9G/57g0o6mn00YoERc2LS7K8MzUEfILD677vgS1A13lSD8fhgS3B4fS1i
YRoxdwCkDO/SzotO4qgOIQaWPoitn4K3Ig7qCBbookVKA8C0cQ8gplt6EglON/X3Lf5Law2oduHU
0JbtaByyj4lrdQ1vdqZ3J+8SVKZc5NbPTdD9+ZMmU6J+3nXwFpgGeVL/39lNRGK325f1SAyVB4eS
wzmsiKgBS/wzd4ZkhPmjFms7Btr3r2Ug2ki31VPOkbQJyWM8zCTrlQihNDZhPGQ7JwmFiO7YNs8+
luGi1Xqyjw8vTCmmc+yQdR6fUOJvX5Ii/acy+nhh01K1H1cc9s3BiMBhVf9/jYRPex7W+JrOIOMV
KUPINr5fA8YHzTfsVCEyZFRMi22e8udptZ2CN4NV+Usg/MDC7n/UHrDapR7PFLZS+uzTIRw9Bsf1
kfa7FFOkPt2WAK46RvvUpA6EOGzdT8yb1AL2D1wSje+wz9BD/Y7LaaARvRwhxSsnlBtXuO9NLKh+
sk5MXYNXgUnWuay9b6+Du3b3vO0pfuOTGgS6cjfRdfTHqTupLYlFMu4O3H2OR+JWRJsKi1C2X6EV
xaR2HT1+h/WBMAhj3sBV+NIa4OIQESG16CzIGFl93qUU9o5GlrNaro85adV0BfjOecDlwobxMKH1
889UBiRd0ZjDnE0EmwZYG2sXyQl5ePa/c1Bzaw4KBnGI5c2DxdbGbj0vOxM3QBAklYE5B/XBtbMD
MM4lZ+35Eoc/dlBgimUabGqDBGd+VDP78crjuaK7Hobh7u91Zy/PBGNJ9ugRqy21xdCTnh5MKc5o
23ehqh9oSxQ3GYD/g0RbUosOiBYOzxIkbnJhHa/8pPBVEiORYzVTyp059agGqGcx64A8Ut+UHjOj
Zy6Rp3aa1xDDsogBO0FwmAEnl7MyGrCA1oYbeJqPJBerzPlcmEY6EY3hMCAStCr50LIQqEOa6gl6
sfQXvR7KNPqscn8wpKiDpo5+5zMUmRyg1PwZkLZ7XqUcLmLrMjyFZRB1Q/9eP41faJcBMZqWfsZM
qzZ/CcgdlEIiAuPSOt/OqX5/gTpPxdFnNBqHQeji1LhUr1qMvkyP5XdlqfrjuaP4aIIjktR7rHMt
W//wF27/E1zxN/Bi4gq7829XhvNDPaFn6za46ipuKIqWg/X2woHa46JARSmI4Nge0XilqS9n01U8
ySs+jlqP0cUpwTxJOBqimrdsTik2S4AnWCKJJZ/Rtl+k78Kc14v4mB1qbRQ98ZGKghwDnNGlpvGS
mAuzmid6QA8P0zzq1LzODKWp9aQimMgza0H4D8+HXTHq9734ajJF2rH9AeWd/xAdFc8NsJwbRtzD
Y1JfezA4cFD1p+SGQ8vz5O0ONbP4pDD4ckU8GWwWGlP2+9FibBsO9IMCykBjZxjFgsk5zVKJIFEj
GXy7qqP42yG72CJ7nnqJ38YSzMN8XZmrjs67TQfcJVcwJcAbizOEPl0Y12Ub1DQduJcvJMOX4lKp
5M9sYomATNvU7YZRk0Xr654tM78uvQFTANQ9luNuH7Z2D6dVN1NODm0AXMweK8QahE7yQRenlkiZ
A17Ilnb8F0pJ4Nq5ZMM2XvHAqxLWvqgd5JOZKu2ppHAunH2xj6yeL8DtXCmCcx1dKr7gOPgPmB+4
X+Y+JAbuLJbSIqgY4psq06S22Gg5QJymA6q0zbLV03g1k9E29n3wzBaG6qQv90KH3JbcwMblT3Nb
HM5LL/ngQSVZMYQ+C5XgUxad1rMKFS+deT12UlrRv8uY/Fu0exbgh40X/TGwtzAgeRVd6xYh8Q5p
onp1P7VQYDqO6uiR8F/8n7gJVxpUnlzPk5Vgk1iULxZQNXyiMpX0jbxSRTzeoxFNbq7K19+GC0Zl
ga1aiPEefzgP+O3WAQSNYk27SpQV4tbrvJuwTwZ8MNXRvjSZJcC0uV4y5FWQ/D1R7cyhXbmL/yh0
3Rirfrvo3aX1o6xsbdvY63Qq9tZF/hhrq0pxbEr/3BuK6eDn3w8rqJGOhX5K+1igPCA4nR3lQgfO
zmIOlWeLMP6yZyzkhv/R0/nxJfMb3BL3Dl5j2Uu82XR8oY1Cs/9N0TiTLXxvlOegRNJGznF9gtkM
e7jbJHObIvwhkNRndtHQ90Y16d6xq7ZanfLRBN6DP3gcZTY+oa4Bvh36V+rI56AlE35VmmqvB+iV
+7H7jFeYTfBoeC418j6GbAFvJeeD+tCSh5TklnDkvGPv0ULXGi3XCMXbOYsacBOQcO3H0O/5tsPy
ed7xWNyX2CJttNBCPqJ2p9x11H6f+P7W52nuLEz+gkS2G1iiILJlh/eo6ue7+ugtoge0l5Dj2SeE
O7X/uEQRFlEDYf1WULM5gLOfVMrFcVQ7VeW035sEpp3iqd72IpN53hrB+lVLdHBhDYkVG5+h9PZo
wcNzH0HQgHUve2XFGm2CTOgv4q0FScTM4O4qgKMp1Y84aqvQcWNtO10hLnnwKImKMlijCl5i3lld
oSnBUupyZMRJxPbl96rpXJp6Ofto1aEtYkl/sdmJ724prsn12nHifvFafHHGF1NxevDUpMtBH9IA
pKcP7fyQDfIQgNMVFw5vxi4yKddLatu3uomF2Wo43RSdSnGcyyE52kCtWnucV/Dke3PHxGI7wwz6
LFcJ5GfFyjDy+BH0T8oleG3G5Ex10V+DaHC1sr6eN7kBEVCbBDONsghNO628oYMyHKsXhT+J83YZ
+ES4DPOLUFe5efCvgA34SS++fKmBXaTex3/FYTVlSzCfsjt4NiKVxnHwNBukJK0QlX7jPecL95Fj
5KcdzR+L0CkVJBLh0n7WE2rDLb7J3i+ar02//9StoiVFiEI9KErkqnNpVMJv+YQXZeaQjJazTSIW
3MULeuW5y1ZJWC2Gm4Nez5J3uHuix7s2XZ/+rA/nFROxQnloGX1cCl31u4eC84CkaJXd+RABIpKZ
m24wqhLhMd+nREyOXxbXFTK0DN/Enlua2fOXSLOqr+Dy+iOqZkApOUVBeEb/oT9RXdPp/jpSnCdJ
nmCNQSQbnT3FYQ3Gk1c2fZPO4QE0WFXlky7xkJN1BDzaFBrqBzHk+sgOo8u+occnqpEtmJPk5LkH
Wv2AgYBpveqyfsL2a8XaHO+1SF4Q+Wb9Cuglx7dPSNwQR7WZCqbIySRaTgO6VVqtjatdL60Lx2j+
o3Wc4FmUSUfH27ktvAe9PaBtzvd96vJ2fAfkAu4myT1Noxc0KRWxTw16pb7i/GZFZoG882bakl0V
3jV0Q5F7Pv+iJJn4mJohdgXpPMvHLsZpFhgVXsTFZ8SBPXeEAi3yYG1r/IUXNIoHnOec5Laof/Yv
QhuoB048MHQqYEReEubA/G9p7wCmpBG/pT0fPjpgj/LhH1Q6IGzO/YnM+m1dcNchSSq9MxVzD54P
iz/NezYYL6f2ZgtFyNxXEeajGDXrYE0ynnAyJIdNA5Ei60PBAxPZqN+9c4IGfrMk76S9taDGEDd5
Tkc/c3yYT2arCwGPZPiuSpaUSNiAw50Ts+zcDkoBPyFxaLPHUFkDKUOEzsUFHDfVwGjVe27ZK8WE
i8fon78ZLr1YiCJa+24rffrp0Hpdl+EP9iy5a73l7M9JLr18rAPnC8lTMJ0YFAlVmbvR/jZYbn5G
Gz5Ab8xUhn1JxmI8LPKiCLPlXM+tFL8vpF9h4RZenMXFx8rxDUPHSCHP7aermZoo2r5GIaA0XhN6
2XXc3TvaMukXQsl92x/an5YVCjLhxmCDY6XC2GajQATKncvqTF2tY1DlgB7xAOQCHJ04K04DeRmU
rUalMDOr9qwFibh6m2hUTCqICQbxwnS9EYVV8a13gVSJCFdABMCcV098nXtp6l2ZKpkTMZoCV/QY
yL4k6RQd4AvZ8kLaDpV9q39iPBxAm0rS3brhmmNQqrkHnuMHAz75c6ml+07zxzkEfrr41ZVBsVCO
PRr4kTo6hiO+Zz6KqENCdUd/SI21xRofAfbZkYHHNAQQwoIJNtsDSJafijrunPoM+SkgXKFFOQc0
uOgCBn/pQ5ryngnfaNaaQimfwqxF0avR7lrf/z7k693UJAxDJICsDA+HbOjNatJ7FmtqmYJWIKQr
m3AcYPD4nqd14WXe6ePX/yzim80EPICZ/w9iU5bin3vDck0SCdRe5Tdb0c891ruGZBTFXAKjJESo
+YtJIRNbFg9WaKG9aybpzJzN1eExBifL8rWHIU7+5xV/OowszqzaM3+RJeBasBHZ8sLJ9kxOyvyT
IrQbKp+gjLqT4e/YQH4k8ufmUhDmM3yyVRDuKb56dk+bivQjcHdAJDrMF21zsDza+nJn/Ohjf42/
TifhK5t3GhWOUedJpLgzYC31M6oH5PLlZwV14MNtD/CJqVHxSNpax0wvR6GUCXdJiCC+eNoS6wsU
LQxblLAJxpGw8w0ISVF5WK//Q3mdg8TPHvrW6zYjKrvNRZMxtuPHdQ2Le8YmjgHI+bvswwTbDMT6
XwuBy8inwUx86MmEy3g8kIMRow/5HQ9cLcVWgaUb0u/V77XyT7KzCCurJS1SmFpywn5r3ghkF/qG
VB9JlPiV8EtlGrlIZxXQIwl1TLeCbVd0I/8G7VnNcoF/+Us/1Aemuezrzuqn+kQfRk8OMkuRK4Zc
AmXaD5l54vOPNftqjUtfir5XXTujr5q/V4/79A2NoyHNXI/onEmg09wXU+RdLRZRnhuM+4I7Xy5G
GcSrj33za6ZKrOpFx90T3R8MfUfyFTJBA3C89kdWUIoYY15meQM+iD6Kls6j6Zbw4Kpuhxy3JUCH
MkOJ0tEPTfXh2jMQ1HgoI0mqNIVhCuwrJUTDEzgO3lsSIi+RgJuFCwF9Lz2aLaQUqJ/rfjwCopt7
78LYNurQuVOgjMsZ7BBpP87GaFBran9f1+AzB+xB3xsW6ukZxHNH+JHs6jMR/BxpNgTxiY5tGPR+
bOOnXGe71uNT8ARO+GtFVgR95g+l2vQt5bdaToLC6UbAf3S9SkpSE4sS/RYpiYiog/iHfOPfswN1
5fF3Nqq+EIcru3k9rdigCxAWgwGArYnzae7RYgvRniUGj2tXKFitt4qgrVvRIThYj/nxWU/BxT5C
0P9hsSfa2Npfx6Di89fgA2imyUReu9A9ScYZld5eF1BPS9EI0990WKwZwTmMjpU3byjWTmJbKV9s
Fcd0nAZ9A/s8273IMZ9sEFxTz3QvnlVJYeTv5QjNo676cR8JQhl/G5pH5RgDJ5F6qzvDmjQwcPmt
7+Co7dLR+XuL+77uL+ya80855qfNaOB/NmvrLsOLDOt427PSJx5Lxfp4zA0lcC02mHV2sfvWGqGV
1MaYYQ174CM/BfA9Khd/yKQZCbrSkdPne+2uw26k9eJVX+Y/1QammkNR8R5reYe7LyoMfQlHpti1
iTPxnUaZIl9csQtOJiYJ1y51aKlj+ITzP74kT8mEtEZCL+csnwqpbMnA2EvDFPBcTDsIshJyY16I
dOFb7RCK7GK1vBFX7AhcAa82G1sEhzgfUogB1yznKb3CFJm6+fgQkToun4k/txm/577Nkz3bSimS
pjtvX/jwcqQtZnQiN7ecqPdznq+usNrP/0un9C8M5eB5St4k3yhTOy/Y0t9auu8HVoRmL54WMs5b
wLJLqICp1V4UQ5ui8SrvhNTTQ39H1KBRgMlP4eLztUNkL3KcSmBFCQE+czpb1StXbVl104miwkR7
eDAzpsDHLUAFmMN9A4t9G7ZFPUNqK22ehQq9WSvBsgaNe1yQfzMhixcFQf5IbPlmNa9m+MKb7v/F
LsODgytnH7Jn/TejUjMcBIjluOXi/SMOuIaBRsThJ5q++FH4H7hnLPVCmI509rmT4OjyjnjQYca2
3+YsC5iYZiXrHaHzgGvpzJQt3joufE7mIXzfK1hMQtL/bPnUVKEraKVARGYQWXkASMJUgU2DVUKT
yR4NKcPyZefmSpF8tcmMPsoMZydXNLxj5JwNpvD2StKEi7vTiYCGYK03ZMpWHcMsrVdXjqyxPogg
rbnXIQACtqQn4xAXnfBezVlW3YM8iTtSmKJ6bc9q4FXpArvlIGpThlarIVxKSO/Z/ZweksXHJoEU
nDFRpcc5ic3LkeiuKEB/xEgoDKkPEPCbZGvA454lRB24VscbA7kzkgyNYcoK8yyNf++n3/uhWray
kja7QmJ6ezLyykpu6hPL/ndwOdkQjFdD8kRkRwOJc3gT7dxRQ0a/FRE9PlkYhu3XmRBdTsNfgOua
D5omsJnz5cJwODJICUiRmYMN+gDETib8O7c2aKc1bLuViVQkAjBQSSAqaPezGY6vZ7F3EW/MR+1j
usfQGrd2W/pTSHHQApRYSuVIULAmzvk8O5Z7Tsfiygr0mWFOqricw9dkQZIfmVD88b1N5rSu6r6W
HdHtombhYJNz333gbi/m4WGj6k469SBL61Tu2Gi0FSssSiyTqnS639HFBg3Ww6cU0jTa0lGJu0tK
80U7n8I4tWhPKdACOPIcxFANSXEcRIAMR6CkCJyPwNc2KZFbz2G1kCNZWU6UxRKyQT6caM1vQ9fk
pbSiuh45gXW68IIZZ1IMk5N5ioConGG7RoQJfLiAHqZhTO9NuRoo/SNzy11KkQS/7DMsv+vd8rcr
hy9TeBNWfe5IvQ2+jzWuMoJ8r5ZLZXiugFlmAmnZy9Ge3CFJAMehYR/m1v/X7dvs7cq1Pu1BRToG
DuTc+IHv4pKaIRdkH6MHCsIRtvLi3y/fAQKUFi+psq5+j8F/DTxUiEylXVdCj1mwAi/DeDC9j4Sp
11H9uOiK9ySMVH9r/tJBL+r9mkOAekYEalY6T+JD6WGfWkBKI4dFqqz7wqdBzdoYmsS6xpSDc4zb
a5WRATxwVGNKrt8JiXphIE9J2JZtnLh/f9bpqVSPFk7FPBCpnfkBZaJH7aQ1PB+J5OJvarRGQLcz
x7v3+QyjqakIydi0xAD/SMdfwcHuLUubrahoqa2GG4a2E8/NKzh8kxstEgh7JDfeaLyF7B1WsS6P
nBQEb9ZNo/89MrEuRKJSOGh4TURNuWoUMyajannRkFlS9EGFIgQNi4Vv7Cnjts8cO5AVhGszzE+t
2YNWVpjqFy92w7vHZEWFXPCuSCGNtDWT41A+xiV1XvtdJDGIY5nbE2ifM4tUmjywtBywJRFIJzY4
swuX+r6/fZbR9nH3+M0fXSPUOMwzufHa4kW2uYqs5MqtQXnrZzeELXgsSCVnx6Js05IcLa2LKxJ7
R4HVNuJ8b2HQOz14ER1XaFvAGgvUGQsx28yyXpiq9jDwGbiKFRcu8emPUcb0rcOHyyzOA0S9rObL
eOIzKpR4k69ZJ84Hk4XjaxGLw26mDObZtDt25yGPIGlEAwNNPXJCnrcrrUtzN48GILOOB48MnnU9
UYSa8QluQKAJQ5HXQEHtiUSp9T0IhYXZL43UCyrJ7sEzIeGW35dI+TDZ3HlC0dTh3uTyzbPgJ5qG
VJpskTxTP7ioKw+Bc5dSgdcwYbh0jYjXGAUd0ekJtTLsTyzbIC2rS9B08nQDOjEmBKvUnv7w2YWG
1kuO8tDP3M9cE2h+bdRI6Lj96EJLxY23+qVKTBWfYBj+tcZmTTKywG0vE+8DfQnIqQWxpas9kE3n
yHFlls8q4NF/pl3qTA+gzwR68nIAM5LkKqzUfKMlUQidTv4X4vQZW8uzv18dwvA9nzd5EeC7Welk
MgjPfKJEyLphywD6GE0z0YRofcke1zA9kXWqxAdx4Y7X24JhbrUNHaTTORlRxaVPhIIfxkpFSN4u
J7zFIIhEVIWjsq4/+c6PolzCkcUBRHsiaDo43UOyiFgu6oAf+jYuM0lzY6hpplsTQb5fuyzDH348
luPQ/4/oR3Gz7Y4wnSKsLH+HUbM9uOYyuWk5KMZxgeyIIHdeEe9+IqF0w+u+OGEQ+3GPPIM9zb+a
30ho2ttqKDXB2c031sfTjr6CGHcR6WNhnDiXw9Wg8gDSbmQ0ZdI8IBO0STTvrao9uM+XBcjvcNyH
Ul0aAqOkBboMUwGnwr1UaQT1YF5mVzuCCfmaF6rSnaYsWHxNEP41TRUaDUMv4K8s5+MQQ275SUPo
p6QORacnYw3k7gavRvk0iTwBHHxyOfOrAMmNPgfmjz/lOV+3R3oUHsa57nTZguN1Gbgks93miquG
6qsjH0vFL418mboqwBocrfxmi9PBlB9aHd5jakRtsEgFB8eNsT0DnRCW8Z31EeU256rmXRYxeQsV
0Nb3230XhaPnuSH9hLoZRQ3Xvc4IXzV8BsM2W8pkeAZXRXixdmLG6jN/u+D1KFUpkasTxCtGQfYg
oWj0Bsohg/vOEgcWEGgr+HwUV+52XjMiuxhlR+4r47UDPOfAWALbVTHUvjJgNvH/WeL+C5ZVHzhG
Bz4Wvd/oTbOSbDGB4i/OcusnU5TSRHCZHbrfrijAsvcgH8aAV0cXKgmIrPFOy5iS/LN4zpLGZhuo
76uDt1wmOlFu8YR5tEXG0J65uWhblFy5K7ZI6f53ryX5CA83mQsYKEkpX9H/EDbbUJjlXUzwaDZ0
Kl+mFK8jpQkMbB6E3NozOvRvhhxjw4aXqznVB39MmxkplJxdpIbSQFYVhB7iiqRSXeKHnXpyzbb1
nsV2lVAXgZWSwAgU+2TNdxjse1McZSA81CqGq8tKr0lqQNwnutrYKuQxA0eaxsiQ/vq+QLIhMoVN
Ja5zlg88/qy/g6t9dACXzf358fstrf6gfBN29Hej3tgm+OjvAoHQcGNevxSX6mKYoo1J0+haXNkf
Vmz3dI9NkeV1igi5xejTFDCjHK1H09aRlsSoNEVmYvvbRF7Gth7upkrfs1lcdh7CTGSGAq13OCXU
WwX/WVc+E2jQqgHxnLya7YdiEU9sxWKFQ9RisF+riGdYlpO409dJSGcVBqg0cJvntirlgQO1uX/r
k9qMkIVztr72pszAfpioYIpAkLSWVWc4j7VPSDiPdnhooQAN1ne28xLhSA4spWm4RH7Ckp3UKMa8
F+AtUgmf3UA1eCxew5NP9cfIbXKaHHjJv8yUeiBJiixY5jsQvrntdGvuKZngeGyW8APaEbjvg9Uo
qWtHKyMgez/gkxuVNl3okBEpYkADAIYOmZk1uJbkWBdJcyYxTF55PAW45D2Na+X+uKpz00lbctaw
A/lTjiq5xeSRrqkNcNpf8fADA2AYrADVSTzI/XfU791tSsVHP39xAHo13ffK6vAIx7NzrvEetfxr
TKbvRBcXvCNKLuEV6xn0g9fB9bBwQP6sbpzML/B4Aqr0Tht0o40f/Gk2FbOqCosnWQnt2361bygk
MDKUf4TxXeOFIgjyPLmA7BYxJn9lpIDAoAtqyjQE34Iwng0AuUDZ9eWObMoa9M/TXb4ITY4BxMgF
a8k8/+EHD6Hbcpo7oe/C7eOd/qzcVhQzOL2Cmg5Sv6+lOUtKp7plE3xvQFc7f7CJhffo6SvCBO9z
1cx472JRlF1/IRxvuyM265ivcsXQobia/wJiMoPlraxdjxlQEs8wz3uiE7VJ4Pb5u/ipmwPe3ZzD
hY/g1IJaGz/vzVcNOvctX0dElRk5Idhexd0t6hDIYlXWrt24xNfrJ1gia+vKTU4B4ZtffrZHDVov
2aZkz4sdGAJMmKxAvvLadOMXYXU5N2aGoc9e5ei5Ban9JQaaffLMS8fCPLGLbleKyHdpjNQIJr0l
q9CmteF9flLa5Tq5wyAGG4J4rZqPvn5MqSszmlq5bODqb9ELUfnp7hfVWpfbG+y81uair9zrVYC+
0awimPOBDVGps+/xyPjJV4hXiwatUwBdWtiHsn7rP7SL6mZPnddFmYpqQnUL1Nb5eUiKDCcmWMNJ
DxwsNXBvneyGcU6/x+Sr8x2fW9ILnvzenfHyNgo9EjJYKQYh7RPfm9QVAMFpA9v6iA3WFOOIam4p
itunCRwbiKjVOVY+ev5A4plAmfsoAS0olIeCBcLvEiGHTWXQA+ne1ipU+tP9bxDC6DjHexsV6fRY
oxpMwzbxsmZhsz8msT9EEc37lzjNmEZ+V8l3t6LWgt+GiSJ6Z+612EfHgseYEtQUFLpnnrcUzVTC
FOlTA0ihtuP9cqNVSOIe4hTP+wzYpW60UC5fIyA6wa/h5BoZqLFCOsFS9PN5VMplEN3z9uRn4d81
KBLSWuyntQWBUXf7xjmxpHQFMIGwpYH8XEEgS0PaRhfI6Ys4M4YTCShc0iAVur1GNvG98WIHts3j
T6DUe5MaKrVwLYt80sZiu1fYORh6fH7P9DByjeZNkucO2U+o8oSSpNhbi2ygJowrI/uJsOv2bW1a
xhj1twWl2/lkAWyVFQEDZbVMuVSF9fKttbsartXxknc5uYi4R18WSZWBuBr39QyqMdXS7KRGuV8n
FXNPuGjmfhZKjQCWGK0ZhO6FwEDDTDA2rNCgGRbR1pIMHy9nHX7vHOpYxx+Q80iU5I/UnVurBhKQ
3yVQCV9y5Dq/cnYkV1b0KzWDKzSImUbp0RGg2CdpI/HHAfEggofC9iZ69JpFGqHi/W+MgRpzHSqw
WXADKBlp3jYrupffxzqWo5njAO1iNiRKETcQ4bSk1q/R6yjQafNlQ4vjJ5n1TZ7jA2n40+xQ/Uf7
WgasotCU2czBnMhtOMk8chuSH5bsybVz7UZXjaDMBHbJlfETeSFlyY6rJ2B9EeQ1ipek5fiEfR/T
co0LadWXrv3dBPeof5I31yBTZ9FpEgAjC3rFk24vIoGxDCoQPNeLUmFXIrtcHj1Gr5U8IJB58Zjw
gBBiaNYRnIexEedfMSglKfuasNeGnzndQHeGZhxMr2HtHkPln8Gr2iXdZi7MkZWAVpyVzHtx+nQw
BwVsvU2aUzqGfDFP/AiY1swOFagIssRvCXzxoDwderbrA5pg9WpZwI7jdD09cIt7y1jRBNSPqYIF
JCN+2GdILGE+P5WBnZ1WaiVSPNsCECcm9HY3TNn2iJn2d190oFPm1Zq0WrnPRo31oX1mf6J29cqz
caxUoJ0TlfzcalGe6nX1ldijdvwcnSdnTaMF/s2ydLBd/otBGR5k3F834DqI3ZecHIjrChD9DXKX
lCbGZIJP6C0QAor6xvkQi+s15SYpUzqSUCqcyZ9Y4oC72l07VnZVzrSu3nEzs+XhuXxn0lRCAiDW
3zh0eyx6iWO9U5AO/rUm3hdVc4fK616Y2JTyNezLVM1lRgZ6qJ4FKCY2nhVXPp1tycxqO8kXyWsN
p61F9RpK0Cf3Fd+C7v3nkZ3BpP3y7Gj50oUWcmmdTCQPFTrfQx8M4cG4zouklEjjArYUpKvBVxZL
vfezgAEWlJ2Fxo9RQZEaIQaT6k+s7IzUcyPTuZ3X5ZTVoUOX8y9b7GrFxEX4oqJGsRqhl2h5Mzci
1erHhce6ysIV+msHtImwVmGB/4YZf7BbE1huiI44vj1xnlaMQrH1wtcUOx/oqK27oxkGUAOM779X
RpF2DIGr2BxwsCkxsqS4inyPi5piafJvFgwikaf/wTSYlj3sldMb/u/Eae/OLBi6QzVUkLbF14ZF
Bxzg5DYtEYh3iVZsrTW5In1t+N2Mu+rXuTa9RXE6R8FLPinIkfhwB8M61B/Pk/OAQPVEuMsIWlE+
+9ayNZX+R7ERs/iAIKHv8EsIE6fKsfGEkTJCS6WxEldFYIcFO89coCzAa27Vvf9WfWaadfRhyz8d
KLvam1sY7hpLT//+nKVfOLxsfC6WPGBjjQoPowNA2aSxp/RlAY/8WVkwe26iC03yTUaQW+RMV4iE
lqu+buwFL9eq3Lb94BMievhlzB80TUv0A6TdfG15laqYyFufSAO7onNZEUIsV2Eo36kFHkvPt3U7
TgYv9K9nutKBw5/UrX7xTGQP3ef1mm+KB/H2WVixgfD5zxBY0phjioksTe5eG5q5EcUfL7wHMM3o
fyJbo1Y3rYPqGUwofDTDk9CnebxzKmwJABzi91NuEAAAT3qiyX4djeDXLmfATGTjk79Bz5gzdTt/
/z9Xlirj4CLVdULs6c05oq5dy9jqPK2QSMDbUAFsvDGIDihoC9vxjEofou+/wpevZsSJr39No4kJ
AnMXkG4en7IEZ1edC1N0kT6FW5GjuGCcLOiF6hUNe0SWepZ1Jbl5aAIujF4J+GCEXxRI82r4WgvT
L+FBXX+wJYXrIz5YHsKAaZBvgvxt3F/Aa0yNRJwhSVneAnlKZA+5aTC9MTeYiI3PxWqjdTiaorkT
d5SzL+aaAzcboBuBbzHgfn0B8BXU+BY7CyvcRzeAxupDGeEmlK4ka/DDO6iwOHh+lI7yo6qa28JC
oSAF2mBr2vvnpSw24TP330LtJJilZxoRNCxzeBxFmofvyh5/YDDBh/sYs5c9S7QfDg5P+bcYRh1V
LxRxzOo69bYIhUk5w57MHETY13DAcKYbNzM6Njt7G1ZlyEQO+vcT4Fvz4KFGzU4i6MLBksrGzUMF
YL8qmslUArWOmKv6TKzElSCEtxhaj1kHOTzeH34KiUcD3Zupb59V2IiWUG9JJlCbvJNRIIkkcp6A
xCOsB8v5DAhyZ+TkKOKNIHdRBbOW9bEOJ/a/PtkJ5VfuXgBkJ5bLLQaBdRfCOt2QgcNcJxE6eThw
mCplzCW/EwDNj+SPAMPcr1V2d05VdL8qOzy9ltG1HAb5T2ToecWM2zrEJcrv+l5a+ZM6IvCzQuPZ
id+ciaZ+QxttmaRKQek218HjKSe8H+xtc4iIxSLXGs0Y48rUACgJfX1MfhkmAkmkawF4tBqyfMOr
g6F3bi92PdYzzYnLA/LVjTew8ZPv158ADgQFfVcnaS6R6URyVK/25JJGmtT2w4VxH/TXjQn5n1XJ
KdCXvvr5ip8H/k/PMHr6CDcdNGV9FkbGyfd6ScLGxljMKq5rddat1HNmF/uAARZ4s/sBm1x/yYom
huUlJ/L9wmf8Nhvi5u5Ao+rioGQmqRJewLZyxsl/HYDBeOdmrKIYHP6Z7HBKRohasUeWkcPuY/Cc
Oi2qmN0LKYhzdNuhtuiySJ6XEdWn4CkF3Tu5UDU/fB8clFTCVve+Ejy29ANp/s7zDWC4hCPfaoSr
UOyBKG0AsvDm3VB283kEIwGilQnjLySBLKEwRd5PjXUKAXrFgIhsupSs/kzZ0XZaxMHzV/JU2mWs
0FrrXh4m3rWDHKRF9xcHYYpQy5SBxwhTyaoSfo4rAS4ah/ejV9FA76O/Qa/kzh+GRyP044mRKihJ
xvzxUpTtI/WsHpYAE7YyJ8ShvVwxrFmS110J1BgofGsgwJqye5ftlmBcVobYedFwdSFEeCGWZkBh
/8VGnmp4vAVlybkT4oiyjrqU7HobTmdKxNYyYnfX5GPWcSClH/ksRm3qhBrkCen4FiVGt0MqEvG5
RHfSOJSaQ6biiBxWKI9w1rIbkXokevYdPHl2eYghTxaR6CVavZO0Zjsia7371+W/LmoSjxWbL0Ja
k63N7F+4s+iOdfk2JAePeUtnqM0EoL0vNfvGgw1VBy3trr2p57fB4GLGii349vEnmMCD0pEJr+9Q
OFfE3ah+FeHMVXpyd6ZZqDfJh7smH3HUus5ROoj55dTjQZZ3MdojM2xhmqHHu7R8ZTvG61Ld9Y88
UxKSRAnxITNqARMf5Dzlp0lZ3w0tUv6fSyzkVv3gEp+YDgWhUA0AYvXtaWkiPGnqrqwbuOMAmQ9t
OUv3t1HJu2RFY0pau9UEhZLLr5TAljvVfCVdRm0C4wyyQbkHN3UWr1UasBu220ntuTih7oM6UfXn
t/8u9HenP88mhQ3CwUuZwFELCGT/sZZFhj78yeEPjPxeikYg/Z0xP3nIp/9vsSXkA1Mqgwaperbl
XzMqGSFTL5aUjx9tJLZhtJb2KMRGXRkpXP9xKDM3xSDO89DyaKUWl5Tn4/5JXMX94HBtEv+KP5kI
Y3EaOcD4pktWPo4CRX4zyDLbAouFWTGYVG2m2gnJ+NH6vlJ+Ow==
`protect end_protected
