--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
eB6aWqmld7AugJfO0d87if8GnT6TngKgAMUCu4JOGjnAj7c+foFnSLozkkfyacBN7WIFeiy5yYSD
Aga/32hcjC3q3ARA2LaAR7astMTbYjSvWPjzOHmfv+kY/uRh/1T9udBNLryRgLRsyjl3R44lt4sw
FZzK5az+gFxxlzkVLSIjfC8gSE29mvkDw5aakBN7/Umxmj/jVUC5QZmYFNu3EuPWuRjbZ5kdHRAp
qMh3WKRsj9X+Z8Bh/1oo2zf0yUhETfjciUHU6n2QgAURZv3DSaUovWiPm5EOLNce88qkBt5beKFI
8nYmiOhyZGaDl9DPpoHzgLQIaj3Ab6F5L/Lcdg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="nejo5KmFxzrcMqtBQvbFVVwEctRU/oAUQiTmG4C3jQs="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
nU2zwtLr+ex/H2uY8NI+5oRU6RpQZS6j1wfhGOf3X8i8NblKHzTuXl7uLWPeLFe6ZAt7s3kweb/h
kI6EpiS+2CARdsr49He7qKYTxt4SJqmo2KW1gpRWUa9zQZyPFvy2DB/Yndn96bJTGV7C+W2Yw1dD
5R+BAF1PxpYCrjsbV+SPeLZJate5++2W6sHeTsI97OTSCW41yMvaXcABUycz2hNPevkTfiGQCOJs
jE3frosAiaFWAJ8FsG7T2pyk5PJ2w6YO3uJ1b68k7Gc/zCF4G8ktr7FYceQVC7RjWM6f4regxdWh
NrhhunJFrABF+g990RAWbObe1xSE5zNu2AUsKA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="01W3Qv1s8ZCLiEsGETrcgrZxgODqmguXzDzpbdl1P/g="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2720)
`protect data_block
iO/Gtyx7frfqd/V6WzaQYeKgFTufa4vwDVxFcc7HDlsByLwW+aAGga4ugwI0ESwVwwxwKB8x7G+q
xltsjDhBjGQbKlONc2hkZaeElCWN+HMiRHpt5GQ/2LzZR9cOHrd/PBGz78mvD6vUPPOyTwaoSUTO
YK1hwTxPHEv2ZrENdBOjGObh+/Brns8iFc47wrWC7D4W26tXgDWAA3ntzeqFZ1qO9IT/iERhxEIz
mXZkPKkzqx4DiPWkMeIhm3b0hHsQQZgnnBz01R+R+IvfBJ1N6GcZHm1qtmuih7LDi2keS6RHwKuS
3M08HC2L4Y1tL/6uH6FC29ThLvGbPEDeZ2tkzFXqhifeHpdlmfDC5OV+IKMLnH0StTSfxirjKxtV
NeAgvECfTXUscUSAAVHOf/9nwN1Z2LjiTKRRdy/GOZr+B+ak+WOPufGcZoRPv1TRFqhlGS7+4XPE
u3/nLIEuKyxFYF+LNEUnQ1TEk9Qiu9ZLIJVj28UVaaJRVw96UGD6TG2dLJaydx7GsASAKdzFkvWk
DuGPs3LROwCAw88bg3N/NovKBHcLIWMkGTDQGcLiSt1poQk4UYH5eFrI9iUE9/YTNwrKXx+rq81p
/yOniLV7VaYMKjeRhzRnWEWot0UTLscRy80Wp/eeCwjkqDFyb4FCBG7G646RZu7ets/TK2nI5TIp
MR/9ImpPYCVIwQ0+3AxgKhOLF/PZ8v3TKwlSL15bgxr8bWZ+i5GgRofQfYRnffKBVHawKmcXNsrj
TZJtikt2ZQyqx6Gg7nRtX2u9wItj+Jz021J35ZHxOrvcGMyM5l/3qvH8B/wkWtO27ZV1i9magL9W
lVApCXrvXQP4vEERzVLR1rujMspJJgdfvVB5nhC+DUGoYoryxWOnNJm4EduxUSGpFlNbKl0ZaYYn
MtMMz/H3lw+xvaGrlsiWjk3y5K5DSmWLho+NKt+FDNP0f5n9Ce66v7qI+9LweUS2pvcWkMhTXrU0
/uyWicOqQiTuzOuTplMkGBLrl7fuCmZzF1aYjiJthR1lFWD437uyG4rjH6389Yk2oOFhF0AYHNOo
EU0rSweuFFiW8/TH8eagJeYFeBJi6Z7DJf52DJSV6eVp5WdPodppJ7a0fxYOM6zNIBWKy11hfqjz
F/n9cSckmDQsEyql/N6I8wVjMt2hPE/fbEhUeW/+uQ9ujOCf6U+GsCaVM0NtaYaLggYNP5WZkVMW
wtmHAbVW+kiNmnDfh/tbiMIlwHOVml9g5NHNbd40qaVWAm7e9s9TMCM80r9jy2GSynu/Lf0D86wg
ua2vba1fn9fnvUgqewyiNmZbPFn+lmkAGbv6UQ6tiXoYR/OsB+lyfvGeMbnvCowsDN11lC0wMtGJ
wL7xAwMaqAoQOZpEcPFiCLhJZ24ShXY9lJWlMbL0e1fe775eeFAB6Vfrk6JWv7DR/qvf7bxhU+/e
AEO5kdNEzZurVawLu4k5upeiEj2X1/Ynws11aPBG1OGLwGq1wwhTt1mMfTREHgsAuVq/Xkadtb/q
JyREc5MXIUylytE1mX80k0SQ9x+PLvl6jZeCPU+SrUMdqBsIEiWbQutRUuG7abdLAj9aXuii3OJX
x7uBSmSR0vliFms65gvivfQn6YdtJdV/N1WX0Bd9h8iltO84u3DUKI/KpySg08LwdoHzE2S611H7
Lq5hYDgxllT4Kh/tefY5sLEP/t4s4nZP/muq++7aAOM2UarZUps7iSy0dpUHDfzTJAQ7LwEn0/WO
wVk1yHLuu9aDW/zr2rgih6g7hD9s4jY3PN+9gdOFcdBT8Cq7zKywt2V4sDuaft1oLMSPJ4g9qhC2
VuagZosBEe6CZhbcedgZEbXBWW1Sc8BGpq8aGXJtcaD6VKRwGWFj8seszjqT09qIRNWKm2uUo4ww
jLiwjdy5zo7flY+QfQvZLGKQgm4isREAPLVhgsLXzSnQCb4UhWNbpDiraqUeea4G0RLjpFgzJDav
/p/ja6vWQ/yb+bvqX3edC9SbDd8scO/rdoWjNWv84dvitaK7L3Uq/W/zv521o/ji7erauGbzim9j
2nxd81hRgGdylj1WTgh5Q9WhW0sV6XK7K2NQWiMIzHIo8QD44o5GEbvANjZfDrVBcrV6e/mF7zMG
QKGsGOPYn3bCuwep5DdRFAKGZH+OZqrw3inY23XJ/r7teccC4yYT/5tzHySKfw1VY/o0G5iClEc9
nrYD8ZoZlAw75AX5z8xSJ1KvfeqhHz2GYcl7iG2OqfALfFJNEiczJTxdEvcmSLNGFhgRcVVUdygt
6Ju5PQ5040Qc1rTFIHhAVZVjNVEpwrPP57/eURLqXHMGCPqBL4BSqpxrcdps8Em1lp7mkAj9JpAH
8x5bQCGshKu6d/hcBrtSHE9WC+vjVNv3tf5/7PEXeOMNURwptpZBIXRq1U/8Pp6K7odNXkPz/IPQ
tqK6z4b+4/uowX6OI2KUgpg+OYiVLakyq11AIDhP1qnsJsezfblLEvGu1TYVR5t7Svl1hJm4l6BU
KMj23DgpJmhkFI36MdcQPgbvCSZJLaJBswhcSCG59C20SH1uHDaXHGQAACwsrwKEoWN8Yznw7I4F
37SqoiA/BBLp7LmNidvV9Ssi0YgwQKkezcsswOQ4F1LiyLlRJZmdqKzLIotwcJiVfY0CowoIfJda
LbkFt50Yr4wI8TS7TZ8xS6AS2uu+Up5yIvoSacVDRYceNZvGzUc1Ll22giMToIwBHRvFkU3oYOO5
bzlZGwdmZshf9Xt5DdugJ03qr137YwzKBiMJxK/6U1g/yPUyE79XinwXRGOeHXIVge4KL9YaVpnh
zwe9uthW1LKT23vTlYOU7fW71Cax2Fx75oEh8jpfZKW0yeJbn1RivjsIZuX9YFxrVbBubjWsC4A4
+y31JzfA0+IZveDdMJSTrii4qM5FAbsJ9gmMk8mXFe5SOnV0jMGbSp1F7Agq8xC7p+V3y6YHMdlE
lgrJnjPjks/wkVDsT1VfB84WqtRQ7Pc89Jrw/z0PeaCQDTiR7ndYh60bidb0ejY+ZPjIwukQijZv
sJFmJJKO1wYC39v5iwkPW5XmtsrMqlx1Fq6EK3yaFU2m9WKozY52RfGzVYoe0/caCIBh7Z5HB5WP
nohSgYDj1AlB/Lfc++4PIG6YP7Q6c3FLl826bWrezCQ2bPISQdm1Gi7uauLJG1TMCNjuH27vWXPa
TOLWgd+xlBXwcLnhxs6eJyHkiBKbwug1VjsLa6AaWKR3acT2BxxSmIHdnOGCVGgB/Ku5sTA+aNG3
TJo6YnG2HtUdUctM+tSdzJGe0k9SUbYLUYu6izJw+WRJIIgOktmr00WMdPCasF9GekaWsaViur2v
Iogq3MwqQlBonDaEDIhewdACD96Y5uqbvxMPZ+1VejIgg1rYi/ezpfafMfi7A6ojHbqWI4woqylV
o9ioMcDMwnm/B+9AUHeEop7+Yj3ey4NxWHcuL3tepYYQVPTsNOGxjw32k774hx2Y6JkTnzfwEbS3
Dkovd83G3SkB0X/75YUkg62xpSime+uNGg795jWsTnz0xfuKfFZtAeMGfwUzx6WNq4aeTIquY9WU
EDuAdOZBAL/iQSC0zgNARctDKPYvvMLkwZPS2PUsyg3D/2eiSVfW7P4=
`protect end_protected
