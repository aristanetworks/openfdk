--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
KySGaDtXA3VFb+xSGm/FKOYZ5I64p4G++Ya/cV0yZIHIMzvt3mDltVXiZSMwAFXnzy/qUdiEOvbv
MqLjNAXzSGGvPRWMj89myyKAgOlT3CsAe9xjlNI4hhAxb+5R87e83DxLdGNemzaBE6kfFGdi/YbD
zImzwfG4S1UOZAd3qPjk5xaw+hqFWxJrz4BAFOrB8WqyxUJUYIKUJvtazYRL1fPh8jBVB5vJJZIE
ZTCLwuKC70LWNFhM7g4f+TdTDVQrcy+9S2zU+L0zIcJQ+3ovEYbksqd807SJYdQFVUlDZrRhC7aJ
wVSxr+aKZ8VhZ/iPj7YZFRPE3j7fo6n4+HLTlQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="M2Yui/Qr86xrQ6OZz1iqnq5uRhabgSQRlELG+V2GFs4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
o01pRoA4Wvwjw2O0ISnZm3bC/2C+7aULb0/90Ez2niGrbeOejjqiflpT2OYf3+AoRJkQv1BMAIkE
SLB+HAxYguN6/n/TT45BpItBVzDVKzCQvQ+4b1ZdNDmGjaApD2tt61GqqWobY8EUInnuRLlRHTK+
R+tuNc8vChBzB8rHbQRE1RIydYwSKIVDCSKDTshAzsF/gfa6hjH9oH6Ce9r+D50tHez7g+4aCwdK
WZ08BmaWP13/QtdRWXsvNIb+CM4O2hXaXhKHsDF23gdY1QHIFFgXaNRLH23CzkgC8y+mBP0WbI6m
6Hd3eq+jrsb1NtRmntbcn2y+DFXeISPbGI6U+g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="AaFWrhy37vzpGl4LN0aW+GlZo01h7/BfMO3A8h3uxfY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7280)
`protect data_block
W4WKboA7aDp6uORQN9BpXyg1FeaJ463xl9vfN8+URu+LCA2Mt7j27e+LdOOFvLF/UHpUAwxQUtki
8rph4xT7362YpMAd5YRcwWkrdhPzyIhfQxAFMZjAHpUTbx/kqmn/PSfFIOn2Fl39JpFgryPGdnB/
lOdZzAP3Dux+9oAjfSc1knec8qPYnZi1PTi1H4YDHF+69T8EXQ3u1VcJefeGhg9VFFkC7iLmUMDf
/aXv2r9pdILjkVxrv0WDZ93rqPM31YYJ/wdAoHpD2Ng/BHFnWbqclgb1WbpwamUJsCH38DDBn02k
U+3Y7fVVdXK663ndZcL86vz4CMTMPn3cUqtd7hBXquw76o7wLBbv7PhGL9Os7VgkqGYIaRDBpaU8
XIk307LhzUSu6U5gxXepBTnVXRwsK59vRMjqJJ3eTXLEv/dc6FxoBo0Cqj2YzFr2J8UyoneXgNP8
yuhKoIIE+0VJ5LuI7CtMdMuzjJWA+kDDCLs2blB9ebm9MlO36mALye+OnM5Ufkp32hz2si2KXaeU
OyKy+02PaxLXbhXzhDdcXD++k5CksizdGjk44stJHLDmJBlFqmOIuVDOu+NkGl3P9t53jwm2Ep48
tBHvTvubGxL2Xjszqv5V5dMg4DNvp+tpYdIt2sNjo8zgjOfQDdB1FpRhEXpnancdGG28zQmCibb0
a7SEfWCXuU4Fn2qxCn6UQJ81iLv/inq24LaXWKu4pN/3SHI0wNrKxPw1jCgVtARO8nmUizvcHpOh
1j/4/NIB/V6OlLFW+WI/Lqb5Zwdaom1M5wiownSCKV/OfEzfvO6/REGbqEGV4OIlMBZtZmCm+pcG
wvSiPutdeoGUvEqDflDSAKxaHD+wOT0oSAxSGZo499xwJ7B3KSfSUMjbRUjrIvKWEufmo9hdGKTF
ClWG2g4Ab19txIZO+k71BfyvCqyHFijyMKy8pmtMfyD9Dk5kfFiVNQmWlnA8mfegx9xDOCnTJS9t
PpDmNRapE3hyECinoG0suZTGvk2a/WAsYxPC/tI5L7N5ZcWlK1G82WxQfBWFIRaZ55DZW6Fd5ygm
xKgbJn5Mf5qEkjWJZCf2yW+n8z408dYPUEFmy+a02kpQn7BHUxHX/xdf70sHGcmHi1kfg3FCsxeX
oylFsgQd4x+JCbJKMvs4VZ6sdA65DEHq8goo922/of/C+nfLQARJiaCCzIOkzMFdJtN1aGKOe0GX
Bm4/U/wDYFnjmWCQFobwHmXSegO+MI01iR/2791z9z4wv8N+8X4/BVZ7JbPlTmesNiaD3delzQPl
/3UZtawC/37iVEPQKF7WP/mGH8v1CiAIT4qAm3fk1gjY7hM3IZTndtS4whVhI05nz1qLl5kCCQn+
cfyFgl9k2qtln9s2WdNiGBXcf/Ch7zNVwGd2kZ440zPeB5thT2J+AQzdtyjFqYqbAx+eaYsb/vl4
XqixNdwwJIzBDyI3zh4Lw/96cSbHn1owR0hp+80NDG9JBGN2z8Fyk1Ijx6wGln04g1mAkbPTr8iu
zb3OtT/sadbKUtfOPdo3RWZ0SBxdbNFXM2Su/Fw1y3iv/CKzBs2lYQ9xtXHIVeqciYvDAslPmny4
gJH6cTL2apFAeE4X5ZOkWBubh3qw8tYOjgym1KUFkX9ZcImdrIAlLdqG9Ete6Kw+EmlodZ4QdTMW
tBchmgxDMGEyyC1CfND+7kWL9BSZSoFv5uptWHAzNVnXV8H7xG61IjMIO8dB+EsnXw318jgBRgbu
pxlgOjyLXj2YejNCHWx7ztWkinyqOPSsICHmgRD9Q5f/Ttfeiqbjml7QNiawHxl4PgUKetBrEqJp
Dhwen98aPk6pNop+r6u1bvVx2XyCIotAIUMLwfX1JPMOosSPU0P6L/mpNMT3CMqRsMMwfo0w+U3K
udZJ9GiKxw0RZ/Ns58MSiFsTjeADrFTJpknTY14CbPwXIBQRb7FyeBWVB1UcrPfKuC020qqQ+1z4
SXb5a8MniKuK6CvSnHM3WO++rzZVch2yqNqLNAGxTnd/P2k5Zns6I8sD2YXXej6ShR72xCAVY9TS
m5s5ONi4/VMu/tAiBh2/0aLpnswLDYgQMus8mug4MrN9p+Sqbu7M/s2CIisfE0vVTUkB6uBpZKtc
eKuq06vLHRHapblyT4y4s3faKUChcl9Xy3Hva+4dcBPdQ0TPxe2ruu9hfpJGFri8nIhm3Ei7j0qf
/dFwU412ybbp6GT4+go119Xm3BqIGx26LowflgYTkB5QgRUS44DouBteklcR9z2hrOPEgDPyxgiT
NHqpDBVMjIwjjx13aj7qtIPn6QwaE6erkLaD8AZsgqPslVPsXzdDGvrHlFUlQG0PGsWLLQ/MqEAz
OD6B3ui0XBlWWQpkYx6l/uLF47+BhnMGMC9JBMPGmpjHnRBxFXXHbXE+JRm0KxkEq0UYrAq74HxP
lTe2s2hVu60HVBs2dHStOoOPhIJDOritTmDENTvp6REdco0ihxEY5heufLBW5+n5duMpQQSB36vh
9LLklMwxkE/OIJMYYJ1SG5KWTNUMXZlb1aMfaXdxznKFzijJ0pKaSBPP6N74us5tjMkkZ6LPanAB
PTSBInupBwDd6M+f+S7ltYpFOhMd6KPKlHv09dgKPtPo0oFZy1e7bRR8UjCYx8dQHJyplncBKF5M
ih1YjdORTTcXs7rQ7CISSGq4WM73IQIltWk/YUeLib7Deo+TfTjrgAfMgQIT3tAQI039QkYoTT6m
QkgfVKJhj2IkViS9RC2N5U8m8mNWuAKtXwSGVLkzNEScoM9CkcnovbYq9rDMB7keeECTyipUbMCA
0Yy7+x/BiN9Gp8dT5PE5Uy/E4okYPBmnrbZGE8cTJnwPrbLk74GjkWsUAukArgEYqxecCklhujrt
HgIPEOQ6Sl1sqYYMV4tIpMkrvMvFx3h70gylAK7IL1zyMmxLh3oXDGIIGZ8NUCxzIwU7RS/sZIRQ
+ZH+fuvTrdoe5mDz9w8T+9YmMt+3eA9h0+AOCiM4CpdBSMW2dA3aebVpfR3o6BpGLrC3nrKlp9IW
jnlUGtDig/4jU8YkHyxxS/gSKbuFaO6p+TJzi3uXNl8o+bX1qzkWhD4NsxXf7Mdoxt9yblQZ+KCJ
b9L9HHLEp6Qvhd0UErbUQxoXmrecJ7F4QoFPhvN2Jsa1DLzYFuZ6j5AcPTtYrZSSbDVvZJDAeuH5
gfg/lMKWRrRI/kQj4M0FaDh2pPGnCobD2ATuStKZBZSpp/SW6LI+Xz+uVrxN1+b9GHt6D2DlEXFT
eqA1UORVeXjQ+foC+53waerQjVP7ThHBhH/pWTmzL2+h0g7CNvj4x6KYH8FcdwJpaFVBOiglr4cp
sbPH3V8zCRXOARZfHjW6qn41UiMCbDz15jqXcz9tx4qTB2uAo5SEl0ByGSAhtSrEpWAx7PTBmf4B
zV89NMbBAvkD1j5LXtpwEpaNuBlrkew3Z9iTM5RBoLIo3EV5SHVKDvpuzQHIi/qImvABMQgLi0W8
Nab9GdIXW/nWDXq8C9NVvJax1OZNgW+Jx1CKGwNorDuEFY2w/P3FSSacHLRvwA1HNKFGe0nd4Rc6
d67Qz5O8mSx2NSyohXBMs4wG0Uj/JCvOKgvtOXjCG6bz0EIxHLlsODLs2xWn8W5Aux0xoAexbDZg
5h/CA1CnrvRFWNdCE6gC71oDKz+8Xkq4/kHBvjbPr6HXmsGGtCpSkjiFzadbkQ7BzN+VONzIS4aU
FCZj+N6D0p11w+VR67HeT0ilCyceaIf4bz4Br2H8fV37Ax1+NDLm4jttAegUhoaOm6EgAc93o+sV
Y9NpsBIVkt0J/shTsoyk9DjSo1zNiLzsCoVst9rH4rao12mkh83VvQ1YxbpBq/KUA/JQu1wte+WL
H2KPv0cekj3911x2BpROJibElTFRmWuroQecwaA1b85F8Aq9shjG/FkEBzc1W00JsImj2w1kJ+ee
BAEfHWWHfuoCiU7TkZWNvXDhfHs939OD7NNNaYZ61ULRq3o/uVF0rA4pKE3m9Sm9u9DkJ7AGGVlB
9sfIyIeFgW5FKtHwwIPCndXFo0EYqdI/mdNsgxMqZI6miEUjiGNdYTWrNd9KZNZcdvLuAiYjnywM
x/gaXLqDcMwomQ8akMZQOB49UAvNTsmDWIianv4V9EH0C31/BW36zmnrwFzbA5ZfDVDLftQD31Ur
RvZVkY8yk5kYfUnACKprnA/FolwPQ/x53DUT4pL/4ZoClWJfGXTapGRAW+feBkY4qlFc7WR9s+LT
OBQ5AS8e+/ODTfa3SgQyolyuhM+SGanN4LfX8f3wHEk0D4+OsShsHYxVWYzd15X0jYSckU1Nfw/z
0RpSH4Z7W9a03OcZMpfYgiOcmYZDEz0MdpUTrRBElQUSBaSef44tsr1CLRs+SeNTIy6KR7AcCU+4
QV5htlofMv7dZb939bKihIfBF+sU1ZqAzYXBGtrkDkuWLqL0HBKl57cghhTZBgfPYLqBmQuqqnOV
6c75ybxNKL+X1TlxCjj9tJpZA4ABMjYiZS9No4wu6r3e8KRazAmW5KHtXpEcBUySuYdUC7sJMXUy
6iwx6rc96PRNCUWLteacsjjdMpzg5OY0ySivQVC/f24HXAOltpPd/bJFBERFr9bKX6uuYCulqKhj
jFLPFOb/m7Toh9jPrdcJpXxHcbpBVLlPj2BsZ2vGKDL/f3zL1NJG9JESBrcsPU6BpThPDl0mo55y
SAt+5jK5owpUEAZw2wMI4snoH+QhO1lw5AGHtC0oXkp5ieXNK16GfDSsqscCpbZM95JkYqD24k8d
rCtT1pC36Io8UtwnMTKi7rODF4ve063ICiZSgUdnGUPyG9A/fsU/lewlH54c2piFNCiaur05cDmt
0Zwe8UPazPBypH5DIoUCq+fPU2Xpcu9iHMMP5ASPf4vuSf04lPl7QIiGUatOPe3Q5we5eWl66pf1
vwukRJbkG695UQm2STdKrHvTAGoVR8focO7XZiRCsCTXExPuk6pZ4oA5ddR4cWB1HXjZeM84ss28
j4APrOg500rtkKWBJ9i2Fgcz+eWpsvmcsCqPZ+NLABKAElnc0287S+wxs54sDBQ2Bj1BToFqqTz0
mosFkAPBjQWI8IVXrt8UtmAMKJv0vYOhLbV6nD3cb2h8dqVUZaD8LmUEyv51JG1yITWMQ95bvmjF
252Ughw0MIyOns/A5MTfoVKrXYkHS8yQXsJAOI8MdHUiaGbdcBPyEsq7dJOXfJmd9F9Toc4pvday
WcM241f9+gTiqqO7xf6EP+N/e3bJX8KL23uQeK6u5AAW47d8CDSUTbKkEebp00bcH0H1B1u4SrX5
bmVJTqyjileDGfpZkR0ZY7aCWd9TMlNQxud0HLPr5zCjg7MgJKt6HYM8inc/E4F9Hfjd09IRk7Mv
18ja2fZeQOKBs9tJjZJJ1F94tDrnngAn+QMiauWU1BiYkImXRwJZIB7AyKhZng0BHBGXVNZKSRG3
TFrMdVM8ZijKQPqMWLWi4MPBqvvtEG1Oj2FYC28wgDV1OXe9uesCiLVGVtOzGfu+AlEtrKYiu2x3
g2+m+8ArYZJThZgla1TYs/kEMukPtcr+//7n1+2TJBp8DftswHxPUBYKs0AhEOWg9LWaO/Aed/EE
gER1UBJsMmcORqLJCoisXEhfaiZcxmxHcc/7JaopiexsMWGgqejaW4MB6qzs/gouOPxmDw1F/NT1
HhhpsYiouw4mCxGlSUCXB1k+d9WP8n+93Q2KIszkrrdHJNhU1lIm+eXXVvbmH6JiCnVw95Wgfb/F
TkYhoRhbvJgHaBlWjhCTXppKBsSlR4JmEDvbW3HlI6JCzM3axo87EMLFdvQjOHRlaArOQAfWr4Ug
XzmRkIUbkE2t0RxvLZUKw+Pvl9iYF1ZBzOF3KUTIlI7v36YO3Uzs+Ryr4B5pMRY/te/rtc5Qahz5
xC4KHYt+KKGZiOzMFLtjp0j9KaQjWfhBDbu50lKFnJ4rx2sqXRLzAJnlvUfAQ+ESiOlm+zpe4Wgf
k2P3TkAbxEV60J1k6OeFKICVGxLrLXjEGyuYtzGG5j4BBlzjdbIhIayCVZknRSqyIp5CXOWxQhdj
gr5DrA2jptLXYpcw45gK0CD9tBK7FspMfnpfCP2ObSkbBIUYNWsseMf/5p1b1JrUWU5H1T9mmd6S
1bit+AG+dR6cMDFPaJ4s3VsUFFUBAgduDjReGORn0BUs5RD53ig4ORseJ3wBmWMWGRxc9giT4na1
lVWBqGnTT61qfNYcL5hDwCBfwi3pHId3fXdDAbWaP9P+YzuSohPiSijjouq30xoWdOSnExcMrNIA
KTf1oECyaWwjR+P+NeejTMKbyHOG9M3lYp6C8iiw+GnJ3K7BkOIDmTjfmN/WbI9IoJyidpKwWjlt
vZkclw8SXWlEO2MNFR0L0YePzI6vObS8msOH34CZRsvK1QG6f/CpkCUI1U9zepIcSbhT58SiKRYe
6rfNf276R7RzJObZSkGgyOsgM3As6MNMNPvWemj7HJhXmfSHFe/MmNErBQ63YJ5Hhc/bwdwS09Dr
Z7X2W2koqbphHyaAsmtE7SwDO7qz+IU1TOIoLabF0yzYovIGogTihGXUfEuZYgAGGsyhjQ0olI8p
oYMezmcM+y1divfHEEdcXHSFHaZMNG5WAAE9YCEN/2tEc4HZhpkqdAUtzvKvz2Vcu2MXYm3+ntPq
3GNeV17I0iAPuaBZuLtG7ZR8vXHfdrAU1xrxoKSzno9JWkV9X8aCOggfoyTj5q7vm2U3B3v4pLA3
NuVBo8Ea8Do3JP5CQ/P9hgKjXVEBA0xE2bIyWuH2bd/9lhK+SmMK28T/O6jy5jDIftevNW2K/+sN
ZenBSPjAYfH+i/xJ2RpTaWPiedbOsv6X7pwSCyRruoCI03KmdR5XU+UA/kAp0zPL+DRwQPZnFRas
zExheBftdHmx7+vEbhxtkMs5DR7BjrM66h7697JBP2JoC6khNwVIrm8+oE3gK5dGfNhe0oBY/XoT
N2X32aha0f32Oyx5A7NHKgP661HKzsjNukZ9qGzOiVtenep7D7zEKorqslHpL0Jpc7QZYEe4zl46
n7m7quMRD1qFmTgUO7rpMtyHjJ/vaLkaFbxyUfqM5sxpC7Mh9mWcQpfQhn12HtR4p3cPupWGBmbP
STn8FkJUM2tqydGvGoRUuRd8wUlVwRjs2VQmzDFmp5ZZqtCIc6uRE7tirqdxFkjO5hj1n6lgRaiU
iIAtmrxkqlFEhtrDiAKzF4O9Twmxuc8s/q8Ie8RfArayEA3G1JT0NJe/jcAMc47PI1Pa90JbV6mT
2EzvgFdTUp5D2/Qo7glhrWrcTYeBneC6hj4gsVDnIdPfGmhIdYD1gGxIEVM9n83xgy+8co04vMun
c7dGRItgN1DdxWVnmZBVfZtUKFtqp0AxnFcqIMfOPoZK3bnAaj0dWNwF5/8s+dxFxM5saq5iCkxs
sTDGOEPyqcGS4AG7XkAxonVFshKitzxMtoh8NHJOm7O2X9qYPhVtUxKGH5SzHiQkqEUZZxdaSeHV
AHZOmVgTXroMQRQW5QZJIV+TuL50X19I/pp1W7iaWEEUjZ9W2F+RfQyQEHHIyK8lHzmKQoDE2qsZ
f4fjZ4R69YDimqpUbRiyhr3f1Pa7pBqHfmon1TFoFkuYxyy4Z4bxP+FrShfgkERNSRCBgRYv+/EL
YvHsfk/xqs5MkWTrbcbOUJnYuxqzTh7ZVFPtBIpc+r9WrJHuAod0rga/60VSvUwLZoTi4sA3Uz/v
seRJUImCftHgBsXAi9P5fJ5/8ywyWgEngd6nC1umE0WP62zUkE9uCNago6LImORocFGnTIu6z8uo
LRL346mRh3kt5985rLId48sJ0LCxM5KYyr55uJYa3PuKWa7Pc10U/qWm+k4/75Iy3hoJkvMiVFzU
aGLHwed95lliit6RGxBBvvnWVo6GLe+011dTm0TVrU35YPLJokX7EGicPAhYNYBHgcnzLkrp88CI
NHJA+hhPFOhFf/Z47yU2ryJb2EcNHNTZ1LCFi5uoAqaclCF2NHEvwlf/W/k4tJOaLOmIsS6ZkTsx
b+oGj6HvWNigynTh1IEkm8g6t9OAGSEoa1fzRL+5XP6hvpwm3KlEpE+Rlji1ifnKve7kDESoDv1M
OqTey6d9OJ7J2Itcaxo0Q3tI6eZYpj7vU6ysX+1eY8c9ZrTI1uN98wOnVGpGmo+eb4li1iFvdQ2T
UqTnWlNOfJ2Zcex61DMW8NbtjB0Wi+WnKbn9FGr+6e30YNnkSTn7gnadAhresXxnjgD6jEUgY5X9
JPZ0fiuWdEJxr+4jsUh42FiMXuRMQEdh26uywgm3ckwaC07Ock+d3xIlrSvxJQr+BSikvjo8EClg
5qLO+w7uaP4FJrEEGdbH87WprISEjOtBQ3CxvtfcUyMHxMpD8SIoZmdYs2OEtsMikIBPBUOdJ+lm
aJ7QptZ4iEJCeUoZCUq0WbEKZJd9ZSM3phZ2TdlUhZqDB3ZArhfq91O2ucug9Lv4heqxtp0L0YrM
HqTAbmZi8Xp0WDit19odACMmGldyRQBiIu8/byu/nsjgv0gvcX2vstay3rh+U0+1U986gYBzG4fo
WGcw3nnXI0QV6UmJlFL0sSPEPqEFpJeqPHqlXEixarI9hwU+UZQxjUwaO0zGCDosi/K7Ai7xqey8
6nPlc1PpVXdoqL7/ncDngR25Non/br5kxvkZ3R5Mb6nsvmIN47d2gd0ioYOuTs+Xf2wPQPD4hV47
/R0klX1S+DzpkgoZxF/SVgcLwhazwAPoyldrkmtdWs/HRcVSosEYn6i2Uudokj5hiQu/cvHTASf9
nz+KofARMrEJjzfTDca55lyoNooF58geMXuRaUpowufBjXabPlU+Xp6SoGPcMFVa4We0ngGvAQvS
xbN1h98tkZ07GthLN+LqtG8cxwLi8oHbAueuiLLKxYRCJ6GN0hQvbkBhyPfTVTAYbh9/wmWzdobp
kyKLshz71w4b+EsDSbBz62XNRXEKm6W/MBzUqwtdEGdbKmWHQD9WejlIa1Yal7hTGqxOHG/HvaoQ
6nE9II4BOSIORMv+f/7zwaO2ejoPaHCstAvmU+TrVU6wxcQq4r19ubu/0EgBKcBge0xhN8KirhGx
4xJhuLpm+LFsbFhL7MThYCo5MuAFFTiTlRT87995009A/30TyAzFRe+1IR61rHeY9W616COE0AU9
mNaMsjhxqKNd7Q+yTSMTU2FvErGv9Uupx0rHkbk6nKwh4bFZD4ueoQQShbyU9cgZ9V4JgwxplZ0C
a6gh3ZicapFSFqgxjjNjSDHlkjRH7KS0W6GGE0BRbpD4FdkQT5QZ8tbKLMHLUCJibeHel5im9FJL
aSwX96q3Ls+WqQquSSK3MAu4Htxx3xVfvNlGLuNPLwp+7OTngKoa20CkzyB1UgNYqGr63RvR8nHV
TCMi/tsgusyjcH08XdSSGW14/rlJGTRYuhm+64UTnLZImevuQsgTJ+Rbo7u428sHuLBMqlxgA87g
ts8zlptGnLU2J1WIi+iM8C5ZuDUZd7HJm/mXSVyrOhNOWqQBXbvv3MbtgbaQiJERMQQp9hz+YkgL
et96es/womzvxHN1JkzJodqckaiVBwqLtGFjkcUaACRSePVPE24+sFIUcAbN4M/AOn8wlerY92fn
XENnJTpHlVrDCKzBmN5PnlPCLBVdrvy6rKY3o/1cdibDgtkYXTOo4bk=
`protect end_protected
