--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
AC6Ndf/c7HSKDAPymKEVBlv7SIzWeeeJPG8QVWb/c5evdWQONbJ9ifmGZFOlzV4tR/2ggUef7RR+
NnQvTKsBB/F5ceIsvK6PGNu+M0lTnE5ScXe+r29CyraGSE4pS686ZBJdvo9F9Ktn8jGLzOPBj/wX
bioeoe3xO2tACIcvFji9Hs2hI6iGDPSOMgQ0nFxVfB5VLsbx3DzCtFZStaab+OfuooUL1tf0J+lT
/vPXp24oNQhHhBnCE/4fWtEEpKFZK8V4CWXFub1NLyy5Smt/nsFupKTx4mroPQZVLZtNH4AxJ/0m
MyjnTN5VKQtwFsPqXhS/McUWPRvi4HbtTVIu3A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="OYEVr0mc1zhm1SAH/xCsdeQ5PTPAV3hL7F/USzB9psw="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
dFrV2KEg3Racl42QG8iTKfCWB+nBROo2Oc2wdOs2hLsIv27m8zz+kRQTPcZSk2OezRiV+T65NR06
2Ll76iWVm+Dwis7MAuNeVx8YTPoGFv7AkFEAp42pP/rTik65T2T0cpMPiPI48Nme1cT7IBNuedbX
/6wuQ6UFhLKFEK563IGi4Mq802jaGdr8aEyM+jw6TZTU58XLEofOr3CL9rNiaTMdLryMCaULobVn
ru4Hi1Vnh98K1fOZnlmv3XiSNZaK0d2b9Z+yCu5opS/lC71lmKJU+SlJJvFtOlj1ik2XMn+QetEq
tkpTaegJcvRJ3Kc26RZsy5K7wn8JIMDA+yo4zw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="BavAoGNK7RN17RjOTdJ5YtkqZeRyYELIpkFRYMGL1CM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6608)
`protect data_block
zzvvzGIZFJ7l/ByWs8Rk3SLwX1vZGllG48bN4MzG/77xy6mYlm67R85YIJAGg5YN7O+s5oajwYkI
bNLn0yFqkDySNS5A1R9YJxIbsGmwZ3wfe3o9sEHnb8BXTHXMQHsP6f7/ScRDRWEQlZpWU+smJpbV
infoigeH6wZC8wC8c8UrpxyC5kpJ2NV6/4X7dGUnmSdt6ZeQ4P4TUwTDaNwVVN72ZKKgEkXlfjhe
XJ5Z7xJQ0vvDrpRrV280cqhEOy0xWXSU3tcSrQkWHjREp8Axy1nLfLLlPK15v/AA6WO6LEfUYBwM
BW9QFDchJBpvJf3ClpbYSw1KnfkIn6P5oAs88QkgDUMAA7TKasnvBcsvU1wpo7l5/34PvOM9a4rV
cq5F3od0ptw4dce5ikO6jqbEhgM0OKpad4bMccKY+mrPJdCjVudNvsJRzAl2wZux2q9IxytQ60JV
c1J7DslAxW5Pp2eWxwazJRGn/shYgmmHUs1wR8rwPOJQhbN3CFa9YdaQuShv+Hh9oPxe9KxB+h6+
jMvv/PX5U2IqRaP9CVxND+J51ftfoP7ojf0oJrGZyAJLw1cJgNIXP36h8CHX3ZsAE+ndzwCvgQ9h
mCT4A+DbG9FPz0xeLsvDhz2OUYTDtl0+o394ceBHBeLpoNQ7QaPUMUS6dvptonY5TRekxFdbOXnr
s0+RbB7GWrYSd7V0nDKBcsW7fyEo2xCp5UyQVUtJvFM+1KMsmivrqqCPJHj5/3zlhTIMp6+YF81F
R4GcxJVM5PN5gaRDXgIxIOnNfh9fLKNiUZhlvkan+1Lj1rakvz/gawRFPfbNUUbgBg23iO2mYwef
8ej7SQ0sdCjIMrA4alC+lPoLSt7MfkbhQdzS9udhdBgJbrkqBvGHbnMkX6ksUnvEiUG19ABlsa2y
pMmCoJG5f/cwojPMq2CDXN0C/ZNb8TGcEu1xQsLs8h+dClvz7ymHNJUM9GROiNrf0xWB6uMcGZVu
8jVMI9P0mbNacGCem5KNNR5SkRKkYiEwn12OoUEHCtHS02uUXwjFV9exfYI7URdtmSVEAiwzL7sK
B3SCcgKrS/nJaXNnRbPuDzvSjlRjKEFoPVupjjKlThSxRPkiqrj/FDCWI0tvmUx6YILLfnX3tRoO
kZbQaF0cM8k4OcGmjyxYjZFJd64TDeENdNcJC/HK/8YdvRk7VkbI38k+3V+BAliq9MCXB2lqohHA
fr451K9GyCy9TPTOspd2nhc0/Q/8TnQRAzyEA8Fd5bIyHpLgRFfZUAFybJMBICBAHhuRo8DOt/tD
bQvycqLHFgeqBRx4gLbYzy1j8AFGiRyuDc86Hw3ud5f3muSTGSG6Rx++UQcz8pXQ9l21KSk0Pipa
6lP4/cCKv/CyV1h2F8porxTeZahk0FFFPUqm/m5ewQ3nCz18GFvKuJ2pGvb3RxYNyHN55WRFY+Dc
tp1iR5PZKd4YQCy8V3JgNhA+vvma9uVibD5LI06LbyBaEB3jQbmPxEW8nfN7vJhq5OU15vqQQETc
4k/F9NnaX2Aett2ldIJo32WiIX+1//zvqeuLJedmQtLkftIL0nSo98WqwA1+3DdcuqYxFXGmpeMu
4Iqs0yWKXgohWRKUKfLNAqlLNKn+unlNKaDh9x10Zh7VdnIEEmnziA+QLT/D2Ir6OCyFTV5ZxVEK
Gjn1hDI25WKexV979mwkgVYHSzh72Od2ihVm1dkRwWceh3bmbVUcD9IneO4+3P/+qcL1MGEtX7H5
58ElOxT2Mi85eArVCLNRQd5Od1gxLIeC8WUgKB05+ASTAuMTgLG/qEDzHaqIa0aB7Er37XlBwI47
01hW5TMbstuQUJPm0tAtGQWbM6/uhhA+qGNs7mcW4rd33UFXZ8l0lip8fxyXT+8YHGsoy9IOp4lM
oUZJZ5sqdLrez+r+xLQN889ns8/pd6WACP0ZS3Hb04Q8dlHWVC+scKXrLqXbS/ucQUw2ZkFSrfG/
Zxo8Z+E0VLHHkmfnTCYcBl+ZtByFuRiCs4olpqGzsfyf8mh1Adme6v9NJQLlGWbcC4rz72tU4IPx
D87qpifWSwyesnTpR+uwZ1zODDJ9eNS4FzXSUE51ZRr/JzZ8wGhcNwN06MthjuSgmANk6cXQ1Wha
DlZ4WInVc41kfwXvhbF4lpf13+zalYfzsSnuhjfIsT+Gkw0lKL5+vrg2RzNuIGwOGatmkbTaQZAG
ZJK1h+HtM/vq712cCuUtvR6r/JsMVFVFxQGNBy6/9FuIGLG2XCnrNmy7vQD7yhjH+A6wyOyHNydK
YlfFvnZ37eIKTkvOAOoKYkrGwL4Dk73ggU3mzLDEeSFz5dhsSJaUXbjnkH5M6dYyemQANxajiR4M
ApsNmH4xWWHaE+NjQaWVIDTHKNfK2Pheo4pNUtm3tRWHCYlt/Zvvmn/Y79T2h0FlXWO8rVhNmcm/
acL3CEbNUfmVaRe4qDZrLp6T4+4BzjGAqSRWyNfO3pSH0xfUo5KbAX7roNBOtzE0bNYC57XICU5F
+RaLXGoyydC0aS4RPe7QrOlLFlkiUNh8t1+C4xp8gl/wxe3cZ1pnA8jP2TX+iseSluW4+jReJ4A8
+5royzEHqkRo/t/oDcLdPvrC2I8Fs6Y/6nT7ztzT7UvJFVpP23mu73o5hsCL9F370n+kO8Yaekhv
WoQThauIcIbOe1lfBcDq91MPZm8/cK0DZi4qXItEDOKStNIt3XyDwO0J0QwnpW7tcwd1isC/vAwc
GVvMMGECpuoh2jtXpbIKVrxpGUaeze7/sxHWuP53jZ5I/U4fp1RZQso5vY4P/Xu7rFiqj8XnSzuk
rDNsgK76HSXsNHpUB/xcvQEBwtz+ks5TUJollY/bGd18n1fmW5SOyZB006PLWSkePj1Bhc7Db2Rf
VvhzSSOJkMHkWn5xyNIVAN9HgN2qXpHJvCdy6QHSCftopdBPNxyE82E003XvG7Z1U4Xa1KiP4Hkr
heur+rRo9U9Uk/bXwdhiZZfX0nn8jOnlJQvJG5SzrMSergcUX74zOuT/BmLKcW6EoVmo4kiEJNa3
S3a/ybt9l8dnkil7emSYQ8Ho/vyCOpBKblG1QWgrqMpeygPKhNU85HyWeCetocESM4jwRgrWvoIh
4Ee9ih+nwHmn9Xji8/GMkl67Fmv8DN5AuKJeQtNYInyr7OS/5zDbHj8DsuIUfTFpPkIyYqFX3ts1
zKV5HV+tO64N0HN7w7WRyWjbrPrWBOe8FXobIDInIQF4zKsUpiESxZPUG21njtfkENaYhHfbFo7M
n4NveKPbEDLTDg/D7GUAh1+7UHDvha5mVuw4pcfu+heUOvOelfw3GWMxmtJ9E3DhTiaspEkuipNL
xnZ/UfUUxKCFWXAWur4pk8UAkcMbQ9E5GHTWD+rpwxCQGwn1ddpmnDhLywEVdk87OQJCWaJKk5Xc
ahbGDnau7dxIQj20yXeU5Z8URreysPagQinuUs3JDP8jY1cP51KHoTU48NVz6r2jQk/Hvu0jDin7
zZSrTwkwO0uCS5BTB/cFaxhu0fEvxTzyd0u89qyBPyi9rOqVuEqdKkQ34lVuoZR9BX7vpuOJ9yrP
nyxRRplM/jCNdeX4Om30+kPa1eemvYwgCyN+Qrxy9Lz5XYGxQ8uh/cGeW7VJ9GCrd8uI1KUZy4wh
yjt9/XExVuNeTd8Z4lflEZdPSpXcMCGvZCBuUMuXRaCEf+DXTrKyZYlAmqPrp8a3Szzf9biRyj/d
HYe+DuxlqtBTpU3U/Sfc0jXeCofoWRXaI34GcATgEyOu1EpSAxvbRg5WoiePN3Afxnf2Tmj6vclq
tTw+4gNUFbPm7CgH6q9rIa5EDB1MKP6K2wKxMiLCcSqHYpnGqt/0PsnrrHopW7rmt+OxfdU23YQe
0aLMG/Xuue05XWpsiB1OE5gtlkTMWxH+GJ5lebTZxyIILrxG4UUCM6bOz6zsMs9cLUVtDcgMqd6W
FIadD4gKxjNugBjkkbZZS6BFe0+KAtRDJPyiyNGDcvbEH6MgkKWbA769j4uj21P1XGOJHfMwuyIB
q6mg5p4OQvofH6QAN7EHR8Fm3RC/ADxbSaZaYBNEX2XmIRROrxezZEybU9mQKMbrylW6nYhuV0Tp
ks8WMqk4/wylZuIqg6iOppTBKhfkfvI3ba6WrmJ7kNkf29Hzw6dYdoijIdlqbhtziJRmST1czg2B
9y3c8meVGX8SCnXEFv5xwelukFV4YBUdQHCvHRbfvBtg2vdTPk7vEbq+mpA2TZqc55sZ3/HJD3PY
5qsu9nX8SEDfVMm9o3RAorLvgtfp/58hLLuj+C1ZCtUwptoVWiFcE4YU0IvQgb0OaYDuHHpUsjcy
ooTuGVQthA8oCPF4xdydbptpAvUpz/XsWobQ95CFRPCFZzdrYs6ZlB5r/c5D6G59dMNjldS7rDE9
eHcQBfFAaf37UBgN6igGMCKFzVtqAoqRo98WTSuUEyRo9aulEw379JB9ERAFO7J1r/Jv6V5YX2AS
6ZrF0/b97xFCjUZkkQJPupZFAF21aQOhWhumVChj5Bsc/ndWf+4v/+iWDrVnTekPsAi9mjLARnCS
NC4Xr3LeZC8fqxKroPHWTw4nPGRos4Hgusi12p1bcJTNt9PKRSJleFGnoBxfMcJh8FDaHeW0VdVC
7JBEgqVkRw4w/0JkoMKGL4/WMzh3otG6vvdo+Zbz/2/75iD0EgIpMV1UqI/Fpewo39RY8DdpoJEk
fBaLLXFg05/C1VOVtNGVFOjI0D/fOCOLgwC9LW73HxZSzUMYRK3fIbPrbp/DM5ETSKkMToOPT1G2
6JoUaF81SBcCuBkOV0oZd0jxzXiLfBX7shLTWByofr7540JbqRFUDJUYAJGyR+6yz68S0KbrqVUl
kLJWALmvwL755AB7DAmK/Fb1oFM54S7fhZGAivvIqdyoJ3sfcvGHoIMaESW7h4as6CBT9MDPcMgC
qxwTT1F7XlY8RzjePV7Gy/y8L+YJkQDmT2R5CgQOzH9i4MO8mHQvR76vy2Mg3JmE7BUUCPgEAF26
VJ7o51NLzKWDXO42G1rilFcaCeIKXdWkKiRL6qYtXMXpigEuHO3PFxHJvhfRHFLGgZty19v3hnL+
ReNoHPydvMPH3aZi7DowTUjBVz7GTbsPgZm02FNp92gsE9avDOZVYCiz8uiGUlKM/pAyIZucexTe
rjCWRkB/JTOh9uQzq11Xjy/FqUuLxgvg+k3GvEIGn/CVWdP4a0tZTIpJwubFqatu9cOUcUzjxIbk
zGWFzdvY+hAPgTl2L6+xag2Rb3V+IOr5hdx4EVkeyCxWwXKtuti1AN1TpBT6OmANbzH3LH1O4oX2
Yj4J1pV5VDfbWJbA1APBnjR0LgEgIoqwcK5cCvgKgtrWoQJdDFqETzpCoDV2wg7sZvEm26ZbU0pu
f47ACMnQ3wYQPqmmuQjpDD/TrSexXQsHnpEYanZGht+cWGvSSucvA1f1IjXt93L76ZajqpCWdRYw
MkYhn7kIlMKj6cT1po+vq4VAnfaZMRthLLSvdm66ClgRCWWO2GdeVZ83tleAbE1Zg6TGBsVODC9f
axRXl4Y4rNKCne7FkBG+Zz7H16tvtpnvm+Xp8mvFtzCqG2y+H+EQUT7q9NlSeQT6i0DM05+li4wD
b2ugJumoGgCYW03i4JQkh5TCLgp9eVDm6odGiHi1l0dUsiPMECxMLrbnPNz+Blbfwr7U/XAjUJVA
g4enFzBXOy5r9Za7RBXO5r7etqC715YxH7aBtsoX378fW8HhGxLtYHjTyFKKlcYCyolL/JHp157d
KTmSFXGvNY25zq1FxkY2YgRs3CK3I8IjoXzmM1mckyRqU9GrctrBhnKizeiiil7unbo54+PIlF/B
qINmNUcqmx0hZisHWL7+FdL49nKpc3zxr2L800SI/UmnRT2JVfYM7M6cUbFj932B/sgOLCQbDQUL
3xbQTVm/gYO7kLj3SrvC1DJ87Kuwr42gKq9Oef5r229Od6xS72b77Rg7PplAUTZSCHGtaRSftR0o
fzkRQNHNBy4Vf3IQOwJ7QxhqnW6Lek3bgFOTRWFx/8JUCv3DyOQ6PzZdcd2NBrB175YHS2CKBiDH
gnjuvVDjOgu0h/+AFye3DqIHt9Fm+sQZNeVEFgDc5SUUE6XcRdXXTF+KBx+5Yl3ylaJl7YdQU3us
Ry8yAjFVSO4qhZojiC9J9DFIg97FTH5L0Ha4W/3jdJUF+fO85heWdQIMr50aCZ9yBswzOC0uCFtH
UZbl3VR2zWbbIuEx17GLlzmZzpoaufv7Qg8G8VLPbVrPZuUK0hVIVI4CL/LuKyObNXaFNaBBwK97
q/R0sMlIsHVfMpxr8MZH6h/mUuqURcYTI3ubZwoYxy6NXQ0Ra6ym8BmC+qRjc2b+2rF+b095zYL+
r29bT/KVYREUQIE22sdfErl2fFrNvT1oqNoT0h1YXtKB7r503TfCzS1XVxNOsOHRQYG1IyUyctiG
Ld7FabtJ5z+fPaa4ktYvvs95gFGWTsEvTzSqhfbUtrjU+wnM2Z5gCTwNpMOPNtPfFgxXUDTZpebI
Z54YXN/uOGCEKF3qOAswe63Ibcg1KLb81HPIQst78Xbj64AjLwTUFffY1yzJO0LqGeoaI+baUspw
qc6LZeWxzTKCkpu5CrWilxerw7XWISF2+tjQrmGvCufQhj69f2XLPFldhpdfkztGYtAv7SnZb/LD
PG2kUvvpxolpglGxIYKkZJAQIrnj/FdpImQygaQb8pE9jtIDk0DxWVwWyphJSNbD6MOBZRoXZo3d
em+hphnK93fIUgLE20foT8r9CnqwiLR8lTjh+yusZBfOUTEBR+a9XQtXZa1/Angn70D8hfFRSgQp
FKEuCulQnJs0InmbASa1w59y+KxXQKJg3xwpqLtrKOwwwni8tEQimNOX8a85ZCvCDRyYJt5Rxag/
diaP7NEODNNma6RR/ktg+prlbhbo9c0FQT8jHARbXrqyNaNEOsY0+mh/tRel9zIkFj40hDbuRmww
ccySqNDJY9ptZXsB4wMbGjatgMERKGJM4rXb58KdV3tG7vkcsF4rvwBRooQhKE6QoyIpGO1sv8pr
znBp2NW6u/9YnWunzwYzwTIGGkfBoKL0PEgNBFnkSemMcucd+Ks6nnBdw1ptBZ4z8++wJxqdQHvX
lsEWf2SYbtccLoXKe2ze0AEIo87mSYKsiW4zBzHUYD6Sp4GkJ9DWafY7hfheJMJTMJLaPI2h6gUb
V853JqRSHzQ05N213f2z1YMuEmjM8Zw6FXlA2O2v4tAqI6BU01/INthKssBnxYGZiUspyaC+Jn2m
UKpbnaYESAtWIU6Jrcyu8qv7TrJTIkldCPUoRugkA0EOsOP/UPLjGg/5Kv1RoQObF496o8wQjIWc
yqTwFHbjIgGhoHG8iCh6uyttR8D8KFF3CIDW4f783eROm3LaqUUqgwc94xGu0WMWqpQKVmn2y+xx
JFulKZV1VlcZIKF2U/BfDtaZVw96OfQiKB09pjJ2WPTYzT2AzoEAxdxZFCo6VPq8UUzCOKGYy5CL
6JLoM4/SnTok1rQyVfq4E1YzUl2ROS9KrdVJwckhrEEYcRibEvUdjUYOqxiKRV/adZSLpnIW9zQz
g7OdlvMcir+7c2CwkvyrKrj+COtkXgZI7yoM7FHbiuM7iPFhUFpiLVvY+T4oqF07t0R7T2vOQq/d
h0GxdtR8GGwBXPeaurj/EHL/Gjt/iK3bz929l/LUW9lqIVdIO74EM6eiQhrqwzGMQ7YdFvFMHaVc
WE5CbG7ibaJ/KVSHLDJ/fWAVjO+huLuZJdkZtJewulzs/urKOmprRdol1kgc7WTu+SwCCy1oKv2w
XJ0a62fD8ldEB6UN+RfK4/JKrsqf1+aM23OeBJblG1QHFhYg+2qCG3DStO8NPsRYAECMse8y0NAc
IamnCiXV75FI7F7X4pXlbUJ6oA6KP0aP8Z73D7di+avRV6Km4avMI2tNTMFTeEgwb16SL1TY3/n+
kXIwF5bwPTz1ytfNzHK/EerleMY4vAj65/3UOnxSUGY8+vxr1K7q+iqs0QKVGuY2bDFd0y66X6Yy
AIONFznZ1CBl3I+2LD4lwGE2rC9rWPwX3twssHYFaB5dxaDMaWyGmi/nxfaRBAM9CUJvLULZ1MRJ
hXze0cjbY5uBXv6StTkTexxV1GWl+0HbfXtkxVrgjSEw0V1vN1jKjvoAVloHA0C1/52uWOp9A+Zq
D2Z0dB48oNh5ozmRqBTMoASsG0DSJC5ahNjlBqGJzHYwWM3n6DZdkoCQdjaQaC6ExeKTc03i9eG9
05FzKLGtLHkBxG5M0gba33HGKxqosUuP5NJxPz7WYpRkaZe+3xXIARu2mfPL4DOtZ+kmw+p3dxJK
rQ6n9W0AfoCTn6f+jhZtPmuAU/9dJ1miyqWNrFj82nwcML/8kFHSyVkMuX8iQI5gH80OKDnojluO
FKVKVtq0Gyec7ag2lRdVIv1cpcZgHtZfY1NrCuv1TBNNCfMIbr5VyaHeJNKvDy8SOJeY32cIIHA8
w+gaquu1KgDHkEJ1QTcKdW7GOorLX7ZCGGgYHLLp1h9NO7U9lKSIbl+PGXEBK+5VS2WiEd8siIDL
WYISFYtReNzbUPjCDB3FpkMjHPq5RRtIAqXwsFFt6Qoa+HDQ0ChWFMaOorBY4fC6ob964FVuXV76
pXpv6z37e7m50oraQkxTq93VXoMLGyBac+nepuyJYfwRZqKxUVhp006bBc6pmaLrJEu//YGXwvR2
Yj2PJC2EaY61iI73dHpbBAiUARptcMeSmityU6EK3VAFYmNrBTeWlksmMle+bzFGnCvuXRg=
`protect end_protected
