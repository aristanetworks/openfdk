--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
KiRb7n7F1eMJYRjMaesIfnykfZ+CfB8rKUXm2G2HBGHe3PY96OGhCM08sFZXuUrO9LTSVViOTw0a
Dn9YVYD7sH7OXXz3dkVRACpyX3csrRv05NUepn8gmNFwLAzs9xqah3mcKVDOgR/jwSPTVCvGYz76
lyQ0H9W9zFnJgkndVOfz34rsb3pIItVXYbScH7/7hAOz3mI7T2cZs1RpD06Cbd4OAXMQmQdwY8rS
SOyLJFUoyTmDVilIXsFVUE/HVvfZQiQI2Sr6+48AsgJqX0LpP1kjQ7olITTMh5cwyQu07unMgFD5
N2hpGBye76dzuU00wpB9t2c1fPbJH0W5rs7S2A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="XGlJdMOVzOk96jt9/NfvvuPx/wfM2mbzCulvP4dCn3Y="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
lvIxKqPNqj3NK0iNY+g299Z9vj+pkRVBiVYjfFLTJJydHN28LBCN3FVGWoLAZOELmrFHqTtY9Tgo
trjFWqyIqd3/9P36Ep8GfK6ncbiXI14c0Nlooz+Q+WCdbDL2tPVaGuqt5bV2DRlbz7HWwQ15wrVQ
kFx7lfhcdXTRDGc6LkZXq13cO5Qxq/LGWZ34mnqCfh2zyjZpj90ByEZf5KsEzL4Tz3A8BjQQjjUA
+5izJZ5FZtziESa87K4sOjU18bfUXQ4mzZ8SdsJK5Fm/ZxrHPvS7GctTrE4oB5pg2x87UFdH+OcU
rfyNBJcq+9dl8G1QaztolEfvrLY4XcphbSpmng==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="2UuJ0HowMNjTDVOqTMOJkeesrr2o06Auupljmt7i8BI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20192)
`protect data_block
DR/Eag0nXHpC5DtPUquT+mdPC2DzbftKAErAOnIw5a+5BU2oeu6lHbKgDN04vtDcclIsRn2yrVlX
AdaaZIONmq18GQ3aEttmW7JVgRM5WdQVjRuNvJCOh/QwFhFC3qlLnlCF8FrNeygRtwH8ke25jADv
vR/BQ1Pp6HzAVsbkTtIeeSrgnMg1cfDDl9SLxhpM5wjUdjxB2ad3eBfhwxWpeFs4AvSplz9Tn+QY
tKZUbIhtlPIa2jiP6gUX3VsYTSKXcSRHYCczig6FALYqP1I8I/c0m42ZdqNNaXz+596Yhn9agpQJ
pyMI0GIhjGSs9I+cRchtZTaZ8EMhG71YwdxlZrHoe4A0Btu5+FBCyCwbF/sOzhbj1RDB0Angm5Zt
V+CqpP8v1BdRakwNXdoip/TQzeq1UPCbzeumkbh3Al6rbKQwsC/IvBGYnedVc14KpTWC/g0nAUww
fhv0yYR4PWO8eo8Bkz/b/ow2I9Yn5c+LIv7kfJFLymWdmp6meiu1TbNk0ZjSuu93f+ZyFgzXX27Q
kAFWbw8PONzUWGFSygYe1SxpCRmfo7KeuW0wtVTzWPe++YdY6ETj1RepAPcP1ihXx49uFqPGnZh9
xtJ9HT9ARTjSZ8TeX2NUo04K+97/9M/+WRiDLNvN1GMm3ena/qmHmh/ECxj3m6P54AXb/DiEFOMi
ggOqId+8MNoEogcwmHKDo0Oy7VLJBoZooQUZDfVmQNSa6eDN1xTSqsDF1Kq4AMokvR4btvJ/LvRm
Vh7I/853CK3Ioq/RgyjsVcXHL3iUx0359c/IDQbuqHZqn/IEd2NHeADfRTIRenMcT0beAqc+9pb2
mfcsMp39Vj8Z8Yih19pQsDOV2KIv5kifUaD5QgrtkuRIcsfdfof+ebH+DtAVoF+HXxxBR/w4cYx8
VCuaPaVaWfM13Ffj7n/+bLyNppf2OMQ+nbLt/ATNGfDebQ56p7k0t4YKUw5y2H3LGrpu8Y8Rswln
IVvktbK5qIQesPIMxxcZeKv6GlW7qNhX9hI4RFzMcoX8MDvmcdodr3hIgxiUw5lCt1mls36FW8H7
i2XbArVG80uZEmMLuXg4JroaTgC385BWFyCDCo4z+m+8G6fMq0Ul8UnN4MJq6ZMSzBFJCfD4JFzJ
N2yiUvCW9uZs7yLNEm3yeHI+Fvb+or0pQfdng9U/y2y7HxW0IagVnZjOvLwMtccxCHj9vN28nx3M
zB0AjwrdIXoii4xdi+8OafzFF42s1nIFwPB8ikQ4LgfjJQzHEYRkHisO2DlPv21Nn11FSkJ0Hg71
UID6huUfjuZ1MUPnWd5SwfaN0tnFiBHOu1KpPMcL2r0h+QcuJPdV32tCpTtHlK1kjhtZrLiU3ZaZ
LdaULjNKe63c9qOBF+V+2Vxo2ck34vtiUfAgSt0WHDvE+w9w4jDfJVGcoDoy6txlYv+aRuoQL8i1
Ls53F8vnyDt9c0Oa5DPMxOqyMOblDWvnmefDDFCkp6OH08PNITcPIN1PYyW/HRQ3JaO/D7CJQiOW
G5X3V5i4qQ3HrdhtlEEzoQkmX7rf5nCwPjYN6xRPriDVc6JXROZ7xO89iM1t5bD3Ej9Brud3WmMG
xBTSVVJTOxxdS/ae7G+JhLTQ4pnYQNMfT1oZ8i28uFGUI7A+81n9NJ1qU+D4/+5id3HwqAYKCgCs
t0jQ6aiyQn1OqmQaprOe6yl0IBxMkvY4oJ/0M1Q8mY2WIPfusLTEGrG6GMgRa/QWjSe3x7W0hkHW
tvnvtYmQzhdShpf6DBR222pF22VkcLZoIvbhj266zcvUluQH6JC9RciwWoJvEt0aoEmP7EtL/8y3
0Uf8oE8pbg18toeHYS+Opol0OpYR3J3BTjBnbqO1wF/mA4WOfxL8iMX2I8uBYbKVhruAMPQ426Tp
0hgTzvjHBCnTSjfG9miWtEiI47Ni5tTEFv6abt2jgsR2fJIJFe4pmfFIn0UKXnQUEP0nDAMqOL/Q
P+dmDjno0/AlsY/CajTFSc7DRgKh8j1P2da8DEBlynwPhcHlLsTIdkJYcCbtqkT+XeI/mJwsaTLT
xon8L1BfC8hokK0D3j1uo3V0BYeRtBTbeBFX7Gh5tnwK13DCST1WRN90cGoYuNp7ahyADbF3j9Eb
oAUjsraW8JxG2EeUhoHNqNzRKbBhNsah4GNCHF/BSUwX+zi5gA6u+RSR2Nb1Y1uNgOpfvCFpfdtC
16DDXAMqWa/GORNaJya1v4KAFuTQJ70cQExq5bK3K5czJ2vmF1p97YA6e+86NTOihRNUmxEXSkfv
3t2sG9DTwFsh8SGraBS+u6hLrgetZPYBTyt/OyWBkCPMxuG881ss33q/QSLRvkVTc0wGpHsUeMmn
djUNKesUwPOumcflCHhj8cAV3aba7XPABrwjHG5zSb1fII9piWbzbAEH41OeBVgeUoXmjzZvABNJ
MgsbkgOuHhM3ljCTn0WA6knspY2J3e/40wZmE2+sWzA+Rx6fFl+epZyVQakD3LLdZQQwu6RBtxkT
UxIqxyiNhX4ug4bI94Ya/elcFk5/CX1ENdu/N0ZzDjQpwKJ7G7K+dkDiuf+Oa19h/zmWwJpBqL6I
feOlsNkZ5tDNC76hRobBCDrOXdAkGOVkgEevdNMeOEpVEHu8zUJ0ozh9OQoCVM36OI7sfjnYHoLk
qDqCntbQ53aYcCPG4VqXluizNRxkEJw3vd2aLgTaLmZ8dIY1iHHALAX3ntYSETk8jQiVeW5YGxXZ
19uDeo2UL0MXgi+fZL5Dyat8nzfh+01WKKGnk/5cyhHosYO2GC14zm+ajLdiz1F3bvyfMpK9rCvl
EnK8OUF5fjGDHHeqwfKvsk1tH2zjOC2g6VNPK83QrjI9ki500GNO90sit1E53Yb3mPW4sLyRWlT6
B5LUWFgs71z0rIVY40xr091q2wEZpc2V2xinnJit7R/xmnYy5G/y9DKBA2yMZQw6goS/Zf8nruQT
Tv5Z0YiopPlU19UI1v3wQPtk9Ti8fOjW3z2y6OsyFCim56y25R5Qvikc5jAps6YlhqT8DIH9UY2Y
G1KNVs7vvL9UJ9nzTerulyepL8uhlylyGGePcztKoN7djdiys/vYzLq5mVe2IEv6dVzRHs0k1slO
ajBIaBIvLODsA2F66hEEljD8tKvHc9ZVnjU+4QxEW+jyKS9KkspOM2B4B86L9TkppYg3T1gsjWuG
vuMnll4qFLmK3hESnHmuNdg8xSWq0solwlbGYw+zrL2owhr1Bhu+2R+vct0jd8ZZYHE00a6DjaXl
lH8FDos5QWN5RdfjS3u+OocrxcxgTficq8O4zCZJIHYq6ZlYQ8ieoep0YNrHrIHeuQgkAvtqkKqo
pYqmzw5daOwTmoJWHYUAtt+V6V6icslj/9cg8xHd3VOGyWkOsB92xk00qO7B5xgOrXFr5vRD/5Op
1dJ+GSR3Pd41HSFw2UenFsqVDYDkgflzhE5z0+DGNYNGVN58yLlcXnaL9tZsUKnCSAP9j37qeCkW
E73njSgBQZR3t0/p9m+DXbr2HeGbYizpJcJ5H6OJNFoRYvuEvGx2DDmHnjMG0LZvtQPoNz9yF385
W64CheW/SxFL4yJ0hn5uB+dbooBFS4K8KzEzb0urPfGhlKJghuZLfgwxOnyiBNItZ8fPKR5ioHfG
3OwYeuDQEaRGDoYeH42gaxy47BJKdlYGvkDl7U3JMhUEKFuSlxt42c6IcTI6HTFdFu+v+xRXqjTY
wpVBGxfYlIaCZpyIuLF+22PYeIwuuhwvrzMR3bp5xxblWcJf22AnHTPhg3I6bRTJNYvDXC3UZJzd
pPZS11wO9viY4k9moM0w3vd4atLIw9mbpO5efk9wvikYZVakh7G70F34PBCI7K4uGA7nIvlWz+M4
ej2m8sZBaMwk0EywqZ01UJnfmM6Et/OhNinV9SyASTJ8Sqgq9rehDRzTai4wqAQD40Yc4Dh77mw0
g759eH+UZ12Vz8pdyu08of+GWGA8cS/yYuRRry6HctVcKXH0DBaAEhnAuWfVoj4o99zrPGU3mhbe
GLtelTNDm/7Wqjqpr6VgrwA0BCwethQsZuJT4sVBrqaBSxmRFzFAqiwas0hCrBw7EdTTuW8Topj2
HWBnbIuMrCP/GULB7tjp3d+mbqPCJxTujoyWUfd/ZeQiGlPGkYDaLin5LoZ5okcPGaZhuaS2hQN+
nvaQMT8u+40rwdsBFiFhBu/EiTEsOPRpTSPccKaxmPFjaXRXog7UAiE1/gZ3duEWmmqf+Bd9eyyX
OUJmvBrEKdVE1A8N7GMMrcsIi9+cn3HB7mA1OOnzEfljZvhHM/UrhmvW6Irh7AHkN9sacSYSJxep
i03R5vRdgD5PsXEaAs2BNGMGqjR89y84XSJDgvEShu8En3yJPkWpzvVdeQbTejHRL7apuPRyEYrs
9Mex4UiLQCJE49FwX/8OgEJuE3Lih7j7pdaiJ8JV6b6Pro49QxqHojdhzR3NuPZiN6p9H2nyu/lE
WPdcBVU67n45B9e0lgsmTG8QXSGLcTNxMdJD5yUoX1u/h+A4pYuyfCOpRP2Kgi6ZXa9h3uOfdaGR
PiR2nEWb+ppKBHcPInWm85yahdEe6AZRZgjNVaykBr2IGZwuM55cwYsLtdMkgGwPBu/3opkJ6FOU
E3N6WdcawCPiSYUCxpr1NXTspwMLWMtlh6mA/4wGPmkZzokRsv7x+h/VKJfm6uZGX7Phx17GWW2J
U75nI74PBglXfT3612lAZgrslaD/7ZKEMWLCCPdU8Jyo2Rcr9GaZ4i2Q8y1n7AI5F5NwTTgR0cWe
S20H2RCyWUAvhdPJwsSHn715dCnUoy8ivfoGUiB45dkihlkD802R6GNAq/wznEyMLsANpJQJ+OmE
ShXYduG6/GB5pboLr++2bW9W+61/+h8qw+e6yC8ws9rvdJ1FCp9ILMOYpu1oUM2IpbzX4nwLuGAb
l461wVtu/A50tz1/qbf7qvwEBEDfpq65qL6osgqX6L6F1oxMAjCeRsgJfGDlSxRPbcJWgZuWEgI+
czlhGKu3sLBq5Rtv2cWraPaN2uCLME5Dp8m5NBUVxQwdt7SOXoXlH28aSuP5MLcEreNOInlCvxAH
h9ud4WHD4H9AuMyam3nfcOb3/XWcEGbGXUI1aSXnDi1EZ5AT7k502He+xVv3ZuzYcr3+k8Cvs7Xb
2mzyEpRvrJ3DLNn8kxyQfFB8pYIKqq2VThcFnNwq34W/fhZD/ck2KfWTHqt1cNIA939b7eWfhDb5
0Zpd/R/y/NbzDGsgn4lXBUxMueJCTiUyPLHuAfbHpWCUdLfVUD45e9levNh8TI6pE6yDGuTgyOLA
zMjaTw3bN/cb26iMHVKntzOzbff0IYH+O2Y+w4Mdmzd84mUEMjsjoMzdssiUaMx45mvRdxgaJRDL
L2d3yn+akapNTnwJ/ZZRp2RGzculaaT0Ci7qk3NhIMdYZ4RznOarIpXm4mbdPWVxR8bYCfLhkhHe
thuDGuNEbKPt4Czfiy4FJA+wzOjwfDQLGYLXfdQDLtSM3nC9GXmpQxOlO9EcNxmX+wKDhwMtpyLV
5Z/g6bz8DSIrXkcBUmz0Dm6+X/aglsgxVTskyXUPxnK7oBViMmHKPllHRHfQJx/yxLyV/ctvv0mX
0Vy2pavy8ifidwLSvX5I8ZlsrJLDyAoNuZF3YkIV0IBRVJGzwoxHCI34026bKcBk4s/K2Fl6VPNt
vGhZnlwTKZaMU9TG2p4WX6HpCJ5GKWh9iT78xxjb9DD0cwz3uzI/QKzunzX0ItJKX142UxjNqjJV
tW2ha4zI5XGeFZYrhWtNl4pWUICbRMEkHfm7jchQVatAqNwNX/xdAPAZXu59c5d82E6yFMFRxUrO
lve5YnS0B1+WSiKMocjIv9vGbJPvK3Yoxm/RsagzvuyNHCSJ9OpGHF1OuVF8sx9GLzQ5TZ5itUQz
cote2zrENrbgnYqIPUfTrgV7n0qoXC590bu6i+wzl6HqUrDeJQd1Kfp7KADxZV9FFiVnGEZkH9nd
JeRvaOtcRhrVvFDcZVX98SI2t097ehOjY6TSq80GmBBBecMo7XCsD69DZcJ0dVX3reBreaNW2nNd
x0/25GFU/x3Xk/z3NdB4hU+6C9UqhexnBwVOPPmr7bi7Sw+Jtt7maUnpV3iRORnb4mnVP9yjRWv1
eYh5jCocZj3AXmy63XPzHi0k3vhrFpvA/8HYnsOi7C5iMDQbq5CzAnSLR1s8uQg4kgnOJ7ZVGKLz
9qRwNr2l5YHRFpaAPzLa5PuB4dCECAl6SHYNP7bxkqqCkC2UWzDpN6EkrpmTA9DiKnBIz1lXDliy
5zVYSau+xdhFsdgpVZF9AmKkx6MGiqvWSiCpijUiVeXdMuCFjR9Xm+Qa7fzCJ6bM6T5iy+yNd61F
m/dykOu5kvnhLofQjnQO9QMsg3/DU8xn7hUnr9F2fZ1Grk9IvsFYtKkxQjeNGq4bQZh3DE4uCk5u
xM8KmeUr1NMu/b9CPL5Iz71m6NBp1sbRLTwU2hF7pKqr4HEVAVZ0XIbctHT/pDHxE5BOvrYHGDse
6nszod91eqNYn+ALKmUy2MQw3jIVKS7V+boyhcevF74b34q3zMHG0TW/AQqFoSQynDHftRqO+win
XLYtTnp98bkqD7D+X4PmWpg6YksNHHJJhRBd87h4NaOjJdh9SrlXbwJsp+4wJudFus949IfQE9Jp
yfHc79tpiosu8zQnjjN40Is7+qwZTA66Ow9cRvFXyn7+MBg9P2zyLnKmZuSMHkfWR7pj/Dj/86vx
PsQk78ytrTrJiK7touwA/naVWOcmjwaqn18+rk/FUlv5aSU7iRl6Uw2C9h1CUW81NYtxE9Rl2CmD
By4NErqrXABO36irp2S1+0Fp/z7vCgHR6rqJZyBpzOI70rkhSXhJc6n1Phn24mjKgLGEzit1xacD
c+k+dpJ+PJJk5YJvcxSnD+4sjh/27+z3/21kIQLBblES1tXJBx/3w85OO0WGhwFedW2eQXjiSTHm
8QkBP0Ips0DR8MzOzMUBB3IswhfEmBfB2HWj9ykblJ1OZxna4EhTC4SX55uCRTODIkIWebj/ZYn9
cmPsjNbSwTxbLLvUcN6lyhT3j+cZgXk3bJSStJ5dLoT16ixk61qZeAT2GRmDwJ05yKtQIZUYb13t
UJkvH1Pgws7VM9zqk1qDLSSffpE4iOEyaU+TJg9QQcxndiJqFg/mehmd90qp7VyGlPA3sHncNkbf
ABDiMPJVji+/8NPswILP1MaO0Sci6WdAHDbvfzgyJhw7mvYSK9ZyGm/UE3WWsUMAkq9PTo+WIFlR
KAvD85nOCCc8Ep84KA3YFNpryXP2WUw67hSmicyRTydwzIg/D4jhui3ZFwomveG2FvBDxNr83Qc2
/HHkkNVJkBHgWXwA8PM9A/EW89mk67eyUf0MQ8EI5ywVxyJwmq5vMubaR2jTaqw+S8LiGwNTV5f8
v83From+7PtMg/LFd/Ea0mq9R5DhuRBhxS0Vq+h+e3fWwfHgFHYRXRwgQfXLX1fOcAyoZyobgzt4
MkSVf9/MDj2SVUnvaxD9LqmR4iuAGkF8ZQdXGSVa7sL9O2tQOvBJqY74fGsTnW+IgQZNCuz7M/mY
eDGdWf6r9AjxwmTTImb3pm8KvXw/9QpCNaiGcVbF8rZJhHC82x0Fa5QfHuio3VJ3KWa+9yN9dLCw
dai9WKEGq3ybMtg5WuJoudQ33woCF3gIQq6RVAkMzSWAN2JY3AExjAsm1MD7TaxWvsym2udsydjy
zt3t1b9+6ni3MZzdbGOkYObuMLKBKsOq9XWiW9PhlfNqkFWgZtbfqB8FilYA8WwGlIsSxDFHYGqf
AYqf5lq8qIEUZsTvQySfJvHuhTgFmRZOwT54OBufRIUDvg2vJHUyQeZvTqCqpQke2DApOg2ny4K+
vkg+L1nnE6ATI2/9VBptXPDqFIgpeIjgkHrOcp6HaUfIQBBjiUjc7O3N4aCpR83EMi+athAonDl7
TYc9zVzbLltMprTWWmJGqfS4MyP7zsCEgFL2QHJfE/1hNYhpETf5ntxtnBkPibPSBHmy2fheNodA
NPVXXE/15K/wtrfea9XwBEY6hVlNw9tjBb++JbXpjF3/+78XLhsBK37yrd0pIJAYa3c7e+HdvdAE
UVo2aucY13VSc5KnFGqIxeIlmFi+lsehMaBQ321DgXXP/zjCDigs4Kr+VV1kf1mKNBrMmlmGBFFj
1IsQgPxipcf3PQF6AXPJIXQv1M6nbsQF/u07Eg5QxGMHm3B99pcnBfrUSUmp6TFSNockiwIcbZfv
Rw9phcHxWeg1wycSi9a0lN1ww3ut5CBG8NVske3O8Anf+CC28w41SIuvxLDOL6R27WTNMEkXQbtJ
6uUdFhY1kNwQLugphFol4hlm/cUGEcOtLFaYxqJMlX7I9p8MwtsbGL0y9Pmzz1S0Si4wdyvw1gEW
JGZGrOqw7FJPnX2NlB2xCJQDrXbc52kuqQnMnYtCtkpQM0FrLNWYYRX5o//Y+hQzCNPXeipryz9E
t3R3Vu8McPEIASIacejOxJyccdKhwA4dVCsKncrdF7oEsorhwMW+fWeggnzNOrnUXAD/NPPFnOVb
fn1kT1mq5IXea/pi6dKf2OFE8bTAtiMZkvmRTzNdsjMiSm/0Qgurk01XqpmXCxh0XxlSYz1FljfU
4D6T/ro34aJQEc80W7Cdcl3zkbY9eJ69SU4fRmBB54RGZQ5e9hdbgc52jUZXNuyj62Tqs8iSRMit
AZku7EYKa+8dVZzxSHaKq28Gn61yz3BR1OBB+70ee9f95rjc94kPG9cig7gZMNgIjCgPYS0jaFfC
VGlubTkKTNDbU73GQnIaDEHdEAsOS19jsBY0yRRiRXVrqyHAEMuhISg1G9dUUa0NWnJKmae4GtIS
z+DQMNstqbobgSD3j6tDOdKbco7Si0bq3i72wAzjSU83wZ+n9bgmEBRHJa080QjK/L59YgmyGkc1
5GLhf3oig9IS96Q3HNUiM0byLdWDPH3wcqcQr3qLvUtrNxDFDf0+/vfWPM4M2brOX/FNcAFR8ETz
5jvLMhJn88SiLFaYxoq7pyRV+kOuWNkuBYcOY/U+A8tedhMloiBdOmhtC4UDZgFRIYdMibL31DAe
kvPpTlX56lawb85bOgo9hlGvMKOqoLqn1DiBkJos3zqddVGsgD4p8t7MemLJ/JcucpmD5DzQKUfh
AMw604otj0Jx6OlvJsFf3vSgKrjfy+10q5y5WF0z8oHlwdvzWZqnN78w7n/vJwJ5FM/yDuWA511c
vxDlUpUYa3VnaJ7UngC02X52YsaMlB0CpKLiNcgo2NX73SOpJxhw0rBdp8IdZmPQAVO6ehPRBOxu
UeCfEmlpBlTOhY7jTpEhQ3wiN0VS2OAThJnLuR/A5CF9hyv6ZTY2GlwK1H8Pr6ujwnBgWy1z0wwc
Y5dPqeb2yEoDqMGYtfRf92K9FzpcdkufEtB3+AaOHvu91nV4eKuqlednYPuo2nxvCRavV1Pg4Luo
QX6iPwYRN6BETRvgtxTbau8tor0Zt5pHeKs2H3ZbWXlKf1/wLH1lQvebS56mlLJ/8ODXDfuyMQEB
AvOi0dLsWl4V4fk4iiFzbEQ306T8tA0Jwa0SGqXbwISMAB+Ok4a/7+FY3NJ2tk9ZAmi53PlPzpJc
j1F9aj0OzZ1Urkv+L3d4FgK7vP85+tuBfdyteHMRtWMjZUx2H8MmGM249tH+zFtku+6MLGsatA0L
xWXHcEdmTa0UQ2faYHAIINYRhaMuiPoYq3Es4RdO5IM+GtFpjaYWuDsemYnehvuM7d5aRwf8CQmW
Dn4fvAhuYKoAzGpbQzX0fFbVshcOA42oA9lJ8tFKmTWVQiwdsWLIYTwG5OF9OTZe11y23uu09phZ
PR1CeOLU1TI/a+a1lPdFPrWEKh/IIw0BhjZnk0Pgmz4nxykdhUvgA9gux40yixe+QhruLrrHDs6a
vPCTf/UmC/zDpLtkKKcTOP4bYkTwgFW5oyzPy+DOt92z5/NDEDICdlh/sx9DiZcFskqB+7/H64Qv
O91WsbmAnk4mSA3jJcuE8lPD1dJEYVB6EAz1D/CFqF82BZMyluyN+BecTtf6gyhs5iDYIsHeeUyr
UlBPtTY6uIvHi0dD5eu+gGIMWOJ1jEbScPKa2V7v8y7wlBTpQFKz7rmF3q9LyhjE8pZFRF3cNYLS
9mJcekWtrNOchEdveGa9CD9FFRLZS0IHkONEoXssFlwZdbH+PKsIUsUamRltrlkgM28D1S/OqXt6
4gafQnZBToXhXYPGeVIsGO+l6Tcz8vRl9YJ7BPMEfMA15RE9ewKqfiCoQs5cQX+Q5w34XN7PD1D9
w5T3fztEfW+0zSMbxJM6QF0o7z2OTNSjHnWqmSL6nac7YpxixBxajpDAYCjiiSUrnK+P+pwVBGCV
pupNazaNDfoPFcZ9YHtMLaV8+16D3BTdSq7n5rotADUM4a7JPWvpBEw4CmxjfEDw0AAjpdaKYLU+
yasNRzFVIHTBEfXYIuHkYJufkzuu1KrRCKbwy7RG9u24u+u8CAoMXIzo0obxcO8iRC/oZogfjR5d
Ht7cjfbi08j3vT29yXjhbKRPYvBvYkDqW093UWE2q1VIqfCbSXVwlvL5f5zZwzXU2Yl0+1BTqAwt
dPRgXoETHu6nO0eHDa+EaI1jiXgNfo4L+RXT8F2yIIRzBtM7ulnI7TWZj3robEfVjOzeFXHZAaFC
e6DuAU1s2VPvGc7Xqh14hdvYvmqmoP0mwqVj9Gank+Sb8wMm8DL4odghLjb11G0SkE5ohqB903dK
QQmclEFPP2Gv+ON/ftz2Qzhs3oVYsNNl4kws8kVN0usWjalFZTXJCONfpQ9TZEqswGkxT1ScPp10
0IJQGN6+du6KIhum7hkMicFDn12v98K0rDTygQiqlFwcYzScHWtxj3IU6wKpxXZcGxO5TcuEcqSy
UDI/U8P8jBLrJOUm20Xwjv088d7eZx+9DFiij33Tqc1KgOu/iyNI0pSkrdsPU5fhWamrXMChcg+K
ZyuTbUs37n88S2/FLecZzsviJp5sPGkvnoSPU92/qBe76MTWXVDdJSMSwb1r2a8wLamcARQsqTQH
Xl43S9mauMTxP33EYpD+OXF34BS1iDSb/ip1JPSIuee5e3Bw/h6ghkTOjmDJZD83gWFvAwhkaAS7
zgE0qxK3j0uxkBspY6OrFSJBJ+toS2MciNvLawcMb/e0LXgLFmGTpHMZwISA99BvRAZ//c6Lrojr
g6ZgvpfMRRFYqcumRrN25MD62TOAJQLpQmZT7b5vWBLw0YOAcxn3oxTgJ6e647DEQZ+hZTNIc5lQ
meRY57FCmdRBWboDRCPrJ5DC+WmYzhXhmVa+eQHCnozTB1PRC3QeMyp63Ez19+w6CwBExrL+TXal
0nbt3JUNwQh4iFEsk6Tb4bEBVsC1/kOrIimWfotNlTfJGEMXJUoQBzzSOXxWtXBUM6TssGnclzn1
uiq4XVIEHoxvluBZtsDMpQmut2WFGiS9QOyRcOdLIa9kTjFufr7/w3sVx9+uD0stDPeKtBs6OGJc
qc23JEPHRpqRCFZ5ohppi+IedAI6XPzQ9+O/RvhBvX2XIYLavztdgHxRILRSpLV6RV1lSlDpWiTL
bnXI8DJeqRlhcp8CbcaoObHV1NtN3GRys0WUH1/Uou3udiVDV4d6lUgYv0wOp6KX6neEpgu8KGQj
/cqjoRVHFG2nIF+RuZTBS30V4qV3iUP/nwP04LBjftgktzvUOaXZ1Wx4aVCDQ5d3OqmU77XWUCoJ
qD6UfTttD7Q2qJOJIy2Y1LaMqaAHvClZx67+F+QhZNPw/SNcX9lxsGSJ9zL3dffUfdS2xjVmU4L+
c5ICJFtQruFWRqPASqIIeV+gG+BHWiZiY3G9P5B9jw4aooLQu6tU4f40yQ0or9wAPC0vvSl4cR7A
QkysYM97WpgjWPS35ln9uLJ9GgfZdiLwS8B6BHc6nzqgy21Yb9O33768LR37tZhZ5LyX006r3OLd
e9vaBbb7NwUcpypKSa28xGsT87sv96wVPDl8DwMib+rG7NlQuDeUuKjl8AuwxorAOH3Pg4CwXnk3
FYieqr15hZoacJTBsQENbuj7sOvMBnQhi8fntyv4S3c/OEhixs6igPBeapt1KpV47SxuqpCvURiE
/x5n/ChEBM2gY7R1uasaffzIpsEaUvJrNgnolwQBC2FNUIwF60jDcWK/nTnaxzBblO9sIMpRwoil
X2WNwfxxnojn/zpPGRcMb4kFqeBEU3zI88uQR5qKbKk+nbaRracKozIbI4LXRlIptZ/43B23SJwQ
4h2OhGRsaJKPaW0LCpDZck/Lz4QW7WAqibexzn0HHl0IVS8in6w+LhzSb7i5GFNNTti0q2NdfKx5
ixsIWTWA9eVvf7rrquzZGQKCuoi1cb7ZQdTOBnO/GB1eSlWWzz/MFD4yphqyEttp69j0eXnaC4pO
Nx/Yj6BmypJVC+MIJncFdDOaByPld1wMBG4GvyN0pfyPJmkLPS5bi0ZoB8ZjiPl3mq67zK3IR28g
D7/8po4U4PoA3RwUv3IrnmX1nIpHES5kibARscBOCNy4ZQtloYAvNitylZewtG8OxM06iFoDj2u8
GIj2tTIO26/0MBuMmWiCxW9oa25t16U0NQ5uANwoJ5N48tLpCm8ITo4FM7RecCfvHm2LiXfbS/uB
JBGgw0REYdalLbJwPh+Epfm2R1uI+ce+DWglyC0MRIVn2RTwxR1gML8K6ukBOCNrYoj955PgAd5b
U6/pWbQovcr0xpCs2HKjHjCveTVGBhaFkltmJXZscsJGyh0YvWONzeY7QyJNGHlzMhvPagIYKXnM
+n+g15KBjKDFSmnV2P/MxcOojbOH+/9iDPsPL9qqtWbfU2Zwzg2Fq6f0U3tm7V6HGvYUtkcUqGkk
Y6MTVXQriYiO2qUpM7S7XBmq2jZstW62J9dDUsqXIUv74aL05XSfbz4woFx5kJ8PLppXcSQ8xFPE
XDYYCVfdE8tAHl+Gl7Fe0MFk1PVJSPxLoXXpOArcAuUCelOf1bquTrY+GpR7sOo5v1gvgqj6fw9i
p7jeITcw3CL+8K8A3bO6PQXCcdzZ6wbpFPlYbkdd4s5T2l5j57FqT5nPGpo1lvx2LDq6Y0nCBNfw
OjsLnQwZ4sufnk6q96jyIGz88Dly1ILBXHMIMeZo4TVkrzFwpk3rryt0FDrB86svepEcXvc89bmV
10tq4qzJdW7u+XWGfKhzgl69/Fz7fs/vQwi8LJKVMVd/9sbT4BSnp7PtLUmXB8kiqmhAo3KMCWTa
ZSimeVHqipv4J0YAncj34lLRSDEYhwDWTyHaJ7IkXnQg2TqjT1Mql+K42Co02OcOh2/TO9COuyxm
QMkwnXtGwUXUNNP2ijnoH/DeZSiswNbsWgG8Xu0MOOdnxqRG8fILo3Rw0MZYdHx7LcGZEDxr2j8+
9v8fsRsesmdA9YlztM9wNXuYe67S+piV4vT43Hahij8gxcVkYkgMJ5Fh/nHA5H5D4eXMUyn1n1Tx
PbgdwDIxys8Hb2i2p6KUsgN0bI2xCiutUsiZ8+arLtT//3Zb5/IwbKhfy2qnzpYHaWImFVk5/lqn
XbunIF3coOD6phTJ1Eo8E8SfKW5m2xRCxrhkg0Q0d2INTQUwASjwm4wogTh7ssyt9tyaE6cJeyCO
e3lFcOs8BNJJZ9jzy5tVi5Hp5LWN/57wHAk8NawClj71yu58BDuUH4X/dYnkZW5uEtAIKh51dsbh
yLQ4IGYZNl2mYkwLMYwAgyMMAwmb46Ospibi63/c2G1fKMgKUkkNP585QKmJi7UGa7tdD38nr5cE
QVPZFKZcE40RYmDTSkLohJV8NMe+NPT2cNO+JzlwypWYlBAFMdIWyClL7EnPOiJ5QPAW6xd4g3fo
fJFnbWPTtPF036QcS6piiRHVD4TEmE04ovw+yn9VMeaJd5L+xuKm05zFocMR8Tt9uATMFkZQt9jF
sc+I5P+opLPSSRcWgAkmkwe00mySzAHXysLzIKZs1y8wj1M/T7W1X1B/WlXnYCbyhRCws578xnJw
i8AP3F7YNnRdu41ql8/wPAg6t9qDwRY+lsnysiu0WztyxZI/qVtIFpg4qzAtTCd58zjcmKy2uGxG
6knVUlB9shCupBUbOb8GE4GgBr8F+dwbb+HKGuCKSV1rBw7tuOjwRLAAh+ozP9uCsH6M52sVGPhb
YEV+u1euycV54ikYNg9rO2iYJmJ+pvXbxmS0ztS/EvObUWl+JZkWjoQp/c4uruFlVDjLTS2GLT++
gMR4hfN1hkGV3GGCm5+6HpWOGlkXsevGoYKI+3pu7mGWg4R0Q1YBoZLmVEa/ke0/N6M/H/uq62yw
lfZaixoIRD/Kvh6V4KIc49EFlNbAj7Wej+ibwKjhqtBercrf5HOtRL4lD35klW/OITwku2rF7CH8
u7BDrLTGiJwQzw9/5IQg/TmGptlqRXnSTOj4pz0NuTwKoFPmaanIuThpBfemeYYQM4sJu8KXeNu5
AgihocDsDIMxFE2bz5RkT0elu+jS48Av/XoDA15KjZWxGlmKBEREpaR3A8ZKz6xnopVe+iNkPeuY
07KAh0Q/3mcsNVsHKshOl+zrMuP8GLzSgCY2YzXwDo8DN3Nn5ouDq+q4pLIhfevCQLj6NWZGs2iY
3H4NgsSK2NP7VRAtHjpWD/fHjBCTFij8Ua9iQOaZzUJPi7qSXNgW9wCxw3gf8IZJQbsvnFPQEK4V
b86vMmo5ECm097VcSX9LzTvmT06pZd0yf2byVHfRK2p99Dz5fs+EsXnK/a1JhVH1tsISbGjV2p8I
26CkLzrUmCiN+j4VBffvTUSZk6/hGeeWJs6+NSgB6LCRmvdcqhcEPEbfKKh6KpjoLVmv+iZgB/e/
Fz1w1duNdDqBUGrIIRkSX5iITxYCi+uSlpAx+O4udwkNb6ZOzahwU7RiPPG1mRDHSciDF7+8pkB4
Rc08twArrh1Xu9dmLj8txemWCLH1qSvEnZWiv3u+MQTwsztmXuqIzcO0y6+dP/+M4q+nzkXBdgQd
OQMKS46yy+YE//SwHuHofAdAa25R91OxFs0pp44NArwj+BH+yAg6tFu+4S+alXwi5p7lcc5ik7DB
UgZ4L+Dxn1/vF3INhsxsb1v2Iy8Fv/bdmJMhd7smOzhCQdbKpE7hqOKLpDBSKqSUiqpwh4kKIpSg
8l/89sSwejkJo5AOhr+4SrhzKOz4u/CT9XM/euyn2WM5R99PYrAx8rd73FjIO1HzYcNuXmoS5goE
OrNIrJTcVoj4XwIJZR8azZK59IDoM03wGLTAv3mzaj+oVHt8aC5aAULcMOnItwOaoXosYUeLUdJ4
IEOc0ZcXnbSbDsbFbdTMo04046eQG8YqjUpQWjHbN7Au5wDolD9gubssntWF1gs9Kae7If4K05z7
0mvsNLCC1ybPrkDFd6ifSfxq+7gamcHfbR4zed/ZBP0Kan1E1ri2OE13Pptp+ntHZvBM7zXoDkqd
p+5ybGAy3VULI/pLo4WBacbmK1Dj1QSzXU6DEWzNNmbPMYdqE5hHNkZscnRcyYriVTVzqLlcX9qJ
AweIBujd0cPBnlI/hbfuu7WghYhVw4FgDY9kB2kxLnbB5eeWUAwW+Jo3EzZsfOzQkZnAkRKGdhwC
vq5w5ARldK6mecQi/X+sJshwU03YLIfZ0HgAzunJaxnbK8HCz0/7egqyUGjrfeNhXTJZIeJbCn7j
Ez3jxQypJa0HPrHCACrXVMHORNUm1MvtVTMH4sm99hat93sIA/MpBEtweWKlmZAyYNhmfhlSmHI8
zVnfvlRZTYnl0BJjLdoDkDOR/GRA4CzhVoqDhiQHBucfx7aGzIlDsrpTuX/wbULAoEgeU7HyHXBn
MFdGJg0Weo1q7WLtCUP4F3XO6ikVRjSf8vwVhCED+PkjLH7/+jGiJkcGrqQ28bno5cXTcQj+BeV+
2dIpbvjLT6IOWkmxDt5wE7f+83uix7/9UMh6SwhIW7h+ZczLszSLKPv8d58VbeTU5SHnowZjkWcD
VvxG/gitmkzx8yzpkyycUhDw14eoSHDPhWGMDohlCpRHti5FT30wViLizKbpvcbobx7CX4N3oayC
8ds0lHn4Tj09V0cJMwC/R3stebfc3yyk5+MBcF0B4/xMKP8mg5hL2nYA0fPjjmpc+lqBP71QkCM7
SgDDUZOyi34Hy/2XkhqIPs4UggbYK6yWVFHYXr8HUxp+l6CdPzyU/7TTsuVU0Hc5m9BqgRl4aseP
oeCebqLmUJCX26TTBU4UwW2UbODPhe36Mu5QQYov5uuMqZ65FAaDApPlevfy9d0qdUXvb6EJJyNe
pCXiCv4v/2CC0bUl4OtaSVzXenklzT+Eg0Gl0NNmco4dMV0tiPBoQR1mUvNn7oYyJiy1eTdM6BLn
dme+ZaeoTiUcUr9vuWzpFQFFuDUfJiKizXRe/J8Tdi5Xvfgila0zwdWD+dyHz8o+4+2T6Pw/K+i7
ghqm/AZhjhuvgLEEn24tpmSx8dQtAKxoHs03m9bt28535CAQBdzwgS25MKYVfZRxnJuUzmZxzar4
NP400jUF7nQAMIETKfl5kF9V9bBIr6lJLPiDL+XMRCGQhtnG6ML52tREszhYzDONueygJ4v2odOG
y4V7AADQhtoiOG3aM7US9PGKbRy0zCZkWhOZHCt5K8vU6IjpSfaoiGp5/ojXpTEFm++oxgAVdW7l
2LX5YLXgHKzHXbQ8pBD0oCDlv5PfDxYdsHyOPl3KQYsc8obuxCpbYuysELEYjx1iYg+5vQf/p0oU
t2DKaDEpQy77PzOaUItbUlEzCBkUC1f0IMuWPNpaKRcKYAOENuKulxYir9kUvDffKvEUUDXLZz2J
v9YjQOincsyAU59zbabbF/pJfUPyAIRh8cT8sgO6Dpa+/2WRzcSk6bEqj2bBKYSTtoKew4OnsPpK
zqlUEQe2P/7b1QTPVPm8cuji8QiUyhpfFlmN73gFnSao7ZI3a5aHLaDUwczz210PQ9gvf5S9W/dZ
rAPe0hUHr5otYs1L9E8oXkqwfOO/jgQNCmXAk8nbmvKcY10/RwoSYZHTf7kBFpiNzlkaECHXX1+p
itTo89MYuPIWB2r+v9uMLhMO9ubDtm9PLlCsi7o3qXohTtDmOz1srrDfTMYzrwd0tlfGqj3tj21G
mpIQPrz4h73+SBryMs56EYcC0vdT4nJVmQX+x2UMNdU0KoDrgyqiYqUd2wHlW+EhrwhSSeOQKmFX
EshjUBE4OqInJi4mOdv87TGnvaJ2/Np/WHQWRPiKnTVO6xafTJkOOUdDzpSIuEvoxB96CdZcxxyV
3UIxbZk3jawnpHjE7bk+TrJapcrK2/WVyFlbfS/f3Q5Z2PFtmewdWKzZRl6vWumJ7ARd0RSYvi5l
Op8De1J8RZMmmhqJPWPBS93cbliX2wUuVpCuZejhRCUqsdzLpPIQP7cR3JsgjU0SfCo0tjh5e6AC
BjMoYZmQv4XeaRop5n9Hqv1/h7Vwp4OF8LzdI4lATkHXdShnp5EX8ac2TC5A6fsr5rlsz8sCoof5
LUYpmGZtpjSGTQ/4IQt3A3I/3VfKchs979d1S2Q6JAwt8ZItTJT8VtlYQsCY7nliYjeKzZocsNLq
WprnqEcdQmkpyT9rhRdyBW2LEkhBNTFJYBtyCXGvH9azXjdp0XKbAhPgBCtQA8Z+hil2Sy8JXMO7
2Lg1lfwEqUM/GeJh7yQgfEoy5B9ok2VfjDq6A5U72thsEhJeEYZUqYXv0bHqBw5ngQb51RM4qIZz
9V24Q7SbunidMIaZjvT21SDXZi1z4l4tYq2R916MGSrjzG21OUg6dlL340SnTuRXszpc94jB3tH9
6dEr0zRVGkp0XdA7a5M3cvBFjxd819cziTnxqkuErTBbk7vbZ5O8DvOnHiAgCoQ6/JDQaSK6jglA
t0sd5qEelZGYvIgWayBmzo54VFp2CqZ+qhjaQu958kRC49IzmFLnwtuQ8mBJU9tFahgaNIuyLugZ
+50VFDcMhy03h7eV9Jvz/kdbI/j0p80J2krU1tPJLCbavd8h5z2vdjmbdRBk9ql+QebpY6FZ8TqO
i215Ee8n4MTHy6FdELVOExH762H+i2iDzGF6rg0+EVx/go3ijRanPlaMU2UjdPlQaFvXXBhQDyR6
iwIFH4GnJvIyOecjyfvxJLRwB6LP4ax8UkppqSYX9E9Y3jiN9hq50xuPKp4nsxZ4rriI+Fy61XbT
Pq7UXoeWwQBaprjiFI1r0QrgTovVAirSb89EEmkAPvStTibcMzfFNQblijK3qqSQPBL/E0GMTWbq
o5YgAO6jv2lDFWd5C33SXSlK8oP7BGJPdOfwSz8/pm9HsEiTU+HHpo0j5qJ0Qr8aekTCUVhp1+Lc
Iyr09rFzz7T+5lEwMihOD/sdWIt5aKhf+Cv3/Ng9ceoucE5fAOsrB6sl/g2TcUeRBYf0HlxyJ5v1
jRSg1LFruaVOft6HTRfLOAC/CznHwTqM3WrgU7qWEK6ktedKqxrmjkkHI2B8sMW5szXMjNHa750z
VbVuR1N4OwT7SxIn0q0a1QzyghARayuB7XYR9BIKtDdP5j/vitDBeE/f/ZM71nFuWyg7TKlsEDnM
sdAdYzerT/WTgzFR0Nh43x8Pxga7ZYwQIh4yu4suav4sNmXuRKyD654A/s7HZj/UBZkIdpdHE5p4
5KDcd4wUMxx9tZqgeM/AwoFs/VQWJbvMpsGXHYEpHmLxe4ImEAtGAEcHfhSXY6crB6pdKmwl8E2e
TPB5awxf87+D0Ss9jPL8nCT/ngIpWa2rDpfquTVGlFlj7sTyshVgtROHZokE0O+SoUqToqpT1cCa
nxdQw/AA56ZKx3ePMGi/CVOhCd3BRp+A4lwd35CY36kNIC4zUHx2E2rrPo8UMTIXH1GDXm/AKroZ
aHZ/fpvrg5uXUlnU6Q+8M+9Tl7IWrUS2T8tlufvJeLG3EpnIlZzXQ21mnNtctj/cKuBVFSxNBeNI
UGmbSLrgp/fiUPUAwNIbj2KoJeordSMiCwCUJlgh3QNx9dxU+vSRvxVptBKKAvr/pDBAqacWudIZ
49BsJeeScnLqEgunQIruUYUzjR9pDo1wPwpUugu+gTPqJ8f6zXDUCfCbiDQZ8ASzqm8oYX5+kLnF
Knc0dezhFJtJagaRsZKjVYZsprrw4YctorJOpTh6cC/llvfovp8yUmE/jC6XKgcoaR+no/fmdr9t
VvwUFKSm+7Y9ZPmTHucvrYVSl9rV5LTlN/16440bPmwbQYyJhkzMVT6YuTQtlxK20lYilMtqknGp
HR151yWdickGgypgeUyAnWtp5xRVT1LIGEDhLp54iovefAahRlzfLv1yiEUU7QDFXUEGgSm6bH6h
GnQfgRG9u/pBrcEcT+sWcNSepY6skywFXVJxp+FGD1E24YGp+hfeKnvNBssm3L0XQV4CTf9t+FFq
d7MGbmrm57n4S0ST21y4RWsZsBT4MCkdt1LFD5h5+P4XLFa2RsyeW7kKZt6EAMaXXJg/peJUw4PF
WUudxfQLa+rCl1nl7slnJnA9AC/ogvnTDnR8zyGHGbdiLZKDzWUwbSBwLJ41vnDrWdytPKvso4r3
+nQOTErNIFvb0kaUSoKaVe5RJt/ZdfiZCFp0OQ1GVYklMmetrrnz9L14ma1Hd3RU6JqlEyQvjILI
izEMuHVnwEBZ3MyNfG96xopqETWcWCTV8zlhp4ILlNSFK+3GHdzpjLA39nH0niRDBKdiwsoNWbUs
+vXdCllCKo4F9NIxVncs1Yo+xtWjfKqCi4z5eM29lNBKP4cEZaMJZkICyHE/rxXuknIlBL/fFNnL
Tti2BHSzR27YyI4JF42uWCu2wdV77ryOmOV6DkfA9+GQy8I4ZGoJgThcM4H5GMxxWc7dDFfXFsxY
Lrq/ypy59jbeIQlKQFZUh/d0oWXy8ZF9R0R4KODHsf3F1sWKdlV0L5yTUysh4Ks6H9ImHUGkQZAW
H/IhCOTBewHQ2S2CtjJ4pTPJWwlHJEO4Xb7l1L0Lm30VpMxshJhwbJj4gmg8Oye+Yauwz1HuF5Cq
ECpJEtofPPfrcl7eJKTT5w4pIP4sZ+19Y4e3fKA0NDglY7pYK6lN27E0sRILKRcsPTKuLJSSIhjs
o8ONkbmTy94EWjYFC1/2DTWNt0ggC939V9pMhDdj4MnMM9yFo+ZLPOEA0+HT1MqLlGdB46619wa2
2zeGCq8TY5sdOiWgJiMjlAnY55SFsjljj7DKFEH4aXAJum13NiTLEWFV4N1IRGtzhkpFI88zHe+0
paKI3uNEmj7C8lX7/NMar06403fawEY1r89pinPnAyy/Sx61TYPnDl+7jlZnTNe4u8QJwbbT7rWX
0nYG1Gc9WTu7GLOT+Z/iswveJ2H2aRqal+5a3NAJ4lDceCLj30Jn5rxW6gcVcArkIZTxEylRfCgE
FY0xA1CiA6Xm0B7diEy5/NVHlfp3dsigy3pnNJWSVweHFTMdiE9a8bW1orr73KsOOvnlbnF36rV4
OhKggL4yYMdUfDEt2o2OXrH7jTUDVb2CNxO/pleIH6ELf+WH7ckxgUqLhNechQnHbKuJTAy8jXAX
k0bMY/SS2y3RbtLEBje4vtROjKA2Gq7fxYrFpsA52z9QxTSYnzrizAfloE2hQ4M22WnM9HiksvWP
cVddGDEzq0uj4AFdTm1P2DpYH/dokwzIJVG2P9KIN62c/xfYpIWriA9kOgv8zU2bFpV92fNcNH2D
C7az3MmzRQSi48DK7JwnS/RBoYAr0KSmtjKCXo0tba/FgkVBb7C40zEYjLQx7lGJ9u5me31FNT47
5oarYlOXD1B/wyv2bnhSE1D9JJTOy1/t+Gr/rZKW9VV6YiKRWHsQiyQUr0pRzvVRUD1Q/92U2LGk
nLOIWE2j7nPtG0PsQGjEbBYqY6lUm8wO43u5jQEzHzTFVOTz/++O9jToS6SNvVtGL6eAPtI+kOHM
rHUOUxtkDFFAMFqnWnAnCi3Aeg5oaZ2Ri9mv40E/SoYF3e7Lfuwypd2LrRt4C16M6lD9kv95XNap
rnY9PaADeVRsCALlXfko94HEoQJYuogvjajtw6Xey1XG+OeTdL1rpKNYD1ro8LgFVvdq0XlFYs5n
K/tTDGcxJM2lmjYRcDiVmpfsaW2kTVk2ysRMbLbhx4dewsVILCMW/TL65ZGuL6OrOA0MROTaSeHG
ZpEJ1YBafP8JPo+kjxyld/+nZ9yC5nORHJQNoAmUT2CAvHfmwRSaoNf0RjAUXeIwWPmk4AP+N5co
8zG5ySpLkljD9I77nJHNwYm9R115S6AxeB+zotxU6bMZDpKvu0SjOcosCt4IqA7dsGWa8C9pf768
9sOesjwHKJVL8Rvz/ASj+8awNB9VXnKbWXUSqmo7JoJQtNuF305OFjknFO2kKzSL7FN/jTXLvfeb
raXMU+nUmwsmot1KS/PxRSpuBmR1F8iTY6IEtzAYnV6lG28gZWMV9BU8Mgp2cTgE4ri6a2ZnpGsw
kFvy2z5yciRIuV9jzEA+a9+4jAFtbiaVz4+bMU8MMzwrVbIToLjRvxSHVU7GWj4akpjyX0n3HC42
upLUXDh4SFZI2gtoccoAPqkAE0+UbclTU0j3PilqJ7qpq8qW/KtcGAblaxhiyn+L92kfNy7T2PRo
NY+wV/t8yia2GxpqAaqwO5PejWQCpNQVKcH9pZDT6K3KGeFKJfoSWWGVqAiMwJ93cYiaTs3Xta98
rRszyLQNV5h+dDRKvgcQq5FpYQktfQM8IQbOenOhGhto2Ni+Fv5NH5WAR+E4WXmOCyO1l9nIpEGx
QEi4sspVPxh6SaTs79ICFDVK+bjAMtu/KyHRUwHCD8Jek2ux2HdPNTvWcydbvLjdAamU1W54+qMT
1t18CPCe2UpJwsHhHHiIRa0UdDF1NaezGmLWWQHu7bdllfn0MIj6w7NNL2uDJfTZFaQmq3/0MA48
Ufc0UbTxv/xPbfg3d8aYdy+lbF9ha+cXpTUmMEkyaSzqisqsD4J+P1oA68IP1BFgQxc+a3K58cS0
VBUIrNKBRay4b0yMB959x4QyjxQzRLVFDSHi6fZO2IOiWH2GlJ2j6R4rEK1ovd2l5PiI04q3t2gH
69ETqEVAYxxP9dko81L1mLK16Ky7Sh8CMdLpdyg7hSYWaQ4B/4+8HqqxIDj13C757F11RaXkkKvF
SK3geOmCUfsLi/3eTzljWEivSF4i5CjtQsaEKHgNUd7z9RZeeMC+eUat9ePPOF/rGlbFC1Fz9sXA
ODf4vxxv8qi3dQWu9V6v6SdmBaBT5T2aDVOQT3mqMcvYJPm8TzJ0YjM3TWpxoICC6Lrij1AcQssG
vT7qKp3vO/sLEv2PuZehBYII2Fqv7mkWOk8NikfEpL5c2XNZ/51HNpKeUbNn+jaitO3BQKvpLIDy
lpH7nL8feseOX2CKWSBZ3Ur8y4FEDZVYjPn+EXLpxsRSxCdjO+23tMKgAmnw4slbLIIw3wiOJvUO
d7CZLAfNjTABvF8eEvVZ79GFjgn/h+Ee8oE9A6Qt7kcyIYV1cNuNkA+bCdCmBHRXk0RTg9hUQjAh
zL7VcMtp53fVOTF/hCtUrfWx2w6q6UyY9/KY4LNTVHwR04SNbAFK/PyeY/66twNpU3qG1i57FEl3
yFNLy+htnGlhRbvtgYWcxgVwe+DdH6mWrML8RC1OU9uWaIOVBircZcDyvebik4LIaJBw1mkP25zo
g9sqTirZ/iGYQVMqh5S9503yFeSKe2aBEraH5x78T+Zys5hYMVwvwu46IjhgMBH5Cyt3/kg+gdCR
B8LTypO26dG2GrTiDybnejnyOb+k2kPJW1V9OBL9RTL3ZgKovrSmm33fqTm/T9C0oJU7ifN7e8Ai
6qWE+9HG4fm7shtXqMSjUor9BFdEL0tgxzdL7p8p1GmTUjiFOrdMtAjKUgsSozKBUVh5NWXaqr2u
26bxEMzV5G8PDDxDSerLYh9dpgYk4y7J5WE1Dye8SjV+LGz6FK2R3lXbpmyZvpr0pHb9I4rM3588
lFqtwuxQZ1ac2UfgEcoIX7SVpQDo6p9hLcmbT+kH+txW+kEWm9YUT9y4O+D8etgbNB1K5JlKvGa7
rX8htmw9t8ScueYrogyVhTqW9YAaTq4w9Pi1qggUkk/8nw1n4wnXZX6neLUkXVqPBt+RXQm7H3z6
JED8dZO8JKQ+yfz335yp85Z1LNtXe9wc/SinxxRFHsLFUN891VcPFef8fxactqfxkw4aqIg0PwAn
fmOjyZb0KYjY9iv3IfrmTNjOgLKOnCviIY+dcxLbNaZ2mu8ec9Ba8s7SfffdqEwDRqEXX82lzVgU
Kgj81x9s/dxdPCuSRFVEJ0hPk5jB7Fk+opNF632fO4L8O7dxF7DFHp4GpBf9XkJOeatWwnr4gIPu
VPb5NDykNrjPaaw2FhyTi79Vkautc5CybSNzzQxuOsqsxcDls8VDpqQMZ2wPbsp8ZNVF1fZcTBCA
gGKdpXAR4Ux6Xqnj8eL5r5mCfZlPbiwtm3UFYCuPQVsuxws6taytxK1w2F0LGVbtDUR6rz7ZSn7z
Qobq6HX4xZ5VgOJn4RWVfCCX4ukMUd5nB740DGFSFNfOdHcA524zT5xQ+GizJaz3Kvmn48b0DetH
zdmJY1NNwOVUhiWD6IHM5Hjrka4ihrbzhjypDJ+6En9d7Lf6y3NDQEWY6a7adFw9j+Zn61kSVHlp
OrZ+UEAeK5bMUp1N9EeVGZ4ZOgk59qKP1uaT1UCUCCsm6EKSoNigXxU1oSDCya1OTBEhbrunUzot
vdlgd8pcJGCLuAqppHHn6/0AhyWyua6T8V7OQdswWhrTmqo1spC8NHj8cIDikVdse0FcRGCiRg+d
HmnsSv0RpNC5BQjbpZmBbUevQWe4vo8z9R8xeZDYp2T52A5QEQAD2JFZmvd1ejG2eM00Z964TVMJ
e+qwZD8Nc73ZipXV9DBfN0Cag1wJzeq9gr9ngKE/Za6WrkV3NBOsdZ7vqcqcxvZIi3yFdN6T1fu4
tIUTAeAWo83rh3f61mcPQUHAHgji/YSEAPKz2ml6G9/m4V7Jc5BMNl72NCKrowA2oI6p/+jtjuJ4
RzCfyHWow7hoPCMpnmlMZYlrPR0Ovyz0lnUbvL4N9Smr+Awy1WsNRWchW9iRzzuzF7eggI/Nzz5a
v8kh/p00/ofiFB/S3n5YOLP+rtEiY+W7lqnaI2T0QI6qjKbZitIhHwyGbnovoEWvXiC2aQoHWUSE
OrqHQRqWGypkXBInDtJkqBMP3X/oYDg1uy361OvE1EIw+rsXHw9twKoEEYGb2jWTMPQcG2MgXMQI
GsfpASftckkyy1NH+GN31yrHuq+RguyHfxs4Mpz+IluSypZXqY8POKRGdM8a3mqEwaT6jwjJAcIg
hL61LGkHKWbwsr6DMKjVxF0Bi3vpYU1nQTFXAzs7weib8nj55Kk8GxgimFbaObrO9vg465EqpXoI
Yueu1f02lNrP5M1L+hKlivBxhAGY3QxHmwv7wpXtZRpDclZngKqZRiXV99fgI5Y08P7TN1TOQAfp
qp3LOH013M74xxu89EzLOrjI/d6IB+k1fD5eT36NzMKRgWNuh4T3YW3ZI08EyAf9w6Dd7RSXh4PW
K3EhHTWCtwYu7nq84TEjPmQHaDsYZnvWRA33vaI2YsWTbXqYNcxVZi1plnyZF6+bA/QAuRvgnS06
KyKRdyhgUhKnN9SI4UFycd/kytwDXtYuT68vv99Saa9mKsyPDLxDJwRuoxMrtzU5uBfP87ADa169
xLlG4D/rGilhurT6qCbM40aUb9OralsKrgluK4i7zAsCXvqXY5OQW2zfEOPqJDvuwKQ9AffXBSfq
xNWg/8cgqkBEcGk2fcSGMNytWA70PU7U6q3zXtS3rcdlv01RAvjjX+zd3MMcZEWBEKyfT91Btg1B
gMN+I2x6ppos3xc94mvuNk1u2RqfZNaS8Y86f4OvaM8fLtvLlnPyDSxcOX/2/rrLc++ecGrSL2fo
qpcov0F/+5YvVm4hg3wgy7rQ4nFEke+e2d5wZrqCdnVxO8k7mTabQWl7TwW/BGkxYoLbOZ1g+znA
HflkqN+QGcWh3d2w3RuzvtkE7iieNMVHNL8ZaG7sy5BOIvMg2m8F7DF+fTm73sEUAOBMFvf/EJ2u
NEUX7Jq1uN69zMP1j28v1pgZMdiHcJaH0KoqwZaWd9xfV7wAOtj2UjJ1ue9y6LF8MJFInPq+htDS
Q1gIrGMCeOd4S8bKVuTxOay9j4Q4Yf2TOTM3mfRYdoz9N4JKMT+HVAaUBlfDDrioi7vZefco78/E
QeMvWjMAsD9HisHhiwjtrvD+Pd8jDq5OVt+LUrhBpKCCvJVz1ZMDLnyf9j8HyVoEQgjfQgXMkNb0
hAMfOBg47ilQ23mQbohzhVrTTeAdiMGirn9vSUVue4qHIhLkuuchyIrEYkEYkSk8ggfqSj0vMJiV
ijWrog6uHEDLtHpp9y6R2c8s9nszsgO0HKe2jNlkB1R4FeQN+KHt0W1zcmHh+HP17nUfEqOevdFv
aUXioZ61UVxRM3pla10kGt3xsMhY+iKGBlLXQPZ76/AP5ksA55CsEjs2YNizCfMd6T9tcRN8Lqae
p+OtJhBFEH6sHff1eZ5FFlyWF7BAPLxXZuULK4fZgzcKK6JLKe1ztuFUFbQaSVqziLVIuevaa3EL
aT7l5/uyR9oREU4Q4ZX1/GVrByI/Uwb+HA/k9HXF1cufloCBnyGEpOwhFyD58voMCBP834Wgimpa
qWWYWppzmGjl8mO5vIRxMkY4Bv94zYXjvYdMT1Gszsi0YZjI05TPDqnjdwLSSwx94E+aj12/KmRM
WaIKpqZPs7wxjnduombp5itKxFSUvIDmlZsbZtKwrBjd6IDnEtsX52yz9o9Yy+VRr4fkGVMW44eF
LVU1R4sfIVzqf6t/Ippjju0AUlAAPnM6XD8p/oGYncYuOQDjTxwh9XXTCvjAZHqfdmc7TD7EY4ki
hf/fbrKIq5nhoAyxNGgXg4PZg66izZFIb6tO891vsoyUOB0m+u4lm1RUZ92FExvH7MXYxdK/X1v6
tzue+h1CPrJKbD3w24SN/gadlNQ1sGGISKjc3rD9eFzmwliUA7BlJM59AzRDmBmSWupfC9lNXSSO
3PWOdzBPieie6huEzvQnnjF6ddEqtzeE3cWz7MxDt/mvbpYpT4nDL+vnkHjkzwb68jP0Qdb9oUcL
vJVxjvB8JIfNzVUeZS8URvhaufRX9CtS10d91dyCizUACfc5QxDeSYx8mNvheflHbkprlRmxT5Qz
eA7EJQWqZZP1xBK8gEvFut5AlNbF1T5dtyzjrrythKLxLBksXlt4sNPXzQ6iBxkwrOj6i4t3w96+
/jvXdVVrCzy+Axg5XII+5XcLI/W0dr1EdhABr/q1mQBgMmRzy+Ral4RG/EchokIa7EZ7wgdaiaWr
USQ/8+mxsrmaKXk8kfOZyzbdqKcReNHLug0SVM3H/paFm7cILpmNRmYg19kdCC9V8NK5h+ihsFAL
gfBdeZO7AaZQLqjnKR8JUBK50vS4Pc+H54DFamADwR7pkV4r0OA9vNbhjReN3uKZyGdMX+undejV
sPtAvpFKHOCvdAzn0kFNaZ3loYz9tvWaCg/TVcZVzkhFFdX3jzxq0H6bQDnch/Nv1hDxVQAbIYcN
zXa3ewsMcuPsif2IOOVIAtHTkO+k2CJWMq0qHZasm5A4v0XgqzJLhgZ2t1/IOdA8buzJiJ5nu5UO
h/uMKpX1FGPXfWlt5WuHWTWEStGCMbr67ax6M/jJ8Nhi/WVeqN7mGCMVSbLAZBYA46U1A3rZXw4n
lQlf/4emlg9QBJIIQQ50KvwxA1hED0qC3z7KBK/eOkQw6Osfb3VlL159B6qOox946qeB08BOr4mu
cvJHS86a0nC1xBnDVOc=
`protect end_protected
