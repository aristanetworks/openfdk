--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
gl/dnTDiXf/9nXPysqHdsVGfAHLqgSUvBpV39MCRkQ9VbNgB6KPg/JjAcr3RDY7yPfralhe4fPRb
7FgakvoQ5whbF73E/7rBNKTQd5CSWi/6jBPyo5hETb7zTKJ7rr8bsIlSbJkBFIaRQc1K+FdBEHcm
iMOtafi/EW8PyI3k+GWe7WSqHejEbh3sruSL1NxZ7RV9S498riWMnKtgYrYSbH1c+eeUwJOiCRL+
1b/ZWViNcPC4vtEuq7/+m+7aZKJcvFvfM+XAnOfhX00s/JDL0SfCPape0OGku+dmSFU2/P3ThOhR
6VWxYd36EOe7AGLLzn4g5dlen++sMxUQkh4yQw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Oq7WPtkQFe+X4HBn6vtYYOxrQtJuBx0rkNkmXTcDOME="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
ciEaJq4bgXJNKHHE/INnF5VyuIDRQfyHWoAvb1s0jQoV2DDEfxamh8S/Jil8na97l8e6oiY3hq45
3M27OJHFpFd2Pwi+n4CiznAu7ano6un1IQklMMSl9kpmGbTS2qUU1fMBFMbduQ2Su4M0P5Zh/uSu
8W8nlRF2TnrcY69xQwcnHxCOFGKXxtT+T6Sui9O73Owb8YOWbDzcT5lv4GXlntqMtC/B7IlF7j5i
XK/c/Zq/ZXGld46qBavjfu/R+TQk84FyIle4UPjaiRMzKlizQ51h23xtfhWrGKnNyxmjXNMQE/Fb
7xOzZSBV7X/o4xQGLDj6YaPJSIj0F2S9/fMZ3w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="GsLTeoVDPNuw1+EigULu0tHAEd6xggLlAp7bBIIB52M="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6608)
`protect data_block
tvgBqvHKeOaEqnnC0p7bTR9gisqu2GrB5vNHZOzmfyzbj2uSszrl4oTGHDvCdBO6RWr83NinddvU
QKPLx1dCuNLLo9irW2UiCW5z68RW4kFzc0kYSQ+cUXToHh1vgRs1zhHKPJdbR3tQfuC+OrvumpJ7
PDcY/m5lT8iJgF0/eVxM9uHg88Nu3ZWbCP4KZPed/f5+ua0ELULxX5Kfpxdsiai+VSDrqJab9Xjx
Eu6Cl7qrLWlQWW8I2Vn+3xse9najHS9conhgvVz/jIyCABY370+Isz0Ry6jBzRAVu0gqTnco7/8W
qoVyEwJgrD2WIQSH1bGbtmxVjp0WYvMqERkygsm+mPKDpAu8X5AkZvndEllaa//LiqV9YHlq0u0s
bYiuFN7KI7hMBWim4bagt5dO3dAXo8S3GHZNEAehNocYyiE/6G3Zjt2Xvb+U6Jt867BfjLzBHw9/
l7b0sudvaTQYMNkwWuFHVp0TGOk04SQghuFlr9E8qJWKdvBbddKsBU+/vq9rs8HmgJjosp5DYUxl
SMTYElaY45MJEpTKBE2Bwwo02GfPMT683HxnYXRnuYDYtu3jrWBXJhHdf+st4S5aQVcpxMTyOd9n
vM16xVDsStNwQV1Twwm5DtpfPpRLLgxUQFk5wsUGG/zJS0Eizz+TblU5aegJNWDhfiIwuEjxNL/Z
YY3gk8yWDwA+nkADhYwEC1269Rf7B4z0EJOJRzlz6t4SYJOsNxxzqHybRi714aBD6tCUYkEhWJcf
PKsGfS5pNo2fqTDanhrQBzsh8c4VaCm+um+LyEHFSea9aZHlykKOt4jQd7WYzBfMZxaCJgqM9Wed
MsFItyPiXoQbybTnDaS69bdeISb7sgGKx9gSDnZtboyVOXNfbgJQUMlgbVkx5NuSVd992kAvoyXS
cZRXXsDAtEb4/gWzG7gOZOwmS4fBdL08uPp8dcC30KqEtaA/th/0SF+kz4S4fu3dHimWy7rZTGXI
03Hr27sFCvYE/JzheM/4x6eOohCH1KmnmLtvYVTUl+LiovKXR3HnAFeXH8glSuSHSWZ7vtUj3wIB
3K0Y+SvId0ErkTdsKrKFOPpMgiVstYyOKAt2AGjkQ+ZjjrCuxtNOzuowHi3Ah2/ldWh2oOy4HMkH
WJlwJJn/gI6lJcGxUdCut+H3t2Qj7hG4FINOeSr3eRBBW/vd2YhryBUZ4zfT1GPC/YS1nQ7fXFWc
ThkPMilOo+gOqtUbm1e5RstI1OkriXyGy87WBBYU8821qy6Z3Tjxl87lOr1aopAF5pyRC5znSteF
yTdOcc5C94o/CrR6WlrAcKC69aVQECxUsZEdQa0Q4qBnj1kUnboswU/xAXAq8GY8BPDYvkQEFR12
t4549SJJVLEBHN5X1ml2lUzWKeOGtuXlQzrMpltHErOOvnJLhYjOeb3attY/kqG74jpTfLWxPve2
QIqaq/nqeT5nAgVZxzaHSnRaG5Sv9CHB6noK8omwWYUfowhmLdbz3y6vdQ3RPdtcpUB54M11gNkM
fXuZ7szLkRrOqXw8mo3Ti5LYYg0DOi020lTjN8+YazqzeQY0tTmL0nhco/j+b9pVfdXiWYl28i+J
zMLomF7EWQJ6LJJcqPtCbCdh7pRGMmDU1LwBN32qVVXLgVHAeZElCn+gzc+DYRyV+1Q8kH6h2F9m
tX31Yq6y6AShus0nFVduoQAyZi7/vyWxyoyyUueVeqCxC91x6/GFGCmn+MTIJtCppQuIQBaheh1F
qSVeA4//GdZlpNm8t5FnYzEltW+KeGAzfcz5NGGY8A0MhW7hoJpQZ/wptyN9rh+q25K8wdIKXd1Q
BDu1ReHXw7agYgxot/BNl7lPa00RECfyoFncEOViW7DVscdbjnA1UIyrGYoF0/0ROF0sOgYa0rDO
+1YxxJizfR107H8lhWEeN4wkYvFSwMYR7QyGwu3GFJl+5BKiV52u5+i2a/bTmPywrHSvsqCkE+Wt
ZJSnod/rN9+Whx43ndk6zZ2wMXwXNt+vHbmY3cX1TM/gvmlIWKUpFLb4weTqSRDLtqCdQhXbkS/X
TB8CIb/eBYryL12Il5xE0aVfp+U3eDVT6lbudPI5omzBCtaNq1dSLcPfPblmNVlnIKGL5X0Pv3vv
k26Pw3iX8cFtu5nr/An0lxuZYPjJMfyxqsWRz2NA0R5LtVd/nUkKV1RJ1hG0vBOj8yn5mmOoCQgP
/+PFlxxgxUU9jOtYA0nYXEWlaXmtoSsFfNQgPpSEr14sflq2/tu35N2A5f2Erylid9z2lFiolI0Y
qf5KxTNFatt2w1Tp+r6hWeSMyhz1EfrVllkI7uJ9STTRxWu7DBxNEgDRkQACwHdM+lph4htSJxiJ
6q/futNSjMCmDlVVswtKCM8vhrB4Kqfm2AgliMX767BvaPKhXURwpEQbq93LHQehzMIv/Yzr7eyH
Fpa6VfT7Ry/bYM5gHWlYX16Gc+ZuHbMYgCQZqclyNVop5MuOI0EVXZkDekm/hdRll9+d2syRd7vP
hhiBZs2Zbz/GT2iJyow1NVspAFDuDhCpskDrgnypXVKAzEo6D5CZLSTcxdhvs11inVsNn1i6BfGy
G5m3gOQVZJUQcfoU0cEyu/eX/Fgyl5uL6dPtPzFEiwEplIFv9IMDDACWY10paqKK4RO5w2hxt/Ij
K86mNN7u/eE0u+0iFRhBhitDusWuSdxVxMuZIy4qyU/Xgja0RkNmOxjWDjeMfVxsgOQ4o8Q/JrTX
7UJvJ8OfF595Niz4c4FemzfE46g6mYJCZsTf9UAwW9KqrwvfFHQYJj1Jvi3//nMQ2gYdxL6RaTgQ
LGX2dzYmQy2yM/RxhRsIQYgx0SeR3WJ0+l1h6xAZK8zq88D4QYR+wiPnLAM4QrhUGlb1X/N3BR6g
qr+aHwhgDmW366u7BTYvZicsQ6cy832CXbiEXcoDc4OoT+8/J12KGCIxyc2idVEhB4aAIROWJlsi
v8y9td1h3OjWzBzO2deTBlR0rTNG5WkS0/X2/l+sHafbPbwQu/+XmNmHmR5GWMx2WkA15OUN7afs
dz7HbzETozhkYag86qhxeIKqMxnNvVNSwCz5D9YW9J1f5kaRpuf+QGjGarKKAVAakNHpBij7zevO
o4kw8N9+7Iw287Jk7PYVsQJnnYAJBcqkYurTZak3F5SfQ/0yZOpF7feB32BgeS8y1HqqgPdZk5V/
wS14/0AfCKImH7aOVdtA1Cogr6YSx0wSmiiVn28qq/LlAzhqmYDtsARFVCQ9lU84rbcmfH4qRqpk
yt5Rb0oYWK23z870V4h/r7xqLTcNYmQ/i4t4i3m2y5DZT/oB49nflcf351SDd4LkmJmMOGZorq1L
IQO4HETmx1kLQVEsmXa88pksjZqPKX0K4fJAXqUNVnz1atIH8tZ73M3jDJ2v9s8EkqKa63mW8Epq
7DS9SX+4a7x2kSlV6g0jfh7VfOXBa6fAvElO0YvfH9rIxqTCAM2JFdAqJP1d9O7MzkkYuexaGOJq
wQcQ5QKHojJVwF2gA7ZTNLLT9sPTA94PSpmJ7guDM2nNnjLNKYstInDyPF4nA++BopYsu1KMNtNE
gnhrVmodcqY0nP/iRR0LJzQ2RmWj6e4Hr4kAYnDDkPodEnyjlOQAL+laW+AgjkK9lfXqg46lWmPQ
RU0GqeYlrEV1I/df+Mb+9VmAV9nxq/x1yCvUSbLPnkQnx8ixid7YctVMzZdNOKAYDxMXmK70KxOH
TifuJ5nlJ+tQoxJfIAd3Fvwx1py7LyGSmcP87gQes10EadMBnoOYdLG6E10inCbG7AwqOSF5tugH
EOeHVzIqIkAzSRyU/GKt2DNbrmRLxAqDRYGr4Ds7mkZ3Syn+/zrfUMrAIZKm7FTPGoV5CLqJTRVy
hNjKo2ivd3qfYC/YBo0F35sfqilLrqPp9dwC9lOxPyZ7CuwHfbOsEhuawZ2PPleWoRrhM+kFecJn
wUhheT/+lDXgMLMPYmpQnsiEMimhEGT1seAeFdb2+xa1oKWRTj2AFLE/qebG+HpD8PirbKh3YITm
eki4FmYNLPaPzJI3Tfg37xSVwYfp1mqq7mngMbBCB3zflVC6oBw5xoEHT8zvwUMbA7bscZ8QSgUd
Bn6Al9mcC9ZS5pJ3fXzLIp9ZiGTzeOnxfwtXHif3u1ypPqdVlQpnqbzBhfwRSqVM9KWv3BFzklru
2FZr54pAt11Sz59VTFAOpWF/gRVJJ2Uzr4lMy4A5Kwg7eYTni+8Dlgq7UYF+tnywU5qRvVyUG23Y
VpiWo5vfOgcDZwBRR6k4PnCo6x/2FDVz2xZslxloS0iNpAUufKNoSHVEvobpmto5FI4onE6Vzz4j
EhMT8E4yat31x/AbDVYWV5xlHPx6RQt06EkccFhg0pBTGCeNj2cBgy/XBzgGsDIqyjSiSFbRe1B6
/7X87iENtZpK9Vyz7pi3GHUE7idhBnYyq9lRB0tftOKfm2lEffEhMFQC0AXicd7kgi4yCNx62UoN
Y8N3uk4YUwXDJY2p5gqTfTLFSZxK7wU1JbS35JoPt9/5LaRUUPYkC4dTJlmIEdaBnee0gbnzdfHl
fZxkhKojFPzwZczg+BjhOJZ1WgTzWEzMMCwMUsDCiMaS76uQQrfaMJ6HkAUfSJPw+N4HK1HlkSFh
saR/sE1vh780Bc3bFChoZuyARzMQtYZUrmkYXJWc/gF0H/hkpCYHpL8TIt+D9p60gBVXv/RjEcRV
EW/NQ7dZo60WbPNYD8vnHQE0Xk/vE3QDJYgGaU9VMjwJS9PRHBxEtjylVNg2QsaS5xzg08nXSjir
u8d9OF/pANTvQ0KlEs0gEgqKzuS1GkZVr9EnfDakmerPhQ8LgZO81slWJKDdFPE4mofVYn8lulgn
/tJhmYT4COrnDPKbvHZJ8Bsjs3uozqB/ETUhtL70GCMMX1ucVqF+gzKz365lpCAgZXb+Ua2CeWz3
E8QTMO4JfK+6nyxa0F0x6hH1mS66dxQOHnbKIifeioHrthbKqVyHFLyXKgupBcH3U29/7OlWLIli
pQMwWyxchNVapuMiB+P3WgE98/NMwe1QHx5r2uQshcMUSuufzbPerPiMlHQBypXQSAy2noLlwtKT
X5PHsccKhphAFhkoGkrTIaLUyTXJpJv9lB1c+9YWxUVqHpKyoSl3tQZYEBOt6ns4AWkMPY5QFrjf
BlRPH9NQUKbH4KeseiVehFhOlzvfEuqJBW5ixvKDqeZsjM6456e1wLgFwhKbw/EsVallRGod8UQp
YajU90htahVB4ywfNm6XMg3cmmJS8EqD1Ay2oMSr+xQ1CJaAPapeCZ+pnN0DfBRazXlbekchI1DJ
DnqExzZyNfuw83OY1jmiPg2Gbb2UMj0ClFXRG3V+XoMztmMG3w3OliPOW+OlYbi9oKpG8QxPPI6y
0lvcVe6b9GP88+GLPl2VqLe8md8w4LDIuPNj/LE5N8MXb/gg3Oe+ZJP/HmpK8Nb1buF7FfW7Ezmr
XNDMIIK914vAZVM0M94fC0KyVH8UVld7xgvy578AmQgLF7BfIMdtnopQg0n+NBHDUH8pvYLf67e7
kie8okKpaAgvevebSXOZ7RL34GrWfjXS6XyNRrw90gEOrRCu15saunrcIqkijHDWdF6n5SPj8vVY
i0I5T/TAkA6IeMjrDWohXfstdNXtJMx6Rfc6/sjVn87EWqzbXBuv08tXL8sjkyS6J7Ni5RxGiLtu
cX9+Jz1aql/oq1C4APctVmkjsQT/8u097fYVmek3uwsEm0bTaJRl82NjalXo6gyc8/E9nlWtT+zp
gKhxnT9bvDGCLvmoPEWQ5g4Ws8RYP5gAv3BuY5QRB2IsouWU93uU5JrmkvwgEuaYhKeFXl7hwE8a
R4JUfidI9V+/VX0OZh0rVWrawfl1+8T4FRDSVQZZDAY7Nw9X0yqUZ5X8+GnK4DKV2/4AdLQejrJ9
K+egLuJvpMfdvwU6hoisxs1We2n4CxYJNqyZbicex0wMf42JzK4GlOOyfMoT0DsK6leDgL+hOSB5
t3wHSz+BcCeiYWnwbmEQ8rIf14EnPd4w6s6PMmptUmzZCzUlF3o42+5PqmOsKKUsRfhCCXI4eLRv
McoN/sSJI9Qz7G5qnnb/9QLg68HjonNpSZZawz0oY2vkcgOSDStT1ooK3P6oeXIxSGrG5gSZo+yK
48TgC9yju7vFA82eHhphspt/A8qLcNG2+k+pNl9PnHlcU12m/WGsRf73/v+Xijhq8ti+ny4N6jS6
8jZcge5HXqO9syhjgLUUZJ4gQQTu1wiFBxlO7KeYh1dLxwFHE1ilXNpBqzXQpDRYgofchhTF6ztA
hymc8lZ8e3DjWCFM0jV36O7vjMDkn3dtC4WvXVSTfnaTD7F0/gmdrvOmJtHcO6W+mRlk0xC86Vvb
pOFAbXHWgCevKm2nu08qTIFeMjxTiEnUbPN3ZDPODXS34itdAUdUIsuKG8xpfC2OlJOzZ+r0BG6k
vZeoIvqPjZnTim0T9ZykThJ5rnkZbmjmZqNi5ofEHDIfi51CedwrwLq5xw6HY4dI2biF7V4Twmda
ITwtVhP4Bp+rjxOUe96TRyhMbr0BjpgD/IM2ozxJwDQJfpUwso5e9ISz+SOMPkPNkt8HABxoxdxw
VvkDO+Mvkhp8XwLvNnkSR60TMaoU+BTsURZBQSmSwzubWjywTRa1OcnFCB+HFtq+Sxr0qM3cqN/9
GPUWWA3QlZ4EQAnRsTeBdAFTKLc2whWez2Fbfj7LTaEztOrszyt+QTtFuatvhBY254CzzZSlfXOQ
wlDyNr67B/0YLHYysI/RXn4bue45GEuifP8ac5DgnjoH7N861LKdlGWl2KSb/MtBJRerNCN7MFFD
/jmIIJjQTUVnyKY/IlbdPAfwqw6n28hrS7b4UI9fJlunmv1WM7pHNrnHCTatY79Ohz+ewUh81gmR
KVtBaKLVbxVjysge30cj8FtG9ZKOw9T+WIHVGMZwXR2r4kXeZ6aiT3UpO0uvN0qT45NANDP4M6ax
2eZDMRIeAYwb6MfvlwrysHq1H6g1taO/nt5BiA/2/HPADZoOfhAU6KjvjwBPgTFLFZZveBpPWtP+
IQ/Xr8KA3tn8G82h9ek16lzHHDMIZiuWIv+MlltkgvJUDPIIomdSQLSvTxiq7kLv6wyXtDCwTwts
l0MLfq2HLFs99A45hitF3AiDBTm+oo55IzmzA/dNdH68VNFmYGnX4H1NKgC8+zKOxJeQPz3QfTfV
b650S5ipiX2OCLN2UbnvR6o+TqSS6mG1C1TqdDAdYLcZP2+Yl33lizWw2L9Bx8F2v/R5TnDX4mcE
ZrOVkBY86vWJW0r8hOB5hyf9fzFw6qgBuqNCwGJfUdE+La1w+lmXcy6HL2i0vedbJ5ngOtnpabx5
20q4mKjjwKJMJL5lzCr4L0jLOychn/2El+h490tL5IlqWuWeq0zb/3BM5STftFEkSeqGcriMlihL
XQlweQmlAMv6JWE8jvbUkGhOeh4gJD6joSIw9ivujqssyAjVJE7AdLhS/ntmh4fo7u/WDCNLQpXl
f6Lz9HjjBLa0cd7453Exs4vgSJB01UlTKGgOgQNShSvBJ9hDHDGbCyICCDkdDb/Hr6wISGvUwIiS
1TQp/w/lznz+aTpKjY8QtE7sBWDS8WsuOf/DnU6wGHAZ4L6fcymemo2e1U7MPupwyB1vo0DKJI1J
lO2NTx6pkYD4t1W6Ub4WnKc8WfhDrkjlDFhY24D/eTJd+842GYBNggARc7iXv2Mheuoj/4Cbkyzg
+8LYycPMAwe+pCeeZhFhsSC8PFfwFmgupfluYuW03OHhb87L6pX2yrPOFTWv7fNw6TZbj31Csd72
rvQIzJ2DslUhVX0OBd2lRRmk/pcg/ie+zlZkIVUrwHz2fuLg4rnGpVk1S96L416ZAs0wotinmL6z
dBl2fppOqFiDTARUSnAKNLt6/amMTj+sgW4eyiTdexRM3BpGXScC0xVeg8yZ//Z8sBp5j8keyKp8
qZvx1sMdoHcQdb+I3btMafKc1AUfTkuB4KOyJY1medx+B6efpRIvsNm2GyzUN4HpsFLMsZQls6cK
OA/PivDORCDzeOwKXg7QUoWNzgM22HhT3ABs1GwatKCW0xCpKLfytetWwUyAS9dfgJYDPTlVfMLp
xWMCECzAnwg0fRgF7jqE3rDbVqYKH61IMJAyoxgSqyA7elcJA1oNfK1xzA6ATBwermQYzaL9nywy
kL8dmdp+2nlWFK5xU0mvNIIeJsPylduDf37M4K3h8hRbHSWlJ5n06dzJJhc+rCRX1o0bsA23g2RS
Nccw2OOOKELFIarkpHkZbWh40IhgTeMfRPAnfNUx5a22eVmsPY2ZDgzJ3ff8WyV/lHxOx4VcJTT0
nvXvHJyEBCcBwkS5TKQ3JGl6fTGylcGMvBuGAieVGDosz+r2RsM/Fsg6nPDrmypvHFA11NCqYI7c
wb7YPgdPEMSK9YfvVE8W53LtXgGOweU5D7hVKrexkczo6vZmCyJiJ4hDpGsTRQUhOR1qWNCfcK5C
Z7eVJWhn7OaRS0Jg2TI+/RHS2zhfvlV8dXasvlDcxkomBevtQ8ibQqyZfHU9W1gUkZOvwvYZWExb
8YdiaVQM8tKYaWsbaOv7ZTPJ2T7D8WSPBu5TqUrnv3lraakgOs8Q+7qE0kn+z/5go/9f1s60jGEs
mz1w9bEaondxTk4Kami8rG7EqymE3w55oduWW5jr9dgBU6D8dcM08KeQalWoZ0oUUzJRE3YkvENM
NHJyxgkEykxGC5FIxAgFrQFrN1vJM4CIFAWk+EWCGPU40dPIBlKymvC5gxUSA39IsIRTaDA=
`protect end_protected
