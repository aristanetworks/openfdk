--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
lLmHio+/v8TfZVBhMTFRmfk0c5XiDtXTI4j51AQ6mmXIBKC1K5jv40fZb6ekxIM/gp+TPiplmofX
6Cd0yfEGVn2kkR31eO+nQJH0tqQgE515MT9KaqPbm62nLUupuTUElnGdluD1d1XohES1rrgTjMKj
/xfsBOCrXW/D2IK4FGPb0fa7weEkIJ1Ad8/SimkmceW9LAWWQLxPdRcWwKLDZZti5vGx79+fwVA9
2VGC0MWTU6ltdHRKzJsm5LLKQeB2gSBcu2Tev4p+ARlH6j8/QvZxbCED0ddugfiMYZAAghEmhTIT
xr3Xbyl18vV22wkcLGUFGcETphIvotCsTBi1Qg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="tqEjh6Sme9x0TAWxONfBjAiOl+u0kDVI47xQg3HZ0nk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
d7Bmwhuc7nuS5ObTJEwV3VKNES2LoQTQurSatWTfFWDnWNUnBFH2JgJ0PmYT9Arm1AXzDg3B0M18
JCwd900YGxL/otQACnH11+VlWe6E8lQu/sKSLQXloMrE9NZV1Y0fYzxieDxEgqPRhPfsK3jtC3IJ
f3AoXSZ+q6LA+cLFHUCN2m3lLgIa983Wknf0rP27mKCAbBNoGn1qZ4zRCE5VpX5P7Ae9eYsQblQU
4htHKIfhTlUjXaDxMTAASf9ZvYCcoUqouWhFerCLWt8OxCAqoHROmG8p3PITBoHR9UhfSsbK0fLC
xZ3V2mlmEAl0yfn1etJ/kyJJDsgTNOGvPJ3kGQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="tjfCI9R20KhOcHScPWQ2v+NtLBchv1Xj9UflQr2CTgk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3888)
`protect data_block
cU6WE/W72pV4yl9gnbfIIW+0iiG0NzToPsk/tI06JHoKXpQL3vSncpz0E1jrkJQuAs+GJZoSL0Vc
BCvHfqSIKekNw56KP5TlI6kyuAwASEvL23bMSlfmk+6EEeiP2OK1RZiYKKWxwcNvdq2S04dOWQM7
3gMXofRqBQIsWPFx/kvLFEJnrGDvKnZ7PLBG+hMGekoM1M/mRNVyWWuvNPuG3oaZFV4p8Et3jZkx
9iW+jGnl7xiRpxPYO5j9PlfiJ4/LjBqyHNxaH2qudDQUVa5T6FC5SCnH6nysEFjKvFgXYOtIdMAF
w4P5ZwBmTiAKgYmSX8swvi8C5tU7hwmEQcPj8dyZRv44Lyxg5XXJworv070OpjgME4Gdjrdu4j6z
OskrnVROcIDxdQbLYlyYq/Z7DsRwTWYDboqK4ngamiqi/cNtP5FzZtD1CCk2roQsY4k4p6glAlNr
vNwGJoW/3quxsX//hnsDuBKdGsPk8/CfDd9s934aCe73LKnx9QfkfOXyensprGlD4BiU2hJv9xqe
4pWIRvKOkoGV8NIZ2GZ0htS8rwHQHeQHqvfQJwP+Z4zMxRQsIvt4Q8NGT+i1LrM3K8qt6RPcTaQu
wb4Qrnw1J5/uZm++yKcia88MdBM03Y6hkh7UJaXxaefx4YQ03KbDDtsdyCEmCIFLVHU3kerTB69s
g5MM0cgBbLw8jbTHwchGPPtF/b0gldGjpz+yFbLDvu5b7YMiYijQaVIrYTmGiJC9s2/YUIzJUVSE
3puZIS9uArYSgZDQSQJscp6nl5p06w2x4OGYxSta9FmnFrcqnpqrb8wMZXzB4la1bMy58O/BAaZY
Tl1nyW/6ae36O00Xo2hsK2sNLYmlIbspNb+m218D6GP/SsIoju0uQ4IjhZb39INz3zIxzo2A2fcz
o5VQ40YtReb89hU5j896O+1LprHfiVrr3HIv1hnDO0HT18Eb3CTBkEf0/7rezc3N4IJqqEGPPTb1
UYZp6ZX6ZpnU/fNOp1TeedPjWc7p+ZMPlwFK9oYxbdZVJhi0dNnYFT1RP98/WAgU73UGLOrguvmT
yjmATtqVaHBiVDRXhiu/WIPgidv+GjeebA+UASObARyzWkMA7hZy6TvJVn32hQnaZj5oy8m76x7T
tsgggjUmHi1D7WLZB29neh/jNmp3GIJm6Z3Lo9jND7PK/RZtDyEO4zw5R2ILML+PsxQ62xalhHFP
YCQHAwioinPyB5Wo6lO9q1OzGuLVQnFmQQsbKMT28lPFsxstS4E5oy9wR1FCvkansc9K+2mLwZCK
KB1u+NNs2tYBDsOD6+l5wpUmwBVvNDomq2LSbC9KKR1A57OK9lWwQeP3VsZwzwKuIQ+gAHeeHI4O
s3QVxioYSIBSwLtL7cYQ3sxDmK0O1Gp8AXGUYtFfx+aY95ISa96FBopNiuK5dzhsiErq8PCEWlew
GPiJRhHy7dm+3RZIuPiuQ3BQr0I+lewxZdGFDdK52kz8fhY5JDpvLnKOoEnhMHvcI1DyWrbxTo4c
CpXilOWEeU2j3rUB36b7fNvhS/gGZYGt713T0byHaV8WLHt7hnRUwwoUPQ6G7By3jciH7cwiwwXk
dee9Lu2+KCo85crIO6u60vtnzEK2h+Y0rKzF+InzUokxQWLyffNrxEBetZtaamY0+laQgi4QAuMK
33SnD5s1v4CngzYgni4Q/iG3n68clZDZsRVpd8C3HqeCSLekvtObtv6a4fSwrVnL2ortqKU2ZX/x
VS3yllN8+vWs0A/yExgxp7Yg1o5pvbboi1KOICbSl2TJFX4SXJEWarliP/NS58c8gc84FBuXDTrm
0B04V+ZDqA/VsUngFkPq6uDWidrhNQfRWE27rQ4ydvTKiDqQILFFTaiLrusfbJBOJ2GywuMeA120
QR9BCzBSdV3OliRbp1LUVqXsOeNxts7+qjhzGW2agfWAL9/TSPzAin4Ni6faCYB3ENPo9WtmeN84
zgZ8mXJtBm+DFf4Qsq1IKYJ+1QW2PeqmeXD5WLOTIcPIC2C4vpkd4iqux68zI2u/YH/XvcEDiaRY
VZK7AvW21ckgou46td5faNLcbha32U6ZDMALdfrb5e7D159P9zup9Lq+f2ysBUvoUO/TSupPHnoy
tKBjNHPpL9Z4l5R8IzU6Lno06ysRAmG81+X4dxBtYlvD1lTigoxJZeWIyHetxtNLKESNHKQcbdve
E/z/FHy7dkwkfkfpjSLL/VHFbYReerIsyZa0R5ONoQu5jAUKnLIik5a70I/iTpINqKGJF4jqeB4w
04QW5gzZVGczfgYgA0Z+iSrko65Y3nGfLyaONB+HZ/VO70+FPoZzHOOEH05e4x5LzT4YOL0iIe9+
GL0ZimjGgavAyOQEMoJcuDEAmnVDPZkVD36IhdvkmEJBKLOzY/6OV3oDImV7C8GPsX1TzOrTzgZu
wqyNs0QoBSrBYFfj6g0Bwplwk+h1XVpHQzZAlaQ3tapiuhaOPa2XOuynry9pUpNG81NfL0xrEgJq
M7NUvxbSNrrRr0MG2HEScmNODPemRRMlt2PIswjHoRiOQpVTOayk0KZKQJuorpjLt00APTWuwrgR
vQfjQj1he1c/xP4o3lltes4+GxhlS3wjVF0415CtJ7e3Er7cOLeDJgkr9LogE6aM+MllfTfFkfxq
IGpfXDD6zIXzI6UPgbOA9DcCHatdMDMIOLf3vAU4fZPi9HYQkyX5nECu0tdXipCyfSUju4u0zZlL
xyQ5483+lhX9qxTYrQ3qs9JEhU6luTq/Yvxy1a2TCNJGLl9FVC4DtKvVpGSVpGLvAxYu7qeLYyMr
piR0FdI34eLguWm7KAcfk9YW+donX8usimcbt9Pm2fkkn4rF0DBz95gm7vR3fcXGrLb1j8Kdf/6J
UxrXTYxTokhabz2fR1ceV7ct6EpQODoP4DcCrK79NPgSsCO+RLn+fRfVgLVDb0hwB2e7nKAZRld+
0nlfjJ4khP+9Df0MkFgVOoWfmXmv4yIcsrMCA4ywiA0SJ3uwr81cItgCytt8ZVpRIzbS1DOc/hC8
JcqB15U5NliBOhif8bvoqUBLXZfsZCXvs9LzQyHZTGdKqi6jpuk+NOdVK5K8FEqRQGB9xpA41wqG
nV0WOd35ZJIiwztN5qe55+KzxmtlIf1QhWVR63QWjFnbtLrnsQ/K7X9TaruUmQptqFFx+t6qKZ7O
ubtAYGNh1sg9LoCxE1NxSpPoTaca6Gqk7CsrI7EyZP6yxe4GelmbakOLHWjhoxdhIuPSN37ZZmym
hI9SigvodN8H6WM6dawzfRpT4KpuZG3LCkwghji9QB4vAuv1xUCBz9rfwK5drAzOjgIIn16LKlhk
ujg/xMfwEceabBHLMA+zI9VZrM7Je4wTmDrdnejcPb4ug+brkXy2V+fCiYrwXqOZRkJwlgzYr1Fk
4f83pWhnt4mHupuWhfmiyZc35kn2MgYARuGdvF0huVscrQPuMvAmmq6NvejMpFAzoZC1awCnD26p
LlrMqknQl6an1JvLkY53nh7/fzy1aTK3+p1tTLYs5frnfwDVGW4EuqTjylBmBCKu0GqOlRjnSkJ3
CZG3TtF25InpHmsTpWyCo8QPYU3UItvk99B+rzAT7MD2BeGVoZBXWm+bDhkBxrV01+56IUFbdE80
DJjq5vMTiRXDDJs0mgd/isRBbYrPSvusqnGUaMIU1mYaqokTnKsWbwFT6lwzgVSq9VGCOT2bCWkT
7hOYly24+rVtRynOxsQEXQB3iiw7lRGGg7NrCtWmwJ4zHDJhwP2Hqfj2SR0Bivo1/Ww199AtEeSb
rkGrLM6gYKDUmdjFzoEZ0TsoQjhtdxdN/DCiXyfrRWSXNTc1f6lEVCf+6OwKIMtmbWB905AyJKFh
ccuwY6iDs/gVvmhE787d/KMCQBOMeinMOx1kj391XIMKjnW3CX15lE97hayT1CBxtowSSPvWUadg
Ia8NXAJ/DcM7yUGcbqhnqGvk/28TGf1ntGA+14eYqqn8LfcTFNkv7A2cdeK9TmA0ZFD9dJYQ0H3b
N/EudGBhSmNFef3FeMVFcIZz7KnmUFihPVCJEwrXdx2Fq9I86/ORPcaldE0aC5v1XougKhrls4XD
Dyl9Z9ztuGLEuS7Hzl7W300OIvmlthwBexwUfP7sRLUKtWB6VNXdPJWzaLI/Cj2pyQQ6yA1rLJZs
qXNwssYvKNUayZp3rN4eJQT+ig0OYwC4OyupAqr0hMj2MA7Ls9Uv6vv3tA4ftB/uXdyoH0SIVeHc
exSf1nZf+zePSDrJPZs9qr+qMjMwK8db30LDug+2ilFmMTfgasrU1BsF0Tvb6Brw8BgtWePxV4/U
+TKYVX8XaD8BtIyjgkTr1+JEY9+OxmB42Urod08UzPVEEqfVND5K7VhSF7VRavQmzWTlJy8iqkns
6a3eBthVkI1pV9Lw04UutgkLvl9UbAAiYBkH0TQWqgl8Ph5Cx9FGxSgR1vCprx2GPyZUtHuEJFbu
UMfDaQefriQ9KXmOqh08+XMsjqFC/6lSPjdfQugEpLs27GDTCOSQBv+XyZKlZ7cg89crq+hX+mMb
+2b3epyDQBIqeT8y58REOJ4tNXODhYBCCpCe3hPcuy8ZhXr1S1UDaTot5deGQfFC9OTyGTJwcmay
zMwSDup2iAh8gjjjDnjVVdZx3nCWb0WFPDV7Z4rhSzbo5mj8ptb/AdR9wP2chOiLxdqFlXGQVgyD
Fq+aI45d7JzZmGZ+XuEiDEufJeJCluwkKu49XQiieB1UUDDoauUHuo8m6Zk9SuBCZR8i3jW6EKdq
ojmFub7mCtdr338JHFxGsrcvVHo103s/W5c/GJl2riX8sGuhqblszwU4nIKNBL3bKkE+DatAkGl7
BQZEMc9AQAGg7AyEgdpIAZY+oDLXOcZq+sYaUi/OYT19jl4a1D4Ns5orf4p49exSoYPRHWh9OJaA
4DToxpb3COEjvoHGy8DkAZ5NpKR20xPCXnbxh3LTGfOOw8DMp9Da5a3reK25bBNYdhPP3U2XfZ4L
5AsEphW1PqplXAtVEkltVjIBo6O+mxDawh0f4Jf/q1kDbtSt7KvuchgSzmzx83mEXKDlCj6lxGWA
IEvArqkkRrkZ9Ahg8kfndik/+9Fuw7/g+l/26vcc0axWmk/f76v6znGukLgybAguKmR7mDDeJXjX
oMQA/qQi8tDf5/oh
`protect end_protected
