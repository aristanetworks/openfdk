--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
fZEtkrlmvdzC5/ljz1etdFGe14PG64jdB2fsPyjiMFloWDAOO8P1hXeP1vZ9xVwv/M9gb0fNFOli
pjtPli5B4pi2xzOM16rkpTCv4WLHb3KvJke9uE2oBO2CTNmHzkLisQRI9Lxn1R/xxJ0e6dg/WWSG
J9tJnq4eXDU5QFvTLucuDRQ3zqeV04sJg8Qp+LnSIDTlPk9Pu1CUKkHiMpF7pR9NU9lFvkIrZMgi
QzbGyp793+rNqegowBiTQKeLMba+fY2Re5NRLjUiR9M8fSZjj9Zke2CQQmChLrEXA0EOEW2SW95w
bTMo2G/wKbDw6RmPtZUEhwSKErMl60tJWMOCUw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="dQhB72H/uHxiCZtzWWRZdZ5AUX+w4ScI66tZJKtGG4s="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
FXoSXXADjITMSkfNBostJJDPH6TWCO2ii8wHmZQKt4ggFpDBl/MCwfCjQfbOD6JjGpcTCnMp6+99
DipvY0oBZ4nO3+JQBw/FmJc/AFHWLODQQuRf8tEwCv5zqpaXohTj7fkQXxIEH+3nGiM1ohI3V2Ql
hyxtmptyN7jBWXYoK/h3lxC0g/avHk7PTcgAzABzfssn+kzUZ0aoJ3V67XF+25/b9TcfG2yM92iS
vKVzqcZ3bEGwOjb/RjdpHwYMbJNarhIYgBG5QpgUZrORnBdLBFepTv3YLZVZ7Om1UubYOKBeM2Nf
L9MYf2ohf0rg90kMUJz12sz5uzl5/f4/AWK5Ug==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="rz8jcTuGHqnqspA5X22zR1/gxl0EFy/RQXvyhW7entM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2464)
`protect data_block
q6G2XUG+WLYKkOATs4YDpJyU0sGmYJ/E93O/7pn6UFvLKCKZIxQk8jzQTsZ8c14Wrw3NSiaGsnzf
NIrHzBKA3nNmOpALCe8RYLYoopnYKFMSkr6HDjoDTQYjY4e8X78O/0EMktqryMGVZdalziH71fMi
M/nSKlO+cV7vf+OhIM9HV+mAb5sOXtd+DPU4x64pzKh/j92ezHlDIh7jCvq6qeT3PkjCLQCM83tK
Hfu8uTZQnQSUQ7x/zoFjQG2+9rfVNY2/yuSlaotPqsZ7b+v7aGnuevsBINb2gtR6JwnieWWosWDz
L11AwFniYxjeBIj8bF7Rz0mlQvhORpmSKIOAZr2fER263wehqADVLP8QmjKNQU7SR1vm7sLBMBKW
/Wzu3/2TN2uB3445S4rx5b932tpdLgsNMM54HfOAw9YwniwRIz8vShSPx/1q4ID/pSymBCELweJ9
Znhcy/oMrtIjC2KuRK2cfepiD/A/PuT0wmRVj4a4YuU95M/Y0i5SGJwCI/8FgWfWKyjY8yyQggOe
sL1zeHu2X4skD3SyN24iuPoHyIBhPmpmjGeJKfihFfWUUbe51cBoHyZ3tYIkZovMs1FRvpfJ0QYl
AJLzOARQDdGR2ty5ojMuWDqiNYVtw/9p4qrkZ1kOgHyiAyLhW1kfuE9DIv/PYQW+8pVTTcnXq91q
H+Kb8/c1/QA88/kw1gzVHwvwgDS/FqkOOmAtWNgEfuyJMFwgxk10S0/iE6aLvdVrR4U/EsRxqUu7
TjHT5n3BYmIsMatw/EJIZHtRvvaSL/qM/h35mHk3PMu/wcAeMtuezi3B9rfw5VS8xoeWo66zw3gc
9J07mJpPwlS06ZEGQidAnvY/W/Laa+ogiXxRa90qL3D1iC8jtUklQ1CQGaqjBkLzzXSMOL4+yClv
4MWPDeTs8kUS8IMLTv+CNC2RnizZcLjo/RRt8/2whmKQH9X8cHNYUBgLprXjtRh3yuY3rlZdsNaa
chPLKmb8rQQCamRqlQhv6EkxGfUyvbYVhIWJVgsYnntcfRAnYSUf15U30IrNVBpEuyyHM86m5Zzj
WvTS/pgiyNWvoBqafG6Xan2s5hwd3JBg7IQa755itsynY1ZihVu5t/EJX8etfJppV2ag3yWp6yKn
g9CvqmiqvgqNOBSbhLHAu/OGJAleX4Pa2yWHMiBtZ7JDvxyngLlbg6AfTyKLwrG8+XAQ89Q8RoKf
LTqJ9SMyFM+o264ObbnsvXONJVM2XXsvjponanBwQekw8tZ4Cvlhar9Jn4gAxsgvencpq0ANTrIL
rUXAtmSfKPNL1AQFAc7c/Qzj8hmPF6T3on9xffe0J3TbcSxQE/w4zq6VibvWe6RNvtXbzuE2kUoZ
3erRc/q8p9ZLOJ0whcRko/9Ntha+N/kjHIO74gEjZ83eobh8EG+wHnsgzDXn2F+5G4GcNBXI3qxJ
NncmqUcUT1Ld/fH/7w0ikIQA08Q7q3DpFYKl9SYoqqx+uWFaalT4LVKGhkf7dKidyMNb/xa/mh8J
hMGA96gBpSUjuSIjZl3RYnNIkIO4z7YVGO4Du9BIHd33UVniUM6hPiMLTbd9hXfOUVehJ4NTXUpf
MxzLjmTr86aK7Yuk2pOIObOvXqGi9J0pxWr1hWF0pP2BgjjMfoqMz4f91Rpbc+kaTaluZ+oKdhIb
IAqZgiYh3ywXCvOfR+kL5ps1mCKebFOmDpdvQYIseJXSR7xlmSyUR0x7friwg7+b286HcmrKr7yS
SRNQ2v8sjW023t+lDWj8vL0YhWHTTL24JVkQgs/koqthkCfoCm6TxSC8TugBEIfqPEZk6xeF8kcS
x0vB585WIUwgx+0uLFk+7IDBKjxav/XY3BwJsD3OgkoF2RP4smrHZCml9KQ+FwbhOXOCeHAYTTDP
SXg1HRwIgtwwZwpNzKYzPrdYnUxC4EBel/Ec/Gv4PSjWCXsHBxNVS77kkK47djsWjnD5tp+vLrVd
iWu7Hs57X+/oUY3sCflgbit382mRFIgpQWEQQ3cHdeFCebUWXUpg0Kq3qrU+9UolG0x/vWxCgtCB
AzGvutFtOrsDM0ZT2IqTSx6ZuBeM4sOdbK9ACUlO9brAV9150lL47wDbGI1unytPK38bRCiOYJKn
55Zezic9bng7ltWWjgR4kDfq+0BWKzYSipglSP7VZfP44NpJa3r8CK/h0M+xqC1bpzD3UdJ0CQIM
HFbDWpG4MEjBJ7UzmfaRCKEgHscHs4MiXReKyMWb2+EDNqKaCof6n/YY2mdnxMNdWU/GA6kbxVmM
ih4q/5TI78SxLG4d7Si9bt4JE5D/N+bL2e8BfjlfuUbWLxnPgP0J6/RxDKtVJzelBN1paqonny1P
c5JSHLhwPRKSocpr2WzfiKsOYmkl21gjjEz31s1dKvKvPGdx3r/ibyEDiurhCpHp4X5lUueMys4O
qRJBC1Ih3PbdoLQF6Zl/uyuSXgn6MyyuAW3XkwkXqJkHsO8KIMl1iSc1kSGn3NHYvv+vpIL7Gtvz
emI4SuZ4vOEO8AHIXS2SD1PdWnnKoAnrnzc44LDGSL6bionpYl1suEvn+M9gKAn4Uu0vD8kZXjq1
U58aepms4JabWXrbDuOUM6Eph0QXynjBlhAiPzOMsMY/rJudL/rgjH9U0qF2AWofk0CXgBPE28tb
B5ShtKO6+fxnDui3s3yeyWkijvpThhTWuERt30Mpr+voY0C4DIu7SdIz2eeVBrV8xu9fGnAjlEZP
lhId9zKuI9KMShOjF95QNpy08PDEfAjC2DMZ+diJcekXOcFxxVr4ZigJtV64xXYYQF8HPdBD+CfV
sAVUERDp63RqdSUglM0egSx2wkIPXFpP0zb16nRUvzYEu3Y1yhZ5XQDHYYM+DhHCGFXbay0wXaAa
mWZ04cxXIrkqAmAsmRa3hCWktDVl2K+7P9p6FHFzRGVEd1W4FRRPWOgs5MhayyVw3AsgiQ/iBOcW
HewYVaiSpAWBSrpzxf/ubZIz5uIOq8C/Ii8O/o/rHgTQMQOR5zuA61jOqTvI8gcJgk8qGtjCzMhn
gslgs5op84dCIvI9ShO/siKuqNRp7B2cUWeqv38gqNnUC0iON5S4xt8kbBpyfpLhD+NOeJyBakfk
a5Y2C/CrNCQxNTtW3ZyFat/IBTyqdoYc0kJ81YZWnQAxRKHN+emRtBOax0R+VqkGBhZMyYAludkm
vgsUXGgCYC/TtZwRdENm9us7syi3rzCopEGBkw4FIpR1Jd4GoTiRmZkofDFU5D8ReL+1quNO2PTr
rWQF5y5Xm0yK1kCybA==
`protect end_protected
