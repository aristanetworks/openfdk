--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
ANx6C+33LfenXHGmom/ddmo1csCOcX6w1M6gGQjcHE9q6y0tQPg+AAlnPxKkPBitAMBdVDfROQm9
0gfu35N5taKniCyF1R6FLdsoBjvOdeYSDVb4ToIg0paI2DO4AZmLb/+T8eO5TVZAEoCIP0GK6SGI
uPQpxtwcjKLjDiSEUG366kwKtx1F9sVB/EmL0RYNEepoYJEspxA+ssfpliVmrNSsMOioMThEjIXJ
3lQZuYP1PNaDj56YHK6kyotwO+K2eUjgoqncB+CXZLCdaiNw3VOWs+sNE8QWoSWVzEVXoOmZ9eed
t8JLFf5TcDXgN40eK7o9Wh6mE/ZlM/9Lop3BsQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="wJwloFDxodiPHkENmLLwreJkQLc/f4SB82dfSH/dwlM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
SYG1LJQyLrd6NEXsIspl6E0vfJOAlbrEbHv6PhAupXxSGDl+s0ftrRysKi4EHvrOnYaOxl/HNRBy
5Lo+HJaP37UsOwBS+C8IqYhyH7HNNIDA6V4TYDW/Spn4slkDPL/QzX+tEIsWB/VafWOyhsNVy1Dl
JpVVDXJJKaI55ID1x7lfLy11NqVgzeleyHxT8dSY08IuuQbn05N2oox9PQYnTDI4Hm4y8LbD/gXK
TTGUQF38fhjEMfUku7mkeoggj3qh2kReFUOA6pTV01X2+/4hsqx4KimqaELdsUvUKzscOd97/SbT
jkBR1kd1t7cX2y8azkz9kK2CLucH4xqKXC9eYQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="KcxCX4hft+H6P4PgQAvYagj4kBT4eFq1FqA9A5oBjD4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14864)
`protect data_block
/zOcmWeToaOOz91Lidyux9gSnmos5XN2TE+rHRFmO+6iwSPm/QQXrkie6v7jDgIPlcAM7ld2a66y
pU3NNIhj2d6F/aD9oxJXYs9e311jDj3Juv1diVVWbvmT315D7hQEIu06ihedwsbkm31QQ4oncEfc
kXNm9UQAdk8dlWuOnjFOkWOBdi4Ln0cIRQqKWfPkIenlwezfCqdA+5DIoTYuYSmz5BnpBTKD5vVq
EPf6kmWXeVrTaSVOkc3Wr+QXuR1TzrLwaFn/K63Ak665IrwC2XkUVMe/pypnyTecLmsAZviQQHe2
NRxttxE5uiAx4EZRJi2hKbuJwcoJoTysmT0NkUMnemT1b2GZb92esoch1+sbgDld2s4yrGECX4ti
jYdheKJiCl76TK/1sMsmVXBtfHaYHv92jcHKYMQ4YckUALOQO7IXomOksQ7k5EzPA/S/LrhY6M0w
sc6Vjp3kNN4EpUKn8nShlDS513DCnyFe6oPQilxcQEghmFyO5QMcai6z9fcWn1ISM5r7NO8hol28
zuYzXhehHYlmV2XrD7XpG5lh5IgIPHJIfUqyWtFhR8IT6WC/ScvI4XHgTKbvVsBQkC6Haui9rCnK
J4Ir5yuDxuZjl+zob4oFZK1bk2Cr2etT0ZyXdn5BX/NYmA/G7/6BLku+o/1pctRYqw6ZHUCwRuKe
XRrQtuZKpMKvkWwk957zGYriwpUhcacls2+lViFkTDr3aq1raZDjfX8cv9kQG0D+AHnXTsaZ7muW
iq9F5IxVfKg5WM4pkBxVkpBNlAD6VDzp1QaUU7inmALCOTu+t/Iq3v3qHdWLgfbVKKxAeJDDGISM
8vcHfdDKeE7PBWfgk2Y2em/MR9f34pU229AdkC5PFXQcPfnF07ksCuvzzXvije3cbBpv9HZK/CI2
27Xq4dUqMjyVAjeVCM+KE01LRPiLTqjrQ/bygHXB8f2uLX7Xl4YUO3DuENFSJTpqnMbkmPjBweIl
m3SnfE2bGCX7hI8JWseavcHO/SsHQzPmFjZAh2zb8x7vF/SDtetixl58H+WKxre+QlniC5ZJGwjq
EYx1vclGUCxZrsSAMjDCe0RKG90mxwHOn9yRiiFmrk9ocjdzfo2pbrFgwFdmgLRLcEy2K3g/g0Jp
HegBZPl8l9nTKsUKBsfbr0S2Q+vyTa7dP43pzgUGcA+kgEFXNZ0Kl7WYIRkaB6UyXXWSR3NBO/Kz
386bg0rnImA6jZDCK9u3MEwOPAWMLj0j6Qs7AEDdw3v8zIMg5rOMovuKugOmnTjh73HWnHXOUjzF
F4BIZxi/Nf55kIRYxrcE+8lQvFhKbuYynRkfOSaNh40YxF5eunj82sIBlIuVoIEEdKIUvzsOgl0g
VYyxvjDyFtcjPMh11Oc6cVarStk1A3U5z4AX7SriDmc9EfimhkYgNx/+2GcWlM3SWc5IkWnfxBQt
AINQYEBxN/0rzvxjIQSHr7Oh/RourS8R3Ie+AlyaZN+z2evxOACjHKORVLPlyqzxn18VHLeRWpeA
y+73DKFHDfCAj/uCLgdhr2QgUkYG9qNYha39ngeb8FCe/YQswfC6QwmvukLL6zOH2NuPYFyd5qjp
t8JfJR4sUi3KyGRsGQWVbvdXM5kYDybPjvYAQvS5Z3yzqxO9OjeDRy0kjfkZVLqXcCKjiNKFEVOK
3klAeK8GuhX5hzetcVdakRfw8Qv2u3qaRSXfxCgY+WSU6AeotuXjd07Jb+Thz8lS7YpbxO8Fk2iR
EuZ82y5Vk5iL5X6giBNEcvCUoLEjRM8LGJphGCJw4hdR8Wd1854mQW2lVFNzM8HXjgti4Ekepyrp
mTkVKJXk1jneuNMk+weJnbx5JDAG49d6MUl3Xqw9bxvYscvE11a8LdcnlFp8NcbqAbljzRbB0WH5
ydg0x2fcLuXWqo+smhCp0T+VMXyMH+bn+3gPWH/iL23cgkpYWnbLz1FYODTWuzplefd+1KVDTCMS
ffJl8VqAz6EpCHHN+vgwaTbaY1woI96hMkEx81QqFOAIgRgCtapBn9w54oD5x/A8czHPJFJRHf0W
mK7OtJNaqs4liCyO2hToKpgZHu78duF9ehSGOi+xDNhfnJaMlFQ6uk4z2WxyKh5kvRTf8UJEZFe3
WojLrMn+9OX64Xc+iwdHtER9Z3q2c0vCGXRdwECDXOG/vVhEYqDmZ8iqAXRl9QVwJN+TT0+q7JeX
WWB+F60rS9nTogbI/iAg37bcV5FfU6TfO9c90XAtbjp4uT7fI1vDM7dSZS3ZVLFvSiOZu3XnCihK
CSCuny5LFzUqRufXIFFFIwaiMXBiVm4kWbir4QbK+WiIa/FGiUBvioO1PysrvyYvrhFNPxBVscvK
tJl43sQELI37XgSPttPb3boVvG7XJ3MejE96zUCrcnsXs4BSxezkIiNZqcOrMZX1BhsNH5StMXKY
nno9efas9godJog1umzcuNpoxwfXzicmw9JdKTzxeplrwR36yh6/0vDpeoNzz1MRi6DuVrtSNVM0
nHWyu1iURKmPNPxvgSypSTbxBLwn8FLl75p5+AATxTx4dY6jat214M5QEqNUj2p4jjIpGe8bCvzh
X11owyBf5Vh2dnTtv+iCGuwUJcKs4GkVb2LSG+oNJwbjl1gN81gUjA3w7tPxhLicDGBrDUMLN3DV
qvzXHILLqiF8Et0c+La3FRu8Gqw9jcImXb7yIZbFC6D3lizQSrqnTCd9kREp6eoadgWuLSe2IAlq
fhSTvEupbTeqcWSnr7FHSI6hMpufUCD0D5A0wSl3juAsED24QVhSRtmHlkhaeFMArX787XqDCQXT
9X9zbwJur4zFy24q3O62glT+5ZLqViY+dR305mPpM+QyLQO0dW78rr33NibbSaft+80dtDXPMvpQ
f8AXciCvb1IM7GLAx6CWYQ9eJoXxZF95jm3d7xCg5pwSV9OybGgFU3BKoUEDZb20dsbnUWWAqf48
pCXjxkyZr11I5ev1wdKDAVua56g00IwISuUeDufaddJf7Hqu/4rW8xN1SKZYqhl/RPD8HwjwIjfw
uDEVtgMtkqfh8trvklrBAYK6UBmX/ZqtkPcsnd2CHOPAyJJMyUQaNZzlbVl+XHGwXKgt2KboV2tT
oH6QP1evPsJtaexD0CnEEJqbZfFeYEOVcWH4JQQ4TnpqJdhMSCC9H9RF/15QABVgKogpgSSs6BkT
Vz3Qwt4NghISNcganRsjgeMpHKxol7dQ5Gv8c8Z00OYUI3YOkKjWv6ZbUPL9yvacQbEGFNjN87cc
BBC4/nO3m+qghusyWhHaMtI85fZqE4GFMv+uDinumqlJ/yrMbKUBm45hw0gUoRXwEa7dwGaClPtS
wWF2okpfogUWlxu7xuzVadIKqLGewrOn4weSluBUhgC5qNf19Ud6ddrGjjhQID5XUwieJMOm2Kl6
DhLry74a0vQ6mIfcNyy+/c9GpSXS9F3ckOhk1aRKmmcvkHgpfoAmS+QlxQ6V2pClN8N0SXQZ2brR
Jum+x+ZZJYWAo6062TNwDdF/97OBSSgnz8IWaeTIBIvBUMsdADB0qZo3hWAhNdqHHlHpDlbVhm+Y
V6CF5/E2hTL2t9Q0PoWqmH+hK1HFJ48jwv2z4dn+ZNg2GScAw33dzk9KqG929xWxB7jIfpTNDVlO
qezlCaxp6o7RqUY1GZrwIrizQt14+CIy9rLaUX3/dJyEAte/u4tyCm5vp2L4LSWJNm+YrVvzJ72z
0tjPd9/SX2Lt+Hus2qcdCYd89JP11JxVnbKeRfL9ZR5sCE3z0G1KBVZSYwdCX8tHitAtHOyEjCnV
7Zk6yh7rrcL0xlm8wtBSIlBY/IdMGuT9G096opM/8pD8WEdcxnNH/T7sBPo4Zm/LnSUWXSr8//lY
BcwsxwD9jhGOq90G9yoCSkM8PFxAWxqlerbyqEKGsjbpyekWsnJvU2B5I4+MdnrSrrHUxwhqeKPI
0MB5U/TH8EXRNuVrjq6z5+b6xZxEVvQvPgiqekwG7/QZ60lLAGy/c/dQjP/QEilHSoWdiPbWmfil
g1rs3p6VBYts2wRPl0JXQ1r4WCrCON6aCMzIo5+KSb6zg3ef/tBvC90vfgerkMsAOzxKsFhDOjld
1LOnpup3a7y+zhOWezUbfRamh/SRk5oNPLsYBC4THykWMJwuzLRuzaIz6iTCIxg4M1++oG7EzdoB
8hPjywEvZreNFEDpz6FODMdgQni1/6tsXLd5wZJ6QeWsa1y4ADBkPEgcD5hpOb6cVXqIsYtM/Knv
ZUiRaxz6On5bHhJQ+kVUtiNvwccrbjpSSdJGlJ3pChuC1ZbpBRNEaN5J2Y1s5HZFZGIqTI5EzLWE
pfPQXIS8dyVgam2RvBwBzyyCqMsvafxuX9naadWm2zw/aNDzqS5Du5N9IV+w8foXYmBIs+pZbqIn
XnigEWFHGZbEE/e1tqu687mYrhmH/JmjB07ajCUm2Jlih6JMkS575ku39N+yhsfAnmsdDkwyCiPr
KQ+okZh6QMlwzOzwTEumQc6qQI4rC/TLshMv/37XVrBYPYUy/nja5rvdEuhANb/wMS90roJpjMW8
OdyVJ+QiIq3fS/pHdbEhGmr7Jug4k+ldDCkXPThY++x8LbUU49J/4e6GaHAzm3i2B4WiTX3DnLTc
uNTlh6VEe+KibPw47hzopjiFJ3A3NaE2IC8BLByPBlI3qVXpxFA1KCOgdop5+YX0Y+6roaNq28iC
UNzV1oRYd+ocbg9wDUBXLaYk4AN6IrU9p05Hrer2M+pt+brLyn0VWGpy2PI6ZCHnSRA+soAwgFqZ
4vcS9g40jJwYyoSwM3mth0diJ/en47Yw+CBtzSIENzgdP+fd1idtHH2F6UMqH5agzMu3TjdAZgpD
YC+2LcFBCPrdjoioPwJqv0ATu71L+01fPG/hKEWi4jQi2yFLrFCdKNJsu/mlp4/hMCOE/gSNv8vT
CboGM+N5GhCEZra4x1wx1H76AbqbKY55qezmd5FpYxyrZNdg1fytMLeSa1TxsqHB7rh9r9eNrZlF
LZ8OimZiUOq0LIrGjWy/wvAv33wxUIt4WPXVmQ3SbUVXx1GFpmSZ5TADlCer8hEzCV/GMnHyP437
gwFtzGTK8vEDXnWrFcMJqq28PRSIzVb5UeWeCOtMC1udg7AN2wAK3+rxNgqRIcy3V4KFY/7IW9ba
3BbDlZw8i61rF3fdgVegwHM2DhzBIxKBpkZ0u62V5s+ZIJWZ00IDGuSjJSmf9jOZZCfldboNJRmR
NcbPOdGW5clSv8zKVhXxmxNzEb+4d1b95rUMdBkyMkUQd8gyvhSrooUvvEVy51PhnyWKH+421p94
wyv59jiP8ENzwJOw3uZvP7TX+idHgVU5aegJY3m3a3Uj5xYnt3GuWDLiqCqwfWrtR0rs5nTgzX3d
o0G2s6ONz9nFcFIZoC0jdi0wC4Ayl7pwKOio7w0vqS7flkKIO3JW0zChnwfSV0265nvv4QK+D3mz
kZVPXaNPdGXS0XPDCwxmxjtVKQu3rEj3eaI0l+LajK3DhvGAnBXWzkng/Wj0B3XcSNHV+ivsfDjZ
bJt4LtZNjMtaToAxpOYZ4pbj7s9OYP785fDEQLMVeYg3Jd1haw1JRpoE092s3AeoPm7wXh843gSR
2lSn0rvh/24bBTfvf0skrp/uA8tJseGC+d2AzqaQRSrfPQvK5i5RR/nMy/a0q4cMCGnKEd0WPqYW
TIYSNd0HPV5/wsPOmb0v6VA3EaK5QNZMNY7cIS2XEh2icM0jQIS/72MU17zR8IztHsTaPQfcCQmP
Tvp3R6OC+cHhJu8+KGWnboXNxNe2gTf756B+xYT+gNCtifRw2G0nyF6o7cS/m0IdIsnCIhJar1YN
yTuvwDJXOcuRAeHPmTZq8bryFNyIOYURXwJAXQwSwHu/8YwZOlWzGS6yoJ9ky6jGCJCF/93pkzjP
8veiwmpMLvCQFZaIiotXcVlFJWpBZtREmXou+o9c4pIxSxvdNms5ARMziDWYyJZxgPgVOd6pJSyv
lj0zextUsOcfaqvNvFdHGzFPJ3zCnobbROx/cXJL+N4+Ze7auc2OxlvQWzL7oi+rBWuLS7s8/QcG
TplyM6gACoNpbuRO9NFCiqesqUv6XwEvLNpG4YktjKkSzfhOXKLqecaXwbJAW3GvRgaOjCm1ToDx
lJpYqYIwVN7lkGt1DWOiwPffpqAnatP52DZNQb69brDyulEHlK65BI6AgV4Te6emX5R7WdIBhL4j
598xgjB8zpSdrUKtsfOrTetDVOdE4ZLMnxvmWTM1BxuRtgBO68uDfrWgQHG1/knynmaOmwt77jxN
s00KAprSaplw49NLQcPchvnqG4crjTSXWSW+uk6jpUXMW2I2HuDM9xf3+mLyKgW7W+wPfoYXDmkK
ZjAOJus4DVsZO7fNfUJ0ohUmZhGAHtBNa7TAGpVtZYbKImUMXXzvcfjxslr9Hp7w+xTSRMFLaNy2
E29O8Jdo/XQveHizZoJ78G5Qmc09bJxBTF2uGO1eHR+WcviiB8ky1VlcBqhTxRenbUt/r5f7yamu
UsqZ7Zfrjccg7p2UdUzzYHhpWNG+WJ5MZm9PmZCjxP656mXzSq47g4J/6RuoGWBwmYJPhzxBMFlC
qyaZA1Z9LzooVbGX4+cQigyIUyIsDaoEjYFcaSEdg7bx5kvyYLSw19u58hZJjoEOOEMYfu54lO8/
W7KMWluPxv2ji+uf8epkYuJsH+I2wYjmXS9Aky0H+jA9yEr7czmQjMXhW9zcaqy8riD35Evrpmel
243Mp3HrpBM0XMgQ9CAHMgaqP48SiNdl7+yNIm6G2d1HLZHzFhc6GxIrlmF71HwyIox9+G/AH77s
j4j1VAG0quWeZk6EVdoN4JD+xaP5LNG1dbTl7mEcO8QZSEto4xSDe1R86pIZ6njgq1Mug0Dp47jw
+RvLVy5uW16EIt0ZG0DvlXQ56Xs7Plzet9R38vE+6HeyopIx9RLxaTeFOwqkCqBvfzja9TffaSUd
UXfSAfroyKjxGhzWQZlB7gxLo64nNXidZqRhob+YR9x+Y7S5Pr8rETX68TPtE1W+Z5lRmFlqixlO
XayrIsYY+GHyCteNgTfaB/YU7IKhsL45Z7sTdXDVxmXkL8o53YbrLSUNQYx22B/BQEmufBqqqxwP
OLqzS+MBZIKRSLlvu6145+V4mlVVEHVK3anBAPJvfbtrx/5GuXVqdUQL7pbNmfEXZih0dh7RVUHe
tZTS3b1l9NBmVoerHLQCxLT3qjLhVqrlvf6jAua8ROCd+O+8JwjxchLjqN9oX/IH1G7IsnRQv6Yr
t5L+sRR4ceQm4plyyfwdagLGEBMjGnHOocEPe7uwf59ILTDgZQpy45XI3qJEXrup9iVLCwchKMrp
cZnCQbCIVi5VUV69Tnz4HzOVfIXldnJhlTMnjDonlit6w8D+sILOD1mGo/qQIX4zhdgB8Q/EBW6C
V2eCP57KXOAVjutZuFqZf75XH0qkqlkaeHP5yVxT0lyNo/VPCH05N9YlA4ywI+0hOXk/4rtSThOo
EtK+POhNyszHs3GroHF6ZyYK9asVSnxwr9KftTekSGmR/bOjapz3VIE0wdvfAepOj48UR0uJhFHS
mLxnxfyTWXjQXW6Bdbu7Qdv/YaENktucOrIAc2jy1Q8PCD3RPu6RmI3/2BwBY/fe+TKT+nNinVPf
on8DdW4nOJpKk/zgFOixYSQcbu+xmdcfPACgQUYJMKWwA/skVqBX9PIU8ekQ/I3kN3o57671Q9Ig
YMv004WHpYD50oNQs+CKZKVNt1no3NYSXitGcGivUFd96Vo9xdbEab0LJjpDiO18Bf7A3j7CtL5O
sdZXzccQxZ6XoUk0mZar1KG8eo+aH53KYWY6n86iFwntkGtpdDV83OrvJS3svaIDw8R/DQJwFdHR
hcvxJKj2ZEkRf23nT6y9yPrQTUpLaPMrdhXyHFbl4DC780B7gj8AwiDtPowojiDlaS9SnvKGNIFk
Uj+aK+K5ry91w/IAe3i8V0Se8nkVg8DdwpptgfxmRoaBmQOPrNhm3qzkgeXu3EVp0DOzNXdyZLe7
ep9hQH0avlm/IiaigKG9lzAmhUl8TFGq8ToCEnbLHrqXnMeBpVQ4GJqKvke+17VOIX1nLtJj5SM/
hDFGRjOLT9YKllrFGHvfB88hu6M00854cx/P6WHP/lmLx6YYyfV/AtcLXYgA3eqXt9/wQdNSulja
XEscrlUOvjbgYls5QTfyKbP5QjyXQ2h6EjJ6+dQ9yd8Tz+eRgmLp+D306Wb2oJgF7ntTFcX0e6JS
NEDUwwXo3fvFc+s07MvNbM3zkR0mtkahGyHmrsUI72p6cA/6jHYwJDI2ezwxeuxVGXa92TqA/3c3
YUn0UL9Gsp9hUFpBuJzWUmBzAiqhbXkkQlHjV76XFuJeo0lCYuEbe5RqkjDpNczhnTuWlyUOQzwk
Rc376PJKQF2VLi3NbZIDxh2xN3Yw1eH9fW780NY3e2RXqJqDCoOBJlimV0T9uF8Ra5KoGgIxe01G
CQBFbBEtKSwFNzJ9CK3Z8+4f+ZuvKBhz+q6Qld7tvTDE6ZF3tm8yZt/nUi36BswX/A2DGese1O9a
IxOu48PyrHemcsY5JarCybzLh8pd+1fDPQ9kxgqciL1bXe6lGFv1YXkBy4DMqeobyxWu5fw1Wc9x
Ssd40fHHNNMXOULPYSraaGTM7P8ZopQS4ZrQN7o+X5gDNa369N/zNOUzGzQXHMJngE4Cv+r9EPzS
zRoRqCUvB041lprXkB0K5BPuAleDDX62HOFyA2vBvIwXNWNQxL6En9UmHxL3ibzD8KkTA50Losnp
u5gg0uQixx1sTiIEXId6//Q9J757NsY63SzOEKxaS5qjfjKbVEMZ6D/aEjYOkdhAwk+saRoYG6K4
EPsFb1Og5fdNggQHUiDk5bYJ8YQrQsRDGDz0fV92ZYa2rSCKolx+vKnN2GKeY18XKI62x7sWgZF+
Gug/GFH8Fhdrkmh/bFHhdIgGT9qLUqAxD2+YfN3qKXwqM0BiBuBgH762vSfVWAPns4rYDb5uBsfG
YA93f7GF9qEqwDmSJiueLqmI5Zxyv7vXgryDAQtSBTWnpcOBVYsFllNZgzbyEDoaYL2J9T1XjIlr
GhNt+WMPFIcH6k7mM416oEJ7AXifDqCsgiMK30TWb4N7DoG7xfqVdU1JG5gXMJW8VBt6inBOoVsc
sa2OcRygW60MeMRFV8sad04N3lGiNmWGjJGLdqWkcD70i1h/JZvjDiImBB5RbptmeLpGMnXwTvFX
0ZfN6+RL/JXA4Iy3ESR734nuy3sKXNly1AuIcuZorCuu934y8FCfuKH7f7ZfAv90POPKYyL4IZ6d
lOoPwHIkz7UWdD2G6ULIQO+H5H5ZZegTi+4OXIpAMXddAMzQhKk5uAW+ioZKCtxxewcPDfYbioDB
Wf61MN3I/Jrc1aIjDIyRDQH5FEfSJhJ4b2yqB7Is9pMk/yOl2cZSIrB5Eb/yjon1su5SmghpcTO6
jx4M4XqoIeFVlGE37fmcv5znlDKZcNVgDI1HYBAXjiOcdlqrq3dfQrDxKaMd6r4pbcknAJtabYrR
/VnciAxjPBgBOxYE4jwQzfxtWjm/qJp3bN0s8dp/LoJ7pP+SjpO8BxWmaqKw7UevHGi4adntX0jU
NCKcVGRCFXwQqqbH2jDQ7Q9W1hNNfpYAqVzwORHstBpn1ub4I237SlHiJzeS7b09kxfVRc4pyhbQ
0ch1DZSnSyiFIZNQ6sCEVZaL2TQ85h45UWKkgMPbMgLrbF4fTDmfdvvxqFTv2coeqrHaGZIwZNWm
dn3qG02dARJp+R83M570nM42uNoYr3/JO3ihJkyDosSx2hezXzXmODuuRTmmQvIhVNxHklesQwdw
3YO8Bs/Ym2ANSwP+VUnXVL4k83r/bbo/mzpdVg5VGzWGE6VXRpcXMBdrZXm74oXfo6NwzqAVJcre
sr2euillpaMr7eO1O7FpnPo+qnvrYW2DhVNUVPq8/x0M2yzGJNDUm7+E/XdKSg0UsFH4IyuqLqFZ
35CKc3xLL7vFDkXC2WSA5AsXmx+EXy9vXyQHJ4rzDAeOBvsr/+OBuIV/4Qess/wimTWqyeZP05m2
mBYDfPuTbDl2orJH8HNVoAlN7xR8NzRtQaPIgGJaY8ah6UAkfmmlDBHLdVjRCp5z0xrN/UxJJUR+
FRTi/ABXgk+5IkWkqVMRPOZgbmHch77tDI0P44rc3+H1F26h7iKlWNO4T7PPHB9l4THTnG4RDB2o
EqcBvlDhJI6lYgOYehnrv+0UQLJFmkTLD2s+xwBXXp9e1XIOAEmdGSvYEHoZD1vcMkJd2R5EjAnw
/kSDAcaawbLaXT8pYLn7pPQS5e7SFntL+ZzdiVjIvS8WgIbysKCJMfoo4TdVwV1D3J1xUasx74jU
Bbxqy8x9+D9esnUON5V7KSJiE9M8UnBhuaNTpk+5RFj3VwLSqFp+X674hfVx9imVG3qHfUZM/Rbc
/XC0hsVc1Gw+BdpWujZ9LbECTKI4rQ4I3oSkBcDJSZB5MhBuyhDvtae8hFSMaJdxaQB2SuVe4K6E
f8kBXCMvDS6JhIwTGULf8jxFOUsn/tdXQZMENHi2o1jDCD0xN7p39hyATeOeqnotDIvU2pJGEiSV
wafaMEB83uSoS1O8KghtH1kCpX+8BIy4jZAATq4R2yomm3eEKfIjg76ny1Il+ueTrXUvWvwWM77t
N77KQpK4Gu/jGjjRn0AxALgZwNnFkTBnpq/0HWJoOiV/Zm5ZpZV+WcJrfAEulouGdMl2/jYDD9+Y
vRNEpwXh5t1NArqTVJ4k0GrvosB1UmD8rFdjg9H1QXvNznEwpsKfXv7NomA3ps986roKLe9kqg62
c9mqeXdcSx/TVzsG31YdlkYBgT1MwFxcVymJmG/7zJ490LNnIpeDjPE65wZdOirvRR5GLu4IN3ep
fQHc2z9er6e0P32szTdDy5W8Xmiqje8XBYZbGq9hOhaJzvp6sxzpq4FdhR0QEsYmqSK0e/p1I4Lr
JaGaILBFG6kzguC46wLhJGnkSAMdGCTDJLdwAn4+/tc3b/mn3aKJEGJm8/HuxuKglNbVp0PvO9X4
on0hTubSWXCAZSBFgiMy/cjq2X5spLgVyMSCezjCB4C1nmcMVkgiqYmsBtzNt1UopC6A+L6JNv8A
llNRwTCONOsO8H1j0XKvMRUIzSGGVsWUySDlI7fWadiN9x/KGMAB9RKUUVQ9ux+wR/huBjDy2g1a
+r3QekOJp11flDFbj8xRJC0+9OcDmGJX2U/74mYLBHcQRbLBdfz+j2iUQQ5Dk3Hqbsq1BXoXupn+
ZxpLv3U9URo//O30ZGFiMdfaaFpfPfZMjSS+8+Ekri/Qix7YyhagSHvG7VygO8m3XOZeR7zEJHob
9RWPdbSGtgWXbGBdQOIPmzKeAuZ92KB9QLOEslDlzQ8SJR32iCdWgVSK4Nv0TBHiSxxsbCGNhg1N
NMNBgUv5syEoik0sdqdUSp7Rx+TjLisiJkFVxxj9Am+7VAdKKA1AoJyfMUrkmfIpzZScagBOWHFc
DPG23mUUx2NEk4rfb63zwcyXBn8i9JaEG1pVYHKmgglCIgqv2gG3XRBdG1k/U9JOmZFScKTG+Vff
jvFkepgGQcNGbxY+DQjMmtfuiCk/+hYlBrNn/dLwC90PN7cjwC87V7ofBK7udJzzYTBWTzsvQUS1
AYOTLglQtRQNEY0hu3eiZwNMAN9+wjj0MXX7XJpr6Eaq/CvdV7icchuo/ODIA3x3B+rOx5VvE3A2
VFRTICdvRK7y6v8QnPZE9438iCXvLe12Cj58OG9Bl2OcgA+cbOWi/49VgYEiswcBgSBa8hbRliqP
5hNbqxu3Fr9p6ZqvER6evSyZ5rxhKnn94DTFo4GDCgko3Nc585VEVKaAkcCbIbQb1B73qsIcyHli
FAKlHFZ3FcrfsHlbVBUUEsWa399vDX+dlcj8eiTEJPs5SjoNkBlxranlZ8xjAg+JTjGxytGod62N
Tbo53U/T56u0E/mJhpMT8OMM6XRKBXO0X/XOiStCLn70bbugGEF0m05EAKehjVnHPBsYNWAg+L7a
RrSmmv8Xf0xMmPzc05y3KAgz+Z6Ex8zT+nXd0dbHllwxaGBRJKiLEbP9Bspp7/G2QLjvJYqIoEfe
gBDabVMgf5PSRu+1Hp7GXnXl/MRF03nIOzVdlZDaMGYYG+aUNFf7Sick2Wxlz1PEYDfp3tnecQRU
ryE5iX9Q/boKNhln2RMM5PgYdFlOHSoxlGdhtiASigMNF1FRd2snpZCiLLYbVUMLXzz0lM7RRJNQ
+20qGAGtAzDQ7JzOCU6f76tn6bd/XwTUnKYcooa5mI+rCfVogsCzo8V2NumAhww98ZTb9P0poCrT
5pFm4wDHmDWceod/kd521W5n5R2PcUhhta4e8DgC08dznJ/NTqVFE+IkxNtXXBLKNI8aJ6oj8TIq
BaTrnSN9M+3T/yiD7lZDTdvKXzjOHAbh5OCbSvr1dohHSayhwA7pTIGOOOsWuXsXSBOmRyTDmpao
4RV6ep2Qq3STvMSZmqYqxaJcJwMU1VTUKEoAwjjSm/9mR4sDTAD8Fg5v4c2QLa520Nv6j/MRqD1g
kTpPJTUMaKML272sHFZbwHssxpM9fgpII/WpJ+urswb8jWM/WqiBhsJURBFe9zWKlNkIqIbNToWM
w+dBrTyhYa7kZIaJX4imkyIO6RXTrXlUI+7tH/BkAfA2obfIPXRD3BKn1/oeeE2m18NNqgg8+PSf
0BexvyGDwCWH3mX+tB9rUg0yJc8WEkyds1KAW/c+ttjI04faESiCVliMCSxUZE6a7uZrEl4jUoX4
lPTz+1XtCzYLS0IZAs8QlsfrSox861brH+qrGHMoLo9tCgsDhtr2r5jVCAVmFFbVhGnu/jZU5BHV
55GS/Q3ydt7a0xxYHPevUJfZ3dYrY6YWckZ8B65UoJq36vrTYbFS35RzJUQmgRtNMOBavC0UHPwl
GTlqxWMShz0sbB5CYD9hUBvgqfigN/h2EtomJ61OIhngh6oLB3yBu4WX3TI7BJzr3jvrZI8Fl5i1
qjP3gH5d2+jpEkQf1B1pb6IgZ9u51J/TYkFuPoySTOwSuUAg8PTMpMnZl6xRmwWpYQNG2XKdw1Nh
/dD9J1LO9KmY21eUe+vI6VMMHsARhCDNKV6QOHqpXZqwjIrbq3nbGTzSEY0DnvtO477gp9RqicvK
sxRZHwI91wAyYSzn27KCtmqHsuLUvdNoVq5t0NksxEQmXT8vAN6/d9QeOK3alk5DNGiZ4p80cj0D
ZYuf6BloF0dSKXiyNnpOy7W0YtgNit44scaXhdGRREfNlKxWLZwicmdyjfg0jHoKssyRxUh6OoK3
6XJUjrQEOnIbKAcFEK2jqfjz4X2s/ipetJ+8dZaxXIHsHprWw1CzRe3+K6QnMoJuOsD+U0WZpUmB
3m7dX4Kn3FfMO2khwKm2dVbddSJX1vGq/SPsd06zKGoluGr9ecfYCsMhUQ29W1HBZs34GvuEyHSV
CHYkfTTptO68TX+KjzBv+AOvIo9X56xyvSdXfHmDMH+bzfbW6roCbDon5aj0qWufIRPq/S2EpCQW
qvDPl4Dti7OHxNpr8HIbRmU2F1h8H2NXbvM5LIEMYTpnt7nGF8TxQGuSraFPHKDcBRVvEdM7bDUQ
49G5ZUOBFItihckKthEwMOR8maYKgofBSfkw2S6/3ehT3zcN+v1N3ekbyBblRpfwbWPSambQxE6Z
WDmG2ppcH9sYxgqs+HNc4X155LUVxqnAplIGqic6Qe4MWT22A2brus4+gisAYOUIE5ryJ3FoZcCz
aUmaerAFc233lMXLGREFbdAtNdBvBoRVEeRmeaX+eQpR+OShtMuFiUfpFwIq6hXZ/WZId892793g
+zW1ewqxtyHN1cFs3GpATmJjZbh7nWQ+V1eb2q39QuwMacCkh/d0Rvy4IOFBmGNYy4LNpdKsR0c+
7PGRF8za3E+Y/qpEmdZp6WY0D1ZX7QOFy6XrGmP5StJz0ES86OTa15/xrlEMDkIQWqpVGjFShrLR
c504EndgU8haV5dp4Bv9RHlJcYLSLRys40HAqJXKgv2D7bxdD+npHrRUbpbvHo8k+2KYFXGZUjLW
btWp69sFaSuHTZWrnnHY7t3H5zE5KJcnvjJh0FPOOmPE7U4bHCxgS2QoSw6mgQTswu9c5P9yQem5
nj4FTj3eS8e3Jzz6SBlYxh7xOe5zmPKCITDq+S6MXVOzWTimVqxNczpp1LOVtW4CESEFAV+sy/hL
5qxLEGzsx0v8DZJE+zcBHcieDyuz4s7cpqPE017Z+7U2nidCQHDt4qvzAX2yqYRJ9Cu5FHNi9VQK
je8IdR90Gwh2xiznnSbTqjc+1TRhSmXaIwxCHXy/IJLfYU/d5L9d2wVSpgO1ek9y5pINr1xwB8Qw
I4dq9vpt/aW71O2AwcrkaYfknMFZUu8kzbIkaAEMcoOJv+lATyqe5pxG52mPT9Ew/wTxQtqL2YFe
tb5L/3BHXr0ZV/DB/9GyEotnZOv9DQhTOGEuy4Nrrt6v74FUgHMJsAN56G6/wnyGpHZn2Tb01QIJ
UHxqn0OV+xtnGfyDAVWqn0lvZPJqV5tUjwN97d181xn1nL2+yrbyEGuORcJd9CFP2iyYCukWnS2/
iKIgW3o2Efrqk+txhuHUBc+A0d80dFfZUC8jdP95zgyvzqaxTZZYDuha2X11PFiQ7agMoBX8Wf63
JiGPAzm0WqmEPSs2zMFoucvdOIijaQ4ILoX8YnU/UlSvxItjGWwBSf2Mk8O4qXwhZ7bXQ8P2Mgj/
1I5u2l/L5ONel8czhi2SGa+p+5UMQxky9fe2Ow8yqPh75ajvWIrNiavKU/Lx2m2tbA/F5SpPk8PK
iHbiHgaoZj40/dG6X4oUkashD2FQZEeKZNNyO2LrdL35FZ+XR0QqEaYoBi74VsVIc3JPIBSLMb0r
zBivLM3zXW5iVteWkmh3xsGZX0cjDhT14fAWDdReBPipOQuuxTX+bUpqHECVe3zS8pWASnX+2eyf
rl0ZwGDB0awcIdDz6RroHP/wXWOl9S+Zm/ekK8geBorwRxkUkym2+A2TRJBQDeWkCEFILsNMPVbW
sUjHpvUdIF3A5h+Iq2T4i2dJJu2VTmuQ6JlfPOwoZfaxLWNGldFAzMW0o4axYgE9d/jh4y4EF70C
WRD76VGnsNvxtaePS3rCEmqud4LffkUehhjSktw9yZBU1zjXECDE958bwh7TxiWDjYlZk/vIwHQz
58UHJAL32+FPrbaTYG2YVrsRBnyhEXiNflTcNfq9lE/jIFvzUyuS0h+9XRUDV4GS2e36Xem67pPs
9pcZpjFFOzn+S5a4UQL3RghJoNVMKIZoXkIjzJT7uIMiybCDVSZg0RSC9+UKNpdjG7wedb0nFwDR
PoKTJ9sKYz/EFFDP6X/d7nT3gxNRxGBGS6w40CfidSr4Lh6uPjm564uIZPmkdYHeoGRvUj7gxDNa
ljlhTjsuDQZb3bljYNvwzm9X3y9Nc84gZ5XHGz853WL907lWasF/MferQ+5hOMu4lMsekI2tfqc3
dosKosEyvFyXkSa+Ub9Km3QJ50bbxxmR+dT+nhyusvM5aSPJd9FiySTwKhQ3e8qgsayKdtK9krby
lVFpzwYEQk1flsp/UKpbLdXYK5keJhL5JrSKGx+7GUYZ1a+htR/n0m9R1G3qHgLqH9nOMSRaygTc
8BijLf0s1IhRxJ55hDReUxFmXKvS6eoMm6p+Go+zJybxhY5QIbm1SkKvRgXdY+8i4eq66XTfiEvK
WR2vL1/ML7n2H+pTFwfWf9uMaGZxNTtBO2qg3y5lJD/oLGxHzEiDOQczKnQxmCIIlMxz8smGSWV7
RhBQPiVJ+/XtnPQ92duOjJ2UWbEZsqQTq9Hg+Zqy7g3zVL7o54oeopZ2iMv7uMcChyBJw5rnsE/w
xa/QdRrT+tYxJWPWObPHP0UiXDwnzfaRNJE871Axx7SnsjNJchpUnPdPqTWXpDBycD8Gb3dsjGCt
Imc6sxhvhsn04WSeX0e4hES01EtG0RvyXE779NjD4473HJK1GJJM72lJrzXgnbcWtS5KJ67bO/Lc
R5Skl2TdyWu2V4INEAbdEBOrJdM/oWqvHuiGpi4HR+96R1PtPFaIta2IjEBKH1Scub0te+h9dzVT
Ln94QMqDCQQ9V2dpYmBddi/iFPjtd5W5+o/wwPe+CSXhE9n9lnYK8Z8d+G+T4swvtgr/9dRupxa+
f6u94nGL0xCM7n/kyaLtCVDq1aqn2WdxaUuOyemw2kQ7Fen5NXStPj9jeYhnC8UTWq5IPbaazWoG
MLdKTzORQjtJ3kGMJKt3lsrDMzO12GMmV9nMX8/YZprYS3YVxVVRiCC4uBdHfOFAxAsFrb0IeAF8
jSI/nvqalMJvYcbSLUdw6AJypTg/GrycQT8w0mXgxLWtuobbgo4V6A0a2OwKmuTfkQCumPvhYslL
YTzGb2UiHGClc5xIrcJB4nsLMeatfdF64IpFCdLbfO9i2JWOVrh9hD1rQrRTnUEhQsmQzhgTRfq0
lyr+5fcm+IgpuUKS14Y8gCQ44IZagc7xBN1JYOt6rcatmEmcL48EQahDdkOec0eBVzHo2W3VodXa
ggTVomWDmBi+is1PegGKL31z+l6nC30A8jx6GOdvVtyYbV64sPG06DF7a7ezxzGtD6M7z5HS+/tS
aNWb55Hnv6bPFQ8QTQoAYQRHyYT7mo6tCmVdh77Nqe1fbtHKi9KlmQciBfeHc4SJ5pnv+QdRDB2C
K1S4CXhENyvJ3YMWbia6AffFtEWZ5fUa2vYc5EN5Lm+8oW4AkDT5nwJ/6I7jxlgEDJvrbL6eR3I4
day0uw4idXrWmYf9PPRw88OrRY9d61gdCKwX0yueVHc1ChCjF7twvPoewyZwHbPiiADF+RP3li8e
6DVSBL+dNMg/ZKo79t2N4WVmmm9xw+vzza5lxIEETK/Oewxx08Z9IATmH6WgDPqhxDHPH2Lp2HsM
hWSTWK9JtACi4kLZGaRQJ6JQK1dnyCoYduE5wFQ0Vau4Bvzi/QOxlyWtTWC+kXybrFArC70DAoGH
dbsXy+gA70d0YCW/6y0lmnxECPwNEPHL4NRErevhT7eTjLBcr00ffRjWXVo+af9gHT82p1TdiKg1
ZhSAEoxOW1mn4GZ4twiyghmRna8rlOU7RURjnK4ZwVUEyxuc5bJnuoLrAtcnMbc0Yo4J3HmxH5L0
Xd+cD807OstnvJHwBo0OqpTFTSbg0gRL7pT6o7J1ItJpFZvwVSaOg6wp9kpbkW99AQ5rBUUVjj9a
Zv3iPbd+VIVG6QSA3QUKTWfU56QjuhbSxGlvkQDkzrSPD4krYxeZ3nGOYMTlk03DA/bxKYnNJAhS
4yz5jOh3beU4f0tDcTgM2cQKK3ymIVgsmaf3e7/RhvDwp+CSWbeiJIo/THWXxuWNobqAn8Rm+5p4
KUojsUEEZCx8yi8GS/06nSj3msYZBms7/Lo8Ewq3w1Su5sE2x0IkJ+fQdK51GVjNH/nT+gj5Cb8q
m22wZgA9/8wDXzjHyfuyp9KQC02SitpACgieYMnMSLw6t+Uf36/HbYF71gmMyLHK8ihz/2ojACRi
YTATc4+mpiIt/KibSCqQ+ritISG96jEc1kKLOYUPF5/yNI2Cp/NIDfn0TolyVcbITKQmtU6zZULm
0zdqK6AQBT0loqqrhAZ7s3gvrxpcenVf1Xi5hfqaP7ENEUftjMKJw6Sc4vFw6mad4cfC2d2voczw
3DLxlpyvfJtyr9xePEcTdhdBkrug6IgKevJ1H/txZw2FHa/5DdBp5Z3pJvns3zIVBjjCTli0TNVC
384favtJcW2lzMUjALgB6aBX4b05Jik87EVjWEN10umNpx4aVqO6ox2DY1RYPypwpmUNnKmIdPhA
MCK4kXIuIhFfG0BcxZ23YlTEB1irPpevYghAlZwtL5B4iO4JCFCoRUKRHnYSoLuqnNFOnCz3ZHYh
MzF8H8iMJriKtyoaM3Pv1nlE60azDeDstgoge9x+sVq6+abPS5M672g9C/RK0X21iOuAsUijTgwI
q7G6c8YH/4NX13yo0XyEl1HL5iXfku8ZUoISvcZ/uIXQhYExiA76vHESwEQd8Z2KKNeIO42T+0Uq
b1R+meEExRJxInEZa29p2ZFkumVz7eSiADV/ce6Tb7QKLpptgwiVZNDZbr/OvYZUTLUYRvIUl6vT
p5VtzZZWOY4tZLX0wciUnHAMrncTF1HPT8Wlw+LPMnTTovI/7rCmtje1FW8HoA3dRKqOTuxViKLW
MYBmxFqu7NNJIBxRXmXxM/SGeSqKGdQbVmPAB75/apiO16OO0zr7uQ+TYHGupAVaAiajsQnaF+ts
pgU0Y4Hm4Sjvq/RiaAVAsu2pvKcjUIAkE4CpGywMxe7s50ZHMoZEDCiihaoBEnh3+jiNGdn6W4aB
MqA3o5Xj8ZczX3/AZgCxE9dfAs9y0oZoEY7GI9No+1XmA+R3ujqQGv1j532IkZ59CGu8AmsllCUx
0t8ePCUZPqohwhgJSIaOid4bA4GNKkQ7rW6R23e2VjejD+Vi6irWTrSHQ4LI28KtjrDGDamN6c2/
FU99z0ZNh4A2HEMCGCFucPstcPBc1iVuNlJ9iiUlmLWUmSjtSveirQZqTeDRHJbniRMqJLvqj0zy
sJwhxreaQ4hIerPJPRpumz06zt64hShDO61cvdvx0lRz98s7zPQjgctDWjsKJNDfPtHMErS2X/4N
BmLvsynIZWgRjZmw02worBzal+c+pJE2G9xqq8TpDJi4cxI22NAS5OZY3IoJYpY6/PGOCOaeDlUr
Y3KCDwBM23ByyfECCuK28fnHoQld0BbG9CrhsHWbXTqhl19GAfPS9vU+AihpE/rf9a8A7v+RYtHg
GE9tc35qJNxK88bMrfI6gCZec4sSCgB9k9di1+aiaRPwOKvlaeSDwfVjlprpkKuzkLGnFPifCX0c
3b4oSvDscsB1lL4/0zWxBHM6mRPEBFGfbc5ui87z16k3f3EIcX3dItKPxzSDueE9XfsN9sp40QaA
H8aN5C5ivCbkqlhVUmrauOA5hLw4EUCz08toLK/W7qnFJJS/gXLX0oKX+UNfjJqgWOz9a1cwSV1Y
zFxF2AMbNY6p24bNB51HVz6sqPP7Cf8tjy0w6Ox9e0eqnXadrlT9wd46svfTAgVyx4kKbCETz+91
a+WTAPkvRcLDcGQhfdz0LKjxxxNflsntrwvxG9koPi8W00KRSi2N5pyQkWhvgp8aEwAvp1v//SC0
RJR/Z2tdacmciv+zVBsRxh4lELNjthjRWd6+FX4Tx6fpIY1iNsI+OIO551RfT7PBR/rq3kgYTxRl
50I27dML5HVYFUP9xBWfRZzA+XZhWesDa4L/QvVKmRy3NnB9dACFcdpLrPdo2auG30JVFbqSn9KF
ELbZRrHgCPnRUZb0g8ofCJizzNK4U1Iu6ic3W8vYn/7r9Fpf6Rja3V9oYB68gBkeVstnRmIbuVfb
Ob84Ma4tMKgE8HMlDjVM0heASdexq75IQ9i4DWAolLMpDrhQ3m3nXh7Ybtw67pMAMex8AHv0ZXCc
AeKnnuvX273ypLKjLAdiwzZWOfzFUjWrG5x94YG3jGD3oc43w9Q75ahpNqzc7jYGnrIdRFFVmeJV
cnzpRFpQIOCN621Fjg9af3RZ3pFXLhy7p2IOeXTWTR1RG9RIxZUSaroXuccKHDMWZw2G3T8+Nof0
0C7MT5uzVfVJ6A3vNvNgKBH9kDphVdabhDDF8EFH0pD/Rj2Jeq69XWL6kuI=
`protect end_protected
