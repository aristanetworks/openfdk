--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
N+uRBpNq49qJHiLipelqiYTjdG/3gkd4SbpasF48hfgfVx4BzEpzmXiIDExdhmo9RQ2hoCMXjOQa
eHP9zpVwKd7FoV9/F81ZkgDkX0pnX/gyHAc5GKTp3vwHFL6YvnysPm2G8ReKt2HopK0R/+l0As9D
NvTdWkNYDoQ+zkSZTKhNxbsQS3+BJJC/H/GBwMcj09+Dz5itrG7ofmMSeK1jUHe43jN9ABR4pV89
ekVuYlhKeDK5lf3cZ1aInJnUbk8+UENmxXsTiUSo3spxd91NyWrboxdrDYMHfM2TvwKteDfAtVPR
9Fss6kBl0aoVL7e9yp5kjbKjjSlUOwnYQieFqg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="SXqgzn4lpMSJ8uh+VB0ORXGkK7DUjtvqzXKbU7YtHgg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
bHDTUAa7OG4DgPcxg0jnULLjCjMS2gXkmFYnRrOElzyDTiiSdOcIc/GZmpu/npubR5OSFMVyBRD8
FJiKj/0GXl+7J9G3UEfh0KatSFVpq/5zGjBrfBAT44ExQJL7cPglmN4IHS5uWeuOy3es5ZnTLI76
lAoORgYTjmxhAbg33KtSkhK4m4NAQQDZOZjeuvhTqreZNeTO1fQNYj3TuNefqttRnNwUE1Aljzch
OdhT0dqX+8gXN3Mx75wQNjgqXmAmLobqTwQd9U7DPt2aOVbsUNbtNuISI6fGyIbRUr4CGlt0ibg9
PlYMn7V/lrDwStbReFGpOOdyDz1dIvwbSoPlPw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="7+j4Xix6Wvw4yIlBa8y76xS6KEtTtTZPMCdKgtQWdIc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2544)
`protect data_block
drfpJuiY8cpvzPgEem0ZtbBbUpYKkupFzvR2YnvCe+9nxWoIwzt7bkUyXGXvB5K5xjC/7NUr9HpW
sp3eQSVJGtGEMbsWwv0yy6DebxDeIMxD+wEJpgBhyVoTvB5i320CordKur+vixRWiZ2t4nAro5Gj
n8DWC5ZGzWL3/hysHGKC+JtZGblrAMjhFBkKw+ZvulCg2TDx0Wm+P6md3tFE+rUel3BZQIRwy+eK
y++gVJOqhbY29SSLnXSjrPnR+0ZPDRHLFIex7wLo6+gABprw/p70bg+Z+mnh4L3XUkH/mEJirvAM
lmt60gCnGiusZC/pyQ1IFZKHa5uUVUFYsQYIfn2QQBKD4m1Tcm9OYI8K0+h6EVM2ouiuiRlrk4q2
/5GIRQNZKDNpP5E7duhozqNL+Y8RL9fLgWr/05tpmHXRz+266pZGjr/68bOHW5+yMMyYzq0QR25d
5gpe4luxMyLYPsZZAD89SBtk/DBny2sICH+nt40hhMGCE/c1lti9KvC7RVEOPrND8BY70VWvf6xV
QFLsrV9fOxAHIfa24tXYdCtqyWAcgm5X7ZOvPdDZLfGKpx7Ag8lEdZjvB/zOhipUh5WtieRM5qQ1
Ev9q8TWoQ6floT14ASwUSqYtMsOy9UoSIiLVJ3EhQsCjyVCjQiQhi1WcuqiNEpOB8PO5RPT3LDRV
pznih6UDi4qINYOXKme54PsSwrjU6bGpu/528k2Av4g48QNp4J0S1WsUcBwG0oOdZwMrUdSb5c0b
s00RlDkvpdsTwtYJickliOhZTfQjhnF64I2uOZ3vkPfcKhmM54nwqXNNB1P6IvCPaV5M5mXqoBaC
tj8uuiUK95K7pB98uWtoykodnzyb5Xt+IVlXWT/uN6jjrW+MKltsGgtSfYCiNafo8ZWkpbN7Zt64
85yHiRpiz9MlHwDXrMMPsZxNxTKZzyD5P+r9vtsqii5XbWmxmBirU8i2mdTNtvBs3MCxLiUoZOL5
7Sx3HnQOiAztaTs+x47QasBKTO5Z5fGxR8iQ9JV5WtDzXqQMkMe4nCnHAW3dkvvi/HpCm1OC+Kh3
FmcKplz50Z140/RHRh4GHWB++3i5qzDMdj/fGRxPKeBlabuUNZu+vvByacIPJ23cZss0Fr/Xnn4S
nWrlVBqohSAc6mztBLJnlaXpIHJRLard8oCE0I1PS2RZBX0fy5Z13u8QMLP06OD9zhuL4KD1k44S
MIhL15+c6VWU6FasCFNuvAH1Bw0/Vln5pLzejmw/TuB1clWiW2mNWB+AGiXK0qf+oi7mBObDcxhT
16gE9iHPg1NH19P3yyb0INCXNOaXl6GwfJlumkMPh4QJn94ZEfcMtrj6juhOZHOMFgRH9/+W1rNR
Bo97VYEg+nAIXE8+s9cAHryJ88BlTTe9TryLx0oVTinh1e+NVCgjsU1/5D7wGm3PBMN/x8GPw/Zz
jp3QtajbYIwC/EWu31EOAM4sKcoPKo/hiacTMpJqWNrcz30QzUuhOW9kk7TjWLIjucFlffqKMO3s
UeFPzRRKy8l7D6U1ZHiZp6dN0oqXfip5ynDsZku6w0mnRlwOcXKBBk+2ir3BHCPRJkCkNnDDanr/
Y234tDY3862BWviB2RTsVr6eRX2CokrEjVQ9rkyXNxQtOCTTp6lWhDeBe/wDW61/Fg9YEW5Xfn3h
iflPso8hFqfBVI/yJ7pOFPUgSsgjxdofU5tmN3JrqslqxUBjvSlQVYLeROYhGFC9FzLk53yBQxIK
IoHTQCunuc6ORurOqHnyMaqstT41M4kYkDEV8iqOE/wZ+4nW1z0QVtYNjCpHLe1kUm+BhHC4v/U+
CPx+lGLzeGxKQUXBLCTrS4O3YUaON6xvsZcSdG1BT1FRAOprqnXTkvfx7ykgJIlQkZtwsvxtY00e
zauvXtGmMSw1J+t63j+P1ZV1bt39EWvIF+0d6KTXWaWa6JTyuGwEO1FOoqz6lTujJuuz9qXOYwmf
jU/f/jsRn42mImtx7WxB1SpNauPycb9xJ7jYsc54UOS5pJLZ1giYTpVigSSgDMWw7VCC7fynHBs9
eKK7ttqanKM49GQyUY+O4Maamc1z4MvYnL77evQhjiiH+opTuzHuXQgubXjqdL9Vu2ax5CBqqIOu
Tx8GW8DYwcbK1jU4GOJ5CpWxXxkqOtIOBEC5VokMJgcu3WwDGmdgZwmnNFwZmGd98X9hGR3rc4ME
cTF9d98jLg8cznNWSH5zs1ZRqf4BFXV0rnL7P0QKmIjSHig6DubWbPzJMLn5SNKE0zdGRtMUhWsP
Mfd3q6wg1aVK2qLUNT3pH51U8aAEQ+fC7QEjBH2CiOO9mhrshLqoYfWpTjQlAblsKALqVk2A0VIi
bmW5xWGJC/veBYSUb03kMgacFrtCm8kmW+orXdKSoBRBYEdwvWT7aEHM3hzKarCFahPYr2YkKwer
W6SwIKyMzh/+quAtGSniNoJBEZa5uFreKP8H8h1waRSrrMd346TkrZkp1To2qIiEe3LhPYTtXkeY
PwpQUsJmp964QPkk+4CzkVbyIysGHF/693YhpVfSZbVOGpuGDvBBhk+HoJDuvtkxS+5lKuwuLpPR
JLdssyBrtHBNekj9YEJG6uPNmaSlzuP0jK0q9Z5VbuNkCqGeAjq8WBvz68DFrANFFg6cQl00PKEN
l1oHWwB5UOQSTsaOWLLfJF+o4cu/zno1aIiRjbfYXVXcPWBVW5iTXNPhFIkVRRkTStYg63UdMgDS
wvisUPKrojZuWx45BNAz26s9QLhIaZ/v3ey/9OXNYoTge+rUWKqwAsXmQbdq0Gqs5b1e2+lOM9SN
bBxKO0quHN8oCmXsQ+ywHVg1j7HA5ihwwtIzyD9Y6C5jALa/htb41KDguDEpNRHXt0wqw/dWkW1w
yycGAPer/JjCTeyyS6ScCEoDXEmgpJjFKVNDKYQESazbWiDW2xBmS5adwFG7ZbXK6NXc7r2SHFZh
os5qSKNIUEn6vYg/zjzPGGB9tTOJZkjLeLEuQlbteYYhkAY6zxHfDtQQhsF1/OiCLDdwha6XW8RO
9CyVf+KAkCg8H3u1GNLA/9RpS1UvXpyZITsh2lCBbconouUsBE0TJUiiV7EnGIAn/clyYFllmAb5
N69sDXXRFy1quOvVF0TUEkti6PLUjnfraR6CRpHbKTDOOOap/4flnG2CIxaTQdWTISjzT7IdKNvI
e8LAhAXJP157j4W3AW5YBoAtZiqyPK+6+b0bbToA+OB9TnbAFDYT3fhwoIimC3ePAMXrPsbkfNLZ
ALVsYg85j/IaAGRXnQ1kGsUuMpR3x/FU7TN5eNbJ3J8T+7c99um1su7vAnWFioifS/QmzVBSbqG3
m1haiuscJlpWw+8OsXKmclpN4HNcqyIlF7L3OkpFR901q1TS
`protect end_protected
