--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
HENC/qV58qqrAcROu4DvEhl823Yangqvt3EVjFFSF6+xwPjWiiF6+/KnnVRcZLX9uAnN0CFHnvJ0
bnPRu7hXVSjM9O38pjhor8IZYWLcodlpyehJKXjsN5HDl0AdCNQiSzB23X0Y1VtCYH6LurisZiU/
q5if8KjwOwJUSobnMXlgV6lG0rW94vrbRLsCT5OKKxS9CXqRXPRQF8wUX31RcGhuD80+21M0jYZl
5f6Y88JgXQqL+6ThIE07Pu1YfijX5DGqiWwYWnV0IkydyYyMhVWBb4lab1qNdPPX9vp1U7w3lj7x
AZx1nEN5Z1bSJtFisscAYoCvdjo4kMovzwLYIQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="gNXaJh2XfPo8pKYxNSndAEnl998ApS7LMI5N6mTF7Jk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
pqi1InwZz2HsS0DmocEKIuZ2VW9I1gYReld4ErIQH0C2kn2yIaPhjG/K/DznCLshfPyKwC86Dnrc
fK0fE0EbqP27A0FquSDp0QkMPHW9qoKZ378EJR9yL3PXHXndX5uIqUC1VcW6Hf9AhvxrDvIBciu1
kfKXX8OEMZJMukPoEkWSwTkZ92S804bsRTw18VcNGXyVY8DibXIkKcdS80wvfwIk0gf3opWls3pk
SyKXBcoZFEO5MXbSIXq8g8rFbMb7wIRVOi9hGIZ15jMQ76ey8r4c8q3LTcrOM1uSUCwnNDsYdEHd
F8Qo3CGP2aVcE7wAay7qTImMFNO3uKG92rw83Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="m5g77CDv7eksjCE8ch91OgpMy0Y+kyTT24/YIZDQrFU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 93168)
`protect data_block
6DoITMfKWAxq0Z8DwWO86frPCRzP2ypj+cLQaNHOXcWe+o1UhO7L9rnmWTDXlJSSF4T9QiRpjhB6
aNrg14hOd+5dqTj5MtEksmqUuW1MKZoE83IpJLvS9Bfo8JNWKyAc/lO6VeEZuHI2pjZoMNZz2XRH
Y1P1Rm81Lvfa094HPZzznsoY3OuUJfHR6eAIjfTibId3DLMZ6vFIpiuAN2VKiEv9GuIkts8gj3vU
mHT8VC1W0U33sm0tbmqpf3++e2yf52mu+g4A1dK5UH2VhD4OjcoIcd8R/5hV2xi3QPyB8Sq+k9uZ
3aVXTHv9cFYKZHIklCglDQzYek23+KeajGC47k4YioaNvEHsurcx+CxVPNsIjKu9Py0ZmWX2j/QS
kjwijBmiDytX1fZVzoE65FYgbUXtv8aXEXbpYayr/4M5J1hUPbZMEyJviKVQuxKrPFAciYVxaA3N
H8Lujt1cZr9GlkIb7TeF6oA5X6K9oKVXHwWulCwU9chb/GO8EC6+/fawLcuAnEowYxDgdjmjqkq+
NGG1ffTRWS7U92UVX66cIPgQUm4DAdEXxhd718Us+t8of3AOdcO0MCwPLE1/8UIzL5Mj8ZLJVV9S
Qa2X0fMlNnxc8o2XYrhyw86HtR6iBX1PNZeH7joe8rQBpdmfuZoxVzQ/hPPYu8tl4j31iOC5GMho
9aZ1zt2dYQ0d2f7FqyinfKzKMlnrh7khc4LPNooxHXdEfGWwv+SJ0PtabrV/LoJ/8NZ+wmmb9zW2
9E/m0zH/J4ZyJr3yDcxoGJwXpRnP204t48IRZnC20FgF+LJWtb5i70QiywwbFd82kGD+uu1aSTEL
B3owMbZEQ1LVIhOSQ+nCT/jkXFlvJSVqCbpj44Vta23b62dFW/PYdhIO8WM9WlqjFq25Emh/UdPt
AarG18W6RdESF4eEsmJORm7ozdt0m0QyUnqmrtLWLHd3its4hrGbu0ayiUpiJfH/v02giOXbg6q+
LI1cml/O3t8JaUEWAehaPYXhKhO1kYtMpRW4x0bNUth708K4im0v6T2vdA9jkPKD5WBUOUixFDxJ
yorIbW8/svWDKhPlinW+ZyeGcIPWQwF9keUvbhLzFfkEovJe6QtvB8egKMfPoRst3mK56pPIWku9
hH7d7Xy6nUVsoBR71fjKgJ642hvtlrZTRaBT6RPe50nOTKcAg3f0VOEVmmkaLGp5X88mWvmszMIG
9F5/nVjww6jvDghCWODIlKPWL6WQi4wiPUDZztpaNmdG1O9/T570s7WZr3a1KAKgJuvYpx3nq4vK
q26uB/nuMGKCMBzIWlLivJq6HVZz6+qzAyxFPkdDw3M/H4SIGnXcPBeAQcVnkgU3s9wkS4ERbi4X
w1MAul0joiBXFSNzyE4op3ZJbnsEkLPy5n3em4eSUZWHTlMpxe3GIA9qCFpGFQFujL0sOk/k9y57
hR2qr0J6olFvoaR2gA3/JPWGc6CW/FWdnaOXEAyCAhH7sdRzKkFNHu6Zjo9WMw4FlazUkNFbImIV
MgFi669i862Hfv3tMHANYyZAbIxSlbhpTYd3e0VkDPgKoDiQBa0mBVM6idFQnrKkAxTlTHGLLR5N
s40vSh4fw+ucjqrop5CRmpoAVecNdsKTVvMo4JwJoI6vEf1ZHBsyfQr+cH280Vq1O61Xn0bRF606
9WcHPjnMu5AtxAILpS5lHxmlYwXNkvCH4UlsbALZSwehkNqRbO4MOAMkZHRp539z1NyhNPQCc4sv
mudVMCIQHDV0HJ6RrDVBhsb/ae3gOM2kHtQicjEtjs3ifn6AGXoISLJklCse14lvURQY+j0i1dNa
o34J9uKGHof9YjgBJ6EnoZXbiIS7lh9KZ2ndU3xAHoKKryljPKN9/P1ehMAhVBE8KvUfXI8RBtN+
er3NA+btBIOTMX4rj25F6fU69k1D3LGFV8XoQuWJkbg2FVIZ+G2tfEUQuo4LybnjDTeQwourrIoR
EERjAVHbltnUZuIsfJGfcf22OYmjq93qFWcQFXA9pnzQ7tD0RW/W2xMSumeUdlX1dT/jPo7+X/uu
qoncis0YDooUDa0dkC0yaUNdtn0a9sPk5kyaZESnqNRQLj/zkXYc+krrm5vis2bjy5qy/wR0qpKQ
CY0RgqdzitPgb9ON40p4LVVjpj6rsuZpdJyyCTmT3rCas8Nppcf9NyJaUfhVTc0cYFjcCgcjwYJ5
sH9q/enQk6EI2tClLUa+WNqBs2nlbQ6f1qxgfCcmJ9kkQq52djv0HA3O0+CMfFvOWIUV0BoeNQZi
UuI4eM7Y6Z/mCU8b8K6vdTMYX70Br9fai9j4PjX1e5k0TZFDMLzu3g0VkFdaUaBpqHsed3WSeuAs
gkGFu4JaBkKBQsHmemzvyQO2dWXsTXdooVm/Wt/v2hYduzXM9auFs5p4AXDHnXaXORCMeNG/mpo1
BRQUY2mEEbeEpE0XPCcZXYgBZrORvm+n+kqpE/NWos9zDP0bchbSCM+o0MnXng9tNJHFXpiuJJ+X
AlsyUncQmo1fm3TFBXE4l6JOOEKakFbngYH0GUQhn/3Qu+0VyP4kvIbXO/27sdzGqfjrJst8NdYE
WJyFeEPndgaqbcRKD3VzoroFJp1sfOO4+3Qruwle1bEV4k1kQRJYdbiQuXkPmjnUPaw0rpvrhYzK
BlmnLnaCQLBiJopvXIv2V3XnT63i0iMYDLlSYXtu61ghBJbYjUP8PeJ67sIamchEA2o0I7tVGvV7
tbVFy57TjDrfRSc1/34JoZZQ0ifRjSlEih4YZc4uxaQ7JXU+O2sk4M+lbtOmnXlThNUlLTHX0gE7
ZPS1Sff2OlOfpPiGw1MBf/1ws2ZhqbMY6YAVuwjXAQJ60Vrp2o8s2wN8ctHF7oqC7kc8ehG4OMgs
GS+HEQ5oPJ7rponW5JTcJ/EWl0rZ66tUUmwIpfSFB73jEHZtxK4Iv6AH4/X2anXFh5nNIr/lq/yf
mJQ8rPTbIGHijNMM5FrQ5IIpbJS12wdBQ/N9mVrIKUXdrLKqYa0I7fUIJA28dJs23Deyd6OaYk+E
G/l2IwmOm2N0UJGA42Onrp85K3NbHb9qIHgFn7Wq8ApU47fQ531RWQq/BPyf7ZfAZErIVd0ApgIf
9pM94iu7QWB1/M+typq0/fCo0j4urJop03TYgRItN6EY61rtjXwlsCNr6JAyoPg5TvfnZZRELKtP
8EEQUFsSIcM5pmW/WLSiMl/ru1pTNfQisnaeZoAPxf2LrB//5ZxYt6uTSuvLRx4b+yASEl3O+PgW
+73QrdPc10zlwDeskUqIxlDixkYPQ7JuBjN/Mu/NABYToKArsLW6dXG0f/8K7wVENWlZjwRgI57t
NmRgDdSaQ5t262Car7Td/RgNuKmz93n0AvFebU8dDcqsYFl/hmPkGBSw/GKWW0cP3DbMQlKJeMBl
LBtgKs9VwcElW0gba/G9r/StH5tEZoSP4u5FMDplRX7+eqwc+bmmmp0uFGUpBdZW75vI0rSiJQFH
fJVlnqKNQ+4ZyWQGjb1pbLtrWmKbTNBgR07WTMbfVELCYmByarc6DhYZExUmDhG8AcgS06BNQgbN
Ww8buEJ27E3f2i/CFX15WZzwBJwnVZfstbxbuqDmj2z5/Dt+V0xf1GDTO+xVbrxFtYx5++2NsOei
ZC+dPtm5SbK9RLD7q3ZGfe5FNS2JCxXNU46YvFlgK64kdrMc3wv7kxfeH7F9qW43DjLnwObKhyb9
nNILHnDMyX9gI4KQFGNDCuGat7G1+maej7ZYSYUGdlbpjaNXHdQP7340CMBs3ja7uD60D8iy1Xgt
ZjP+J8/mIYtGOyv9ok58aVIx0tV4EHLiVc8EvZyPgrvSlb2cGBdVa8ByT+j5ZmQznQ0Lk0SlSHSw
yoZ/1kG+vh2bCBoSN1zInJIJzRlbQn72/cj+QABMXam3ra+9OzNL8I3ZvHoFOHfe4DN955S3YBED
0VrI89tS9Jxw5bfreG8DerXezvtVc5tXR4ST4wueUnUhwZLkaxSRHsDcKM+EufATQDpq4hDrznKz
Gby2lojeETF2xVvJoj6v5cbS8NtDwB04uUr4CQwPTW2mKgAbyidMTu+xVf8ogOaBraM1RgYDBWSH
OUvYLl1Q+Rc3RulKdADcuacEZt4hmEt8YY3bK1eOHrpmJQwpUDRmnRZWqz+ZrKrzqzqlZIaAtUnx
/n8IPmeVay65KB5UKy3m6DL5oIe/fCvFKv2ds9RsZNMLtQ9WYYEfJvJ66Yt8/etkc/ma/GJa/QdN
Yhhaacz1QEzEjscajyU3pgICAA+NCnkWL0pOCVcq1H9T/Ro8IglOU2WtOSi8oC71JobmvvX3KxFP
dMF61WCCZeSPCM0PRWmNLrhW6bEyaYOm8fFLy6jThqf+YJ6ujQ6tSzXwYfsku5Gynsrc5HoHPzk0
VAQtVB6mPcsRsjnqxb06AFjNWrmoYY/hzsDlg/AWErI1ORFjZxDCrZijBr+Z4FOlvSIxErMbGGt2
I0j53PK2skcT9vxzuPsY4WnsfUZG/wDD/g/Z7jB3DxmjDLZazOWDC0wDrmhAgfm08w+PSBCV7gCx
xc/tUKDaGpzj9Ko7Pqlp8biuIkZSEk6DIjCVd7SBOPzE/jdKem8f44tR9l40nIkWuqee73ER7i09
CnhEhBBhOHj5KKzvjYLTiFZzgPxfe3BlYbqR0jSI5xrVCZ1jGjwk+R+QVtMrL+DTnsUJX773RnKN
nCLzK94EG2Quzf/g1PmgCpKonmYbfQqjNbgLZrdZBxHS91sBVKYj0dky2GK/V8LUl2iYLwQwozjG
QKo2xwCpPiI8d6VyzmnuiG3DOsdAj2UK7LDQEPKiujRQ8KHbKxbWQTZfi+w8x2x29pXFxlKau3/p
0C4Or7xEFJ/n2HhPUOJhPWcp8gAhNZkZO04LbdeYNLHPZ8h2cLGkG/koMuFO6l1BhYpoU+8qgOgV
0BbgN0ybPXa92WUoODDIC2A+x3KItOVotDB+P749LJgUTH/2H7YI+g6+LlX/xj7W7YZchzs04ssQ
ZxYR4CzjWO1bd4U8vfyOCG2XqdV8V08hAS6o3mymymIA1woC/lBFqLAFkfa+vZJ4Epx4cjvs5NFN
qntvi25GMJ8l5UlJHOOqRXf97W3x92P/GrQiukGJ2C1EgVbwQvXFXHYMFl+7yFndLJV5TDu6jGFE
z5xmY13RNWishEyUQ3CzS2FmIJQL5Sgd/Ah1c37kf9oltocbZ05KOid29uZCN+HpRwB3UXuYKm0R
GzrXIhkekDQ+64m2bufJ/rKCb4Ys3ESYBaAKFCaJyGfzfJB4HUmUjgE13K0Tkj0ZVBsUtBdgXcKZ
zl96p321zy5p4Uh4WpBtYUtJC2bHQ6W3hIi/cGlwkAgG6veXJmSNO+TqwuoIijhLt38+lpe1Hz+v
/bCrCAaQV5B4MiQ1i0JSbwxMGFLnsrZWBk+mfdoijGrHvF08qjkwkH2tSbvrkJ8BlTEuOZtcRLBv
/X6MKCLKpi1QFovCiZovObHOJSNgl+VwbaZ70ES/4xcx0ZK/xwIhGnWu+eQb/WFeclekipU9Cr0b
6itDfC00qDshcEf1W3gR1BOBj7cUP+QyYY5lpdBRaVEr/5vDaXfvYILTSAnx+hInAckVdr8pZEZS
PwnOcI7AFh0eb/VFYpMMhSEVKPtGSvZfS6poCmAsM9LsB0SIdN/glDxQXLP1hQVX6Z7r9TroGJvF
iB1KPuFvreLT9o0qF4xQa7vyfZ+ozQg0nXc6c6+azWrZ0YpS/FS8OXHbdI5bU6+ISC5+iyxtKavJ
bGqSQJH2cZGhYyalB3Dyogc1oM/yCtrGRt9sIxdRzDZNZf/uhRzMFt2pgKgDossrzkCNkA/M/Hks
Kr1OitslFemMVJWwP/+tsJt26ZeIboHkhSNnCbXta9r1fyjjC6oOvokWkhVZQPfwEoFDqH2F9Jtt
Uro6lInSYZG+rpUsj2pd15jceIemYZb6wRuxaQJ9g/ngLdQwgyxdUdbeZXBDF2BI5scRUT60aXfP
UzKzo5Xi7DpYg4POMzSSaflr5S/oHqizr/YhK/dnmQFdxBepf6YkuvcCI6RrZLHsXj+mcWSJ1/7r
XpNCoGK1V5LSoAmQz2olu7Y6A3cJ5KJXGneb/pQ414Qh1TnyftipOh2iS3trOfbWr59HInIhiga0
MAcO2/XJvRbzwvsBlADyWoprP/w9OUHMz/R8zotbruJYl8NZP6x1Qwt/WoJM6a0ZL67AIvCY2C3C
Tu/sLZJGcgS8+LsucLQWxFW+5txdBXPDCZ0SL27+uLwkcjeGo6QB8bMbR8mjwSw8mo1TIfHPMh9i
vReHf1ZYaXDBgveJLFjrao6j6DqRZr0uXw/w+vkPvStduOOFRvcjfqjNLHxIC8+pQrmkmAG7fP1F
YEBirzOqOEnSHdysZ4mo9D+sCkPGACBADr7OzBeNvGf64hHfvNXGMIf1C+vf4/j/Os5mjQkszzfT
KDnp/4nXHZdREWTiLimSFMLQBZ1USJADELx3xCv/Cz08y4SNnz4IGqbLW9YHCp/Nm4E7cm/Nm2nE
SB0riE9GzQMNIyYSh7ECrrMMaTh/naSxgpLSVZCL6NgHKm8SONyFXfc1+wu3N/rkdfEKH3mWteYT
vYxkwpBEU8Bgt8Krt1BTVXe9+ytpvJAgxs9lPi1BQkcrWidusad75YZlXIxT1KRp0AVdAnMcO2PN
2INAcwSUOsVePNrXWzifd39VvDMQxDPTYRFj5HTyZliUq05UqwBF+1LyRQhHJ2y6JAZtCpEZJ0ac
HSeUDODpiq73q6SC8wbTSU9PkRxyO3TUqKIQLlqEZNs7GRHeSmr+l7j3vtlz4qHuGo3QSxt4ulus
8aEIic2zfZbmtGeOPqxhitQ8oczi9kSMtFzaR56CsbuxnspwQBAW3KG/cpAi6uOqGY/NGSFMXuuj
23DlQEGj98ngfb42WAXxZarnLTXDlGPLSau9jMLiX8G3ClI/JvK6v7OVOfBls/TJB0T4wK79RdCe
JwRQx/puH66h9CRHK6seQie7YUvZVShsRW4igh2fyoUMGXeEXJLn+qmPeYDynALyi4whV+86GRkG
HmCFgjzSUZaSCYs6w7iIjXSUITIm9xpHQynSjS6s5LeoTMDHGEnD1PL1XJ4P5BwNzlPY/wCHI5io
a6eBKfldKKpmNiHVWQmGIP+qWM+1mYvA4kb2Ib2+10B/iuI9WNYZx9jYC4QLMty9Zl6rHjqOS7NQ
/hIMP800PjusYT+DRaFpxjEIMKim5sVx/QjTuXneLFEBzqlt/GZEc8noy1LdEbUzYPdjmhOii/iH
wC737rK2MPzPH1QNz7P4e3crLeUldPRNxWBNC/5O+cCKQ8fUIwukNsTBqvKsJiV/L0BfxOwEx9xA
DnmC3rjxGxQPCgIBxJYpiL613UKLiFgb/Vhj09MuHXMQM5bzYxTzh6uHMxR7zMhEg8LLluGIiXsT
s636bc9PVy3vrkF/lzvbCXH8QSEC+JOXelYbcRa9ZPRlXgc7ZNlXrY5FEZVxrrjjg0/SuuUlijXU
GLqIToex1eG3wMbKT5xh+5/fJPSZMlFD22znK9VrjePwBZDeRTcSyClpwYXMZrmQtjRI3JwIarhp
UVBJM4oYCfFEfAUO6XiAqSyvFMPrOSohdK7eYNfdfF5OEo3F51QYCFDb6AWMxTPDWCs64eU7w8kp
ZPwziy98lKJts2Z8/Fsk1VmI4/OvebuTlelLCOVXkaXrHJiMo6662JtnbgMJzU9CGFl/duTm2t7e
JkgFTI9bqMPdqyVk5dMtyl3NTHAyUFqy0i9wbbYBcPZHiL+HTaW3XQ88LfombWAqKvxbFC3u8XrT
2SbDrWUPbqaoytgtFTHeQVDSqg4XbkGWx6wIUnxwRspsdM14w+8BQvZ+nKR25LxRHxL74H3savsk
XskTab6VQHYO+rfXrpXhWIK753K3Cj2ZuLiD2+mp/kDy7V6dgNC/WDwxfrZFpqxsfC1BCx1IFNq7
kCKFMmqpaIzB8c2R56OqXdIdFxwoKqs1O0Xr7egtFIxiN5MOKIgDqhMQgxbiq9QtvBAIcposE6Kb
eP83BjKDzsHZ48hRN2qRuDbj4naJwsen0KxgcsWMPRwOlTc8GY7grEVmEohctRLVXSi5eV4vqgsk
EiQDE/aLd1IpBVEiUYtuD2+0wQs5eZ4+XcW/ogiLirJIgXuqwa3GRqW4xljIp501H7vNci/qYyuC
i5Dz0gbISTN5ZCNt+mbp44zwM/Oae3a33uiobe2lXPI0Udr0tCpKIpqs4qjX0rbUaa+bOk5n4rja
pssz6MdNHwAX4Jp9tqdUVvacQW03JHMp4bCTSF6bEmPDHT0d0ckw84CojPcBNE9NHGAW7iIlezn3
4Gy0oXEJ4viGJpkb3Yf6+fopUgfqW3nassSaWdZHOhPrRi1A3MUv88nVqP0/fkjwc92UyqSTOVB6
ZXXYFaZALvwklk84fxgC4bEPUQ8OUmQpMDnTxImMaou7fvUe16LxxwyDlXfnElXdyLEEjJ9WlsDk
h3AxLlr82o3kq3e/TXzWhpRSM6dyTd1ntQ5wjR/afaqlQuhuLLfXad9hotAc/ZBolmJqqsxMUSpL
glReJJvBxuljmN9AHH50biNLO0FjKC74tNC4u6w+ogSVXXT0Xq+66dZe5tbHrTvx7ePw6c5CUViW
NXo4I7DybMurmF7omLPRGFusWWR7I2OelCHy3ySRz/eh9HhyCNFF46JrTo6q7I7ekIHEtGbyzJCD
Yy6ktdVXqV5QjfSs2GWtGbThxvvJsvzNaPXe7cBxnzBijZOO3Fxz2ySSRExZDrKYdasPKvI5F6+P
OyCJwLJFPvXHtzmJRGAb56tj4VfSwDAs8eL5qhfTZFcsTz5y+PkpUcrJf4YUQbUmuX33CchhXzUd
86hh/zHKa9gEvrulisRlEHREjCZToGsiib9OabZtyGO6FmtLyT3ZptolTqNw9dwWvzfcq/h1hI9i
sdcQqDXtqZtoYkSaX/AXuW+D9WHHfaY6ZrQvB4OUZXP20NXPGotWIEAXKTTcYYuu6DCPiyigr8Am
pzgEze4hgQJtuMkjGY9wifevCSyTVg5nrN732g4McMb5JbY+LxYNUbD1NG1ZxiVOGiGYlaYaoc9a
bKI1Cv9WuUOBE0V4ZjcDlsWpDbwYEe+nOVsXY0up71x3Kwc0ncqiJHdANbT/koDxDZNWK7Y0wzhw
9On4bUuqbDqKPxQDLepi+HCD9IyghRXQBP2hp8O8fPSGNRk7fuKLghv28wLZLreHUiOa/LPP9E3N
a56pwHpF77oo6dYGBzY0rSHYkx3FtiOURU3S3X1Wn7RDT6iZhKPRu4Gg1saJKMXIC+pyOvakrEuU
Vk5g499nJLkpdBS3H8RM9viyq3VqbK1CdbdPtpFqSzPveTHXcOtiRnggDFeLfJZ7GomdmciW5CwX
A7hAszhPzkviYg9Yhl/csZfauobviDXV8+SQqJts/V4CYCERvxUyv6KNLXb0BYlJJfIyKOI+mq5i
dKtAf5lXjhCtri/DQ1X7eB5r4By+QEXwW3J7droVBekGQHwG0wPb1hXpfFsnTGBvNkLIcOHrO8pw
3mqf+tlQvJ3l/ZyJ9rTUpQRio8GebDyy6zRUfQFfctGMpKQIwcSsNyFfYi2LW6N6ndlDPZ4rk6vq
4jFNT/J/SvrcPnbyjoymVfRVA9j8FPZ21iaLPGChfhYkiHMetGZiz3nWyYHDF9gDzA+XJOmHaGE9
btwXSk7XB7K5aKspViH52l0wTyLtpZzu01OYROeC60JlNJYTxigOdt9TuAnfEXK5jnU77iGHN9sT
e1Vgi/GW6KFUjeRyHFLZjZyDGfvcRC8uIrUwnXYMJaQCqKViQVAZPeSFo10V4Gp2u+e07pqPaJRN
7teds2Yjuv9KuNfEbl5unwpmsOTWWNVFEX78w3zWEB2Cf4v4SwjY1256pAsywquAaymPN/nbqRg5
vHJACOZqa26OThNIvhfvpW3P8jgQV4hTA89GIR3Oda48nSZrIzBx3ESOYsa+VuEi9hvA/o0xYnCi
VFPbzlOgmd8uWuljn6LbMHwcA/2SbmK9s5fT0mEldJ8/CXDA/sxsjKBOhZg+EUWMwCgQJPivKqaO
lI0+SxmNyWxaV7VaR91/ZSq1Gm/zt+MU2F+sxHDXZbbeMpnJwZwEjh0VosWBa2AQu1hsOa67JPyu
aZIIxlrZaUPvnBBG/A9ocUWcMvtbOuaaHagLogON/UGQhmUYJp4oTsqsGvT0iMXmpjrnl0pGJHuG
Xo/ndEXRPP9LrSDSq4GwsHn89j6VkSj7qCQKUfaoxA/SkWq/kJNvmcLXbgJ9Vl2xYpf2wasPHAan
YptaUqUUEgJhCc0v9x/UYQphpj/uru1NrKdjZEjhvxaZhvJ0GUBV3pSQtjeiRvcWKPDEk97Eeaz1
8AFgS1TJfr1hDvjeqTFSTTXrCnZkXZJXKTF1CHzGPJ1H6RsH1P/yb1wWs63Wnw3mxbDh/eps5DM0
QIiCCGvtupS4yMNgg6F0GqRvqRjQaPpxVWLcjboC1ZK9lHEAZxE3CQUDBUnTgv5tKfG2h/A2D05X
E9QHKEQp4rQrX9ZdGyM0M2SNYlwuWpARHIt02r+URer1Yeyco9lbo//d9ZSbqYkiEAYYtT5ovk2h
H2y+tCeqxK4dQF/sQwboqL/hHXbG1F4MGCKByACIuqOvnmlz93fj8+FcLUntaCO3AgOZNLJrO7Gc
jD+oGMqYYrYxOlIKIoCTDdvcwcxbBYwOQzkKySbYZdR+lecnfRMaMRVN93lMvEsgEQ8VMu1K8U8m
sxqMKkE5gkjZxI3+EduyGLxDmD5I/MLsGnEYG/0WKMElzrpcap/8haqT/5C3my7uPmSwBoLQYcyz
BHtw6t7QaIcCcqdQta4Brj5heBbRNsL8gMFPvvAKs5pPk+Nqy3ojpNB8JCd3RQ2jBVfGYYkdmuvv
FgXOba/c+2TY35v3vIRKxQiUeYPCAJ6PpNs3DU/7Kyit3EOKQlhzT4uqy1mdGbG5A30K2bupnO/y
MZtBYpRv27/aeT+QqjUuVLuYwc3jCCCPvxJ5dbmxBPVfgPALWevlsZQjbcFGAK1gAla2luTNiGlz
H52DmiMZjhpy20XCRSsgKu79XVPK0ZXsj239JNWp+ZM87JkawLJ2COFCk67iJ5Etxc6Gtz2raOrH
hi2DHpBnzPIvXcu4sgacWx/eQXdDMGMYlLJvHzLC5IbKWDdT2cHlt1eXEFLgHVORCRZw3br8bPx+
zCv7eea24GPwwvDTL55e5TJ0rPr4QWbUXai/QELhYZXL9r1MQ75QWNwJgFZEkpwuen/dGUODaN6a
HsdJop7hpUff6tdUOO7LvE5zEbV13IDVVyCusQ62E4VrPteVTFJhGKosXOu0HRMuioDDn/e5Hb9j
7zovzsLzbh2T+ffxErJv/m6nwrKXzaAtzxIoo2lrcJenS2Lf8pF74oqZXnDE/Cesz86LhlNnetbn
Y54em63EzH2GK1FiymR2J3gA2B1JE0nBUsjTYXoexw5ged9ZGcNYgCKijRnee3rfS6zZvjsg3XNK
0vTfQLRgKGtpDC8TKca9+VwcV1seJkEtucetMgzLfzI75KJUjcW/siKnOgj3g8FjbJ+Acw31hf7D
dCRUzqMlWTzRYJIebV7JULpdoPBI+rg1DmE9guf6y2bp57m1OAXWbVsN8pa3JDsiUEf6+bQHTqAL
NzA4cMErfQqkXBehmH6xcLuV7abo1JmljijgyuU4VlnJehGs/1HJwZBsiSIV53+ZWj+Z/1mm/nA+
yOBkr0UWVaBzl61sUQ2+He6trRaI1XiBKZHQoK/F35UqSlFkDITW2DN4XcKq/AsJdRud8R4PlflG
/xzRY9Qdua33f5TeisILylEHtg6YW0dL66uBZB0wS2RUUQKxLaX6IyqfiiKO23CMGueg5aFecEQZ
4XUc4foIVpSjoET+i2/Opt8tjnmcRvQozQjzJIEOXC/b1qFC9MIRMyQG4rttSlDepUYqh0vqirTd
NX2MMYR4q5GpQY+ooA/vs50bBxUK5EY6Mj/XRO38fYCvIgqtvBpiY64NLLCOzicol/r8Xg0yjHfE
lRe4thqeEJbEb5aYLuZ+OzYhIa0RDaPz/xO2IiDSxW8YaPfGVE7IBqtTkjBBsIJGr5o1QAmNYvAE
FXYoTJEzwjYTiABexLogKW2FBUqrZDVKyf2/OC2xGuOoAeag8YvKli82FEWtpsqT3boAb1gvnTzE
Rp9s3lDRNREW9bzi4JJdkVF9ia7TNtTzyKnH1Bb8RXhVwUqN6uTvtFKpuqTG/Cs1zqX3DhuAXRnz
oWTDj3XOaBTrxrYeP2rnRAEh+3mK6xdZ+Cqwkq24b1xY8Ugo4J+EFN/BB/rsPQcweXQpjdAdqUcV
tMjMKG5yXIQsW7yUFmpPvDO7Ze/gGeaT1cyoXNWDgK4jJquHYCHIky8p2wKegJoGiqUkr6KZc0IA
ngIkA1DbrzYlEsLhwIOzmEHckeUCczGR22C17jVIjOVbBRNh0aDHN7mPejSGg32US2FkUS3K6Qc6
H9WnnNtqtyrUEHBawO7pDshgVXtgP3x+7yrEjbTkzVAZvEgdvr9FFVc/KHpAVhdTMrliCFDpe1Sh
8A4/JFahQXUCCkaR+PgktrMJcZtTnfJ5lzKBIff1eU8n4cIrfx48FnW6m+RyLNsl/ja9Tw63rT1j
AzLkOSNLj2V7QsxQegb/GtGIDub7DoE53fd8wOxyPr6i9YxsRhyG2YKfJ224SzgyQcI4eMCRzno2
eKf/j/Y9RrSZ6yjeKIghROq1Xm58oX7bi4oiIfPP/g4HWmhrpwJ6vp6TRi1mlKvlNjd/He/wuS5E
nvimmg3bnTMeeGkdvY54SWSI5Hy5uN1y6EeTwBqGVPqQcBq3g0OSH7aeubYKGOF05M3U1k6JqbZF
Qx5WRY5+Le6eJg5jy82YKjVlTNpTjKGJhz4t6qwP0PPHAR2u67xGJFsD7hDdFFMrpxrS3bNqFOWD
xF5CA3EGPIA5DeLL0zDKJu0+6ki90EtfXVxjpnbOKip1mjPJYc8Gh+lOglTBhGhRaWb8C7Q4ScJk
gI7JYVcrLh7QyU5gWAOv4BqPYD9UY5awvmVqjTqusB3zZhFpVDop/48ZYL37QKmQE8awyRjtmwaA
2ja0Hl8tJzg1AwnTWQzWjE37TBS6qcQ6tYnGCU/CwmjzDu5PI0OxOO0ZGF0YYoZXb1GqYPgK5yVd
oWLxpqfu0fklUL25C6waUFL+PZwxqmnwVLudrqH/riNaWkjQpoq+/pRqv0YxH3CAo+K5mr5YN3Ob
ec2AL2u/JDH2ZNXTwsZS95go/3BnTdycygNgiXUtDlP0LOmIw/OyRm84yuavrFtEzpDSQLKNeOCz
1PNsSoRjbQtI3cLUEgLn4oRWmLaJVgyWDKnmCA6OWzRN0afvz8v2VbDjjrASzElmOqpZbgR3w2lM
JLBFoXfcpZedyu5MAgKmn3m37WGlFl7/pPnC5YZx62l0HUTYy9thjovSxn+iS+JlVRGoHqScos2p
OKiRsSXJhu1bcDBeGtCvekAssQgiJ5u+VCj6tCpDRtdlBSgIe3B+u05zT59jsAgG9tjjIIMyj4Td
OU/q8WAiGVw046tFVMrtZQCUJhPN4ugNG5ZH6ueY5V4YD1sZWDRVrYtoUoo34bAlrDOeCZ8O0EeK
KmLZBM9FvsnY6o9wc/IHQJRMbJIOQCbwjR89tq9JWuxDpaQXNcB0WK6McmcbBShDdWXWr2GUHy1Q
MxBBfAKeYDqA52VvSNO1pDXa6veLweush/afF+APEkPYTbMNalzVrlBQecRynN3vcER7hhou+J9u
ljv1oXzdxEpR7NIcJn69XbkQcxkoXcFXOY9AZPp1W1aYenoI9wb7Q+eZyAeSHzDqO+hAZ0A28jc1
WIqnF0eny5wML4L0N/kN6HsWQ3ribtv7qACCD0LiPc7idr/IdGFCP4TA7hasu3Ve2Tn8vTgiZ76H
LICMBhevkgQI+PhxXUFEqxIt0BFhqp56hpScv+iHm8zm8I3hDISTxeDSn3dhg51Kkp7hySd5VcQn
9zNi6HZoJVNAGFkcpfqB41ScSVuxTMesQrVCdV6JpdaJhm2BD16vHD+wn7rXRkvWYJemlOelBJZZ
MPaw31zm6KOCdpXjD1uEWkcIayE7K5FndTTGJUFnXG8Z5JSwoBIc1p6b8oHtq0+YfBPp5RtZbPkA
KMfV1l2FMiuFncV9G86ugAVKVZw93ygGZzyjh6XzNYOv/3aDTB7zJyIV/Dt5bOnCLeTVcAzbsok+
DfkAFbaRuY1wjij2Wq+IyJVvTw/KV1+bw7J8VjGxWi5ShZQNVoXW8z39qhgOhH7V4m3IEH/jJyEQ
+hft0RQJijYaAifPStjEiTpRyfDzPgoPye4+6NSSxXv7Gpdho7ZW/XnfPG0U7DCT9yPCb9xQ4e0i
RVM+iAgEGfJqEKfiRZpjxpXifWtAOXbz717emJT9iPZ3K5k8/8jrG6T6uvhUfcqQkcSOOc1E75es
b/uWBaQUhTSFTFFP8Rqt5aeY1yTA2Fk87a0c/nsjoDL0H2C8tqxHqhIch/vReUv49jl6+VCHRkKM
6rnQBlR9BDkfdQdxSUi82JTlXyJy0DCQXFCXVrJ4zcRZj12JhyGGH0IyB7KFqrYDqe3bbCAfkU8i
SGoXzeiAZgwj/bGVHLEqG9Einr1Apcuwh5YanImBi1RWhD15b0Nq82HMqcmEUP2OHMYR9Iyb2nHK
snW+n74lNzbp9Pu6B/rllMetkQNgtI9EGH+LZ/zqHI8W85j1ew181Jqk0JAG1rUqOOx4+giIRWfw
ksOzNNEimMaqLFaVW0Fr4mltkQ3/c81qrwXy/y3yCNHgaW04a58hND+EW1h8umTABmOZIb0TG2fV
Q+jxWY/COr0H+j+rHVtO0BOw7kro/1RQTIImjq19QAlTKLqnsFJpCgLhsQHFjYyRTqOr058PLV0j
x3jIA99mUauy+TEwWjcDSQJeggmKAo5oIfnxQw48d75re6FD3YIO2IvbTqba4DQk49i9cazVDv8i
qJyBsnVbLKz2Ykqxv7Wbs7nNH114NXPVNsSnndW/LDeoVJhcMrdLdfR1ANdINxNhzZzvvpMCN+y6
nEue9BpdSY95z5Hcg4bTBtwomAFvjaO8sVijpBGydeqcsPhIO6QZzscz1mBU1B3l0RL0obimX4Ww
Xl/9hDNffreDneDotWG9qsEB8OQm2Hgcfopfs8iHkNMUxRA8pkKcIqvhxLEpVOsxDrXEptljiVNo
vxTF+j/dzHf/A9siDHRl2GQAn9giUNooIKIbynJ7Z5K4AIQXKCg7ovJ33N+ApFnuX3MrQIS/GAwN
MHmvriwaLRJv/4xwTmS7DdCUMDumkoiDpbDz4GC097tBZXoiw+2TWwi82ediq/UXyyirr576+qKW
MP/Vt44nVJ5l8XUVlSgEUDrzWsJPWsuZqz1f0Lodb/nuFI3Ju+w5ioBMnnGDpmn4BNDf13UGB3kC
36l56la/0fDoYK2Sb9SC3y0T1JJkUW6DFnV4fHwylx3qpzKC3up3ay2q2t17Tx/o/iLLyiak5zpN
sa/UJDdMDQ4Ljgreh0eEvWmG2xQ2lmQdQa6TAoVcg3w/f91MI0tAT2cGRidNknoioEkotWOiXJ78
xKZyinzrEmn7/DiI0iQ/jeFfel6tpxKNDhYXfVE1aYExiemXtgZfTqXbpj91sRRgQ2AtC6NSJKaf
JMXR9WE97seIXvN6p4vtm21xNVr3GHwvTdup72i+s44uWalxHl8Q4rq7nXpizAXXKxKxaLq5eYHq
+UbJx8S/aniBcwzFqCJ8Q/VjIpDKgqBbb56VF9DQ4ruIBnpY5RufFr9SCsbSDIkkAooMTVJo+ltp
yPA0qzBPPDYLZ124/rsZPDxCMu7DI6y04EmLB7g4TnKSA+DNzaXTkAnt/NpyneeVBDnAjuZ1Ckx1
69oxjtTfclh9OTIwKeLiqU/b9cFe63Jqi/K/tmRxrklbrSq10mjBxZCVZnLxbjpjor+Dv2iOI5Ig
Css4+nyJisDC6x7JrYnCCqr2uVbst5ss9SleTneLSSu+zjRB4F/g8TyQ6l50R9vSeY1Ne4h7OJwZ
0W8r0X3FTO+ob3lAYnycOQx6zqCAdt+EJicpHn/ZZrFZf/qsrOyyvQrG9uqIlKvsOv6ZfQ/s+S5g
3LhgyZ0mz+QuP+9sIk77iI6Nnswdn5tbXkPm6f6sTG38TObXVq9616sxCJIH+alg+C+sTdkvcClA
TD3JfnKfOvGSeUJKDGbBvO9roJlzTPyIdC8B8n3gGA1Nh5cWOeDXBvDVwHTC0cnpZVxoIaX2g1sG
Q4qMETJgmwxAsxgXOUbEbgNkVgStm1YyKPG5Qa+Fqfdms9Qc4lROiBk+DlCedlNY7FJf1/0CNxOr
MhcQvFOAw6S5wKKyGEQvlV9tQ3tu+Xe8uT8EAcvLKQAI+psdyfAcIouyNA6Kr4bWR5dwJjzUzO5e
zzd5n1bVYE02zw6P2Xi686vQJcLico5F0Gf3UzC6diVJ3VNzNOBzn0yzJpqMc+EcHb8GFcZ6QCZJ
rOLLoWdvKKzT/QdLTfB4dil7oV8y32WCtvgUOH9w/fvm9tJU2MjNvWdZbpvZb2E0hxTSXqirm3Dk
wCzsaRGuT2iGItkArI4sKnYxWzOIndgH9C1DzSWjMoGNXMkBf5IBa/5EF6b5yEuZsA3TUqwSODsQ
b+KseuFLmZGKBh+E/Zu5+Gje9d+vk/L3NSLWoL0HhcSDYQ2ijOg71T3UiBgaObBiFvK/rYkPoTY7
nHDfu2DLxrU1jOaKQYyERpErlf0yKItKYWm+w99nMpRwJulNRwprh19J5LJ3UktX5wesvxjlxfeR
rQsDVXQMH3BabYJssFZmkVc7BHltIN//lMq2ujbwVvUgo9s/uiSnBbKdeDiyCsYOxdtg6jn4+5y+
O/EWKTd9xTX+bOanCuHtqvnyNPktObddAIv7dhdjjqJhUROeN83HBSmAoImifmEqkiQ4QdiaHnoQ
OqO10OZRPpFr6b0G1lSTw3UL3zsxbVAjjyfMPZPAsC6TNFu4InLSiufQ1lWByX7/aluhSnarV7Jm
FaZdwnxXPZ712gOJq486aZRnKuUfJ27o2eTL2v5qwBbFNzCXvc5EB3XLGQbWpFUYAPTI2iucw4JY
TYpuLVbldvnRtFUhsllwRL0iPK2Y2Q6tbxAg6AzMgjd/+2ujk/NTvppJdQTRFMsQn1tm23hY791j
Lt2rnCRCXiq5MW2s+aRIgscZl6mAGYJ7NgdStv0pQZ5KYb6PKbCj9JYNAcZM6XYaOmRqPmTJY8EN
7X2bakSt5B7/PHGk6dWdMSCoj5rYwXaq2bYdvdGoMA3PDS/MGipPnEinmv0ky2MELnJRmf4bFeEB
2yTeKWvW6W9JWf6i1WOyzXs8J6DWT0nSojM3EQvEtYb3h2eP+AWi2B0+nw/wSTrt/kdKy8FZoy2I
OKL3pm/OuxqlYr3nkL5D/xCMtuxKuacnau4sHCLpmCFRfgCE24ab9gWuT52ditBeLAQMjs1VZDNF
4w4NmISEYKJWGYKjW5o9pNq+p05PTcfO1na6dpP6/KSbK88hVlBw26ebi1uZkcJxwPiS/YcNu2Eu
FklezEaXOxAmEyjKy/c2CBEe8Qi3e0CEyD7PVIsR6VQB5U9XxcAglVSjfJmyK3BPrMhoEeQlhHsC
uTgIFhSsCVySLPOhNhOwhXYvWS6t1r4U1inpeZwdmisWrS4jQvqRWR81G1ulDPfm7kP2zxBDlB2S
hEwrrDMhnf7bad/UzWkDJZXS7SuAUJPGt6vjLjYyVsV9MM/tnoUmms237CrAyXStKvEqHjFNZXbj
Xrhu0jvM8Po8xmu+MX8i1Rbvgyx29HxHoB6be9ZVF2XQfxAytiDVpzBDRNBjxUuYL9WSNVOiQpe+
13MiZSXoKCnY92Ik5P1S9Tw2HW4hEK2IOVlONbCxDX7pfqeOy6rTA6By2/DdBRitt9GKUC9haXGM
4K8YhJbemFAPfn9XpHReFjSNyCcieOr3Iht0dvmgTF+UWz3enNQWMwy/1L8ilVAiYn0VsNyMKn2a
u1mzMbrPke898vEmELm+1OvNMTpsuKlC8AChBt4vzXsIqQllcAB0NWgV7e0PtpmYa/1zilnTOA78
qmTkvNvLoraO6lZyLVpmifqxQMjfKGjoY0SuUri2mNHEOfnI0P7o0SIqAmxdoqq/UY5Swuv56Ic9
oGobuoSzEgLIsrPx397481sWXWZGtpBAtYrKWYk0oh2NT4lxji8gkttTcDjuRBU5SsEsekD16f/g
9bmoP4HywFggdJ8zcmg2j32EdV6M0U5rEf1KMVYlKqEGJCHgu97l36cLU+F6bsqHQSq4YGAbqdtc
jsm/3NmwZkBXePHNW7RoOE4hpKAFkGTQXU5Lv43bHlQEa8Ii+auRzXJZ4mbpFFyg1AEDDMWSVdMZ
QmxXqAiW/iOlzpqkxwMnQ8zoB9Ca3RC61r5nRHXWaN8junZTxfddeqpLaRfQPZk+mbYz97acMq/y
zi0gweHn2xJo4fB5EkU4EYUdOKl95HSo63jqtKjxUvy916d7iAm6PXs0kHGaDC9W/AHY2xoD0irm
FQtTnfUh5SeEEBpw2K+bJMT6gfWptzJ8/UFM3P7R0/eECczRrQW1j1CV6s/x5t3ipUO+HLtPhYDy
2sDHpH4ukLp4WZI8wnMOsyapIg6NUd7JSyMTJiTPRaI1kES0jsIrNMKSLgCq4IPnG1KwJQpppRqe
h8II6VRJwro2Mi+zXpus5EzQmMD5QkXt1hHNlWEvoLD5tpnu7eFb29TTv2w7HxhEimMBhEJYbZ2j
hhQ2mZQJ0je22lgylWNhQPOGIgsZdbYpznqFq/F+U0JFiVd/6/KkRhMNQ81HMA8p2ugSo+v7oWij
yzFx3tpgyX8DGCCBLNgZpnRzSCTIGQqD9u5wIuc8MEBdLBqQxZUYm+FOB2heZxIbrqQsHiwESTf/
DqSsW/f1JLSY8HysiMVZcnxZPp5FNa37HsybGyAQbqME/KxkM/+TDSednwtrwU42s+PPs7w1rvbn
Ncq75aIjrzX+i/45JUjeBpXKpEFeY9aPUegS9jMyLOblY4lS9H5bd4yy6pos92JMz9UDfKgrETz0
tuTdvRmbB/G2ubRNkX6a9g59ZRKOdLyObY1FwES+7gblijCMajK2eq/7PrrDhVlTdwtUqGEXwRLb
OFpSQkE8/ALaSGxqaGogIfqqDDprBrhYjUV+5H7wCDaq83gffRLqbe/90SqZMf9sxrT8vp0wU+dm
E6l1G/NNXnse9JwxAiKSdkrCN8CPdhjmbLfrAprcIQvDvXsNyLR3Q0WkTEmD7GbTGqcrICQETMPQ
4Zjalv1Ys6brTA3X4r3A2qM73oBIme1dLKP7d3L6Di/I9HDDc7TlCx/7aSJ9bARg8Xe2EZHNgZbC
x7R42LQ1oMHum5QhQ7o5bef9OkoDJmUZG0PBUF5xcYk+T90Dcj4gJ2FPqGOFmFxXvuk1IzjhHVxq
yijEEdYXNrulowIK6cOm6HYXTEAB+OLe7TfVsiO8VcrIMTXkn+sdVDi/xKR86QRS8Uxn4b/uzcVx
syekHXZ6ZQI03QrUKlNebOZ1u1cMkG5MFQ4oJnOqNxOTSMX9q0tHy4or3YiF7lfzRNtt0SQLDZZp
Wa6NskeYYuI0xZ9gf3/WYfLUJuDNk9311WWwlV4rXpqJzBy3GmryANJHyunhvAPoSpy+QZ2raoos
wi2zb3Bn/dJ17/qtIePQpyfQVczA5a+KQC0Eyh1YGIYU6sPuqywLCBs0ksH6qi/lq//o4ymyseW5
Pvfu959y85vDTLXOn2GH3of1FHH07hMEQTHNR1GSRrzIjlO64vvGurOsg0X5cHZO+uHovESl6845
w2cs/B9d03Hrh+ABpO4ri5BpGEKSytuj1AAOuoO9b4MhYJcz6mFjX0BrIHkLbyZ1TLhplGu8x+Xp
9YbohsXfVzLAJ/KGTD3IGw2Y6nhBOi/bR51nJ4LZGHbYJmcxafQMiB1x/9Dxsj8uKKVepTNFFM7T
F3n590Dprinpgruht4FUXg3cvjxf4rozSuoINJ3qEFh5kOtWGyUDMIPuVMM4V2g5wCb8a/lKd5ei
C6mEcXoAUJUjTozFbUcv8wNm8SaiQz0FfuZ4B0QyaHJtYmvld2po+cSw11EI6pcECmZKAKa/gDdu
6VeHh9KB3cEKk+RdkuRNn708ux77c02eZZOBm1ZMzvik0NEZyBvXH2cxwkcgC78jnaJ9LTgGVMHL
63+ic2rmWwtvT+JO4T4IRj/3yh3RsexCGGs8Nf6zrk8H2s5LAjSb8gh60lDSE6ezlluMkgnJVABM
U1A2oDahB2eLI4iEB4rH6gsG+/1VTWMAPA8b8gE4KWCFh37ozipMzDIjXPGLt6wC+xEGCoqjPo16
9+sJkVHZVU4xdd1P0QCHXJNwlKCatNwjJGriWC39270B/cRQGseNY3F2E4C/5BaHglZxPI1SzFC6
llF7ENt++1hWT0BcbsdJyMv4fgOQJLxT5b8GZvUN4O+qyehpu+JBLRGv5XNKnk7hbwks86/U3W4Z
DU43yG9rrQYDxZlS7Jyx+t0OlhB0EAo1Qwu88vlpLQEJ1vWiMMSgonUr0fUOIm63X26ZV8FhO3wc
8RdPOmvEfWK8zb7BJN9vp95i4dvzQNJgUzDTLyHKpl/XKoTih0WngcYogxN0jQS+GqFVwx+9K9ai
HY4FIpiu14Z18HFBsbry0su3DbZGnws1z8CO75eDJOauLrTL/GDSP4iilbHrHTZ0ybRipqrYfUKC
F4igkBuLVsSZ5eG7+cniMneRYTfrqDwUwem9JH9JYbFdVZAPQ9+I+PpKUk5AnUfUNJQ0yXnMv2vi
c4tzTNeZ4lDMESoVLU/j+XQ3SLhdNSuz9y4K53S62mpU8SSMiEZnFFOPPa6sOojV7wdDzSJtWTbH
6TQVymSNNGol6Jo8bViS8fXTtOSPLRCB6J3V4EtW08ujGY/Nmc+1p14BX4H/rX4xTy5lr5tlip+h
alf63Lon8oXodP5Mx2YtmWaYUCvWxeyOi7H7ANlRrn3Nh39d/s3MAdcZRXVlXAqGtMxB/gecernJ
8lFkt3qtu0L3SWOSZhUFbAB9OW8rsPZaGK5ZxWf/GR//btgZfu36ng3J+tma/W1+lH1SlNV435Xq
cje3r3MJQTMI5hHN1heDqo6yHNRr/lJBUt7MkdkZ84TLPibzcfv/VqrNulCue7YLt6AvF0jZI55H
MrP75+x5Dpa7aQ8dcxmzNMC0YEY9u5oHlqKtGz/qsRvdFgfFaKNQgK0sfFJfQMa1mBfj2btSwEbW
0JewRUhtmK9GbhRu1StXI+bQXLSb6LTP9xStnbUwQ8Io2EzhF+PdyPhgtO75bq5A4A1PHGNEdg8z
uR0x1iWVrywmEIcfx63gmhMmix6WoFZETWmJ6IlgbZDfGduwUqOV392qc0efJSujznc+6ahqSvww
V4Nmo1UZWzo9qko+GShG5WbnBGCrA4iBwEp6nbjZznORuuJxyTDLbsEt99EGtP4rWH2WzsYZCqGh
dZxKHwl9SDcQGog0Q6YtJmQhuGGM7EtOfX0/R1qMUdZE9m0JoLVpjV5XA0jaMHMlSeuQPkKiiMx/
DVr+at+0arui/bN39DUwhjHV6leD/bWdWTnRWDfils9IsDoCkDumZTbQjkvwcd2R6ziBuEKfk1Tc
cmqZIYIboaHF+mOCt+lhWj8jP7Y97pEa26i2lt7/miLCE+2nf9RhNufY98Bb1vuDgIig/3LLrKnX
xM/zENki4ehh7CLO5e2ROHdYoW4RCHcABQ26d4t+wiMIgDo77WuZ3lggDUUvEMM8vX5l7xYtCqZo
cph8JSNej83b+YJvtFZRJBTVfoZZbvcSK2748HgQ3WVpKd1TZsndx2pV2wDuTIP8jLMqZA2tVas6
MZH+brR9XZbP6CNezvYvj1jbBodmZRmmS4NOxqrowzrMjxTV4GvUTTFpITTWbnbQqBTRVmgx9q5f
4XwVQd452SvdjDCt4z1PhvuUSMbwF+z57qmzXGCdB4CLhuIGVctW2R4Q0AAq7vOxOMA5Nek964d/
5cMbpKBWpXuVsE51OMOoHdYgmbO5NsVD2E7yEqM/6ajFmIeUrGt+ufOULsBIfAfPlR2InsIS71xQ
8vyFJ0ST0SsYDccrnid7nFe3EhT8eTkmpScDorf6I6cXgDgiG1WIbas4Sgcfrfem90cstDHGV983
YT4uQgUuF+SgHCqGf+62cgjgTr4vHcf+6wNTW5yOzumxyN3H9/w9QtL34FJxDIvKI9sKJk91xYpj
hSloCbhKV7znkQP17XXioABlO4NFwPrrs5QcKqdJPi81djLJEMX5Ed3292Q+nDu7Po8lOEojDunj
Y8ODzKYB45XsBsVGx2OuwFJ33rzdXnUnkj8wq/aoJl33dlmy7mYUPe7T8JO2TYvheLNlLwTHBaSL
iNwWMjd8AT5weBKInxG+8kexcWZeTENiWap3JFxTnG8NiRf6wNsx/HeyLlxy938fYRyzXkZTH0zG
3j60Zaa8ZOCGFrahM7UKiWEWgYVIA7H7u9rSM9zc9kWNv9haRZunI6T5f3j1ZbtY0KrA2qT1vNsX
J2R6j+LojMdQHmhKqresgjuRHsUYzUIXPTCj0hEX+NKSveXWDXcJjWvyw1TMBYIKbnryqivuqv3B
FpPT4uvkVEi9Mwv1ONxciE9euJcYgJLg4TlU6Sms4hjawRPrhqxKFPgxSF1HkIu8st0zPh2jcYr2
Q0h9cLdnp52X9U4tADnE2j3+aPatwVxJG/YhuvwsHIokNuEvxsGce3H9EarpvemnLqa6cHsJiGIH
CuWNbSot4tubGIO7Fzp1OAThtP3AyIvHL1BQ6/hVZzk6yOFz3qOqoeXw5XZek4y639RRvjZ/4qWd
I0sMh5vcqxtnU62PRFLh4iD/3GEA3cXG+w42mEIJwFU/0QFJXf/EI0oXxqeLN9NocoDAr3JDOZIL
2xRE/pH0hYUpEJUsHhpGjqwRBrwHtQo63kCO/ju0ZZDKn36NqjLNYGecSgz7MyV1ODoDHuz5n8Gn
3lcK+uZBaMx6NrxEogDVLj4eCVOUtwSiH2EQXXYEtS8U1du7exIWR8Ue+gNvJIYu/w8iJ+66eTj5
cy0ApzbVxl9CUzBZsS13VpAMeBJqJY7zDgtWK05pC/s4q1LODUeqL7LEhFwi1snBVJLh6nA/TqC2
Sm0QW32wZb0XkGOwHEqExwEKNdCB1mdO4xmePbjbGMyYllnpDot78ItyYzHIDWF9WZXuwnbNsk0M
qovRpWAuqbVURXzqtawROG3ptEiNQZu1AafazmSoJX85fbeYdNanr6ls7784USpokJijQy/wpT7J
BP8lTeL+Kcjjtc5wSAFcZjiG07dJWddqLLIUn433uEzGqxZmLlGtm7qOX+8nX1K8C786QC0wn2Lq
jL4Aps2wVP+FVNcrTBR9xxtaKowV74vZ4DX//aBc4Bh2N0twAwQ1hiVUItWRGRWH18IZJPyg2ICg
QJ9ZLMKA/lp+DLTA8Ed1BvUaBQowvwpn2qjxmT8vbMupQaYv5x3BE7rPkXb/6OinsfuubMSib3gH
65Sd2zxwn+9gNMZSSzs+VWYsyJusPmxYdZr6vYT8pJq4sUPGnboTGKmx+MEu+WtIGVFwD1zeeqel
HAdjMp6Iny1bz/25qRwTbqzfv1WnbRKgJoQZW3aW6dt4to+wVg5wLMZltXrz7IufQQR1hJdrst7K
57tluSRz+Sg/OUv0rmw9J7N9zHNXMQN2NYtvldM4wCp54RtVRbq6PY5N2LV4XlU4JHlM9Fg186Eq
y1oFdDVLE3mTfK3VBYUJVA5LYTeobSQ7EEGpqy2uuVb19HasO4O8US4thFRRNAm97ujoMtxziZpI
jJmYzp5v9OIkm0MRAKUGCDYcyJTVcLVG8eLJ439iAzrTgcMxm7O0Ct089rF45/zN74civpzdrYMM
Y7xcH6fU6LRcMjozWF5V+pFKraT4YOwtPLoORp3h9Y9YaaNbu/V+FLLU5HTi3/WS0egaa3kO8vD8
PJh0OKVVaGm9F2+vau9OXACYX/HnH77j/rbpzIlj83HUosSO7e4ESQWv3nZ+U982O9wYlIndoz5q
KJ6ixGaf7Z8bmVMwRh7d2ASYso9VTb3I+lg4jZv0FSLu1wgrZLqIxoUIMRTYdavjVm+6p3aJQyUR
YQSTcdNFWSXNgITVWg/DMkrbT35AlaVJ6M7uVIS2c+/29qnQFm+30NnuB/c/CT2/3ccrWKX8NQA7
7SHo76uMmQCyUY0282DQpd2E31CpTiiENNQB8u6XtT03OsmOUt7CFcBLkjJmu8floVU3z1NNx+o2
PC1Zr0Ya3GkyaC8Ue6lUKlg7UthmTZerQVRN2ENc7VCy/eeD+97mqxPZdoK9LvPw6ChglHS1M83h
b245ynmmWwgfsZz0wWv1Aeg5EXJfa2LHR78YcHrhnTRJ/8nx9NG28FAAHNRrWnq7keo2fyWGE9lz
DHIJHuRtGoJLTSjWigOEhTiaT95kZVkauyOunVnBcpe7d068GxkscyLGhWzCWY6WyW696eCSG+jt
odEacKRmSluEl8t2BhGhRn5tnLMapz7Us/4L+6grY/9Qx/jBO0AZa2+cYfjBaRjHqpkbiP0GbANz
wK4SywKtFHlX5VOzwfqA3iPVjq7YW225qjumkQ9IPZ0cxrQ7DPdiAZTDCXjLS1h+ZemqU1j9Woaw
XdpG+AJIv7Eb1o4oirRNQmZp9VPgIJnqRwRrDzFsGRxp7+6QkZGrJeC/Rbe3iWPYt8nkuz9s3y8C
Oj0+Zf1HXNVaEksZ2ro+y/T83EBnJJrv1le1G1gGy8v1zRHohURH8BbyVvW3fSI3CB60wtxdf/PC
Lle7LGVtgwk7YJAeXR992jK8loHCZXu9VdUkXpNlxfLx1uEG0mzEEQn1toFztXAMXPQ+a/MNKKTv
ITvfRu5wU7n25r6IGwMChzd58ZTaDiU3aOBvljw+0JnTon/iKBxgztxGcrQi9EhtBBLhU6dEACQE
kK71t+Ml8ZKRBcM0svyuBu1Ga/LEGnqxSDQb5c398S5aFb7sOrIsqj9zpO1eSTkdhSrBh0jRXwpK
7FA8ycD0EKQBOcgJ79WIbmitI6USSq738IDaViuSbq08izaYSkO9cUXFXFIn5kOcNH7MnAlJLmL3
Pl1WCLzYiFSd5kv1TZHWDWGNg75hJI3kTP523U8eLeDFtgwYFNra2C/6VKF/9dO1CW21wOPcgmFj
OqB1wp9B0AyDIxHDUPqYGkLYkm6w83pBYjH8IxynibTXLCjAD/MZ/9dq3SWwjNvrB7IGLIJXyb9q
lnMjTkg2x+RnrUJTaEsraPUkJVgdjb26MfhteNYNe3B0dNwXu1TMPo6r1yIZZ1MBZ09RgBoMbp27
BRkfvI49rrGMNkTrHzpSFAgqsmyM6kKxMsnCCIzsksTd70LgXby2WgJ3YG9i4TNJREsLKTeHC80u
O0wr8HlPQPTcLc+gB6n6uv93J9dSASvs959+aosZTzNnlFjEZyIA1myA6aN6M7spqg+eDu/YbmuM
AvfF4JzSGuZ4Fa7QEXxBJOCno7LfZl4K16y4L1ECTwDZZWXim7g3W3i8wI/T5G5lc2taCD4VA+ia
UO9MpTHoFsgPdb7ZArfj177c+X+zZJnCjgPu+hViWRDBrt9fazNStdMttIDcc9RRsh9gfnEjclGK
8cE5yzyhsnWCiQdo0Eq/RO3e6/LrLnyqYzzqs99Srq3GfM2X9xPk3VDsUpzZTpc174RqBFrFlqOZ
sw1bDVeXkkWDqmecZaqFpe/9NHh2/psRfffjRWti8BEBRSwPgj5zYkNzbr9Va0lXwaCyoMUcB9nt
7gAKmoHIH9d54b/fdFzT0UChWU7YB4YJOgmKrzDFTvtTOcPD/nMi3i56c3IWuEcOlCRX7pY0iFP5
UJbqOvl6huf0u8fLf0KJnrag2yBoJY60OkLR/ZC4yLyLy1GDqnqAgU/D8asdY/iOWvUM4fhc5twI
b69NsOkSbheChV1LYUp94y0tNzVq0T+ec9Jflx+TrxokfBIBI034TWeLfn0WKBEulps4jocWgfgn
LTgHV8Gp0chI+QMr+6BruQuIIZ90sWIRdheEYCvrP6gq1Bp1izSpeSjwckCn0QnHvcfFNSJ90z7N
A4SyUu4qoVlg8wVWWikMzFIVQA7LgGPxlZgB+mkP+EYplLN8x6HNXL48UOFdlmXMBArbVLltgpaZ
eTTZOdMcbFa4SC7v67XC2O4Rn60bK8n/I2XmuYzfhpPy9qwYnJnoHtU8XaYOFwUQR4cbjI8vXD3V
lvjhjaLBYQu4UYNvdwRErXuX0LxhF8tEnfTVGdjwHMmvpnXytjckKJaosDLv6GJISgKC4UFaFNVS
4Tyvo/a8fu+kOcRTNzJ/iz0ObfVeFeJkkik8CA0SP8AF+DknsXrSS/W8JysgUCx6/JvScrJnabE0
bCr46LY7dU8Rhgn/oVLlBAfWNn24JU+PLxCrmVjR6chJ/z3BXVsOwb0wQgUOv2MFzw1gPMJrJMWD
Z+/AaTIX/W10+1mTmlcPpOCCc/ctE1MxcOXlPG6gSTlP6X7qROug8JaLJkjULW2BSQDqvGmRU2wa
QlSLpldfbfUwr0JEq/es31mV/znB4f+zSUZnfsqzNoZbAJzR+cPd29URQN2pgU9CsuRywV42Khb1
i6su/qpDibFQbsH023+7WPMjkASo1CbFSht2x4R2isq7kJS8Na7XUkDtEKJYnWm7bz9TO8vo0OJV
pVRSu3jUpycJJUBU28mnB+ll7+0obvFkqhnNhNMrGTgmSSD2ZCLGsQKsoiqA1MH+xrL71U9wSPrV
gCtKNsU7QUGUBOWPJ0BcMcaR8CKpy/uSdSzt5Mj8cJpBg4rW+O/oci3s6YKwnJ6uaa9JzSQXNfL6
oKso+E73oazHwMasEhQ6iRwmegREu6QzWo98MN7IRoplq2OGu0kFjMyNviL/0JsfOD6Whtp4XbZo
TSVVnRPLY8t5Y5LmdPIyeeHZO4rkhkYjJ47hSn6+99N1sCnna0l8HNnvYGe2bIpS/MSxfxswpIa5
4eYMJRZDKBObD1VatrD7yMPDJvIOcLiO5pcdGaiumTJ4nTjEbJOsd+aPsvOOXRklSBxJcWdtWSLs
UaomB3Sda8Kw74rmzzD2jXSce6UL4W5yxIUKuJ3BREoRHEGlPohacKazzCWjzISubcHCnL/nMJdF
9I9cHgp8msT0Dao2SA1v+K3RK8HPfP17p4xDX+k9VbuCyUXa6SC9tLtpRbaXiopky1RspWb7Pp03
4i7ECX5HsbYgjc/JLNXVwiW1pGpsqYvNTtNdwyoUqH/na+vR0Nbhldd1pVJCfvSvOLJilmNVfTEf
YsEXgXM1b5oQFM10UIL3UJgjXg3upbFXImI73rz2iu0txmR1gxTffm8lpuq0PZ3QzbGqreNucpLD
KUKL43ah5HHwfjIVhW1zg7QlJeh9Dqj2Xf+a9Tu8ALFPWWdVJhrZ17Zo80alUndhTky+KEeXQ4uj
RXx8lS/RtTPGQx5XjHUPTGgaic1hJ0rcFZFUyPUCbWn065WYneUlEWNwfA9Vz+i2Y03444UHShvm
hEFF7q5mi5gYKm9oz/yQx1AoJfBN0snucU9tfLoypNoAu9TjVwJ8HSxsYK1z6NfsqgwEaLl9RDDG
ciAeWxamsx6oTIbviAztWnOU54AapXeyzyXaFqa8qunhWFeJfxzF1Od6N1Vwhd/LSMd1cWdj9KGd
2e3sS60S5HEkX3DO1wxrxGL8Bp2MpdmcqZx3cAWUuhPlm65ZyfHUVzAvpJq5qRZWE8Jz57BVtKD0
CgSGeq+4fcqRLHPSs1ylGuRjOAQ4QNPXvB6+gIoY0sDxYIwUpn6lzed1pbERT4L0u7n4utEQjuqi
saNF/HP+bb0vYwaUdKE4izpUq6ME4g4IwolFditR4zkeaoFF5GbYTGfYwt/mSCWNYxDKGAuwFDqc
UnrY9+qMPfmo37FtJK3f38cCVLJq6ayF/Y498btu1Uml1ifcEeZgLoxcHIMHj8aY7SCrEzSqQenI
zT9TkSZAG4uOEnuHC8xDyZmmU7HbczDbz0oHQlFZcYx+TCRSzyL4Bw2fFdJlXHSYXH4P4sjE9KYS
Vb6LSRQ6gVgAmW/m8whIkvnnAwbJJnxR+aFuJx7Oe9CUrj/GasOk7lEtP3CSOGcryY3T+uXhkv5n
AsJ5tL6kUy0GScHLbFoXiXNCpOcMkyymEtMM/IB2vRYDS9tunet7hZ9PCQ6uT3bM+vfd8MmuEVow
roRNx0QUI9TRzceaaz2EaBsLxnTIOuI8tt5AZNW3TujAmcE2Wlyx5nl8RvHQzS1LUsHXdztuQ+Hj
NrMacN+fCNAw1YhITQbNDSvY3o8qocOneO1/Zbz+J5T38QlAb7OHZub3zQibPpDrR67Lx5j7Hn2H
GlGu1gbVAnwo8WtiPNAg3LdQ9XdfRrzVu5B0IhOm07p/ewhjOE8RDaRYvXpqzO8d1kGGsrvzyiI6
nSJ/4UTQie196Txej1LsTRo3dBHPFhHJPfQ1hKI5sHHI03a5Cil801MJEqbmdq2L6wjaCMGdmVbC
RLLZuZVZygRVQDsqeoSs1jwXKiP2X4q6yg5iaNais+eDM3I04Gy3NYSKy1+y4DxpucuNXZdHSJFj
k0jjDe9vcwYkcs7nVeJ7oH/EW5PO1J9rlypKLGJTZrjy29+rLJB+88PO2rIfaRrsrJq/7kkGwfDt
vZR0rRFUCpUF1FTx1p/AvpptZVVTHD2c9aW0AoUQyympZ2hhEzpkghoPxqlMgRyl3XcShVg+Ag2d
RhMu7+isckLYwnILz02c2Y9iVbfCPSS3+DbOqSsq35CcV70Ex7oxEtYqTfyEns/bEnIezTJIKfPw
aYvp/kcdqA1EI3pymKVzD3UqygdgxkrlgEhU5RUwct/JGHz0RKx2FTiSxW3SL7gvKs25sgPo2rhp
V1v1gxhbI5Xb+MZ6Yyn2TswhB3sAzU3iRmZ2X8eiez4/rNMyA1+ki3lvt3JnQxx3Oswgh6+5IoMz
+v9l2k4mPy7ne2JqmbmPpxftI1VrbvHsdwsaAUzmJecPC+gm/2/2BNLP6ypWqJqsG2r419Z5gPpH
1Tjh4F3WBJ4R0R0kqTjMmQCjl26z19O/pIgUglRPGvY3lo1VjD9IQhECQKU8gUHiYEAY7Jp0nwsi
A8fa3HzUUckVgWwq3sw5XLayKSyh/jX0EIsfpbxAw/dCQYmtxsnrZez/0ySkHIgRYGetP8x6FOLL
IiiqUa7fX9qhQZZro4qrU2df2emlRGyNAmGr0VMDz7KU4fWilmIqopc4jznkJdGa4aLk/EDre9Im
UJSaZAFX5COCo2IaOD/TpaMzpBxyXfj05OkDwi0rL7mb7mqdqMKDvARomaKBBIOLxk4Sb3ZvUEWM
gf7tAK2G8pEE1785L6aWLtDIfzQdl34VifiFYCh+PevmF5q9mdm2EkEV97gpxAv8k5jm9QeYS+DE
lFXjy4kywpQYNDG2rYVhyKBdIbqofT7ydQ7HpENClDgGruCIDLYf/AZAvlllRTArejj/RbG6wE9Z
4k98lEBnOoQJcJTx5acpNQaQ5HkU6OFILFQaRIdU9Ly3G840gVlUOk3EZrXWeB+KYw+zp/+TfXl9
LvAmv/kYUl+Gh5DvBeC9DmxejoOzOBF8tZv9peSqt0DpXEp6olatsQLxTUBjqL8TNbQAsfGgAfXK
5ufm804mH0ByChWmQvlZCQKWYzm5OyLIq49t7eV+7jxGHAEi9NHTPl7wFBigTHSz78b3LuYSFkpZ
CRjlrA3IDCUSS6N+EG6bTf7OXDBiyjkh3f5F/DoX3QVWM1XP0vOONyGCRkCgwLFOsEe3aWP+eBJF
eZPTzdMzK/sB+RwH2dvQolBcdj/h3DRbOAWD59xoo+n+xa/0+4dLEImbVgkkF9zPfy5urjOyJQuD
f0tWo91YHTiwGBYb8kb2RCr1jH6eqyF1ma/ZQfKEHaNHT+A7gUsF7EMSoD7aEINTEojrqe0JGXM5
yJbIDWwfY+wE9eb6KzqZCLyU3Wm4DTk2Os0E3MYhCU1G9cwVJSq0hIZyTjRLEvnVzeqmDWibfGHs
AGgs9vMSjb6tTb/UziSrHtSPNpe9cv8xb/eLV/Df8jykOH0PQexArjfMaVxoAUk+ga47+DUGxY6L
t8UVH+m50wE9F5pDVKh2jwbTKE4pIRojNv/3R0Oy/Ccyj+0XU/U/zdWIDyz4QOwzuHlK/JjmO4Ul
E+g5de3dYzUWkoKQlZkNe5cu4s43kwNyed5m/Z4BipRewr7lLZszBY/xdE6aMgUza1zgILMzePa2
GODSDxxt5ONOWODv/M7c69ViNIiO2wLbrsxYpGfBN4rBnjChJYJq5/vc6ql63qXTTdz9rQmWnMoM
Y1vNB10xMQlFCrlm4k2nN6rVDpCTkvheNjM1Ygrrs93i/TsHGtGI/fj0GZkgNifwsJSfcwydpMC4
+9wKhZ+onXpTTYNg9HCHX0sboNGKXDT7dBoKjFK5QTeRdv9N7q/8c8CgJPnMDntiXyLn6xZVK3zi
MT6+Mvg/Q8FRh4cBfZlPn3kx7oILZmWlJNd7QQFvCDU20Y07/qX+68w+bExv61yMSyHlq9+BYLaY
AZwuihZ/YSwkLU4fJpqK8uxR9wLVOMqtT66LAtSQi4MkDFjGfSOTEf2LGz/D4hDNxT4DZWSXteoo
WNkcU47bFXW/1LtLqGnE4pFjGqHxF9Xw1BkzrodvfPMOL/J5uxAJV1P1r2NdByjlYxyQ0P7vyhF+
+a+tkFWsa6wdO1fk/oIMEqf6PxGnrbgRrx2s8Q5DhOi5DgIuMGZFGdHUEjD7mpfQIopIaWCDlI/g
cHU+5nkOZ4ramtbHeG2qB5qCXSel4c51pMOsXSk3sZdhJJ+mdMnE9EkBaV7XYuKrlv2FWzqtcnjO
gXHQRQFw9M+MqDcqP40QtqmNWxTRzriDpO8JBsCJQXTKSMegQ70IoPN3MfSvWL8dU5A5LSLaNNd+
bUkMRuIVBhNVuu0GvEvU7Hl6OmLOgxMI9ZXy+4npBNUXsM8ogzb4zHfbeWU1On6OjfEWQD5izjBa
Rw2vuOJzvSh+D3G8TGGla/BI3k1eD2UhmwmJRc79sEgVVBKhakiaAMWeap3fPO3aEyvqw8hm83ha
c418MCdfEP1AMFBxxmQDbFJJdtrkaa5s0pcWopBmSHj2OfsgSwcz4oAJ7KikhoiNJyC7q7fex0B3
r4GU6YH/BMEVzKZOvkSE5X9O9AnlC/10uQwAX7HGRbIn3e63t6+y4KNWt71VS+uYU4wcveFRFutg
fQ4/t2Z018cb8eZC+xaHtsMQwGjAgcUXMys+eOPw7cEiB4wEhsFmkjhFnSkDV+jXBoQuw+agrc+e
XZwp7fPVIYpyz9LpNnoCZtnf8HMM6UKOF+cfSMjNLXLZMQHwHt/ThS7W7ZJazMbSqOGcTa4y+a7l
R9j1gJA67f0oSDxyZ1YxKcTX5Yp0Cf+LytqfTY09GCMwkeNG9VM3kHISukuHa2H1wvszrxNA1IJA
snCyjTZWKXgZMtT0xhhc2ojST/9BLD91EcQE3ULeg3Mot7ZNYvHRhGRJ9xXj1gyYycsir1V442E/
E53I1EoYxt/ndcHgebO45ysGBJdoCbmCL3x4ktbl1Uiiy0ZIC680EWsiLJ2zu9w4GWv7eZCMK2MQ
O15bSXw1V9sCfBDRtTLdN6cvtQv+VYKOd24Ibvm9OuAwzSgCkD6u/L6KxhS0DMmC7o+WvvSRDo0H
NaxBWUyTQBPr+sTuSDjMrM9apSXAbwKSdBJHn47yYmRrWEP4HISn62MKS6UtRQ+LiWxAu0gQUDFz
uTeAs9h/YnBCnO8sql8kgR2AMCQ4HBSfzW2oJGn3appxGleB5soUWwmTOhOE1arzcngt2OL3nItX
KIi8sdstxrfuHNBySN92jtj1TDfhnfZXl1ay2qCymuSVoH40ENIyFgWHillW7Y02MF5SkTo8mZtS
aGUmQd73Fp7biJQxZYn3t5LR2dhShfKyRDyJ6inCC0BQYplLr0SHENIEx2124+/QlXhVE4VdMNvL
MKhwehq2u3EsMjm9LEmamRrL+AMjH8C2D5N1JFiz6Sj3E8R/+aVY6alhmyJ9cfsosAefaZ9xCDyR
xHJ/wULmizlioJex2No1DELl2hHPEbqogTKT3bQ9Vdhmq0dPQ9AG7lLupc8EO5a3QGNkkv/Rw27I
jRarM4TF20Mk/AB/Qn2n+PYo2kMp7MKNpw6ObNShjHFJxyy2wx/dLAx7imI+KX46tr8cCkjT5UgW
5yopb1lIhMbDon1vcjjLd6jsRSH9zCNpQgmON/pNFUOrS+dyN7EOG+BSH+wMlL0UYRLaRPVQw/hp
aM7aYJ4M+peSG07PeqnxFR7sjZ8pgsIy9UFo1vhuCCcPs8biVRXcQYM+3UoQMGa2Sc9P/lh36h6U
jD1NxAliKHOL2LOmXRF+38koPIU/M3YBTFMFzUpDeCXmPt0t6PHioUCsA4lG4awTmv1dRGAEMxNb
D3YmHDGINnfstZOC+x4Z2vdnRjDMWw+CvZbjUS9u/ILfm5k/CRxi1fGorMBviohE7S4rNQyAZIpl
AvEwpe3iRtA6gz+88PHvN6mM0dZozE5myoX72Q5CcM87tYzPwFO7/Gvw72MPuAFIcdsTrhXIB4e3
y5tZTDHL4y8T7AqHUcHtC9DK1TjHhl3xSJCX5fpS4SpdoPKVHb5aNrlU52r199WAlVpdbp0ocK5O
Z+U+m1weQuIci2krj20YyvxID6CDbbyx7V0xshdXuClq6lAHMdlArPuDBaJpHMPauJp3AsJXHm7K
iW3o7+p2/e5LW7uI1SfZPQwMRTt1B1IUYFVv6lJBsd1pN+8t7C96xHmclnTSO1rg20SA5+ltMyyD
o+j19lkUiOoBXrfMcKWmNDsFmpy4vrHYaIsCCalVSCOv0BI+0X68Cf7oOh+h35bJxrrTVFaAKgvg
qxUg9wAxtcMfipYrFQ3EMp8pXLlXlSekdNfhyRw4hQjMWc28dJcngPqwplu7F0u400xSumR6hj+H
lwhvvg9s57Q/UA+KgQMPlUslbPNdaQhtOaHFRXOVmZvG2F9DrArEmVsbOhkSW3Xq0qYxlpUVBzkc
x/YrJB3hBUjnMLp7fmeKKjNbhUDa4oFIjRXzOhAj6IoVSTV2gb9vbv1KSX6+raJwlqfPirlLm0m2
qlEfujNZgib9hV9ReqhyD15V+cyyVncM+AZbLPVDr1YKp+PHnD3FP/zCtPYNAh2tST7EFQ68TOny
OI7dNyCFPpx4hb0KRuWpOl39UXt3j0Oiuf5bjZJIQ3bgy1oAK9Un3oCmxKRQVDoKQQ14U41ivO0F
FMIYnpnun+f87yHj02kiJivbKNzo1w3kUMZpdlml0qrQOkN6etOP2yMkiGnGoGmaupRXu/gjbGt4
l5ThVy+srsZnhN/Eaq90cR+VloYbEiaz+nOwB5vmL/yRjaKIcBh4CUseyve4nEYaTCYjEBAVzlj5
pOOHVHVpuOY8L2/tSoVOuPw6oJLPXdSiLaIqC7c+Kaio/XpxYZKFdIn3jiUZmdpyZdBN3mC5fqF7
HGAdlghbgOgSh4PIXoil9gTPEs5uEcvwT3kzf0FvdIezdvseY6h/BbHEW2WfjuffCld6mavwwiu+
4EAXzscSx+//f0kKyD4glm9WmBQBMDfpHA+crzCxkruBR0YcSsOoeJ4BQ+55nFeWkyNSVc3hw9JF
BVj+L4ereDRpM/RiOgurXLTNd5nveCPY/I2ZV7WR9GYiQnC4k1sMVSELl2nzylyCywFz+W1RFb16
JTD9505CVxwAI8tEDrqKdBBEwVdeJGiT6fbJoLnKrCsQHU6jtybMDHoG+I/JRI8GOWVZYiiqK7CU
zDAIq8jpnFrei74XgRcYyaW8mxGzz/9qNc3p5bFTqzLYLulhn6jr2r2u28XsXrF24lpkZdHdcitE
niSes/k8p9FoEiH5cTyQJQLyJTweemlanU3JVIvQFZW0ANu7vlvzAMwyi+FKImgHQnoPhsyvdD4j
Vm4+kklKSp6mS0WoGmYhhWk4cNaB+OygNurpEndOM19iChoobhuzyXhfeDfRGJ41L+GNJkfY1haG
55rLC+Uqddhmjl61C6E4K2hmU+fnrOiL3kXus7wUxghhAQWC31tt909MdvWWT8LT+zClYFU0ZzBF
x29czuSQHLymVxF8ljl6cWiZvye+KKdYUpr+AIbho/VelgGqcsw+GkL3YaGb/tjl1vPJ4MS7W0BA
FfIFNrm1XwPBvevBQ1wD4wEVJwtjflSZjkT2+MqLzmrOu8syZwx0Do+4/igbDwPyrKO8gpMzJNGV
SUFecnr480YRX2qy8wm9Z3BAoEsaDFC2LJFyHezKSyuXizhZKBa7B2AS+7kRc2dkJ6krCAnme6Zq
ibfcZVMZok4m9q/gmhjPzcSLXcynj1dDCEM6AAvicVIjcnH8IR/k45EK4B1jKCpYHabimVcL88IT
+BbbJkPeCGnFebC//LoclvZ2NG3lsRk8BM10XQdrkZ1yVFOEjen9kS1IeCdfIGbI+9Tp2hTRrT6F
ET/tWEHshG8vPTN/xSOGt07gvQb8l/R0KdUlRL1YJuhWwdnrj1RobUYNF4tQ+OCcYUYTbO3+nEeO
leoMUy/YAhLmyDIy2j4CgOgthSsjdruiNB6ni+9/RINzLOY+oboZCVWeIt2JW5mx2vLAS+jeFfsZ
JzWQAP26OVHvvc48tAjmOpKdMzm4PjL3axO3n79e8vH1pMd1UGvqax4t39WF2DYjwGuBNhbp5zzc
WYEn7bVjEizpMBimELyyPZrrjDA/uQj0fY/hrMKlbuUwKJgUSddDyA7w87XF1wJa6tQafcYDSuok
4PTMid4y2rfOUrpIUku1FonOd9e4xoxZfN0Hz4/eAEaQCgsghzJnqzKAM2zXCCDM0N1dpbpTGtFx
QLNIyqBjkOmechUqjm3XeJvj1mz9Pj3MjINc711P3Eo/EBjXDEJxvPeoohBskeESml3RhvDHUK0F
frQrPatgr1+39+WNkPL4vYMQKf6hvnPQZ+AsksoBeSG8h0BS6LSGlY3UVzOMjVCaysZa/dmblRgM
A7n5pkFQkOR66H+sLikz797ExLTWa7U5JW9syVwkIkUrk9j4k/jI0Kz9QziKfdTy15rqVNr6GTjS
icjcPD/rRdD+p3Y/T7EBI0kzzcIPUznZnCFkcJ4fxrs2IeJ+8Bjz7h89VkNi+y/z8a2Lh3uCwkTS
6iP9CbnMAHFT+khcrw+b48QFWaUq5tUehw7juCzrtr7bWAI97nDI+jcE2fX7wFllQTeQGg58YBcU
BgZwwgP4U1ti+M6aVGfoKlhnHRrSfAjS9odwvtsZ1yHppgbPd/Q/XaERc/aRJ5O6yx8vvP8VP6Yc
Iha34fppHVT97hMd29q2ZrfnN3oomHkp8wcYMpJM4Ifo5y9eMePilx1X71ctJrp9ngmJF8PleGY7
bc14y0mVbJBnXZr4eeXqIhNvUrWig7fIhyNu/Xn7CN0t9UtE8iCvHNYIiIJBmKf6HChqpSd/fnzz
HGzVuUnzR6TEgZG1haOsrAKc/gr8E9+lXtiQOzMDgdwIrRF8799uzRzAobSCZvNegudIe6AWhX0L
/6mEO48Jg8ImtVQ7/btvef+NpLQ9I2KkZO6fnaBV3oXjjqsQnA5cfAn/Tgtabdx+CSDJTVVPMgKb
b8ZNDqHRTodsDmPymHeNONw42sKISliHlzu3Z/01Ly35O8O7Lz/gOyYzK45z/CC7KUuKGRTxs3o9
FLs2X8ttwh69wmdj+BFaYcTltRzyGTwenZVCgLQP0tlfeMREKW5oM8+e302FJeDuoOQtkDfpod1L
GFogtEAdHnMMjnkN0A5lpO9vEpCpnKt6OtJ/FuIj9Eo74dQBxoDuJBO7/uC860M9Ct0ZS8x9OQxM
8bEHDY5hk20+7vwF//uKr3WceUb54/zZ6yEI971A6rpD7l3BteeazzVW2RWpvdf7LoyzuOu4WT+7
fkAZgT10HKiVP3la4CIeauT6fsGhSVydEWf7K3N45rmD0U9uKcbtc3S/V6KILDEdALmsmBssVffs
oi2w5OebGR0eHlyCT+kvdMzoEQLruWACyGbHUvC9S+A0WcRnWDdyUYxvuKJgxBF9VJYXXDj33cag
mM/tZ8VtaRJFn1AsU2mHoMau2lj/xAHaLbXf/ghqM0CuH0sNCETJplz9EOH1iA3KxcAWEuNb/JcL
sJe2uIfNgPW61kl1kLLte2BJVOsfj/cZDgqpozxfFamv1RLayd/C7ptMEAe8N18qWC6l9DxaIdcM
CHhsTKYkRWr2+NCV4xbdfbw1v+3Hzvxf2KDITrZTsIw8ADwBOk1R2vSfh6/E2qhHHQpSrR8HoNn0
q1JDVtRytIKmbfbv1R8hB62033fOMxDfiZuoRrRgG705q7FgMAUKNplzj6cM3khEgHqsVvH0tq5j
WUNzNHDYY2G9Z4bkDixDn+RMuQmP6CFRNokvUJfbqrFZrNw1WMzQQDIZzNcxynrJiHoG5Tg8jDNf
bme7GMizz+xlY5LzC+LjCNJ31HA/lvHr27FK370eWU+QzrEUGJeFpebwvAVD91zxc5vYKEwgbMPt
1kaCZmayaDcndHtKH9es1NKUeNcjP/Yi3dqmgunMkBMLT3+IBHSrj5tm3IhLX0x+gggIcvnc6e7p
XTx6uiFW7BZ4imaAWiYE+OoiHDy37PAMdg6Kd7MkW1VZuQD1c6wKjd/bwGK6g5rFg4mJv70lwdrd
C8syBrIiQuszWqER7Cht3dPpIA+f82emH8ZroOJKeLlTISJiM+GkpkcqDt4TDowEkFlrIKYHAEwV
t14RQ09yBbCgRw1lsXW5PTbg0Ew/oTAnyBTLApS10yMAJSqQYz1m8SycUto/y7L7/iLdkfLvfGqx
FzWZYUoOnMlaewt6OsV+mtvLAVLYfYx3C0Pzhh02CNdKfqgyww4AP5n6mAR/+h5UgQN0QKQsz2bl
srcxq69H9kUVsOnlsCLQxZZAV0mCb/NJaKHSm8MLVZgnqFAlhgaZMNFf82WNpm/6VSeDJwK92MdA
4DfcpCQSWvZ67OIoSc29Ddc5Ci+7MuCRhvXgmYTHIBgfiglFtwITDvpeI2b9g6hOrDcze+CBrKiz
RTSOacZR9WSbQnzMCGdUmApv5xrnEJz0bfKud2JLwGMYvOZm0fCPxm36/iOHiBc9WhS50qvv5c8U
F9pqZ19aYugy5vrE6zleJ0rt8w/vpDpuZr16jE4XzpiXm2tbgsfyZBKBgo7aYFPwFfISu4aRHozY
SFIX5nHm8NHS2f6hWZcEVeecowbSt/0IJSQ1tLY42bczDdxHX8C7bXMDSFjzSCdhY9g9XqFJzxPu
F4Zw8QMp3+pHO/VsEot4ionT93viw0oke9zabpnoEvopK5hilxz92QtD7od7zD7kHWH152434Qy3
Pl7KUyZKXMrzr9oMBqpxxrLZUb3Di4PbdpsqTEzqFwmaWSCLGgZbt86UpDeHq7a7NkT4CujJxg3U
sRnjqGfJBcL9SB82qiC4mfaslzjDIZpQhCxHnpmzolOmcLAGIu5JZn2W9eS8soKffRt8K0in7Cb5
VqcB37pGVuXMivtxoddLenU6JRifpKYCAgxc+YktGpARvUNZ4PC1iR+OCvoMfZSkam4KK/hkP1v2
QsMuDPX7UcGl/3txUh/hexv0Jnx4RVZPcKoRcPLl2dMBcT9p/JUifxEJVejQUuirKS8Pyx7eNDhu
ERj1LoCioS9WNWhhEiZE3+XP2iPCuU+KsKrROKMMVAIzcHuzM1USJTf25N55WmfDGxcUl1Wx0fpf
aojQkokd5/VNAMSIpVE3TNvp0Snpnr/WWmJ/xGkbQDCorMyeswAB1X01Jn46rdePUL0UTVEbQgeh
2HcBbeYjWpg4J3p+FJBw7HJ/6JZDeJR/eelPNvQp6DGAyki0DamE5m2dwcTQshvgLfg3Q2Q+EguQ
5M3ZWF4xu4s+vRoPXI7Tpu7Su1Daxh3FXSISVSJEGtf8Hj8haqDJ409KGB16QYUJr4bY1vJ8cEUj
Rsj0FPdBmn4mkc3SPnsH8Gfb+AIEhbNrQDX9reV/WigWYAEg/x8AnvBVrv3VBQu+ZRGWXg8JkWQJ
0wxaqoUZ+im/DU/uW7hB9KSYhHNZrZq2hwwc1yWbdEKl4r0LzXZ6xeFJ/T5MYiSTCpy80ocCZ9ip
RAYyGoKiFVFK4TNxdaXJgx7RJXC00aEWfLFTTPGQDeMix5P2vMZX8XVSHUmKnlUo/AGuMVexuMXx
QJwCe3eKC93ksH41EK/Skc6GV1o6hsEjFzyYytAQ75DeGeQ7qnNY4fjCxH7abrMM3mjJGHUQwX/g
F8proZ5UnL48MlOUx2f2cTcPl2gvEdNCVv9od1jtIVoXFCCEUV/gYIMEUNqrhUe01M6c2o2oLRTy
YXG+SoEkhJ63sCN2dVZ4sPZep1FCqWA2ASdKrXml7wFef5pbno7GfoqzCCqL6ek1gsOXDRWLkBrC
w4CW/Udubnp2ug4r1tuwVyaRpC/Z3WTNFYNCI/SbU1kMZl5Zzd7UEAhxcOniebfpcM0LX4Ec5lAC
E4UsaxtkV9JChkveQYNPiWophoV7VBLsmC7Qkc64cW0s8kuVwWUeOa26HaAYnRT8ktf6JHV8L78N
vCOHlPBSVPNtY9a1i1hb/oBDyA51+kolsnXhqlSBOfW8B5eLn1gZVoJgMENQERbWw1pyZc3HwA0c
eq1L4CP0OKUJctYMX3MZ0zep4Z3lqeJqOLwWXNE8X/a9KuTHCKAW4Kl7QBQs4VxuFNew9hPWyapX
k/qofttFGBkqFP2yzpUP0TQh0TEVvAHx8QBTBE4RVs+GX+T2gWrSkKXvkz/K+HZUd02ePr9LsrgQ
2Ehvl0IaZc/3g+WgplUXBMEiu0VYHf/PvAxx5k/X5b3idekbiW6mfK1hFG0N0IWNaGx+Vc+oSNe8
N8IyLPm7cYdlcGxArLiP4lOXsJVmQPN3xMrg5DMprQE6BLY/RfGuAD8SDE42lU7Qg+eWGdmvFndi
VXut2PHQdxRpFPnEyzN9w4I3l6GZklvfGbXyZgbRDDIvzP7/xKmyANXYOgPRKNyC9TkcGI+cLmvS
1fGzJHdElRpnjEcjGx/yUOCxiTFmdsxVwm12DtmauVwi+ULpXwN7LdLVOfSCzxDE37nJUZButOnP
Ns7YF7UwNXboOFknxNy9jMDyrm6pjsmUNxvD6LuvvSYVmEvw9g/jBkFBXNBkVLqBBjewQKg/NED9
FG8JQtYBgu/F3naMcsYkmydtj9nz+Rt2lHs8WfXXKYEObpdat9F8qnt0jEUCIrdQYoi/l4d8Xefa
ySO9QdQhNh6midiUu0TNVE9slvNI4N8w5R4hmanO+W+0SWuXGcdsVOhmAIj6i/2NTnasMYjpB/pA
5y6UzJJhWRyU3Vdaev1NyNC/fBh71RTpDRP5jQj6OeaodbtyUB1YfM6i+RU1BnfBIsvSpqRSgsbb
TKGm0lwaANdzxoXj2qgz5qy++wcqlV1PTtzdDT8x/9qWm3N/76lsIu+GQAUTgu5y2rAhdnmaptoA
zACxhkDkehJm+RlxvvxH2YQrP44aL57ex3ANE4mXWkDTOKjkhNOzk3vryZVTzsuA3JUmIbYaoxh6
gMlensdt1dW1G4CHsEfWG5kIsHlEULq6zZYb/Gok9vq8upCpW3HoNyIINVVJlVMw4wsjaA4iLirH
PR6GgvzpctT+Vnmv2e4ljsqnz7hUKAgtY0gmFrZ4UvsDYk2hrdDI+uBSJpTzRK/QXPBe1xwv3LJI
/kFGhl8J70kRrB8RtTetxen9lGtrDu6u7BVxOoYpfsku7/vb7hWBvt4OrMJHZPHWmqnv9sez3Jtq
sjddQVv11tgMzOZ1hKam2W7gdTcMVkfvG/3f1b+fSdStqnmc5LltBN5Bb5pYOUgFaRvWxhJJnWXa
LwaLgv4ewwJwD22n9O9ScGYmRsEg00WepjXgMymZXnjU5ItIVzkIb7m0zix/5M0C/os6NfsSDP9a
oPVCK2TQig1MCSxcEhyzp3FmvJfGgA117PRisO2ruj9IMhZGv1HYgLrLVHVSsZ/MxQOwbdgXutN6
cpQ/EI40mjAci43iCt/LGn2aLqCNxUjdnf3s7uDnSVNZ60AwLy/ngL7n3ikAZLY3QIne7ooryk+5
JpewSFT+y/U1y641dklD8UD8Vt8SCAJvg8B1qrVukVp7O4FHCBuVsJnKXOGkWiOrDsdpkI+/0FZe
WQMJVhqdjYhrjeAA+NuYj2muUcujWF3gbUsKYVqhLz+x4dVm0sYXECBygA9LRV4i4Q9zsx6DIN/j
B2mwbSSfHP2crqh/O+izbCt0CKeAIyOrkea0nROPiwHPPVs/Zb/OahoLCdV0EQ95CM8NmSbLJZFs
cHTUFJp5O6lygIBjHL3tB4tGwm1+h63DG7IqoWKuwrIGuUCe0HIlQNVR0mX7Q4qWpN1wTJIGpCwF
W7QU6m+w6qcNmYzSZy9tlBDpinMIFh60VAUb0lI1ScqOJo+WBC6Gx7WW4nT+nwfBXGsRmav4hGBf
frZKIbubbCByXB/Rvwj3MgLNlzNsqbpeQpDpItfOjjDqYN0V0ptVO3tL6QDcxbiucKr7h3VUrt71
jpGbSl+6nJEtYxP/CufYVc4AUhIL1TFqvnl0SSKu2/jnnJqtSsKdQts3rHJjyzR3sn1HBu1suO6c
9/f2FDaqQKqJqQj1q3DWCkEAjhPKCPyMTAJcaPU1ZQXoMC9WXU0syHr0Q8nlibrXY/WGF+lhzkNX
aPi982AYcP11MNZq9lL+pAb+W9mjHx17UZlvrM+GcLP03kp1nlEHIqkB/HBLkZMp8T8oKWcwoquV
ZSoBFl1+GwAif9SLEiK31AGPuQhEUl6B+J1hWwrtTp46wVX0LVXvi6wdgNWhB00KnjHu9/mRrzoN
QB+dmI9Ca6ncvoOfgkT8V3vvF8cmHd52+FSUh0/vmzbaQfK2QluCRXRm+FkWI8wFCniawRrEJSp+
l2wcuCXhD4LVHCUkkvnquTu2ZK0cNDgQiLkmipepmO1+9ia+KJMK7h8Clkg2BDv7eZW998q7Fw6h
Jg/z9RwmRb/79iPvDtz6iwhfAOR1ULa14lX+n1wyvEBxJBWS22Q6oV10ztP3Z4zhPZtWkppozQVJ
DiEfAEk1wfSh4hUctRu5YVAh13GTB8rIMdD8FJ3VN9vIxaXraQef9fcbfdL/RHR7Pc8+ko7AFCCq
qOe5K6HGXsz4PYQt4gwWLTWM/j+7GEJJWkO5l18v9RDJs0BKI0UnJleWCUEa5jp5ZRPoc0WHasxc
ROM6J753su52DRLdzgMwSL6v63BMi8VCdcrmVJlB9EBSiqmsQgKAfEUi18iJAhbglR4C5MF4d4Gp
JvxU+KDEp73svOu9+wCYEqubOjgFf4t+xKfxB0n/7EbVPjfqnk2QO+Meltqc4p9ecrWCTSlOEQF8
iSXMYiYmZ2X4MxWEhSKi5lUiFZQ8hx/gkEgX1QIUvM8W4b4WrNHi11GA6u+tawxJ4bMDFZTWKGu3
BC1VRl8DI/10jovHf7FIQ0tTT7b+AVP40CaYxpFE/CPAvGnA8wX07jyUkhrQIZEHt47zk+zFnjiP
NQs2Em93bLX0b47kEJRuteaS/h7bMcaQX7wxG/oeWV1WliOZv4c8qTLcIhBApttEoAyFqMN4yXba
6FsX7+9/b9eDClEFnIcPxQOmZLJLj00opDESb7cj8MBypLC1T1Fn4aTnmj43Rhzq04ieGYDcMIsK
mRwXoXxPnibcYWzzAj/C11U26Iavi2pb3OWt6JjZmLCG01Xsfo2qJjmfUxSFBG1jzzceSmrcltwv
uGvewMwNl89UxJYHB3OnqLfY95vx9sV+mvAIOuFNVPZmvg+SCX5y3NZmggFT4c/3+csfBjhSOO99
8Db9Jo5/18M4RGDuLVqZo/Ff+JMPdgBsh3ppc5t8RkYqIdaA7f+YJbjku0wA8TdEoLdEiWmKO5pW
fL7IT3f1MMrtcRIaWW2F/m48J4Lsbe7xFfkqMU2zUWF+1vxeCi7STfuLUO06gZju2iRJcCdZwuud
oA5gqo+pHRq9dYWijjZAgUoJXWgJYtdsFWmNLap5gKYdv+581Of9h5ecs+pkQw5rwGnYX3FyHxp1
KTY7R/ykrlMa35mptA8HXQ7qij+XHbkEktPJyGDf34HDDkWoSVI81ezPeAORWgcRZZe5Qqj79aZx
fAhdmt7QxJjExiiUJ1be8IuicPimrGok4P69ZXBlU6tiHIKUHEE4ymCYirpsd0NtgRK/3kMR8zkA
9ACO04n2G0OEeADiupWzLH3ZDKTYZbPJ2JhIdOKnRBBkmHmhRiT5NPkwpk5GgKmxJLVvmRrH5/N5
bKE93rhBWf1hH5w8+KZhLISu6De2r+Akx8mCslqiJVGmDV43+U1FMCg6NVn4Fa1Ir1HVri7xE7si
+FnvlTyfjcTXISnwuGaPMhqK6RF+KniSuh3sZmpuZMqabOSyoH534kKVhPveVUxzC7dRYfHaSpi6
iRX2RUi9IqB3omngLUZyZvnOwmeX7m0LsqlhgGBNwM/Snhtrz3J0Ac8aSCUM4lh3UsaqxtMqAmrg
XcSwzb8JctcvjHGamQ78X0VZuSTDTUYc4ObdY0bk7kbXTo/tKXhJXeo9xnWLQybdTYfs04JPi1A4
dZN9y2Rxg5U280+WMldLiNEk9o1X5QS0nbZvZ0nmvRhpItt+QrzrNNmFdxJxaGcsBqIA9nLA8OTW
2kSgeNMVaTgsOq+o8s1L9l53GxtOiLJ5/8tDC3JdNDg7TCf8bnBJ2H4UdA7bQkx7Z03d94WYs0DV
uikW2KeeOdhKiN5wjFP603V8KQD2x1NCz/MuvydJYOqjadpJDTuwvhqHtO6pJlkxHDbD1Wgtwp2t
CuazUR6PY3L5FEwHLnqHvRZZ2sHp/tmFbTycFZFtwn2k+uh/qdJW7HeGZ+W7YbA0LD7iodaVvav7
Z8v6L8mbhxSlgcQCj+e7bhKDBVNJdnuK/s4kS1UZU7YJwFms2dVeXvugHvSr6QOmVVXfxCBgBbEQ
Bz4TDZVl2evr5dn7Ti0EPT0ta26eIXZ4O14GLEGWRu/dAUF4owvUKGaBElgfNaqOknfGByC1XK1Z
+hvAF8jJg7Ls4y2C73Sf2OXhHVpeT7jnPFJnkmrFJ8FMVY7qhCsTbfBrapDtQf+pOEZikED8f7Xm
RyQFJlLBToqm5iFv4WKQRzgkJNBUWsS0duhmt2MroY4fDi8EDtv84AjV6Dd97M4+yYYYRkJYgLjh
5/HlCqzcJuePCdOOreJIYiBUDwYVejX+wB2uzma0CSFy059zgcCIAGT6L5GwfgrGMwq3okWogF4a
91E9x8K7dCBa/hQiBB9pCMeYKVAf1r7qz6d4yxmztg3L7cM7ex875fhi2Yt/TA3Nbw4HjnuHHrNd
q7l464pd/zwfDrOo7xqMdpHhQlwcfSxax88w713yKtHmBkxHUCn1pMzOSip1c6AwghV38hq+cyKp
vPUEDHYE/p2XIFt6FAcl1IzotzLMxSI1Vfio77WyyXP8z1ejcm816q+DscWEtcf/xG5PxdxmBhmF
i79a7QXdoDDablSSm/b3JA+s+EAuQsfc1EB23ki9SeUFsm0imuNpMbf5nw7bAQvNaD0jfT2xyjcf
kKOK8tvn4gp7J1sdmpFOdoWfGDUidvresUOHXXyGxujxQxUXeTiOs+u86f4VL+fllhPfvENy6vVL
aBO4AWhnhDf74s3BTi9QuKhzcYow0zOeOnikHRUcovW102zBTRBdaGpGH/KWlz9HGZELDVAJB9d4
JFS6qHi9/QHJeVQtWK8uKsngRCitoIjkpi3WQVsw048Pwz4NyiY8tFPqlTSERDqRkkCJgwGLGo12
6rp/+YAmKVpu4TejSr41FjUS++DJ6acGLrXQvJwaOwqJyqA1+M5rWx17lXGEw77ZqfADdtOlcSu1
gRZVNxL/H95mM/FuiSXbfV0+/C4MbmjcWeQeZsllFiCAb3nBfjxN1L9RUL9Dlcxec4orPe+oC4tT
KxywPLFkJ3iVG2EAT4Zv/x1dcY7LDxvCqm2BJpCz/5nJD0ah9cJbQQmHXw9Rw6sz6n4wJ6U7/Jt/
r54+0UUxP6KneHoMBuxdZsYAOyYMMWYR5gFOayr/bXbAwf/YTusrWUh37ganV5WZmQ16enHXCjzt
gSeDqfw1Sc4RWBkwQ09RlGqWoqD4RqO9CrI7V/sXnN2WxXGV1zBkouogtJQmPhwP5lvtcaf2ZlCa
x6JEWQoLjO+6RF6zniQVazd9cmsKOpC19ECkbjMSrwaejz3XRtgEqs/I9KR94oHTAXfyrDUR6yDL
JpwT4mxkw89rvYzqtLFoT4omkcqfLFVe4a1EXoiDyEJKmxLPbU4+1sM5/rVRaIHOz502QjusF+AR
aLuKncprYTTa9PrTEoAoh1hUXRyuuWOtkakCouJuy45l4zCfhkiY7Kvv4jM9wYwXaC8EXvjPpk/2
iusWAmFSMw6Dgef7kDqF1VIj987Dt8OKu7T7ySCkXbT/o0HBu8OEU/UdtlePAmqI36ojMk/BGB8b
adzlpvtTRKwFIM4hJs58ui3khoiJgZKs9Cvpx8PbEU1oV24PselluKPY/ruSoYEYbG6N3v0siSva
nI/oia/mJehxcjpfQ5gr/eMuPvCMD6q1iysu/QSK1FsxHylIWed6XODjQw86UIuBniMTElxLTKux
ASj1mHWoR6UY6wFD9YvOFHsDuFFf9FeIKlYhgHrcWQ6z/bRjWO4Mx68PAOnNfUs8wHd0NsgSL5Bk
LbSo07IFGFrJ1lsTQMaMobz7wDF9B1w1PnDvx0y7kLIT5lS1l6C7dE1aJwfE/GFgCul4zjDZCvFZ
wviD8hIK7VbAO4W/4/UJvc9R0NqzvNw7rpyy/hJN64Z1Cqql2Go7um+dh2x6CW13zspJo48lqgre
ErF8HYxw1guUZ1r4tsNv2iEgBtD1o/NNeEe/gNNnf8cremnbvJkOWCU7//OjG75EWa3h/MmUlz1S
YUdIzJALZFwYZioLeoXOI23coEmty2SX7cNGAEfeNl3qO1rg2z9Q8yKngTZQNfbENkCKPcKJjaD9
2XOh8YuzHupipbBBBYpiAHG48an3WoIB7s4ZuKZMwQ2QVoRO+GnWVE19rj6pRvg+Tz8EmSkTs1S1
SOM5JemY5304BoHF88g+dbOkbWoAIrCKhBfNMMlzlpx7BmrlVtE/tL6j/58hrvDITITQfJwQkxRu
8PfiVB3PyetPtCVNHiduejyb1zT2uyKMhKWZKou2dZzW+n/eGOFFgkm+kReCvRQw73D4NkHC0gwR
1RAClHfSO5BH3g/C1wxf5lkzJS6md2/HxzVJF9iMANt41Zh9bRWz2QN/NJY9W/7GHO9WoYFGDRDu
zYp6RCqOQlz1XBX8KF3OmmYc+4clP8WxiwnsSkNvxEKMhm1FX3EKNc9mrIgL0IRzy/o4TZsd6qv4
C5BuYZGQhiDhEDPcu37+h1mCJmst+qiBV9fRbINsFaOiJ1tvhAUt16nRdqlfC1XtJMcE04ux2G95
bUvYNSLLrvGOXAdo9n9qTIzIL2FqiLNRRiKCBYkGzsJ871OeDHEThcGQraZYqWQBR9q6AI5EkVJU
/1mfjEzrOz/4qc0c0sZYYLjsN5cMXhuzguiip71K4AldJsOowBa1xyCDV7ahC5q34pGVE63VnCku
E4GJtyWAYUy2QjbrrnBtswiTF152Xbcy0f/KVQI+L4HtQZ7zzz90w2MNVCtyrcpjKjLRaDXujtKJ
nGpSM9x1CkpHCWHbACVIqe48fe+poMeZJ2EgcG2HZfwUMLYQ8YSThFqmoB0IgMn0ATggzPt/hNqF
j57ba5xQkAaZPTTkxXXJHw+ujSluwiabL2YTaeFszZbYzjaTYf3sV/JhQU/eT68c1CqiYD+2yUjf
f2IrBfahNFaaSMwzBbeajz9ogjqcTHgTV3mC11l1iL+YrB0gqrcxnzGzt4rga2nM2oEkfDiin8sQ
9lqA4McnSIRe7uBmoS7DCyjolfo82Bs7fbUdwVQaEjv/fIwJtVZLUnjX27mVkWi3u1xMHZcGSBId
jQCCXRrwuzf4/1QoFMpaCBoJ4k0dwgxshpzRSz/Pkng5HZhKe4eIF1dJVPqg+ymTUO1U1r+4Mjq6
vvBG82WXfJ2uFvZMGllVmpSD+JAvRQKBHPYMjhM7fu6hfW3gXTCkghpMHM/rXu86EqtDwrBar78r
rVHtGdNM8z8kuZR71IdNAjYQ3VVjA0rG2TZoDR7K5WMXg6xJTGJOLmY/wzXZ1+L0I6Q3kGc++9P0
CZIVb3EuH6wu2nqQuidzAZqpmyxKMlESyfHYtgbcfkqFKgb45JR9K4TtDkKGrldNF7Hm6T0qr1G3
5j5wYId5I6Ys9t7vI4INuC22dSo4zGPWcs08pUBxp3zlPVOwmky0KQzAZv2Pcp7Flx46jBEMv66a
KyWZaxMSLPcH6bIgWSjFXUhp2AmlB6xldz1t0wYtouDqPG/kyRbsEYmsUCmWhpX4oVGMdl5z16+6
BCbSVosueGrgmvn/v0A7384hmr+yZWGxrLYxosJh4Y7vh+TCMOxrIrgpmS++ojnAtU2B95wGS4Cx
zbnvRlVcRcDhgG1BOEGal6vuXVjiGltIZ5t+7/KaAwNKtnd7+Oq429Rj602b0Ch37JcqH9pUGBUS
1v0MS3b5NkV86Tw4P05yoeLWDZRNZ3azW4Or6Z529MIJouwSMqR+48Bn3cFfiIOsZVacu1MwKVw3
CSCsQNNy3KHwU1mxDPkijopyJ4MhpQRaum/SKKzAPr8N0k7b9rT7gd3U7T94qXIgUU+khTjI0heD
vehvhtSCHwVJHTTxAiT5QBEMST3weskxWVKncIujM8bVNrQj8t2LlrBVEwh3r8wJxsm4d8WX17mu
sR4RNA3Hpk4oVdRD65V0a4RUMi31OHm+RKyEodqm/f6MSWEj5MvWKQcZ+SkiZ874NtVBbzuA63Dw
ALM7J1CHliFaUc9wqZchxppEi7VmlDQLdhUEWZ7C8+5p3y4yNx2RfuGOnX/1wr+XrfKJmvpYKM5R
Wob3ih7BmsW/riTruNU85lA36tkjHaav+oquz6Gm7FROP9P6eAlaVtpY+EYPrVYDnKbSZJNL2GXN
N7LKcT+MozhxYBT2/8LBV1xcmc9PcvfwZsOngzEuPqwFTDm8VKZ92Eymt2QUXaypJoSUAT2RkK6Y
C7lRnEZ+RGlTFt0u0kOd7btEkJkw5G0p81ARiV6AGlvWzMsSzqd9Lfvt83XDapXXZf3NeGKL6Bm7
ejl3DVSe9JboYEC8dSknQBWxiCIGmo2I2EZ3IlkUOhiAViWFc/2kwKtxS+CHMhzFmdDjQp8nZaPy
Zzf45bgKPhaioPIv+YS7+kgpWskt+ThaF7dsznimZrLhvXcc8YiI3HgKd2jQMQsaG8Tz6nZdGi73
DKqxF2qJuVXGEPLAr5hwcHtQTqj0N9DhJZmSG4qgr5/bsi8yR2Hk6yf1dvBkANWCrmqZuk9McCKL
DglrwdifsHg90EauH9z1zpDeh1CNl7VLEjAKKWLWy0WyXWu+7eIv7C/C7vx+L+oc+WZJvhMHxcRP
saJVAzHigjQ9loOLpMjhzEiR6C3yPJnchWlNQDSiU3VNRomviB3YHXmXkZ3BpUzDJLVRdpE1hrqw
dT2pLFxg9bPHNZb1051TJSkmtqp1gHCES3VBP1KtJiArMRc0vT3sLiGPIkxXBbamEbKFUtN8SzzN
lmzw2ZwF4rpC5+C/YMzimcx76hkJ2NI+FecriJjGlg0DL54KLxlnaZRPLE5F1PTE23h5pMLot4K8
+q4bw+E7A3baEINUhGmUqwGc+c7iPsq9EclY2LUstH0cl0BxQmfnZEoSGdyCulTOGzJK/Y2tt0nA
T2J9q4pJ/VLXbCvV1lof10JE853de43xMEdRYyANTiwAzCCOXbwVNQRZ96XjjJuVd8fR+dhT80ER
5iku71v9aQ8J1whTrqT5S9NxXZhYHGXhyBr6N+LXeQSFug8FN/bgf7+Yy3fAVl8RzgjaCqxvNVXX
0EGZzxT+8BQ8K+iiOlNQcdJMfQFDL8dwcuKAB7wSzJpczAxBXQSIzSNYuG9jjSK4l3sTASR8Kd20
EvcjYgujhWUAXVD3Rb4LNf6oNiWDmKWNQXsPmibNUHzN4TDpJSn1HjHfuLddvauBmcA8DdiBJnDE
mKII+cd8SMKv4v5vNy6//m4SyU3cEwR+BYVYPHzN3m9ci6o5QlHLAqTGeK8uOA/RZWe0mi43VsbQ
55YncH7ojVhiKI+DakCjDH0RsLsQilRUuIrHfIt2ixGtzbWgHGYF6pW4FaYNCbkuiDra71FfTQKn
HIjH8/aezQ7RRUiWoG4Ko98OR7o84nwrNizGEmFpca2WppvDQbeyrvKZ3VJVmxkNezyfvD58v7FZ
zY/Wh31VPiGGs8VXLNNzajWMDhbojO5eFQ9wQCh40H//RA+8M5aYLMDLCANBCzOqUC29WyMee2Jh
kEMFJAfJ8cjSxQUFPPW4WrMkGGB7mBoVWQJfvK5AaLUSIDBdieeCsRwDVuO8LLLttA1aYdTB4ycf
agyHSKR8f5MFjn91SqsMSlcp8hdzidZk/JW2hgHGeCEX9946gY8oeh1guTOGge7GLOx1koesPOqk
wSRNDcIl5sCnICwnRm1+EwrH0yi8+yAMlo63aGPVDOm6mPQdAaXOwO63NzqNCEaSGZt7nCK3ImVo
xfq/hkTjhDZuycIpMKx3mrR4vVDBU5Rj9L5cvzfbHRycz+lDmzmDiXGXFiCSvF9N1t4pQx0U/Ksn
T5vNYnFfnHMq4L8YE/zFeZGexlBf2i73aCMcTjIo/B5JMkmqfYC5o5A4cqvxhWJBUuX1a5K+fzN8
NLVAecHrhitNGm52vCHRZCXhQn5T/WWV8u8R/5mHtgdNQEjxwzP43ws1y0wHAfPaMGejkB516yd4
DKHJdj/o2hXZ5Vw4t1VB8xUl0Dp0Umac9SJL6x2HsU3TNcIxzwwf05YHnABguUl23rtcDd99hscI
eP96ZklyLa1PQ0QiVQGkY16wApNmmv9m2nx230RPk+lmLr+ixjGvQeGq2k78gCzb//HWSrsktryo
yheCZytFWRlw9z4ICRptZ3yW3ZDv2yHvN8Gs9IODE1UPgtE8kHI8i4A7ZZjv9Kdc6dA3FtZ2VbEh
r5MjKdx3XSaWuKEwiijMcPzKFnAMNGY7qL2v7Bv5dZB7QBKdF/OY2AUxJbsfMz3UxldDXxRLD8B7
RnJm2lx5dxdt/yLUQ0v9gCVEA3vSQ38ViS1nHJ5quHIzEy9IahRp50/6Todf7qSGehdbmItfzdNz
skw+nE7rTK8/1PZKeaoStgxJIvwwAXpg4sBMVmrpAvOTnaYba1YDzAmrn5unbe5t7MG7zhbyc1k6
1PqpUg93a2r2JO0Rkgm9yTjiFgjQ/n+p18HmW0U5E20UZSyHcXDUNXkDlwvxEFbNQZu+MTwCcdsd
GNkYw3e9xiEB5Wz6W8z4ftrnhj44KAvDKKVjFkBKyAbCJczNq/hNsbBusV82eQIYYvr8MnAOV2qP
/eB9F3PP9vic1RpwxrkiLz9SPRkGjgwjjsy57VPQlu76t/aj5b74BzHIDVKoxbCtJTHFDRWKofSl
GljhRQsXkaNBlG2R0IgWDr1wNjj/4tBf1jhAk5/sm8h50PGpiZ6BQFaa/vDJqD1QpJp/6VnlyGJi
5mxRLl1m7FYV3LguqSG7Y++HBFJplRzdWxGZ0nqI5H4MxuStegytHmni/IUM7XCh4JF40lYHd8m9
um2CtHvl2jMD6zV8mfsKbfJsF9ncpUJMrRbqZO+lajHRyi5K6sIkoa8aTEPSHYa1stK3vfTbmSNn
3KXKGLPUpYcsVOJqftXJtRMlTfoAnZQjtFfCMOzl2PqPTXHGYap8vzBICm1Bo54PbJ4ng1Tkkldg
qVcT6SSCJ2axqWhQbO8FxJj6EClJTqC2nQpmiSGyGmVTgX/AdOOjOgwZJJF0jpqAqCSiSSyB9RLl
x5EIkNTlrqioVHIOYglU2Asx935ii10cHKXxZC5Hg+irZl1bTP58ck569t+bpiSyHGxpM41PVxZW
TVgL7JT8n9bCrwmOyBXIxu9PsbbC+dbkXUtvqogMUAKQPG/LaMIJJUDpFsV9rwph+o9GONbbCdVp
gnEHzRwlN6CFJffBJbl4O+eEaAHMOYsQoagZ7gbH40khn2QRkMFpY5ctW/12trQSWZD8zHEKg9/m
E32+/bCvrmYDSsAO2SAamWbe5n5ngoFneeZyCK3968qCXvRXW4+CjRudjZjw+zCRCLoDV/TqavF6
UfhatEnb4a9s0a1R/rcZo6QsSSlcLlntJv+/NOpdafufeQanVv6E68fxpIaGJSu1aXRMvCGPYZ/Z
6JsSHoRzsVFHNjxxjh+QimeTG/v6iNHly2LllDitCe90RjHj+fKrJGT+iO/npYNLt/qbNisSNnRh
ou1sGg2OIF/aCE2edZ1DOBN1oDPMpsc12El4X+ql3YwhDerI9XK4+zesL7qdS9Yj8m4Eq0ZHRGOm
Bv/DbcX6FIDTzShknodRkIKI6O7EKNhpm88uWJ0yT/YTrbF7NFAl3h54sGBPcnrvLuk1z9481c8f
y+8p6GaX0Q361hA6Jdelb4ILDQ9D4DhJUXvJMcQHSUVu16ciisv/uFJLEu+IMOmQ5fTltFpFakZA
gF6CcREVWxKMyaW4wK2AjgZjb3Jh4Lm00J4I9ZOHp/6c+/0IhZ4aJ/NvMVgHzeKlj6DGiNOC7vom
quFwQ5SUGsH3zPscyUwSJX8gA81wjGpvjntFb0aD5wcmtvkHEBM4h/NoKcYHDmDNTkdwpnDOxuen
N9AVew30IK/Mydj5527FLR+VgNSCNhYfITNC0LwzsbHU6E7aWnphPPzQzpiGZOCxQFHLmUirDuTR
JVn1dLDO95WSMxtjRmMB1fyW8fwOEbMO7KalphQXnlXMt5jVgcIGW5oxxslVbkl3SuN0WJDlwapJ
ymO+Mdk2VP06LFs3DT4IPy69C9GCO1nxnVbdQe7OyH9dIYJ5HjBryHQjMsGJrmZ26Vh9/UgjV9Bt
UyzAQy1B/HpoUugexLMi98QNwpETUWffNEChoT69SeLzujE3rNNpgYIt7z7ORIoD6mTGuleEt+WS
RXfBkkDF0gmHK+VFKye/eW6nB1MlqTPvkM2V5jdP3lkN7e3WcXQJn3EvTSSKRVNgqVMMZ8Ukhzv0
1IB68ZUwolr1znctKiXUxNg8RTdUzOXVUn7KTbp1KgbsW9b/TqTGnCrP0IsTGxLqYfBp0HHE2nEv
fFdcgaCsxfzwLwO+34RNhKleUdQBi9kG6sggrpqleh5SX2F7udMoinCW5Syjx3hGHikPI+LhwpNp
wsObQOjOLx82qUySRWUH69aGZftjKifLm+TCRi8yLY2snbiOhp8ncyUXDA18U1rPr9D1+dtPzmOi
HBGYskyySmjfTGz/dbq0dHeblmntOzkX73hi65thi7FkXFY91clPQLdPbYjyWmeWIPdCG+4OhKQ7
AzITD/bkqgGrLE8LEEYSBpr2WLsbImKHBJOPlDPBZNXnysRTmn0cEdHRHoCusOwJOqIPCbKSqac5
1A93rR7HFKUkjPOpivWnFE0vFh1FG9PIxcDFBjQL9iVnk6KPUdKaIYTL1AQBT8p2gLSArzINGhUJ
M1kDIEWQ2KZMQeRyX6bFeQ7c5rVK8ne2WvsGPdS8bU92TsB+iGyr9/pK+1gVSaCrctEMbcEnkeeG
kbY9aNGHP/oBuoIxyNdZDcMQvFjKGWYs+R8Usw3zF15LsmN8cCatv1Rk+EZrzOW3ZbTmYOVsMA0z
hovpE8z8gJeWaauxDvKfa4VzVOK3KnuGP7WIxeS7kHqnUD+6sJhSez/jAQrG31HgztlKhR2cEMaB
rgVSLY7h5RNSQkR99rtfpj4dG1Vn1006nRuIhX2PrTjD4CaSzi+1JisezP+B3RM7QZYS+MifcY7j
oXNK7ade+9qzfhR8yMtw5669OpfAIneFg/vh4b6v+Mt2FWyBg6ASZ1z5fhN69iPWAeXafetjeZWi
sUrHMY5lqGdX9sxyE+IUspjO0i1aO28wazAT3SwlREqvlgj6f5BfzkXYoxNz5G31yzQhFas+M3/U
kL3rDSBYqrI+EMY3pwbBMP/22t9nV+qWrI/LunD6PrQT/434+X6FSbZZIqceFfWVkOcOi9g4QfaB
Qm2DYesM3IS6HMqXnYVDIW6odlwSBwNGbRYZ5OKAp6K52zXICH7UuWPLCgIdDVBwrGYH5iuT2CVX
WdOrFEEsiXUiFn7HEB9B93sVx0dbMQb01u1qOsU+cIHMSoyKzdWIIEz6YpG3JjECOU3x4r7CTAiH
KLwJ9+QnEHyBX7S6zNI3+nnnGibQqgq6i4UWNCYiBNhJGwTp0+RgapXtjIbqsNjM+9UKr3SB4rh9
3ypIMG+LgvVgVMUjhwU0uFTRHcC0JU7S4vOhiSn9koat6VT+G3E5ENo+KBpH4ZE9063SE3Nf8kXf
RPy1QVDijpO/EimxZgPgiDx5SmSWRZYziI3wVNO4RXXwUgX9b13aN6VGMpfP5Sj384zpn52WMGqE
/uJ+EPZODGwPFOYGfTdWHVPIcA5wcuNP7JoanO1dxYNgy1RbQyUERiCxRbCokpuIToGW+dAP14n7
24lI6qcfMbmlIoGWlJQY16zs6i5boThYk4zAJRRXYw3XnwTb/nzMEJY9wOTUOMLzKBKYbyXH7+HU
72jIEsRQeFviCq7MVhhoEySfAMqzj/1VBgqRUs04KcFS+TD/RYdzU/8oq+ws3g3kJ2s9gs2g8iGY
LyWHoRfMXCs0yE5pi2nKCd48/nrDP3uBbYK9BPo1vwWtARY706jLkKFFz2O6ZKSCgfXu0VN64E5S
OZJKbLP5HETpOcuFhwPApLJ8NVLsFkQpXrXkS6kqZ1xFuw6j7QGPdK36GeViomPi39PerqssgpSE
5xq0g9eUs30Ikt1Po6pjtULim+MD3RjPtOvvORJ0I2VdxMCP0uml2wQYYUEpNejI7OMRgHp7dUCW
QXbrXHFgIAQhEfd8xIh4DBmyVl9Sv5nyfVX9YO5Oq2lH7sQOmIdxbk+F7XyWhdgy/7Qqc6f29tnv
daZOWRXEPpIPlN5VG/N6oN1Tfj2CykvC+l06qzxnvBjR25HQFBcsVsD1zEzvYr1dRshwC7/zQyqN
gx8FjIoA1oNXpOgfgeZgS5THDP9J67hYDgeYpMBDRTeColRXyU3Gt2UNX3tyy3rggElZWcEzpfk6
NGyBp5iA8Y2e04SBSO4exfmllxfj3AFMmk+79g5ZACKgZnPnGYroF4+j+PaEOVOa0YF/99mosDbU
ObefHP4JOG1/O1+6LogqbdPEQ1gFCLZ/ACofGoTe1uxRNrPWShLGGe76ceKoqtr26ljFLdKL8JeS
sOvWKMaNCO1GH/TFtHF4GLlKIyFj0vhdCOOwuS1CMCPtRM8cOWTnH5G0j6uwsFzTsN04DJIX/iUE
CMZsZFYet2UWMN/j90gWsaCb+1w1G0/R9PzlonbftcpE4hg06P8wyVaqmKPx9ya6MEuw0kevmtz0
MJL0uXz/RtlfkePbIPNW4o1X2WmyE7QCMimfjV2rG23PvppwNrBxXaoshPhY+b9lNiRUJRy9NThG
m6JqkWYR3uKGppCBBlBTB4L3xF1WpLveZnJwBR8Xdo+eMjmdo4sZHil99lwfqS80xDpMyxN2LUW6
qUAT6Y+usIbMdq6OUNKnT1XR20JSS/WHIeuqhqLnRReNBaOPzNOyneOIs+/tXXx5WLQgW0MIkTuB
NsoRvCVdKLzK7uYqZHlXV//MflObJATwyStwp9+0x+UKOJiHzM4brFsdZKyHFhiriVveULn/sWuH
4zp0BCbqsn1NNK2VwsfImuhCQceifK0ezLtyT6kBx0Ni7K6HxnxBufNfnUg66mRKMBNpzNLZMz78
/7UwefqjDnWHOccOr0gY5NKnZHgRIIe1wbwTytF/qp3iNgMFdF4dp5B61aGp07s7ysi8i0oG1hun
NISGDlk7I1i4qvjQwVaS/ISRYUGD5HYKAUrM+boZmhPcsMBO3MBWii0DtbfiXRURhm/inkod68F/
x2LwOh4yMsoJI7L/9ZJU5aASI93NLFxol7NR18RnRYy0M+PX7mqKZLH5PMJQBe+1HiCSStYKxcRt
YMmrwoJKjDsu0iBoxtFoEHEdT81R4TbbhA7BQZTTE6IZM+10ffVuvDNQ1LTD3IqZHhk9xqGgUWZ2
p791/FSKrzRrnfnh6d5aCAJXFqgLftcNKV5sWTTEwe1QZXmyL2HjQegQqp/Q3ms35UrRw1r6UQh0
mFlUateKRCYK166ZKW/xyBBs9LySmnBAWJIK14GAgGK4dxoEBgNEPk3Ef/uF9o4eEij4rM6ZHxft
CDzL+8+KFRZGeYk1IwLktZ0ie+KnYQnqrCRfwFL2cqm7On9B5iFZUVKyuREuCaWuZEy6YkHTmWs6
n4IvolwwEs0pBUlIn0jtG/RtMeQEyM5Ysvc06kI1yjjF7rH8PMY/UYul0aeFP/yvLVGTIUN/y8py
Q5A/uvgEEqOrHsLV/yDfVqWv8OCyphqPiWyg55dIMhYiedGwXSJzU+FhBMIUaZ3xkyysQ3s4lSYD
U20C6kmGTxfB0KuLEnCvzbWcs7aJBem8WIVL40e0IhzIfwh3lxss6yaSaKEk8mO0GtUEpjorOuve
Pu/2Rl2i7xNMyGPf8WN5mO571S895cLxnABHKhSG74dLV3kcHTBFodYkrKne9Q96zfEIqyrUJv8A
couLLzaBb8/RPdj/VuNfpf3Blexrg9hKjsCceCVFOLCxJxMqqgzj84bzYlmmQAIutXt452lP4hSJ
tL2PYVPAXp1r3rpZndqr7+yPYbgbBuUOhwhDO2lhJrgOVmipaZTMQNHfdCYemAiND7txhlW3Q1Hn
DMvLrwnFDph6QCfHysFVRL/ud3ezcOIkYNZ6zFmHowZKl7SmXSjrM1JTYhKExdNJkh6o/n57Mwkj
XRMvZyMzN/aMPcM6PNYYcRc+18bsPUu42ycPFM4qvkVMDrYjiVF+29HFwWeW87h/tifMa51lJXqK
Wu27sRubJJWke0jk2LrVeqyRyPj2lOHBjbclPmYKwUIIhhSJugmMdbq4OLs3uxxHogFnysKTSU+o
TTHyqpj38hX4yN6YD1wfojTEy4fzoqwIdDHfQ7Q4XEz/zAwqXMKj+9+TU+TJWrORpfFY3RAMJq2r
D3XWeRXuvu2AXAh+cMnlRs+dyKMzS93Pa+skxA36406CkDf1D7/4xtdHCTokkbKcsFbFDsQCWOtm
Qj2F6pWhqz74tzhiwIkRYTDEz+CdQh9ZaBpKYHGE8yM3RI6OvB7sF0EW9uC7WnGKZvbYsy9STErD
TQf9M2F/amiHV5bRFOw7GWRZY5mbfzO0ZbVdl3rgH4I8obTdDuvi+Ii+nGdqwdv7N6nVRR5HezVU
k9SBoXqyVAQEa6Qt09SB5yQekXkoD81z+q6ySLYWNzOy3wG5K6Og3POf35JiDK8nOeF3aK5uEP5k
ArW8tNkCs6Ak8wHQyMSHCNp8Na4eF2ZMsmS2B72TPOZUw7AH00h8hdapdJVClcXru3z0M5UG7hq6
jLy5Hg0YpNsBkZloNSTspPEkWJex02UWjREhEaufrvwHRra78FvDNoj4VI8/bhC4LZftNJGbXa5Y
KK4ZFKKF7TJXT7xfwdLAyZxqVfL7d2qcZzNW5++4OtZaDJgkvVvt0RrYN2xWFFa9frfFTY7prZV9
jABwyC31oe2WOS+zd9feKA58WolwwW+1RzEFmpPKjhNWS/CNqY7wMCBUxm4miAGxgWNoSalmU6hy
LVVqnJTPhPRvwhbTODELL2xvXNowu8HlN0EJ0dCe5OigXMrAj+0l0+AkWQl3NGp96D2cnsO9UiBS
RJWCYeW9U8oPzN+e0xE91lMtjOQAdWGFOayHWUOoiqki9omCGqbXz5WM2fcnOCkKuCq1gUSV2d2j
SAzSNF+8LFbvEe+Ewo+HnNSkCOGadkQeV0DZDVmYjQYvGDqq0HZgO+ae3MqzlnBuKfPLO3SXiWEh
/Yn5kfnXbLonU6mSo2ZJ7ayiZCIRVHsuAUOfOYd3eCwxy6Fh9y38u1HB6uMn0D96DM1hVWEf1L6b
5MvQmkF1fN3ni6tgL02CF7NYGgHbsh1Ov7f5xED6oJ20NQhS1OdQ/BFwKeGxu3uLKKY9rkxFwEaU
55I+gR3J2o++ztiFPoIAae+Dg4eyRm8O3v16CMnkqi65WjwPoXKBnADcqbncVa4+UJp6jIGJae70
KziiOHOwb+3BFXygPPKiXUrkWwyvN0hGRz0E3egY7ntimF6ORV6NKtAA5XxvyGxr6MawXi4KAQ5B
nFZH7TcxWjk8lCn7F5wT1DcYSAZ6CERfuV1KizCTEtHde/UgDvtxwIHEuoozsK2Nlo1SvKV9qbZu
+kFl21ZJmLGXWJ3T105XUDaM+kAQkeIsUOInkWiO4ICBvXIC+I4JCkBdIi6jlToquZmM1LP41yVM
jd1ShITaQn9Ta32pyyjrekzz3aN68r1/B2LkpzLpTnaQWf3xb3Pese3t11lQ9DCU9pdYZI7H7sXX
mH04+/2lay+omdlZUdq5M4v9Hx1pa7dxxyxue6y/kwnWD1tvCLnz+x3jO4tBVS6CzQdMNcq9TpZx
4jDBqTmrqVMsZoZRL6kwIgXxt10qtznVjJwN3KyixL9Y2XnbYlXoJfrHRCmUTB4wq0IYjteR7YiB
WYrBVQognNZqvH7jLDkMeSx9H3OfZc3Wyi8T7AE7KLiP+mob3k8vlr+VrzlbmBjfSPBvj6LUGSU1
WE0RaPIehcJbH20uIxY/8azGTsK2EFFPywWLHc7cxe+LJFKoMefMe3BLp2StaN0RoG3JPkSFMzrP
C2Hw3pSB5eBOi68D+4vDOZMzBDhupN0utfBoCmGLfVL54o3N4h3k2Lx0ih9f0R9zJNftez3qwMN8
4pYap3a5SAYdB4IRZIYRifHGI2MvzCf2/yU78QKCOwkOdtuJnfEynKrsoMJiqRVl6qzpAFErmsCV
zTnpZDZ5S1uQKTjMtBNqxGXG7KC9yZqZ23ha79taKY1VfgKaEl+v5a5X9ocxa3FPtkkxLvdIB+DO
Ec+b7aOm/dndt0N5og1psa9E8itn8jJpyfuvZ2pZWvmaV8FuqDQbE0cdsEQllzfgkeR41F8r14vY
jGc+YR6A0A6Gcn9THuMnid35oWqM6SKc20YcgtemnHLBb96Kv7bb/81Z6E8HT1w1NEQBX37lE4H5
W17jQQYngCFUnN/nF5uUx4Sh3pL1p8Wpjh3RbtxZO4DMSgauT62r4vcu0O9aJjc3bJmdK8LxEutf
oG/rSDpFZrZi3UufwU0XiEXoI7zzFpwD0/MbRTxietK85VufgZwUTy0DWDFaIW719fW2lEu2DrzB
fAG39WEsIfghwHyfa6jGSBC64ImsMMBk+T1owgYVxWW2R2sjirsl8HoIIlW5SXqre+rDrCKYlg8F
EFgP4Ql1IPD3wn0IOkzxH6tfKT2Q4HukaRk+R362e0j9IQI3WLX4tA7armheSgV3sVIjMrrz1XzR
G6AGVuO2wd7f0lVAmiIhSW3mSO9OUCgnGcaq6HRy8+guiAjvCr/h+SjWiSHwa1wQaHMHqAEJe/NM
F9ID4fmWUPQjyYbtTA+w4wFWCPR+aIAyOp40Ar2uqiX7sSmMj4PkrWEZAESn9SJuEraBSOLj8GaV
OM+0m4K6ri4POO8eC8HNPq+YXfOnC8mn+261sKZku+McSe/pdxgyDYONYJKqFga6GMPRy2wZRIi3
+7TX1OPhBNbd0xBN3j/fhAlH2eknDek66IReIEScsW3JElPaKqDGef8IbWXq7wT29vu0UsNGm8eE
KbHsTHCLQrE41dA1A3w5Dfg3SAU5SeSsKGyYs2dxvEcFlCi6lgtccraEpjer6ki03VDwuHJUA9+m
DsLzAcQMwPyesrFTum4ng+0iYc+uE3o1t6cHQowpEphDK9xkc/MBc5H2ZRziKKOEDRnZ6KCigbgV
PmyNyuH8tjitX79ned/VLVcTIpgiAAizJhDCkKoxCNvk2PGqEI8V3vR01zMKn6yElf6xWlBSHSa4
NJxacmFqAjCT1+56hJEx2yla5pW4Qzljt+pD8DQQ9nDWEu3i3Wnpz8+mpCFAZHaqqhwfT11v39Op
7Gr8Rlj4ay0MUVMRDg2Ge9+TE8uoJdVbuz1IdN0uqVukJrIJ3cT+teLLDxaa+Gb23lLq022bPxqA
/IUKXvuyFX1MI1QSSp9G065JbsnBp+a0ukV2Wo4WZL7Ehe5NoHwqu5OynN907MCkrVcu+7uKExae
SFDKJRpzmKC+gJgoVpslvQziOR5xR3GE0rzGeT+dOy8eJ8VTCTnPCqQDvhuWx6PC73TCqYFrc1hR
6NTBhzVc7rE/NdPHgNNGJDpBNxY2imRShrVrhPk5KDfCQ8iFg2voEVwJ6ONI8TFa2sjyXE6fQ6Ds
insZnSBrvJZFK+VhhNWUpsdET4ZWrywcLA5BSOXJ6EhwG3+toP/pVCwtkB49JEyI0e0RIf7kjxB0
YS52K6VVDSEHMoJg+J/kTlag2kBdQsNtTgZu2UaIWyUfZ3I2m2tI3HCU5QJQ3MGxWY+2qd368yPj
GA/wE8/+psWP5uout5W7CThE/D/kRh0/uVW57IqYp4yzPd7PkpYQFytCjbVbQ9FKQeg6CVq/54Ju
C8wv7MZpqxijfJMwQ26u2Ki8hd+3vf7RaSbKUjSLR8fMxsFMZKRJER6tEZ4K2aryWdVT9s1sdnOX
K8L17cH95I9v1VgH7cVCoD9sYzX1Tb0hbNxJUrmpYxYVhiuqH2eDKaxSTVKsvbpoAsuNAfonA/zR
tez8HtNrbYm7IofYvNkziwGN5EuYuue+EVJtBPgYO9PJP+XpuigK4YsX9tUqMW+3jyhPc3H5+z5A
6YFMYfkMnN37f2r0lQ/EoAXmJNRuWJK702gLWB+prNATxHWhV39oYd4cBr2OcgznKkC9kjSc5DBf
rTMw0tbsKGaktfUNoGotFORvYcY1E2ToEQZggFgORsTgqqNMD/x1472kcpdv95bPk7ccQp7iLfV3
NSbHK3J+uyn4WJ/tayqlfMscpinOxDvNkDCkBW2Z/iqC1FoVLwkxhpGrlXwA4t2flHAux3QuR4cI
mT5Oo+RQTwIy94Q5U7oNYjREsW1gI5uZ+cIATcQ0kkke0AY/nh+kwD3HVxhaRbGTr5fdO2ymrORV
1v32W+OmEa8K493aSjVGfartTo3gJdrbHOBDQ6Qw3JLS9zj/y2GWbcSh6tbPUtFwGNjReKaeCSiJ
agohBjo9MZdK4EitBnifhCTDHG8o7ohpRw4djoggPACkOY9a7YT05ZnOz7u/xmR3YPDq2UGGc7Pc
C5R3yTUXx5GSYg7XHuOTBXiu7GoNY0a7IyLcEm7R0BCJWvhX+sIeNrqb5XZpeIPQ0vo8NOPRvAr9
a3jnGoBK+dWVhD4eJRk9PiSlYX4Ksd97SIgkeHaw8gmLdKvviTYlW6dX2x/5z+q3MQLBMUQV0SQo
uAlG7XNwjAJr5UUZD/cB2qbCEztflfeB9wlppTt+rSY7e171IQWzGwoA4CEXGQjRJb9MnhLVjlZH
NCy6Rw52cECdPx4dpMRlieKTtZQNi5P+quoBjJY3EPxP/bI7mblzfXwvINBU7zKHfAdZJB1GnBjo
8ukOHOjn00UqM48x63+Nj+KcgA8DSyBuEA4QAZ8X0CSIlORqH/pOD70r1nUa+MFZ/t9NsXQKjTqS
7ikoHflFBNK5XXK4lj1VhFvn+Tjt7WV7TzTxbNpc5ZMRYOwpGyKpUMcyEm8VjPGE6evHPuead9Yk
gF0k5upLiCzIqmSnU7PFDIkLMdeMSDazAULJBYBGJQPS1DJ7VL9WgaOkqLZGX8AB607EhwND08KL
qpUjZqrC7H4w/syEbS7c26ANy1AMq+ECHfXdk5sRQTTiZnjiOw5XatNbBRC+QjeAVglxrC95OORc
FCZkeItikb1Q8eDfqDAoHQ+QNkPLBPazKJcM0eM92wD9WWRPn/b4E5WmjStAVYWWqlIMc6b7YB2s
XuRevQlgMSFNy5vOjEdkj8n/6zCR6vjEIiQ2jgVgwzO8CIGJGoIhGjoSu8QWDxVrLf9J0jhYWf6I
JjxT6wtYk332Y9+i6xFkl8HHek7l5KYC9/5NJWx0tMEzVdvA3o2vUIPGiELK48GDNKUeXHmMQ8xQ
J8KhIWu5xxGxTmJESVFIXcp8LXab7jw7WHrIunY+7+ABkQ+NFTs+/68l3df6nsHX8nm+urTqlqWY
4OEaLU4RgMpp4VvY5UyuJcqjTIO+qaDQOhUGeBHtNm3NTZc7re05y/LgRMDiIBA2E4rtBwlT4m4O
1eFR1RQ/48oIijcp80fbLgEbz6EbIaWR7AsCELOzUj5aKuVupvwIdK1vSww08zGMGNNm9cbyBlbB
5t3wJXeD6yQOQQME11ikl5vCp9VXQjoPLEABDovmuEw3XCp5MFkBKoQH5Ym24kaVZIVd83iE2532
WEoeIrLYBbYrAjiCaRRg3/FEhJ2yZPdvXaCnn9Kp8xmwG01NLHZQ6OXqY9xj/yRaiyBvvlVY35du
OlQXP49RNmRC2wOV0vhzoYxYA+IhcxtPq9FLYNy+ebxJ/3J9j3NognFwGBrZ+611IRjdHrS+5Imr
jMcjgDcd9MCS2fPKY4H7m4U53x4NNwDPBfpO5QMK/5XU6c5/LEdbRvZ8E4eEBhS1AZfY5RDCuG6w
eBEHwdtMy98YpRtvkd3PEG05POJu8JVbhJ0qE2Dc1ZvYI+zJpR7PKxozfkpi5IJtwqo/Du+XAycA
wGFV8jm4ocl0AleRQUHIzqunNjRKxEDhbVTAous/auI0WcZezwgGkDqdc0EMEtfV+qEAoFJvaoMf
hJi1kRCpXQRnvdKXcXMULDZy2bDxFsi2BsmO4Im8X8cnOCjsgLPM3p+h1UST7k+fKg9n6grAiAiI
HyqVHi9ub3OwZys2NUFH/q0QyeacACZTGdZXCSbHHP2bRlChmF6cwxQWEL9o/etNPj8CoBSe9ihh
bim1iBE2MDTVLMz33kAyjHXLJvwJHvOIRtFYvq67LqGNsOnH7gDWUkYL+Z9kOH2Fd4YZ9zskn+yZ
XAy6N3uGOZQ81wq03lbKHMc+bs7mlL5sIpK2knbBoAdJHNyqPTTH0OD55fq+NQ2X4HCa/a3VgOzi
dsWWvtnmBAld811QOTHb3oFUpppJTyj0SPO3PfGhmuKJJ6IgULWIS/QIXzVKOgPFXQgtjXsMrL3S
5cV1FACHrkojV+HB2EtOZ4jaQdQU/jP89wIKRZDPdF87/6rfVU4ACaFFEFmDQMjPG205IrX7yILG
AjJcZFJ/26cZwVFaNKbVYycMRjRUmMFhPCVYujXhBaN5v4urwJlnQjn0pwOa9BJJ3IT5eeRCtiEA
TZnhTNAu16TsaSNhOIK5Wfy5n4jHlfFutT83V+vV/LYBLL2Ql6pBZ2C7l1bHMTtxezO3Ym6fO2l0
vW4etkXbBN00Z6pFs/CK0PCr5o/mBD+y0g7wFTIiodYbJ/KPD2yGDjnXaP0zDKxV7ZhDyktlhkvU
ryJLfxQ5jSgFdrz4Gx2ftVp40UvXdIp3i/+19LJ8WivaTldO+l3muTLXnosMc39a6DldiPIfeRDU
ZQKaRfmrQVQKsU0IFVllE2yZkHGqKlJ17Ig2gOKZLCsQuXjCtyD5cc1q2JRkG3bbzO+KhYmmDJmO
EiC2SrI4MyQsHLYMf2uSQSSTbfjLpyCKjYK26p9IwlPJFY8c30xUBY6asWiImjzk87brORQGGHlu
yVHwkCcf87qyTMPghHDZZ8pvMsGKnOG4T31pzQtQMCJRXF9mH81U8+tC8jnGCQE3aXCSIlHG8miA
sf5PohkeIpzcNI5mgamXJU8bXdIK0MPhfkrWSrrDBQ6ZnWqqveBA5ozVqGTsDASKlbRPG9K6ajFI
YJj7xCaIwvxtFkuKO2lyP6zKmQxr7sw7TYHdGh+tE3xfAT/2zZ5jtuyaGhSotwWfWqE0iSKwXkYv
QlFT2c0h0wZPzcxC4ySZ2/A4wTRkkKenUFu8mSZgok+8AtYyKpeJCU9qnnXtx6Y4z2E7cWnob0Xx
dCJe/y1QjvVoi9AOpm2SKEJEx1V6Y3NAk++uMrOx4wxilHH78uN+5Ds4/BGcnISx5yJ08JB2AZ6p
IbaB6uS+YJC5hF3DAhd0AXTYJnmKBEDbHT5kpVmP1ImZSWjHBcC1ciomkdOriI10ARJve9QUoe3O
MvCd9rAHb+O7DEbOildLF/xT/3i/xrD5m6IlwGnm8NQE99WaaKrDTu9Ecf5amc6s1nsbxjRVVeyR
TQttlzFFLf6WU40nB80YfA5UvOXR6fvnCiRQJv7jZBrbavvIhE5UTNGZ1OpEq/Fgc7gr6XV+ME47
4P+97LbleylnDWfSV+SPcKK9oRk6xwdyds8AOdP5zxix6utkZ/NPBqyHedaTXa/jqQ5oNnOtghAQ
0yQb/+9r+nqU/s/fZLZwR1clrz05LXEdBg+7vtA4TERhut3ucD8KizbkBpHki8zFrqlZDZHftZzX
ALZcs2VgfnKWH7rR5uSHlYqIDqxseERZvAChkFSMr6T9znWvYBqVtEQOj8H/Uc249jJLsq7ONOsw
Zm3hXTw069hWhDFIje5Bvfktwwsbdowm4uymUTKkuDVKwEcRiRd9jcSSgUgKJ7Pln4J16yY1hEJ2
4YNjPNV1JLxIfUea+eNE0YtDwfFanmfQ3Snd+GEq5pLKeIjg+6hN80uEBDqnMn8/cyzdzi0ew6sI
iliETfNnvsjFemUp2G+EFytmlIuRI+Yl2LgeapyRRYXMHNfP5lPKxRYKK1B0Wt+MQdfzYGfiUN/h
dtBqaT1vQOuSL3rfNvam4S+LoHA4P9sQehVhFSX+z2iHTnuRpLsox1cdXXmFMuLspCgv8d283qzH
oLKWCNDzNDa6Vh45snh/9D+Y68nggoTZNcGK3mRbr63XRh6fVvBFmQqXzUocXM8nXdRycP/KfFl7
PGEr5kfaNSKJQ+6dfQEfmChW8D8iuKecxIzAygHohmprdAOXOH1FWHj6IMzXy0iO+v1u8v8XZ3LN
qdtuDr3K/Oh1QdD406F1iUeAASXecILydd3hyCKQlo6xKsW2nY6Sk1PcqtinKF6EWbINu3yiD+Yz
c+nkljKukcvrErrkOE7oULQwN1c5HAspCoZ8Dp4gC39cmJ8j2s1hTvIPWwm65NJ/qctFVBi0ujZD
93U2vuOM29nOiKyuLGKX5c7UHDXUj7zxOEHZujxJSP7D2JT7wtEQ//e/C2tr6OsPOlAExFlsHcBg
haX3jAGQ/olqGThH5+kz8tkphfdvL0rUZ724MXbv0OnqSydoHmCjRspl945q0uvCjwc76YuDyxV7
oDdXGDFzwK3qwPQChZ/fVg927iZkdR8LENToOoBnHDEV6xJfoDKbzNBO5Rd2x7mnwgkoEPeE8etq
7an176qGI/sTJx7PdmavO4aQwHV3KD2kOanH+FmWnM22RiJkL8UpeZRzNSyoa6bjG68RniMiKc3m
CprYBBW+dH73pQTF6mkar/cBh+UL9STR/Md5LwOIXpRGUi9Wg+hnPowjP1D9dcCiKpwRt/LpFqpI
M5NsdCXBC+MGA7EMHe5I2mh8X2k7xnMq5ENXH1sZYs2YmD14JTfitekKtxfgW49/d699afC2Ry5s
WZu2vAI9IkbCq8fXQ09xA1SvxPh9l2uq4MQejy919qB98bl9Z01SFBaYM8OFRyPBQ5hWHw3hZ2Q5
VU2OifxYQwRKdR+yl87DQz10Tm+SbZPP2VzEiYA4VhEjPjDImhssyblIwCt5t3oE8fKRjWzQ0BaF
WAhKA4Ami54VRpRNwbNN7sBW9Cqa2FzTYZBRFP+6rSqHLiq69utM6mSj8y7BaV7sgpVZaal1l3HQ
BaZSsomJa1AFNtfJkTvtTuVBo7fLvBIc6uIbBSq7wZCUizp3m9V70I8ohMpL/V/R+IjGqiltgfm0
Efua+92Hn2sH+YvNc9gZTbNJm6YJfLnBrPcU1wrdbDkOe7gWVJsJl4q6TTmhdbUNlkfWzaJtlusH
dbQePgBe6ie0VQycvT1OsVuE0nD2NTEZTj6ocY/dRFL7/LLvUnB3rBsPzra1TjatLYAPve9R7J+5
bZPb7CrXLHtGYEJQnyT2ySGfoSWtiEZAPDwQJ52XKVM3/TNpKwtjP+d2V8U5wP29ED5zakoxFfiC
ZBSCoHlgkgPhUnRZ2xsIm1f+bckjNCY2Bg3K0XTezhGbItkfch6AOMqaAPKH689NW6ino/TMDuYS
XQEwOPDyXe2y05DfK4UJyX28BEsOWZXj/TbXj3Hcp30JjOw8thu+LVG8OCfuGVINsBWbJhg3xc0O
LmCl+mAJ4k1quFRPUosYx6DAAvNYuBscY2rFCEDnaiys0uf5xATf1JZA1ZFp/+izbTLsRwMk6PqN
TKh3ArBSpbAJsNrtnaNtU4es4FOan6Sek0DuZ2aM7+FNC3vQJORcuBSMrelxP6fpoxxebmYoLzvS
Ok3Y574kBAIs2gfhHHgHSlZ9MAbMhD3w+OYZ4nIp49c+y1U+tK40tCh5Tbo9iuG4TzDm8tAKXcmT
SHhKVdVmboUZtV2nh2jS85fL2IGpYqwcPYp4A58GNzzEx4KDipbr52Y3tiXbsUiYntR2NwXXp47q
Zw0cFa0KbLE7BpyUk5BF2MuugMO8SvUeJkZhqjc8OT67zzqTJKqxvdu2OYs2khQyu6tldEQsED1e
SzmCHx3Q8qYmPvAqm34O+9NFaVVBoFM1Y8MqiOfXKDKxWVfYRhhjxgwD/p8eNxPvKfDge/t4Xo4v
BD/1tLyPNnqwtelgMxLsyHYK5Jt0NisOM0RSe3hkQfWnHAYE3AmwIILba2ZQ/XLDjHdPQRYp2KSf
PUr/PkUqGxB/6lSZzKJ61+fA2rNLAYmI9zpcKpZtpGe4V9Zam+bOloJyZLZ0b8JNgLHTk9KQ9riq
ZILHIdT+Edw+WPXVcl19Qqy2PQ+XvvRKqXsrvPgbTUulFJ/CSnCctYmaoRGpWBdFWvsb5Q1qHxAp
0SW2yM3BNECAuOzH2pH9HYXDUnuP7yFKknPbW6P/9Ch5NlyoYaOWYgYnz8b/P0QiHfgabRRV+Can
he8DA8F8126/mutMoDVWDRnRwhDMYobPi/8kMkMkU5obosQvNt0qFHt34J3qiOeLu05Pw5WFPe6d
9ifPNT4EVOjRRZ82hB45SXWSrffsL1l+Vjf/+/k5+3uMXVwgla/OoJccMmXg+V2+kzCmoUo4Wnrk
xFlNcZZKGZBouQdzUEiNntx6e0ce38L4OhZdAV3idLYvaSH2Lu1FuP/LCEnT9knQE7xojhN64AXI
XQiZhi8zCg6ANqQ67+l9NIRJHvk+3xc/3yS24hv7FUip7XCXA7ON5SRgJ7I6Hs6iCsoBTqd0Bksw
3yKx/+1AtfOx3VFGwY7w2zKb2ua6zy/HvKrAB0jjAH8ZbtqnUOKKdciI+JnNNw6/0z6RXvkapcDR
rBAsJ/0VmyeWZltKjkmz+rOSqKrn709J9M6fxBXv+ruKkPksg4mow2PRTVsfKPtTZKkBGRyP2ykI
mDfs1/oNGewZ+d0QkAtmqadpHI+E/syaFF632osnFjgMqnZc5mGlqdLMGzuPfgepia4lWazHcLwn
/IzTFrNURoV7Xf0Kb/uMQwi0T/SukCIJbuYm81Rn3arocbYcImJMjcycCUtkypuHNz3kY6Rxys9q
rIzV21HJMKq8cdpJrckZWlSxcazojlIMlWxpOKJGgW9chhWih7jEdZg1kbA1fbQqo0iRN/fktFyJ
1Xk20/H/TcvlEDlqsOBOU5Db5PGTV+N9tY8j67pinPp7c+dz0ZhNnb1tEAoNO1AZMAUxshL6YQyY
/flLgIAyZUNGN4GEncujULTSP/U4PJZZVtbikmB8ihNSUK/CJexwvvaK38QVnX7CyUTPWvrqovFl
/zQ3IB+f+nkjV+14RcyId4B7OFDKD2cbyvPKl08nLlbJwfY5PBRofDUDcqlqASR/HlBzkNieLLa9
QmL7zC8LkOs2h56uxk1r59LAS9h04APa+bk6bQTcrmhjy0LV8TkEBaMiAQERqlGDTXS/7GXbwtrE
80BwG/nAvhypcoqRDzs9gIeUqI/4yakfrU4OXvyl5GzIb02dyaFdbwOHs2PC1R0u7LxrtDZDzQXY
J3qPmZUznPA1KMaGpyv3jVtOqOFQ7SR5IvW/cz73JQjTG+U61nH1oWcn/nLxdX5RqdlAg++0JgMG
lrSAIN1AOTA/RyL1QU/G/m57x4TinxPdUl/akzmiFXY+xNcXOuc0u1vaS1dYCe9HbtL7lLvnhxhq
SuF4xDuglCOPM+Ogk249K73nqbsJZ3jUYQPvM2uwwLKEUMyCKMaNaeetzMD5aipCcNIuvrbF7LcL
Aa4Sm917YwrsidKzY6QOtmaXJTNTCQCTfmDqO7kYMk+Qe50W4gJFbWVgxd/FQlp11JJpxbP5abuI
DXLQ3ZVnsRE9/ktLU4DDJKE45gMOXXv+lQ/RD/g/swYRJsC41oqqJ3A4vrh0QVJVtwJPpRtSE2Cw
5ujssYTkJgSWuBx3TOhBYHqcQXyDd6zEpfQGqamxG7+9n+ZTceuHLCgImB2sOPw7GqvFIm4ykCiF
YmUDV7MIvFLDMPSc/Fz7M+Gpo3hMgcvC0oYvs4XDiby20ZbCz18TgVnQU685vKozn+aP/FUTPj5O
EtncsrDyPKdL3qnn+hue0S+o5+yF8XRsbn2bSYMP4xdP3OGlZlj1yUzAh3ukkMfb9utAxLrLl9S1
ZSRlBJlLi4zNZvgXnmdnLWUDYy2fMTcwPHPSGRYRVOJJfLNo3Wfi17AL1o42657iZ0AnfcC2UT5J
aSHG9xg7F41+cYnzDqMAt+Dhws4yHg3+nW2S9p8XZkftR4ZU9vBspDL5274TBJMUU+zp3sx6OvXd
L18SuFhlR0GPbDvS6sbY6cGnnVjXdyDx/Z52MAYN/QeSrHA/zrX8C3Oj/mrQPpDY0MrKGQACgx+u
MP1MEDKUS/7rd1YJNB6wAQAQOnyPKZi+FVtaAScKnnN/fsJW93KUjTCbTLAsbAWPtgD3G/B0tRqh
Csoegk8+KII504R0EJ8TCduN9Qa1Ef3O+XClRanqrCRY8tDslF5jO0y+XBCBu20AwKam+r/V0Wew
yO/COnogTkN2oaohrhQBtIfB5iSPedliJPYfrdYRNoQuuMuSYgHyx7SBSFwBCByaAEVvE8ff5HxN
nb0Qcj4d/DODIlUg3/lvBQaOL5eqG61zbcgJSFfes6vTjnvM8GLPVUU3WznbfXo6y+XMqWaf84ih
fuKehSizq/vB1VqDHUD1OcnQzbCYamD1j9TXA2F8emnEFjKhl2bpzkCLfIYMyFVKrHg3eOz9BRXW
xkjN6uPFc/ySTbFzQmhQO0BP/4jkWHUptRa2i1pSJaWIan7KGgfTA+50KSDKBxD53oblmSmBXDAo
nR/SobhV2pVqP5N2+Y9Om8Q6BmWIrDLXtn1JqaKtP/P1iCxvSmTw97hsCcB8YToDwuoRgTUxH+71
VXYTf8COxhP0wd2MpSB0TY5ZoWp3TSCUkwzMPRPtiqWKSSDjoFV0rB6/E6eGVbHGun65gyx9J7RL
sGVn/ATrPBr4hq666c9eQ7JaRBSzEcP4QhvbV2+KcuYlR+b5JBW3SLc3smOAu7kgji/z19Lm7Xnu
dib+aAnp5sHhyvDCfw8Z37dWNTCEsG5qG32X/NvuS5k3wvbxCJeg+EfRGWJJURjOiM/ce1ZWqSLl
LXwTMlIymQwCKIfcWfOzfuakDMIPrJg5TvBpzObZHk8uVDn7weIJxcy6LaMd/WkNDJooiwvSEeuo
hnTExewXTyDmFuduvBNnATJav+bUY5OsLMYasDK0DPrbphH/f754ss5B4Q7hgpJexQ1RlDzFw1jS
Skc/FC5sKOJHC6hkBHAMCSWh1Z9l0E/ZF06SyDXRRsXGeylBRNNuMJUg9uVB7dBFvouEw1b1CT2E
AsDyjYBkaCGOG8gtpRh/JhixBGbcs2zMM/h7WoRsRWjDsyDZD1sqptXPeeFLks6Gl5RRf6gIFUGS
V7hcjthLbk7rsv+8OIofFZruWooYO14gBF3If/Y+osOiWmI9DEWXdWxAPgjBXM7d3l0n49uRCNio
OhnxvjqK+RaE12B5MxFTM0NQhVUrA7VwRVr0sOROSLhHSy/XTJN90/TiYEGIH22jGLpcrz7tj/FB
LKo0Cekza+iSk0SP2U3SnQ/ngAUNjm35gbWZnvIyWzLVwTflf1DcCrkcYyNHb1cNGx+i1G39ciXT
0//e/VD4/1cZymkB5hFnqd7QmboWSMJg5O8NjuZNGb/ZMvzr+jKPM7alvwcT2bGY2t1aUIkAfCIV
2FnLWZIVZqrO1cZwQpS/7q2hoorsBAn9J/R/pGwq2IXOsnybNQj0B/9/TlO4VHZO3+QLx41TXXYC
TgyvpfBXNJRmJeSlVRl5MN5iB0DDSfioJbQNIiAjLJWzN2TZUGqiFFJKAqGE1n6T+VUZdg4A0UAu
0906P/qKre+hYb+MdAR1QDkOc+QR+xVVlHfKU4qSD4yoeYTzedi1kmXmsGA+Dhp+LTtqyiIs/Naj
R4IZVi8dsogRyH0bb29WxwLzwD8vrPNxuy1iYYFYpZHNDqYcU6i1sdsKiWxAjyXgXaqF0svJdjJv
mDymL8vqdzMWzV3lYMVsL8qz/ikyG5PGO06Y5zcybmD4cBWLC4sMPDczCLuWBHKgcZwabxv00pDz
jecv9lkFNDOcp+mNpRRDq+BsUA1OwqfafYBUNTsNyShzae5gxwq00LnaI9FRK8BatD9H1Xj1C7L/
r58mKlfJ8l75HXYHuYdAULwsp+TqIm7mHmnsVWo+4yfl6KQhz+am+pdRkj6sgJdH7Rk3CeYxgDSo
fFGw2mjOhdYaVyq6oDakWuCsFZGQMuvOg/U5B7+gf0l+AUeyFgB+sFECICuX2L38OLViz2hKcdk7
GxrhQuePw28smF9cVwHot9iDZTp+xN0bHqvJP2KEsIvHPlNU7bKh+mQK25kuT6Hvdh56SVfA+zFB
PXmOsP+h33j7jyhf8M9R22fxV4eyxfk+F7Nf51JM0g4IZMo5FW6pZM5zYJJcNzikwk48FcdQTT83
+8r5xNoYa9azgwBxcIxaFSh7DHHamDsN4wyVe+HjvHBW7WgAcTsG6Iow68FtvNn5pcRi/HEbEk+T
W8OgYY/RAl7wkxB27WTmwYcuLx0Y0ILqyb8ck+cyB6/KZ2+Baa+kyO5kHFepxnpP0Q3Zdc5bei4i
lVdvuMgP3n6gG4pjyrcsKlklwIYB0t1Ik+PHhNk6TxR7pED2EGv7zFynN7R5fmt4vP8cW0dITWjP
7I6CvOWD7kVKTx4HnQdyviSzQXae8AfBgcWE5/rHFrKklSPQhft5/fn5MOlV0nZI+cwLKUUmQw8Z
ybqpJ8MDj6E0vTWVskO395UhmBWbadI4SgWwQ2sOb+vPjEDWmfNThzuyj0V/LkheXqate4yGVrZs
bsVX93LpIhKqeFKXyhUpTOfdtCTrbOIlxNqrlCmubv5FO6LAji4vNpHHIWDauV4Qe9tTpsbr3Zyr
4QEerRO7V+kdL/WgWwhhKY902lvO6hB8IdVbIZ3+p7fRtL2Kl38eCq1KV9mcIozG1qgYydnglSs1
ckwiZ8HslqguKkPSsScbUA/UyOBm7z9dLYWrDa4d0KJtAUMuUx7BNjSIEgBfD9YjOx9kdIDULim5
CRHcsSGFX94FuN1uUfSA/gcAtAjFVngW9NoIOkExqkYjsm+lFxlIramJm3VVI5asE17AXtemz1kY
RM8Ls22sntGT15cvtYmdIpxo+veMN2nxN/InHdHpBjHjlx8+LWF/qaCaYN+4ToM5HC149Kaxw6mD
x+WdQsUaRSOl0xyx9pxcZITE6iRDUzFq4yaEXhRKXIzRhGCz5hfNg1W8k6IPacwTaSVvil12i+GA
aNi8WnPTwlbc7RlLZCZq2/R1C31taCAULXDobmL/FP7EPSL0Nc3xUro5RXoLIttTI5VhJQacunud
Ys3gEORJTfJlPNSI+8HZKMlCSqrVxK9Ncqrc/3S9Bqh6kQCpuIt0tUHgqJagaP5T3bETnFvh9OPN
eFoYvVdz9kgQ376WqLBo/3g2k7ziX+ygUspNzo6ICUYG06teT3tgB06H0aJ7nk0aCAK+vNKG1cbz
AQpGArUAxd5+NSgpbioPwbtxbENT0VGrFP5S5n6h7aPZflpJtxLiR1TO51CIvnjKNO+yvd6TRaEq
K9hRCE215N/bEJVioubYTAm6Dk1gwnz9LJAgZr+5q8T8hWVF/+bTP0SU0DtQpfJYSEXxLyis2TQ6
9Cb/7tBT7Z1JEZMP4REDOpGjro8BaJY4gz7L2j3HOy1klRue8PM6ZacWpoo4PW+e7iWlcNIRBHZi
TMnSiU91yRwuxQpkq6BlifGO2yEjzgGxnqhqy9EgmJ2chffafI6LqUSxKetNW+cfWBoywX99ogmF
XRGw/4zrXntlyhXhf49HXT5+xfgvw0ZrCUtoGX4MTC0a7xVTLEVf7NXC1GXAn4uORr/FcGnINrGS
VFunYoBPBoHSR7gBM2flObHkC2apvZoLVJzHs+01h8eEPgM9Q5QWpTp3Ad1rZzCyADN6co7z/5Pz
Xrb71upHfpsssC1SztOQdCDPVuhAtSbD9Rf1H5UlouukafvTCxA5uyL0grI0FVI6IJuNcsPB7Rii
KxngZTnJNqcnD5f5l3cAXwSvLQ2WZ4/7bBE/1Cr01zlbkpcypc3I9vV+FPp4kjTgmDrXmTpLgHn9
iyJdDNkoDfHuUKy2yH5O+MAsK3IRzBZtqTry+eRFACtl+oKIbG2Z5ZRzaF5GTjP3KCinhURPxkIF
JSWK1/j9c3Dx5dPLqgxurzUEDrhuk6Iiod0omvleSb5dUpohLfghJQ7NKvfdogtTopGHjGkJmPFo
Yx917ubINKrtREZyRkcBEgZqmF20PnsMVgBD/fKqFaR1pj1XUYjHIpFgKJzjgQc+O2CS/iukwFwL
8IDPcTpKfzQEkhPAqW1rs81AzPYC+8y+sHycnD3X/q+uofx9nj9QlXS0nxQY2NyykFR/Bgj4Qlpp
19tYGZos9WjsusVa+CgIPmtNd83HIKttKL+AfDtfCBCCI8HDxewgd0DHHjrEDAgLGT1v504HvBXN
cV2mh3nQlGihPo/gSu2Dg0aJ85zZxZRoiCGPWBOircE13tOdi3ou8+alu+Z2d1oG2PYMaBzJkBLD
kry/9r7jjRo/D8CQidL0CCat4o1NyhygO1ifsmELc/MbDrfJCs2dXa52G8QKuMaboq2drGib730P
PgL0jHLZpn/YbLg9tO70Tf0f2MB2B/O6DrLJNTc8naMu3rIc1mu/UzFf1kzNyAEd6gnKjBrmAmQE
E3Jkz9+1MOHqQB5l4TD8iz94LH8qrrjnpBeW3p4wLSEaFe5NSMv3fWh8HNHPkKaF4bsNObg0pvY4
CyXKPqIV+V3ZT7a8RQycpMKm8hEPSXSvmAU6pXFwUNL1JMKJPeMJF2S8CnnUK+VrB/uqUtpRxEK7
0md/CO6lOZBrIZgXCa2Et8clxal53YzJiO63pMHGTvDEI/sMVHUHCTwnVketilylxNCsAYERrtOL
11OFUm7HqaHaz5fu3Mvg/PmTotyuihdk47kvD1uZFJnqzo8dmRru8f5QyJsAZsXDtHwsSHsVQ5kn
+09GlsbOqIsBZKtQkYgI+f+YdF/UDaOgVcWxak0BBfZ3zcKqWlv3gI+rS8/EjnrPZCeiZN59BwMR
XL7uf4T4GZNySxkoKb9HYd7+iSbyzpbab+WsAQfyaj7PW7fexSHP7IqgHfAHlJ4TyYpx/SXd/416
wuwy6j68Zoske/kLvbgawWf1eF8IhIAaBsURY0X829mY1ErpCvbrPznar/xnqcvwqkyuiRus0PkG
o4QkluWXL41yfTVPIqbaDTWZNYuvm/ntxYXQeb/hI2UUcgLuyYeElL3eJH/Ulir2XFq3EaTds9cq
jUnoR/a/Yt6gxmFrr3Uw3Rn3UU1WEnCnTRan1Y3TWiv48zdBZPCFQaoHUE63Yz4bnrnuJCOfHK36
AJiR4+3GIUNDrBw1alyQUewzwPj4f9ulR7+rrfhyS3bdxW35fq4c6Ltuba/j6uCvFiY7W7Q4HkHh
vbxDBxXtWQyGffcERvI0gF8PuP9HjXRJljs0/6dRaVvpmYaFqM9TwqujmtNouItgzTHq6ayUSpKX
ujmPtjPCDq0xzgwSClWTV6P3FP1G/ZQt+OOvX3fRN+ia25kRg8o/6rJ5gyVcFv3MMhTN4PC/YzHN
HLjevWNmP1bXCE/Lod969CdWmRvxHtrHJCtFVbJXokArnIBkUrcz1OV4PV01cT8Jt4kLwy3zfhyg
hqM2VEruZyTe4nazmRVW3ZC+3y6SS61tlna/ntSeBRUqAqXdbLybJsWzarMCl58FhOKg9HFkqzrY
H5xcA0MHk6JSNOLRi8bfPpZCJXnDH6NNjWG3BbJt3uzPtabAMfhRfZrBR0tP6M0yA/MW1e3c4OnJ
+LARtn9gzQC9G2IQhaPxz91nXs3aEqrSAuBODzshXKsuE0Uryua2JwJqUqUqWCbWGb+F8NrS+bFU
8kL8HfbELVQuW3yaDI/p5wXPyZ/IYi2zk/pfA5dr1xmitk+Fh+kdqE63oaUmb2xWrGCQRVVzMKUA
9cYTv30E52fJ8LUMOhuCr0wGyE3fVwL2eY97X9nQ2F3pWmP/uqSl8eAgoIekuj9ZUvhRYHDH0+CF
QfTQNSCEe2LFAr0Fmq/L6a62cvbuHJ+JBesnqw6GOg0ezAVMK4XYApgDQXjV/IU3ylPFa0//nDM3
ij0obW3w74SdB8Z02yk+LbN5G23ViohwEe/7QHl/pvk2PJk5g2nzWyrs30gQAyFrG8WLRkv2nXVJ
FtNryx7bybtSCWOLU7/W2gLj96PtnmxCsRY40/ooLpJdfm7w1CFvCPYRzDYFl+AJd9gdsDxzmjTR
swEhyEioX3yHfkZrlTefoXS57Z+R6aTOJ544Lcoxzp++F7i3ghOtXiQSZ8k8xiMognuDyKnFHwzY
soV2V8GO3diYNb+8kLm5nsRteg/ZW4MCoaJ54X5OvRu1QnuS3+ThBn183FNO7uqXT0YPoGNeNkST
Dndh0zMHIdLYz6PHGQzl2x3LpLZpZE0WycTS4bDONgyZkddPfK/4187XrXYucfCxylGMIYoDMU7E
HnVrQ+1bMlshpBF06hFXeaucmiLmKQdqwv/Bx6TNt05OigzNntkMFIzfkQ03ff6rLSHkX2zIAN2l
2iuMWJy3wJBdt23oxlGv78+WsCEp+EOWTgG5Wj1vX74ZAKMYspJhGARtiqn3qSKBPKDBJlBkvCVD
0z3OhBGq67mIEJ+52u4zbspIXSeELCBus+3cunzSZ70xWw4M6MofqnPyXNKFAr2s5ijVWcWcx805
e0M8pKoG43NfzXlw5nS1lOLrHuCYIxMd6zRv6gb8O2gPYDKPUIvfQCqvCbXnj6qoRzP2XjBxG1FM
PYB2DKnPUc02Mu7W8QXtnCoChkGQP5Hi9YtVjNT8sal9pflTMpGnHOcH1GZvhtOPmKo7dMoQfCcI
WasBbu/OuxbJ04U4I6MfQ1ro8RpMA2p6bsKLE/QHN4nOwQeF/rhDrYYSJCbDIyNlDdTjj4Er3X3H
XvmbDp2e0Qf6XGpxEGU0pEiPXbKVRBJWxklHsqT8U6ud8kGypFf/UjaQuUnwPq+C0j6//Pee/zes
MdU76B5OVS/hUCtRx4nNhgMTm2cLno7lV3YgP1GtL2M7N5JDbv5RIBryRtza1i77Bciz8v4in2Od
Go74341c0uhSNuQXrQXTpeOkPK5l9vMYLXkQE+UFOlNESjGjg9yoQkA278EXmcjaTwvY/2SUzQsw
1K7Nv5Ef5am3/dOCWE7Z3RgOmtjmd6h31CKyawsb1prh3rE/ES3f6TmLQs78aGtT32bRZQxb0ME7
P1bva4iF1BPWF7IvbDyESsST+6mAxROiqGe9ZAoTa1O5l2khqCn/Cpkyga/IWIP5/2h9r/kTgsd8
P2jHgLKwu8eH4t0t/iocZC4GNma/Yq7URce729TjhrXOUCSYobcOfzhHFWpWemGLDxmOeL/alSVP
067itPd+XDkBuu5u/Q4sd2OCYThrPct3pimveFHXYTzv87IIwBtYee1Qe45Vj3q66LqBCNR4If9d
8BAcKeZBRIjx8HK84I6fdtj2T8t/rXM5PBuF1X81dhxLpLlvJUgaTRrp3whsCNwe0f//rtFwhG+C
hM4yQUlZ49U3P3KWpc0Sj6FyCQ5m0Rg+VQ7ysTcz8MCu8FJ8+xduB2htUeyVw4pOgUhKL1QHb/Th
nmuWFgMKs4Go3l76G8RoZqdpcGuudJD7BS3U0JSLRBc21FM9M0V6D1jfEuun2ZjBVq3QrazlEkmL
TIUMHK6RwYnsj6NnvvQp4Esl6HqOgZGc1VYYT0BQ4KDLskSQ2Vc216+icEirgUEFx+xsVZpZc+XT
KcFWS6PLobQP1G2Mc0xde9QYuXV5QWnrhYZitWaLMh4r3n9aFFKiSb2eImKErCSmOR1fm5QgSs/h
A+gnz6FkzkxxWXW1FuM3BoyvYrmKGAW/ZIS/LRByKE6+aM5LcidMf8Xq4YsrP1zbLfAqJSu4/6e4
7FgcoDXm5mx2Aaesxh7BnojnQuMHgbgKbzA1tyD5wT9WGp9Hv8LIrNDGDQjHf9lm078pakgOeSut
fOCJP0C7nDscHoxoJ6dZNmuHTzAyp7/1XIzAbY2AG2/nXsGWMHFEINtyN0jm/Gx+QcnUKONOVWdv
UXxIJVQbYeK65VCbLDn8OIv1KWgJWazzEJ1OKIBOo4vOWMet4iPBcVhNtz1+lmEZuWabsFfJJsSl
CrciU7UKUhF8XZvHXaQlsf1oaaH9PeQyCKXdMrRig7wkfqqNsKQ37R9oXknRy9QLKe3XkVGTZ9B7
Zjh9TLDsfXs2vbZI6q+sFXxsvpHdlJ60/hbVlcfJGxEsvsodpXN8d9K22TjG3EYynX44vTn8eMye
wwzvoRwIY6MSfA7UldTY1fCYYuo8MD9gemQX96utCisaCKMlXOfUQ2qGPorWb8QZdanR26zq40eA
2gW+eTRFPDloIVc6qnIDvZzRwQcWXzjHoebn2hrgbdm8vRXh5X5n25xtU/B1twovmkCEd8y6wIfs
kSMKzjzWMTU2WIdBNpnrfSASkneaS8345P13Nd8icbkAOYNS69iAMZWDCr7YjHrbDyEOIXOkLnkl
x6YK91RQxexSxjjVAIruMgO8L8h4aUcNEFleoJ4yXSujdvnrL25CXozDmfqHGWfclUmxAPQLXI/t
0nLiIDliLlGOGNpl66xmJRJTz/5gon36TlNy/6FGWplTOVS+9wv1jh31IVG3FftI5ZMOhg45hwc1
yRsEoYcUd0Q/ScY+5Vq3C5UYLksU5CkzrfXuHf1RuJt39UvUxt9LCuIdo8+V73FI10BZxnw/k2s6
QFM3if2Fp3i2jpxDtVCFWUMiMlfqu3rreEdXhqeNvQ/uYo/Bv3zErDwvmmCN3HdW9ohCTZkyo9C1
IOrl56Hks0/HGN/DnSv6oaJE5NlYoKMOHTrza7lARTwyY84VVrTPJUs+GBnapIn2MYotIb4J/MSt
hFwPb7cb9/7najU49S//ycXfQwKAaOYRL8lGarDTvS711lYVpZsmZJPi2yWlSNOp6ugt3k3cCLgP
4ziaQUdQUeYgIZWyCNQa3AxlxZ9FXdd4AVEgkWFYjvGtss4OZSoehUkr32OhM/jDoTAi+CBgCKFr
DctuDRhPn7cZ/L4+nVkNL8fGz25lEsiaw5u1PXjA8bJVcdH2KUVCfvwaseKy0b6/JIM5HOxqu9nb
OxNWq2qb0wYu4LTaMZRSyhx6jFUSdRlCk9FgIdXN/5KENA1LcWAmOSw7UEagELYoTL1rZCUMXGZX
/oRnTb79EfRYnqjfvbVjuQXmVphDGp3HsM+ZwKN8etHbv6VFJzZS/4/90egzPPXT74DYPBoG+5ZU
oox1g8nwiGrv3A8cDOLgeRqHvsOZejXpn/8P1X8i0jzvNh3IM066LxrthASAiAVKpfJ8EKHBXPDk
27TBDfmyjacDW0bWCzD+4Gbp+YoiNJetbVnEAcRbeo1nCZOKYAt+eE1/Aey/KKQ9jjABJsKl2YjQ
XcnYYahvN32+ezSoc//J9wKQvkc9vmEZIXWRq3YkeO7YZN1YhTJZS1p1UtOIbLA9+Ey/uygvIjPf
Dmh2u0GpqX0TmDHoRwZpeUUdSUKF4kRouBZfXSTzAiPVuBysXxBPv9+/m5u0sy6Jr0c2y67NwHo9
Qzw5kUxSgYJPxU80HmovW1GLeNS056RENvW7mxp31Pxb+75S5YInNgGpE/8Pp4rlJYQ4kzXal+Xu
6c5E/s09BGPEt/KgdiEc3nJk0kzAlWPCHsUh7q0G+Fl9X9PdrTzKErmgHSVy6xl3CylwXNVkaA3C
Ho3xy77QMxu3GUIVpAqQJ8WZsWzFK3+Q74SXybqN1WyBw2b+g6Zlym83rQkPzxNgcm00D6gxxVwt
u/lpQieGKTiIftWySRoqV+OPWFBAShVTWWHycN4VpX8kr6buzf6TPslNmPSd5z3eLXqAltYxQJi3
aUD/KjkSqTFWJlzyoq7d0qDLRkTAxfgSmLIdHa4nlslhSVn41z47XTJmNQbuIDFRit377PZtKU3g
LFSr7ylP/xCxlIr+q4bKR63rRFIetmZzHnu+e7URGZecVTumhyMudRP7eHfRn6gzOymO9XvazdJT
HIY4WHmddK9f/VGAtFKgosUZg/KKw+4Y6mPSKks5oMswdKCuUNB9kzUvteFcSCNvmiSvOhY62dnz
sfK3oxEpuG61/yR1X4fr6I0gKIE5a/gm8FCxCR0k1g3NVttrDr/iiuuwb/SO8InPkTE8Uh5E/G23
/xp+QlFB5cFJ4e3qcMyF5/ZY8DTg+eaSJKVrcEmg/wdrGGvaDETN1wRLcgu66fpqG1ZgioN6RFCT
nlkXEGTnDNLvIVJs3vjo8lBFmRk5DG4NvCTGkwS/zD3mbNRyVlR3GWcW+yl82EhCihLz4aHC8GSY
LgAGEAQaFx7tEQTy2YxR6a+WGx5mP2z+Dlu7zGye2ZZ16tF3UiCk1NBMt6U3mSSJ80Q9hxW+VzfR
VqMKCtNlGEcrGuS9m+N0CO09tcwWthcwG37q6cfjmuL7Co8/5QAEhpuT7lquqsgiFJjEhGzWlFJ5
GnGJYjFvB+QEbGj5cPT3oAde5bKnuOW15Am3ORnhkKlNDBU0mLVbzZbWEn/mdQFWiNidv3U98yNB
vpbgK++TBHCjhC6bx1yEZ0vPw4Sz4h0Zv8bCUlGaPACvk6EfzAPNjks0nZGuOtV7z/axBQ3pG7zN
A+AWDSJOwVF+GhaFoezT8+E730R+B9C/BX3r540OXigRnMgwE1KPYJuFWriQIVfEVlTEcRicHqYz
2kJ1ptvWMhtRChzHpIJP7vlvP4r/OPOjM4TeCkPsvKjDcpUTWdV9qiremCRbI5Rp+DYLvG0cZIHQ
huOneNY8jgiKrI7UcDdEOE/OBt5xtXuMPfsllSKCSMYCnupGIOx0LzqUPL8bqiqra7PKHXzEcSBC
kyOOvC+tFU06m6BM7OsGprxupHXfgVhZR3mOEI4lPhpallLAQX8vk0Jg001y1pPVZcqC1LDFSJ/e
XxaLRan1iTu4UOSPQcBZzGOvhoPMhCdHJ3DvIjqCWcFGfNG0VpfbpjthIWOZOA9vAHhlpxYJ3MRv
W7Mm4V2lyycqlLuUTcU0l/pzc2q4CZa7g+JCgJw/GGhjSKyVfUB3ZNaWambxgqkRK/YapYKVENpk
C+4r4sbOOgOxw6rptUGJGWX9A2RLENhWmqu1NKkWNbSnWxuVyo2oloxGXKa3X+QaVgmxofq1GD0N
mPmXqgLhxi/4AETZ64t7YMoyXkOb9QaBFs08IXkFUf4B/dBQ278QIr1MTvohZEl5ucJHCi9Czjk1
0d2CrIW7ZPLDJADOUMM1byrFtVaSsQjMuzpJg1fP4ubPqh2COXGvZWGIK2pXoLVTWSQX73dXKgvM
ClerWD4FG8pSh0FEl7naf90N87XtdFJ7/32h/8rF6jWfmeAexfgber6xS3waxhyrPe8aVmEcKiWN
H9O812+oILjf4prwJutJIPadqSsVKWvSbhym9rBB+hYZwEv3HF8avjl3FoHOvK/nEn4hi5NPeheo
kDPsUW+POFTGbfU0FUk7jRMFEr5ZSD+FN917+S6VIANl7rYnRZSxcqG3Dy5l0U2dnZA2oEr1gcId
vOsq78TQ1eAmAGQk3D9CJVdKYYZ5wQKy3EGpp9VO5LHc0GJ3RHK2c6LUToafKuXD9ELryWFs+pf+
dKZp2jlC3dbAuvOFlqi2ttcSw6S5/u/FJegt/rO8OWSjsRGUNNa+IROr9CSfRtenGK1f5tlGX4W4
RCKeY+aTtX4Volz5cIjqeiH59vPBQh0Ancd2c8OPCs3E1mrvNphUI3JflmEnuMvR7+wyfTZTzAAM
q/r+91s8FY/h1aSzWRFjMS4R2E7Fycig4vs2BKQHrGqZdQd1ImqJeWAAZFgYX0yQiOaepR3m4Mo9
dD73fLXAH13D1rpLIOr5GcI98KHqiS9pAiOB7T48BqjVi6SWsvcEerpdp7I2/ZzEb2gFoKUxqNby
7Qsnl+UqSSycGdnft7gV07E+yTXk3tU591AnJmH6ZWrz7OV8b/oVNPdYsd1NyZWwdx3NViI952ah
bdsEZDkp6yj5IzV7UF3DsIkY6yw+BFKE8bzNSytUr8KvceEnAXpD4beih/BijajkZomMPue+N24V
TZhOsSVFXg42E/mgV7SJZ4GLQiF4vIepLL//TkmOaHq7N40LsjW66ba3fUaoI3lul8IJIuGLXvaA
YgW+gqkUDVPXJoJ7fe1JxCt9BNAZbT7XRfFtqhX0eDChe6ahABvXkOcdXtaK9f095vH8Fctyc9u5
nOt22R+woMLRiDER+jRYr8mzVolliIrBBhQI2reToMofMkGRdlOX64XVKciebm824GVaocXCXmPp
WG9jh90DyZff6VmXH7X7upoVQRKrsm0tnd3R/2IWdejLhhKvSq3a9t8qiIvMh3b+MuvtICBO77cb
IGmZlQ8ZsIIFQPq/YTmQMc8dat45e7wn+asty92n402o2u2hfE25q7Op80vuWjG+vUsbqhmLyQrF
1lXelgMRCGosyj8LzPkxJMlaJ3uV++49eESsNXGk32MCoxnTv7yIwJfjJ8soZHrRDknunDT+MKVl
svbktFUKYyOLnOX7YiHpjtMecsqibqTThwykDumz43TlmejM4pnqP/PXhNoMT35FYPleqg7+b/Rd
eqfa8oMOq4RjH0gURJ5PPl0PIcPZ5fEUKVYukKS2xl5MxEh4e03lraZHtK9aq2k3PaGaRIqcmF1g
9Gcb6iSP54JeHucJZLTDvFGM2pyRBIZIMdGmFktDlOWN4JJUw8HFTa2z1HReNV9tbc5xTu9WorGQ
YPxCsUieJKKW/okDL9kjjln5WDA3FI+vl3U2Qz1+Iq+AlIZJ3w56LNEXlF0o9F2Vcia2fIdvGjhO
RJmUd0rxol7NthrIXDSHUUe2Lgsp1HTq3z0hH3EzCAKvxABRpLYWRQetDf921Bm9h3QinJXvMMSX
JePtuYP6tolzqQG7FZ0JkHqPNeqBTejyrVQJbpwdGoVWnnOD+cAtXukUt04bzOz2bTEjnf6tGAxY
tNWuTEcGm8tTzlbN0yLCm/yUnGNQRPEDA+r6hSgWl6GLgO0MGcpSXpaXYaPm6b7YKoWo8Wu4xs/S
j11RlFaMaksLnhia0yjPVvbGUu54+zr9/ENPY98unfTpJrZJdP/xxlmpzmHuphPG6228Y/MiCUcO
bgKETZ/HW/hjW1Z32injF4YvmdhTQ2kg2FQ5/MgUxGu1xmo2jbQcGy+opucUivSXwjK3GawCpVRa
0T+z9prNwMlbpHM0CEJ78AP/Ei8HhJ7s0OWgky2zEqtg5y7lWF0qL4UbfnxaoeygcPxioSJdwFeA
xykM4dmgFTvqIPhf46zVqY1/NLjfP89wnbakj9uK13fWGYh4LLmdA+0U9G7hCcFzIsWhiimrQHg+
OUDiuz/+CsDbsG6Bs9JTQpNYNM5iZXk5hcC0MqNgwm5o4Hqk8r66Um4lUjWyNoqAF+8IJiJF16Xt
U1vVnS//ChlA7ysDpLOdIT7FKQ3hs08FrsbQsA7xbnciP3TfDvLay2gq/qhMJzGu0rKZNMNVd5um
5JFtFarT/92fnAtNgRk0qzTn6W07Im3p7qcs6IxKE3Ar3dOUkgroJ5cg1IYhLEHfgmdh9EU/arx6
g0MNCVL4M/mhd8bnJzRYhzKpPtVHFbC6nf9qg+SvhpaRXzk/LIilyP8dg1i9kFVXIL3U1b6IsmVD
13aSXPc9TPNqL1sCrrvs9KwbGWuP78HGg3rqTLziVznekFkp5lgKOWsJtTvkfPmZvBd8RbXF9fxo
Pk4wBEjHX1MHuqdnGn2r7rhjVkbexNgBoy8sugrAL/cp4HPGUs/F40kW78vpWhqCNL1wWcyWDh4c
2ZhfAS0YygiQP16oCx423qyR5F3JaVhqfdVGLh1GffbOkB4xROC+LO92ereQWfTSBiPVOGjUpj30
BIoX1no9q4C7tUrj6K0CK5oH+gxD0QMgkqEbV5yirDnGpvPHuU4Cs3zJMOvzRzP1UXVJUcvD6VIm
Buv4fpHmVCaZuhcEGZMl7sSF8lDMj67wmMJEDL7UxqBTh11XeyLmX/3F61Lh5388ZoCxtnYZu81k
h+kCd74fPAesob4U0TSp5HNst7EDDDq/G3OzXfjxbjLMQS+X+pH5/ICs/eHTkp8hYaNTn0gcFXaB
h4PkQqd3nFu3WPnIsedhZmRVR6jQAQuocMtmbUUMLvow3v2OiUDQrg5ZE2sBdOiYj+O9FzdOw9aM
kbyeaEvMbBn+DScYIoRG+yJtjvRXs5q4w5nr+t8R+aoK+HAjkeYys2/t18y2FbukVweDtoroWOTU
IXkowoxpX9DaEntLjMNhxZpnCBTWjmJRoHMYeg0OQH8+TlzSaGE1dtmx7kOwin2842fjS//C5aiN
MV2FHR0fYXxSYpClWzsARv4YUvjGxpgO+TIgUNuZoq7k9koIHf3I4a3EtR2LJ+0ArPf88m6T/iEu
xMM4gHOUDn5diRtaEipqzXgDHq9TrvupKvQGphixWAZonrzc6/q1QbjVpuxXB0LlTui+4evyHMsV
b8nJGJMbpqa4wIKYChc+gpFncTjgVoH7R36s2XmhdIawsaM+hzsIRVMdMIhDof1kShaO9twDO3Zc
+IBQyu1pSJmhbAp6tMtFtdTQDWDHH9FW4DTb4dcE472hYiUGeA/7RVdu+78/YH0PrHNNAef+dA+n
DiGGjfJ7d0x7DiHXlQwkxqa4hHXBn3X+Ig28zubV0LtLgkc1dgKp9KjEQhdwFn3b3Nkx+3HtYwkV
xoU2XoN5XUbC+jaH/fhokBQ1p44SY40MojMBJt9YsLZLV5ttADIvQA8kvWKsGS5Yi7uMNhFhPR9i
5Hl093SRicXXaiOxxlnLWXls8JKpjhI+lJHOGiERaCefbv056iFC5AA57/e/5RAVJLpBk2KR6XBR
9AsZbCmlXSDoMDJNigVRUKhNrLn/2zcEsYm1s7z8gaeq1GbFe9kQm4ybWf5TJnxqnv0L3dmvovqs
JAJNbf+3bfgU3FWO+43jdfQqonP6z0Y2wz8eMIyfWK52V0p7sXtM9NzyrZmY355z85OxQKtDeX6i
+1JSiNShQ7QWnpLrdlZPtJHttlT78q3pcYYQ5o9lKG30N6IH4H2VXN6Dufqei/s6303JDLzCbgLc
n5nAfdiZIMUMyijKHa7DMy50Dp9g1UgE1YI+o9VUDlVxF4PvvN5ykWaEVn7shML+5MnWC3yaZijh
rqs/GVJMT8Ec/WpauBa8moFXXktyJizWRYlrdq7PgJLICa3pNi0qQvm/XJfaxGqLg8tXTnpElNKu
/zf+M0yt6NHoxSq1SB0FfXSde2R6EqIUJXJrDZRqqMlw80zG7PlM/WMe+VVGACOsfzgQTsbfBLix
I1A8geLcYOTnJBCH/wkWiNWTCu2IQXBQ/RNlGaffbX1gpyw4GA3cKmf6/AuboNCKVj2IN4n7OjJW
oz+2qi5ae42fyXH0b61smDUwFWu5b/apa9mUofEz/rvPZyyn1bf/l2M+foJqmxweOlk1C/hxaHSs
RJ5woLhKVHUxZMoC+e7iLlju45Wi6tAoW2rrMzOvk6QvimDZohyZsu2wmAYC0XPwJ3VZKHAkTffD
6Vaw4sih7/eD3Ck1TNfRZIj0/Vzci6Ru1qiCqU7eaOYl3mtVFhQgAL9xRDMN4XgcjQJO98DSCchc
g2RvV7SWMDm23Admi0JoIzKsZSMg4ftNU/Jjyn0GSv5COvwMbGyN1TypIWOAw+Yfkc9TBLov5Xnl
0zFwBZfdWzEUFI9j3BOLPh4mjcN3nKxSAZuXky51uyzPBjlV3t29MjpyBFxqidoD6DVM3gpdsA/q
RPAtDmUVVgpBpf4w9dkzdDZjxuktJRnM/LX1rf1S73aZLjfYmm4GQGWam1L1nIlNvHVfzeWRhLb7
wgsk7m5hAXWVmByeirPrpX73D/W4/s4FUd3hPbCxHAVd5937cWd6bWMMmy2QZqEAYp3b2ZKm3soK
GlgH0aZoQB2d2xZlps2XRqKT9cDCcBsarzcdPdXrMJk9CyuLQxclcJ5XYC/ghsjrd52oD1DVV8uT
Q2fkyR09zrKHdQsHQz40lAaT56svAUuoXPmLHzHA6M07BWzFPyRNJSU5YCn3Qx017u3wezZME2C7
aQuMLy1Dj7z2xUMtF5ezJe00Cd3L/pWwW21wiUMkSPnG47CjPOmBM2dxxNIhyjtOba0tr7ssBdc1
h+n+WPD2EmtwLG+oMKUcvH/Pbx7UHhichppdH7RV2lHOrNGA/D9IJVgRQ0cY8i+Jvtdxcn42NBJ1
RC5gaI6B2bVkuVB8qziGbjxCa/XhMhBH4wBItvDP8qGgX25XFgMS6tMPLswLIUwyyF6FdQyGcDf7
qogIDgQ1Owwt+lEfEJ5cKZUXB/XbotmDoqZp0KRLQnMi8xgpXfqZXv1usny8nRrit3qt+W7HieGb
UfgjOb1fFmUoLsS52IqTYX8HOvkHfeXYrdlDrmFt5KlThcUwBdMlL1O+hiRPJHXZhUeYVffqbQ9O
V9jccWt6bX9AJAZbrhO2d7jgjBwpkguHArEljiBPUzA39JReCwcuKnrh6mUOVNEgv28qI2AepTRQ
igdrAi5BDYGiOGccfsqTOZvqmBc1oXvjiOjC8DH0bxu5iIkba1MdmzGTIezNo98PwkFt08moX01c
zQQD9R/GcEjDUrE0jq7s43x3VyzNzQ94zMd4lyqg7mkWxM92BCM7Ct8ppb4qu3SjpuPHweuWU4Jb
11W+hGPgZ0QamyDmQFGrEB43US53Rqug5SjrFx543whve6i5KmGw4tICqDz9HSsPgdcM3nSAVVRq
9nkpWVdag3xkkNcMgMSPOZZWyVaY+IHSxpjz2RClMSQA4wXCWaDxqnNq2sirJrqiuShqWFRp+LQ/
t377gtE/AhJ6q5cTAt1gSJvJbcvsbv6i1c/wOwGU4HDA+rsQmjs4Ut6f1mhorsCpLT5BoD3RG5L2
A3urVISU5wI7H1XFlBTV1rz6n8kOwzLYlqWslGxLOPbUHppe5OPREWj0I/ayMquJiL8vM2ArPosc
iyWJju8Yu2Y6uTG44oB3Xf+vPWUPOt2XybJp16PRk50uKRW8xSmXxQbk2IRhU4aVmZoei+eL1xU/
eAO5fV54zjWRuSjoOegw3joIxrk+9sw8JIbdA3uyrtfdW7JBwSX9TNLvHpqKoy50jEIQpThqJeh/
561eEBS6njJXZMCU14YC2Cx0IgNlCmcICOI4oEIIFiUlT5HBQ0kcly37y6atiZBmSneKAI4PnYp/
Pqp+p0nNBz2N0DNrTK+/lF7xzkSHrzaH4XQ63AV70d4eTwOQCodum1Ti5OQkOuLxui17H5QntkOh
C/ySwajUpICXhqEMX7bZs+W99bzTr90m6OzxsfIrlBlAC6YghUOS5vujPfYpPGfViPRxVv9LvFsN
fkYIbEcqME82/usGqaK8Dqb+cNrJT8KfpXihbYyY6R87/JdNUqL5xcG4nmrRzCEMjrNrV2Nwd8wY
Pv/2Mo/0fTf3uG4M7lTqSzhJHvWzEfqijrVwR9BJr9Ee0bZJl7oGf9H8Kh249jI84IXvvDnkZTVI
LeT4fOeeOYhoCoSfD6NNnMysvfSWg/I/VSt5Ge5xbnnaFCVNV4vBcQZ8jVSSRKeuyoAbDXXMgh2f
YNi2zhzJWWJ/corXuEfM9jFRtd17UsHo2wDz4JOJUTv9DwcGGiWsKS/yKKFydgicghNLEvuX5Vwo
gMe0TTMYe8YEU9vZn/+GOA/bgJTa5I/d8xQ1TH8HXIcPBOgQCgNuLhfLUap4Qy4Jacezq1R5CTv/
+D7OItYC1m28lbGEsEH/sC9LIk+p1wy3ti1J6+11dAqFvNrdLip84HuLpoIo5BzL4A5vuooZ7nh4
XIysvnTHHhKiWJHJAVXJj7ZNJ8K+tU49dGdLv4a73arATl7w4eewp8m4Q6/4NLdeh/BLDmEemgxq
RJuT69mukKjSZok10OvVf+5BK3qpcSXpQIUwLqYzhpqfNBzYGH2dbZMiOhJ/UOLgPJu0fW3VnSR6
Zzwvh74lVx0x83h5GWJSRenKcofWZmlCTU4AO52mCMYcpvugDubWkAbCNmIGifTl0rw0JuuIrVwo
69OdLSKv4rSqa1j7I6DlQD3WQJg6YJolHkzsCMqn/zi5XWOevK1w7Ir9wCZs8lmUpU3ELg0nd7u3
EZNleY0O9L0NU8WaKw1hGVCoMqxReu9AGBxpOrpy3l6Vf5/KTGsoPYIYK9m6yv/XWpRd+bOEO9/g
JXg/lztP5iW+cB2mth+P1FhYWZ9W9v76dwXhFSkkwtQz5wgUwjmXX4QGqi+SQb0ycu5XE2I9LfTA
qvvSf9ePvl0FRzDpQDbFLF3nHs2Yyy5cM0mJXQDr8N6cijgTwZTD1/wXoBuwtRP57tFxbG+/99md
F7PVlVp+7I4rjbLbxjJgegzS2U7I7c3y0DuyN97lmwNBNSIjXbskAiOHHWdQYt+qPICLrxOUaDr5
aIyMIwIRg/tjLCldHZxYhK+NTaHKzWt8QjvTkmg8e18Gss6G3oUFnqzZv3/Ln5z5snfPtyMnP2t0
VdMntWCkXBwtArUovhLNGKNX5CJBmI/AzL4SqemLhqiMJbEK2UpwwsxX1cW8gsZDamseGTbhW951
IjZ8agMUEWOqWjQZxpqPwEmmAdGosegwhVJHDmVvg8ksLKVuudH5jwPrhApEwVjaOm+mAxWrzXiK
fN4e5xVlu7qowW8QJq0bt7TTXsmi/RG70p/O9DOOHrbN+2ZM1cXOwOa2qnowfUigy0XYDb3v8UjD
AmoVSPXAniqv95sDti/VSsWdDclKBWXjNIr0Tx1k8l5fXnlLB2RvI1GRUV0yr6PvJY2DtCIhUC4y
rSBZAMIkuCZsLmJOUjOXqugkHrTnqHXWbD4qoLJJXUckAt0DnTT3QcNWv4VCv/Cx46nNJJFxYaw+
t7CMz+2MpcSwc1EbG3hWXA5h4LOd4oQRQYtdfkJ+Rd+9Ka9kwfMlO24TA5OZerGCwnlOQ0Q4eHO/
X32x3jq0tpMtKFZz8yVMm+Qj3eRrtxpVLeGqgpX0dS5LAl0R63VkW2MhMSIzo+ylwEyg3AGHxIcb
QZMW55DTYBN8Nqvj1zAchVWZsnwix90wEh6Bd0cjMdcapFsgQjnLkui62U91V4YJZSQ+ay5I3n6h
euD/CTFXXs/+gdsVtq9UNsfQYkvGOx0pdQLAJK3HS3i2La4MntLdjEFZIu/Ny5yd6vgMEzVsMi13
C9gYJNt3C0Ov3BXcPge2ofI7FtyG60qa/TawxF9w7guYWlhHdc6Jupp1oBxpOu48JCvMboT0qeNK
TL9gK5sZM/XL8YRUkP8FjvUzWt8REJcMjSgGNrjmcv23y0PoAExYDAXMn8fHNJZ2BGCvAps8quJg
gDuDgm8mzjbVqtW0TUirD8LKJzeIR0yf9miBFeHj/wJWNYsc+F4i4KeEcIDY2uaVGx/4uQO95QCh
WtNFzQLVJQ+hliHZBhNp7aNlP7+u/Cnu0GodE68qsw6k8ndPRtnNkD0yoZDHGA789jxSH1YByxMQ
fEmyG381vwgrzzrIYDUcNwDOoDsuIbi1kzi0jdtAAkHCRaj0h9tJHtHKr1zCFZCuotFkVkFxNlzD
2y50zo+oTr6TVQCUUtjAlZqN5BdrqGg1nXzYmB6PZgV8N8POD7s3/JXFM9xPvQ7NznvS+u3Hyt54
5HdBZqIrTyvITAAny8bXT0dknvqbNMfzDD9LDHdM1/oCxSz0LP3kRKR5DJpGpOVnxItU9syqPdVZ
45ETeQPzXHrVDgejoNKRdGCwOktVrCx6Ys3/bSB/19u0/tcssM9tf2PigBMw07VYcp8RsEyeZ/JZ
MpFNwkq2TOodicE6dog0ezJ13/d22Dp3WXBjDrwsni4Mj8SawKKNOO21PfRJyZ8NyTjMkrZyze7+
XebBSeJQ5qwo9eGQ2vxcnKd/Hwc+uPCxsbzhofElyRdb6tZYKOstt2YbQTdqwZSLfoSW1Q1+jXRt
IhDG6DliFJZqcukXDsnc8JYb8029nEme2BiOxrUMuTkwbUW2lbrbHfHV/oBH/7wV5HTNfhbrytgn
FZV+EDH/pWmyp4TQbDFX+ewKWsFGtBL7J1h0O9Oj+7kt79G4/vTQmOBuhjLBNyN2cY+MtuUt0lT1
36b9/Mmvg7fEiaOCrYinsh7OjucC0pnQzq7mLEugv4riiKV3NH5R+hEHEnR5zLp5NU+EmckD2atl
aWHDRw7tSPoLvaKG7iNLfMT0+Xn+FQjb12Q+Q+9i42as4MQhqsORtMtS0YRM2wfF3IAp/eGQGo2F
s7g6TES8Jeb4LCsrxKB3g5UxALQYYyh1Q3ojglbAcfknwhhxHAhhM/dgx/9NR/bEfytwaAehhdiv
tiuXU+3f/MWV5bKr0k2qzMFzDy2Kek61s9usUq0p0Z8FBTvWZMDSE0VqV72CpAtZKk2C9QxN2Oj1
hVvaKT6U3ClVKz9YO72B94Th+Pg81Is2ZkpBG0/m2AaYlja9eDuDurbscJYAZNnSvuSODx0/AMT7
NyZokJOxt8IwpJ+N0ZZftdCuCbeRphk2aJjlHI5WcqhBl9sYOPoM841a6fkdlacaxpotyuFCJzQc
RTbsMofRH41JbL3R0CcJe+LopbbcIDwRdpxVQ1+vOOldqmyczl69MbdkHAtm/KXwGGlxSnMw1/aU
IZdBA67+j64FezIpOYaD3jpDX41tIGy8gySPURyRMEzvZtPPiLsd9TK2W1MpegeARJRMX1QZhUQK
QqhjSzrAbSJ/+dsr57+lQ9NEVtaEyoMF9ubNM2CjoR+sHHKwlg+6ClcqBMXDcfPzS2WKMKzp1Ohk
eHbyq8UaNV2fxDDBtmsyV3UIsFCw/m5nMCOsoko5UdKeDIgb5zUj9JucG4pHychliwouMrFVTa2T
QDqE8HG5WOH1TA8Peb8NeS10vt7NztAI4r4bZsHoWEjKbelPF3XQ7XhVKSOFo60sOG1FfEnntzBl
gxSh6vph8RsOkhylkmxyDuoGdqeVRq7oSTb4npf4/FO1DTUqlDz+NqATygZf2vFCEQS4uqLEHFcZ
UUf+3Eq9OtY07rt2DCQrYjh1R0n9f6jmJZlRnS5Zj5JYo2nBis2N3fHSlmxrN5tHnl7GdDrIXXA9
jR+DnLDYkT4p4g+i6ocaReyMrTmpqqIc5p86gjSSd6iNsaanEZulZMaFEa37OtMkYfxJIvFBFIwX
8ZkrZXBqsfrDXjsYM/SSjd2ncJeP0Wp5YcCVSAtYxTpHHiEXS7zhDovcybBwrRbs7di7NdzKTNot
HN8VAlCnm1jGH+fP7Ht/ioJT397xzBgwCeB5BkCM9P3x3FZ0TNwK1eMOg+mYsk7DijT/ZEUQ3FQB
ZfpDOoae8lDcyPKHq3P7DnpO3No3+z6PJCqutxY6rz82Z2/Vk2t8AzoyE8EXcedEIuKJPjZD6+eb
XVGDVpMNFJyKxzHu7oFQhAwS2+zc4j7sFBHoUsBSCBWSZQ5QMDjgbKJb7bQVUmTveJeaBs6D53zh
y5LMkc4IGP36hdpotKPH9gRXnZuuqTKz+RUTddPAZ0+PlNWmafLqh2yn0cIQwgVrZElTg4T6z6TR
PPZt+sB6IZxHu7iowVRn2BVou+WE0XXLDZZgLFYt/bQEMVxF7K6ykgEZNmwcOHpBXmJvCAcnZMJR
L0shGXjIrNx/FvJYS9K1hel7p9iFJ8nB/81COgu6BpToiFtvbW7Zy4Ke/KGi+QUnrpP8HzI7e6f9
+/VJbIuFTQXdqX6AZmUlVTntDqOJFjm+D9SzcbgkBLld/YtE5+AbYYjJ+RK2NHbEftMofGWziy+K
0se+beKKfntmWh/NWEBmsDDfwEKr+VUhl9FaHf0eniJoLidtt1AU+rdgyPmXm3g6kzE1crkm4z9V
XTmnCaC9im1wzKTu16f9BGfrNhHTbB2sTEmgFw0oi3lwUlfRkOHGVBoUfdhy/a2KjRTF95VkwYUD
ljXvJaowia+1rdZ8t/HQbO7lnln3Ad6cuyVjvKFJmY5cZrgzppWqktqVybChBIjpzjzy3NlgoFMx
sJvsSDcTYi/MCSG88qmAYdbAeYbB4NivK03t33NndB5SvUPItFTCdx8SBWFmXpmRXxRCOzzzd7Nd
kgT5YQccCS6/jEMIMVBBR3aEwMkQdhOx0L9cDDhwTuvF6iwLO9DkdDq9g/MjDsKfl4hvYd45u3el
vMkhgAOhXR96AsMzhNZAhzgek7Qv8ixOSPr8NzlS2KYY0xt8eYBROqXy0dMnBAW+FFaiBgC43u6z
AGWjYTckKIwUigo98vFPM0o/nc7+AH7W4CQNJjHnNTyNjdDf/RCGFafu35ayzkZ9mqYKW3GkoBuS
p9s5egwMAsLF1xFPSlAZ4yCsixQ/T5LdwvedB4FCX68+wiXBfzB8krmtJkj92/McvOB8kBrSrlH7
Kem3IaS3o+UcPL9TQd0zsOP3FoCAslUYAHFk55zNZ2KqsCb1C5k/eOA15Gfkh11QzAD2HIjgEQQ9
tl1fV9ETTYCbwJvKFOOOBnf8ie4SbU3oXdmhZnEGPB5Lw3YBh+QJW1M0nJQZwOs3JBPyxE3q2+FC
j9qQr6cEfYB++DEbiksWhDWO5++IOAGPcu92pa1QG7/V71+Bnjm2dnPuvXml2LGUaICaiZrb0uVi
6drD2pqg1uG9WblEqeNJgXuYhuJyg7z5/T/5vxutUkPITJi1V1cEPtlBxUHl5CXDqVlvtNXkU8O6
VYH3q1NbchKrt5qVpd3OGjX/hwiP9Aaci9yMMSWU3vrQqV/EgFQWSe8tNpANoYMBOJp5h2qWk2+P
oOPBzPtJ6JN6j1sJDVpClayCPeg4Ohh2ejcFpwbxoJ7VmQ8pAuCY4VbUpjOS9HnigDFnODl7cfPm
KtHJyJCNVyUWlI/Okqe4mlFE6TVakGcT5cR6U3TAonQvJDnL+bopVFNf+sbjea5TdC2DK+Qx66LI
HHFsjWvm9jSsGJAFdzWloONA3UCytZMKm8BQcomeJQIV0N8EzmrlxdWrMEYy12uOWvHyjALb9+lA
LFu4WBuLGGGk+zGD9Xx9G875yqZ5tgTVpPltBYsi3hQ33s78ppVcaXDlVugY/ux8dGPLv6kCpql2
lZtXqWJcAbe/ObU0GVTfPZt435z8MxCRNjQtRc6gq7iSEvxObZ3ik6Id8AwzBTjojA7GtOTzfoIB
fgj8Nx8igfAhD2p4bq/KoD1P9ENhdYIY3gllAerWjH+hHubWZZ693XUTlAPcGJrxDY5SbtJ+6PXj
bdFTHozZHIHwJZhlahZEtmuN3kOug4qWt/F2DAYhP1z/QtdqD9oRir2uSlcjfHK6JHvvp6ctmuxi
rP2CtsAwgZ0kg/pM6xf8/dSyL/BjnMU9BlcX0Y1PzOXF8J1X5vrz2bZh7SYWzGQzjwkeAragpi8Q
3cqU00qqKt5IIe10F9tKxJAdFIeLKeFTFjRjVxxxiXCruyehQYRc+uXMcRIi3c7mKm2G94v0twkg
+ebvo5iaqY0dcHik712FAiEwvMuOfEaYvrdzZnIPZvvi7bT4R/zQPTM3fmxsEVQb9PQ6dUrJqItv
i1RMQich/R5Zp8xo81xqQ21q9a9Xvf5m7Kf5X1x03713tlmahS5CJTPnL0wCS2EvxZPiGHUTR/bU
oCLT20sgO0kTMKGKtuF3bkF5E8nCxKJW5piFuMZGzBlnuNK78+sb1uPXWRUxoj0EFjudvwTln7mH
gs4ycjUu/a4owEb7gP5TqjXza/DZTC8ZPUJIC11/BwLyviXj4G5QSpq5ed9UK9tUHeZ35+KP8MEN
AYQO/I21xnsD9ItzHjWeGtmxGpTlNsB5XvmfVCMvY4Z1n1hj6WrwNLl74zFXA+eJtUR6+5V99dqL
EJmpgNEZ/aZQ3iHMzw0r0FFTrpN1OAfMuhaHFCCCq3tX09XgaIAj3EmJi4jOQQlRgEEwTvE4mbw+
v2ejzv1JDmwJmKjBkMYO7cjtCp0FzJh1aBwDZx8ktzy4ZBu0tSKXVkZ5rBrwr7IYU0lOVJCMQcqI
q00bxmXjDvosKjQ3QBmSMZyLKpi996mj2vluNo61SqvzPt23ITyUuFvKDpXZvCcR2xSr2Y03nkyJ
VCQfqHCoX7mMDa5iDzzvv1ArrUH5Yr7zLz7X+XmUPeZFAzL5hUmDmvuZtEHJkq2x4zIZTcZS+lDx
wFH1neC/25pca+/GQPIlwMwIsfUNrQ7xF7N1MJbjrwmdc6cOaL75JZr9wVkzugn7+nkJ6DbjYS59
xc1qsFlq07JCM7vqkqIIqUqV5YFy+X0zdbp5RgrHq7ybT3KLTxh2VrDeiyHsMb/XnOwzOlw68KYC
yrvtnuEapAkz5zj8omlJgt0zJRmD95cqF8vLseltcukTbrfPZ/rwgeULCN5YXYE+w0nxRj2REbp5
LL39z36+6f4hGpp0Z5zKT19376fNCQtgEbQYvoe/R9AZ90OBkJUi3aM82VmmySK8R6XeDHBkn00L
25jfbngWzrDOKuuaKsssXpYzCjnTo8nSMeRIIklw43QaN8xOB5kJWpzMwLaZ526HbraD9LkPOpNN
ubpy8fJkoNd2myieNBR+IPOJOuJPW7syf+A/GWXOD5OPIwYpqLmXip2kUpQzrBZkaNq2TS+JEUJf
LVgyygUfmKSqsmjQ/JtMFpaPGvSPLjT+qSdQu8kvATr9bhf8U94tJl5cQD1LkVN9a7eL5RXOU2/t
ARS46x/nzKGBq1AFfv7TCHtdnz8Yl4jCDCVnl0ILSoX7UFg7iVCtD3NHDU8Ij/04vgluw2PE5XAH
rneJAGT6mU/0WZIofzalinpGeaW49wt4+ZSEFOjLylBY5VZsJDmzeIksQeW/67V6jDfn6XM5tDH+
zPo3ybJLl7aEtTHihA6OFFXIRzHtLo4bNaZSx3zorXgQDHtaB5RlM4KyZe+dPPpQNiB+Oxk1YaP8
qrXkKcgDPJZr/JYVI9RSo6yI62YyMIHUXXK0D0H+mBhTN0eTREOmSEQalq6Y80mBOh/B4brVKuMa
UrvMo3GWp5iDV+bHfrmnQGzQXPWctofB+zEfmAGOCfSVa4APmhrmRwLp57CC2iAPAitnkDlRamQu
gZMJ9hBWE7c5iqDi3SrXJzBvVu0symsZVUAQQVNC5CeArrOpPACzrCXtv40Vd5KX4IuxPTKW9TWI
Nx46b5ixGQlh/wGy9uvzs6MeQX7pxwkJXPVikLzJJLJY+aaE585RvEwdot2/05NZ8DkZzg15iuuf
o2N6EeC4txcAb1VFE3WiH7kNHFpTAQkLIE+pOg/CJJkoMs+rs1Q+0fnHJVpQtPoehy37hIzcLoaC
A6/3OIymbZhRu5bUkVRYhqAJcQRHmsRFqDYY1QQGQoh3nnVye3QOYu+FHHORAgqxhRyXObO8O/sO
KpTa21iU5aSzpYEmQgKpUqMFj74V8aYor9drWIoSPeKU6lZLatwEBBodK2eF1IpZX1TBZIBBtZr8
d4nCETSVGc6C99FOxtdargIsLZpvqb4L9DCuwKN0+aem2A45CmxqGoMyvSsvAGd7uHPo8TZ+eX6A
mmk9fu8T66Q/osqzjmpM5siv7WGkCPduxwr5PMCODFeq8oW8FJHftpsR312LJDcwFFKEZVBJ6gyP
O5y+vnVTtzOBFZmhPgs6Ux1BPZ3q01rGo81hNKm76bLKFyJZx3dSQsdVEUkn5U5rVn6Fh60e188R
97kZ9BhNbSIrVEuq94ZdQ/6u7nnFBrW4xqHgriCPp4KjdeCtWnR7ZSJOhORjzPKQOikoMCTQ9WnC
IcFb9xP2pCxgpMUKjQ5d/4mCVOTmnAvWY19Te90Y0pEo8GdtcdPvREgmztapQNt/dfHDM/HQhA8s
Q0RBt7eIzgq3d6m+GekYkxQRSBleBgEqLtJSMQV+7NTLjQPE/g4cqcfmgvKPsznTUTOPyjZON1IP
YCDA47A3TTes6oQ63FOFWfWLbJ9ew345uR005mqDrMUd9N4OQoZBzQ8p6apwsipgcCx/YbSsG+pz
Jocoet7A39CF3YV967dJqNzTWVklgGgBMO/Cg9woirhIvVV6q9IXC0sAVawUre54JHOBp68WIKR5
mNra6JldPk/BMVz1mkAclGb6iB142My7vX7Nvoo7KYRQLON5zkOaHpC+LEH1NIcSpHIckmagKqIj
Otced5P9sK4uXaU6BDkmy9R2+SXT0FXxDFgfzUINiYEK7Cr1xL4XoewTbQHCYLi5BJQaoToxGc2M
TPSrhWfgwrUcmseBVPU/vrZfBPUcU+4Vn2Q82JCNgZhHfUehZUnUn2ncARLQxQu+3BHgFuQRMD9X
w0Zfytv/bis3u5psrmXDjDXKua4EEP3P4Mfp2lMOsd3mAC5ZEJszZjRR2Mu4YskvqlUUeq7iIUC0
G84jrJD4Og5T8PwWMvelJTXNGpP51BwyU5953NV3ispZPCb9DPzVSoDmkGT1GJLYcAx/8SrJXHOc
c2eqdtcPb6OPgnZjokBZzaljjqqv4ecMNHh6PWj9XwC5JgZLY3XS6/vwUgJ6l8tHdDKq+LpAxw2h
uL4vAKpwB2Cp+/Uls5you8uUgW7xO7eArb0SemE+FR1gLjkSwQ17x5k2BlGYwsG5jOKP8pUDpEOD
Ihp/vXnbLg5icqBm6hZPKsNn2WFoqlKZ+Y0o9GoQjsoX7sk6vkw0/WRAy5WbnEtFkTJOnnifTYu0
hIZPQ7smGLNUB61uFLsfU2kFjsdmpU26IwfEopbfTRug1D23OB5eWmol3yNigRGsfCXoD8ZZmkfK
37ti7xxvcnZnDdYIMYgd/0mazVhtKpBJYr6oEbLgidemIGuhQ1cBZlHBLgt71T7YTcFvY6FFEvT3
JwpYKMW1GnjoxVPoxu5XH7BuDKm0lP+OCxPbtF+rSJOd+JYogyoNdUikXBeGNYjene6dQhtC5T5R
DIWFnplfLe+LVskvhNF46yAsqYw8Cpcy6mXZgeXwNYDEEyCy917pFonwPsMIuNvUnjfHn2C/FlPp
9biuuskmiYSkBLpFwaVd+tYRUebxupJyNKHUNjrQ6t4AtlpdAl1qV43ovGQNDEyVHt//vkC0CgOg
Qz8FZn6i0dDS+11vSEu859/Po+zNMk8MRb6OrJVwpyexyZ1/63g/Tpq7uL9QV8+AEuWG3ccRbyha
vFm9jalIwH/c+05hg6WLsPFbxO3Bo94Dicmk7Lnvs0VpglhfEJ805MtduaoJgb0WOoVqkysVtx/z
KsU7vMLBE3JyeiUEX7MaO30ggPCQmqEiYZt1kJGPFUfaf1i60JwxPaCtIfPvaEgmNeHz5axD6omr
9RHIn8RowoMDj6PcAEP3adL04KYizPGtpScMZYcHCBThHYiGgZxSlfWmt1DvuZt4l6l5AMHK3uJP
M/74tM75u4ihYQC3+aqL6UTgFTJiXnGaDtg+hkPtrdTfBfuehSGM860vMTX+SODGhJDxsalat5co
IHHD5la1zFO1hA5PBT8cvxJ0QwoYukon7r/EdRymeJOs1e5oAFAMi+ADBTAB1/UlDdZ9K1pZCWSj
iVy6MyqXPJwbtS2pNZtswmeLO21ahYBNGr1Scpwj7UZ+EqhB143GDaLxeqDPNZHY4SWmHksDEju5
qVdRzYDIOR2IpAYbme2TxIyR/uUcfwWLcMXQkkqCWMX5rCh/s6/mKnCdpvRgtt7W9tRCVt+fgV0X
nGwtIaqc0r6nH3sC8WAsUokdlMSb3P/2GFi/0k5ZIeYrxx/e3quZJEQa8sTaaa6msilf9d//VXvn
AdR6SznZPAP4barPqiMaZL9/hBzkVSrlybfxCtDyyOaISHlRVy0rd49Jg106Q31dWyFtwmKQV1rw
toDekoMy6mTZp+UGdEx/Zo+yIqruMSxFFbJ2XZ/KkLG49cx9idLdXSCPfz1V4Q+tfgMPViOGGim/
tsa3wWcFuEBA8o0GZ8rgeYcOWPkIYmYBdBsr6sQnMVpyGy2b1JVt6VDhoryo8rmdNPstArYmuh4m
dV+RRiRQWb3Sp6MeAE5SUKDIzIPLZ9dcmN/bOMb+C8hosQpBOS8hY6qbJBYrZ0u6UU8mtnyoUAR9
/w1zyD8Ys4aB3LzK8DWlPyG4OKdDPVOs7GPzAuCq3QKoe/guLWoUUdX2RBdfjh223N3uM9fWMn3u
1ZNUSGrmLm+lNgjmq9AfGf8gAvwsdMcecCzRzMP0Bu+f4yINE8ypOwd9Mo0kIOg5KXxvxDEIbpd3
wyp6C+T2yMfmqqkva6NUVHPTM/eSGcDqQ35Xv6Imn+z03WN13O7OG2kfB0lk/E4Ti3wbXD8cf14T
ADppAfvh5i7VYxgIOFJcyteLlf11T2LGQWnYIueyRnXNMmU/D4PYQdjgL1+SNvfDp7HtY6oVM4pP
KoRY/ZICF2rwp6+H6Iwi8GsLsZ+JlRBjtUNzD/yjHKS3htPkWmfA8M5pShFzlqYGZx4wRrtS6y3J
zyh4YLNn63Q5efUjkvFhop3nZr1A3UeGx1xtt4p4V6nd1yON5TqTtBDuOydzeld5aTDipkAA8xYb
NFYEipy7OXH260mjxAHVecHQdSAwhBCNQ49CNz5y8CiRP0ST9m+Kpjv/r0NmCVOlPsjslKrzTlY6
ot24Aqt2DQ2ljOU/atHru+C4bqgJQ//1lIX51ItJ/Lo48UXoHmpNS5RxOCDQqtil2Ibo2W1FJi6K
Km+ptnr+aeujqWbYhsXqyYn5gl9A3BZ1uQhyqfRD3dVG8OozMLbmL57zna2nHZXaUOzpIua0C9U3
iB4oDU8y7WXNCRydRivyY0UvcAB+rvxNd3mnqi9XHRNze1LaxYLWdqGPJZduMujqPj7SL2b9UT16
bHur226By7dD167Ai54RmURjlaIYfrZBSA2uwWytdqgxZSwBtQNUQ/WM2ZoB3ikVzThBOtTpTt2L
QtAzU67Uu9nNqdt4T1Igkb/mnHyIPVloXuV4qo1dR2rPAUuaH7wj+lF4SdXG4l1P4iAW/HCn/YRm
nZYoVOB8x1e3CI9/uCTjq3Xkrq1ULIk5fsfUarLo7dXz5EqkIQ3L52g1i9tqowqeo7iHhpouMFRo
6PqAvNpWBWd6ntF1M6Qhhzd1+V7TnPIQVrnFRddWicuiO+ndWSHLmaUMk08yJx45pkQHF1b2YSRg
gmshk0xkQZG2IOydjznaaBoCHr0ea0JKP6XgPqvceIwn8AwzFBlwSIjPt72f/jT8PIWXthK16Yv6
J+RNGAZ3sz5wh7Ujyx9JoKyyRUwaGFlRg6m2Mwwnys46h8fIdub3cXZsuWQF+S7/qUPKHcl8u4UR
4f2sgQLpQp60f4MbB9H8nJVCjQEpBfBqubaOZw7JGff7OQb2NvaY+a4LljqMLJ/PPYkrzdfiJHaO
T6XRRujL1l7xyvLvMx/QVqudSNFklRDD9JPtxhzLJGe2O8DNP4VJVRc8209wPYI4P39TTNdC+zgs
MMS/9V+e+MeRRDRzmEC/9C+rPokCYJds+ZoU1YPX+OP0XLwFxEuO36bBXd1lyg0pu4/9JfVKqZOa
WjteosrOmqtzGxs4pvnMD9MKKubbKjeO21UXf8kQ2yuqCzWDWo1YT/qjQC/CqLsplpD0md82Cmzp
Jmuo8nHuw9r/C2Bf/wkf0XoHlKGBoV8wdjx5QVbRHW5jpcNaJne18xGdCd5LPKXUHITxzujYGOTM
tBMV3aAJBpKbRMqKHVJTbPLM8c+WbpJq9KL4ZaBLNc4dq4ZEWKpaSbXVEBADpFsHKV2eAV0hvZS1
jYpYdcEnLYjIT/5A0E/6DmdY5gRx8oZBAT/ypRofLTE9BYr7DuiNPb9y8DjCJXkeqkd47XrbWn8r
Q+YNZQMfSfr+IYEkSUYramZ08CKaTZpqO2gWxz8frEU7MCJExeODhCKbsfZ6AT+VE4b8Jt2k/FOb
cTNKOsfWCc+0H4b1YuMQYMSg97ZheS/YHz/qCe73P1UsvKoIQFldKc+nH7A8zyfFq6taGU9gQnwl
2Zp5Vgbz2zqKntC03NLAcnQK6ngstZ3CFBH4LR3gaaNhZtQwiW6F8E5gYJMBZR8f8O87dff4n+lb
asBu3A93agx54P63OGhnkUmP74XZxi/qLIETKGF/3MuzEAuh2SUyPx8ziu/E5QaMDF8q5Jzzobyf
YbMiijxQIgUKlY4mRyA80YiHQlnuC1qVFVCcnMUfhRGP7PUdufUiNLjtociO1LfWavbjfrY9l5V7
gm0+k298tKXZiLE4UnwWUFVMy9f8NIjL5/I7sEDJPyK3a6rxVaoIjIBYoLOvDJqvDA8hwK5dR8c7
c0mmNicgHEgjLEhKvG5ynRc1v32T/dXgiAufKb9DSRrRceEygpoPhG6jM4xTwcGwufzwd8NdqcRz
mgtHD6lemrMtvd7CC3HzAOPz6iHKoDgk7+bNlIkX+dQIKn7zO0YH5wigEZMmPoU5QeIwDYB0Wkuv
Pm0UsW6ZykaxhPcaqLrt6LhhMsY61ioFL+JDt5rjS3luewXz+h7m4Ujo1zRxg0sD2TBVS/A8cV7z
csNsrECpczi3vYUyY6njecbLJwPAlU+HyAoDJX4dX5SXoMFuLB0tYlvP0s3gYA0SQVlR413p0kET
023v4UYXXJ57dDaNlzq1oq9RUeGXmS54rrfTL070qjYUZuqinzWnXOxOXbOZyyXvfmR24pHHNL+s
/jtRt5UwCmaJm6YX5bsVQyHcXT/n14lI7e5Ks9lKeDhQ1IyZW4PRSyB7ntRZ+0aChukD8hTP2exy
WD2nt+z767ME7CiQicvAQIBbnf/SYAlaQauY6GSGsWsqHY86U59OZuPLKIsDbjLuvUghkatWNbWI
Ssbd3O/fftyzkRaTpTE/m83lh26AQ8ExKZpYTXw3k/QRsKW/MC+k34x3avPLPBeUXac8EAr/V6tC
KL9KhImGEiKgwaJe0oOslr1j261BooVC2wWQVmypzlUeY/TCEM2dhBDSbeH92Dbq3XwBt+Ji3wkW
IF1H069p0siYgexGpwxkmcePUyXSK0pjYlar9vPlpjU5YIji39chAKnrkFSLqHBuGJVYKUBOyFl6
i5ktU6C68bK4YMBY3c9pEtzu/uEYrm+7m45102d2ggYMVULHvx/FqOB8fkZsQWm+j4ag65c6tCam
fjhVNwgl/4xWPpwMUcunWK6c6+lhjDhZv5ZYLJHXLYxbny+6Dx0WBkRS1lW9C4Kjr72RVS5t/w86
YIFhPur9BAcfTSPVWfnv35VqJzD9vlVNoI8K7/bRSLa3/WN/r8GkjkJeTiqAVTwTtL9/evxgr+YE
7T5siQWmK86LNs5PW1kJIyXow6B46EtOIGcHgeUxnH69ttow4/uUL02RmoZN0pfZ5JXb4VImdck+
ZxC9jQ35kr50+uQi4e5YKEbEiHL2JezZMlFNL/xvr4kwVqV3nMDC33krXhD7Nfs/4VTuCz0ENWZh
Do7uXXREwZyytA66Q+oaURo/f9Dt7wLhrB6fuUgQ+iQRGsCZ8tqQHGbndSI8j5O/NXRFBP9wDjX7
3XxzX6sF5srBqDZTn/DPmiUEUDDVi0LfEwHJ1grqj21qp3sjqd3hulerL+/33+gWewBIM6IEnAky
HWlBxbQCmmynIX3F25W3Ym1/cfQwSOQhh2tTm9nR0HGvCMMVIbiRDpAd1lab7naj1CkaKpyQqL0K
tTFLPGlKnrVCpECRWyR6AXiDUCMurB0N31MZdL83BnVd6v0Bdxp/Az/uOKd+Kr2xi0qRNOp6g1/E
h1/jVOx9Wp1pdYWEvkCTCc3z0/HmgswDKYKlESdx1EFZc9Zhp5DmU3vHK6oIEVtpGzgmHgDjFOnp
5ISHtY3Gtep2RXecL9NXNVADGbsjHdIPi1cSa9UslAUi3ZhjnqZKjF9+a76NPJLeP9kfn1Hd+ZxE
Ik9gIc2TnqKoqek612P6lAjCD74zsTllsJgaOHz1Q2ME7a8Up/OPSh3Ahmdy4oDaTbZx/uOAKm2j
jWWuw4OEfCYJiQmuhEiM9P5BKXyeCZ8V9vuoc+7PD9w7xrIKg0tfQxVEKvYMT2w4LVZQq58ktAdN
l4z9sbfc8HSov19hPQ7RdgMXRWb/6+DJSycQGqK4FehJt0hvl0uSGV4vuLvydKgMH1uEEjI+AZZz
L3yP+NnEMgQaDsTG0z5M19CCN1+UhcBMfi2M+p+IuagMPW+9l5yTIiwYffRs+bs7OzRO85lWpMLQ
YeZvhncB4SyUojjrmZlZbiW9XEbpx8mrlod907Du+2J9dW6rSvIiKho9l2zxEoUISbh6J0lNAhQf
db6QH/GZHfeWTN0/O210LnOFI38rcXJZwF9u2nd7hnilHpKO5FHFxudxUhnJdK4igDxOX6EoHKPl
YtQjeeth8H96jqa6ERdm22U6paPnH09uS+ujYUSxKQtXT4mZUcKdnMHbk6fIhzYVf0vRzs7IpdUw
RgHlogHbUDJYoRnU68eAzs9tbxlXAZkHMgKspIp9D1h0NDqaTV4P3gQGmeLwzW0fHOsUfhLZ6zk2
RyxxJ+RQXRmmqeG/QQn37LQEcpaphpWR88tSosSwze3aHuP4Oym12fZiyLahbh8Y8euZEaMhmxLl
wvBn54TJA3V6kljb/t2C+DHNJF5jSvdvBlg3W+lqefaZPOoJN/djZDnF9LVPqRz0m8hfNG+tBgeX
ItplcdkL20fnMpTZTX+YQtWA4vuFP9p6jEmHuG2uCLQwFIuaNafdrat2cmh7vMbrIlctfkT3eE1b
ng3BbQo4YGMO3AQB/oxZw3lfpqSREkdsHtaTcUGTAnqoQLpViGdKgQEZJ+vZicZgIPAh1tji0XG+
vexbggN1S7ykc0M8ANL9lzStOp0mnLAc0/161oGOOrvsopXz7adZziyiNIdF3qTY/JvdLRzXyY7y
hRQdgEf6Of/Nni51Ah3OKp3jXCn7tbJHqEeKtNCJAh/siuYFbSue18hG6vBfvgZ3Ng4VIKbSpaXP
8XQXTKbjukUa/oHsMp6FOX62O7J422bCQmDUbuZOWzE7A3NxGM9OOI95J/kKhtzA46fCD37bdn57
prVG0Xr1oKSOYQv1dn6THSlGMbsVAjiTpnSwxrK3c5CFppkrLk1Dimov87L9Nwzyhqf6yliiHpqJ
XCqr7hDpsUte05EsUIflYLuYOwziqjdP1sxlD4k6SOMR/1vREcfarz04iFIwuWKbTeNi7yVyX2Wz
gQDPbVw0leRYKbtgOSSTVeQt5B2WZNv5XXI/VmhBhQ61DxAUQmIoaMIh/iwHrY/VpzSQTgox+fxI
r0J3yny+MMM/xspmpRASaxx0MWtQm1IiB1KV2nfGwRso9jjRzUa7BSW1Su5csmXm/hMyIM9ijdjt
TRnbqO+OvyRWOjybjdtY0ARVd7FanBFyFo9rS9S/RSN/c13zt7+rj2k0NmuWkAp9yh0wvun132F1
1oJC0O/taynesklalePnYt9FMH9KwUviNZl3nre2I1B5HxkxcaG852/Lfy1n0D1vde5lHRoBkpop
8twRcv2YeCnncC6q5yR7KO6qbGl5nXFUvY8AFtrGmlzFSUPC7QmpD57Co6fLCCvt2Qq3UfnMuQ69
yHqBmHzBzoUdP5CpEEOEUz+Uc7TlImCUroD/A9VjKJYvwg6ROk/ZuI6+djtIqji+evAi32lhLAL0
tw8OL9joWg9HlLK6uJ1tylXFg86gxi6FsbqCH9omDUZNxEvFMo84Rab1ngmcAAezLBlSgaYK4KzA
Q4vk420zVD3l1K7olzf9E/W8kfX1dSFsXZTO40f4dDEpmLa/exJ2Tj0lfITg0Ik+Z8VFsve0Jm6w
mL69o75w2cdNoK275Lj9khtm5vp00apPYivFMKXm56lJAfWtudjnlFVF5Gr9j9ZEmN/yiXj92wt3
0vIWP9kvgyAozifiedk9SavrGZoFL2GAFkrwjGnNyens4ci+ZVGVKLgLyHhxROMvT20Yqe97cegX
zhRtD3Dbq30wqhcdJMhmENs0J7dOXqH5ca0Jb4u9dpdBh9wwLt0ziK6IPN85V4VjlW4cI9LyjX0n
ZbF173QYDXj0FAevL9aRkvIDyKZZ4SvXVbsHTo/epSe28Kdsb36oGSUQoZ02e1uhzn9JNJn7Hg+A
qTT3QjUYN+YKHvHTirRfRsmassGUm+bnn9MvFtrqzm0zienHujJMCJOUdvqfAFMHIauXj0xJsJd8
YZNSyrENzRnrhRjn0rx+ldxV5HaVL/ftONBJbh0XbOsyhbmPldc2H9YXuvMi3MTF2dZf9K9wCc40
gzhd3E2kACJwJnq+xqEiYmWtrSzzisedmcODEjTb4Q/Q95lvt60cctbs1gqlNq4j4yd5Y83RdZyI
sPp3X6cBjk+xoIvVFj2KfrTqotwpyx9AU0Ntt5WekdjpYHFktpuVolOl0Ayabj4YHF+kpiUnuH11
v365fqzIsYGI2M1WtpObL7Z3QOJLVXXTeM7uz+et/YDPGDnnCIpfDLlX7Gu5SBVpwLHSm8GgT9Sw
DR1s3d3faZUOSZGoAPooyDtZC7bf7EYTBuQBCtr0semOOsTwrjGCAJAHXPJQ/3CIYhQFk3at/Cv3
IVRvThr4EkSsUKszx7ttFP8jmmE+4JNaOewXNHaQED/MXHb2AvPqaBhwU8UZi0XfuyjDfSwesl8F
5BP2FS/j98PjVozhW9m0Ck0Yi+QQzUn4Vkmtx/3pCl3xnGvknTk8K8k2JODkhXzm40LBqlLEEuf/
5Y4CrW2I/tFJIRr2wl/ztRVMvs0d0R+T6YkoAQ3EnRhE2tXK/N/wTCP2bKaCkte/B4ZTpeMMinAz
heWdR2JAS/CiCh2T7sx5nRNnwdZDiLf5xgs6MnCNBtjUz181v4iAjZkw+PpGy5beN1GStmpLXt21
zqo/j8ebEw3GIHqSA0D7FbWhI8BZMVVSsQgP6TIXqSoRPvz5AsuWko30m1dyrTS2C+6r9LluiTrW
eXZNFw66XTVBp+7rrgdTPE/nR9vHmvjsaY+eypEAFpkByBWm3Tx5/2rzy7oY4kVSkLilDfZvr5k7
Hq5KrFLIb4bwdr2Y2CEigjkhx60F2YHOPjdhSVk3FyCs6FDh7ppBK6Rp4C49tnkuUPlAF9D+WFsX
mCyx5rsYt0Rye821b8nnY6hJeS7Qixrg3Nd6NUne0076HnuqHlgZcL73HBgnwtK+/y1GEZ+ShILP
fKW/GsCJPb3vPehCFMxfMWDWskFNYJKz2vU0BsaCBVoYORsTiJfAMkUA06zMpNSXajvhSNkqT7La
2i0AtMOFojz30R611hE3zqOA1u52Mer9SAbl3Safc1/xxg7fxZqtHCkEPiszXqPwDmzwTqt8q0Xo
SoQt0tmb96CQ64XrR0y1uXprFUrTwimk/+FthXwrxDhb3OOjIdzNBJ0aDf5nqYgg1p4HGh1yiZ3V
/43bYhVrsG3R9PgsEboV0dC/D2V2wWn/JdSpAdTpvVRk/+nM2OSdb8xWZudEg3FrqgBw5PPs/DQm
JK7cWx2vqb0j5Ir2TKM3dCimWL8ucE5U+s3ucPDC5vqE1zLvGtJOGkQlowRR+qizSxTzR2tjMBh5
6t6otOJ+eAj854KhaUvsOtMXTnRypbzZQp4CU1eX1bQAKtOcXKKRnoWoX9p6wWJYocxC7C3ldMCl
aALX0AMcnZbL4tPzjSBDj2xwkSJZqb4Alf6TkiWRI/4bZZ6yOqeVFnXrA3ysaGhoxGmWx3bGjQea
CVrS/WJSrofMAXgjNZuN00rz5wDhSWVbYlXVaKjKsqVtQOZL+Pxi6Jg4aiHdTnoqVyaJ2f4aYJlO
rEukxA0IdSy6iY0GPBEdZSM+U4iaP/JEF1N1uwxFOBY26lOOXPTx+9S1VQI2y7+Zu23XEuDD2uhv
GinVVLI4/Om0UpNBrwW1MyuTgrrjcQElvC+L/uqAYAbxDBYVYyce6zyw4SHaEqn4cyYVda7cZd0m
6+XNT9AlHW/QQu+NOA3aeZ2lHglaJaxY/FhiHWozPDwxJnLsCjRuftdmhpVeObsa8QsY5KWebwZK
JG9Yvln2mD434I5tRLSNcN1Uq5qtBdXMdBTZ48Ua+PJz6oaaKhySsX/LP/A/36ZcxT1jgUwFVymj
BUnZq36divixrI0tMdCVrJhNP1lRRkVIyK0rNMFjp7I5JC/JaT30j2/NgDjqDZQgW/696QIDVtyz
O7xrOd7Jy3Eomwln20OtV1LTs9HXJLQfD2I1oUiJgaGACnQplo89KixPqijTPfKIQmn7Ray4yNYB
aFfA8iUIKTbQ5ws+Pqlzwxijrg+kvWlUNOP2bgrCwM6b4CC/WhoOfAQB5LOJ6ztD+NhpsQa0fl1E
aJF/keB3Zjc6rf5o31zPbslP3oMWZDC1TuGibKJvt4GUrkrgP81onIIKdILXvrlLUEmocaT2+mBL
je78+dJwn7zpJQIxwFD+gg18VUpegr+STIvsBdkPaQA54jMV/YwJQnTUNIF+3+fcvXstwry7AM07
XKN2p0c/zRZWm7x1DOLVDFbLgb5nJvRvQvdh/1bY0nexGJHnZ6Bc/0RBL5Uu6Cod4VtJ6Q6uSW87
I8nrT5ySjDVU/5OS5eiicQ2y4Z96QdqnKWql8bwNERBtc8sQ2EYVHeqwNnBI+TmHJzZhwvX+3pyl
agNpKY+plzZBgDpt3uikTWMYr0b/uxOGbvWmqKo7DzX0gYmfGHuMaD0D05/SXUupFhV0TEKfCHcT
fYgaaaWltjpZYEaEkRWXs2mcIQgZWjK7+vJ6Xvj+9rvVsm0gwTqC5GEO9orT9AEIM3UXmkoJXnlq
gQcULCyjme3czRBglzwr2yookAlb1zMKXZW1OxXGBg+l+PK4UNCtYIJyjxYJyohYM2ZfFRpNylOJ
/uAralqZKDPH/C5yV0lpjiveEGaCgxrqniDM/Lz3v4QUuu8+Lw6hhanfYBjxphtt3Vn0EX4o5jio
2Kwo6sMSHg4zwnJR1qYCDfYPgBqUzUqZIeF26XAfFZEWCIbajzvUM8P3puH81CB73uVj2+6iD2mr
IiDErrBP/Tl/398jFxK0PWE8sbEbo+OOa8KbYYKawxw1jzvGHtcF1Btx9buXYrs9DwIVJFe8C0vD
yL9YjoL/CZGbCy3cPO3vAkh6cepba3zf6yegZP9dbmhNgZFSQwTlrOUZahQO7vHJ8w852VIEQWdl
5JCe67dIbNFW/N1EvWtoOIMZaoLR6z41ZYvGe26iormJ6Aw+lkV6IhPIDNFwwAZqJsjPyULPST5U
MTK4KfTOOfeeGtxUBfj3dSGiJ1nMUa+PATrQS4E3WwvQB5Ny1ssgLCKbiV5UsZO3lCIW/TTNyVMu
wMUANoU2Gp8hrsqAS0z2p6TDRl3OUIHOyXAYztXoe8NrVF/5YH+SoGiijFBtMZyPh4C93ovQ7dNC
/NVkAvpDTLExt5BoDuPvJt9K7E9Vy2+950kflfwJu8CUcgEQeQlmG5WwquT3jzEao2v6/iVAvjrM
M1Va2v0i7y7Uuacu86wDWDbNgbUHvzed+zxfcA4Rh9LDIJcMAMNgSWRZdHmo2DFmWx3drnIzX0C7
4ANDl9nFZOg+lzYOkK4VqE89K00AD575EpepN1pYUs3rOVzIA5L7iHQ136OxfMa3bQomOc2FcvSX
jM8AapdDi8Jwt6/4C0/C8IWsZW8h27oT55QFNZAl4snMOji1/ONogl1bskcQga6aIQdYwNFgox86
hlimu1bKEBGbGn+/OJl91OQoPyxBcSaE5hzeOCOrAGpKMwzF97yIf1js+vejs7pUWohXFvaW4hVT
djKBS4icsTmeadAn415AAsR1GqSm9qIYQdgViuqU5Fa0l0cMcJHlTTRQw0udxnGXchlqo+bMRyqV
NZ7Hm6CRspFeC8C1X0TeGPzrbvaCkBuagSZ+gOeQ5m2gyADHCGE+0HZnxkhNMP/KsDd9w7HgUcQJ
bkRiNZ3rVAikJtTS4dVxL6IaeQbEnUgmbwopUIhGA6E3a6jSxt5JYcciOojzHYZDm85e6UpmHvDJ
J9STT3ivRZpfCxDgxRsCL0H0JnLQBpqWWsTK31q4eGNOELn39DDmPHmcN6JITX/HOE0mVY1VpBlh
/IFhZyL3BuYJFHl8FdnDjoZbRelPx1oXrpUYTtVXpEaoy2eiyFtYfo5iqwyz8k5dzXEl2uGfKn19
0N/Xt2BafFoKYs7BvimzH58DeI3fijFN/YpK2dR8WaIYyMmf6dIBUprp4LAH1D+oMznadepCn3o/
jjBqS/Dkw3X9uHxuRsfShs0RHUp9Sd7M3BTIDql2L7a+N/q/GP7vW+zca55sbekv6cWUBUQO5xDo
0ueWow82UVzOXhmholKCMtyUupWnGyT3j0N99zyiRLgvySSaaTo7GJ2HSfFJjOuKrOAA1jTxa0PQ
MUtHEyOYnerFN6rwdibP/huFl5I8Irr6GfBZkdmBCBgvDrJ75LpeNZfkFMIlODLb7zcx7D3b6XNx
E3cO050XvV0HgvVf09m/wSaO9Ty7O+Xz7rxjmATHh5LoxJYuaJofTFU4M2UZOnSWENHYMQUUW8fh
VLQoJevWlhqas5NzJD5D5bZWmzA9Y1B0/1RRnlkqCin6tOEkiBDKg/jSg9dr3n15JlIyAmayv33c
qvotCua+F8pOYuP4wdbzcHy2JScluWN3S1nWP4+IpQEvrw14DAz16DAowWxEy50TCttzGbM872a5
hi69WAzs6MYSdf1HEz8AWJzIemcAWrNjCZoAAb6bhUT+kFv1Wlqv6LTYbEznVq2WKQknUqcdWafX
AmVI4zGY+vLL68fePpxAaHhZHL0RSVyk5JHZuFe/TL4G24aNSqMPSZPuxze5ZNDOu1chwAjAlCaF
S6lWWX1NwNDd8tUA1aZMkVeTLWgWPdVu8EPvMp2n+usoDmvGl8Jj2Oi0SG0jkwJOVx5F1xjm2Q1o
OQJRse+jETBPhF8ixwAM93YSAjZtxfvgNvTXW1vTIk0F4ykOdTtohMjiokmkOY/EgF3mkQ9PifCO
nQFSmwqU7TEJbN96jcKVJ4tjXYDR8WrAIqj5PgAx6PvCBbk+aEC2YnMYqd4tw2Ip7xJtSJydnskI
5ZFBJCUGWZU0pTd2yk8k+T59tbifEhX2dYv5IHcdljGHNgoPF0AvAPWq1u4oHYUj5HjyF7TzkpWU
Fl54e/93FQEBTXBW38w8yd+T8C84xtcGueuo+XDn5Sq/SYp7XxsxaxUz0pQ7BD1BWoTzloJf5Hed
5hqV7/exKF4YBb35/A91jpxws1ZqTrdH3xpIQNwzDI1Ut6G+rI7l+UdEu+IHOWbuai/Wr57SdV4B
ymr1Bv06xTCyrqX2e20CdoLCb+xU9gqDZc/dlNUDc0aVFcb8DD2lsyySXK8/Ax3ZTUN/8c5HKsEp
9uu6J6zH1uBCKIDIpntp+iQzBYMzxTA4gqMWrWCTP8sFXo+fEG0hM9iIHM+rjPFj3vOUZRNELxua
dxe9A0nrNieeGUnGc58lnHtj19G+g7bQPmPaOrpKxpWpa9xwSBZR4yZzV2tDijaMid0/ADtkaotv
+tvqMMRpnhZ5CfVqRd8M4v/oSeKXcfs0SYmoNIrV/FCPLkbcZbG3Iv04RmvGN/1duAt3yxOjBwE1
rZQRv82tZMQ60n9cae1qkqYFXbnMddRON/sbZFVS4oSVtj7F8K+iFBXoAb8K6aizuxRDsqFLAxmJ
0Kk8vlvqb0zSb79kHBh/ip2s34RNP5U04QGwNGZNRHcPvI1Iofo49T04CR/BGV74pJjsdi4aaLHe
uGYXp+hOyf3iigBPUVsVnF8bCq+UZDcCEuY7PLaR3OBHS8T1RItPrFCbXaW5iCb30utM4JoTQ3cG
VZH0cXlq2XM7Hy7ZVd9XgbLfvR+qViRMnahzurpYvVYEhW3DtHfj2MjuST6M9ChHoa0n2QOJP1IM
jSj8hcm3TqaHfTjbFRTB/oS2Hg59kfxXTqPmzFt3U4O/ygE+IHgCoKTQNJu0o1akGlys+Vr/rskR
rLgxdbcd/4QFUWaC/W2WwgZctMqSYiXy/GfAaaDQqZIlMVgAI8ZATkyne/66Gixf1LpLzvc4I4yb
GunarpmJSP8nn/jaG/epapWcqWjtagIdOsQXTa87ECJXwU8rkaIPvInj9s51MojJ62m2G1xPBANU
IbAEGhTahZ4qkL0R+8sWz9b3wsWcjzdGdo4eKpfJwcRak/IXRmZU7cODzXHXDhrj1iR/t5VAYbeF
22Me3GxPWrSXPzV2G9HtRlZJU+sx2rSOsMfzcaYrRMC2B2LTWFPurz+5yQ9fZT+WpCA7FS3Btt3y
qtKZhPdl3K9BVXSbXaQB65DrYaZbXKsh5ac08kqRY4N5GCwKi/FwEJLD9S1V2kuATh0DdvNdhQhk
a6auoBpg58mB3vF5fOmiI5dKbyLzNcv/8C1k6QIDVRz9LT58EmUneb7S6qHhTaZXQrJUO86WdYGh
jzfi9DITwK8HIhnDG2QBWgCJWRPI+8Z42cvMXO9GU3/uE4PTZ19XP8HMjQbeqTkZ8QOMYiUo18oe
Dfra7b637IUCHrKH4oV+HnmJglbTt3SMcUHl00uXORww4dtMwGz00HdoXDbzYkOrOnG/14073/zH
TPN/S/silmKXG++MxDoRi2w/nlBAESBGF/4oC01oB3CVC6PNU6U6JgzG0v5/ctNwyAdv85GhmJrc
cN/8z82CIoEVuabb6CywYA2zxWRhb9Z3S8Z6+5Ltb5UwjjtrEvlY7sxGrm45LVH5WxTbIZWvlwse
huoeZzKQ+Wu/oRX50OD/cQl0s4pesYJjH7G2vbcxWUExk4i5KGjReLluhp1rznA88MmUWCAIIbbi
T0ZuFVHrq/2MxjyoaJngQ7sjeARmrjV1/uEP1D+tIIsD67Oe9exeJr1eq4YntxcD3uLpEB3F0QDu
wMe3YzIhSfRa2qlmeAlj+JIxTRhRRdLQRzWVpaHgORrOOTATc0VQ1hUxLDnlKCOfMOMUfc9mJTGS
iKk6rBTrbLBO7E2YoM6JoUvU5l+xAlM3gS5BWjQGp40/cD88lZZUMZddbw5d9P5LBwFf44QAIebe
NWJPovOKZExwwp0uE3xsKDALiHY42iaeld4annnGJpDFIHIXu9jVmFRTbkgAb4GbHmie5jolSQKM
DpawkTmY87WceEHFWpWPArqJCdTCwwWQV3MNdfLPBclLYNb5K3jrOPwZrkXmVnHNR4BjosiSSAA7
98BhmPC5PAUpBR5aZnkLh3ewrQIdLnrJ+7h+YY1DdM7fmM0gOGqWu1HloU/o12opYohtF/uU/pMO
zODYQdx1NlVsQZ5SJfDJpoG8y3oFx1W1Q00WZnmOWtDmE8RWllcOgUNUpxUaNVaOr6GUNSswqBR2
3kXWVUl4ucaPPbrwg2RP6eiTcgSb3Xof+iFIPBs1YRiGAsd7EdRIzxld4hhZpeU+fHYyNGXAVG0V
DdHsJ+kZLZ+H5S0nXbiD6WeLgZOGzLkLl5UoXtN0PxDkPhdAkOdZc6umcE5+mQKHGEbuzYtt+vZt
nNG7KjY7LtfDaD2/nMBRSOrTzWEW3otVQNcXDvjOXqvIUu4xv4nP6ljCj8eG5eMWuYHWCqVFwR7E
1b/DxOt5zgIrEkDXtGs3ixXEwMbOs8u19ie52g6AwL3iUD0shGEORtNLeJ3WDewMjXqm+5Q+yz6z
aZ89npTpeweOhGsyGxo7CSp4thcBTEBBq8w2ZbHpyZ7wJDZTcK2srszWiXZba17+gzv+sGIN6Xif
lBQGLLjeu19Vclbrw7TDTjiJhLYnRaJOh1C8W1sXUsBY1Ot5YeBuNW06Vz+silPiTLJdj2rSCss4
+PWdw34EdLlXuTC1Dg0WYVqAsP7vEF5GY7/ICx58WBN9td7/QgHbBIxBHbg4ugp37awG2GNoM3YJ
AxKxANZ4Nhna0moKpnkTV/I0Rl8JaQBIsHU9w3rXxKUM0zs90QhCMRq2fOkFiV4/D0PvSEzJrt+d
i3CWpXCZKXQBdz22w17naFS4YspxcGheefUWqPH09hJRrw+pclPIkVDIjrQn0o4t1hvTu23zWJOp
auf2ttwZmaEihQRUUYlnntt9rEaA9sukj8yIA6izk4nmeZUOwjbxlR+AfVkPg0073rQpM6IxMIwI
BlfLPoun9zLHbR/hkj47oguc84mqP9Yl57OLtco6Jeg5SwV9XCA5kNbmilCYJ6D8G9ketqAXu/2S
ikV1CUnhdRLwntQv/IUik6srb8yl+ERcscNX5X0NsUzio1glHLc9NtbYAFh8lIrSXhIKePMRITvQ
NA89RFZR7Lacf19MaR1xl28jW9/TQGb8GqPY9AU/4BjIdHd0QFqcxwv7GAqJKBCNZtruXAqvMn8o
0BcXdoMNYr2JrxmBlstC5NGoVdABwyacjanonBaYQ8TXxFL+ZhFGWZMiD8mSDkp0rkcnWbFLuJt4
NHV3a4IyP6PogVlejbqv0zXwxm011pus3JM5rMbmsdELbvxDyzIn7oUMBi/zdTwSb46bu2ALq79F
EGtlHjvlGrRMr/3IOlP5mDcXaqnSmOOyzniNFfjHf2NZqTG0d6OOmJFo+24w8F3RkoTFQya0ZOaD
Wviq57JSWZ/80RampThqC4plWC6l7OTkN58ODKl25r2JSAq3lTFcBmeVk9RDH6VX+BKYatnyryUW
dnhkaPLO9Ea+uVkz6/nHLc43FMxNT/hgR1EFA34AKukvM/31KiI/8r3g8wSRTf1B9qMM13dMRWWE
ZY6KBlMUooBKOi/0DYKLjL2ishCnEka4R6iQ+oHET7dI6TS6UhIpxGaw2Vyin25odFDYteB5KxfH
ALkITmqmHzclS4cl+UngpbyAjD2GOfoCDCURklNxInWHxg7AREU4lletFdqRXVhnKErAJ4eP6JD5
TegQ4GDBuwAR1PDHUidzZe3vVtusTcqeGvANLmUNZM6pEuBdpF/0XzNbVqmJzc77pbhl4e9TRgIX
MsXyiQeMm2Cv+Iap3wlrr6+AuBvBtjfdW15g2Zwi3VWLTegnX9acsQomVocAxLBgw9vd4UbY37ov
evxPCQUQ1AEQsGw44roVY1gKB2n7I5qOcKNNVbf3TUrlrZoUntgOwIji5AWFeCd8xikAdtwLNqCP
+ewbHZrhzAq+7NZYQBhWY9MJcbbS4YilGaQ4cvM8eYfUrgMLtvBiIXAbvFdgu4jvawpfm6a4csuz
U4R2ZYFtQqKCKQkCsto2OCoiZuEr9ZnEZqW+EvxbOyJo2dTbQIiAl8J+rQbyW72nIGO3ZHDvEUVZ
+GRCOueqFKl0pSarpQpocaEkAmjII6QwDeb/h+nNi+DoImbdFLnwjUnhe6wsyseSvy9Pkd+8+pgA
DoQh2mFbsuWcYsB9QJVVaPrefZRdbEtgAUd70dTBUG2Z4MbFqNGieHEBVdYL9sIfY/aTK8SEc2Rr
BuwbosTmytBmBrKXQJHbOvRTX6mlqOk2iLmXFndZwlYVFCG/7BbouM6fvijYRtQ9TbVTsTaada96
3UtkkrFIeHadFj0SN1vmNgnZGlsXDovgh0E5UhAP3E5zkliyu62aZ/OrU5iGChTjiNbgu/oAtGDl
BeHKG6DCo7yw098VY60CgZdF/p4rUjSWwTO/GYZ7DU/WqXXWKf1mWAnQedUrLRoDHP/9wpk6rmkq
a1wf55nsOsISXVdkAKKXDR0WaERxjQjw7kYqdEF42mq9zQXXqA+i5B904UbGM5bV71q1zfsmUU3C
SMczRJICGPzoH63nku/rnbfIIIBYhx78Nh7Pp51cpjdXE3ByoIfVfPxDcETQpSpjx6Ld3erW+jqJ
64lLVFgWlhTOjOlJBW65Ck72GY/f6s3OuAmv+KwVygn8Q7o0y7qondhaZ6noHkxKrx/CrCogJM0q
G3mGkPih8VAVYIInsypXeUmGzUpQeC6xnq7LXnsc0wotphMsZG4GPb8Xb3h0JXc1NH9zZ5GRC2nE
K4MpG+Fs9bHPFj1GqPZPAyGEzUBCP4W7BrFiMm2rOW+mx1Bt0jhoOWHjbpsRzzlB9vb8cnyR8RQy
bv1LfTAZcKMUihINYXu+L6sYbtWFoFOMqUVNCBrb6JESpAQynKwt/mzPIFj52cS08v0Hb1MCZA1X
BmP/wvmOlcanr4304O4LjJ40zc2h9Zocp/FPQUkjeAPf9I8irTBJ5DNpJ9OHR5XALANtmLFBdLDY
Zfh605ggfeAaIjQIrz4loqU/YJ1u6hk6fU4cljORDQHeJM+fAspCoJFWA5VUER06pgSqjyn008z0
8+Ush5AIezY8SZhfFZ97d8G0L1UcqIix3GqFk6z90+TCTM0ci8tWJaz7vGCB77Ul0TsegBB1MK1m
CT0bLauokFiX+W833HatiG5jffACDigm+GWkcw/VP1S6afmhlidGkLQoeef+fkQIv//UreI65pca
t9+IaanyD/py1+28Z3Zw46Hwq45JjFNhZjj2oDJ41xYJWxSqHv1QRkofrSZEy6jeBtJGaKt7nuxG
sFsgv6weR1kn8h/kvsHajdoWwbONxCJST3vPjAFlGwX0V/yAEyTkUbzjQc3yzfq87on3iVb1h4PZ
UeJCTeWwzj8JfY5Pi5zxuVntgGd+RJaH9VdqfHyoNc6oppEKVsp9FsScfl8+6iJ0PshBCrBF/IYe
/ocE71J7+2wYMaOjYR4hdA7TLhznzeMEmGb4QfmaySVw6Bwm0ZJFXECk6Qz3cf6OzSLO+jC4RqRP
UxQy3jYNhR2UWDDEhAtEfukmSu2KQE03l2CDfm9MKD8lXh/cQj8uEV7Su0PxguNSsmB7WtA9XZI4
0lhQtxvs1MZXnctYSBbCoZbMowNJ/dR4WI9YbKDUMOA6A0n6H0lk0vVQ/d5yIc5R7vZ/4KDX3ywG
W/f1VVMhu2h0iFgDKAbOJvvOMvd77zYJrk1jG45L7Lnmjgz2faEvsmv6L55bUJQL9zL2fstYjlhN
2lzbdLuVoljdczhx1aqzWeDrB+AiUzBmiMLIksoRd8lSS/Pp2cbcmo8WqrQY2v8OANkoi0tL9+6S
GxzLKK6kzWqYdz+iHk2X87g6ESevp79qblKnvr3BGTJ+OvSF/RsIVt8aqTTUTolpMyznnRjWaD4V
Gau45lxDw3+plumlIo8ICqmIkmLcl5OlPamyqHzlBLsiWd0sNWXqDrR+tNhEFkBgXBbdltHqAgc1
j31up46zXPKBqU8u85QNoOtKxjryYGi/OYu5gM2HQ4BeEhYuxUPn6jKy/BAeym0u8QEmxBCx/dXL
qcqAaUZ2wSvcUXSe/U6er463LndOMmmOqXG0gyWooCjbbThg6Wraa1gaQX8XEzJXk/xl/76qmLNd
wE4kzrfCkVU/ULJP8XK1cCqepSOBTw+RQgK7oEXmqj5sWVwRnwTYoHJIJwMWedS3nbQlSUOPLIO/
aa130aWIorkFSVFxzz1XHUmXR3c+/XSqCpVRD1jgHOYPdlDV2ft+2hoV0d5NuED0+q1DTchK0d2Y
Y34kdz2tltRifiQXWcBBx6x6RTJayVHrVwEH3kQQRSKohlkmEXSORi9angqEhMW6ksY5aCFRHTsR
ArwffooB85Xxr9G1M5TEtns7qlGpkj37p5yyWHeW2rSZbZypaCqzfLw6+uv7NLva+YFPq+NcKNP6
Cr7g2G0ilqU+f8zFyZHKtZrEHGioeXkdam1ycfD82gY7OMU9DRIm6iqQAJV7fF3oqqn9n5gvB+pb
1Ub0gNvaV5GsD7qfy9GhnGWKOOORlOONZRPVl0OaAiUyRtEY9zVEBs+vQMsWBXIFCNWHXyayy/J8
K4PCC519CD981OAK/in7/2MlBBD5131RqCX7euyj0bkDm+FKKWXVr08Niy3x8WFfG0eQ33uz/DC5
q7GqjaZS5p2Q1712ZbEIVjnoVC6o/MSDcPL3XOaa6ZdQHjtCCxVRxnJBc3v1YeThPemKhND7ugI4
RjNf09MPhja16YFZOjSLGo5xXuTtSLxo/85+seCQgR5eBBvSTdoUAnuyUU5AHymqF5ndkWAJikSv
E9x4rcVzCWb3UuFP4+rlYZxE4C1VA2lWSAZmtvIfwO3zYuFhMLxxRlqfJDJPEWwL2C2+HY8XuPpn
eSvrwf4UcUZl6GYU/h1ORogGMrXo5oK9zuXkvCJvvR9EyK0IZ1F9tI6Tvt9T6cVjO2MmIXlVZyL/
1wG3pNH6iGGCrshXbOyU8vZMYmFUipkr0De9TngjI085+YqudgXpnIturOfV4rAkKb9EWJINFHQ6
kJ7AARRLi9py1Hrn8+a3nmP6SO/pl6VWbPsWYzZLvecT+hUkXaBaBHYaRpW3bhUvfUXaSkx4sFRd
Wy3eEJ0yXXovKLbcQprSo+W7ujsFxL+H5WaM/NrtFmfGqg3NBw7XsNtqQzpXlR5dkMdwBfvfJbc+
OFrP2w2RxTVz59zG9s3M8MYAvC+pzMQQNiEFKs6vMukg8kfyW/BCPcmR5+nESDktdbIjUsjwro8z
aFXkOtGh3yldLkUmCWBnGYEN30o6+TjhAKHQU5U23xHxmRyyVd8ZYWA2kUIPDDkr3LJyOy54dm+u
aVpKB98PI3zVSVM6vdGHANka/FryHvgRCy4VSrXUsHL4cgy6ZXrbA9pDEEbpX2koCmxdODSXE/89
kXjd6tem6xh1HgDbhaMd9D4qeHodXYl1vqoBGu/aWTtbsYj8RQkiZecTdERFiS4UUoXRSs3XyW2z
fp2sJSETptJ5r7Gk/ssOQe/xFV1f/z69YfxfEOIzgNUm1Go35binapHo89qLw5EbWv0SWrrVnb8w
1nhuFa/7Xw0Kc0Hpid0dpTr1TkTZDBW9zOPhjBdYGGzbmRSdQbHR0FnQBWMFtsvOsnhWvz+NmPTS
tYZJa4VTXBd/7A1WbiLbBr80CAEs5AFfqZdnv1EbUaXfL+YdV0Xe/JkZZyOcLEvnXFM+9Amo9pS+
aGp4TRJmBaNae2ai9Z2rodzN8GnVnjzoWWW1BChsGBlKox6MjyrqZqW1An+ltv6q3v48Yjhdzogs
GxMOhkz52TpThU7cU1kQ13OhrF8/16CSV3hK7+Y0kvnTLFiii2GeCA6VtP5aRwyP3WkLFKEnxDpJ
1lvi3s0RRW+ErOCVAo0Kp9Cm95L3B6tP2doHesQbWRKbx/PvNJoUW9N/ZgqE8ypfwsqv0wedltRp
VmRHvzZAxA3zILPexm5ZEYLegxGRW03gkQtPKoiS3Gu80bIc8n4RZUA/M1OEZpaT8EL63oxad7ZT
gLjCCEwdMr9m3643lMRWgLVlhf6S7DF5l8NcYxqcrDWFew7IItVgVKWWdxSmZAiitaZgvVwtmWGI
5nqpZXurANfH/CDDC7Rjv4it6cydD3dY7iygPRrI358T5mwOGJ8szj2RRIHgbNOY2qjfBPLiVMrG
z9KPi9L51Tw7TzUNutYy4ztKaiKcxvFxnErdJQO2oHQwX3wePAHsyFw+49VLv0uQtfSAEkuhJvKK
Out/EMRHkF9f15WoBDzbTrTwcto758RsH0TkS0TuPQOQy7/SsZxG/ZkzcNCPBPgc2SeU094Ky11V
BX9kYOyYMvQKih2LwBKz7Y249taZQIWGcqPlC65Qp8ulscHyMLnszJjvTWziU8X0rHF/kLufvETU
VJBBuTMihvoNEh8WyKA29Ue3TkyITvJDHkDr3e45shE5NaSiqLExh2kH3BOXiuS0OFpUwOAfibD0
ZhmjDWz/p99UdsG4qXhuKKE2UwhUUu9SJJ3JZ+9C+aKOqnrCr3Orkg7N2eNq1raSWlj3maEwyAaf
razGuLHIKAp/o/uODlyrLVmtJmf5Zh6p17xPwlNcx1ExOxO10JTB52jT4Mm+2WiwBdiFGtfWk+TF
FxQSlCFgUDTWgHk06IfmzpAZImaArvhVcbYg/pWmC3H1V/tHOMo8xRFtJrCt3LUpMboEb6akpPsT
DJJzXvoQFp/GfEdJL1won5Ya8eH82/S3ZPI/2zvjmloSgOcRqIC+34vlnKdmScQlxe311mqdCDrW
J2w8oxJ7ze1peSM5mdxRC7qzCiiyB7g7Zsg8jVFLwD41jdMKNnpzOnsziqR+OZ84jNkxenfZ8p7e
HJIXUVpjaob3f560h3ILfHAqWW7YfyvB2quvKxBCMOu06XLO4/xxXE3joE/hebU3Wnvb24v5TSza
3ETich8jqYAxjGWfdRWSzaQqNiUUIOVScZ33W6L2ALmXfCTdkdhWwfmhP8MGwXeCqxzyu9IjvqBb
0iTjHWmha97qmncMtjOgbgiTuZy3qst5sEnvRe3WlWeIEQx2qIF5DqJXvNpHO0v/CJlksFwsknlJ
6utp0YfjrAt5lM6KnwvyW7zOCM8qogPLQH2VBx35Gfla0Quz71vBw//mhHZO7FQjOkAG98uCMRVY
mL2E4Aw6Yu0/UfHZ0RhZNynkUgUovIjjY/OrG/eeeBGuEKRcxwRGSZQ6k5CVIfANIuFeYsK3A46c
CGhdW8Ltgm2Tt5cMyKbLC9aug0BKV2jZhwOx+aBak8weC9WuUG4ocvXbpQqzvA/g80D8vXSXyp0Q
vRGHtu3Zg28pZlp9cfUJYLJ1EG8ira/PryP0KNpEQGi658gfvDvbqCWIdtPfzT63AlyqS63VUzVb
2dUcPrl5KaRbe/zEeLUJ2kmEzSOTiE8GP/ruBom5zADuDJ+6OfC5PYcS9Vdj4U55DNgtziRIkWDR
y0uX9NeXNsl3dp10y4CQnbb1N8w9gT8iGU0abU9W1XK9UBaKQm7h28NERuONMgip34AqI+63MWZY
4pzZ5X7cyFfzimKObA61Qsxa6fIwDMjwAtyjBIbjcUqAMhVWeX9l5Mya3Lr5btaGmb6KDONWyE2d
50qOe6RGz0Th57kOyNqGomXW8qbI7vtF6whGY0BtjDpgYaPM8+Fe8kL1iZcxb7pI4v01s4Y8eT/Q
+LwAvnldxveDUTw7wnRLmFdXIApDEV3JpVUy57/M2rONQlYqUY01RrXDveaNBr90BOG0GS3Oe/8H
FoPAZS/HqlacoscwvD2lByuRXcFnpYBL74G3A2cKdof9Jq9MyHGWCaej2WnfL/D0x85TTZl9pLKK
MwPlqcdb2EEwb6Akh4ffonDBrTPviiVY6GOKrnf9m59VVdgVeXcMSl+JL/tPdZopImTaa56on7ok
kQdGHbUH7BjL2cd67FQjJe+blOc4BruAwD7lUDAAcYm3KA6kPLTgD97Qfw6ngomKLzgbbxNiDEgw
3SFWAZbi9vRjicq+pLM2Tenyu5sYAB1yZmIBoNdG/cUHS9Jsyp7tHloqF2YqmPA3QPhidsdUTXnu
KrFMo6k9OFjUltYLo1MxNAKmBU7+AxR5vGbFt3UIs9WF1wl4qtjgW8QCXY7CiDQWkbvvFKLi/k6J
0mjTQ3rh+DqmPewt3vEFuBTVr+8MmcDV5erFz8qnGzggF9yOcr6T1HkFQNooTC/hn95A7VF/VYic
IIwD4g6W/49LKok1wPll6GB1vcgoPBLwYDIZHYq5mVnCp7p0djJxJzVhBph9BOTUV4ydMpWP2ak/
QiB0L91qkGu7XoF1SwwuCUkFXfqUfxbNayp8bBQ5HXMJnkbZHvguuHwjSURhdxBXqCBU14PeaIpn
3qT6FjKIqcp5Sc75M9Go8e9iBLgp8ZVvdbW32pz91sH1rgbM2qcye/a7rqH2ecf7fjflhYIMGmKi
ug/3ThvthoUxq4Z07OTM+CHaHALQppC/TjB7c/KUuFm4HzD88JqqIv1pRZ00D7a7+HUGj/uIof6E
ZeCbB/5DPqaQLozLQqIg/CrEQ8ot/R8vwtXmd8EJJEjEdXLf+D+Z7DXwHLKagecg27Sk0gal7s03
OcibZFFHo4fpWR7mGb+FJm6HRyh8LFGNu4gGVDHpx2um/MqG6G9t0UdEA8hy1PhTGPCvxYfjktah
QBh9gmMRzgA5nYOrPdfpzVpXW4Ckj2KWc2NWLEXlRUnRgeJ8MNNLZdpqBfuj/0himowMyWZRl5CW
UsKKdgDK4YhxMfh+xyxL5fkdOOamWg0KvZyd3OIwBTSCylydZhmWSnTrldjKOlsFXfitnDkZy9in
T/b3OL3cZqVNp43QprR1XYcDod3qruSw+ctsxosrjLxkoKfXi9pB/5mzDeNFNRClIVlmIeUhWlKp
o5QdUhB70fzpYWhHXkmTJtfoYqRtTXENhyNpkIa4xOxS+7jpgzjEggv2wYWgO4M25SRvPUdAG0+E
8fKGWJOsLuQFFjahipm2jWts0HElRnpi/mM1VZMHQp0YD8VaVy9lPJkUbmIazANiP7++nMEibLld
Ut62nks//AkYGg0x5zoq03I4NMGa0pIuQ1Pdn1WNbmynuMcWPrOKkR+ue3fVcazj0mDP9nhAsjPj
hsx/QmuI1IH45wqGMRmgDaXqzAinKCC0nAFQKduuF3IXCen7qbyTTZmZs0lBYkuLNMsiDmC7Gz9j
+p6y/A5JYAb6mcysx9qDPRfdiHFo/uVaH8Ao33op1jHDX+Q5dcdqUE2u0SIWHxPjKhQC656Y+Eav
hIbAfZVIQt92FCgboYvc/WmBJneP12GtUlbGWyjQGdj/hsSaUN59a1Msc+76xPaKcYN/FU7Ba+Fo
jXKtt04KMrUi5PdSx/eT3k58NL1je19b50Ue/+o1jN58TqtcqNYzmIKVPNm8utQ6w2KhHDtRF7OU
hxSC19JIT7nVGG45MSKuyHmqLj/iY+L9UEhImfPTg79S3xr7a8C7+FQIcabvFqyvuMzRYKNZI2lg
+wSwuQaQ8r+mTWu6zonzYGfbZvW62JFc8SaMiXhQ15ya3ZvvisxoUEKwqKyXDzcn3PKJqmIxBmIY
UC0aKRxURZPfgdvZ+kD6AjrnuDcNTuLhXlxjH8N+mE03SGU5+DV8d8jCYjclSV+jl/BPuuS9TluT
juA72j0pT/3tZjR/KGhrmVyeex8apbEPg+3Ryl2qcExWDwyo2EvzV7QGROPSsL7I2yO+GWDSH/Ms
xu6h6nch+3rkd3dJN9pYUayStuxTFa2kkxazEctdnky9qmafjXwtpoEcZTrQ47i045w2gznfG1TO
mAMNWx5uKzzT3sukIlNFOB8Il/YIywJNT7l5dX9bBr2xa8zY3u3bh6rpcGwkAajfcvSpqpjx4x2A
igcfA/xng16hskBXsH2ypWoABYnGf8i4GIJwxwcKfqjP+QAegmxLJFBN7mxaLferAN19EpyLQ0iy
tKprwhU+Q9NZeG7E+9j17uK8HKnm1OwduitMgGrwzr0OhKau+BnrXqIUCFycnbxt3V1MbqDo/ex7
wOY+6uh9zeQxK9E0bXBaQKz46qMHeSUl+FrtQPgocACJ0gK8NTQknLgFsRGInCcRH2kYBwx1Z3/Z
5mYu3T19B9WF9VBjMS1ZdGMdXWVbuqa8UZBW6XY/AurjTD6iR61obgK8CwY25Yf0ob0wDjHpLw6z
yQK6lTiNFNq0Ha5dMaHzj/+PtWk3aeXc8MDJLmwbY9AVSbXuGENQeWkYqs5kwdGC/cE0Jvm4Uvf8
5fimyvpGEhGpvKY/7Ax7Gs0qJLAXm132qPb67sf07WvolmgBG6QCpUffJ7TgcFeR7Hz3gMnFBuhG
wpM6C7KDckvp5FnrqUIarkSh3Y7nhdCqrVmn+zt6F7VaHoJt9HEvUWf/rJsRxavxP7NGnS8US7Qm
wBM7Me0EfD4WXKifM87VibjtNulDufHn7soy1q81xeNdev2NT8NCgVlKgk+wxB7YTCddAQx7p3cv
FaHleUEftJ5D1X5Fo/2jRezAnI1dZwLp6F+2+c9ons8bvStWvd3hIXQ7Q0IBruSeCUFQnjkgMQqm
RUo6+oYaBr3vjBgkCRg8B9QYGt/P/hcF4lS0GEMuPtbS4KGAGz0yB1t7s5wH2AgeWtc0J+ZPcOmq
NhieM9Fw5Oz1y2N+RoS/7sD/2Q/6aq7j8iLpvzD3W8bKHvCMqgBUedm4aK2v0sdEB+AZqHsPhuC+
shR6lKmerkrkwQTKESdMvZvZDlTaHwv8ND8hUgjnLE+qitL0KcKfJNfziaukM+YM+zo+k5ASwPRD
QJMUJGmoEfz4316nc5Ag+rteJ6X7hXs1NVQgTH1ydud56WhR01mFWRc2KGWCpiDCsGKFEoZNoQke
RIizxt7ubnOF0N+nb0QqGszK68fYmOaWz+Hp9WKYAs94APhqBnL3mEzE46vtPm4CgtoPdKstjf8A
wZKlorFqyi2K0AKoJ+RY+UQr1ZyPukchWLVD2Jf5AMqDNQFPqq3xZSLm2Z2sOAOv08RChnNTOY5O
oh+Bw7XgeBi5Jk6cGMK8gzZsYib8n3JYojHLCyjxuGg0qrYxyE7AtkL1o55tmiRVmlPlOOqbeaVg
M9etc1hR9ljyqmgoaMB57ieQEnk4BvTyLcWD2TaepI8RIN9fceuu0Z6kKN0QrwCqsh0EJmeVrLq9
8/DYnE1J2WaWE1nDbCDVNlKAQqYV5SXUYekCdUq4lPC3KUQ939k3n497YC3xVmmWD+KAzvxVKo3u
j58H/5NM6QcV3xd0d9F5GHMP5YV9TfaTw7cOlPwpxd/0f+spfFVJ2h+hm/VtIwwJCw8llZULB5Y5
AMc0T1/4oeMykV+pE6lT16FZJZWMED0EuhWqYlCLy4GdKm6XzbKS5qVmvgcooxFnhcCSyx3Dpn9j
CvXMvFutgm+YTk8MgAJ/titiYEvVMzezNw5VcDTW7W9Oqe7o+i58gh1ZB+nwHwf7sT9CQzufJtmH
2h/dh3NuV6+NxlanE32eTPOPzDQ6TFoFnPxjiD7kRR6wlWXljIuBtaLFLpdgKytEnqsUjKFKNGAn
GEJTUQM342DaOHhtNBxBZvTTdtYfQdKOmFLj0iIscwVuNwberw1atdwOuUs6jGPsjDYh7ytvdAD+
OW3qrrdoVhbOwSbr7r+33OOwg/JbrYs11dRJ+b+XRTAaq0rcikf+J6dFVmNYTmGzy73NyOruQJzt
q/6oP0l6CPkH6ccwEGE0H7R9mmIrfvFra6po1NwFUFjYs8/cvq3wBoqoi7q9S3z3aFItOne0r/LA
4R9ozFamaoYvMj3YV9SUWBGsKG7t7Q4Z3RBKApfzznVGWS9r2Dl/3B2piSVxV2UavF4OIApT/ph0
pcKnYhC4ti7+Vs0M5/REkLLuhumqqxJZ1jKitneDxN9SzTqRm6eAIYt2eSdtj7OdLji2VPGoJNRl
+0mWHqv4/q9zDcpWam3S28L9Xr+bsCUo4RVKXxYJmw9mkeQySEP+95QyD7T/CblwBij8mnNN6X5G
G8JdJ5kZ5/O+huL85GxVvM070aMqx7a0IOyePOr+PnXhTAvMXsNbsNtvth2MOOro37WuO8DoKeFa
JHCewfeJwOwoNfk62fzI8w2d6AFlx6dhphZIU1qXN1DhwTjsN/Cs2TYNmGOLdyG4/oGFaS0x9HXG
9DscPbxCH5vllzScI6QfViXaKI67q8ZBn4u3Q4+jWCo2MfBahyw6qfp34YjWOk2h6bw7fuOTyduH
Q4fXxGKs7ewjrUJee7MAAwS68ws2Rc6lJDd5q/YuMiPw0G8zdVCtOtk6bVw8P6gunzjgZyGv4iI0
MUUVqp0/PIDJi4hvPmVA0xVRvxffg07zyK5D7cZx7H6bLFzCKoL1/ETyIFRDjWYXWLRF/QcfOSgj
Y/QSnH9/jSI6AneqF2BBYdnSkPjxOPCQ1GkKkY1GNeT7lqzJEArXv9ZaD2RVEJYb0SKU+86y5b/b
a2BSwpjS6YDglfOEDUxNHDADUuUS3oOPuN+1a+5/svWDImA9r+4Bb6Mz1TKfyfc+aZrRTXNV8CYn
Qxg95oVzTN2EILU3KljGE/3UUhrq/yROmJNYkiDmXBbL/8cq3itVp5Q5r3bTw1zsFQSqULYJnMgS
MbeUn2sdxL9oU1BPoPAAazUd0Wb0IpLr9xShOapPd02pxYXbhqEUo7ZtGKfgBNYlYJoQ8e835TjD
CkrT+BpSzpDoTspIYJRx6ZY+qkD1Iy6PZRm6Ij/G1hodHERvC1sze80DKCBbSWwPEaOtoPU9Xypo
3JBXTZ3YkDJnFRaB1YYHhoLJ5NbAWV9tSfI/CMpRVVvgjOOvJy5fjolrn+rvNn4f3AiJr7yffp2s
NqOKGZLfKYOoSGUP647b/YMcLHh0a6iwkqD9KBWny9jZ8QUSx3Z/NbIx0p1yWIhbkc/xXJchuaUk
k1fBTXOi6zuL568sevos1KrLm2PQCmY/aR2jdArkWgH7pIiltwRfGtErRBj5A6msZ+pt4Q4KLh+c
BH5RntJgQI5lwF1DVxqDa8tLrKxRTtTDccPmG6InMhuT7mvMenqQNEPMhe2l0TgTPg6qvxT7B1/Q
+wTGFiKTX7Qs8mE4+hH5yRoH0kIsuTuMr3WOeaU3C+kSL1F63s/X25K94Pa2hUZe4hjkaK8TGh2+
lm8VhFcvaB0bju73VyKL25yDm7JCzUqXni3l6SOOxqw73+0V9Mn88hwRig1GyTheTp7qwSvMKRAb
sttre6l+tUfg6QUebGnVmH/WzfMEfnZsh+t28jipcqRHNmqs/mO1xSxJH6v6eIIQHw+uCtubNlwx
IMQlztczDqsYMeF7mqOxktWQFf7MMR/MvjUpgveVieTQprhlWu2K/QNorcN0YWAPBADZshkD1Oyz
MDbdwBwQara7+IYUmsk/b66bwG2P5kXcp0a9RzfU3z0DP4aYuum/CQ4shcqkINyJDrO6b1nnggwH
Jtu2fPbkmdmvoL3jTWwqpbegrxjrt+I4hiZwTk9+gQYuJL7xrSkQG+Iyp2maiSd62/zXlywoJVab
PMHR6Tjyzv93zGGuNaaKyF70J8IE81JUgQZkBtRsXMYOI8DzjiWuyfz3wfdgudIGSQsHjukyyRHA
FxTU5sBKuFOx2Sj863yxCiKmHnjiUx2nOskWdOVjnwRVfLIUIuKiSmp1eF37JMhJ8fPm4xeb3sLI
kUJk+LHZdejaIrmlizChkCxXeVWXUHZksOZTzbiNP9RHXnucJBHCrVtjvPAuiDnZYdlt1CpgEFpz
LQst0IsgnJXw14aYWAIcximxyuCxsGEOnwP2I3YIOJQdhK+FVCQJxc3rQYw7u6fXaNHARKkwDS+8
+9saXv5mYznetFsWZvoB01oWc3VZBPyamFnrRM/bHksHTuNYPE/E55SWaTqzIu/WLfWurjZvR/Ij
eaw0isQ6AII4/spPGkqzn956O9M1P/It4BS9vdLZ/FvrAuPXk22SF+aHwQf7QDENXJwCKZEUZg5x
0zp8URr0dxEFJukLqGVAvrDQhT4tHc2oZHnEUW+aqlo3MdDnASbmA4VKcrtYuTbwG92ZiW9J//LD
XOvypTJOFGtMJV97SDuRQI9bnSQfS8KEAS8scP0hD0M2AZH/5UTaQugknSYlE71w9duGg/p0F0Uh
SCZ8+UElUTHBB5RNOpJEq5oRMcyND9jfAgM9wLpKZ3zHZ9C1q4BtL/OlSJ+u8D2Rl/IFwlZzgrL+
ACBWaL+ADhKvfpzd/1ZxO41fIs+T9Sm074kro5W/yKJh/Wb8Y7OkotPiJ1rLfXzWNbFGlHirn2xx
PIxlhLjfu8gb6qiO4wiowMB++B35wk/Do7qxYiL7SgEILply4Odmvf/N8ZKoMFTzjx2inUafiZDG
CuPYcj6uJAStBWDTed7L2Q8n+m4ReWk1m+I2DGWZ6ipknmsZL9g9AD0H1qrX5/Yw/oS9pHePYfrg
f2/NzPAJnIHR2LFMZ+85fBEGkNTd3qxMDyMr4FZ1Esjm6pJqU59A/B+auwOVezYi3EmyiAOiSRvB
1B/zawXUrGyvRVXtjSvFX6THrINfn8Gl0m+T4hco4Ivg+y62+SyaBXZdw4SYCpsmMbtfjqjqoi2P
5T9ZejrlXnGXhFxEOFPMPAr9I+v5n9eXsoWqkPlyQO3lhfTCOJuuU5yd/0erqXVUYSbwAhWlrWq0
POQFB5rlDYpnGC8e2aTpKh0KeQS7Q4UV1GBgcjyjmOv4XeVZ4x87NhCzg4bdjRwEM5ZHXDHSx3dZ
a+7lbEHfx98+5h1gXIffQF6if8CExkjMmvA0PQgzJicCVMzqaG7KrGC0FXdymYYojybSc/szqVAD
Bweg2yVs44v6l5lLSS+85FMasNDOIf6zSNFId/TRH1y+tlCnqlwRMxnO9qkcI3gVOVMeAmAqmRDR
58FvpgGQfPfq5s4HplsJHd+/wOqOYjMzcSw2bwRTIxoN7IXw0FXjBKFCMyrGvS/UDf2MwCYVCZhM
xT9x7+8NdURIGlrGpfo4qZ+ttmhCr3zhMBXzoiiXFuTmPkceNMpvkACRyapFgDwTLNyfC22p1eOh
DFjxTxjIqohZeQ6JCxF5ZuvOCrf3NgnpztN+SeeBOme6tEBRz500+YNQ3PVEygzi/yqSDDkGztTd
2A72F0I6P0JKKz6nkuMeqDMqSLYBmwKm15fJDg2neuS/+56O/2tj01X5M05c+he/gIwqEV9L9Zqd
R71asOxnbVcRvsnxuhQagR1tqhkEGF1lw+RhCdXOudsrRfILIgkqqBlcCFs8uFBj3VyW9H9ojPUP
0hfqBEVOJNYavticByX8+ulvot/a0X/QkLPzI9N94M1Sl1MX+6L7WCcq13aCKsWuCxWbs3I/tfxn
gs4cixF0HNRYSLahCOh12/donepxMPXynTXddnHicQ6VV8EXVCEL3k6YqWQyOtvObtqMDA4PR8p3
S93glaQwrfSSyKghyqf/9Ms58a6qeX5Xa28sz1OdyBDt+VXt1jXu1OU0resZJMB1NqhI4fuaFXfu
38ylX4O7NL3rIiJA1yeexBsufVqvGya9yySNSmKYMqYQ+ADgggcXJwSbchPS93cmABW9mnQ30gCB
uNnRYhMKKIpbFpU9OiPySX2ak86vEDb4HKxuf+sDNZkrrc5JmJaTf8foYQlqHkvdBcp7YA2esQOm
HVo7MdKqGinUbwsjkke46k6sHONOtB4yDTleI1thRZnnWne5HIRkfF2kcG4zhPJMNYMYsJGQAUYN
Gj70FIFWl+AVbXNbRjK6uMFXYAr5e2byUWzIts9wvuyNG/qSE4pmNTcZZMYWb/WNrybKqjAnmTjo
WV2bFmjQs9C3s7Ipa+qu3dlw4YgyhN4vMim/jntiq5XNOvj3mtczEWQqwhmh4NkXANu1v7A/Eq6v
/rMfmxasaqczKw3AJOZq8kcxENAzynZLzJdxBwHT16C7fPVS9B05kNw8Su5wJuEcfHSs30AQNpBg
ghOrydvYcg57iP1OfbZDvXMFVl1mkJrgAhUZwTteiRQgQ0rvaKZxMO3D9wydZQ1mPK7v8/WhBIXP
XQ0j3mXc6TfaiYLJn2+i5E5v4B85XWnhHJwxK+nV
`protect end_protected
