--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   duplicate
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
PNkgre6g/yT0wQD8GrDH2xilzn9jnE0e5QtUArlZI1QLaRWHpQUcTy+RH2x+tUZ511x1P/D1fSmE
zjo1QVHao6DHtTmz/pFWFBH+BA8qgf5jRR0vB0K78RFgRpPmXYSV9I8fOKIXr+0TQ4ZSYd7Ke/Fy
GGPUOFRV+up0T59nyGQGIbtTZ0HMNYaqhsXI1egEaeFxjvFrrJGwBG3hatMhzmmgKUiNHuSN05uR
oK1jYs21iyO7gqLDN+LBEFPlzaOko+s9oTegtVKoXWmiTJYEvWR5rDnqN+1wOEV4Jvjd+mkITaaw
IXs4ao3+xHGkjt7aD096Mbdb7TeNfG57Ql08jQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="HM/Hnf8dy6maypb4BI1ZWFZScjp2mL/+Ujv82TQ+kzQ="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
IT2ZIQQn3x4dHYdMECAI56oALP/YHY1uPbf9OBwkPgl7LAg10z+AEqUUzPfyyZGWiR7ANIaz86fE
2xSLTG7H/kFVbAdpVsRjLPIM8WUmX/RBNFE03qxtP2IGf1lrdFoxZpzxJ3E5mdWFnP3madYlsB3q
Y4MmaabZ8860BNPk80fnOjMdK5ATSV753rqEAfUg0TyVpzV58U/NQxOGgm3SwGzFQXBtulWIwhWi
XOkQAKErgIP765FOVXlXGB5syuPoLY9Ou89Jh4/YAFgrSsDjvOGnAuV99spiL0h4unBO0E3gXpzX
lr5jHCKdgtK2B5Ef2c7YM45EoOL4q3zu3Ecf+g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="MkOnvkWRUm4pm90e5SquSuJSGhxboSR71MDQeHvfUgc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22704)
`protect data_block
iqwT+4KZyh+nFWfag0B3plkMxzJ1SIaQK6hmZlOhS7C3gMbX2Ta4vAkSHshep0MOsalgm+wQSFek
bTm1WLfjFpTIV9BZdro/787tTQPyeZLfSXT2DViWSjRCbIrmviF8xTlTdI1P4H1WHVpgnbZAhehj
KXMYF3ZIo6/BE9a1Tgxh7sB4tfnBYAcHEZnyyOk4IyU9H03x2RgW4HIU2Qvo7y/bnh8z4r/zDi1B
HUcQOXoWZl/buE5EMHMzq6arUYWPpDDiz0dBIE5hoRd2qNR0MrutKHAvqXrMbSW/MMzDJS5EJKcU
25xFl76xW5ls/Y3dhb7mpfL9E/WJsdGpATshjq0ma/+IwmLhf8IEfml+9G+yH9h74W6HaBJrR7as
EqARXa7l9lEMD91h/PNVvgeY5pxsrc9UrDCH/8sCmT9vD+3ak6t54NqNwkl30cohfGlp3CUj29mG
O926Xxu14wpcrG4IIMTbfrAXddGqsMiffq2HsC5a3jJFuvFzdwaUd+OiOEBMdguB1ZZCIRb99Z3e
8HAv+RvvxzisXcFZ4o8wwm5giuopezGORe0JjeF65PoT1rPN01Xv27+l822UK749WSExx+olCjTG
v+72n2UPWEiTPA2K98Bb1ynEFMvu3vljOFEej3QtogrjWmnS0KwjhXT3zfq50o2F/BP80Ll0DSNj
b0tUSP44OySw5/jzUhW51I1hdXS3HBbQIPiBHtl6M/dO2f4BiwrxguVxWF1cwuBJBOFxPD+yiuid
8teq2LbhspHxcImjiIVNgkZ/s0/zPoVJFFIFyjel4D2TS40fBpW9SunqEv9/of5gcUco0mN9J6+H
c3krT7MeHgIpocLmHNbqOw700hbix9JmNLuov7sJpFZ/vfj3aikZf5vm4xvf5ea8Y2WwZCLOBlPA
4h5RlAJWJsrsuyLY9hsvE9DFxCf8Lz6zETHqeORZB2taMIg+Gj8tnEJsaZjKC+tCfoErRqDdC1tK
Jz22tDd8+q3C92xsdv7V2SaFfiYZqX0GD9UYH8QUJlvh/2XAe6iaBd38LrBCte3lWGl5Bwuxb7le
ybjZL/VDx97jeTC1fO6hu8g1rxzJPZulJ1A5drUzsHVsPJrz8HgfLACFdds9JSvdeIs1imjHVtuC
Lmni1cIsEutweN7JpczLAAdySQOhhAbxJTqolQR8rpAiac2Taz5WRAELB1VwwIri28gBfGj7Jxp+
JU3z8w0xzIC2wJR0jf6OIV80/kPlHmBZQzO3X2yiCQ2RTSEn14SAc83YHdKKn2anz1Hajn1TViD4
d0tStmmSA3U4ZreDlv7frwYviMoTvSSWcjEyOpmQJisMVZJYMvYWI/1cgEY7YyxL3g2GcgPNz4Cl
AdAliKLvJBhKgMbFBjMxQFbVkXGbOuF/V1hCLUUasCOe7aHn+wg7cWYinV3aq5KzUeU28ebs5jiD
2H+dPi71faAdKzdYdMlds+dYbEomjSKuC2kDmCeQYz9OFiOlGVcP9Ou0poVhwuPEEYiXM64U0fzQ
GH5XuunViYJwwUWy1Fv+FOx6uQLhwJiOQS8r1L5QldgFhdRFGT+GQGw0w1poBMiKTotOcB6rQoSA
61Uz8SVi9PtFOC7sSGpe5E7iEpKKWfQcTRkd+LTUK6/BKvn3vFPtNZZwKLGFgaTwuhFrRNnyPuSD
ydq4e4iKdoDOolxgKUnAIDYbFlVdVmCi43YSlEPnPwkMqlX2xOr3j0BC6Jw228lAcSxvtIZ3Puy1
WrVJb7TOwgL0or4G1HlOqOXTp62nV3qQfbsJlFVZd7av4V4AD4dvXHYOjWN9WV/+oGI1KozQOFIx
e50NF4EQtwFWUghichZc/BqwvShIyK4jV50nKrHBdby8dlaW2Dl2TIEWn/1CnI64cn8fbRtW2mkj
9m04o2ljzFNl3iIXlhbSPY3gBv4x3HTl5RQ3497XfmbihrkISOPJHZJtkCISdec4ZZNG5UERXXie
ix5v6E1Ofr13FVmBtNihbT0gciOO9uPF3r3Waz1848AjOF7/dKcwmoPp/SibAg4wXzorippJmvs5
oAc84WbAwV+z+jShh6u+7LibvcFXPhBdGuDF9V5hgTPxMimscHp2n9Sb6fi3hzpU6PLaSpdEGkVq
FUFfJdRTjw7FGwE8Tx98nhsukvQx46DKLpr4PCEyelmuDUB80SX6LB0bkE3Mw1pLp+rgPNMvF+uj
CKYjVo7jr+jDYLaSc+dVqk6UY4erZp8WlSbno1nCMzNBq7BkPkctFc9whu5PQwmRKjRD4dQMTz8S
ZXBsIaHHoJNoAjrkK3VMb55lmTw0LcLq7e2+go1vYGvcg04GWehJgHAYYop9uS1R2X/sN8qlT71A
ts5mtOGd2ozAYf7WIwODSqVVkt8EmESFE7vUM0aVGDaqojQmBoPkgG8rgdySp9TRA3IK3uYwy7wD
ecRqO3xG6CgWcaHwvpdwFlEiNKplq7Gxam3saxvuBYQDJJJ1LQpgoYzVww8WnCW3lbbMNbGU0quo
g0uQMkJYoY4RYYfel8dhX0S2I4BJLnaR75wSS4ntGl0/iiqfJitH6PD8rBkO3WArKiIQvtawkKI9
mFOriJge50GnZv0rZ1RTmHVlP+VzinkAeX3BUSXMp/wOK+f5YC7r+/rcMxZejuPTquJVU25AEghT
nxU3tqWnr64Fy7xBBnhPcArsWCbNiXiWLny/7D9wdRUW/+XTI3ZVTTZ4/Qyic4Pe2WcjoMRSVz7m
wfNd4UKrNxs5RK3kL8XaOl/8ELFzQyhA/K2Xm2sC0f1/7+9KlBYUfJ+EXzI3TWESW25KZ1+8ME/7
0r6eOhf9tz7DF+AsVzT9pNe9xKBMwu4qrC9pNRebXGIz4x/j0JwYsM8oDgsBSV8nviZc4mnn5O2B
0n3r8/LNNvLrWnOV2S9etp64mWo9TkeZ0QejXogLV20DAoa+24PFEax/2taHJWqpGQVCgM0thBdw
AWBooVIhaX8h4xDXzf+xdxbDLjfj6Vxrii0XFvrvFmgZ7LKWRNtZkCyGfxAf0+M59bsbAecavSVL
Wo4KTETqoNz7d5tzBKHonsECfetWH0Xz6gfAUWWB1NqRNdjfSgqKcab1us7Y8JD2nIY35lLRzurF
026h8vAh00H824tQlxiFtQfYIeMjNS2hRBrA7k7043OBrqp7/585V3MFx6zSSlYQce6l0+3nBFIv
nIf0YfF4OdF7PSl786zAmmenf7+ef9old54OBFgDnHgljaASkvbnfI2mm4yiCXTw/A1kOaoCki5o
e5bwubYGN6vp3iashphyI6GxiEn3bAJjQEi4de1ocLoRwv4KD31etpi0mopmeYXagwnZYSUyLJhL
HCxeDyyd4jBYbpUJVIYTqathOFCAI1SXjVaA0+naC5ZYjoodzZ6XTB1/Uv3dli6cbAEuZU6np+ma
TZIijamu9nCWl3DwyPClhkoat4ddE0MeBsKbrp4m+YvTmeIaYqXJzfXxlP2/1r5b/MAtcxjJCTtY
sQlAs86c1koFUYaeM5LQx+TJraVQtuVdlorka2jc6T4Id4RskL+DmCE+JudROjAcV0ns8DusHS36
K6hLgdhtxyHpF5ymwlcED9OjnMBO3ZxSUU3yddQRQ5NXhPpIux3hVGNpR/t5GSGoQQAnZrF//eWI
Y7xGk5JpuU+iGbCLIJA6lsuz+1vi35WFjj/W/lAJEGtdr2yy4HhkZveCvOaPddWrdoYDEj3foJJI
mjZJWulyIAdzkANa8ko2nC6N98YHXumDdnJBwyUmCp2L7Z58XkxdYAh7qLqb7NVb7FqCuDjT6SqH
+ho38wxk+aVR1exfG0eXYLEml0ZoQRwEzgwRD9BzvA6NqMxM7DdsrFzO2j9KXFnfZF3T9KzbocP/
eOxGLX7vXt420akLj7IykccJz8R+7w4IW4Gg36CAWJKq+PRfXCbZU0m61a79ef4ezwxyDkm5Yy4t
XkzTQQTmGgEaZqZ3dWFTWx3MX+ZAQ+ts/B6w+y5e0QI2kg32RvdUKXNZ2hkgZJ8HGuxWnTKEVpEI
VFcNFJrhfIRf52iBSwGKbDktBADgg4ECJKrPSKfPdrZEH50SQGAnkgJ6WkNTxclJ26m2yfTu8/vM
pcgzhL3le/MR9VcbYIC510hP+uisOh+kH19iv2ddXzGiQPcT7QlDjq2/dptVFlODHYwcW6ipLbJs
FoIF+cJcnP66rZbmSZQwUFGBwkuxZR1DXackcAviqWKXE3fppvIw0e/gE40IHlZvMIcBUO4UYDof
May1mntT4sm2PfHTyHYCtdwKGy3c4Z8Dvyes+5aa6zkBKs6Bp9tBfYbaTf0af2Vycii11P4XjSE/
QuagowRVck2HDlwJrbWeXmsGTvwABk4K6dpMg/LO+T3dwKGLWcDaMSzpliQbiq6j+LJBlQIfN0V3
F1B5ZwGumivsIiqdP0sFUSt8ha0QnHniq7qK93o08qmDm3tAN8jgE71NGwfyhmmabpRue2vbPyKz
mTWJ4NQ4QePf3iSqcPmyRGLCLxRrk4KX/C0Ny/dyjYBQt9tyJ2PRF6Pn/FD8HNfRVz1qHr7cXLNB
6xKDz4IadVncBgIugtW5hAn+JOrJ3EbUFy+eZJNnvMpofseGN7/g91PNMoKPU8qHyA8el97BVdNj
Idik8X3nplm0AsOXpkraC/hvVs29NhU1LxOZ0DKBva8OotWSpp7MrFPNP2Bo1WLdX3JzQ4AKN89U
XhUd93gitownOXssQ69twPZ1I5VerAQ6XHRat04ncHK56WzAYbDbVP5KH6k7ayHLBUZLN6H3xM1K
W6cs64B9rnXBY48ZgSXxIQFarRYAGj/xhze+MaSth/slwjGpuv25tGkdxyNASVcpCK88cUUXl/r2
d8x8su7d9d5lysgiPzMcGd/y+d57xZ+WEbx0+WcNAaW1YEjhb0cFAeDZaHvTnJv6cPBwpEWheIVn
7vW9h6ZLylYo8WJR4YV+j3vTgyZ5RjAFKGUZaBtzRF5lplLhstg5KXFoKNSTelP4j1DH68O0sUtd
q6NAzvbB5UEwOPb5R8jHz6kinsWQ9RNFQ1KWgaUfx3KWiHspDYdCQ6sa/NYrXU1GVE/oIqvGo5L+
8VcIDYUpTF7ffpZ9iJh7vnYFQImxVNDLGtAvThhK9h0IB3GPIdaK1l2Gf7InGvZjmWFDeV0icadr
LNIOv8yoxuQbB8XvVQPqWKA845Aox7Dm7DORs0ltvfwpDZJMe3b/5zfiX1hEa0n6w4VUfHCZt5XV
9K946lVXIjOR40WAZRHCb63kb6JGW2PBtlKSPFXS2nkhFe7ebGY5dz7/00zra7MZAaHdGs/a3usM
dBgKD+3/3XjmL4fDg5e63lFYoVmskKCANc8DBhXwU9jWoJnAt0lEZnl34KduNyV8ZL4nMzoCOrKZ
V3IkTZIUqear5fLWjYzer8tasp2DMWVd4KYordz0iPTfOYi8rhhZGYghV7AKd6Yt7ePbOF99MwbY
SAaxo5Q02bXSrUlvahKoPp3A5TiHLS3WMBfZraiPllGvyKBNhBim0oW5sdiwZyZIijFRFVcKgO8a
ztO7Z2aaXixjPCtyZp/SQCxbRvGBgRSsmuXBL3GsteLjchR3EbHi95sLyt075GDt+8mBDZMPUahv
AZUrl1Ng4c0THdBr0UVkLTrROf7YSOthJul5dMiX1VI/d9CkqJr1o24D10ZimjVMCsXqmktS+1Vo
AHPE/HlBVfT4mh7Sjlkjl1FdRyx5Vm8dm9DnzLVaRsfxT0n4NMYS1X90EsCqVOU8My13JJXg8HOZ
i/i6N9vgB7lVfN5V0VxlWGgY0WxvN2ZWb5aZkPoj9rXENZCX6ZVp9wQrmPysXTsMfVcU6oW6LLhp
Ei3G9XxHAZOs7I/c3O2P0HaP9yU48fcNLc92tvrpSwFfS9GKEOxTF6ADHcZOC2GY1xn+rgUNeqKK
q1xhHuBdCFAmFoeMrlgwQybwEnt4urJFWOzDpOTEn5naOobKq3E5JhsqZpfjIj9UDFFxm4vcdi8f
rFKkpEvR8Z1d1kV1waul3GlP2BBHA79sE2eFXoNvTRF8dSemNzDb+OdcrDJxWBCb30Diyym//eid
Jm5ufwfDanH4/4Ugnjie4WHLtRvBbcRdtFnaHcBoNdXqQXdPVHjpjKAyKaEMmvDwGGhm1UpiM8SL
mfZwQfpafHbxvG1meCDezjObSw+3rhoKkM2GJ84VeNFHnetXggjmushTZ+cU9bvOuy86VUm7GCb5
DdU1IOOL4mCYqYM13Q27w6guK4c3uqYVHzmRjtV574kwiM1K5NTL0Fh5GsHMAg/9eiLxPhRl7dV4
nC7sI2glpwIghDZXDOzPiphOX2hr5pn2FaLRochPjssMPBzR6CsPpYtWWpJELyrDxQ1b6nfalvlz
zyOgf9Gv8uYe/bAz7FaEIw56NNhijev+oeNvYZ+rsWFrClLndnznMTJaJJp6gQ4/VMjShqPsNc0o
5zhQ/ugQeyhpkDyqp7IE+g8jI6YvqLzcpgxsOHWjQliKXHxqlUj2HmIQL4yI6KmssKocGuDXGptc
yEnrjpx7DJX2QFnybhWJuFXdC4AHV1oene+p/prp/LFH47yERFDkd4GMYeEVfCVtXEEsMrHWeujq
mVwke2POoEghTvc4RK5DbzL/0MEpiFN9iVnPsZs/joqB4W5d16XZLOLU4X60SlriG8qGTft4C9Bl
7WgeZAk9YNi08gihYULCsnGn9kufvt87sVkAgcUYVQwEJ0wI0ufzRn1WINKX9XVpngVXqd5PVsyR
ky/Duui25H+ZugshhLGtd1U24wftWoeC+hOtsHxhKtdo7tT+0RRCcQ/5s4j8KsTKyuQX37Am0P8/
slDPId4eXOg+kLq5w53CBc/Hh1Er46mtxAZ3DSBDGPYvxpNWFjmMJxDLXFmAq/ZFcUIBxEXeGo3B
vbQjJOdXRRGHi2cTGH79pXwnMwho/lMc1i8p63d7+v0De3MrmSCZLllrVpD1JbbrYQ87idQk9Ueh
kz4mzbNbwnrt3Y01ToD5O19NmPv5VNJTndeTGsAClvFVdBlJQJJcAGxRhIng9xhM6DjAynX+3zla
BGyIJyw0fTzvY7YcJD9OwFkUcqyA70UiAbZutjazr7ztobwheCzj8103pketCYTsH5cTt8aBN/Cf
z8GGShXvFeLpL1rHC/OdQ5BWbwVlZ+yubK+mPz4WSYQmVwjqg2ak4JjZwAyyik+a7dQBAMWZ5w+y
SGUyopi6Xp8mhjrfz5i0TxWuBsAvhjqewxIUe3OeSNJnsOHCj2GrEV/Ns5Ay1O+fnQw7nGulSoKz
qaAB0TGqX99nHCLzkzxAG/snfDfAov7SxVqwQeZE/GaW+FaE6Az9TqdL6CRmJnDIuyx4gcyaaQe9
IyvkaOpS7hgK9lQIb7fgNqdssFNYHUdct5wzdXTU0X/P+kK5WQCZTp/bvb0DgN+9hWeWuouiZMPA
GgBbrSImyU1VaO+tVgL7QCePOQsWfK0Hn4SmbS7dRoM6cE7xrPtNBVjjyqrIAVSTPx7uDNr1lEut
QTFe16BDzc5Dv0AmMwBCCxzHCHFTclgDfhBOoBEg235fqwC/zh1vAggt7GUIQUiv+vvkyQs78uuF
Iw2VhEMJ2Tl7MNRz9xa/o6quMVp4hiL6MnpkQMTxuvNHqUv5/QwVyIBW4v564iL168dlAJ4no/Ln
PTDiPwF/qOix4okiw4v13ejnjM7WiQlVjCL+26MS+FHQv03rOK8nHpTVU9OaU4GmxoqtXUFhqvKD
tB+pz8h3WyQzKDktGfvBHZxXgvRdal6mWysArUI3aQeRldoU1hVF0e+VUmcj/RKQQOITLUB8qGOo
4Ofdxf/35zeZdLBtBoBjMvXWihFwxTzamso69/CHDDGPFv9OjLx7u2dIU4z5ki7+cOaatQ5SHLs1
eCsTw8QbYi9O3nW0dcLhRFcgefDt99EHcP9eBSWw9G/cN1+YfY8JNqZs5wcpUkJK13lcMbbIgIw2
EzZACXIqnYkHL6JppU7v5yLcql6nba1sKhz66hk/gMhRqEXIByylkeoT79pm2f6ys6adRP6lY6vH
NhTrpRyscOaBo+/oyLAjDOXnpBI213VW20viX1/are1FgsHlMvYFmiyYDwsVETdxkvkzT18YtYAk
n1x+jLKhhTG/Ct3brfOruzFweddHMAxK82q17tSurWnWxn4GsrQYa3SJj2/8lblHLvF6LbcVM6xz
et99EuRr5J0+w/HPlbKLgOCzWb6gEEjn2tQoDYbvi2XN9tNVtU/xhSqPDWhcFSspiFyjkaaI0F4m
Wsv/BIMnXV+jfV7N8IOfp3nvXLMKWwrZAkIukzczVukJi7sqGflBIrVTG8s+GTXQ7BgrulJKFYnV
p4nKnBmC1svz5DTerz558UG1ME2rPteyXLQDfV6iTNjHkptsiq2NvUMElPsSNjMe9s/8DP9KbK6V
GXIIEmpY11EQCo9krrXvxQU1YPHgaVUF8ZI+JFDw45ECRH9Cx2a4Pf50v3xjcc8g4uelWwPkC0uX
Tnqa76L92uSzUGCrhfGykpet0RZ1v4HZY+ZxKI3fPqmXuLuhjCP+Lz+os084SE6p5aW5iGsQc1R5
n0Qa87jgu6KvfmaeZ/tgqMSh7IkUtR7aUSK4yuuRxFWJ1wWetMO2Y/FqDQ2hE4pWn1r8ynihSN7s
BEefITEKTSLrVcetYAOjpmUDppq7bIEWX17iISVNOIkTOyUv52HkLXk7DJzh0dNOBzNtSuEEYKTZ
rMoN8bTF3NopA0uWDuLKdgZwtR1g7b7OpLPFrb95JQdiEabmMHHZ1izpBtQyNYieF17b9kSt2ep4
B3jYWp0BuBJxY3WiHr+stauNPnL4zK4s5hSNjwKXtqSP/wLTyB+gzZeO7xeJx5asyQ6MWs9ot4p+
9f3X37mi9yUXe7gUxChX7NEyeLxsuPxYPutBWMLltzEq+PPAhNM/ma8HP92yHHgSKwzlcGoARwzD
yuXSSYGNtCpOIZS9eIwcPwLHkq9b3bT5IvPawasqju8AwhQ+4G0zDQHM65ImuxguBjp6fsy00fqw
OYgFtVVhpLLJttsRujs97zFqxPOZMhzJV74Td6VDWs8FmrhjMwPK7K5tQmf4Arq2DkmBJs4+Muuk
MQM6vAy3ndMtm/qs5CF5Y90furUJF2YeX+n4kWsiGJ/LCGjih0600fA6QDY8oI9d8OXJGjPg+Az3
6P9XVfQ9eLcX2fHOXpk+FUjgDzaj7k4WJ182itrl4ZgqT8FLUD+E6lbAOk4CfShpzL9z2Fr/K1zZ
v17uvro1gTK+iJkk0Am0j76cWDrTYafded+wmOpeJH8S4HklZ04gIsL8pnC0kD5l/kTl79nDKzyJ
oJPr2lZg9tZQU9OKMvp0w0EJGK9/D+LS4aLmHtztx90KR1rKrx+orm5rLgPVCazPd8uI3bm/IGEe
s240PVZ+cGhNPsQaE+jwS6SJmVRbzS3LBG1/QE+BeqfWyk63gar4VeKHEmvVLztZId+ywpXNT+KP
61yH//V8h8uMBOkDj1fLwkEHhHnSncFLfYZETdBaM5qI52wFLZnZQlwVynotmn4Lh5qOwRrDlyhB
v8xQsNMQ0oeL3Sv4cYfbxD/YSCEdQyIPx+vgAva7gdnYzy5TMzX5nFb1//Klsw3yLhhQxRwaAVTK
UKHoO2BsunBrIRpUQ0+Sg9DWRYhRnFtO0niXjsYEGEZ/5UV9tTA+kegdRiV03UlAsanKAcM1q2zU
nenVQn+w1VRKE6uPOOAjX8pDF74sU7dNwUpIJBnKgqmdZ9AEVvTliyHFQ63K6QzyFacbu5PxtU8L
LKM+gmwZe6KUkhrbcsLANcmGRdguJ5030egFn+xklS3csOa+IY6vdgEDZGDv8aLOYnOzNoffDnRw
zgiilHvX1Jtlq098nT//aFC6Jvd5XVwrSP7zDr7o/3YWyBTiQKJ7pqC36NPWFKQvik6tUoDgbQGu
sljmwo5WQCBgKQXE0s6+0b1zdqCqP+PlfBiaUQhimfYlBHkb6t/+IjOnHyCBhO9zuwtQKZv4djyY
zSTeMymRdFAKR+55hmk1xtwM40uDidg2ZEhHwQKXzNWNYlEt5VLoEjDS8EmrUcz+SN8l/0QHy/Ud
W0nrOi6NnM6bebtY6xsl2TjCJ2aEFtLDrdDM05lvXZnD3C9/qG0PcgqkQbQXt7CLxHBMw6Vfjn6s
HZMXsf1x18vu0A3tiqa4bbKhLghH3b1wDC5FOXPE3tz7LjGEbIjrPoZnFNQbV+a+LcFUhr+f3rvF
/85vwkuJrM5fxtqsZU+5zupZd8GZHkR4UejztE87EJr+o+WFM7B7sK3KGeMOoJARu5AufP8r8sGO
x6d0S4G56U1DLBFXIKwN1SC0Pd6o5BDND07vml+51C1EpaoWkA4baIcmIQoyqalhXnQ3+c3ayfpi
4UShqtpZSyurEn5vWIC2ZKl3+mW0SRD4nDCaggu2UtSEATXZuSC5mLZVgUZNHwShl/tp/N9ORqlH
+lPJBjnnT1ckQ2xa/aDN3kkmwWmgrDy+64YAL0Ep7IEWw9grheCZ5vzb4d7MOmeCif9qnkeC5sFg
aY9oEpyi0ncgYHiHR5iAr/qQvXrkSoUTOkRGuA6/8pBVp+th2SsruKYPF54/B0SqHe20Inhgw0YM
vDGIU8sAVTmfTNMu2IdTQ2VSoWlWO46w/O4kJRE+zdt4F7skydI1Y5Zx0A+GZiMDFVwqzupcSr2I
xSHloSOOYSV8M0eqRDBCUcusT8AkXoKNECHZZU4kEkLA/siSr2oe7iLP/XEfK0LCbx/oNAi/XbQe
qIbqRCgyji7qoJviSi0gLMRhkAEztEg3AIxI/P5xRDcOTcVZ57gVVyBlGiJUGQTCuMcRHlZ5vIUN
R+0jSx+xVJvO7+anjebzwk3AHy8gYRQo/PUjs3IypQYw0HoXiLOuI+WVht/NDpOd1yy8tTAVO7Tt
Sqnky9RyQ/TPOzXLo5IxHkBhs6MbBxHFUpwGp0P2l+djY+JUsq6YfIPkg9Q6jMJOSMpYDbtTgwxD
TpFiO/lg4+IPfmFzmAv3fbCGv6qDS5RX7yFN8cHy+Ct0j27X2nGlJ0kLpwzkzBQ/raQvV3hUVsYU
Jg1YkGEFBHNfqWvmKQ1QslyufcOb0KWIvFO1KAyQm3yi5VP0CyFIdHOKvFzy3R2xqPs+h1B3raIg
om28ddPUsTn8VVzxAaehaSUPt2iuPd7WYs/B296gXIuoFlqjqGJpDrnHF4VNbRZxbr9FL6+KePiB
PbCmSKUO46M5itPnXzMoaxlTw0ARGcU5y/hwnPwsqaq8jwbAuUqbI+47YHha6jZxpOQe5hICW4KS
7eAF2EysRBycGbzsT74aq52ojZQ5Wf/D8FqNb679/FJPoHcJ9qEyOGt+1pJl3cNzqomaIfrxkDWw
tlsJ11h5C48b9bWU+Gm60r9CLcKhPulnefs0JH+oaAtpPUZdEV0ubAu561XDMTUGjBwaLI392dd3
S4IWSYSJTrWgyJEQthEBlBUQq8jJUz4EEvgBFmbWeHfuWLiqH3SHFJrMrkIiKDFTfbmVdG79qHY8
4nLyA/oyki4S1ukU2GcJcPvfH1/Faa7XeheMjJAZ7v6iVL9xJ//L6CshqdTdOq/CAqvnuX/YS3qB
SqIQKSJAtamuVUWrFuEsCRgnvqLL41bKo+whRm1V/UyPPLT+qpRJCKFtSuHq5u/zCeGkTkuHKZYq
B0rITuHbgOd0dlOf2OPeMgESvVJionWTPvGGn/qqd3IrdlR6MhIY1ZdKU7xDRzrwlyTTGy9FgoJD
RPTe1npZ1MooJAveboP/bdZHL4tkwQANGLjaJtWCZcSE14z8+NUW2ymNJ9ybuihqHS97vaDbrzb3
vS0PL76FKgQsPULTC2W3D2ZvK0rLweHDfNl1WJQxBi9X6hgi0NkwqpXlqJdI3jAQE4Ydqn/wcipb
6B18UxkivOzSODwpu60cPkvHmS03xEsKN1iQO1s5+YUh6yyho7RN3C0exvlOIAnQenyeg9f1aj+D
cjdW01k0RYmpar3kUUx9W57k9YGaPBahAdERYpOUlwMs6vl+1HzI9oVHvMD6LWx3QyMRpwuiiaAk
ZPhanvHkk/CFCjwkwR1xdrRFLWyhPrAB8CdW/jboLxWrfQcvv6x1hbvjJ/QwSOzi7GZ7rYTXnQva
3PPRZqXg/TFLBlIg3WZVxXfWo5YvwmNmTMYv40PTrmzaUW7pBwSjDA4Jl2NYzyJ+yD7O3vYnsaX9
jSPOT3I7jTF+Bse+TLqzOhCTiYpAkluSfHCXzeR+tjaw3yWkHtPI53ZAUxT6F1FqapZGkNIVMNz9
4GYGOr4cWOuiIvy91hHJlY965E1kOoYOyjYvaCqnxHq2LsXjL+cHTvRrrfRfcYAV9x3B1aMpK0RH
RFZ1zFr+TULbIsQvfKReBMZdVHbPhFY5tunKXGVLYlqLLnSESi0o04Rjj5VQr3v4LsGjH4UQz6Bp
bq+OG1ZJ+CDbE0DPpW+/npKEjLdnshBlCO49cUq0nBVNwAP7I9r1s6Wx9mQ5mHZbRJTyyZoGRajM
9ZxQIE041uaMyn9qZDzcn5t7uoTVTdVU8c9U2hf3oW4czCStKFBby2+8Toe6MHwrW2kWwzNEu92M
lgGHWVhJLqHsSZJ3f8JyERxUkUMj2okj/q9luZVOzRREmqxLtTqexdxnBwH2OKJ/MeF/GgUEd37I
tT3zqhhdz1kLyZ/7ZPb2dYC3xrYduPC4fStwaEM99Xd+LLdyZJyZpJPCENpdaGVDbDDleP0L3H1i
Fj9QPpWvea64eq3knq8XkCzkyBpYVf/vBEkSt0hIIrfaaGo2X50J77j/4neyWZhsetArD3sD1xEY
P7rqYxAyhtHO6S5KZXYeVLSgFQb1+btSsk7uE/c3ZmrdVbWiE+ID8mmxBpe/nsibaSs/AlmckHfn
ZNqDpUs4Vs6FNecCBrxdXU1zfb+YX5MfPKOgaU9UYIA8+GGCl6q+1JtQ9nq/0PhR6+ItUc+zYasz
O3tubQpHo+DbScmMXZhKq6eYdjyAwkJUbi1aTO1ExnWboAxHiw3i1qUG+73+8slT8aWr8EMGPV6x
LPBlorbysSClD9KiSniNPkmwFZaeltvDsNuxb8NM1w35v4WXPG6j8bXMde46hmlzK9yKjbM18b6A
Bcstuhjs5l/6+3uldpSAxUjOTPG/UmiJk9hJPjThVs0FaJEGM6AYWXFMT+ngodESm58kvLuI7rhT
RHSI/dNqLctltkXMhILRUTKvmynJqu2Sg4Ay0nHg8vqD21mD8SIE97ieYYFvqIaQY2iJ91WG9NDQ
jbW0siLEH2CfxkeiNkl2exlo81F+0s1WH5AMvBcdYreYGFxY9ddhS+InqqsVbYSzJnoUWWZZOhcF
Ia29yMM+533fnpDGOr3tsc67fT4BzvXIpPA5/0T4+Ul2boYdFT+24LIgbxUD1vKI7AfwQnSjb8O2
Rz6eEwghiCj7YnJoEK+9AhsEUsyjffGcHnKkyLU88jQaNrLCqOhmY34n9D0piHR5EZ/86vqUKLKa
H8JMoxLudAMrOAqK+0q1K//oOc9cqv1cPUsM9IRPI0DfuLE39qnNSqeYPrnVJMVoaczxtx/HFUMj
uezXRjJjOCyDUG41ge+w2t1TlWxRsplaHAsR7+tI2AXsGWhYFX/WHKL7QoDce3mQnmuY+gx8AvrL
uQWL8OdLhRPeR13DkkmT0xxKFWSVa9x1ZFq5S6HBSeIbo4GY8RepxSALAWxqOYVzpFK4jrfKMgXH
2dDR22e/aD9eJwO/EdNR/CUnUGErJMm+s+yGHQwT7ntxyvfEARmz60RtRdbVPMAe9YuKEPy0Lydx
91v3dbRogUhIkg5BMJ4jHSd2AAy70aSRzkPotgqW9+ph4dpUusXRu4jbHY84IYq5Hqfp8o8GH/DD
wVuYYXPVmGG6MK0oKh/x1blj259ZQXk03jn5HQucG5PU6MN4YQMOEl7igIdulZ8/gYPvRxFPDl12
DSSfsL1/cSaLAHUZi9Y4z5qv7UUUuPEuzbYO+nU87RRLlnSheyulpf59zMIoYjHPZxGBJOgyvaxD
lfeRpYF2WH+PplQhOL+8mAOpT1WAY3XR7rx2F8eIa5JONzR3WKubPv1EfTm3e5ne4IqUTy/odIXn
qKbJUuCSQ6WRjSnUs6I2Zfh3tWmi8N110CMUaUwP0awhn4lWuCgqnoD/nDKhcJqoX42ZcfHUAcyU
KYHsp0Hv1b3Vp1co4Q56XbkFcxkUvW/o381mhlL8VkvpHo5Pgdk40G/zL+8q87pe5XRnENCFJW28
fCbTh3xJOuLWMNjmGUbbxIpEFNF5qyik4GaLoVHx4NMiM1WtWfsPCIjdNCZM4JvlLbiXUX3Cd6Pg
ad9GSq5k24shXFsXrLdyRWQosM2GQQaZFPuMGdph/pSGcN3ApS55KTWuB9J4zfogWup8Q4Tun91/
5hFASCCjT8YU5xBfobgGRVZSEO45tISENXOX3WntxZoMcufKp1wSOXbbIhmUC63ke2UdGHE+jybq
heeqCgt7Gi1kio7oV65XaMgpX/OJgqlbBH/WnB/z6Lnmt34jKpCZDVV1sM2mEjMs/1Wb+0sonfJT
WLrClim5LXfMp7ACKmr3rJELBxOnQrzP8T/0CK0PLqkSAE3Yz3iiw/Y9WdyxuCS5njywcRh48P+G
wCk32LlQvKqptvPOQN20oCmPvBzKOgyJ/cbw4niUOUws4uzRE/0L3vwSbibhYZOHrwG6ceWr9PQY
Vv5WajGxwzLrfhDHHw1Qrei0Xr/o3AcJUU80ZcV9ZgidfEeAuhy57Lf0tR4Tprot8SwR+XBzkw2I
ePCxG06Ng27q7jnrH7BZRaDsCIbKnN30acHEox/gml/J/r1qCgdTLqNXbZUxxwOtUSKRcvBxF4Ep
2fTA3aVeM2cHGz3Cc1+vDgBMeVq/uScfMZGkfUMTYEAnI2LUJiln7dCSIKvFF4sneQGsK09D+gsM
8tCQTXaCnrYOwMkq9fhSxwCDfcddvs7V0v63JJ9XwVnMbw/lLW4xrLHoPgU3UrTIxpXVGSRpj0pD
mbT+C+K1XfoyRvPU9iFSPq2yycIqR02z/28t/XvO2r6N8hmAaNvaKYlziLXHSElfFJtVsSsECZzg
ctuIkjtCu1rakIQM1DBq55Lq4oe+RRUw8IbWsjh5mjm09Aj2fRFJhtC3G/+W44e2WJoAnQ6e6Yvd
YzJP/ULc5UK3nET4Sp4ff9pEIgovKeGBNfP6sWj18tiWItYOOL7oqmrfTH3tQqkt2+7BHhgKWWmP
hkd9lh02D6w+uDzJ663g5+c/vLETE5y0758+p+JP7ziLNZwjG6CA+UQLvcAUY5t+qMB4RmeJE83S
H+Us0RIzo7PhsaDN8s/TF+cfRWYGsU8nj4CZrLEVKhI1042o50w2p5WY5h+usw6JsHRywtpCMcN0
IJwooIRmBaR4y4LoVR7ZTFuxs8zQUDVKSwXlM9ofZ1e/ANWHggrXlvdtm4tZUZXqW76q3YePvK2z
zQSCA/XacwYUrcW7JnMJW9ZADbUBzSAx78cYevKIxGUZt33VoTnM1Az1BP0SuPuJ+D/wacWypVKt
QJBP66RRkHjQ1j/sDGqph5m7kCWMpTujvAQREaLp5pkeEk9SLfyByzRPtzF9amnl3bxEyf9n1Iii
8LnpcwikpST8f159zuczq90jUv5K1jm/tjWjskXTZJEGNiTTANItYVfOjv97Uwzq4YdZm1kTMMQb
6no99bQgibBUPJDS2LqrVbRy6ZbDr8psgID1IMwvZLYgi9YO6FvaT/vM6yJKg5nKFEmXpCK7dhsg
kmP0Mezc5BK/Nps2d8r+viXlBuetTf20kduhUNGZOzOB7Wp2Q7ggW2jv/KLlgr0gjk4E1nvqmAhd
OMX2Zwuunv996aEqzZ4Wa/7rcUWg4tP/dY6zXMr1GRGbQ0RPr/F/svtki96CUM/lxWTLAsJPDRv4
Oi54Mabc2fBY19lPnm5m57fuGSzoqQBB6Xi6YsMCABKsI/EVrJNCln2XAqkvSAjzXQerNOrk6CYj
Ekw2PTSUJaKTytcgcFe7knA0eYW+O3Gro0jB+XqqkQhZINheYxy7SiSPuvfEmE18awHdZyYdginP
AY03SRXNefVZS+6RM4w8g6i46JLtpqmffm6q4o2GN8lKMhr7QCpa48/I60yrsgcGej0dEREUr3id
rJ6xunVXmbfqVuXWFmX0Z0hN6naKwByC/cAodR6wPYkAGPWFnFhwDxJhL3rF2X/udGe2rkJyZY/Q
7tU1kFyPSoE/xiWMhWX5PC89HoMj2zHntUlgzqRWEJ/u7q6hQbCi7VaNLYb4/oFxALU/yhvwTLBO
0F1RkZkBAZYyA4avWHXqdH+V5P7BmH4yC3mDQojCs6xXm+JRym6YCwMr5AYUH2shZVApZIg6exFG
/oLW/9VPO4A8GL92QJuAesvX/KL6/5cK41D8kqSbYXIxxy8tgHugAj2P4L3qne6xPm50RQ+UlR9N
Mo2yTUfMGClkpPcSAuXDlD2zXFgg28g/I6AE3mDosn07oCYBQVz0UTjVmlWTDfX07OH0ROAjVR/k
m01yPjDTj+wp8DQ2Ewbwpfb2FcfaQ1/xA1bPZ3ooEYZpIrlM7pR2SSMr5xSIcOYzMPqyOvSGJ2uc
X2On13BnSuyg0k/skZQ0fK0ECJ+foFYBHMYM5hwdKlvV1sfSin1nYbi4mFY/C49uccNtrBaRSFB+
7JyiMXcQfHK9ewyvoEZIrU5B7g62v37gvSrt8nSVTTpxU22tlRCu9+656ATyKO8bht/BrEbuej4+
u+azAV0ASdxW2TvcD7EpmcCquqBMTNwsCW6BYTh3Ee0N4yFxy2SPo3eP3VGuVJbUelESo+2+I7nZ
hhy5V0R4Rn9TQqiTnqmrzsZdLNM9gRnRCt1W/IRxLp5+POyZ2Y4WlcmezNSEmjcC3fiEnJ1RTmW/
fqnB7wRUlmytKx3qqdLJGNUxRLSt8Zbz2I/oY9yTXDx9jQe8CN4yoR//RxHyKG28unze/H7EyoMh
WH3mShNtQ2s65zHr55WhYtPl1m/bHIlwHlBZ6CFHKfdUEIHXcVLWnlqx3tZxTcReyKrLGaXZI9uv
sEVZJCCjFjFloJl5AZ5pXxEIgpLB4ZoX6nI+Q2NgLpiXhFC3AU3wQzGAfp2JQjB6j55ZKb5hf1Oh
Z5hFAMY/I5TAE5NYIS4QvSWMlWf83yiUWG2uHCjZDOqKJKPzVbjVjCumZC6e0qIRmUgIXg8R7Eij
Zb4uw/FakhburXtWx3Q3nRYm1sGOU2i8gZgNTKLOGXXN2jl1Gv/QXI2JZzdF4tz7w2FG8SJfmgyw
GsaAlowYFuRnLk38/dX+QJ2eLwBbgIwY0HB3Q78Eqcdhr+38yW2ZSjdxCfjpoQOo0VCru4JkmOg9
ZBY8HZPwvBR71wA/iDWZhxBFCznExIlAeY3nkggPt2CQjL3FqFFnDsDMGGsaxDFlkmg3KaGJrQGv
DiJ5t9zODr2X5k741r2G/cQVccfh7T24rBzDcglJfCFb1gzDb266pqNQSSelVkOtoMJoQR10pKhV
2nYCYFDUpE0B1GqFpZ9dXuCnsh+WYqFnRp8NQnMzqkqkMScJ3qQngk9nuzk689XzIuCjmr+khVll
mKYavN3h6yaS7Gihqx5SqYwLMGmJUjkNzo0PUIff7Q+IV3Pkg4XRiZ6hvAU3josjla0OFca47Mm5
X7fEnMiOJhLEwhhrWb8Nl7i1gyVHCCUCr1x9JhulZl3fB9neb2s0eNNtaYh+xYK+WrbpXEXM+kki
vTnxYvA0G+W3nWyR7IRLTcqIp8A7eJ24B608VzItwefy45PLKvpXehH/hBKMRFRCkHvOil/vK96Y
EKMetG0oc6hJK6so6/4UUffYIaLTs9SJkiLMerGVIuFJjZ9aRQNqimwiuxMtf4LuTpQIbWXkpbiR
CDp65/NxzYec0rcYxECmiVQ7RDY7B9mYr0oSYGJak/Xm2UQ07c4QDqq01CKYDh8oCZKmIl6ey4Vr
/3tkXNxWGZ+VPew0VDjxV7NODEo2nWvt/ui7FCfoh9Sl2ddlu4XcEoKp++dX5t4PKH6hskwX2EB2
baWXMR1RHhjIUDFWI9mk5NvPIMHoFecLmTkNvf5uT47ksWiMg4aPoSo5SVvuwAQVHJOxxuMgxim5
NiQT5bRG8Mcc98EhWyWL5gC1spvk/XBXvm3aSMw7FzdAfhC41fg96Od60MQqZ5gI3sV9B1TlLMAP
nqKS0xwoF7TXnXH5JFmk7OZFcVdIVcKn74hLwWwwwbCLLyWOlNtPpFwRT0S6pv2K0u4z7Xz5RwpO
DyMK9Kz0zg5GU4I956HUho/VtPB69d3egz1SjbYQ7uyFVaoxxdyurihxidKOZB9PRV4CS/gW2Yhl
UGvuFmslVtCAVtbunPxHHEoKMohPWHG4a8bOlt2Z0JtCEhQxhN58DRrUmngmLRz8Oa6+r4GYUpOt
utaoKtbewrijQbkyiZZ350qzloU00U7pCxD/BKxeC9C4iSfBkm0OVxIMA5GSxajW2xPNiU5RqTMP
Ycll57FDpmbgIBDHR01cv5EL8UlDsvPmPG2eHzQMSC0PRM7PpB8HoUExtp7b87Ioz6GAC5jhbKGZ
evYXbqwsCr7VT8tgU48TWG1uhe/ntyy5P8oiclxU/1XmfkaGkae9EBW8GZAExaQvFHX76Crixl30
4DxotfLT6KW3u9FdK26d9NBqnTIzgKa2h0FTyGcNggGPDwgEtr1G/xcQCReFvy4kBmsEf+Jpe+vl
QpUut2Wgi2N/pZcTR5Qp93h2k+XCxiO9uL74XRzA9xefGVIO4JGUJRaVB/87LRFTT0FQfTCkErGN
phyqLtwORewqZm7nuvmcmP10zD+5F0+OiYqpMaw+sXDqxQ6TQx+ZlYfQvI/0BqW+DZdqdSDU2oww
8DzM/6MZlnAb8eMTGbVgLcpTumjRQKW/0CDC7soGlcpLwjpI4RWoB3D0Boa3q/te96nG3bhhqND5
MnfMHP0RTk+MEU98PH8uef0VN1wTzwojkwSTcrVCd7LQQAfBVlTyMk69fCWWCO+e9cyBAeGyMnAQ
blaJo3k7qEwvAzvkdlrGAkIInjAbaIlQK1aCyN1Jg6IM+3kqzjbra03fEYVuEvCvYfmvknb8M0dI
iEez+L5bbvpuCjucVnZp3s0E0UywbGU8HSg2pYXVMcw0n4a8r+TSsNvQCzmjgrYZw9eU35WJvKvA
+x2hRz59Mrd31ic8nJ4ECb5ByFhwiTqiTKMS7blNRigr+NyWuiz1gLr2VgcgpnDhhBNNdPZ9/OjU
nRCmY3Q1akRZoJ6UdPYraD/zvy9oToDfL3D13uj0TZEam3X5txtxqDCijVHcvaIGKLZRGLeaL8WM
91N/WlACPjxUQFCQ7ub3vF1jJNcjGNVAKxYcqwp3iVeWQiwBRBCN7KzBWCA3ZD8UAdcXLaitKKN9
IJErOndb8+nU3AbKlmDwR1rc5k2wd5QjetdhqTC5yaREe+OyXXYqoirWi6Ziy1NArdMu1lbuzLvf
lOkDaHDtjEyPT8hL/o6qWwC4N86Pq6WEDz9QJ+0WVObRkZc0RuyLUw1NWkfiJ+jUDcJVl6P1EQhx
omByYKSkLV0PnNmWqcpDSgB9jZUPtGKdoXkgUpploU0c+KQ32rjNpdf5wkhc2ds+FPfo+2wMIUh1
XqKPgJlfYbFnAcP94yNAu7y2i8wpxnbc1rhQP8njSdeH+4AIZUY4/YJ8w5syf9uKWxj88PGmK9TK
g578IRTSjdvvmkZRRHVfaEmKr7Z6zIkx44nK7TA87MsZUKKoZ1zlL0OYLnqyh+zsS2npuU0JzPSP
Zj6eMZnZVAqOF0mxwhBULkzV66cF97Te7ygP1T/asF4xveH79HnX1lIZLG/o4xPt8Pa5sfNNqNUu
evKLXf1qc+G0VVPHmN7asy4cufK+1dTDY1i1cdSyu6ln6C1JmeGthYdWNJho6tWOPVDUcwZToIJ0
5jf0Dt9ObbOvISBoXr1BLy+V2MDIn7IpLGuyPpsx4kAieDwVW429nroyFCHNBarPhdD/bs90UfZo
QEwtfeUtYp6s2DPuyPRPpoURh0Vc0LKRq7dphqYI1E7hw4ubTNQy/iyMs6dAHZJJdyk8CtwSqbid
CwFJjroG1nuVY2FpQyXtmnTP7XTnpXcx5IIE0x4/llE75xPbrkoXOn2gS5uWkBewfHDLjHSrPa3e
T6rmg+TloutkZ6vp2mnEh4PLgoZxlRJA0rsYEIr7UwxdBGoYgKDP6x7Dk96paqjhD1vyfB4a/Itr
FWGdpoxgvbxywEM2qpbseDKeZ1DIzNnr6kUFmpLEv75tewVzTpWUd55jCOumm23InanZ7yb5If9j
6ApahbS+FRXLrXr8uip2lGOd/2/GTNR75JI19Ci0V35lNobn9bNfzBc3uAZ2B567WVpSNQnJU7+U
+Si3dlQUJbpmNBvvMlT4AZy6N/J+LRmeSBfCisiWzwOUYRFo+VXFIcbNbfPKCWwIihj/rVXMz4/W
jf9Vgh9yZxxgmLwf7dfKaKNHysNYqIZMEVfWlX4011GC2xJiH5COzx5muxIrXkEMPYxdNTln9msi
xLzvq/Yt9tTtWnhNYgcD03DSV1IAPVtunfd7m/XOfVnJBMrcrY2X0jtpdpzClagh0BA+aT5KbL2p
VPvoA7+01lYh43i/1F1l8gluTB/vGTV8AswWzr3yiP73HpeQtWVKKCPiOkMwcdsETR07tTYw1lIP
B26Ck73NnJZFI6TV8z/GkSQ0mA8EPw35/r6wLSOwZiLAToKoj8BkCW4mEQOiwL045uXXEoP4isyj
EH+cnH+mNUuEnYm2nGEtFzQYfV78seRXPah0aI9Uf7bwMwYm8DnmCwC44r3ba45wzM3F0FlZhr3b
IaG6DdFEbCRMOcrnOcNuxnXbuU8z7m/zhXM44wWrvWOlwu+ZaP0845+nQAFMqPYEGF54PoObUTDr
9OHzWBOBaOx33qTxY0YJcabRSosA3leJNBV7WicBH61o06o832JA+5BD0GVPFbjUdVaMk6X+7oKc
EgA9Ejk3madh3stkWz2N/omqKCbyMuHcZ/t0ZcqBprOc96iJNtE0u2/UWSviKvXMMZw60kwRL8Va
y+dTA/Z7dXgs17MDSbKYhyTHIG5anVNm18axUNDv/klVp8HcmyCs1JNwS1dqHqrSAZAEWXXWU/wz
H6XOTazidCsiUURisNkJEpM7YHqVf3/83lTpLcFy41svJkbL25wFQh5JsAk8stAup58T2ZRJc7yB
WRqDiXC9TVcZimFN2OwrxSVrthJphKp2eAX0G3lxJyCKPz95Hgvl/jGJ7PR6enJpKT+oQw0/xDSn
b1QCbjLGOz/rkx4dlty7wvG4CGxd1tfZ9Z45nvB901gWI6fgrplnbarNcIVEOSd1Mf7sxtmKgq9C
dMbYw6eK9380PbY01BYJcMS+a+8IJcxezlCU+6iS2oTdEBqPvtZ2qvjtmGWPwyA06FaoSFEGzapY
mbn8X8jUhG8BVG2XcLgynv3FyWcfXAuxEFAC9/Xjzw3ExCvfziSH8qmVdUK1Y8LSMymvIofVXJVr
qZl44NWzxNoK7aHeyusBPceO+ihnVW5N2GE20lez0DJvuf0dxDnH8ZiKGX54vwweBjqtS8XHdVdg
ZKUAQzUTVSD8KBXPjCsYeq1dXxOPJ/UUgrzsVF1rJmm2yEXeRxtULahCa6l5pM5SPxg1o9psDQoK
+0lnKoG25fn4aeSL2g3UiUQKvyDELbh7crhgKeaiOI5BfwZ5af6N5RUApsQNL4anu2kNOnB2dvrF
byYSsRNdQ0zz2UdXqz75pdPBLOfyjfKeJ1/do7dViUhhbLfElVEKrfxbtdfef2Fdz2iCAGbCXI8/
UfX5Fr5mm3Ym1T4q93WcBFYB8mfPWTIfkREW/RmMHazkLiF85Kl6+avvZRKNlxVdjEZyCvfXk/81
dSnoIsgd0XvwFGY7MIxxQYMfZ3L8FWTNDowgLtMMmYUobY+YuF9R1hQMMWSAVL2635UFhZ8yAHu8
J/SZbU0OEQI2QcLPnC/S203IjkLis+r5bbhOlxPOHnjdjtDOv7bwHVFhepFlXCfJYGAApjEBMjbB
Utj7NloUEYjq8D1EyPS3tY9ENWjHf/JkA7R3aLsYYWdV7SbVOmEFnsUl8t970CJGLV3F5LWuAYz3
b0AY4VaCIwPsS/X/l8tKWEurvoYh9aiRYUmgl14QyEWd6NO7t6wM8LkwUociXkpmPBoaeNPmydNZ
x22o5DdnaZbGn7hfU5sbzu9g5NJ+sgrrl2MALpIn+0UPh3Hv4aFC6KJud49fbW/Rq8DKabuEGcKE
8Eb5pLsQM7i0ImrZzsy4j2DV/I5zKHW6qFxjnEaT0n6PN9TAfqULtofnNuxsPuS4oXOtqopzi8eK
KC18adpJZK6DhhbzECJVNtIOYwbyJA3/sCc8R0s4jEnqVRzyhBtlL3h6CTzFp1X1hrNd8r0jQA+F
vQwGMWuOMtI90ExWSuGXHEx7PjjATxB/KHIRRITMjYKjD/f8a35VGIluiRbNRmtRDDdQVDaqhdXq
D9wmUjCjbQ4X/oSaM5jleQTtSGlzn4LxnkQP9weidVFhKZtPf6+qho8/CqHGCCuBglV3sga+8dUp
vqbVIjwStd6b5rfQrIjB66dicR9LHp5kH4q4qwx+20jEN/Nznd4XJpPazuYxyxFHnpjTUyKyVsWJ
aKv913R6QjIhUrLNoWNlAFAg4H/j1vncIwo/UR518LqXWuoSS2wssphllMkzYsEbpQHUnweqBFt/
NqeajiOQm9O9AAU5G+cI7q0EYqGcl/VRORCIVph0ixxVLJqDw4lVeXpeOw1enGnsKOFfN+O5ObL8
MzRnVkDnwcMMuufyZFUA5N6BfAA2wAZ/wVN/eeUuwONwDwUhLBaFfTV/k5zmufNB1oMXxSAmBexg
7nrTKiWs8YhlQ0Jj2Ikah8cZQhdtnhZA67VrfA7SIfVsZzHnmfFOv7JG/F+WIgzIDmoYah6SE8Sb
pearR5z0z6C4g2cZgOya+mf+3vtOmDQ4hyc4eOo9T+UDkzGvSsR983sdQGuIzR0A02KtpjHNcvrB
Cuw1BV91p3VuguXEXMo/NpakK3+UDD30Ji/PD+Z8GStzfnmxEEiukMVbtuaFxG2AErrNKw7GEK67
/7I4d8ktfzp7UOkTfzGPEv+T/CvR30o4r8+SgMcj7SPw9EQWqSvFi2hBofq0vj253j2HPeG+diVI
muXEVovaJLdSaE9AY1wJ+tJP8FzbReBmP+UdnqDoVBWRUxkmcMCMyu+dQZPg9VPwT9FLbl8ioDrl
J2pyTWu9P5wylkVwAh0hJIuKr7W4nDbP7VZSnRvrGRtcgMHC5doXGaM38BNNVB7lV4y7H3ZSDTzd
qaQfhINc8dA4dP5hryAXLkN3scplFfvptTi2UKj3VMqfaorwEJDzKpvDoPgQlx7IhTn2wWH8T/yx
P0zSdvz6vlMwCD65W2wiyxcxvWt1A88SzzeiORQoT4JRKYdm2oT8Pa7PfNnqhC/+SsoXtgYHVsbj
WafPinxGfAaiZZyp8tTdzdLSAXqFIol2esT396rLIQzIeLNZ53kkXKVWHf3MgaAfUNsJF8XBj4za
ehhAGH3AflyybHFOtiY3kyFiJ9J4bPwZaEqbQHOqRYnjuPMPqsEnRbgEyYzMgKnqaX/W5GSgDhGy
yFb7IATvdZmyU9JheG5QIYRmvgoz9rCXhHV26dZlIe8ahzeECODaXd8lJWw1rzBHOLljsWTBp3dO
/CMzUDYm2ediK7gYc5uUxR7pHNw4Z1xMvobphva4sYpx7yR0VtPtdtTacYcaNfXz+AvpBaus1BlY
ooTj4Nkxb+9S0T6oQqJksa0xLXopHMPlhDyNutXORjrjr5IezW+lFNKxFXBEujBw2IDf5jSGKVJe
FKVUAWs7g/XfmJwloSlG8manvr5HF3SHxrcgxr2c/ncbzkZBIMp1VIw+fDla5tHDsBQEJSUhL821
Yb4hJfif470HOrkBPPlkI+dCJpu1HSbhrpB5LCIJEnPQVAD0uYv/iv86lGw3DHfAbuqTzV4WI89x
jnTmzZhDN6btzhN01SlSeI6f38Qm2KfVxjFpR6MTlyGyQ6y6H2oYFv5q1auQtbHozgmfe1iC4ftm
wdwvyiGS0YwBKZpPFViYZB7V1vZ+u/7iwEpW3CRdASFQks8rFWBWssQbjS39h8gQpXCvBhB//aj2
R3ruES6N6or7fMLLN4TB0bjLTDk6EH8CRl/i9yldxKw5LIXX/VCENVs3BYi1EP3LSYkStmgkb3uS
ostXWcwWbR17oq0xMFdCjwXEbz0Ed/Ejj74+g1NmBvo7VpKhCPjOE/xuKSz8u9DCcsS5MdDEdiIK
4FL1+ySeVV6Ic3mpEAVo+eDq0C0Y4yNM7sH9usPgs0ml75RcnGweFwdptffIYDX3IdvdHzVgbVVq
eoDmu322zqEAiTVnGllGdLNL5bZn9/ySZpWtjKO+4DPsCiHl+pTt9aJeJCYCQ59SUr7yICy7BzMv
moYwCn86mwTFDMXPD8h58aPfvyY1GIy3yhnA3Jrd/KCs272w0zRPFcxcYDVLAZXvtog0geGWOdH0
QBaWuap2cJ1DRuUhswweLn2xhcKxMNEmm8AuaWIpU/oMxQx3ySidcl1w6y8yfqIDYFiNq2DsrKNs
UsuhS48nlO5Bf9IpAzW0m0CHbvj1iiPOXJo7Jm2rCzz43Q+P18p15lBK7aogBfSANcu7W0lwBpto
oPMaHqxsY64iP4bekFSE/3l9tx6pLLUxA65otP6tBcczLgC2Yxke8z7Rf+ybABlKuvY8dnNSz3Uw
LmGV3uVW7OJ355rRLwH0i9fv8zX/o1Ddf/C+PCP5SP7VbB5psIwtU/XVsDNGqVcfD29SkYY5H6OK
uJsYUiSzrGJxfZZ4LEsj3MzIQuXyB0oXxl/w5Mpk23WnVTJEGWuDRAZ/qozYEHk3STlxiIUDqW4d
D5GaI/zdfRbBKAxDAZNvZ38/vG6AoVzh11IicwDyiWh02QiY0j5omFTzVMDn2s3JA5jqXhzY0rLV
KYlpw9WOA+JeqJ4gbQ76VMCbvGKJ+g7YtupA68CDh3BZxx8clLWXi9eoKVhpEKDB/B4SwFWdEniV
sim5xLBfxwo8jlq3CpVidgh3Gt5VG1qPo7/vOv9HORpSkN0dWrCdmK8/ly7JKOaYL/0tqA0WJqTQ
RRigPHmuLfRPOAQftoRZ+rEQ1wdlbF+/k6CMTEjLvVJ3oQouuvSZ63rkwBMuYd9dwyx4RVz2wG65
Dim9h+KCociasWkpUtieVF3s8B8/mJF8ETU6VuFmXXSTm0UL/dFpCRfM4x2BU+ksHabDZKXm9CtQ
4ldWhca9vrq+C5pFhJcoGIDtYksbMF2xYi/YaIKmzvR+Vd+Y471kqup9St4wQjuWPrmaecXJKMNr
IssRN2gvf4jlH2dKg9pYLX4DXEaf5BROgHt1DIGnkUQ1SpJT3zytt9sOQfTIPlNACYJqe7VMv3Cv
ywXsdOGc6kUoWzEXRA/65M0wWGRlcks7XhlscuF1CpCZSDeMyYADpj3DNakdParIkLgpg6cbtKXm
XrRKr/lNi0CRqjTYxaThBoO4o+eGSn+zcr66dHkupQ9kvft1oljHynoNppwdhWTHIJeJP3gsyX+l
0YQ63z2jze9Ns7dkacjshwmOOzdxxKDY2TNX0+2f1Tq3PS68xuHNjT3gGjQlMdzJYntKed+4gGuH
gW/5XAdrLI2u1FmwOK1/Xyv7U2YFAOe/Sb3978T/3ohnIdAcjFbt/1eumyBUCdD7gn/xSNIIf7rE
wcMa/Ryg6EpXJfvstQB5xBILnSxnTkkZn8q8W+z+TYXOWmsVaCYIX4gx70RtZ12NKCxK/amsi6BQ
GVovAzQgJ5aUzoIWm8OmBgIyd1wqXXtmIPWISxuw+0/ka+6+15hU2ojjm3OdW5DbPXLGBwVcgBvj
JjXibOMZdMykhU2pdZjuWnez409+zMnQnR/VQRkngJnGwBdc47LZOsviR1qw7QVShGDTLJJKryCo
0xANhzaPwp+E0h431WUdGBB9ZZRQf1OoKQl8aFl5EBL1k8UjXUhd1Nqe1svLsyLc8ODQ0T+ixrBY
2oHp7XrWFT/NLdn9fkAbQ76pdkcGvPcnA09F9iGJ1ksqrMNGfLTKMvmMN3kSggCIsa3maWeJRD5q
wsT4PJdBhxgTaWTayj8FlSw37rGSxce8HLsxZgh1QC27TQnM88jfSBLaFM6rcWlQZuTquPip1WXL
5e2Sq/OTffT8OmN1gGFlh4oPYirmep5HEKRlNxO+GuTYpG2xF5WW4z1RbKYNPHWMO6xVaVnG7SU/
lL40h2ts7j1UPgrMadWFaUwmJ7gE6GIXMhO//RUjEybKzvOsqoM+S6aJjQz97ZyxRJViB9jivrqa
fstmZNpkIfVvhhOxwYKdp3HzQbJ3Fk+Mj7DYbcfJbkrEjIVdZ8VxwIPfaCY+S2CjmNkzd61uINNt
0q7K9/0ISu0Pijp7TrQmprATVa25FLOqS1s6bKNoc5AMFbSWOlE7A71DxYthdfz2WpXSVPlP3hLi
l8Cnu3vDjZ184SGBQApQwlm5WKV2JJrjGWOVjOuQ2Io4KI2PGIVjn8Q01xn9YXgfm3eDWpIlXgRE
DmsCpxu02lOoZqPblpicWeHTkTxmV0WcrNjtJKESsMyg+JMmIgCLEommg7ry1vP0HsPZpBjRObH7
X21/3bptgwgdjDm7Pz747RVE6+yqLr3/rSgldV/aY0LMLlCaQ4qfSWURJgkSymhDNEofXlWvBvGz
d/Vsldprh3XHnB9Y1NmoQfrmjQoxMlbBunGEA9f8BLl4g4eyMx6di7qqnfbWyPt31U2qQSzJGUpQ
PkZAdSu0F2GJoUQQac/X/NEl6Gzj8A2zdALuWa8YOEBafEtB2UnB8U4ACyKNWMvu9I/fv7x8AQv1
7tZxx8o6cuLJIK2SZ3YFQ2DgemmtAsHidp392IJ+N0xykBINV4Ce6CBdZAyKDsQoGypp2bVI6JvE
kEsEvCzBCJoM2ICYOAZ1EvqXMW/Wcp2FgS+dwxjwqECl0nM7V6+lARRUZRwoHfdtgJ6PFBv4xta8
xrCADSxcdA/QpiMJRqSEPNtfTX4uUYcrXCLTO9g2wklc+8BRSg8va7p6IRs8SZb6Kl4xd+nWHweC
IFJ+Zt7Gp7dA/D5EQ78ZhvrhZAgB4xe4DMQBGhkvVTCA3r5joCuprJhxBZUCp62q6k+rtGkKgazm
jeBmvkXPP6v0GsMQ0HzAUF9lbAYptR3ktF6dVKnQ6hl9ylhPEvbY1eDSVCHL9E7qLVFtPPXbnH07
alOOZZ13rhlvmal9ik7W5aEiJhZI4JrQ5Wg3WRox0BGW2aZ5jSs3lDTrgu48sQcXqPvPoSv2o9q2
0iIRCIh4oO30QxSFKXxTsbFRAzQs2Mx6xrn9ICQm+zDUduxto2RpeBDD+/eD6OpMtRkpv7Z8WEKU
YdyGSkvtNhbFdzWNLaanYYWEhICLLHtb8YgGyVCy9erGy9PfWFmEVMum1CfeF2FJKKwQcD1MMjFq
e16TK9jknCLpELCeBrsHiuCt48T9A05tjDF9Dz5Ey3JH+6Bh5Us0rxJyB4hAJ+9hgUzp5ydf7D9o
gJFknufUDlDxijAzvGs96LLrQZDlcJmI6voxPczTHfzORDZxD1ZSSoqBCJZPd5wASBemFVgrrPZW
SeS6S8NIcNIbjZmawg672cXxuLULNwgwXQwonTLVmfO7qVG3LuOPZ7qPX/zQAfdAi6656lGbO3+Y
s/mOBg3QY6DAWQHTNClsN6zr3Xd9A+C3br7ZMhCzsaX6geX7TNh7UnYbXpyMgB01TFVl2h64L07G
VZ9Ya5HU0X0gQJLCgVVsGIElK50564cTgA/bulOwXQx8uB2oitAO6ObQENFFYZpzZhWUQzszOvhO
glSddOfDqUemCzCLzPxr9aq1Jugp3g8/aUtqjKJoZ2oCG6lt2FFFy2UaHdjgK9ZjJ/PF+wJskglH
QS2mxKU4bnd2gqwjQ1P2xhHX3HFGiVjPNlLHjT8QM85MVA+hK5ZuSW7yESNdDMUcOeCWEBADQl+W
hISrIHr8jXLSH5Ht6bxisgg0lPggKbLXogmScVGpsMhyHEm//BUW0MR4CxCEWkJ+aqINCAGTBSUk
s4K9RImKkpV5M9yF/f4xnsJrSeJd22pg2iYXp086ResmNMYdJ9EPjFN7ROrWQ0YIXk+QCtOD/MqT
fGrWMLe7hDmbjTr+1K7sRuKRiW4IQydGtdrt8G1wWgPJ2z7M0RI/giuF/3XjidrJvSF8E6jl8qbF
jWEVn4rOFaWQPaaXwmErWE1z0J2V0p3hGkfjZOGUsWDPV+5zpdmACjr5zNCS9SgPOA/uv0qqkmCF
XuNjwoO00WnMk4Tcg7mPO4jZDpls+WcaPdr0Yl+2ZjuGi2QzDHXKKzh/cIsTuZfHysEbLB9iVsG8
BDpWIk9j1O5bmO4IXLlw0eMEaCp2dUyVC12ox8ncTSp1F37frA0K6EprboE0NHWuJsbXnF3WNEvF
w67JvVzsO6VhZyXyY2tzMbYjSR96mLeoshGP/v/UOko0tE99NgWOs2Npg5wvv3FiO8dCeYt2mRom
UvtnpgSh4tE/eLD2PQLGhCSIyfE5QiyOSCsozndgXIn/RGgpfKioP6cPSzZLPpQTeobtOBxhQg0M
27kK1C20QAXktdjJdsLfYe9V5WeNtXnSWKH0abzPPp3Z1ZUz/E8Lc4e/GV+WLJ4mUNh5biDEAoEi
sueLQMHWx0M3E042JDaO4HhhVBCH1Vsd2iIBprN0OIP2Sr/srGfjkDAsJJzN+/QuXcEv1zWIiQ+n
80aHCltNmSfuTDpB/8ifLwYVFQ6XGek6jJCKJ3HUhIgkw2S9IXkloesWxmzou3B3UuFdipGxm5Ma
k8ZJ/m5DrQdlq4XowXe8m8w3JJIPuyvNLuTYQYJeHqqpP0pEy194zpG3GAlA56iR3OZTraryN/2B
9+pxRO4pFTcoUrp6YO6TvvHlXGtlTr8wL6L2Nwoun8ujld4D1cDjix/WEKlcX9xl1RjeVbeKbOCG
AKTx9iC34rFAQfL0cd+h/ka/OJcX8WZg4LI5P29ZzTvtduQpNLfHScaRSE6vuGPCC2l3nb8O+9jx
aMKNQcLDJNR3TMoovPWnVsVv9I2sm5SDhkjMfYYRS00d85mwRIWLXtiBeoTM0z1y+RxwGNdFO6H3
Cu0aFMaIZvXY10l2ewCldlaLaiqUAkjBYRLmjI7CTAHRpwZY4F4UZtrpYvbECB6HOutf/Pci42Ui
6mpmy4qtgwkL24rPL14E7gDZf2zHu4BiXj9Qg2y/DEhmFHFifvS4f+qiqx7cKRgVTI5weAGbsaaZ
TZ/SqQufdnBQndKUR1Kl1fuN6tZLq85SkoP+ruge4TSH0ZmXCiO0Ii+ccj7PhPtH+XqT4qmMaVH7
mS4vMxNaObXEx7qdvwmR9no1ZBv8kz25eOlqLE5TOPnjdoXHwgGCfXO/3zzvg4CWdtQylQnQ6dpX
L8odrxGAO3A2t5PnYSRBEycP2AkhWMreAgCrGVgJJ8m/jBOOqOWXB5ylTVQ0wej/HflqCwwCzJsl
Qf2FTEB/dGOyexZSQKgr2wMOKckVh4pZihhHBiJcxIQWU7lBDT4gX72OJrtxdTp1JUYWiMCYagi2
+xxVjkOjdkSGxsn6eUy7QGxgQzQK2Ik3QtSuM9THg1B/9efqbqh9sjXVDDxlFLJ3tb5vabTpB7t5
TFePRCUgKMl/qUnvPkxNbUUle6qwiWDGUy1AinDG/G2Va0oe1LMINt/PWm7XtDkjvYZxqGz5VcUY
20NDfbOjC0qXwFmhkwfrBNBmP967qPPLGJSumM7MzsB6L7pk4cmrP03Q4tQ3JeabU0a/xzG+4coJ
J0q0P/jF3aAoFofaYDWRSIuHKcUhZtf0jl/QOJzb9H/welCXzwfhhzr5GilVMSSMVwH2U1LGtV7n
6SJNRGx5sW94k3b5xYH9VQg1YY3UjKrgQRzmF35cWaRgVjQ2LKjMCoUiDQ2b35+/DqkjTI5cs7vv
03BzWqu60FU2LuVJMXH5omcRw2usLsPm5zozfumC4KcIkWDDhBA+OQyeJNMhysCUG1BuMJCvCc/R
4N72eSexLadSrcIrXBF6DIBrQmeiZbEsNsGfPGjpLzt63p/1QbwK+zeXpyQclKFYv4SkIZp5XXwh
fyOmbhqpl35zAQjJnf60l0WM
`protect end_protected
