--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
iYKAgzzRNkZw9aXFIz/YrLoCOUN4tektgy+siPJlSAg2b4bH+7IlzyGC6NaXdDg8HGasUjn0J2NV
6uGN2q7L/LBnD9a5do7LIhpf01TDgc8LLlAam9OIKITWdF5EhFuhSJQVVnxMdblSOMCFDGEytIY+
WMu+Idwwv/1iFuEkCFnIyxM9SUf21HDdEywm2vhF8X/IrZD6TUDuz1KXwFSRN3pEZaEVt4sDgCqN
LWgxfXW+rK1DMx0gADYkm46dNLybXXqBatefeqZ1EP6m81dgXc+fKDyz9FAjHcL+ObPS2gBITNY1
4rzTrk2ClU/CzpXPP1ljRmx0WpW0msHv1a6nMQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="qnCDOU92gbAUk1hOqkbyNH+J0ubLtJOAQYl5M7edXVw="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
p20qZqkN1Y+QODaUIOVLMJSUdsQT93x8GNyA/sZzGv4RJz+WXlTvlks6DysQtY87ywuUpXKBKB35
D1RaxS32yY5IKAKlOOZUDRLzm2DV4unlhU7JslOieMj/oe7S5q08WfQ/gWrplNJMzDdEw2zeTU9j
7xWM0WzC1Vtb7Je/u6kqm9wrLtK8QlUEolfMGMYvdYPn5Njpyxl4LEFThuxsCTpd/POSXycYlgEc
cf4nvbzrr0HNo8KXOm4wbHAgzRktYwrzAPgbEFVdZL1Z0v3UjX3EkgTRWbD4/pza5N8BZbC1MU1A
RX7twV+dkvKH+X70qquJf1QdK+oUsFdfbG8Zkg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="hg3Hvk/HaFEGVjoYKSceSGRNxYk8bDgD9a3C8OqB0CI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 29168)
`protect data_block
XZDSZDAwPGeIx8fnpg5hKqYMnt6htKPi/0h6G/4HPhvBpvQY4Bd4Zw6501CGCHa0dd1fIW8r3CSG
W5lTjU6UXIFYMTRirdyskx26yqdLLseXMEutjeSAl/0U9WRxwB126xW+i/wG/HVpbQMK9FInB7Mq
T2DSBUSIYwi/0LjBe8fikmarWImywlUoAB6hsF6kOOb4QJA1rVa3v9jyU/bs+M8AvCAi6fDJ3nUQ
2PnQNtF9s34KAEeqMv4M+Y3ytpCAINOfqSB5vt/8Zf4O9ldUnD64higMhz4mWgePtitNtXbH7Ps+
XITe5+5X7IaGTcW3TupS3AxG8rZ6wFo6++6XgrGMco6KICqaM4XQzKBnshVqfCHZ8m0Vy50Dhc2/
6f1Jp4OXpGH623FdKAvYpXFFEe+9G2F8QbVDEFLkR3vNCASpfKL/NoHfeTzoT7zf+KDySh5sGSJB
mAfb+lHCsQkucBRvUelkCoXCcb9HYHDBETjYgmfLVp5gFC7yIh3lCxjwN3MTE8WJJ5XI3k/Z6QfS
+e1Dfdb4LuPMUjmZLuQ/N2kkqCii0tQYWqm55ppNFsjq7PJ79cdnnKIZLdAN2d54RbKxCt/BbhnA
lgcpk6v1m40FZg5pCLtvXwoiDunenzbV48Vs9olIHM+RPobPA7YKI7xsiOn4pNTjQ8oBxLUc4Luq
9dMG224fMku4UX0LpWIK2k9qOG5CUcF1vF2l+lBTMHKahyExKNMpgqtz4py9SlPCpsMWAtWae8C2
ZsgWt/yElnmFzuXSmLd+AI19aSZELAJTFovAjNrVTceJV7gl+IC1cw0KnwAOxugezDfp1BDicXWx
zWXEvmFiCgh1UG8E8tcxUGGqxMwr8lZS77nE7UxMMTm5Wo6J/ChhGH+bUDo6oLyUCOmFLfO98rI+
q5hQcM/tyzugElfw0zKtdyxBT0DrJ5qpY0jdq0N+zKH/eTRBoiFHNaMtRzgUp8hw3vVAPIwVXR0e
xiJ4JHbn98E02IBwxptl04eE+A6CSDETWG83iH1Z3DZew+TBVptiw2uuc9IPrJjp/eAOE5nbRCTu
SXSO4jQnCUpuTuMNsyG6J1Q37F46EEPFccKS0I/RTp78sjiVUJbU6LtvSdhxvntnriOPYpD2BKJs
R++76XFbRKvELm6fq1CWnyWGLHkOMWIi9xFXl97+OKD8L1EgWjvITU9IL73ZiGfeiSNDsEd+A8e8
u2xPSuK07yF3c1NUzYVwb24D41D8iNQCwQqTi2CgUC3HjG4Q9SqROQXYK2AmNs0z3huINfgfRr80
43sqswTHjK5v7eXwCkzQCd7vpj/aqQU+UY4l143cY7wS+qXyxnEScQnzSy3YHpOJ32uKct9Y3O4F
C7MN0gMzmiOxWXDnWrfo6uIOU60EF5fFZenukhNmNgWq66fEivNbiZUd4FR2klJhxMYpC+NL/xIp
+84urQCMb9wZfuNrAgDf2mmDl3FNWOWlg013xr3/Q9D9EY/Ab2qPFaktNKUCVKawBMbU2L1c96at
x6P+6qlLtNcFf5jP3ImvKeESu+KKUWWN70KmAAMxCZFggmSU0QFxwntmJ5dOqCamx2RNkP5b/Yu5
bVGjiuBm0Q/zdf1VnwCJxCGewf7+0Rn5bKotM1mFc3hI+nn7bmaiTQ6p4c8ff6YW2BXTz1ZtMUbq
qZzb3BVGfP99wnfNh1Lg2ArYa8KGw1KRsxb3hXaR7AEcvJNi5sfZ0XBPq/W1hIZfFhYbBpq1lXuq
GMo0Fyo/iCAPONKV9EdSRTUtaQJoweAGIMXtAk/QAZ/uxeimPrl8EjroNnf4a8nH/XZtZOvRq8I9
Q98akGUd1OiJsmLqeSC+GDyRvdmkrgDtJFH/DBZzIw2W3fHtkRwMlCPVed1zNQ0gxOwjaFqmBCjD
LZ4cCen1ZjwLoqdm2tiAR8hF/eX3+xzYkm4pXbp8xCEHxWqRiaBUszftS7Bg7c7+J4CBR3/XCEOA
n2YFue+smT7sb5o75UnDrdalBP7Vz84gzRa5dFJeq2lw0i+mQKoizVLsiuLd0thyr0CW3TL5hVrf
FKf/QxeMH83iEbZyIppefwvGY2XcNDhksGiOMbjYyrg4nqD1PjEpNxj8ZfLU3MRg02oZQNjUPUAM
Zhut0COWyX+mg63IVD5qOQPAKQV5FjKtqd79dtoz3a+D2HgV0dfSeADLUe9jQEz8f0ICPE3Y5uY1
65uO0mEP86vi/nZpWBeT8fSnbcWnWqIt56nGQ3lxzxNVjxtGZ15+HFeHdnKTabTEf2EIN1CpSxbJ
VsRzAKAYNeNBLUJBFVGwwOHow0qGesDtA4J7WhrvbDPDwmue5g/FNt8X5z3h/X66ZrV3d5ZcMxNW
xlTYUmuaNQWRD+HUkCHL0ZjX8QI0onkit8d3l0RMMK0vw/zR0LlV/6l7ENYe+0K/cudwc/oAZc/b
HuzJGG/o5Q4yDzUJXDptM8IQ/UJ7I2ept0MqCWdRwAEtWfeuB8PVs8q4w/KwzJ61m6U4CFEQ0jRO
Fqt1PBNIK5ZrBqBModsMfdGcBxbKjduNITdJFOQx+VNASAyirrl4BDew6fUp8K97WJyxAV/ThZ03
Cdwsyeql5yD10Ez6hanQFGgqoiMT27ZftHkKkkzZddDzievG7NGL9yfcz2g6Dny9CoQbVvUYSKpv
GT9CsXsy/wx6WkPr3bXr/HKMcmFOWXav2VNXmRFVxC0+QiebXVwCGhus8f+NdgIVLXlXBmr6O01l
FrfwU410wpTRNd1Fy9dkWQsUNz/8BnOBngNExNTMsmRNtGv75Q0MRk29WtUx8LxeHJo/CupUj8q+
8I48Gx3QcrVkExDxpMFCYa2uR4MXN3zybLBg/svQjMQN3p0lAnHplrn1rKSxY/xrGK+jIF0U6Hj/
9PQbEGZiPzs2HN04WHSp6X6tWrKoXcJ8cxNGmbRashdjRrIOLH1X+hUqEzqVYnrQiwvcii+NAtzr
vmzHrBSxiTofePzPwyaPv1cnzbivWGHAEq5nB8CoFONOonmX87LgZDBzBQSrZspZPFlW2PA2BSBj
lv/RGJZny5D0a9HW+5CyX8foH6BjWz/OTSsSp1oRn55t6HJtGDJcV36cCPmT4VPTht8+c833KvWM
9VUSSfMLvEjXL+bImASnh3zIUXeMMbXnoLOaXUMndRX6aDw2Na5DtA4pX2VvFGu48Nj1UpfV5e6n
xUhAR3pObBYlaqwsAdahu5UxrGaqYURHC/1JeuTZxwCfMqIvqXvTZpQb3b1isFNKDRcI5RGd9g8y
DYZXh7hibiz6KZeev+w3SfiXD1X1X36+vvACGCIpTwjF4JCeaeBqwJGXvPhmWzYZA+h0ISYhDELN
jShMFmCbucy5TmbGRvt9GdncYxDjb/4dVhUIO+1//UefEwWJvTXVWssgc0aXfdaTtTEwM++bNDbj
0Jz089CRsjSUCpBr7qohmkBagHXlBEptSKwo3YS8Oo33W9flW3e9IzrY54rzuaH7KqDkLsiJqlvP
7JYQ1GkA3VtT8iq/7AaugNuLjBd6yIHZCMBBPDK4tH9KvVb9MAJ8OMS61Uh/wSouUimNZ2EqYEws
fFRVwr8bTnYd9g0MHzTdzW06+r6a4PhkoT6DqQFd2Ib6DTkijXHZPBHwUWDYXC5UhX5At7D8NBM/
1q3xe/CRboEA2Bbm9L5GW9LptWQI0hh5ZkwuRe7z/4TlfCRbuj0DIodZAESxbfUBV30IFb7dTp2X
/fIenWhwbC76zSSJR1MLqGZQdKKLEJtybZuAQDQC9r4kQAe2y9EwIXp31Su7MGillStVUx5oDkr0
ol+XmyU4TEdRkzF8cdMNReAap6OUiSm95epDwmKiYwKn6dj7xk70f0f5iuupBH385hHnEgEEjvfX
PdwY+qNjT81OhkiiZQVEETOSe1ef5rkyQPV80/BwTeq+e2pmAb1bfTBpz33OgpTody98sKi6R66k
A5qHsVtsOlPWVcRsKtZ0aKF1HV1ooUFcghaiq5R/18x6Gxw0G5H7Z2cyHAzJ3Is3VFjctHNV+xiF
CqqmiW5SetDilNBDYg8MsSftKW9rRukXbpMe85TqEbiTjGEfQr5G24iuk88hBrxrDR8U+O2oMxoF
9WDOBQhy3o4PxvfLWHE0ody8RMCxY1PrzMPMhb8V3uLOEHoniz3HLUsLnBW0SmYihoKGZ9RuUc+H
0fIIl/oqoxCQpo/VoZq6obkfByTgDaU7/fKLnPngKCAuQ6wjruU2ynQD96S9HtCqeJmPOaat4IS+
NAuvo2KSAZmAvRj7bObcZpXag+jlavFpn2nopa+1Trpq41vva09P1G7VSXABAtPndP3xpXZ3OVJa
4UIFx9Byy1Orx7EOYIFpo8yABTbR2p7sj9UBfusU8y7YFymWhgoCc0bC2BE5W8xqSETPJdFXjYIP
Vd46STvzd+gH78ZA6yexuG2M1lSzNtrS3Phndb9KMIDSh0KwSmlMkDXMarQEuuo7El3C+Q212Oi9
4paQllfowWT79F1PH9SJ5MiMu0vDSpcT+JSjgqAmARqllHH9n0I7Bek+g2SUs93EqCJL3Y0G1CAe
yACAyUn3sX+LbMYMkyFn0FZnjRZjUSOtAdXCjjEiG+v+AT/WiRrQDVNlZ9KJ+IIfQZxEzadHs7Jk
/L49ZSduub/MeAHcHDh87C7TyO/0sjTgv0M15Q2ntfVRBRHqYvCx/JwpWoTo2S49tcScwVgu+A3l
U5/3XNpxd3e0qloDj7zbk1vEP2r2z0eJb6W2+/NHCDTJhSvTvInCj6qLDnclLdoBh++OiKIOmZXp
EL2BOKyKwsw9LtczI9oT3ssTVP9qcP1RaiCBYldfRDzYuWLTNX/alQxsETEw0aSRAuzUlSRDdYev
A3XC+PQmdrzXOXW5MHFz4Pcuej1hEsNp7UsIO7UruEsdrC+t1FPDqkcFaCd6CSmp44pz08pA+72i
ZcKmXij9tjGAadkhr30S3uOm2tBI/dzceaFp2O9D2/znPiXZu3JM2oELYDPV55x2oprkMrCssbZV
A0K9fhoTwDiu0q5hwhS0v7qRw8h1kMnSyEy3y0uJrIFD+nZBI5EEwXngxUxgoSdTI9VW58WjT9CN
Dk/yTMajTWlRDApzRGuvcpGWeog0XcQROPIifUXlmEpxvvN8iFqK2b6Snu4zH+aUMX89gezikRvz
vg1A4bSG16TUpOAAafUch9lOj6YoClDO7Yn/pTfN9mAB2RGgWUVhDeTRPBS30xemQX0Nh+w85Veg
gff1HVKq4gE+QozUDK4jnvLkK47NQIubmQNtGV3jz7O5mTkbvGffZd4fZ73VblUFBk7xlMvzICKT
0vt2o27dtOEf2HM/zWLYIZQoTf8oiYkub/P6rmdR3int8lSKMgr/x/4c8qmIw9sHuajpRQs18jTN
TCnWliqY15uIvvGWUS7ApKk5agHAlF1ss+K/J0hZp0UQvJ7BGP+v63SsY+ZSP7CnQL8Ls6oRt42K
RwDWl3CNHkHTGqINRL5buF3N1WJV0+LHv5py/TMTY+nLqekDx0xoyDgPEKFQRJZLfybPAeg4aoz7
cCbpurg5K6AUQOWMuN12ro9LDvwkgU36H0GwTq4DcMCMIK4OZGA15p1JFHQH98LmgyqfAaoAdO3c
a6Mw16AuEHXX/vdOxEsxPfseC/OxW+OnbrLFpw9s0enZawc8pOwy6beq8ZB9uMjqCjjAajFjUV30
Bd3wn6fO8swldptXQpXoLMmvmmnWzpDqjBqxmx85o2SGsavZF2V/0iGt3kFfW4Sc0mAC9xTOyUZb
SKmYfTAB6Zuj43wMTjLJnEaF4qzQSmffaRQKR7By22qqXKORwDyQD7XpXxYNWKu0wtl0AQSZzWGj
Hkr5VMO3Hj/Vu+XDfmJX1loW0UiRnpW3ERrm4U0Kzda0WloPDQimHm8B7B7WbHY2f5hjNwALvm07
+eF3chld0scOkHXHv/zi8eRWFVS2YyuBfBPR01de76+X8vWyKe6rNzeW/Ogf4sI+GYvQ6LSv6qnW
BXCd6f9rTlU22XEsSvdKkFLDDCaUl5GYJm36/bloGJ++NPipLaQNauPUbG82dbLxTYBvZZBAW/aH
3zk5/hgFrJ3gsUd48go+eVxEVh07CegMzx0WVcTcVI+x5PDzKoGEBsHw6Qn1jys/IMEY5z3oIcAU
u5yZ9ZRpphB1EJ4kUxsZKLYmn4+Jeoid86glNjuJiadpuAQ1KKHJ/3cGMUZqQPQURriB7+Pedp9/
D4KUHg2Foyi84nKpGwQzbCInY6t50AGcHdn9q3igrgzH5jVJnZWkqbZV10EhMdhhGvYM4CtJJdUV
B7punruLHPpJ34Woe1PfhFm3Sx35mCDRAGo3u7aNq+1Oo522xubYWR0KowCUIVYceeOhpLwoPzT6
qrQmnqKU8cKDF6i4DcPGdYe/FbMEKsaXbqQr+3j1OoWTHA2jR4R2O1WSLVqdqkIcIxH/VvCaFx8P
66WKAN9a+qAL7TsszyPzxit3Mi69yDmQ68pp7V6JHsKR5OL/gcieR5ov28rwKiLl5c2uXsSGEkf4
iS2rtERdKiPSWQmqcI0lAarqVfUqXMc5RJxIKnqwvIUdyo4XPOxig2G2n/Jky0qWRmhvBBd/U3b3
LhEo+MD4oNeyq0kb/AP3hUIxAyaM7DpSwdVYosD+Ts/hyvof95GUgYztDyMaR6Xr7Bl+nxbOkYFX
l9Z1u9luZ1Qb3hQyRz0nazt5KedRDNPYATrUbdm+UF/6jF2nE0HzBsik3EyH5nFZzWKckWaKZPrd
MP43aRpl3xS8AuoN78pTzq+DLHGOHbu1Zx8ds83G+Y2rZy7dwvXtVieXQV5ofeCkQAukN98Z+2gg
eVJtVi4jmL/Phlp3N5IRbl0SuwRZrCSheAMNqlGfj+KHFV8D/y5WcKwXEGjadF02hnEkFk/QJS7x
wF2ZAzlAt5k4aevtKFMdKLrGBG8N+zxlzCehMHbWtbvZpOZQpvEceEnAF5zzaUgoLd1ZaaXtEVSx
Sjy1Uilk6nveP+emd+FQYgVihbq9ILrUn3wRmGSnSHyrtGNUuyNuim8Yd2u4FfXGO4GwwjXuBj5j
DTPi9jCIMW2W35C5BpZFQKKUtutadgHX6ETDzWt9wXpMp4EZXSjCyigCNk47xly1n573C0tj49LT
oNjDpTN7uNUo/bTATMKMqc9GhqX8mhvLw0lKUauRz7iSaggswBoZJCkSFBCmZZEW61+GIafyfTEY
bwrOM38tmcItw+XUvfzym2xwzwVr6nloemWOUSngtopZxksBx+MeX92cpxAEDqr+UjcgROuWBvI4
Ib83psRGP90nnGISqYtY6TiIwuk7tOrI8hHBbsVAfpejOWULoxAVWz3ClCFu5toWEkPGII7z6u1/
+72q4tJ3KR3OUegh8XqrL5KzHy3oSTTF2VjVXw1woKoo01atvLrp1WnbKGIdVED/hT0SRgS8JtHV
/Oiilu0a9eNePHPw7eLfdiIDBFr3Jd6hOxN4WRIgoly6aP6ilrqeaaSza32B3lvblGppxIWSL+xF
wdDbk7HADURo3M/kA8jgJ8DkyBbIdObVWPxynoii4ttyvaw+6egvL+9ADxs+FCAA8rOiiLgYPukD
hAqMct2RfePeBgoYQtY6BqqW4LJWK2SFJb8IzEjOLRAtDDYkvlOvbPnBIpi5eTda5u/JHqHAc9y7
BqSNdAZ+Zd46m+nHU2SEY+03f0Cg427hfsTv555T3JyRAibOO6UMnNQGuLUpi9Z/8SbHk0v9iMdI
xZCSHFwioPAsqDy775Ts5nHhHZp74MvKl96CQP8PSRugRy4aIo5wQ5GV9+DbXpxi5O9TK3LQZl7w
DvKtMOdhvelZggY6NIiW5Ee8J8e2eY0ApuBznHhAZsxVChxU5sCyeinTDerzHZiTABohoHKaqgKu
Se/qpI/kmiarY9ReP0DeYlTwSH6+7uD95tksOFquDdP/YRIoxNKXKrs8WH/NFuDOXhjW5sLalAUv
JMnG7T/E4ReMXY2vspD7KvRIUPmluilq2Q70OcH8oxIUrQ3MZpiwzdtYU5PDSaWyokKbwlrtN9zO
U4wYIVl6tcypsq8ZZGDg8/vkwJQnpTP/Br+1cBdvKyhOCnGcEOLI6sxLC2PzY19uq6XzLReyrLOi
RjtpM22uC2EikYQzLqxgZG2EUFBekxP9enSPkNCzHiiqrH562HTGBPUuyiAM0r+TXKnVAQ+DII9G
RcmtEyIboobIYsOziMYXC6GvjmPmrlFdCDf5Wbgb+S+DLb8iqWwOvrsrQWj/kXHHN4RhjL4Lj3pG
wK4qscnXwDFvp6JoLG9ea3TmJJq3gmTXQ1JbzNSN6MRHWR+2nfyhJEWGHytmhHP2t51PZI8RI28f
rczlmlNon+cScxNafcIoNQAFYHtw4DLmlH/fyjRV6LQ6Xc4etxe2ZSgABm3uLmkFuWmnjh83EoeJ
CvPWh9E+2+QF8752za/MdTX+Cpv2u7gqXZqyngcdTrdG5iZtF2rRmJfwOT3pxMgF14ctQvH6R33z
8EySbwn5V3wMZAfEwPZrkJDsFvw2q4lvI4k+jzRb1pIxyi+HcyoRi1rVtuep9qrOz8jz6TuPH7uH
x3UydVKY0txqgegCqnqOrWfcXkdhvAkHvD+EdHwFvswKHzQD46Cwyxk23lTiIzWVh/kubiQsCBbw
IZoASZD7KU5P9sGX7p7/vJ7tr5jwz7JXjNhI99fVO+njLNeaMcQkygLAGJyxDBbWEUHYVKBlsIqw
woPpHAbnzxu9V8nV1LD92BcNwWBH7w0c8JC7fiXpTx2SJ4+oemo14akcjlCwJz/fbWID6196igeQ
QhMoPbsTRpd2w+0ax18tAv3Sq0UWwwwHEHATLlYFCn61c1D7y12vbDx7eJEVsTfu5iXx9lbTjuHn
QKucehBqDrBslCy76mKLOr/+DaoiChiiUeJPEiDF08cM0Xv5H1Bqp47fihGl5WLcEMLntYq6P09W
5nk4Ko/sRQChfjowUUPeQ3cm3BOto41uJyyEAQNvY/+ESpxNHe38UeRaaB2zyS1cNOv/oa1IGAf7
Gt89Jau4BEmfamI1MExOGY81UAZO1NO1pxBNqmMginYjWDbDIo7SCgslXAPBtI9JivK/hiYUpTKC
3aFwU9vEKuJoA13q4tlvp/NSa1WgVTtbNV6C+Q1XOYuV6ojDi+amWgSvDLVHNjKxjDvgS4u8lgjU
mCYJiI+3bjgUYleZYMq7Fc5MydlucbdtmwfDXsnCUJhcCxpKkJEe42171U1LM/xcjiKnqfM6ma5r
iklmiJrAkyejnGD9+0OIp+I+3iiVvbwwEF0Vr8IOuTgbAvHCRipSjaokbIp2ANNJQnSbRrwrNLDP
F49Qqo5/5H7n5sB0gylaZNy5ge44W6LNvGIwMKtBwmoSpxw95UQOUOcM8UWaVniOHR9YTdZSFv8Q
zUKG46sRgsQJtEvaIbIca5vSxrujW8n5i2WtFqH/Vv6Pnw9xbr3HZjHCRQrW+tLtAnUIaLoFd5sl
QJ8237X12akZRtPJZbJyvfIMkN7W+tK3BiyWqbqFJ+CUa2MU7KbbWzxTQ/skkO1hTF2WfiOr1b99
R997RDxRRViVb1aAd75LW6iMQRY+Q5klgnjKWtm+cZ679bOdMkOSxSLuw89ai9i/v7eMWst5PaF/
YZfS4m81inDAkhCWoz4llGSIJ0KSGH4tSn38j+MkYmaAOYt+hP8T2coF2zrGbSmH/UnU2YLYJJnn
QDDT2UaEhLgotaZRteRmUnuH0+KYen/F2F2F8N3crga88qssIsurRumESI++mLeqkQ1CY/MIcy77
1S61p0NowNilMAHpbDT/nQlaRXEI28yN0BtlhrLBg0mhCx6SIShsqvOhA5kvreVTV54DBHICAtxg
0DGJuKxcZ2i4Z3MCb/OJYpDkbdUvuhIJY/bKjADik+9i/hreuGj3x9LV/YaZI/EWAq11SCjMI7HF
DZCflWEFrWWDVXfFTOHhk21+LhxrBOm/DBWnF7KjhMDkkzbSQB9HidpMIADF7uEgvRPTdptXwp0t
Xvfl6lsTmEdUbhZnfDUI+lxKZRhbakStwtE/piiMoI30ZSPOWCjQwMmPw32pbEPuD7syHKrt4YdI
BgDyouVtt84e/Y0WgcKBVen5TF3Tq8lV9C/RBpevKewjyQwwJ1eCQrFtv/88IgG72CeZvkgVAM9i
BgBqzyyTWoLF/1Kt7zMfZnejjJnODUbrYA4ZXR9g7eDq9fwOw0kjf421eNTlnLTrS5h7F0VKAOuO
mTTuvUO4L+mOQwDQYrhnmYuitDouHRRvamcUfhTIgiRmv3/WBAsbtaTxqQwQwcrJ6zi3gfgaL3xL
aMl5jkAoJumI7K64Qgn4qfoldr+gRm0X26etZpVj4FQ8EygTp5xHVD/JJZreCIWQ8YAi2fpqcQ88
WnhIME7VrXfLFdRetsoDi9vEKUQid4bx+N0dumsGy50b/jk7UWDHVeJ4/x2rwz6zHgekgga0l5G0
oYUWVmbjuaLt67QTZ/fxbpbZHT2nt0DZDahjQIeiUjuXkQDbTQl9IUGMMIEd6YVPjm6Cp2RC3UA4
MhPHAuC4lG2UVZku+eOLdzL938oLrH6nTZwGIZ0Yd9clK+BujgMKwWSxgfLMabkX21GqjoxSoFsS
c2A7KTm/so2u3a4/FwCEdG8oyMRbtW92I06lK00LkcivZmxmXCEaw2XX0Qss5TzWBOFYsocOu2RZ
sAgs9zdFQyIlXgHca9qZYfJq7VaJ/PFMeXLsT+4HwyqczcnzKRqWl9i3Gl7FjGjVif40hE4S36An
JSUjENEtR/TbQsXtca+oKuBr7Tkgg9t0nI2escwQGKDDv9UfUz+skCzmlz4S+s3ibcaaQCGg6Yzb
vSiVAb2dxM34DpXF+IH207d8GA+YrFtvQNbaygjXHVhsBrIDFz/u0xaDeLD/+U+y5Q0DjSAdsK88
rMdWJNadwHrBdeKumG0Y/vDgqHYDxX4D3HRtcQOl3ozaQwUXf7/q3Jz3Qz9bPFedTlA7JjolNMHP
0sQNxiP4GIPJ8ZcgHIpN6j3NsxMrnEYH1l13Dnd0tvflYzR7lY4qShGD/LFN/Rmwu/3kk6vexzPZ
BKdNiGZCABqXvLKt0ax/VnCziAlPhHp8+cLGL3ktpm6GjeTOauXBi8f304fmMay8hyBfJQBxgzTb
NadNyCSbnimDxXZVcub9pf2fd2ef6FYSF0BRDy8wHwT+DVg57PVy5+h5w8e3VUv7MujBkjVVM0CN
kY0d6cHhZgcaZoT1cAD4Tow+tAohKmnx8C3bdHfcfMm6j8LNZj3YLaj2DU7UjD8YxMcluTSJFYEm
mrWCKPdNvwBdcbydPSZJ84fQc/M1bvqzXxelB66JU3aqVeso0/rSLVE/u7nhkkkygXW/esGh8G3r
wd+Gzs08bv9dnl0GSKqu3q2Hem60Lk43jHBA4RguyfGor8qeOYHnQDGL6CgXZeejQ7nlBMfPxpeZ
FeeVvd75dwuGsWsTcqIvXCb5QbncTaN0QS9d3CgSgD7ETKSYkLLjV2p4KoMzE9qJSCThRMoGjo72
fcrtbQ395N3AVhtXtI+N4ElKBbeiBxwTyPvcwnaCC/1Qi4lLvsRMv/7i7O8H1oibVjFpGHrsTQ06
meN15BdbmBWC8NDFcu95GEK7CiAcL0u2WKkqB/LDyxrdziQdxQBKnKe9El2LyDUSzuu27lq/1hNh
QIhWD+CSzrGXVTh21pwvjUC0SED7kg+o32f2mdEae60Fjwng/E3PQ9Y5Qi0V0KM05WbztNFzC9/A
VB7nRtEtxkT1wd/y93Nth7PYyaxZ50SZcxxzAB22zS9LHDLxfBgX6HRl/NctVwi3FArn6CVknA87
9JZoRS9owlUXl1eVpGifSmJUfpXrdBn90Bslw8IegL1T0AZr+0TmB5xkINE0j+XpNf27CTqnPtVq
OCmHKWaUI72Stu6eQ4o/S0nxy4HN8R2BdRrxl9DI/3vWR2tDV2V/VntmbUt//eICeQDp/SrmpMmV
PIlBM+hxHun+sX4NKASYM5D8+zlfsOSa5GsqXGqi82HTpehY9WnFvKhyOq35PaJHqAA5eCAqYkE/
FP58SaTiNJ+gbRfy8oR/HsHka1bAm5FIjXdsXOuFcwuYvhaqGcftdzkktnxXwhsCdBlYWcmvYTgB
EWDP7FHZfDACuWhpQw6Q0EPyqBc7DDsxkUObwJyfOIsPPlC+py8/78fVFlYQwg3DweLBvbC4VSb3
H9tc0M7Dpzu4iwwpk1dhBlUBx2Xh39clkeaTgi/KfdlJr/3Csk+gkNOdGmmI3PDkpkKNFq29+Zu8
uS4392fdVxqvkIOXVQXlx93K63zauS0B8JznyAwftzQKLSVpZyIN5Lr4enDkwaQ11v8FiuwCCYUR
5POH70U4MZ2/EoHcbF/GY/JzUuJHg5ofaoUUqvVZwCZXQgpxGN5NxOYRjR8YaHW3UPhBLw3IkP9M
bgYSBoGj4DPpkmmTPlsbtayouv65VKz3PCx65aOuTMEBTTLBCNOeI6n8MGheWSS44r3XYQq81RLP
1J4bF7de/mO4js/7VWHoRiJfme+z1J1dCo+r47hN3LqykGkRaOZrFnaSGcPJBWrYU+Jt/VS5O7rR
sE99MFa5HM/pDeJbt3uSAirOlry2h55h0y5foRT+Y1O2pUZj7wys0xGOwqLcODJGNsJjeZ1otbMk
CiewTgROUpem/Gh2c+9OGJ15nr8//EQZkZJvvKghrZdcNxQy6V+OP3Igap2aHAxg/c1pZMZoRamX
L4PmoWS0IUGQ+WzmkF5RlL3tdgwQokH/sdXhVnTY6lUkBBhGWXn1sJvdOlLVn3XYjNy1+ffujm7K
Su+rIn04i2ESkn0wW6zRE42L1v/4GHGGVncpauuEAIylAttUyzRXlWdgHQCOYJYbSNm1Xb/NRwvw
yvEvFgFkrB/SsMrYAL8qXkTaENWqPV+qFkROZnZx08Z06xlxIaaLGa80kIsMTU+iyjzkSJ38Dlt5
nlB9E5Jy/UQUnB4TNnC/MigwBmovALVeqQZzuByX/Dv1xhtO6hdzXzZN2QDqVhpVNOFYDhVOVTDP
nHFhxZIZXMzkscrD6rptiAcbHyjVk2waBUcmKrM5NTMC6PDVWYxzwnUVZBMuoRCDi6zXeyD61Kli
QL3P5Ucr4BX/Jd4Df6m0zdyw7tMVmhmzmz1+kARYdI/ExgQiijows92nsh3SD62vCqswP+S4LBns
6TLBXXDzF4lSD1sCXzC5YjIQv9vdhC7kN6yRUS7fF0wPrQQaqhvyKBSiajk2MEwNciL02QKR8vgD
LB6WXktf/MCFUSGHsJW31tA3H6Fh+jeWd5smQlOYf1P+CmMG9eQ+XnM7J8Gml+OdTU9F8C3n1x+w
VKA2rVU8jFZsRbgO/onkl7x2CPAd5WPT7Nl0WG7G+gxOaqLyQRqrNf8Sk2yBrFrrcXBAXMrnrGVf
ZIiI96nR/oY7su0w/Y+KL17TY75DEcvU2EDm/ForasB/ZVFmjoVMybIxZRfsrQh44JlmvLYmaS3x
2eVAfF8Qwb6hTplqvxdklG9I/HuDgRTB7oY4qUQegKn8qzgethRVa7zxsYDzS2Btp6QjrcHZtR/X
tzc5ymn5dFYpugTGep0px8tuXF+hCaKYC7Yiv/oyOE1poj9gVp8Uh7jyB+ox6Nx+6Yfv6heFxtfM
apcGQ7Ujg59VyZU9TxpJN1T9AhUMNUajh2K1LzMDg/vHy3YwSl2UOtF7e9IFXIWNfrJ7mL8B76QE
Qf2SVM/VRyzbXGO6rJvEUgEw5PMndw0gIK0et+VMU6T1f1SCyGuY9B/qOtWrOqAp725OkL3izcfM
nN8Fl3vXDmQdxN+/9Rqpy1Xs5ct8SHsrN4MtBnoUd2uTsYFInCsQ5GCZmVBDqCvFpy0bAtHEHXHr
85UEV4PxvYluMefqKM7XEr+E5yzbHE9NoHyFCnpJqJ21NlzTowOuKv0f8izxn8MMH61dtAL5hocf
aNhXSoOxV09It4F0tJ+h8dkUldhUHaoGKf/A9P5JQBz8a7Do/PMJG5x1fCuq4+1pw+18u50myiK9
MkHN/YYXMi0NhTEROUxfHmVHIgxocbOtowCCcE8xG68LkUUW0vFb/tSFZvaHRb2BiFymAedeZc6P
cywv1aJpgnR3dve6SUWRvCyk1Jtkac0gaHYCB2Oed21OFV96XN0tPYy+kyt/ytCbrcNxNyqW503p
ARs4AHNBU6lzBgh3LL7qPJ5h4UEqf+OodDtUJL+4wIQMF3f9PseJZf548I/gj71yMrcZrvEtU/wl
1VhsnMm0Eh9oszgdi7Tz74TycMovvsvFrG33GAhvt92/LWsJOdl8b1sNmvdKzV4tlg7KtEib+M/h
hLeNcTzoThc9yUwVHe44ZgVWwuWL/sum+KPiB/N3scsnHQUhsGUvZftfv9H2YHE/Q4xrhs0RCYUU
MU7Ofju5a8q7GgU53TxlaQQ0ssIM2dsjnJCwq2QocqX36xtMH/3YfxtXiz1G3H8YIU3cEUHyU5VS
3ZaWzr2T79tgplLWzRFOhy4CPLsl676DJGKbP2KDN1yTOcLI7UTdCngljN4PhrPE50dlFYcT3Ex9
eil1OO1fVAWeLt6OuyUUMde4c1riOJLO2NXK9QpIisPfZpdDZa5XsufJQtLeRDxs2QqkwjjIJoYN
IQvWn3A00bx1/jEdjVpTYlQCCmOh0sD86QMyfW76nGnC6gAk9vv0E7Zp5Zwnd2e+Ba3taLnBZ8bt
gBGXTO+DA1Ci9oCm9zqc6sApAXt2Y3AOdweMmC0hbXPPqwKFFkqNt3pZFlMT3HaWVLGPUURvWFFH
KuIZyjn7lCx8mnHazVla3PdV2AeKL3zy2CK1e6Z/SsZZPs/pIgVgiHhfa/yQvThmT17FtOMveEv+
dAX/H2JGuJniuDUEccl0TY5FV7yArB0Gt41c9HsBjQsDM6elJymz6R5wuXlKXImrbCVoVtIcCoEG
WqRQ8g2n3By4Owh+E2QxMfChG5pnYN2y9jZjpJWe2xUBq62MTA5IdFbtbsa/52rDpZOXtT+Ziez3
TpTP/CGyWgVMEgrCalgyyHYQBPw6qyN2J82Vm2wNrXgL6ND4oVqfm+/vQQBkzo7K5fr7Azon3zLO
myAmXloL190UdHSunaoUlEGCPCER628mtrDtnFgUx/JbBBSgTt+Tvfw/w8uSP9DzuxEFOXYfNt/P
nmYP/ZUmW8tZMtHgVppC3fg/CNmSOgdFMsYZEpDLkZUOsH6eb0BE0bIVreRr9MWFAWnUyXCrtjCx
rDzfYagOU7tp7tHNwN3ifAGSHXvJTJj1iuzpCNT0/JTT0Sw8j5PQrSNzyGSLnPGk8nR97+C53Fs1
bltz1zg4JEw8PXaoj2TsrAwIlfCnSnSTukA0mTa7gaeIeacJxGYvv7Bqap/C/RAKpLXpN5pZ0xFZ
p2M58b0OnKRf+l53e0VLZp1rjUVLzjLf6MYtPOFTjZvMFUYsx7nuUiGxCzpOVeIkyW4D4z1GGmmy
1/YmLPb2seIzlE2BQEUnP5xJu/POhBOX4FD7fk7ZK0RNhpfD8z9OU6I1qOAK96jvERRJCkFMY7k7
s5mC7in7N9F7IXGITfOr5zm4iF+PTimkSiPmq1hTx3CUn0mugHNJGu1aUpYCW3qgzjPq2TFN9t9p
ZRbCWE3vBBfXu3Ol0J8RZeJf+ZwiIUcjOL2J9sIBA+Zs+Rsb51pmaOiwgSTS+BQlGF9C19DGNOvs
MsiRKn7yzjMrm5GizxWuJVF3H/fAwmcXGA7a63VLsSqeFIU0FydD5OwRGGs3Yxuu6xQK9w0bkqsg
/pGMUw2RsjZdjuZIKsXGHNDIUl0GyqqOsfvnggr52rHxtmo9TQdMxT5jdhyFsRUMZ3prP9AT7yb/
lX7JJV1qcubjaX6fVmlK7VtjAinEGLPKJT8wshrMe1hirB4vkkcX8KQBDPDpJxYz6vnhU99Wx5rh
g+jCqQKNlPZmULVcagGgtQ45A7VmuW32HZCYpLsUh9y7R0Fu4Qj05rTt6K+qetPPCD/QHoFZgHO2
2uKOjR2SKqgehxbXQBROfBJz3ircU5+HvIlpi5EbwjAP6rY+48wVJ1BF19Vn3BKhobQZHSbb8Jzz
fkAl9Fim9tXklJwo9MSATRNND/n2Kd+lBytUqNPB1pxkWXKeYO58jK+KJWHXZ39GM7mxZDAdAsAT
bfjqkdoYAp3UxYL1xRRf1uUZngx2FopXhw6ESTRCQ1lmOBA402+OS28C3U/9Xqm1ij2q9a4wKwZQ
ZAKT0TbeSoDdyIUVDThGRjs0JYkBM4IGFaSQ/EuY7UdwmzKWvceq7txRvaLZluQIUA0sin6EzDUM
uTG+yk2asB01iHaoC/G9Q3p5gDCD4Y2ovrQc/2Ypi4cROj57g2OfholOqvl59cCnp0KmC2QyMxY2
HhRtBuwMErY8VmDqJ9T+DQyzaRZQHQUHKTO7Z1T7lkM0JKz8lGlYVDKQQUplM3yM/98pbc2FTCDG
6CBvQrX/KxfcdqxQgMBYhlJoFSzfzW8GTU78jXcuBreE3ZhUkwgGlSV6ZNiPUlPAZYWGPOThawKG
q76EiRIqw6uuBTfeO8CPA6o2M4IF/aPPIqNok6dJap45qOpPYjponqtuQSw7gnXVtbhfCUdSk25N
9IcTkJSDRCaJbNivPeMYJQxmhrcIbCQbFvy82A2Hvz2W7ulSOLACltFvs5niMA2suGdlHqo3DXHA
beQtZsq5Vf7UkRhnPsyKuJJiz/DRxB9AKKsrdlnDeuF8x+vw3ayrR4gBEVNHEql3JcLB7akh2wpp
gomYTuiIBvoz+CREh0ErbERjGGM9n2uhDCqxAnV6mh9oTBPG2tnIg3/9np+7gUFpwH1QR0K/XQd7
ZWuZInqWB8/7UX4Kq85VOgTKvOmUDK0uqNj0N5tO2miWy3nx0q/CxU3MhlwRSBtl3Dlrbilge2KT
sDqsM+X3i8mKK9S/zftt7S0xndSf2gzfpo0/hNfuVKUtbuhjSPaypdi+YMvUgO0figxEOTV2UGVV
0e6e7S9wwA3qpmEdZ/yaxjgoIodaTXZFU2I6HkxZrOEQ3yBPBLVo4u4ZCtrG7/CfNJLjojdjmHzn
aWLetCaQo5MR69hkHGozfhi+Ti9sy6txgAqPhsvkvxr1Qvu7VUBtTEyyKX1+Jn5LKFpNpcgElM3E
EsBxFaljjJDODyqtEpeaDqlaUb23mfn3ptzZA8wWyqi2KEPBHf1KZI4EbSera58LRTZ/dvzNsJlD
HgEQukzNkPZHlrVnWuL99AEUmY/31ErNb/tXa7ve55IPNeuTNFufoFT5qH5RbMZV+0pLE+tjZyQJ
vEgWRMS/P//QRLNGLb0SUGcHCeT2OoGkZb8dWPtME+w2NsBDlkfPwMbhyYFkmCAtAVWKOQYqYEas
UXeTWYvNKUyXwwWrzcLuY4gORoCPUoNsQgeiE0LYaRMprnzf/Djm5HPW1iJ1SxJMpKJO6BRenrY2
yoFjG13E6bFq5eU3NugOmxni9/5F0mIQUjqdTxewXfexpBiUYEoXfBTNv0yYvsikCCHVcmye6ze9
rZvQ82TuJxSklB8bdbYRT3gXlhT2ozcSjvcIaW5NYgflFvSvvT6mWyuI7IH8Ua/YRfWQ4Tdwk634
6kTyvpc6cjjodrIKsFQVV/zzVnHLu0uYjcRZPvP8K4iBn5au6tYbbQ1jguuIwVO2M8+9QAoTe1j4
CT1ZGbVLJ7k1/3DBKwS/VJOxw18v+46ht574aOcN+KmayBdaKmWDSiITqQDl2jdRv2TzGlDLQ+rC
ijmK2SPagOqGTX9lq2ScrkCtqjVhLKYLPvaEq8+TSBfqBagQAfDRXZ0CEqYipwR5HRq4VEytseXj
whJKoorPZmW7u6sbZpJdNdzIcT0oLm/1jxVLVk1UxdSAu1Srq0iQ0chgarcx//QS3e/iwTgBxnQL
VGTtJC1eNsiicGsWeKy2P55op7mjb0zGqxCcV2d5d0JC58t2eOJ5tAH9jMMUd7F+BsU1Q2kbiJYd
UjGPsn5GEBXdaepv09n/cqYt4rFURWSEtgmqnQe5sQ/Mm87S6K5FPCfjawv6NFlDHkBCsc/SIcEH
FM8TKCTkUGFCMJ60En/VkgBgQF9JT+2FlO3axj9gFRjKFxleJQTKs5CghCnJlrTwcyIB12GmzkDv
D4tDWzO2UTaemJxNgeIKw6NxHlFfXtcCjZ7nrG+giCqGL18WNO3PtnCWxSxpnUOQZ2SkqlGGGly2
QyExudUMg7+1pMrRUtFD4hc6qMevr5TuiWqzdPwxkEj+XdPmYpPd4Q+656C0NwX7FqSJ+X7Ac2ll
MJcR/fee1krWoCWcMI/kI7pTNqqeU1qkhekT3Lx31V1lH1sWdtAdpsjCx5XszAoEOTwquv/2ZJcN
yYGcTrIhVBmsRmeO6BEKF9TGtWXubF8U9u52YZVALd3RGwBmM0C7UMLDg7UD6TFhM31B1BrxFlUR
71XaJCXbYToddEq+9rRdhe29VOboetrkMPjhghf6OnuNJT1DwW8HFM6dkj7yXfCJOuP7OQ8o0z5I
hGdsWQhu6JngnTb1OvQ6pHZRX0R9dVVllIUL8p3N6aap06Q0mN2wPR7qaaK+ekgwuX5mvW5339dh
C1I45r2/Uml+1M0TRFEP8orJEw3cCMTezcUYesQuxooECNg2R5Uy3CjMUOP0OiN9jrqnUyk0l7CH
g1/s+aYswBU5GSP+ih1M4Y39OA2t41fACSbxxSS8tTnCZ526jrIG1uDR+VNRCh8WteKdzvJojqcc
6plJk/9sTi210o4uO1sfoRwCax7HCb4igmLM8bdrKzFD5IqI66+q2aUwdvHFFDEXI+7cbmzWB9bH
PRBcwVRgUil/lyBbxkGaOHaAg7PPxwxVgwn3N84GpoFAeiftCVwDGReBSVzo4YUqjo1ByiW9/1h9
9UmTEKaqgla7uGngfvzfWqhVprzGQZIDJ6lNK71eIUPLHSFOGF5kvIGzMCqQ2fd9yyN+yPVhe00v
msjaBtovcG4wCRVBbrcDQKWTKMgURGLY3aTIsFAupti9l8KZ8GysExIrrVn6J+UI9kvlF7yYcDfx
aev7nLB4Ma1Vxd+6BE5tOe/zZbpBHkUDsOiiPajgwjlX5YXUaVPLJH2+iAKnjDgnotYkhP/64Ja6
HR0ej6AOPqg1p6UVeUU2MlyIwkXqxcOIjvgGs6EVdDMG5aIzrnPaW0yjFTc50UfXbiantTDIBBv1
KwYF4Bt00IVKD8uOSIhxoHyUhuOo8/jqO1Rc9l37CCuoEHre4NnJYG+YygTjb4TJANz7LxkmVKTa
4AjTrytuutvK7s8q/W/zEvVDKZep857LP7HMAefBluKis8efBhRaCDMYyCcb5+ULuptqfBREA+zq
zItW5ElXngxF/Op2wHk4CaHI90JSAX95/m7ksixvyJbuqVAqdbDBLbn/sI9HcggxFcU2yevyv+3F
VfPBYASCgjJWHWNJfGqcU6oKk79k8Pay4AVqtHB950PA5pJgsouBHGBdjkVyKtldJivvmFkTv/9o
BKgiQhAVuiifgd4+IEIshy1edSF+ctrdwXEoGy2XTKjFYakzARox6sMbpQIQuvo2inurCthVsFML
duhfM/JIjW2GuSiu1M3GEnV6D1cvgCLt/23qNlWNhx6OVB4K8GzL7tIsJR3jpcgzhhAFkUmZmyGZ
lNmvdhvRUeAkTqXpB6ni3+L6MAMczKuZn+yWjoMGS+eIl4vENn8THSQJdAhiyZym8vfiIWMCZZda
LyUHbyr94uYniom9eiSrXyYi7ZuYPdh6ncWxunGHUOcUCh0udTU00scVsYRSfbRNVTkWvSIyAtyB
dZnJRJv12DZIA/sVHB2tdTtBfw3IeYqV4rmDjjXNDQvHGjSPGpewfWHv6PzRJ8NM8AIyRwFm9q51
0K9VEf/BqBmFrb/D7AxX0XA985K+pT5TaWX4tp52cYGstHGmSeqnDjMuYaY0/TYzPlC6qk2Gjorp
CS7u7KQ8RiHm1LusJWJGKgo4VtlOk/1WwCDsVqm6CKbOGtduxkAwDhyjUrkB8do+fsbuApgAHicj
mqyqGnVAocyk4aBQJa31Be/H34Y/8FcibSz2Vz027gLrMDN9jDkh1y4FOFu4dHpdOJEiXsv4ixIV
38iIy7mW8pvQcZk+Zsj2ZnbqzbM6/ZqO5miTSB1gYSHSb6EdgSAcILbh+7eyHdqbA4jHulDdgpR5
ocaSNUD+39Y/2XG8n5Tj1sn7+IWX0lGTC2RWdmlXxSEgUS0bPfnoZQ0FcTLqqseeAq0bZZ16kk+T
smBOUWt84uhOKIkjZsWEtk7VLH3eJpDadhmAEiPH5ppxEow3Lii+eVAat2U6aeMyOIw8NkA8ydgj
q0rEnbis1eA5fQJD9epdCiJaEp8qW9GEjPbVxBn0tnHLJQI+TTgpB/nQsaCtsGuD30tpq83hvpiP
EhP1oQEWNzoW12ApEMN55JHkmyBhW+bRq99ged8UIxmOnhzip936dmundb4dLfkH38vMyO0oAfpU
HHNa4BLxExHZ5/pb1Un9bTsQU7BQktm8PDVIbedMKY5scaUCRrtPGB3U1AFq/ENE4KxX0MABb+mf
xyRkTwF2vGYdv+gs2JBklhnrMqPuKMfAbYD03uSsTKDk3sz3uYBpWDuO0S3iIX9wjPGm1QvSVOG4
S7tkOci6RKtcRDNshSWl8DDjqGcWFI+pyD7rXJTsanjLIoifZaP0OacXeAoUUO3yOcb5ErH5FQG7
qPe2xvWe8tHHoVLBJuY2DOScrrLgzPjEwRnoQi2javXfK3rOSh5ccibw8aS/SmtQRjx0EEaZFjGW
v1KdM8iVfhIaLM0fGgJEGNAVKsnrHrzQdkSNGGgN186pomODbP/yDFCrK+zx19/4mimr8qRkbixq
ciju3yhUXbFrSRZaFMIogxhdZNLEiCKyOMXVxXjMNgce/nig67zEP95uaee4sqtAyUThe8hZHKxo
3HQstUnxAU5rNYJ9nO5ocgAr+Rphv5hVOMmS+GZvv7Gj3BW8xUEwm1EY7NljOMBENTxys3jRUp0B
yuwhTIGzd/jAvOnQUwOjvWDXinSb/Mm39qCYeVDeFCYFznohP8dk39qUHIokp/K2wTwV7opGAx2U
7REAGBIhXe38FAPkeAVGiLvKZdMgZ/ONK2omwSjYVe2snG6pUe1fN9/OGnlXG5rXryr2Eu9wfRMF
vOm/MbeERS95z/ChTGZCKHTSL6zIe6fxYo7bi3kNdWGZDxeRzgmstl6KlAQ6aaHxd2m+oqoovVnV
teCYM88gXbNeX1sMEDr7eMSuSWrY/94qm9OoIxRisagB/0djeYDF+5GzrXjlnQTEPILqRXpJPIOE
WpI4b3x9IIhma5qYgN2XmxHFGJkiHqDgW2beRjG9dHbwIYA/4ur1iDWTGmszLtBjt/SyaeY/CNfm
ek7DKbhESrtXO5Anr2iZBF4g8u4uPV2J3udcXP2DIR1Wl/4XmfxrZBaLJJ1nq86553XTUZ3kWJnQ
gd8mwY2uDudcGwgl2b0qMpRj2dJ+T8CF/wwUYu/eiO+xdyrlIUl8sACSfRSy4fqm6oB435H9ncR5
o9jqgZu3S+E9cy1ICHyDCDbOPDv3IvSoC6XfpQdq++UzBZAidyV/rU7KthQCuIuh4WV2myo04/87
omfJ6AT7gZAKM6G5nxwjksuAHHg95QjWe3m1q/nwE4MTKyhrLurL3+QrV5byaZHGDws1CrHZHcnB
V/7AIGT9c3yNJ7tDfpwGNxMFJkdS5eP19x7gf0fuSijM1xILoF9VqQugiU5LViJunD0/P1DberYb
bOGROnVwZNnKUiR3PhdlAeK6occWHKqq0rVSRgBGJntXY2NqFx0Ut4FdrXtJNemRX14zkP4ql7v+
ZdXQClsYRuNoi5LnTxo7p67rJcoqBJEGj5bXpV7Z+0SGJ0hNvF6WcvoEW9RbVwY5amMF4xGk0k6T
3iYyFq5RIHUnkJAErkaDBYX3vH/WA4FQ6ICrhrvMZyk3lG73gO/UQCEmQCc/XGYQDXdmjHswJpFz
T9EE2ff21Bw1pKeQbm12Q83OzkCxVMOuhc4ZfaBLSM+I7ST5n0/xHrFW5LaEZDGhcO0aSCRO1kIO
MySAa3JQB4EqCO6M/j74LMLT9maPkry1ACJ3TYsuJZkRd4qtcqtVyqQNR0EKVdPUg7w2nCZXEPFs
+9efNdH+U+7nWQli4eei+g8xeY6zG/XAX7mY//vwGjyAe6AOuC7IS0bnk+Lys+cDKBPXxTkqlT86
RVeG/PE9Q7+W9hin1tiEdzfID/iagE2KaGPx1qoxaf+4TcaSO8l5ZTJd9Z59jEG4CG5QRBiR5sQL
IXTb1BKz/k4AavQ8+12kO8bDREG93jnwEAIidnRXQpVeB4eUxIZK8Cdft78UoNue/6vaVGa7Q6ji
+3nS880kSQe9zNE/GTV0Z7j72/isA5XkmxpgF0qnPle2p394jgBDCbdaSxYoCd4YSu47/2RgRQRH
ofWo1YLRSq5HXFjX3qXlqqLHWf6hpvUTONlHb8s++8B8rcA5nTEcKX1/ZcslrbUk+2CilLLiXcr3
GWBHhISnKbZ2H5IcYm6BSGI1v+qrKEQQnrTLOawi31UeUfnB6HQqjlP4ltczjFCiADGnj3RwmJ/4
/ggxKIzhZ+eeZVqCI9MeqNGIjfxL1kNffKKfGNdKIZJZCvSzATce1vUuoPJvWiROP3w2PkA+WOHp
mTsERnahNEfbZJ6jJdo5XuXGrDmwPWFfB+Cf9i3vqCvUNuAg7PFqyJ4jcubq+bZ3blaXlb3+FQr5
BeNtBhuLb5QuIKCTN2A/9GbWSb13zu1LP8p876irA/tvK3I2vwtFMUgciSh+1LOW2Mv4td+qQfjH
R9w/zkqTtQSO7ErnTvnTdK4NOXv0a5se6AsyAvwgGk60TRhBQ69jE6XvCpUiK+DJ0xqKCmouCEs7
QU1PW8vmSkyB2G06Z6Jlic3v1POWTu6P/vYEVL7JUWYwchi5yiAzpk1EbqC9qgidFnH3m5HIPDyi
6j/bWaRgtlhEsDPQg1apqIMnW5uEatVjtHQ9tUYVfRkzc3t9XbQqGUAqcfHfgsD7k8b1DXLLiaLp
WUTaCxj2FtV1ShXK2TYHpI7VQOZrdmLqipH997ehAKfFwYM5eWI4jiZEgoq3B25KbeHMNRZLOfgv
mWAP9mncGByFwfBgIW04D1xbiucgA4ba2/dhnJhfnMHknbTNWNHJUuTkkaJlEvgz80HXvEcJw+pk
t+qHE7yMLe8WAibXN0Os1GA1WdiaVqzaUntWODudl4s7pIwRka3RS5Pd0oCysjDa0bFRcNbS9CbJ
H0Jvtu8e49csy5DhUF0mAEZvOaChigwEIcLlu0KniZq80mtMelDGAZPo6uJLJGX/SZW0xo/SpAIA
DOvoLKXCLSKfF6tz1dwA20B3RQB57KTgMQ3MUKtMnZRBCbh3iiEEZO+TGBzVCll0Y27jkgvuQyyb
DGVIddVJ0ovh+A4TKAfjLEv7MUsGJURrk/xtIjCB7278kV9ASCcsFKd5LXdFGYf8TDxxy1MF1bub
Aw7VME4cHGM1UIKa7R+wezA5EipXbzpsKDbdfKTjRMW1F9i4K5cqh34a5X9iQbFIEsIC3dHNZZ/9
4NKGkyMrSW2JidmG/H1RHBC1zSHirw0jt/Q1HEnJYys7hqqI+qLypgU9j0fAnyw2CJQ2ebIibF0+
IB66GZxkBSHA58YndFCIfHMqE/w3PH/zVUYednftdUj0Eun5PQB+iWT41xSIjxksJoXE77esU3RU
rBLNpr8PxTN/+yFOG+qOkmFWMXD6C0mrRzgsu7iPO4RRaBNY5VEWLObWDSwGgGL4lWMtPMRf9TOg
I/I0yF/QvxKVYG/NwYL2kB2KpaKGvJeUkgG8SXN6GlYj2sGERe0wm0FXZiSPJ158DcJ9/+Pbwrn8
lEC5HhT7YiQMNrJHVmMtnssSai+N93KAvNH3ljuSFBpZ+GeKFFHkhSVrNrBDedzIH8RhItHIcTXX
DoNnsPu5Gj2uRIg6vkzYTmwEbVYVVb7afiZSWAIulObHbUJqa6nT/kPTbbpRveKZYr+aBu9ptDG1
I5Deo21949wwPjNrLXLLPA5PRtW8HeUvLsYAEcwhdixAP4OzJTXbU0yJ8cEWDkmeDi0q82/r1p+P
ATH2MKx0E4Sl9ALTNqmgUSFR2qmaLqhA1nkGPvP/AEG59t4nil5gxNkzCxE+vXSvIoalYuA98a4a
UwVO11IfY8WfHuC/0eU7bsAsCMoUmGVvP4ZI50pZapKXW4CE5IZlD4iEniVPvcfJqBTvUPdJvvgW
HhyEJf3GDEJAes3rnwG/8+Tn0+hTIQ+Vn3ARbl2Zv2NHJ1k4yHBTuZp69crVuBrTNkU4I1Lg864M
24IoV1ayT8cHYDvvAE0aEKJssn4N62njAcmAcKIecTl0FzxurUFrmNV6m4bKUyak29hIz0rk0Qej
ngZFKLw+4x2KTCDGXatKzAS13ryC3Q4s4YmG8I17TX6onctBXcz9VKg0KmyWE3oDUAf1Y2AOLD/U
UDGwgAO2tIjBvfddWj2WmJpuQZnRA3DNwgjJDDvF15p7Vq6qktQS7Kp7Ii9Vm+NILdeUzpetF3EW
gVWFyPlnMrrrHST0P7Mb0Clg1xXUuTVD53Di3xMpXfdezIRHy9qMMbI/dfdN9JNpfdIM/+/dsijt
Hv681VYj6OGQ2fN4Wgp3eBuevMQw/8rNZmzw6AWSVsE6Ge0FqBJBOKIwfMhsDNB4dRXQNtSRq23i
3h/0azZ+ae1ThEh65brZrkey3ageIT+J+Vtqn1Z2ieyijotbnp6+K3szHIhLYPcHMUlcRYQtmsKG
RFLgskDXn7MZKAW5LPO7YV2m+lloLadzq+48aRJus6F3RFsfjZ5zTDMaGhEgvAldH48EHxD/kvXw
rBowhbXOCwdZ6Vzo+//GMtnnij4AkRbpyvzxGVk1jR85OKcMiHfp3cS5vbzbfxHYf1m2mBqBg8TC
G52S07sPaNzTpZ8eVpdUbScHHlmGnZQUhOX1+ZJxYJy6IStBa3wbHtc3I1wrc0v3ZS7kcgOs8TTf
zKXGE8Jz6m5n1akiE85rm/JR0x1rWRv+rYexGLZRVb0HHn0JcJX2LpGvapfW1tDz3sxohp38psHe
5OjqBje5xyzYpTBkTLoN56HkrgZYhPjJyzGOYyM92FJu7BC5TUVJTT7Spqg/MjYsjxx2zQVeDvw3
sD2WZtg/bGh9CeEQfa6PDRaYmStkbB2fNo7u9ZtYrb8PP4rgdWZnbLh5oG2UWlLp9iQXfVGQn/WX
BmcBkv2lYepavAHBuBC2DkRTzpKwH0DDShIWcbkM+vTMSC+W3vqSx8f//dmXHJGrlOcKO5KXAQDL
TGFMNZ53QLcccD7dC46mXMWrnC89SVTZtbSsNPn6PSlaMJJoLdqGwm0hhHRROdG091X7nsese4r/
yX6ytxpg8Y4mdCzrLoi9CSzp5HhYKx2SgFpCdcgA6bP/HH1RBjKWQ0r5W4VisWM0y4R7fx5kOtkq
afKQt6LYucBWYguezFjshxPpaxSbo/UVOtufHkW8IWz1g8ce4ct/jQ0GwghFuVbD8iYFHDB+ZdiU
QNyuhsbPbwz3o2Dl6bEz6S71xarS+HHM7kB4wx3FA6RnUu4jz5I6ky4Nncrjw3u9pXMUzTBW0m8X
Uriq+CnetDB4ZuOSk5gmnomjJsSpY+U0ClDq5YMNQdhQ1aegs3gEtc8U0keh7QzIxr6gbo+Jb2ky
Q65o28B4dJ9s2MRDXQisILlewuEX3zdwZVEDJb5o8yMZogtsoXrCsy6eSBRIHFhbb6qPtBFmezRx
qZAuGJgmpw0NPLb1vVvQ+jWt/RsRvRTU/eVlUw3rJI6bjpHuoNn1sHGFw9y1nJJFzRN2YQ87K04C
fCda4GCS8sWOh+yzb/N8BOlX0MNPrINEkxckaYxvE6fatRRFyXPYwAPMAyjn1GFQGcgIOkeKc/1l
UAsNV5pq4ZCXiUyYv4ZwNPnOodF4DWxozTFc0lG4rjmRWudZfkdIPuxFI4fOLiKjzfFVzWHgN3hi
JOP1EL6Hh5UIH/La0J7j27SoNyS8sBy5ccQ4Ea2BAy6Fr5DYh8rskKhTr7JNS6BA6vNLeujIhKIC
9hyP+FngIr5qAnxYvbHWf/DJZjBH2RN+YR8Wtuaohj3NuiO1Yp8C+XDvvU4XN37ds9UquoJfc50n
cd6vJ6WfI0cEqGVEGJe1v2mqGhrcTdf2ni56hDtBBDRpXygk6sWdGpnH5grM9BZENHiogTZDoyh8
spc00fdShE1f/sXaLYGNf9HPNoRP3U6CvWFEZHRciTe58ivZaNr/vRrrOvVhARomRXdTJ10NOXwQ
5TINNRy+I/skShOOK3mAZVt1G1P9s/KqUjx51ovnHVpyuba5eLs1cNmGZMOL6xzBLn9xwatT5Gbs
7saYrvOW26+vWYaEh54/Q/VCHE6LZtVX8E7mrdKS5VtIMpTZrSb9bS+nJeCVTXahtFeFlmQPXPus
PfLUS96px5VlOYeDrVzdF/0y0gM03tNFCGFiQAST3p0oZRHIn6bBVcG8Lfuc3Ad/0bUtysLjz63D
fHBIeSPV9/aNKXQquMCgcK7nF23p3r0XFWKheneRDLyRDc/s6x9/0vCw0fTlBXDe5q7Cn3vdJwhA
8Ga+wspsr80EWb5hF+EDyG0lwtRyqvx1iOcBqdOhmFkqb35ZSbP/PaWQvyRrNg/wKmMRkmxb/cC6
E06lEqmNde+07DWNRn6ash+NeHApegVxM5chrsaPRjSGB7c1lHMADJEycVy4SbzA24BQZV3kcDtT
CUJRjS3NHMPnie2IrKArFNSYALxBfZyqGo1kjBANBqw2Dfzy2UEYqTsaCug4JFdwPaaA6POywjgT
LdCWCR1zy5n04uSyQvRVxnUioJn++7MzcK9WDWkJUS33o/b2j+lfci/1Sbz2gEvwI4S3EjA7XIB0
EOH73vRxxGfvVHWnszL/AGV6RFv0VzgQiY3on+pYJieLDkhPz0XaqVNaStwf7iY9E7viFz9OgwXc
rZh6TZqP7g5+NplqhOwBViH5IYN1Re7MfIFVqjophmKBLqmXyGT4y7PcKH0UpPNn3dRSpg5PoBdE
+HNHICkvjoXFIIo1nZKAgOUKPZRuXokFJBfOWgKJUXhnL19D1s1K7cXkIiHNkIsABf9VjJAfGma1
IbFoPcWGSmZyh2K6DfQpBIZurdphpUHkKLL8MTtRTNl3XUCaA4VRFdr4MOcAFNhrPwGDfQlaz0Qg
9007QmY8yXhN9mI2rRr6tR0r76pQSrEhSqrRI8K88QxJRrUfTBVTP6FjJ9xJWGXqEcUQBtJnexO+
McgILdgv8OmqEofP80cTAVQumN4IwBn2AN1CzqRCScxqen8EkaNcfHTidlsqZK8aMhgtPs1cJS6Q
WBswk0ivi59Yn6/axBNqtNUlFDi6g/bPIO4oz010W4MoJr8mgusSCjgDxUUQt+beVNgg8+eTaHKO
uhY8XNciWuyOZMZVyYti6K7UwO/TYtVLeVFkADQ4tp6UWfUfGk9IM/pigCvycuFqvjrsXCSQ1gen
T0MxX3mQwCOP0NYj/RY3L50uAc3uQ5pjebfEmY3bKKidzcTlfTylHLkgt+E3tX+u8g4k5votNPl9
SKpcBV8dP6spg18njCAvkHwn7ArrGPb8+/Q4kvM17Aqqc0OELVcLWHWc9GEMr9/2u0MQaPWrtYyG
wMMIpNI7UmDxPJbNy/FHGhoHZpfm881IE1usBitFKF9p0dqgXmX+1Z3urdUVeFevpj6tOqguzRJH
6g6K6SHOmbLANfHM3R0BXNIA6Ip4I3UNMP7tJTLK+epPzKyRK3nvco0anDm3hkHsFrb6clAlKd9n
fLg6Lh8J5J9SGq1RpyOKpENS1Y0FIIOis1H6jspbVPYiVdk0pBE8D1bih5PaRB2EUqM8hD1FziFI
H6pICX3G2Pfg0AQrIo7Rv+ZMMIzDq0LHTpJW6jI4mFTIlbqkPW7Wx26QLJ9AvOvGg+kxfiJ9sGqZ
yg32L1t7sm3qDkQIIX/KA5cg+FWdr8ktgEWo/X0Wpt41VCOFFvJDDiXN6bVQS6kXrz7v2fzVqeaL
2EUd0BdtkRx/fArLm9M+lJfOEpl2Ph+GUX8tb107f7SzBQOwPILZXOz5PPJF2fYCyg3gHKTy2vP6
ikm3GVvrXGHb5WvI0edCSE5kcEDsX4PN77pPggnuCAocrZx+/L2XWL/Xs7MvxFnjXFzyKjTBPbYo
dZGtoI/BJ868X+1nLHsWW1YsRTkHdpLi8XaAlFbn4NqwEqHUOlIO3XeYu6XbVj5Jz3EfW5R/bdyL
ZdEIkmYUb6b2qT8AqIAkfEWH57SzHuODYNaXkmwC2pelogcjZZe26VKRSkDHHPDLeH+EV22o0BiV
8t+oPplExrJceuqOEjaHUEFJ5uezyqkTaYFgXTIYJA1627kBFcEgiJ+r/Zg1kkbVjJbXrUuV423B
qyD8TLvLC9HbhFFdMXg7RzSFImbjX+br6jXcWcRPqLI4ZCqrYEbiofDGpcn+lMzHdPI1m1aO8ft0
oirNJc57mhvY2EgWTy1mRZc6/sy15uTWoXn0hM1tTaVoP/ZEUggQC0uIbvvFTJYuynb/8y33JNmA
jfSQTWNFxNCGRVLfYnKBpoXAGLNQcLcOTX3PoqLQxhuT3ZD1a8Nvkdz1SocnJuhTkkG3emPLXstM
BikGSLskQ5AUBSz79EOeLzTxLm6RyXQkjZTdl25q2JlKijt5R84vLhj4LCoTA9XzXAWJkmZ71XT1
FozkH3lw7beZ2CJ3eHKVLL0fPW2CVczQppms68Y440w+23vnpUw1ga18JS6QeVKvMVWrED7fBuWZ
4H01t0Kz62MQTuBUn6ib/PXu8/IZpAtPZhzJa78kDvMUKyaqyakNpU5y6uImNn2IRxPfFdz3y89q
kSE9uWS39gaLAsKHVFKGchLKXIp+2ncAZ2cwYnfIWc3UnZlXNhbi+9EjVjc7DbSXNQYsQGzkrBVi
NLkj5kLPSMDXjXlGpaijDfg2WeWMaVNG28pTjeU36IuUV8KyzgOe4CGKqMU0QgCRfk7DruenjERM
/sJw1LR/FShL1+V3/FpcgymlzEC9LTeAteompzpPhYoewPw2guQm81VcKdIy8rwbkpuxd9y/UvBG
TVKwONAam/ONEJcjqfqhBID7Nvt4/Q7ZZUX5iv5i0qW7QoWRd5udqurbWhT88tEEeACssEZy8P9j
BmVIHcXSPm/gFyJfw6OQKL0cgpPWK/zED5E38px3og1JEMQ92LsY2iejTXTaqRWNdoJJepbrVyJ2
xmQTTskF/OlDH2gtD+qwLV+Ob2Ipmqo7ooYX9HQ6C+KOI3sv0lCtJOgNYI6XYrlaCCgHkTIOF6Kd
vCrluxWjciIAXpTkQH2OZ/PZoW/+DxJWLqhzSOL6g5MZO8yDCytLOn++qj0YP0CMpWU1kWvWYreq
jIq1YhvTqop4Ck4guxv35wR6lAdGD+absq6oXyyc6JwXJmRoPTBR0WS3h83Q6ofl1e4URfC4nJ0+
dLhfjMWorqLRETiEuV9jlAsGQzWH50xssytEBxZfyEwhZJ19MLS75833QFat+xiktrwknBeFFgQP
cg/D5meV0pp3QS068G53H0iES+rOlM2cUyv8MB+ANUkeXCnsWXclUrkQgKOgpyeI5dbq4FumNh5m
+f5l3244K5OWlB9m2n6DQqsmtL1ZyaW1+PvO+7IE0wltMG+qypDfRGwD7t7zsZy0CE1hfDdvgHKh
WKvMle6qaMX122I+Qfy2uHUqjkFtI/hy7e/CK9M0NEbXlKcDS+2sSMMX8PfjM0p1M0yp/dwynAWI
w9UTmrTKmwBgJxnwq7SCi/h3ObjH16xDHRBNZVC/Lxj5ne+0aYmuv1fjU2ILicrn5xoRbiQji6KT
e1vZGmMnpY5sRTGtEmF2IpPf9AjmYhR5F5KEYGpDj5XzqzxwwWPQMHwuU/Lf7QZq00X6WRwt1Q4h
e+qhvJTA67BpZ2i1rEUq2rJX2ybv3JzTpK1CBsWZR16dKao7eEgZLQ/yzzkavFMMBSwsld3hMG1t
4oChQSj3IFE+QyAqMptm5sGqBOcuNbng2+NhqXOvFM5uizORcWJ+0twzeqq8kqn6doSXH0jF7PGE
uZ01zHayW/pIJ54ALrqTyRIoaML/APK4DpV80czv8C/3uDyA4jc97Lsx5RFGuzi1gtjJIi+lIOoC
P/wTCIEI1DWn/r53IkaC9/GabsvtpmMqUEQtH6YcVDyRX6oarmrJ1B7EtlyrNVFx2jHl91T+plmw
hUyuw9DtfaD51ZqFFzwXFZ2P2dg86jGIgLIOUUmvEZ02F16b6+PUmMZPyDlBwNiuStfzzXIcmILd
VCNb9MYZVONhnmPmi5YAlmV9nog68J6KmheWWIJG9uMsNsaWLVswcXg1ablwcWD8pm0Mjm9D/C6s
YFacgdwkYqc0j+PlIaN96Y7/O2syKR1hGFeCh5ORFywiZE9+0d1YtFuOhcROTm60EX7JlPe0G0m+
pb3zTFKvHqOWpSj2fjRjUbeTiCRZ4IpnRbEKmMIvYwpFuN0JGH+vUZ4g6x71d0gkuvhjaN00sKPJ
taFIrkgMbypPHT/8gzGiJp2dl3dLwFwU0NQvYYWjwocw9OS1ngaiiefPy8XnTxIqylfWnb83YFfx
ke4jFmtnyd/5hbP+koSxnd2JlBdvuQOD79p5AP+Wy/3KqRLmP284hB2Dbh6Y8e3hcNs22ebAZDNl
cN51UhOQ5et4lI5GCZU0vckXSdCPaYR7z/A3gc7wNqkdLxOjY2dfKlo+PJ+E3Y7oJLtdnJlHTsPh
p31hHDg8d+6ys3jQIyGNDNMIkxp8LNnbTT+r1UTUZWlBZGvCaNrx6wz0P3vqjRbwDV7N2gWZWyXH
zRmFg6j3OhCI28HwRrdGV3IhhHcjUz7AX0DunTxjXRGRP8aU6WftTsSoCgRiRa3GyhjQ6+wZH2z6
2K8J14uUtzJQDlEjLp/uxB9zxUpNSjtQBXpioTBrRs23j54pdnxTE8Ip6nUjo3sV14Y2gnj1YHKW
W+dvcDdkCE7XuPFVYuGJM3gKiKLfzOM7WNmHA2QGv3Slhs0Sm3miSgq9ArlrUPEpxbCWixSs57oT
0M0lAmFD8Y4u0YSa5TQwW0VJCAR+97mtFUsoylogP4EkrNiYd2aX4uGsDLRvyk4W4oRYUxIE1GuA
Y+g8uhv+TA98yIE6GE//hAyao6myLymBrgE7wVTKQln2xrdrcVUER8HXndPIZJsQL4kxu1IiYNo3
M2jfL63f/PTzpKroHvMbi9rYCPVDhdNQtI+viQKn869Tqw410IGQEoBq81jn3V2+hOTbtytFWfPT
R9WPYnRjj+xr+WvlG1YElujVd0r3KAVU3qt9OSbxBb7Z/O9r6JWego0O2cY5lQVQ08QI+wn8JMBI
yxChO8FeWRXLe6IEyqO5yRpSTBglOPSSWURqG5Gsq0ZFb3KP3jfeaRiwd0C4CjPu9p8uIagxvAtf
/38zqBeQ6gwS08DPNPGD5m6ZIFgAnIjFI5Z6plPjfQ0ZSEAujzckuTsqb56tgGB4i54A/zlH3mMm
VkakHFR6DUmwqnGdblJ1P9H+lIgLQtM30vF3rBxsbggbULWHhs8+2Aye9CQH3LFGUoJVCT4en5LZ
OlzwA/evkQjUHs5rBEyZsPw66UxVc1yz+uTVXOPa5aXjCpojH6473euLqykJtmie3HlnObs8GJjl
1/gz9i/XdqI+wiXJ1djL2nUXNV+Lu0jrZn1gTIHhFKCgRY/RNUAitQp0kh2T6WvQy6S2qu/N4ePm
Ww/IB/NuLeroJ5QMVp96BLz4j0KZtgv29TH5trLSG1numlYD8aUDBfCyW/UPKd68RvTXhM0w2UH1
9Peihz5/Z89Lj7asHJmPgUeVukqH3AeO8EsDrWh6y8DZZVr6U5Kgc1J3f5ou+YK9rySK3uyE80Wk
3Z6QYqxmixPS4B/bkDjZjSVm0g+vOnb8YlK/tifgdGXhYYLCs2suHGdm3y0+rK8pTWR28vW0JIKZ
HiEPCWEd5e+g6xK8g8oP66lfMkzhAFK+sHPeon7W+x+FzdcVaY5NUu0L+LvK718a2KbauRC3RyJw
5WbxmRofunpuKMa3dUcAsXFttUg0f9BkGLIEkscrEuQ4kbto/j5lbv6oe9IQi5fOQRu99j0pZ2uj
hVLkNaShINGfoRhPaMH+yopKw4rXnMwkDc4VTPDvoEbukAcBE2sEDv+oHs0hXo9Q1t93n6ebGqoh
9PaFPjtCHihVcVeSYrroBf2e6ZM4gluQTJW3Wb0Ux3xwnM6+edSiMDp/Y5gSZp0Yq/dONirz6T5H
xcHdY4SAx8F9JsxRenVRnNto4fB3oLriNPt/lsUez4TzN7LaebGvdcfsgTeTDXBKfi8TkP7m09+y
i1OUPotzVP6sSAibWKND0Do9dERxjva8drtai264omP1hQL/aaE9kLvpj6qo3wWwwuGQxeXwhoxI
79pfY0rda89bLdym9gt0clxsDT5Uxf8Ra31xQoGaOM83DlhwBxtZXQk0/SOc8Mh4kixEuL8QOAPC
rLB4YVRmAwPGjq4Pz79oMPOelhLVToEQuCE5hgmAjAQfuoulah9YLil3iBOwbqvWKh5uV52DhWgK
H8vAPRE05xSDeavBeOelrG8JpUlUY0e9kziA2WXHwDB2R508Qp15pQx6RMRw7muM9NFRJVfjgsJk
8TwRKlAVmXVcgWymSeAcL+RIZ27nMmzbjeisjHgE2ILfwOm9ps78AE4CakOfs9FbGtTbtneRMk6f
MSDX8YHwbnDRIv7W2zphgDZOxzqn/QHH7BV4L5K4D57WqxfLpHH14dmd5Nm+qVOJYi0pkFTtxywu
WnvPb80cYjq+DAPNst0ViQ9QyeRf1pqoRmDRTfb7HvPQXFRjEqtN+Zr+DczIiOjtiqIBBOpF2R1j
F96pL4qcaHdMbKeQMcnYDPkCKaaAST/Wzw+lAFwFEzfDZdRm3myCaT2p3Lh1dZPEKtHbqRFupIZ2
r2l4btN5iJmI37nygvMsmRqCG6kcnlcOyySuIXXGhVwb+w4MPqw8roGc4KF1aRggQONMCIol+KBP
oKtLbpau4W2aPameOyCvX5tLb3ahoYcStNDWMaYZFXX1nldr8p/JRbn4HXiAR+FLPTB8jQpMWwtK
GJWO7YaV3V2uXn0efjDY3aaop4cHIwy2o+AFywE7AtDigwoFI0M6tlYGzpNfIGPxlFc97CrHggAQ
qW1cPQgiGpIIIOTp8jcHu1jpH6zryEBTPCkQD7UsUzONwvLvZ3fgZyOF8OQ16S5GA+sxtRBW6ZXD
1agfqvE1rjSJDjtX57Sa3OH6zug1tBLrCjJg/N/VZGpcu8/hV4yWvrHVeodSKo5aj/h5vC3kcl6a
/aJzn2TSVbYYXXQVTK92bF3ppZrYv/Tzv9WvOKEMQBrdxXI2/xvJ9KIR8i0sirhE+lJO9qUgFKmS
KJ5K7qzSU/aINLPTGDfYfAXJ3R1DRsVFNpI7jrXkerHn0Syy+9iKJKC9suweOZfXnLqAfrV6EXL5
PODSf8QJzt/HDSiueo2kk4wweEDtJucAO3ORjgV3RXfVe4XFdbdDCL8net7QYGjhqtzvnSeSdCvj
OcN0mVm+tA3FbNJsx3sk6u/axmD2WeYk5ar1fU2UU/VlJaqeF4c7ANPZUiU6Yr4PpVfY64zr6nB6
yX1MtUDQLOvbXpbEF5XfschEvsmiqVImTv1xGTcua3uuCnViyzVu+PzBDKk7rLsjK1npPsl8Fynx
Xpf7V0v2CxB/aGrtR1y5AXDerUZqaLUs8C/zEzRqYviOFM6TCvndetAgChmZXu2NpJnEEiRMxZL/
ycrRg9G1sVDkFMOeLoNkrKXDwfoGzfgfYnvfXkddr3+Y8xbg8YjA/EFVmRQMOEb9BcZcEzp2w6q9
DGQB9rKWA2Rv1+rlW118eUjji9sv6gMpf6J0R29Pwi/XfMZNmlNy1zoN8f/uUbedgt0X04f0ChF8
YQCo0Sdn42d6dQlxZktZX3/uwA3bwcvmK5B45muSs+BOlEAXX6jE/rvcjsMgFRg+r/Bh1tv5f3a3
6l8Zsb0rQl61LhEt6Cukgjm+o7Bt23Y3tI8gyf0n15OfC648C9imX3z4F+KmOAOu1vmF1hAY+Dmw
lyLXT7lebbF4+kegXwohGGBKHWbpJt2kzvlCNPZXlohHRFBAR+jCBsqmf5ahfUIgLOFyKgn8VlMG
7WRh9vB93Vb3ykJdBSdcHLqdXzbsFW5R6RvCdv4B3XzVIIyzAs0qDwkZ4U6IVXZgaE2bZ70YFL6c
aBjYuumfaBr3VegliWx/6zmcbNmeqQCz5ScCPpPYxww2gXyyw9vyFGluLDvO2bo++jx7aOSAxYQ4
ytNsUShzUPRCx2k7Xo5046KOCRV4OH7BP0UxCQs0Z5oPXRa2sPT3fPL2IAU0CbjdLQa490UFxqOQ
tGoYhA0V3hejxsc793aFZHSG5u/pPFV7Xo4OuOtxuNzsOfCVAM7QYoZlzNdmkmKAerNV52eEIQTG
0midXR7BJHMGHQrtkKkMrfh8Yf73EmTRdEgRzMuqpUj3Or/EeyvDWmzFqrlwS23iAcz/nRZKfJ/9
KkHw0fBx9eNtCLii2I2F/a6N5DOXM0Fi0Wk8a3avBzo3WdQ3qADLuTqls7ygAtGX+qDIZtbMkgIH
HISZRb7W1twpO5yeyHFL8VDMlV74G2kyYTRHC3BOSMdbapEoBZ3zetIyk2hLhpKcJrcOiqAxSU3X
Ds5Y2/uIZfwGMcShxDa5Nwk0axFmASGoNSD1d32xZ28QIMdvDPqoy5HDXRAMSNIYpl7SoYB5CZKW
zbtmh4BJmE31hCyB10HSLI0s+7Eik5cG+tZHtPJ/7ehXQDaR0QWcHDJsWe7S9aVZXkUfmkQK/xzn
5RPJXQDV7LJfi4Np+GjSGXAOpgd8t0VvEDLb2u5MPm6W+/zzqmMKWh7OygCv44jinxaLfIxNlcGu
pDUs5H00CcGWMwMFfHXBLiwMmEia0iheErFX+apzdpD/LgM9x8eXgEOytjm8rds/GNYpy4Th/PPV
nMMD29sIHTW0DsuL/Cgwm5lVv2veYvRdxlNWKYeWypLTStP47Vr+KqbagspMwqn0BneUZFvfwGd9
ZWvRt84sYJ9BpYMTg9PrRvDNLP5GaMU9kIZwIj0Ohtw0vJJUvcT4428PhAStnegwfzsQ4B5/ueb7
FlEzx+h7fTAe7IEaHIphZqJUZR7b7Ygepk/Z5lYl/lHCzrqvnO6Wqug14QUierNgRXSWqUM/QKN6
YcitG3r4e8xit1/VZ+YPTW1OIthzikNKg4suSovzk3+HDNpkQE3rnLMs+Y97+39rrqwY0qHe/Qhf
zTQnPmKsoVKLsVjcbN4tOXI3Wy5pnfBp5G/XmHoJma56ODVRz+8NbPgNqALbqALkdxeNRvcjDT9R
TOGlShU0UVtWmha5HaUVtOJBktzTQuEsOkxg2DP1+PkqVyQ3y2hb8BuIs0UbFQ4pHnXCbW4/HyS/
7113jHl1dcuHgL3ILOT33hPLYU466jfwlN0Q9QNnosHrnIiS+OpFKRPuWRZGMzoxmQkTXHQyI/KT
RJGML3CPQXIm2VhDctH5P76/MKI7DcsE0lSsgqJ+4NN4DZmoOYiBe9dx2KCygLEkDiGNOi/OOLJg
qzk06BydoKlELM47hSZsrlB4XoQZjJb0By0ZB2pRBbOlWpW4tMDg3xt8I0mo57qbF8uqx1RYco9L
CDeVTES3G+Bakrpegg2VoQ0BNci+LuikORE/ltI104km3oe7dPu0UV4NRutiL1FPMD1NJdaMrThk
FTpofNvQEhiw/1OpkAlBkXi2KB/Cm3SQdwnFExeK8NTI+10zBE+i25RTOzvaiLnCplx9DELk/86c
iwHZNt5bPwIo3tbtu2KuLojkiRyix7T1OxMp6LcqtRmsDG6sAAJYbXzGd1QLm/XlNdEMSnU1R92a
dXhlaJg8CplU93uVV0mljYnpU+6ir6/npCxMiwm6ntOWp3ERXacvLHeBYbsgTPeKgXaSRkj5DJrY
ZyBEh7oJ2WJlxz3CvcxlsOw0CXAKwaJTFJQVoK+uawh8gkH8+lnc2f0+WjnDKMLHW2zJBFTFkYTw
KJ3n1yBZ430KwNRO3YbKTvASY1TfKUdKqCg+SmBiHyRyrTCVOPwlfJf5EhkczkkKTXIuXFL8wH6A
efZ4nfaNv8X915w9tLZkS8RSYhqPWkidb5JYbej2ueTBpRvgwKTOrLl89ed/xARX8oa9n7ii/QKV
eD8iG6glPp0PcU43A3XmaAMwq7GEMdD8MYF9CEBuXjSmk1H0qxVClrzbKE39hoJL1eS4us7Ml2dM
rF/DAGSHYQMup7t1fiI/9NDe5/qNaGFwGzwr2tR1fodbOtQ57tGbOSN0TmFHaSROUU4mpSE/reCL
O/L/4TFBNDT/dB//JV6zes763cJduSawDTPwuVGPuzcDQnvDsy+C/KFPtYqzGPBVybtHvsIiYP9L
7yIKra+DM06O7Ac2NE+LEPZyNg0tqyoEpl305CZZgqPYN4RC3Xqz5IEL/hiXfW6Ysp/w7sGbBPlE
WfMH1f8GqlUOyvRpy6zQCFm/wuTf1/qddBPQy3xJSImHiAtN2h2ImDvulfplNpogUrkR6wBpK8gW
8MYFM3Dwhn4tpTCF0mHnFOeVH0iwiQco11CF4BpYXi8+DA48fe1Abh77hESlX642CFiGP4EfSwKj
DWgUofl/GwjrPE1rUTCRWVPP73Ng6sPIFTD/wZJ+MTmNabMtGhgSBrc4lqHUUoXW5MNGYfvEJPIf
dyjxuP7HkuyRLBlkvj2qR1QyF9tYI+n57c9eS3+mIZpwf7sxnsurw7PpLCAx+NRyfEFLGXHdf4Kq
udF3UVzBvqsYZG3htgb98tui1hE5BKHSDTa4cKgAfwk61QXrgTvBwBfptqo8IZTKpajTf3No0UMa
9lgRJUNxsp2iH+9iJ83KrS59ga/ky+wKObi0fAHBybuD4lWwfXNzciRRune1ba8vTr9cZawQrL3q
0uO7TGEQg9fJ2UCXwhH11bG3frklAAyBaF1jXBxLZJZmrkN196Sd/KNO1iI7yyw4NCGfAjL3o4zz
Lg/1g3ahiVzoDQkZyFxpaDz6QlfYy6ovAbu8debYem9iJ2ZCUYKKeTzwAubY7D5mMLxyNbUNfGtM
azuc5/JbKhshbmbCEWWTOVvtyAcEFXRIQH0ZMRbodDm40pdIFDjU9SCrY9mJR+umFZljuE5GwxTh
kosYKk8B/eUkuURKA9oqgM4OruFkHdkmawLpB6LcIeOfiKE4HC5LiXwJ1nSpcl/FDZJ6R3vlFmJe
c9SdZMP35Q3xUTAZJOffPj3JN4TpKJdQN/bamtIz+GMIxOtDT0hbEuONJ9HYr/HPi0NovQfYGAnV
D2HHx2OSJM9CDQEc8BiilMJC+sOaYCnAteTBEJZFLaxBakZHE5pnrxrP61Q5Fx/uWIOlnqffjeAb
6T69WEUT61dOjP8gmYmvfM50zmeF/94hR24F4l1KPbJjZINYJe3Bsf3ejMQ5ZfhT6iamfdht2w76
Ycsle8uAD5HtTgsTGaI891VchVQq4Dgc1nFIjcwbZjAl900OIEPeT1znzkDZtsYSi4iHvubMkTym
kd6LAAbVY5uOfJpajDqrsHM/wKRqktD/Om1K2w1SA4sn8qFoG/DfTej9Q215DyHyTsLPWg2DMEbH
W1fy94cSeS87fRzHh0V92BNXITUFP7ClpcOCzHgvaWN1nm75PXgoI2vEMdk9RjH6Xlbme/yU8siN
cVUaWQwks8KMkEKNEKXOzeJqC9ng7bEoj25v5z2mq293PppaH+8mD1CMOAqsnB1kAn+JQmm6dNuB
AhT7UoPVV4OcK+hcLQlK1SqQrfIBGA5V1hhxYEWBYDUsmw2K1ly8eVvACvS4LNn2q6NdMbcTWE2c
tCF80lZzy+x4LF6WyEEoc8+91VsXhMzZ3doVqh5BubOSuOrJId14pu4txupgwrzagDveXYuIeewR
Uasjw69I4Z4wtkONfErgy+4aVidkI3pcVbn2He89NmXJErS1OEyk6vvyaWdRutUlcNqEKvFwO7dJ
VkJYuFJFrzdH8f9T2qqSXRhRViSp0sEKD3lh2PDsCUtIbFxWVCJG1/VN5/J/wVzyh5lyRi3TBU4u
UcMx3qnKtmzS+e5WPQozvdmcItsT4ycXQ67WanQbmGLvH8W+Kpiv3GfWidDPlr5faTJc1QwLjJGj
/95nV+skNcI3UCE2BXSTI+YiIJ6ztOaewkwAXdhhUvOmfLT7wLoQzkzblucpGl9rAXQ8pYpNiuBs
hP2/Gj6IgdTtKvE2l6rhC2jhRANgxDNLlcTjTRTRxFwEDh5XRTWuZjSa9UXL4Ma+gTy663o/Y8Gc
2r++acRonbUXZOLmsQDgckVfsuS90evJy0fm9R6KU3hcW2EOxN7VLm/2lsr898q7sHs/lzv9ZjjW
468WyEaSMYQUQVFguDaOX4wvILEnoQhCIoqjsV3xuLdTtziQnfu6gIArphbV0I7Nd+CZl5cJxQed
Yv/KXZJTafECd8cdvQ4qvoSiVhfJakWuZhnECNqIc0rqOn41TBBBL7rnXMLva9IZmEjZLWO3KDF9
ObEy4mhHd8J7cDTVf9la6h5/3jlpktt2EwwoGHhPIYbsTc3N+mlMPh8bOlEi6ZfqDno7EtA8oEsz
qegSKANrxBgfdqD1Nscd5Sp/+EFzZcq0oCGr5n1+uXubnNb0RgNDd6RV1vkhldlXZxTA0jnyKiEb
oW3AEfeE9WzZlhBwIO5AZyvBJgkWofQlTIHN1WgQ19MFD90zy/04mP0=
`protect end_protected
