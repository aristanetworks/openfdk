--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
A1uJtMHy7zGuoG88vigIeyU0LdYQo7tW3mJv4Ec9F9ufoFSOYPuKoL1AnZrXEjtzvtqi9yzL3JQ4
HGko9Z74yUd1J1KmcI6excowGcsE5CP5mtDATyI17aLylZZHaIf/ZDGcrbQ2i586f4dF0D/AAkpy
/3xWR+U93/xJ2gNFpsHaznGgMxba+eZw4e0d6kgW+cLTW6Y36To9dKbUeMD3vxijyibg6xIw/TMT
3jHNh3bOw3VrpZeR8UgU+xtr2Q33NWKIujahR2iOCMMZfdBNQ2avW2NmJic8wwZ2X/NWF3cq6ovA
PG2tBkRsgHxGfSc30VLR7vujLJ6fZlHPXqRzRg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="aaJZKC7oBQMpVnDC0jvz3NbO+M6vOJmht8xbBvZG61U="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
jZOTSl6hBSvyvErkx5iDu7wKchwuSCmdBvz5424LBI+hTvs2neKEiBJnzz4dvHL3ojyTflNnHVCh
0y0Pt0WEv7CLOBOrqZ3Z0JfFkA808ujAzn0YcIboAhkDP2d5EPdWRssAL+2sFcbS/+nleDaT1KsS
CF8Y2Dm3JNwKvfTl2Tihme+mtg79nX9w6bmYrNtqT2pdOydN3YSH4iSWFBHYOwmdECiRPljMsPxX
c51TFgDFDPDYoprIsAxCQ95ew1cHOizn4SFZqb0SAp1EL5Rjdecx6wVXXLzIHKmcGr2fEm2pryGO
XcEvuwYRkTIz/DHxUEUhMRb+Ao9LR8VMHWiwYw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="9ofgWyXtWA6ubrmRCuhsDpLpJbLWi9faY7Gp+N3maYE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`protect data_block
dkOarUg+BkXvnbIQkzXmAUL1Tl321I9I6UCcqydpORuoQ81fWe1vln4KBECjMoYl5rlbOrQ+tc6d
wPgd4lFP1I7V028BtjWZFRBJafwjtn19lMvs/wcwQs1fHL9rmH2LzvFJZpw0NMBKzXFyh1zrpz0h
GyRsCnItTl+6WaRoP6xzUxZY+1S5MhsU9vI7l5k0NwT166gLk/7I6LWZYTHi0V0CvS2D8Ug2ysiB
mzNQuCUEz9l/gCuEjQvcmlDdZ3MHGOYxY1mApi9Vbe3NaxGt+3wiOleU18Yzh861Wqx8ZiS66zLm
WVunUkBmWH7s3JHoghjlhS42bGohe9ujAANYQm+dJlBuL5kI6KupmPp4bQvM3/WjoyCOgBKrwJnd
7WBxDyf4Jh018rHeAmyzOTWaZLtaBmayDDweBY6V6CPDolY2Q38ncUbvPwZZV5bBS7yYhp8ryDBd
b8jDRb04U6bYuzMiwAdvFt5JFRFbQERsOasjjNnIkEUPIADDmbgf4WHVT1dkzPkIwG0KI9Kew9ic
e/jAp0XwCD7NGupTPtUgLiStcub/MR9kahNSIkmSB9v8086IA5giLMuyf//FnaMu89rEumpbOmuC
W/L6Xdhaw9bQOUpYBufkZhGXEn5M9in6wj0VmT5miTY0tiznF+5uusMfjzAPeJpnBlR4gpQa1ZG5
3Ete8qFXmgOXlN21YDluSU6vLTXbhVEkKIrEdEB8QIVSl3GfN3H6N3pW4s2NPZnr3vs1eCeU0GGm
7QOOBFXp7Gek6KTeZJhlumSos0e+kwEMb1TFpF25BiHvjlXHJX+X8OchEIq1Fq1i8LDwlIPi+qR2
dw/LqqxYwdACoMQPmn+fprB55/SKHEUZuaY2FXXquhr4irUc2Xft6gOJA2hOcJa/SmTBZYfYu4xr
3ZWCfvXyP6e5jLpec6MShkLBjWSoukOs1b2+PIubdyxgYy/W82JWaNZcNc22VeP0JtooOGNzPfpV
0WO3jcua0nPafkXYVYaJOy6WhdVuiOWNH7RPsYEArXxpLokqW5msP/V36t+Lkp0ZKoB1FeY4OPyL
LEF9k7Nt92yphjIgBR5ldE8dY52gHWpdEXhchI+xeGHb9kdJ6/HqRcb6DZUJq0N81r5yDQF/sGVf
JjUrnDwh++QY9UXRaKgc/er54N19QKvhx5mqRw5S77DaFCFRsM/ImkHyi50TYs+2E4hmP2AQN604
SJCsjDs9TrseWFlgfpM0kmwk0N40eFh3svpCDpXrJC6BfVlRUXOVdZLxdKJ0Y59JSh1TRISDxENr
YO548YfwtVCRrvuBgenewTdEjhloc4xu9iSp+6y/3h4xYLbgZ1S9x6WfGUtHGPJukeMMvVNVOJ2N
6sRyaGrtbfvaO7aVHyYQt4yt2Gawoxb/78n1/TzBjljM6t9SFLAZ3NTI0aeyz0saDs98GU79eczb
ZDaGyL3SQ1zJ7ycTIvCBI0inErL125wcnVl98MPaVxAEzzLrcAvVnuTQdFXsu/AYcXFWaI8SLDK6
eSd3chCns+R++bM9wUYqYbMcfp4QobgoHKSWH/vT+6Hnkl6xUT2qs8fW4SeHttSKVILVZ1JA2h7u
HQDUx5OaAY4ztMMyvWY/1cIGHzf8xXO8PUWL6w/N/t4cnQZWmI3JRO0xJ/iJ16SB/wSM2zJUq0Sg
FYxT6Y24y93ugVPii8QekG94mSNMRBE2ueEZLP/5FcN13SU6DhUsvrfISb0UyeXPMemjvkLvyCmm
gguoiSeVsBe++GGBAlLdau740Vwq+OjlPk7q4zXp+VDA159yGgjBCe5fYkgzc4ifmFhyvlkQ+YwH
/9eSPj9h1NRMf+T1kergN2B/FibalOVictVwHAF1nnVbm+DVQn8jtmxYE2u5tUyG5JTin5O1P1JD
/M8PEqfAdUgcTMoLekGlbTvCRaPKUeRx1igZiMfCCgCSSVdne4DhkJFIkQIftNQolVyLiZ01IUF9
ijTjgl9qXVn5TPaSmHMpQQyUxYEoZAlpK3NIXthrAw3FeOKG86LQuIUQU5MpBJ+X4JMQPtgrvof7
IVTYCmu+TG44zpL52o+vKtTbPb+ViemZhvh7jH/HAZoABvr4eNmzNykrVH/0yd14QOa5/n0O1PHZ
K5u1IKP1FabYRBMT0hVdJ4jtyXIzzptGB0Wrpbcuqoc7slVz3CtjXE0BM92ClH70cmyXZ0kThNcY
MdVPeZoFyMApsdmaTeiP7ER6KSIoRmFlfPTRR/l9j+wZ6eQ3FLrpPsgvkoEf8o7Qr2SAA0HKo+FN
gX6Rq7Ki1ISKMZIu0X5XkQFt5o8WRcHnImnLP7pmOtINC2+7YhOT8EW074Zp0A1V3nz5Mc4h0Jpg
7G9rGnSuO88tss3GZHTw/2cHPZVzufkk2UYEffMzpghKNEKrci958nFwF7bCDC4+3mjDV+MbMliH
wZFEdoeyY3BkMnL5EaFlcmUdJHtOSF5omKD+EcOuGpmxbv6rP2r0kFaVTl5YJQ3pbheUdbJop725
SsZqtOrNoclIuwXwx+1QH1wlDJvkDwSdN9PrEO00A0D7FtnlGIvCJLqmv7OIzhpuyuhE1K9fWNC2
U1bqIf1HxXN0irL4sZG1aD5OmPE4tvcnUsjiUTzOtqHKWdt+C4cSJHLpjlPjqgMqkvadaFy7HOe4
wAFMcNoV2GP6ANdEgpC6tPj32+kPcU1FxzeCM89dEauJdgBZIFAY4Q8fdAZeD3Wt03r15FT5B3iO
yk7BRTp+4tx7vLbY7Yt6FvNx6VGY3mfPPfbXFXivH+6Vx2GHWk2QEIp+02jzDXs9jP2X1eLY44Ks
OrKfOQ0lIbRF19heqh4YLAbCsb/VsE/N/GQ9yyhN/uZWixD1ejZ09M968qtmfv7f8IqEgu+vYVmQ
ImkzWavboC1AvonRLxfciK8jiJq7g2qfGK3aw/ihiWM2MSYzSvxlesUTKNIfrIRifF0sZ7BGiGD3
VuH33B9u2s4TFyWsuRiOn6aXajM8JOon5vbzzW90dHe1/tmA72AomENd/S26dOM/cw/asnwRGzSw
hHwxaouaCnyCrbP+szji61o5KuPWZ7PZBYtDiF8jbEuveVSjykl1lWbqWrh1AcIDmWWZnKpDIGk3
01af8IlRDGe636k3zfsfQhs217+Ll1r2k8x77ISI2JxzetROOISlmQuS19xcXXUwQPiCAPlfBPqx
vc5L8hSSnKEL7YRNLw0gxJvNGvf2qJ8fvuoidVs9OK02831ZXUhdOLqWvgcUQ+2Xfsi1/zFBO4WD
nYmMVy5hbAtprm6ghvy3vLVgAIsAfNidRAxJn5tGznRAy3H231F1WPJvC7XJimsUudSoTn9aeeih
J5Y84U+jnkmVH6ot2ctBFll0PyneLsq5e5jUWYRdJDT/eTsEq32s9idy3Xixg123/THbeKwW/K7o
O8Re4Qz+NaKZs6OQUEPHoWYCuEJXX5y4LQGLcrl8bCEYfWxhwQBCKp6qSSMe77eMu20WGmGiGqCX
xGItC05jQ6z8PBeJohM9VirYxCy/mrYX2eoAzNHbzOl9ny1M0KaC6hvcer0UeZ7e9BXeKs9ur8go
sTFuh59K/SJiPbIyTDNj5JIsSg6iWFQgs07p9SWbqjE+2YwrAEG9YKgtysMKPZikpy8xPhUxEafj
j1GlfKgNW3O2vNRd4HsS4PTPCVLZj0qnXfJSfFbSy3gfG8bCD1wmQFmPXjhe35Nra7WBF3XTW/mO
si1Uflenyk+9WhW2mUhXO0xhLGQbbroQABc2b9p6nVtqDe0Tto6lPVgU1EpZVrx+Ne08KDJg+CTd
pBS9YqdRJI+/6qyriOqiwhM+3OztjUzlQDA/ByNJ6p7mPd9SuNaumpBy4hLvOrs8thFMG/mychtm
8+PhiB+/Hg3E2/qSQ71dtoeplsQqlg//T9XUswOYB5xAcRuJyvC7CTq/1tss2486smqtObQnNvX+
aZYO85QK/yLWQMWgz/IDEMjRh4Z3PATmULOEmPolztddoab92j0ubyW2+TrRjfSya0zgQ1wofbEO
rdsmMXnX2aznUQGZhiVg8fcYiU1OwYtlIaylYmA5RlMjgIutXOuhY5p6hnkPLJsILwCkpg/oPrGr
XWWrwdNp1PSrSP8JEoX6mFJbUfMhSnDKeTpH0EuhgJ5SjTdbp+eSw6t1IpSm3+hOw+ReW1rbsseN
vz1kg1Zr+ZwOy5R0dG9EIi7gJbmXCicQkUpk/GBnFQvc
`protect end_protected
