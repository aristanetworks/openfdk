--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
hE9hK3EVMLkaMAIKrULlrXvRwpqG+QL9LuDPhmZ4VOZ5Rqym1ANiaMaXlq7UvujFG4WNc3QUUeVd
24CB7jQh1zsFIeDMUHHXPvR+WiusthT0nscsvvi2KYRg+LnDAnqrV0vkH65U5pNrypYU7WGYbwRw
3fvB608NGPrDhBeNaFARibgeHcdwNzRtK186Nr7J+8g+2AK9ayxtKod2vudChPMPk7wZ0uVQc5EB
4nLV+DyxzR3GedbfsZmlBlQhdAkXb+j8lx174zI4K4UljOYDQHV854/1BBoUxmnrDszVVxg+PgVc
K89wyW2o94AN3KokUnF44QjsRtW101W+zQvqsw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="znt47RRf21Tu2LXLw9P5vXh2LdmI4qNtH2frk1srDOk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
Rgtp3tFZMhkU7m9K4voe6LrblT8ZimxGqbx8ZpXmr3Ne9Oa4TbZnjj+Svmbxk+g/4xr2+wTMOMjj
M6IKK9h+L5ZqrkutL/e8w4jfgBXMx5jWt3XWIHLH8xCkUxvpDyjPbVgeYPug5+5GqyyuYDMZWFfX
LKGPQoYKIuyGFOZxorkIj7sICSjZtVgzLYxPlQ4N97+fk1Imcc/Lt3jNklYxULvdLT3juSK2+NWt
CDIjTuZ2Pzfh913RmM4m9UtHGFZK2OAYciJYtmhbJ6tmOzTTkRjUxpBDCH6GCP7MgmAWapn0IAuk
bjsiZvviqCGQQmsRCV+J7Z33qz/IG80BsKaJ1w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Phw3w7gB/K+6NRR99Uculi2E641+cTwnlvj79TfuGSQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2512)
`protect data_block
0QupUQCs1G5CJypsrlqB6lPpId9Ilhu7EICKRbJHA3+Lg3SNHP4peE6VxmaszkDG0hRqNpOcrmQr
7YMvnqrfzPx5V/2jI6fERPAdYF38GkEpvjMzuXtwy7rLTCEpLYGm8PPZV8fF36OwZy49rhjhnqRV
1qyjFQplqlPOsnx4u+a68Jr1mnB8gaGAzvUi5GXMWviygz3heQlSCF712jDMKwGNtFcTId8dE4nj
pduJDJxKW/+F1LsfkXmqnEZC0VkIALvdHbaHfAq/zbgQehDcZVmd9zfw7xqb6VsBcQts4UoEu1KQ
oRkDgYwVzwk5B3nu2I+HfZpt1jbhJBSX5NqcniNAH2ItfQq2Kg2nbmf4fOtvGFUQ6C6GYNmmQDc5
GkyZoPK9o3LZZd188QEjz+eb1ji3oCyKJqbY4D4jMzY32gM4A6Gjxn+e1XuDXtNWSYWQZufM4kBU
m2IaEbcSRMc3xNM8lYGOZEDJxReVczdbL738q6iSQsYoOmb0EEKPmGUc4+PiBdYinryyzSM76s0Y
zqzOk9/lxi+X+MVhnOqF3re4X/lm0TVBWBSBH1L2a1rpJ5qaCA+lNJBAk0RVwvsmvSUqSmdWrqah
+4M+wCcSrI0zWmtQvo8NvOevxL+gaa8Wnv7oO8GCPjLyGEMDtNl1Y/oW8HLl/M5wq4uLsO6WzbKj
4rAvZol7V3ebcMvIH7UGZ3jQwDjLSC20U0EZqHtYA4zi5eIjm4TfCADu7OPoNvSwgOtzErgzeOTT
lCGNijGe+G2CzI9hRe4Y0bPs99RNc8LFhy1Uvdxo5qu5FdaiYi8Fjfvo8V1RGmT28zMIVeSKnJ/T
kt3MUOOyyqsLlqkxXYNZXfjZQ+eM5lR2PnkSln2uck3JmFeisb08OA/Rv2Rv85rSrgAWg5ICwqOL
hX77KToMxltJFnbTbpAC3qqu/TkSi+NTA5iEevjZ1NxQnkS9IoBOGvU9nn9068rYj/Z2yt7NYHLA
lmt2vw3JGvBieHeTB02vYKv1MJrfKL9fRZ6TiY1HNBldH2DGcciCHTHp4Sib/1qqRSi/1/DxZCEy
xxcuj7nd6KpeGq2izCNnaRPOKDqMSVfSFdS3ceAzuFgss8odBbJxXzrUMby1qUMqHS/ZVY16iOqd
3dow0WCFcpvdUv9089aAin3I9Fr3UO4DgoMrqGr22mTUoYsi8zmSYlYbjo1/O5Vw+fWz1ChYGxtn
HRmCqYgVrZG53S6bqA31xWgUM+7aXN1UAFmgwhwjzp4ZBR+0v4nRj3E9hvS8eZju4bzCgDfSKPCX
Bs1WmAN1sUrMgwP4o098NLHgG2Kg84rFxl2jAkOMesyOZGAByv8yMcP0vv6tzgXzdhLZFyGShmMl
93uLsZ0d+h4YCRONnWtfX7/GErZ5NxW7nL3wjqbm+bx3iHenOezhrg/6GocFqpnCrG63W9ILL7fv
LlTpnnX+9JqSB9rDm0vSCTOGTUIQy/liIcWnVj8nmyT/qkK67mEdRb8u3up9Z8FT7Zh1umQn/nl4
YhKtdPxcnBamjRH7H9pE8tBBcnFo0I8FcwELdLUbFhdY/3SuN7Ri4yvFHgHOqyWA5KukjpyFFsye
HhSzl1X1uziY5aQqqC7K1XwIt/QuNcTJj9ICbcmE45Oj5B0uzAh3RtPBKX1yQgFxJBb77GfHNOeX
U8/JoH/1HPiXM957PpqtRRvZ0QCLURaFKxX4yHs0MInQGHI9KfFZOB0yDtA1NEwfUd9Dmuwug5+o
WkKdhjR45/Xhx7qPuCiWDZMX9N7a3T0JVlXoulaoH0w1PnbGRLdP7vVxw1TSySH69jvAH3LkFraT
nzgstO5X2gx0Q6nEoVisW5MCtUzmtJS0KcF/irY+Fa1IFm6WA87ue1f9pPBs57W/5VPaaB+guM/L
CER6yzi99D46klfmLm2D8rwYB6HdsYkQnDXRWSrYGY8Ezz+MinzCC4mwvG3/ptK6VrDf35uVg4do
F/t3SvPTG5QR7eCwm+Bl4Pfc6MyLoUu52uPALWqPd5VoQWMDYWn9xuXPVic9QCjNjyAt1UBbJSdC
XUnK0zXyiwzJsrRhHiah3wCP7M62MjUewG7Ckn2AZi7/+4YrQxAF4r26Rf1THPGrCb2rW4DRgWzr
T4pPsuj5zQn7s+O/dL8esaymsCBz04DgFFwnEnC26DcxbRPpJ3XPwkjfspAftYm2G5aBNO1My6zG
St8yqIJiviwd18UImQaxILOZeteDa/hILaGdcjjJ441/xPF6G0ypyY2MAhNM+86AyHI6XnWsY7u3
UkSMQ4popNQe+CP9XHbbcT8t+ZaYykr+91KyFPQS62U+HjPf/pYCj0CRPvLWgB0f9fvejPDIKbOQ
rm49t9RnqyekqjttPW5iM5i7B97UCfEFDPaJcMZ0IyMXujgLxFmE8T9bsDZ8CuBBB+c31EPWTW9+
peZvz6MiIToanii0z605V48u+wxQ0xfrXo7EYI+xG6+9Bx4rqSBeG3fgWHjcSrLr6I1EsNSFt69t
qO85TWGs30WQ+tsaFXowTFixITTCbQZGHjbjigOJYrk9Mm4kGJ/P8kN6KxneuW5TrcXGS75vxsLC
OZZ/JRenZusVseTZsqJxPYLMUIjxXZYtg87Qq/LBKL6tfvhqdlXHJ3e1SiouL06hZYn2X0GVSWoM
0J8JVygolXCP5xtnV9yBh2/er27ChQd2ktBMuXLI6TDSwHcwaoqDEkiyjwuTODgoBStHzKc9HMkS
AHhoTmGAlEXXQmcS2UOkvj1akrJ3ait+L1AaJymOHBONxDGmU5xPC6Gw/eECPO50ozFx0w6cOTQR
ETihwHYhjYawZuTyMY0T92ZCQPu78vhPpUaqPyIcyaivLCfocvtj6tKgsxcHCVv6tdm+jgH817rS
ocKGrpSbg1aSuNb+U7kFD/dk1kXHdbr11w4rQzMfKVKXxYUg9yXNbHYIP2Wad0L8/upLXF1Ompme
gOjqTORUpz0UNgSed8MTZre6fvSRaEvj6HR+97dyEdeCG9CHipYWvVItWtOkYqUZ2DojeyEV7a+L
/sjRBFfEm/vR1P9kqUM7+Y2ko8rusTaIxLFxREZS5OkPQKSmW+3kkTwTb02wP6+sqnvQLoOewg37
U4tRIItGJu2MPoDHa0OslY9OAjqJb16qBZ6OPKaWhT5G3GHJ9yCw9KDw1Eb/ScVX9uch21mjUAJo
dO5Ym1EuJutU/XDb6obHYOHJot0ofABF3bjKyoQOVxe86lgvY1xbIZ053I5D1ZNnaPGgs+r1ACLN
UTEaVBeuUwYFki8y4EYUB7nmmJDFrhdzIciKhYf4yIqABJNjSdu9+T71A2yFMtbvD+wB1jClM/26
LJVj9g==
`protect end_protected
