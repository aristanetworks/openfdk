--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
ZAfw+QiZPMVMu0cMT7D48TWENSngcGtXiUepcCPY/sOTePfFNmaG3Uco8DlkmturhNi4XMmlPc0D
t2a26CMGU0By9m3SoUDrTgs6doiAMaLb6H8ymdDorIskBXUT9DvANOSyKzlPky1ilDYXtDRS0Nuk
QtdE4uAIrGVVJ+/xhPl6YtsyJcYUoiBXBf46D6qQfKrsglsjCDF2hJEEJdjfZGWjXWKg6IVa/eSP
1l4/kFxesEzx/pecePp8cGrz0H+Y0bbaAQjtaGElt23hO0pKHLaVcv0a1qvzdfGEMBrZWHl4W7jn
GaPmfBQS3apGKaiPTC4OFLQH32z/RZKaZCO4ww==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="a5ZBf/GCeCn3iNqumnST+SyKrSIp7ZUCHhlOy3xgi+8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
QDJRMkRF5x5TaDClN9rhSOlfF2m2AS+ABzwy+LCwKAn78iU5OQdSmMZk89LDZvOJTgW9KKOZLwMw
Gap8RCkA5PODGQ/HBZJN6s1ljavlr4cxt3nTEOTpb7KALt11KuU6XtFx8PAm/xxRVmExLjma3M5d
B6h001ivwWlp3Njdy8KNAY4G4roX42/CwEUkjLkDlTIaK5nE7Mng10b6QidbN6loZ4WTDFnwiRo/
WoBqfi7LIOyQZl7jPwGm1amtpJ9RvObYtchQdXYZUNhWSXZPtUFybUwIlUsWJsAvhI4JUIDSxGrY
sFUX6UptjXmccgWB1O5NvstuOXJfJB+pyyR92g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="MmaUtQDYPzdeYB8avEGqfBQIPq/3JJxS0nCaaJZDUbY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4016)
`protect data_block
wjOprJIfieA36XKerBRPWnW7cDMP9h75edi8TPWCiZK0YXCT8kJHcrkB6LnvNF22DW6U631W5PE1
tS5DMEQcyYR93ztt0jw8KyFm9IoI5F/tEThkTlqtDV4nrNXkpwrLUqyVzrrIy2s+puYe/OIZMfcm
KenO21PVQWtk0ZBUg+JfAe3IuaAvXIo2MinRANlekRRYOpWFWL34jrYN1UCrgnDuVjS3ku5Ue9JR
/ej3rhZdJzusrMkzzyZJq1rZpW/b6vioamp0MX+8O0+ZbIfxjPB29n1thAfCCWfCKWD5ngDS8bKX
MDn6wKydIVdGTeNizNAYcYUaBcvVJROSYPAbJpKO2I/+B73hJATIbh5A4CaunaUSCpCnxDGIQjhj
K6gB9BfQc1WlDvzx6EmVIZyDDwdMTq3t1KxAdbZARmUTvfERuKBN/fnO9+vj/c6w1EFZ7n0o6Hg5
4vX47+GiouXfY9zAyHzNlt/dJzEpBgrb9fQAzxd9yvLOquPxxmVj6SNQJGzCqUVaZW8VaxsUvPfO
gYI3PebnpUejo/s/QuX0xHO8BmCiDyWGThNXLFCYuljEuvEiQVrdsnIu3i5G3qd8WJiMSzAN+yrw
aNFug6nV4X490xERF8ZoFyn2LZlZGEIgpHb8zJtJHxqwKbs0wPOtw7wzeVp3+zDny1uU69ZKzFY6
Y2BI6yn6SSAQQxzHDG/rlFkUTy+EMNMJ+5+gOapNUbso0hPwWNmm2Dxry2e1L6NXQB/axYbU9pgd
QmaAtYEgsLS/5AR2pB18Uj3OresyGbOut4xD6/ZRe9EnYaBKVicjnKiqrDkPUeiHHoX3KyqLOxCn
lb2YhRRHvFLVkmMeOC8LKQCJRm7xnWHU7kB3JAFyHyZI2Zi+UcxiXc5fQ2ogsDycHfOpQ4VeDvcl
2vxai9JCAUWVj1P7K4oQQRH3X7xJbGE21YdT8YvgDabDfvjvMP14SEcjyngblcXChw7ER0J5VIuf
0bzcMyz0GRRecSvMUPKid2218+WxnT6QevHfmZ7mbsTzjc+JpmviSVXWbtMzFDBUlkiZoArQoMAG
x4cx2G4NT0YifWQQtPVp1eQxpdNFz3pg17hVbwGDu2bf8YFe0hvYlEmbOnLTR+4YtDHuMfeb3Rnn
HgIX7NUa206bKnfbtEoyNdiEYdCGTUStuDOih/6uAPVfuKHmgqv1WR7DDMndymTMi1/vo107FABH
BnUidwzPUgmagRL1PscQTR1ii6d2prgyidRu5aUMG2QdjIeIaMDRPeLMgCbFKBmIfS7Nb7xxdzsM
pbZLN/1RUDV4NgI33IHJGgkZFF8cSfDO58/Iandn5Q8emE23mQ9AfqA20iPLJ63xsnadUvQXIDcg
1kgzH1ARZtdV+0O5re7Dtcx0igPPBY51/+TCo9zwBpc9V/ZrPX4Q3BCnx7IV695JCTvoA/CNc8xy
vuNdyZTY3fs+twZitGMa7Vr/RB5mpGPm/kXzUKVoNDMauJldOtSFUkZZcgtkGYzqYT96k2CewBKR
fn4EZ+FzmhDgI2GZcbLI+XyhCv2RKMyjkUOz7Gwr/W0rmAGnYH47jMM0xR2lOau56nnATY3cQ2TF
RAQocPy7Wpq3U82FNug/p3Wz4qw4zY0pn1E4SOhOnsaZBbko5po6DP9BtVTogi13fVqRs7ROEcm6
XNym1c82iruzLctqrQ3rtuamBMW5uwCkPJdwQaY1TXTljgjSMLy5YhOJqPoPQ49dSsIE74ouJYSe
oCBBZufJmTylMiRx6t4IspaGDOGTcHPWoM6zZRZmD6lGZ56Ff+OP9HbZGdh7FLW6C6Vt1yT48uIx
jjaut3wg5aSzH4essKcCRZCXVBPtnCVCaEWT8bBYcB6IXgJW86mVgVNJd8hu/flsLeEYF+p7PnhK
1ELF7jqnGLsY5bIVhaykFHLcfeNwxjH6mp7ErBp+B8EWviAx2YMmVrnyH+PXpu1WwzOr2osW24pR
Sq/nL10aTrfJX+Jyo80QZ48gIr9H5gPi3dkeKLFRFFBPi10drPuF35UIedQh4ZhAlVeWSrv68ThB
12Xx/Ys3TT5JrLSI5RKdYTBBTxgO6metNmgOT38PxTA5dnmHycK9I2HkIsdU2JRNlOZU5eTVlLxg
exzYTNXGTbB5zsVjHsGNcK0zeQTpwLhe9MZbBtocqsXbfgbei4NhbrlKg9Jr0uIogMEcvWyEuoAb
cVoqYfqjPgDYs8ad1LZTOGq9JYN1ek/G79y3MQVXLoxdfK8l744tMPs7gu4I0nbtdUzo8r4QZsgw
+oQpM4g5GmyaWPaQIhh9dFWVo3kZzrpdkXYjczDlu7HYcJXK0+JPZ8oKHrLskn4OXz5+aA3qepnP
6NxXVRlOsnmR6YVa4OqBg84Qs8K2Zwf1jkYTamJ8iNLWLq7drKNXKRyjw6MMHM/hd2c3asGuPYME
LRLansP8naURBNBBnW8Ctf5yduhBTyX7HPyMnbu6zoHvsgOOBV6/yI3udd6ykqHHXLl/bSYsdOIk
GrSzNLF8zlC7anifTHCLd9SwbzhXyQYbnuc+M35mGL/6JGjBDzYV1bFeocrCC1Ukc8vB+W4lc/f9
yZl2FNuUXkLg6Ec/3SZAx1cNVwMyOe7S3VnaD4JXkHPxFNTG7dG1VAIsGtm28I8KDYsla2VgITrZ
MKHeZKxWX8E+Bg4aBvV2N1UMcc4pzSFBimrXgAvq2N8qZTAdxNJruPK1+raReas0AkCZKFMZOoi+
Z2VfETdeDToqRz2nni/TxiYDh3W/2hBCr3bNjv8d5XYcuq/cKaVjl5936fvIfkNgtzhlZEs61ypW
oyGpBVrKbVV13B+QdgLzaU7QwgOaBVBujzU5TnzU+pYiM4jnCcNBs2VqrHe9UKs6kLW4Rh/6qxz+
MN74mDkwzmxRlWRR86WlUJuyo8D/LwuiJjDYsnxk97DtNiyPKQokvipSmlptma9OUowqKTWR3elM
rw1DLKWGCiEyh4it7L7LMzaz9JChTvaxvkaZO7Kk8tSxI68PJM/9jMIVa444Dvh5aoOBpRximJyO
q8U2mbhr43x6j8lOaALFnCDvONfTLb3kSoE8v0GlmK/wYreCf3yrVGmcxb7UELTsLteP1US/Wwbr
TCTUILXfAYFSTM7xBPcUxQcyr8oMXep8yeMgy15Lrl2XS4sa4sUIYd8SX0Zs4Q3TYE0Se2IwQSum
n4Iuw2ZGkrs5ZuZiwZmZmXYP+wsv+rJgeEiiuLZsqxgTM53reoLNiOiJ570AzijW8SoYMmqRNhzs
Jk5+RmtKLn9+7zg/BQe5maDL/0ArKfGL4Ko7MmWPWDX6iRLOXMbxpOANYfi8pYEXHv5SvZVo0dPu
iuQkzeJxsZwQ6/YFBc/OBFVD8B7vR8TMSVtS3Ytyou3XBcriKapKp+t/D3GmegUfrSDedwx9zwE1
xy2aI6/65yglLGm8gAqxIL2t8Kkyzzq1eDoPVqwV661Qd9+AqnUqJJN8z989/0iNjALo4vzfQ/rm
eEmpkpJmW9H5cbdJQdl/UKXeuuXCDdZtbPlfnVKpWfpwdGw/VzSfagWOQZzB1BwvIqEISNGWPFhH
JROOSMVrTYQWdAf4W3gRtAfRzl5UUMcjiGQRI6azCt233dzbuaLMDXnEcFPIehRaEYgsbUtd9/gB
ME+vHPJXWI0Ykz36/XdhBCgyg7D5xunlprzHv7dJ9nWwjwSK+/gdJju8mG2Zh4enbDhsh/P2gLiL
7icVVpikDkfHbtTF0fh0P8nt9A67j501dC2i2djy8U52Hv1C5NeT5hUjZlmjl2kP0c2QDLJMOav4
xLDnDheWjJqQsw2F5+OblM0wWIHuwc6Jz/tM7R5CUhic5PPLRoiPO7N5BTdQYjEWFA/FzfU9erSU
U4jl6npVh8SqWWGOstAwO95yh3XveSQfcBJ/Bs4p7JKOn6FJAsZADNzBO0H5eSaAlQZV5U//sDBV
i1OYjcqpsxHPWOu0PTtjwvMrq/IeV9TbygGqMcLwbEH0R645Mwo0AhcpTFihkiGFT5wimp4yXpni
BafZB6TjJzResdaQP/MEBNb/TUzodcaX0iqtKIVelGgyR8bpjDtCBBq213aGl4fC2dQX37BAkzEt
7VZhgh1rH7iVC/lFD5Tfz8H1jVAyyVEiu2LzIPYhOxsW8w1+17bAHJSXLf3aeKambN3gU3442HfG
F/qrfXCXlBKc0kxdYxnNMQPYO+1v7jOMR6OgVoWWY3PqrS/H1WD/2K1hiPEj2acckm7d5IWSefxS
MceMTEgGP9B/T1pIDML+m5Lc1Lv/Xd8/smnSVHkmfBXtTQ3hoDbl8AeZ8SkMhp1bukfWEqnZ7Zr3
OFEgQaTjUVT2lWS8LJPYh5N3Sk4NxUhqGoUnuEmNz09CJ6atP0fmvmjxVyrvqz3eSvjQatLO8NQE
DWiQr2rJKGX1XESygbu3xBPV8ozJR6Ozt0pJj7885kaqhvxucDjj3GmHBc1/LhaGszo/izCDf9CE
ajJ65JtZrQOcPmmmkAjPszeY9NgYphAh/TosngK3Ol+Ik8REv5LanrlCLhCjdyGZL2SX6dDnX6u2
18KgkBhsWYkwMaAjXKBbk9mJdq5W114xvgex68mDXGzK2gx9Fcjj4uak/WkZCWbLAUe/bfZv1lK5
D1vVZ09ezCbcxl6WuC55busynUtV7u34XVnKAHy1y0d9CvlW8eBRiUH3T7Kk2S9U0lNxm2B+8XqJ
hHRoHNe6UKIldBvxrH0ko/6i72MAKhqyHcNTOOEHURuRrlewge7RvwKle5CU1QVeOd8zsYO6YKrH
EtubkGAgu89XSzBl/kasR0XxZF4I+Gxbf0r8cAsMH/eY6NMt9vnogsfcBWT70c988RNT21jmiTg9
sJ6AJJizrDImb0/el108DauF/nvk9zK3XGvf0Wn0uuEK/N4yFZfzzHV2IqOP2o3jhnHPxqhnxpwy
3X6Wyp4smV+95UJDj9Kxj6C4EJJGCHykQYfjtAczDqr5ygFKcm6wcRXsFPaTNuF9gZGJJXR+N9oB
S6sz+R9/9t8cG73D5IwCWa7pASoUwIlSV2FaCpA0Em8thViQBworzGl/oie+qaR0kQ+H4BPFlbBs
1VX1Ms4/r8F6NbCrNUk06WBxplOd3pilx4f/4c6k7xts6hRUqDoBK1UhHbrkR4nIRKF7OP3IxTVk
qVFyk5stOw8+oZKFfIgJVaYbhSZRm0qipBagP4w0j6zQ0IJOYXfvgrCe29PrdxE9//1iw+H32Nkz
qAyMSrOTddOIoUiht8HaFAUWC6ZalO4nBZHACw1k+B78uy7PqtD0WUepYUr7j7nDfjMhymm157t+
e2awSDO7IQ8MIhwcDR0n3l1mczwVUyvQEfY=
`protect end_protected
