--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
TxusjnbqcSA2AoGIjw6SSpXjUq4epdmcIcBbrFXVdL+bHbKXrN9X6nRiM23uTviO9/SognNQLD1d
c8lJvYgmpIcc2TzpHlxMyWXeFXc/eBK/5NMGX17GCsFjVrbRg9jsnZX/TXS9Q1Fk/fUniIRhNC6p
aadJZcDcCSMgaP31cc9xNZqzYqZeXBFe+z6CKDWBgGK2a+j+JVh4VakfqlVqhKugLY4kNCrSDRPb
iRagVWV5pwOpRJFHe8OoN2ZE1MEG3nhRJC+W16TjdPDye9y12PtSX6vdn0MRl6Hm9t5WLsA9EPZc
zYUzrpklVKeZnqkCDS2najWRcQOVDXQXb/LK6w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="IIvIIixSDitLKc0JDheaRzXxElTA8D5LORGKoQirST0="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
H6VNYvqr736W8OGEjnSjO4uIiLUBBRRGL4luiN20gB5GOteuqVR8ZJkuTS3R5D+3uqFtY5oy/Mg9
0FjHi1+F5jmz8xWg760hxnNA3XzDdfj/sU3xVZks07gs4KJH6ofJ8FrFgUiMm7tW6wUtQxhbeB2H
ufucmCVGApl6uFV5xYkV6jHwMzV/+k/Y5WXDPAsTzMjzCmUbioW95uzcXmo7mS+p/NMdyKcXjNa8
kTNosX6rWZ765u0w9WlqQnLD+ErF/6ZgdvobV4vnl7veQM102Mf05uWnu1Hc1DJf03BvdUUr4sec
rFmnVjv9BV8VV9XEJiX8Msluq1zcMl3/zNRMwQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="fMjGaRq8WcL3GA8Pd2DKOTXJKoluzyGoW7qFQ19fy9w="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2512)
`protect data_block
sADq8ganwEX9IvVZShWRlDMaPJX2Wm713q2OrASSUsNdkz0AjDy/y6WBKgpHUI6JbkCjf89Ii7NS
yezpZQRcwn/E/oglgI4Eg2jI9eiIWM8ssrjTp4wcf5RGegKYk891QiRBRSWLo3daed6thQihUcsL
yAV9UcQOBYLD7dTOcl4WnGbSDPaQrTEXxa5TePv1aA5GAbyADXeYAf37FR7MSws2w2ZWWkHLoTC2
u42LYjFRVBFhilbuh3AF7RauiSbJmmX/VgeWQNYgfvMlagKiF8u+dUyxj1w7Tng0UfwSFTjtkQQ6
OToiDSamkGbAFl2EFxcpHKPNhjTEAJyjd+vufj4qOLUTsW/eJif9fxs/y/9aYSR9OAXQuqUJSAZR
xo8EuOXK+V4OzFo0CICT0CZGU66JQpceqffdpwflKp3jMIOJ1m7Ra+pHuiJ5r0enPb35CwOuJynd
mgxDRJR/nn1bpeNRs7LVoL4yPTlJNHgfziOcbTpOhyScnJMzfWthj3AzPML51ZwbZXY9y2FaZLKT
TIezZzXouTM+5/ltmUUgbefXbVcM5RHghp7Kw+IkXebLh/c8BQP9he7FiHfMjlJYdJgECdq8ra0N
S5ozqGrD3a6AsBLXZWmvyh7AMI9rP6YLR1OBsty+y47b5fFdrzQymiZ39vXwHlnu3ns5Q7mKlplt
hSMW3KVQICMquvU1Lz7UO4MSPXcjraDuJa6TeWacYz0LXNL7uWw0tZKlO5dN1ojN6HN/TaDvYlBX
0s5UzG64nQHv9d+xm/QCY+/uLnBv4urESNNOQfrZnlbLTUcbolRsK0f1Pr33s5oN7QE86gXOk0F7
1yOsLVdyDY0BkiRTRw2WHv54xQ1PWx3lp2/wqxYnfF/G7lb2HS//ouiNuc3NI95PDJbtbD8oCQwO
3465SOjzHkXZh8yP3ZvExkheDTu+Q/W0HOkkQi8p8/zLpfcrqJUIDGjhaiUJYy8Dqbyr/ui61nMw
s4pPzT6IPVzNvUmjg9Zcs7W48EgwKs7kaM7l94HpWjuXMEnHBm1MJZqyc3Gq+OOE0yOAld3fdTTg
u8Y3B9nAQToN/QwBymQpsT4P8nWXbdUs9m/jkLsoNovMJUUjeH/hetBhxnjUnkRivTgOpXwL/ghm
rjaJ791k5hl0F6PAdutwJVJhRh0xyfbQIs4cCKjTAylzsTm4WVzS8QJbkFnR9IzqVLzKffurh7+D
eGyZSUiZvQLhd9rApFL/aMphWvZikViRponRn4G5/z1z8KYjb8FSOYmeAJDQi6V9Nb+U2edfmq9Q
j6Bsny6yH42lP/8SXodX5mlHyA8N5DXho9TeKrCcERNzkY7Que/JUzZUsewFXXLKz+xbnfvyFB2A
N+Lw7sh6IX/F6oI/1teGTg6KBdyF+UMQtffkaW0UmGSw87ErFJKS4PWjkwrSHyFtcUst8DYovI3G
1WrcRbiQlOR3KmUt8QN9ktsO7jhEOGh95yTJ5TmZT1mGjk1M5tMYtC2mFywWgtZBlyaPIw+d46x5
hBKXwjfTwbWfslHfqw3Y+yQ6Y/zkGTrFHcZyCLevWJ6y/YrmjdJA22h8N43oBP/p785kU1YAMkVp
BcXA37V/IaEHdlXG/uy5qLvhKQwMdgLhdCdg7u/mMw6mtdU06VHw26mu+KaiX2gboZ1faiZl4ZGc
ayYHH9WpjAhF9aaCcDpln2TTICz+sF3lR3kP89/QM4hl6E7U9t+2mAnV07jozqOk42JsuJqIHn+m
fHa78Bjo9FzgpTHKgpcUFwQvK+xhIKOFdGULLisbVowDSABVbtEJ9ZrKReHzvLV3ZfH5ri3trBWe
noA0wonz1i8gJB9mGbxmbtiwP8xDpC8IuqovCmiYb5DF3PP8MLkKm+kz9wrh8gSFTsJeJImYRUbO
vSWdJQrCUohNd8U4h7rgb/cie03gM3mFDk2PFgmEXXGofNf4wZXz6e9cZATkoub25e0fj1L96eP6
H0ZMTKQXrkMAjnKV88I1ZW8phpHz36knkV46ara1bzOoPJStzObPeAuiJLfLcRdISfV7iiee08+r
3+WZ4eT+GVsuM+9jdxjpzaPot7x7w/pDrxmKlUislHoB/e88MAf+Sizg8Gy8trmYUbec3sscXdmH
gqeVj15m9fqe2nTE5ynnbEO4zY0lVVu/GhTM2vIRCHoQQA1hg0C02/B7sCJc6+/Y6GCi6tjMr4Ar
lyM7mOUh463TohvSAuwL1Ca9TLjxpxIc/1Gtgkz6RxfmnBG1NR6UaJBsulUq9win4Vu5TH4LKuTM
Se69yoQGNH8uSfIF9vHjQs6vO5XRWMJUvavnD0IYmP4/jRTRwqY8fDvtnSg+DCXcNEp7MBckdCM9
7xEgI7zZccgjrDDXKDXng0B3spc2wdebMeSHrX6Xlq1V4J6ND49SWr/zLV6dP/Ywe2ohiJpJ1oqt
nc8NcDf21QlBq6VEetzUmi37I0b8K/0wu6+b1d/2Urd2KFJir/CRwOom4LxRdhiu1As845Gg+wIH
Xs3Iw3q0tmt7hOos+Rio9BfmUfLK2KNhZl47rfyMpXpxBIGYHBe8i4Fg01+wNNmZC4EYuD0lupEm
ugHU5U8W5u3Q78QR5S2lTi+I1G5W294j+go/MOF4BxWzW6HPicQTc5JrXQISJYvf/FF7Z+/jbM0C
+d7BFzMA3p80OLbQF7E4KU996okjeKdB/7wq/yavtw7VPAHq6jOTW62e07nj5NXcIebSGeuFoihq
USU3rjbASVbPamouIkVw1sJxQzEELcq96eQdQDceGGgVyi39xETwbCzaDH3JWfeK+E9NV8nQiux8
8N/D44pEniIB9/4FqnGlCudnJVd7CemYt1auMplk4IUK2bGYgnbTRMslJeY4642ldWSFVmsLeOZw
FCwPaH0piA0LUzYH8IPAIZmBtG2HE4EDrgbD/vq0i1UXowcwpIzAApid6c5iJElkET8NNGcZQ9Yz
EsnTmmFOx2HsD7P6DV1ta3AsrYhRJNu6RCmo7N6jzHrvU4PLx2F0YEMm78MV83QkVKP9Y0adaMHX
DOysMFfosO9jcT2ZbNJvQX//zwBeJFq9ezkYkwxvYBKmYL/vV9dtUj14GSK3Szt7T6A3K8RT1UOI
yG87Han4Sz+XTcgjLE2fKZzTLRm5AVTPPVbILTlLyJbpoLiy3LnvK8nAEtLUTplzz/TCHvywaLo3
WqaO8bngMFSv3qQpw1jlNHDRuD+V2ngVJW/C2repVGSlo6yPhBbVuOqy3l6kSyUnObt/pdR/+Ywy
WxlBt4OW1ihiA9WIRh7+lPPNFsnJ65gqQzBC8dsp1vQnX54tNxTr+SGoOQbShDhVqwLYr8MH5aJi
9Fen2Q==
`protect end_protected
