--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
VkML/WEkG108uBKxn5hbKQdEwDZs5E6Qmc3yWFbEX7x2NBdUZfcXwbRDa0n15aYU2+dsr02QBM4w
3mRUe1IQHMX6Sny2d1zXU6o3ptf5RmT0QuQPwXjWe/mvOG4X9I6keGlV8IWih0NbEc2GalTyKV2I
jsRccZQIzPu138ajL/v/Lkb8RCD2/zr8632uZb8wXSkpw71EIS4bImDTFk1IStcAESHtynrAHhU8
IE/xR+rukoXqFf938tq43ZUJ4o1moANb2ucNGMbqIJ1SYkUnYqFNpZ6Y4FFL9zNYTZN/PQ5vnCf3
P7wKVyooMMpzG1MMOMN1ccJ7SfJ/zFtC74yrqw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="LIyUOZEmYVPVTXeVqCWeui6gbsbYS6pxZzYCRjRzcTQ="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
spEYcG1uyKYdMZaMzomAf6jjH6TsdTzWlxCFruNRpMv8+9Fi/YCUAKCVu3UA85Et8Eo0Z3iaj2Il
V1CeCMmlqQ2+tMfBjXqsqJgu+h47dPlJYx1y9YHCSVieSaKJpTy2UxwuzMrteeirXHqq3O/rXH9O
duKsYouZi7MNyA+9M+v+hDLr4irAl8E9C4ct2dSUCpNi+0B7oyxBNQ7H0me0E7eWz6C6Kd9JdUNx
BMm+0r3MvrvcNDS2oAABxBxdqPS0Wye6oFzorjm0T/U7mXmNCLXP9S+wtqCRTJgKC8AiUeoTsugI
C1XIk25M2Fk3AeXzUuDl0WDV/zqprRAe8mIbZQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="GOY86EHGx0jC7ehAelJGBkfORle45PCgAYfTBe0hE+s="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
0YFx1U+T8aQAl5Yg3Pfz6/iO+I4/sgGTiHAhtXuab9Y5aHkSmhK2G5KkHEYuvyl+S/Wkl9Ej5csN
KG4GAdA6U4Ay9l8Jinjq5tMnE0bCqICWz1E2QOZ+6zAqEDrsKadFXf9ADmtDzac2fni8n4DNY+V5
1cNbOpKnRELPQjDPIjEo4Dfpe3ExvgXljZBbbu/7GqlRCEhUGWG9tFdCXxZ5EYKnuTm+4ToFdP8T
7hr4WDBRgNidYgUGEbITiv/J1MLXM/6Knk2BEDBzrlc9d9j1Lc7x6LXA81VwyeJhOFNOKL+Yst9x
aefNLX3dY8u7rRYnPbhBzpCCNZVik9FeZUOTWU/cnH6rVmU3M0QYy5SdUhEudBFM04vfFce40OQg
hUY9wh9nZB24LeLoCo6Oix08T7RPxsNynt4Ub7LO9I1wo98FPKRPYvAuyYRe2oYliYZclDc/1agt
VDH6BlgDaEIPQ6/TYcjTIFwDmbuI+nTiHeeAevLLKbYgqlA8tSSvvXktQ/RsMUcLqb/Jcve8GocJ
F9qidtrqQWhsNAu7PwgB8q5s2wOWI8uYgw5awfoTP5AXdTtocPu6ws0DN1zKrMqx0EQSdBVH9ghn
yICNFlDAJdfll0owAsXUjQcsHfovpK+BJHPlRF42QcAy6ZfG8LN1kVv2iVf0RKxcOFFi9LBRpUQu
+yl4iJAeiw8qpHbFmYPN5yJWWr1J/vmuDmwEk4uKUwQLlvfCTXWg8d+VgvPjiuE2SlSkCLlWMnkw
jhYqmvz4EqRb6lvjvoBDMF9L6XHOCllIVI7Hh8KLYMcK9cRhjrqPIMXH6/e1spSRv4aFkP1k2eRz
rRf44BTbkedbZQvfRe9xtSDWd2u3qq8CGw2umLy8KqgN8lsvbXiMZcciKn/wxdyPf7Fihx+VYspW
6hMH4E1FYxxzc8uGPFhiGrmCv9vFTOdeeNsO4Llsg9g2gC6WZnLGQOfB7Z/PMigpqnCd6ln7eDt6
u8YV64oGUtkdzt29O+BlWdAVHFiX6wkYj9BXmdTv/0eOJeozu26+MotmgvzaRt87aeL8sqRBSSsm
V/h7vxeaIFJWJW5o0mMwNyFJLhFGBpxNu7eQZeW3DnzDL5YBLLI93/L6lttdNUij0WOS4u6YkgJg
GNeBLbUOuTpRGsw5n4+NnRNcJW4fBZHPjBUbVuKc5QNGbT+W7i+yZP8Pawx5GGkxh/SoN1qU+cc3
euSqEQtzzRBGS/u/W7KRAP8tOZWrvCD1kBUcTaDoD7Ct7MZtCQBz76xY8m3OK/ZQHGWfpM3u9rmc
rmVQWXYm8Ron06zufW4cZZUi2l8lMp+YdXtu4nxAdgVekZyfvLdO25yOHgWGOLjaHS3PrmO51I27
0sTM+1UIMQEvDSxT74pN5gNVqTta28qanmb1zMdrf9HY/7sBb2eIISV/R4npqBm/9K0gHBv7fdu1
1nUypeqF7GXayTxnvyOuZnZ3OG+oSzjgzdZ7M0mZIrXCUDqQNDeX20Igpha87zFzRdkcQZ9yktj6
9SQ+4vMa1AJrmFNhhqd4phO4+7t67dmJ6cqzpcUw6HeS8gXpaoB1qPUXbdlP5MchU3rSiVFubg72
fU269luxZQuMcgsu12vbooyWpFtv0Aki5eRrLJatHRpid0b51AwAFrvVVZ43AAp/cglU/s1jv4F/
Hb2KkGyQmdYY92HWSQSMBF04Tu8f5yDXjjPPlD3mvaEaDs7RCrgsmSqWn7WoXLI9vy4zR3q6jUqt
SOpOA26Is0ljUnM4m4P+ZOmWpPbPL20ROQc056dD7ROhw4alYJh9qlU+rXRs0v8CyUCDlXAhe/BF
pc70bdi5oA3s51qodZIZUE2ffjhQQbph6hgiUyDW8RBsc35ywFKpSt42JJ9TEuT9QJPK6IjyqiRa
qBCgW2Vpu7+Cagh2sd5dH1IROKiwL47yaF6fZgLadzJ3QtlDCTt614E0MYJi5G1cPxNL9t6p280N
3HX7SRNux88sj+wHCls0yU2CQaC0cH8q7zK5wlF/vFf07HR9W70Sk73tgxGohYLN5chVhM/3MFSu
ZcG6cYWoU2ghpfszH2awpO9aT5XF3QDzws3YslgTk3IqoAyo8+DjzQBLmN4b2YpELi9TJDCREJNy
1Q7Gq3d/iL9QjNU9mK1GCWSwfCh+5JoaOtp9Agzc1bhQx9NO650MTr8vnf6X7PmBdKrvwTEWKuBA
Atv/s9CEtW3mWrZLIpU9GKMDODsOefraUZUKG9u4CrJlqj8vnk9rrJ1OCKvw/JER3czeeRtQ3oSv
0zrA7FokPNL1VHpZnm2cApoWzzujSzlofbTOEZRiXE06anM6Fx1ZI9KnfkcJTKTNWEyPk+eTdDNh
sgDBDM6BigsrLB/wIWpq6DvwaaJVn7PZs+N76GE+shiaWkAuqlPnIRkqNLkADAFqjKvPZfeTzSsZ
pBw6Emi2PS8t6uenhCmq2mzsVAYa4yvAn6wF4/D7yeLqnBIAtUfciYIsshmnAkVJL5Ee5WBJ0BKS
ZsMuqHQYe4nj6gqTiDlCeE0NNFze8AgZHoIlKfMX5OPsfepHZNWVHn+wspUAq+lr1BY87+rswgtP
I+AWudrJDYGdXBXKzPNapMp6P8nRzHKmKcorIwy1D9zt8HLE+h0njGreZ3iOA1Z1nii+NVAcbP77
V3P8BUafntYc9WmNpcpmQ+c4jlsE5x2N7NoCd2zHQgeez9Q1I+baBO/E4LSUPUNRA0PThhMv8Kv8
B60bnIHPc56epICZj8jONW5squ7uqfiJwY5yWPD6WBG8HCzbzg8Esl82zArAk5jid43S6aHaYDXk
dr0q8uwMBVCa1PuV1TdSePHKTuHI/3CG1KEX78PVFjXqfLnuCxdbq5vuxEmDmL52io7pD2/Pc1tV
2naRhdVL0iU3Io7oFX1Nhu2Bkkp7z+TwkWgdFAjjS9UlUoIvqejEboUb4jcEY6ecszPxfLa2ijo4
B3T+vSmnEyPre2VuBqUH2112+iVYq6JlTlQa5JQZKYLPCSMSg48xgpboP3NgSEScPDpenugcP+MU
aA74J3216QocyvXRo60N1N5vRn4HqyHGWDDCiinajlsXX5ZL7GPhDi/OSjMAOMi9/Xi6oI2pNws+
uvUmj4CzuNlyuWWzk095TCIoMjhdl15zL4tvS0HSFxvYl3/PocICCerlZ3t0rgPyufNPO8NOTaKL
J/RvzkIX3H1Tyha6jb/Ft929RXpiGvDo6vshN/+Jka5nha+xWPjJ5XWjuhTGkJBiOcgTOuLyADW6
rpRx9GcYrHWYToLwrlqasWAnhgdnL+cbZ7pa41kZuIKEChs2xtvo7bfwz+6UBGVkFZnxruIsV3Bf
SvINS0+XhgDlPjc8marIdWGdiV1i0EFNLIU57iKgCOqn6G18SMeteIAJZ4G5k9TNdvWObm6OZXkJ
dtkxim3NNf45C1IFBMwP8DuJMMVa0AWEWbf4nuWZ6LshI16ZBw7W/7s3Re/hVnrmbfWahBodf7y2
dIoU+Lw5MMQnZN1Mkf3Dj92oHHAtlEqIrsuzsqSeweuziM3631XuiZTdE1OWyAy3ppgtQPnp1zrH
x9LRdUH/J9RH2Wq5/G04OttZ6bR4I2mWnU3H3FuDOX32j6nQloZLdpl1F/ZGzNBAkDtOySaDVxeR
GSpNf0sMTfO1LHjCVwk9L83vO053x30FTJqSSzUvvgqKrgKKeZco9SoAsEq/kLxp8snBD7nrZOnx
I0AkqO0u0/tieq2rTc3032Bqzdw9om+m0FwyWBYqDUd+yk5TEQpQIV9w21E9xdxFukQ5DYmVBQA8
l/WSa+AqCJiHLibTV3lygcCNiitWSk7uwt1xb0hdrZC9IZuhXs2+I/2ZxIxnYY6UmxkLjKRo49bh
fH7N8onszLItEa614i3p7NN2CCp/bYahgwKhsNRTkouEN/LDdiDqaSaLV4CvrLzjb0atb5hmTQDR
lfWmhalzxJrPlNx5/cQxIYOclZhYhE6ROOScyQo3R67vnFLg0qldMppiLz5AhfR7xs3fwzf2kV8H
fX1UX3Tq/9ENsFe2LWUYHWEj2MXezYxExChb1oynD0S88Whfndcf/KlskpAYMZFnZ9dnsJ2NjWlu
00v98Skx73oAmGTWXdHykztxXncmDqBiNFZBy7Pj0FsNwXwFtPY/bVLkGmYw/FN7tRtIL3He69J0
yeGv8PI6mnT1u/rO3Y64Luk0+eIwM/TNFl/7DZyCUt0DDHSV+WqAltVcLnZvmnBsoNOXnWoi/5aZ
3cid4IXct5VGE2RpD6k5Vlf4VOPiSXt0gpQcEmHM2oMFoiQ+mGlFaIpwSHEiuyXwAZv7DGotK+Ht
h+7AEbgZQpi4k4rvw49c/I4T4YftYx83OmobUDkBN0VVj7M7f6B5cSJonHWnozEgu16uCKe/p+3i
lAPL7POr8fxtzJWcBn/urnaj0Pi1FYUNpQDmF4gspV4ABcqseocb0yoWs7v6W/Mgzv2oubmFHvAF
arhnduo2cUQ+1XDEYU8ZeLPXflRDFGGphIR1JjnmIhyDZ/YUCEv5sIGkrC1jUdZJKqNKsem0tgTE
XJtna+/uSxVYR0r/zgo4IUavGMoPvyiE4OV8lbH7xgLgNbZss+EEAAQ84Su/9TXfpHP0pTU7eCWF
zQ8RBYJX/3/3HVnrWtWmRYc8mda0irftlcHe14Qt/6yl4OPjEfeZW44aGu4ztJDnqvA5WUN6herr
ec3oN9ZGDds0Nqb1omzl2KiMcCoSVCE4lxXUUd+6rN+iUb3EA+Lhl0heJjyPQ6E8/mIXxnSW2kAU
fX3c+68coWM/JJygOXrWfgDh4Mv/5owIJdLveKx0uVF+DY6ds97ssiA0xMcAIFuVIR7Cqp7qr3wc
VrCi6ilfaeDnibMPi2LJg9gTaqfDJOxCghyzqSOJsTHIDGmG8SVLYEZDI8O8TVziJnPUrARJ8a6O
Tl3vj0XWEbKP1RHVAbfW52DQWK/UTEzY/45SrwA6avYX+S4w5zxuVIB8aXJXmxx2H8dhG0FHbFFh
E6LbYFRwFkzhASUFZ55olqazqH1yB9O9XZiq+SgSD16ZVlzbrhPfT34b9xiqlOjrRKGKcqpiEt80
k2XFpP9+7AXQso1EhTA1B0z13wPMJ/veIq2QziHX2SK+XIia/zUPFJZWP1MWbwgVR4oYwP2699Ie
arLqhUB3o0axPjJZeDNYOM/TPXqX0im7qBcsjb72W7MBGRKuPZqwAP8TMQVuvrgW+qOfFBLFT+ya
bJ3ZIN9sUO+kjZGM6I9ngm1DvGxNwg8GGEObYP9K292IdUV7rOhEMkvpmdAo1ODvKfzZlfdu0WW4
u0/Zb/pRmcrZolHr1jneSVgFoS1XHiIl8GR2WCJrI+RMVIshWaF/jXLiEVfYM6H6OiMMek302hHR
RU4RlpjZ9L/OtOCsUoePIzoh0NvZiR/GVyYL9qT/1qqPQNXIy2J1BK6LqkPkDIKEIiknKwwzRw9P
DaDnemW1LSw2cCW4rTtWVINLd2tiEavW8IA8ZxxWsZ5v0JBrEFnhbb0WNuZxRr0fKqSIGqRqigzM
isc0SBNgFeoDFunB7qAVGVXYvqjHCxyShKycbU8xbzNxzkE4EH5/MmW/3LlxsCjlT0+lbJaC1cGa
RxvtHg5+3d87/UrspqndPFTEg3EAX5SFBxWUK0pA4qarTcgU+rxrhQvkME5LlXuhk1tGzqQKG08E
+V/laS8dzgqNufK7iiz6LRiZdsRCOKln3lTYN/Tlux3qhlzfPe9EqotikPWLNmtLLiZyV3JxKS0X
FKgoxpv3erPXf+LXFaZ7xtCeIV7E/U5UTPL7UelcFeh4xeYsi8tjhO5miFqDyBjPzK8+0xtpatd/
Flbvy7nXqiPwKpKHR3kHp9oXtUAnk9BM5EKzbsePM0S6ex1owtPV3mK8O+rzMbiLNqNpsY4x52e8
ugWYZsoG2JLU//gzoYT052ZWiLEjk2Q8tcOlzg1nUImm+/IG6B0Q5jNGzSGZcbVf0AU8a+dHzswx
IkyWUvSk6S1lAm1HCUyUBl4Hq4ptJcqX78W+55C2bxy87ZXxksBjv9wQ9mNSI0XBD28mM5H3AQ1m
EJ3vytMFp0JanV8H7wb0BEuDI8pR+mNjPBVHg6hxggcfeBYiaRZsjcCGEe84p/31YbYco9gluXd/
TrjLPf48Ecwix2a3GDhZEwzsyZizKCGq5h6/STMCbb4FtkPKKY9kO1r9TBeABd00EZPQrgWi543O
UjebOvSZXKPrRqFBAbThja2CksEsA2nsoFo9SmEgz7mU48iKUFrL6dF6pZe8a02z+fo8y3OHO6Xy
cFBTp0bRAAVbpEyOtvSZ9fTtYQSUmMQ/zSI/BKQZKrHkZ8n+D+7PpvFnint7HDs0HewdbwXCB0sB
Jjs2OIqa0JzYISZtToAlwVj9vuIi1uasVdREWVnyCgwHEe1N1qu8VRjGtUatqkLSfzwgs2UUX5so
1mFl+kog0ZisGf45tUkfSojbNqHRC4HCEgCS+D7Z2vuTB4nXdsQ0SBPylOaiFW+FTe2nd2rsuS54
78OWNjIm5zQ2Itxlg811IGIfYaYIh5ff9Vzl27xuXUD6T+Z2rscYfeNCOTBtfHRwj+tlm5qz0hrf
ztnnYEYar1SqdqH/wDsUdfvZIGWPnWzBx6VX3YdETDFDQfzk//qtMeU5ANaO2+T1NrBEznDHab3/
ek/aqZV94oATVHX37NLtE6vAWSWvPXnAvwFPVQeZ/xxyxNFSDH5+y4N+S3QZ9jgOnt4II80wM/Yr
EuknQo53VNO+NyEo/RTdiKMNzeR+uWbpNm+fUwW5gJ1D+wyaKqjgnSXTRxbI9HXDMI5BexbE10EN
Jwc9nRowqy/dw/kc1JpB0NZMwyKB2d2fGn4a7orWhzH+rQ4ICPOELqof4KLOpO4EDy/hknJ3kQK/
K7rYc6VYOYkCDf0fQgWLFGn15PbtXohbRKa/+yYiX3o7Tv+8x4kNJiU6U9Bih76c+m6qmlW/C0UI
blvqjwPp8oQoBxxVT0liLrv52JXa5I3WrRk4Xp7i4qjgG7T/BKuzWcj7wJNGc6i6l7wR/HnSbJiz
cLGQECBR+Wr9/7o=
`protect end_protected
