--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
gbrEl+RhfeZvPe0wL84n0wp02tnFHbb2072MCH2FY24zwAxIY1K9+PqpsKkBnbcsSYiAfT/mv4Wl
PaaKsNNz6v7IUqlhvZ2CCtih3EHXwxoc1HzGH3a1I+N41DvOI6FhRUbVgY0hKMJkf07vekeXoePJ
93r9v5Xaq5Nyv9i1Z/VWa1yQpRzzzIqyeMjSbhUkOAHIp+VArauP9tB7Nxl0t/GC8IhjxBUsmExU
Ph14TIf0gDnm1dmmx5l7AU4+aBEPO+jZUTPv/dKpVvHfvYsLpFpw+cWQjRW5ZikY7ZA0o108ehiL
ypnz0pBUmg7boCHX5TOOxX+IE9wcNO1Z2ettYw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Qza87G4u+9dSlbdLdMWP+d78dS1d29OFd7fCYApkh7w="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
m0y1uieNpvRNbh0p5WX5AqVzGm/2oovvb6zVFLsNhUmF+npwbHsvQ1hbe9RPWeufCLHmcF/l5/Mz
cOeWOnjOyHVIjusty4FKy2LBS2ZAJ9d82QfZSYxzVn3zBvSf/tHJl1GVDL02r3FzxpAS/HJPKZW5
QzgTHtx+hDmcPkGFo0bu2RJDdgWVP9CUtP1PPC4/emgBaOVLMS1TtAsn3iKP+emdUd4otwcxeJ63
DVE1Ge0SspKN9qyY7Y3kHEcIJc9fxS2DHR1+KpfQjgQRY729xobQeT703xA2YpL29/QlKzfR+jrf
290xDDbV0oWUvUwuNS4I2UHzVXh0sfN9yM0p2g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="NChgbCeDcr/DP0qsZkq4xaTO7RDdIiNkeIoc+XnfycQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5024)
`protect data_block
VmgZbUV9Mf3HTpK2dkRfjjoKoOdP5iOWglW4LUSIvDBs0khJqGSWJM+V539I2Eu1tMyoNc96OlDI
TXuWWh28LfQevCDJk5aSUGK1/cjlBly0obVOwppCDSn7Sf8oIa+XKPwBxLTyfQIHh4XfEkuPEouc
EtRWhiwBhkdVwxJ94o6voWscA0biY9ySl3LLWZh3VsNCIdtSx7Dmqdbtk0YXmbsIpn941aK0UYOr
8zORFZxAioQ2po4oqfQ1hop+7AbQCPXCw+Ben+eVmv+E/t83B6meFZU0ylaWIc+bYXNhXfomF59P
icplnb+LLsjeNo7qynOPFQra+BZXs+kj8z+nZkSQuAzJam9vJ/8dGeVlofBjMHCvrR2D2aX35UsX
Ir2LjIIpSbfs0QPYEUAFUNRTAdkE4eqqEyi05LsO4kNSS0MsJbsARUM+slMhjRMSCN9oEKDhcDew
uQSbvTe/0vqeBvNCIRXl8cjXHvDF5SmoocR+h2U/unvHyAMlwF4HBCdHgdfZ4kZHCxTDVJRSBOWT
fjftJUVlY284BPR7zt0edbJ6FAZof6SWRgpTYFf5oglewWH2uB3OTTp3vFJX7yQVpfm5vd+0eAua
nxJmNfk8pGRcLrpsm0BA4GvSoOj+MI/gzPuWKNoHOSqTQRDLlLgzWUOeEjl5IGXWljQ2OzmqDUN6
JSYunkjSggatQZqhcnRmX+lhw0coCUehIhDEgfnhT3+pZs2OboTufJpLBMChQPQ4t7coELnLvjc9
s2yqxO8AvDofJcGZVWYTArzGjM/AlREcc4VTE6EAnwTUYKWz0NkcXBJtbOHwraUIErkP+xwGIkqf
WLe0/htKtVkZ5vU+e2FcHTVnWrh/CncSTrzWr0c7+1UcDMYy4HCql9YDxZ3jYJA21s59LdC/NivP
Zm4AzOK44xY9JFN+Q7z7AuCHbTlbFfkpXo6OMct5MOCLg42BzNCpmA6XlRRkUTIbtdWHyiLj7URz
gr/lafJ7O8kX86tn3m9tz7oNG1ZfIZ3QG8k+Fkzgr8tGJw8EetW45mOkN5GYRu/ib6OfAw6F9mcV
qaXvfHkTw7yKSfQdvNBy5lcaOKoY0IovziNUmCTp3YRFJbR5gkXdEp7P2Krs0HCF61F7x/bHrd/L
DAxoDf0/X1QziiCnv17dxBtTWLwDVb1svmpo1LLDfzeb5ECiuY6dPTcsjhTQ2+GuWp6ue3qR2f77
/gNU5V3EnTn7F8dCItrja6ZdcXS74+v4pCGGMA+SMfAWATy+046QHcsE5xhNsRS9lbXoAuq1rWeA
loOBWlXqjuyxs3oB/Y8yL3HbvkN4ppSA9+7ht8wn7t/26ZJHg+m2DkqpxqCnGEfkIYwG+PvGv+4A
RiA++3nwTd0upaDvTHYVGdaj42terDd72WOSq5XgmLZAUfnF7IY+vILGYBP9BF1QsgvjTQ2/Wl71
SqFR8Oh08cTXWI3jLQEOHbs0QJbMVBG9XeeaOAf1YktUUZWMXUmtAgThPT9j7LrLA7BAZ8zalCe9
oSpvwQfr+U+359o9g8OTuaRVAaSAWdHMUPegLeCN0mTJoWZaRAqF2N8GWDcNx7EgELkR7NZBsBbK
A/ygyFle+X2oVW8+5HCUlU0W5S1pUvQ++5JdFEQD2FcO7qDiBHT1rYQfS9BqnDUczSPZb251y4AP
oSQg9jP+BbGN93I3/V6Vyb6mX/cgZE+dGOw69SAYroEYIPwE+ycp6ifVa8ogTO5sBtPoKofdyMfE
nd4OFtrnqy2gn2a8BBP8Bw9uzfFndZHIJxqAsBVy4Fuwsc4L1P1CuviOU2tEmWW2Snh/r/1xxX0r
g3XEYWZ9i5r+Uyc72BKgD5/2kJRTaee8eFvcKEBVIUQYphDuDDhjrqUqG52neiFOlxvzJMcIpcei
0HU3tq85e8B0DptDbiUBglDWUjeQ6vfag8L2ByjAsURy7m6vNd/gfC4yfiEEKevLdsrQpaTb+MgG
sOLEqOj4Xf9tfQzYvqwo2/uHqCQF7BFsVWDuYn1Mv7YomQ8iU0E4lOBi0xiMwOmz8GTVv4N/CCo5
hJnkzOhFkYFRBj4QNL7GhITGrGEmP9WrrR4MU909mPw2D04F0rddnzWwZRnWj6uDQIKfjHNQ6KVl
u/PRmKvVtN6er/eVIFtYMg2OaIgqoFtyznYzHFmKnCiWtsUkZms6xP5i9bTtGuLB7LcTFZZXKem0
KA4ZVRt3IF4oCHsKEn1MILEeM7/UcW/F7FAcOlNFLmnmPE6W8W27Y7cKedCe8vf3MxyrQ/JSxoH3
fESW4qsh8LumVJWLnseDf5dEZ51Eds+13iO+yKPeXiD8sePqT28g+ij7KpWDJ3bqGdXBPOxd4qVo
gy+OhwVVeBHNRSOsRF1K7s8VBt/dMKuAMtdkzUdIS+uYtsRLx80cGINCojBQ2dh+2Y3l9cjfFpQ4
ABfRSryxq4XN8lLHJUEx4elVFBUvv4DIc9q24GYSd/7umeVYh3mGsBODS69pcnHHAbX+kZv825J+
k1jx/wjVjeTunLG5VdVOXp1L8SOx4B+GnONk1lHd4Zpn5AxjoskkEDb/3Rc74dWMnxiQaXr1oAoN
tWoFEIhfJY/xd1SKtn4FQ7CSX/8pWBDluFAkm8+dvZ0lamPvcMfMLr8GpJy06wVrNlig/AaRAQTG
j/ACs/JvEb+Q50uvC8G0x9OJOn6X7fIRfgRft2l8uU5OPMdBeYj+dhA4yElEBg/niYkknQBJ++4L
TNKp7SfP1c4h0ZbbpbC3BYRW+hHr8cp3kmItTzCXO/C3qVcWkB8d5L/NJITHo4/iMArqcTm2ldJI
VveCRyU+6cIXgOIFmLiyZR3k6C8KKFDNS/3ZRgF1+uFkYpWwuV1bC4S+CD9FOvSllPwXLDD32L/g
Gt6ZNg53Hp4ZX5ZMBWme/mpunCAS4kDATrp5lgSQZeuysRNXlzGNKCxxuVR7n8Igl06gN+5dEzwv
UFNNJJBZdDbRLTCh7G6dAMVRVXqxINAx67y3lQ+aMSLgJNwdIYG8ivJnGgfS1Xp0FEX9djJk1Qdo
WzXtG4L4/VuejJKn7aqynHqlSu8wC4TjqUl2nWDBmHawEot6eXZeSPeTGmltNjxgY0FjGiI3k//5
VMlM4I9a8bZucDgSJIJ19Rvlvocw2/535C0POdpooD0OoDxVHxvSi5MC1WG21bgG06xC3qi/7Yue
SiAZWWTY3gkcMDxUuq0a7jeGbb12FdUmMZzrM39Kci8Bj7bOvHsanLt00m3OhbbVjFKpFGpJdC69
V83sSzVqdtkVu5QzwCz73iJ9TXYGLyZsm70jjxBFVchhgtCqtpqqpqFZpmZU/+EJ5EHqA2n3DJK5
367qblOikPbEE7jpuPW4AecxwByE0i//KVZcm5CYHn0rwXvOlqEFcfDoPmOMe8TAouJ+D1PRPXl6
y/XaHRdyBM+HuIVxq9P99KtAkAATuCGXexJsTQem3OBqvLPQ4NSg2oQ8seXocoG9GiCmtNQjU+te
S2mHQ8gSm6fxmsur1ZcA5VqVpk+qv6ORCPi41nbROelBWGSPOZIRj35d4fhgzVpB3/qLDq0ECew9
gLYJYRTzkAM8hzqIYJkpQOd2jZRD3nsfp6+qinxVFzvK0JYA3vvB77lRi++eFxJlqyINoVCtJM9I
CPEeAVPS0xPjFSsNY2TS3VO4mAITO4/sLb2jABdun8RjH0+Jp7gBxMIiIaYabSWqdnOzSQ1CoQ9i
PEPyylyJicTtK79aKNFpLh9n4d+kfmadJK33VeLzj5aMm8U6XzxDwvFCg/nonWxrYh31Imea11vw
vncBQ51H7zffLc279ohcfLJPe10hIpjlKaD2omX6c2NA/jzqsTHk2vhBidsYoT/kD9jgNKpa9cSg
QWeMzCUWOXYSnVB525S6PI46npjSWSJDAPytDuUw4AZzFnfY6q7X8fjGUGE3ld1rXRiBSlp1BD7H
weVvmHENTsZniAKiNRAPPdToNvyj5bjlmSjFQN5QHP2UjQ7bJF5PxvrSU8PKm5I607A/VU3O53CC
bYg8AytdnS4tqgzMm6CgMttT43VfZIXXao1osYTk/NNWVGFE9dJ8ljDYJjp8jRdRS3NSVN2YAu0Q
M9YEsnaCGVrUy7KBawA2fzB5iGVDngcKJIEZe2EYw9SgUUo5PMBkbCzXYjs1/HR84JQm3OdyNhxy
s0rOCuBgq4TSHLlNAmJg38qNSfu4pnrEf+MOj2M1Bv8JuDc/JHeMi8ykl9fRqAPvIf6uRTGukxZe
KBd+p62hxwXsZ0ll0DVzwBbHvvX8Wp2+LPVz56STsck5Os+rbv031MQjgL9AVXYHAfzqzv+XNmkV
+Q9nTHAImEIAkQtRML6uWyIkKYKRnBAXiJpJSJhPk2q6HqeVOQvclnCjdkMYSNBCThs2jCAwFBPL
lcrBxBAevgg8qKMW5iYibgpAXD4YInWzpqwW6+SC9F/6SAKckwuHyMagwJ9e9oIZJZppnTFhDujT
3yFTP/7AbSCHamszm8JWyOp0qoiUrk2+jq11q2Hgywk6TYthzC1BRMEbjhayHYg1VKQVhHJaqJyI
bIz2SKtZxYzxFEj7fX34zhk3NMcx6cVpet8FrM9fSbBPIzDLTe/1EFe4MOXv9DmzBnxCuCHdxNmA
lzUSWLccHqj1xzDeOaLNcbMr4awFHDdTK54Tf5aujZQqZFpcg64K3XZbGnb2cr1+gPuzJHnt/SEh
QUdXD62EL9Ib3f3JujOYCyJa0CXRiNzkK1mXlcev0F2y5s1K4qHo22BH5SFWWBydqKe06/T7VHl8
kkoFKAuCdvfqOp7enm7Eo0s7ltDdW7PYWhjJlicJCr5gnDb/HbPaUWN6qEHyZMSHSppIaE3Qe0nG
XF1B5PKqmz2R/AZS5gpNrIh5Z/9PbTedWluXWL0O1GkgeWZW/WCJADTgBWr3Vh4R7auKb/fbLUTB
ERRV4Xb1zdAyzSHIIG/2GL0ORKMxWh+jv/mQASCqLi/rchVZ8BfCJW25g/yr4uuTlbjuxBzeg1Rb
hO2xQdcw2tsNZrnS/MzJNHg3iGYZzWyD8rKSfPPIS4pwp8nSENs6Vhjm5IrwbV/blQKMPw9vzsnn
bX0L2rJf2e8lhXu5BXXxBQRQMZnUcGTBkxWdJEjnuivmi7l21Lvvn3ajRlKfglqUeuLvPWc7C5oh
BUNnBY2k9Tjje55f2Vj3AVjA72Fsc3n9V4Wy4Zghu2CVrCLVeVZ/VwQgmOhktpU7GbaVPgau0ntQ
YaQHNno21UQ0ZgqbjG6w3H3hUSy1OVq0j+4v3uY+0tDRaWWEH8XG1A93xexQlQEq0+j8lBXSVrUS
LXpLD9Kk/1R6CHp5uaVJG6JtWyAVT7OLg3jI2R3ddODV32QDQDl0oX0U4aRaV3fBDGAlxyjFUPtT
mDJelXZG+btprKALISuTqGKxWTRAum1Dr+5pGAreAl/YwvC+hcn0V7EHA5pFCMV/UxLG2JLpqDOR
s3S9aoY5k9W5Dv/GE7mk8978krNoAfofafknLT249EJ5tqb2OiHkPcj96Ly38h6fXn9GtUhQJUJJ
5IK1qlHB/Jdh6Qo6B8qzy5ot7ECLAHFDQiS2uVIAoF47Uk6+tJxpzi+gU/qAPBsVX1e1q1UR51El
Af3X3sT5PM8oQJokk7/gvW+dWufOZ8e+vSzfobv0hsUZk39teiUIl+119f8eVPuwZ4EJTzm1qpqA
YTISF3lhvnpSbhm9HJptEVzm14+2vuJ/jD/5oJs8hneZdM625hYhVKYrwGsjtD6GuBqFxqJ9TbUs
irqWuoIPumsShhZaAF9iblZZ7Bbm+4E3O9IiZAeVjbhF7SXLP7eIzH81cFBcC8RNElROzsh8ielY
DIU5wP2fv/mDCvWbzdMpvHn0RkumsVMvEbAluMNihLsFr3ir3kq1FiWs2FCXw8ZoTcGPJXkvVQM+
KBnEI8YbaZdXlpdRQgs6KEod73xih9spQgogaPktyd2h9pktwg1EMi7T28AXSMHczxHrv+U71EbI
t2RfcwQtcAFOcw4nDI55ME8n3bLO5F7PA1krVDCtrtznPGxnRDuH4ZGT/+nJ1zDzUTff8DLlYgzS
fNIo9FNisLrAl11ZNESwt5qkcC5h7IcEHbimwX45EMZ1ySI378M6vuLkyFT4s3Wthxo26/HCsHFS
6WZz/9EqR86tisPE9haihKOyRpGW+FQVTwF7jD3ZQifQligOuoxfC2BkxsZrY3vQv9TJpmVHo9Up
Rg85vnZjXKvI6Fz5g6yNwC28uLquJrrvWgB2rvLEkxMl50kcp1DWRvL58zWRK6wxJnlqMQUhV+wE
l2gbZp4t2gzltubg8rRzyhEvM8tgvMhaEny8JQQ4LmzcMuSGbK4tenlVRNcGYOemA+/x9XFEJI7Y
IX6mR87SnumVcpmLMhrXKhC/o/fOqSkSsE7odVu+XHWbpNvJm278qQRMwLlYWKL5oC2ia/gxMraT
Xo1kvM0m9KZiQiqDh9IsLE33jcAo9YNEb4KTfF4sS941DDRghYi++guSm4zYhY2ejwfWmk0pBffC
pYLMkOH/vrFsvZf8HnczgGnb77llCHcz1lz9Qbhr//47q2leAwTHwe6rpgsAfxaOIveXLi9OljQj
BwOetoiv3vSGU8OkyPgJ34NIoN+ZDGpz5IMLx3BSb96WfG2iYqfjLh2HwrEiCwQU0VeHCU2ALp5K
w2XPvG11pi8=
`protect end_protected
