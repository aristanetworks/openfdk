--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Hof9pSXlwHdnNlBgVqTgmblxQEkjdU7N7dTPonplQ3YtCYNaBB50ZVu/jZ7rpoJiJ7ZsP3UaOTQb
NqRluOGP6E09EFXo3H3kZKElXCEwzh+I+ZRVZ1nLyzp5PYZzd4CLj6FsIQ+Cdx0Wq6EhaIpmpuYI
26xx+QOlhyZ3d9N3fMjJLcCXqGKyDzpM9WID++2KGyBOisCC6U/gRc4Lqs+dJmaump0GvPE0ZFfZ
utRE9+vp2Ti/9OXz/3A9FswcfR7qa+NueWBzvh4MMJziLfrlnH9E2rXwvYoMa7DKbzX+6SP+wzWh
gFcG+pJsJ9baPUxLRvU6/xGC0r5MZZL1YGSMzQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="poZcrqRfrmStQtGrUpyIWaq59cxvBxJmSi3lFgV5rL8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
ZIhRyWsmE5Yi3J8RbeqZmQctAInIlcyW+1Ld5naYwCiZyh9OcPq4KlHZz/Ya7J7nk+Ut+BKWRxmn
xhHLlCzY7tq/txL0YgsjuvJPO9UiQIz3o0cvC6fEHVyPf4VxEYoAsNhQOC+9TfQORWrs5VD5bXg9
r9AN+5FhMDiS9RdGVTy3nDdzUpjpBhjVAPAIPW63h3G55iH0JxHZZySTfuKSgSFuplKc+EC/GdYY
nDjNH69YZ0vjxI9/KxLTri+6AE8YnU0j6x9+bqol8Pi3SqSTh+6tIZLfSrJ1a4MfpB/RC71ZwKsP
g+6ijClX7sCuVdAemjMjoFTbzmb6i3wo0kjQ7Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="HKEQxgD/5fVC1+jX0T3gfG4fAZ6M+c5jbiujJzEhuqM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10912)
`protect data_block
qFnqYq7SLCYZwX2Ks3ELul3b/S+FHcUU865UeH5v/FxRvzP4jZbEZfqjHY6Sq/mk8/wKEProDCbo
Y17jwCNqLJUD4ThzUPRJdXbtJHmhwPdaIe/rS7L8qjzTLsGNJXljBBHNaaq3ChArZvubW6mnDgBH
dS+vhnwfkusEfK0/opWn47Np44jedyOFvueORFdjymdvmw8gF3Z8UIHppAZPG3kidoXzuuXt3TVN
T+swZDmW3/vM1NpQDnT++s2YpI53YrGL3O+TXI6HcVszIeDpoUEi0WjlywAdY8ukn7NjTGnxX+d5
jEJlqasFHAhLo8ZcCHQSesxXWsMEpgwG6NOu/zrNPXjzkfaNrW/aKLvzqpTpvf+4NftMWURPNZ+n
88jHUJ4prxJ8ibEuW816a4MCC/oUJHkv/WnclZrQbx/c7if7nSD/Zjym4UdFRv+lKZklZB2uzN3i
xllYA8EAjCPCXn99AX/pAfR3DInWQkhj/elJIOdxXX56K5g/J2mMtgJURyhVUj87Y+/D2bxNeEq0
QQHJwwM4zlGE4mXpxE0GhR0q8NkLw41yfplAJJyiYe7Jj7/Gr4XEgbCUFzNtyHHpGXB8jvr/C/xB
bZf2KxTk/Hmw9U8Mzjs9O+QDNne3/QOkBY9situNAcTn+xlRODvorv9leFKEd25M06/y/aswB2iv
NuITxoH6JGKEm2TQ9u2m9FInr2zYmwURW4r8oGksBRkqaYZZiqMXjRAUPb+EX6DHBGaWrszAJIt/
uGObLuDDR1hWyq2eSh35Imfv2llHvXUSZyLOnU/ZP10nu23zK82Ygv0AgLicNy8d/9Av2KHPCgw/
0qAEIZTDzggnjwZmYF9WGNnW1x2vocxNf60vW9BD/RshOvW4nXtjjfSxURJlnemC/kRHoJR+GkWQ
xOe+joq9bOv3ReG49d+Fwl72SqdkfXZuPPsP/IAQXg8LCLTpKlF6bcG3Mkx1yGoJAhxHN9QdjAbU
/z9AMDT/5p66RAI5EsTKw/Onp3nxebNIpxHKUJKgE1IfWprXBlhZOyHunNwlrhJEq620sYNRDzWZ
NKq5SVuKtARYej6EDlRgdNfqMGG1KpE7Y7heh90mISXMpuxYASmwpdYR+P9N0aow+Yrf+IyW9Rsh
jX317eopX1xkAK/nBeMKKLOAh/3uDoDpZiFxw3O80byYo2JlfXsSNe7dSiecCj0SxGPQZEKUYDF4
Djb4Xvan5wn81NC02SrwgCJIVZsS4KUKV0jZ1zJDTbwGOJYVlTgUt/Zn3jUsxr2X3ToXnwWYJCuj
DtCbWJWaTnSlk/gEe4wxhSaJWQUcfyAyE5pBJJMtpgXtGdhNYuf+xEoxdW5FM6ex2v0hSpLwBdQN
MzauQr+tF3lR804eI5K9ZNH9x97NDOJhtyudXXUMmbv9HHZFEB1rv89nB2o3jht7r92eWdorcizJ
FL7lUxY004YvmZYyaCW8YYeaS73nay+qML7fSIdJJsohZpMENMTdmdoXRxIbK8K8MHAR4EVylp3R
QWFgN0Z3PJfQK0iw/H+2lAEilHNgK2XKKV47b4tShQRg9MUpbpkGdUu1Pzb1pEork6ZLVgmVdFpV
VBIVpCj2RjdPOBUNqffbalOKFKxXJVLR8lz2Zi7G+Vnps8B3sUtBmFrb7K3SGasOjETDUmsCoBz6
06oCdlMBXhFdrJ0WKbc2i8DU8897yc1fQudwyipTLkJwxR6+hMsq30XHJ/DZjXsyYoCi3KNyBLAY
cYgUl2QkSe0iHOl7Du2dgY5LlAWFQEOm4Kbn1zoLySPmuWvRl9ng85S527V5REwDYpNsGBU69Q7G
H34bHoMnduHc0PSn738M9kJggYHot+eyC1tFqHcE74Ccpg2NMcLLyPRc8SVRV/Ebw1wLQZ7Mu3Gq
KaNh/OwD2aTI4+mrJkpylGUzj7dAIfUl+Mh+2iMHhhYmzi2GLv/hTK8gQQ0Cb5obWknZHz9Mhai7
UNa1PCKoCopW+7Ro3so7jQai8OPtgSGeRYJ4INAH6yPEHSeiuOCt9qfRf4UxaeltQ4fM97VK78kk
CyOi72PqIaQQW0Wtu1IzUGk5y8Z4ZycOjSx3I0CzvRYnSWmEAHbJJrIwxCcjQ7PM47P3+Shg7i7V
Xol1JIU4vS1usllxZYMd15plGUvDDVjX+rBN7JOXTWnGq1tEsrnw0HLV9ThupweVkh1nePlP8RPu
z6QZYCpGv7COZFVhPkPZS6mycutPPpaRI6tnYeME5+8OJizFDcHuL8kE9TflGe7GAQpFX3pHn1SZ
Qssi+urJbbQU/dZQXjelHSzPK4nO+6ZiFVx/c73ox2aH1zXIs2JJXqHlz9XdhXw6ZYPw4svJQhCt
EuPG5vL4UFYgzK2uaJy0vUwzA25mnyNCnL4EowgxL/UyMGN8CtzbvJDjLUya5xVqPKbXVpKQzV7a
AskO4VSoyTjK61/iUbADr9cvtT4kRSk5ph4xbr6pnp9cSt420VXvXLb8ByWtPkSh7s8w2+p+TUCN
GNhRowMH6CNo5f7Hho8Jj9qyODevK8WLHAFHaVFq3SCyAchyYLmrUtHMGO3548UWxkNUuiFekVFR
5reT+A5hUQ5JF28xcqHno+iQekSvkuoUKt/+MtdF4cY8ikiwLZVJzHbmHALZEKyD/nhlVY7YLC5x
zWE0I+lww26kA6uM/JqpQ+9G3i/q7VJAESxtAjMFjxRwfXdAjEZP0UccPU19bakb/B1worArWHod
VUGm3DPxkmpCKkBWu1CrENVl4epLSitRfpBldnjdXuk5f72I8wrlv+iCPY5JWAtkDQg8trWUOUYo
CS5IRnMRTnQeJcE7T+fu9z/A5BK/o/kmxuWKBAxgKzl71i55MOFZPV2zFnwfbdvKHV0B5hJMvYEU
Up41M0/PIKvYK2cac1i1TAoUCKmuUNbnD9COC6lK/vKZnfKbrSYo5rBueJ3XIX52dAdfc7T8x6mt
nyJ3XjbZffbtSsCkZSIpYo5NJxk36oaiS8ULg5BushXUlsnEE5twE3Q2GN0yMimfJSq5OOjWwiIt
G4cpJLj8X8Uu2Lz0Q414QOmVf64JKgNanSCeBeUvOMLUOuamB+TKXUrVMc8gYl09fxwojp5cAAyR
K1lPaSIsQt91yFF5rmk5z8+EDZh+5MjvosdLhVjvrxi284CQLckmxkOX0n3Zl3OM/V0HCXdWT71b
jRIqLXW8CL+sftSAFXF0CGL1ajF9LltCJK4MTMt91X6MXnGMFgM4nbcU1EG8hiENyck2GMCvMPiD
uh3wtYHjoxt65Se4MRUXA2yj5W82Y988AdivIaMxD+LFmzIQaIE0EO/vfbbousrZ9H/IdJx70SoA
19pJ4gRJi4hozkr5KiMf/f2gITD9gdToQ3eqLgVikdaTjm3cfeZevWvmETl1UDr0ck1tCTiQybbQ
EASrLH92RKb1e87v1TB2THXbwPYMIiq+yYzD4AM/l/3LioqyNytib7jPNeyyHro7erWVwE6sslU+
qOaClk1aEIrfG7yEEkLI/teUu5F+p64gyj8Le1hPtinNQzcmhb70C3PIRi4joGC1/RlM+6TQR6Qi
zIdo22EuMT5KqTFSHHLZaYuKfoVLZh6oKO6Sys/dfHRCjGAi6chhz51eAEHyPd62Hd5ljUwP8Xgo
Zw1FqyRE26RHVsTCbEvX/D18XQFQ+O/kjq0UN1tcGw9G9AX+OJ2kZQ2WnYm3gBj3EfzbFgfMoxdu
QB2qR3TVenMHr53ooAbM5Qw2ewMWSUBp1himojzigRLDTo7xrZYPNCJlhUv+zPIvWBX8vuGyutpg
puXOlyqi3dkMNoIScL5OTZjB/bSvu4akqwmAe631fQK86v9fVkWpjBdPQWw2vkcpzAdZ7a4O2SOO
Z6MWqz/7wETNFcd2f+RFjnAPSBGTZy5owEsQgV96i262lilYTgIFZnoywapDaJoJ3XFd31PlQobJ
xqidoisIhGiZU6yRHetykExb4YZ+GBFoOGNG61a2N6Tpid9673HRv1uy0csYAESK2L491oYR2hWt
rg5q4pXpi8jph8obWeFTkXQ5sqGgbqBCpsF8lRxXE3cUTL/pKB7as6x83z4sPcVlMycrejxygxML
OVAHeh/r+Db77mCx6YCJ64o8W5XxO4m8SUrkA4QLtDH8kl+e5cWhZb/LDYqrbKMMYp2YrrKoNaCP
eI1uNfXf1w7VkYTcRMJHdJBNYTAqe9H75/TejdZNctHpAyIZvlbBDfYgFHNhdNx8MK5Vs/FK1ost
xaHYF+UTnQwITtev1KJdLeZRcYrfxwF+XaWz/VuF8GCRxyPpXJIrhiO6LBxyEgD94+5JbQZe+d23
zVbtBYoXN23aKUTLNs5o7lVeq15LCZiZEqu7oRihZy6pZErfEPSlcDUb2Uhi1jRMs8FGFcl14UVo
enPhLdTn0AXRWT03BC5+g/x8KN06Sii6KvYgIKtvy0/5tx2YzSX0sQgXYcg3FYBsY3o+ZTswPrtk
EKDus31Jxm/yQDT0TbN5hfnn/34tJKPkZrHxRdvJodatHtZrzGHazYZNhcs4HZfrzwtY+W/gq3ne
y1hCMjgGiOjZBMj1uXWdPJncT43dMao4jekDAzbno1KEHCIcqtlBKFvKFyGpmuCJ3qi/DnWyLfnZ
oFCbzMkmcvCVuxrWZmUuwwbX1TSJZBaACiThwnHHLQDE//vsXaP1LNOXkvLiMHqDL5smgUF67UB/
en+lqnCDdEkYLVHPLCXXIibcGAkO5bVBtH6WvEkKq958aPy/CyaIdiSj302xMnHw3nnppDVT4L+v
kPsPD0UsZyY0TY4x+uEwEBv/tLu1MkBMmiINBerFjJsdFR0wed2yGvB9B1LNspFNkf7xbVFALbzF
iQQtqgqOk9CxKL42gtLCRNnAlmRL2yUhF97rd5GN22h6CLXWu2nyBPxIOLnurdIP5tb6s8GXCZrV
ljzc5lEFxio2UsIUOCt8ocpID1tsinxCC9wZjTlK0CRNZVzoQmpwVB8vZQuPUVWDSaJmnElVKBZs
8l0LzOtR7v8RJtSB9OuQasyH06Bo99OQPc/+vNINVGZb3HgKoPYvNBH5iPpBan+zkguLf/m6Qmpk
PxMNHgfWrPJNXxTstG2eiYTnXlPYyGlnf0yBn3AhttL522KbKz7in00WR3P0sTuzkpP5l9IFKX/4
eFDbPINlxA8/dFuHtFWcFH24H689PgFU0Xrh3GGEzLx3R3yUyy/EyC476CGHehxkDuxptTVlbzEm
RWSRMVLZcYdGZvCTuCTbMFXmPccUmPn648938V4UBoT8GkYCiHTDAKVyU4Kg8YoV7KkSXOqdU4So
4e/slg4xnueoU/FWxQjrvUKa9DXjkRpTnP58hbxLpCUaumq6ODFMXi2irxLBLOCdfMqUx1jSA6qZ
ZrR6I5AlDRxjpA8Aiw/21valeallR9Mci3quIeSEKAk8+DBpvfzHW73cq15wP1Y26Tms4qN7Brho
onvBCwOmvLfoPzVxeRCNrTNb5b/tlslPDMDeBQWwn74IEf1plm6GjgzJrUEdmiwG6sqk12AU7kDc
iobaxPBIfbrddo9kqO0t356KlzkdMbq/cYpLOg9Rh7ueawIxkzYt6ToZjqihwtXz01QOc0uCWPJT
+2NcxMkF9I25h3d2W+H9qd3rJ3MZt7kWVAHfzuv/1oukm77v/KaX749B0bofV5a4NTUSa4yBzLIO
nQ1T9kfSNS4X8mslwv8DSmalEJNq1Ct9lVwzYqYnoMcYACQKAr5HmQN7wrR+NI+nOPlrYdRHMV2K
gASUEDnsGf8ad42oeqZH74ofK2PtHM2UJbOxeWKchzNMw19ZXzfbg8YNuvtA0Lj841JRumCBEVIu
oFFN2OkGPkMyvXwyf0cm9EjZiidpWMSzy+jedzNve9U28A1L43SxCPJAkoY3ZiEfB7NLc8oVnoYr
2wJ+YK7l8ZqewN6YEl/KK7COLIP9kTPva76kaPPUSqBPvFgLFi29FlrpfoBJ7hiXg4u0EihhWBgM
p18EAIcZERXWQLSdsuE5fhasPCtbQhxSPVUVullXsi2CMa4Np4L8yojJS5zNrjJNinK7qxUC8LV8
oeotxsidPa5nNvSH6O6oHHH3uBPat5jSdT/FgFnNkABeX1N9j0fdasp55GoRh2oOzHS8/nM4asgW
CS8g7GJiQoPBphBMpiBcjAuPUtiBDtCYqnAT3K4pKMhp3sJ9mV3dH6QBZBQd+ywtaosVlsOgYPaX
zudXYS+3xGwiMfq3WHfh7H7+X2/57nqgtdfT66G3ybvcW2QGnmuXzXtFLUaT/XXM0pgTuSHUwjlC
Bh/Dl7dGH98VB7l5QJZMQuBHE6chauyp10vIQjVt4/y4KhIcZMQe3d6d8ZgSnaiIkJrb1qzXl404
8No4HuV2i091FkWOfFdmmxlbqEstzZg0JIcysUoRmZ97AzOzRL8gYlczhVSDpNHGgR+UHOiZQEC8
OOAJlmpiTKfdKbyPbZ275SJ0OCVFyOn/fnVYFzDXR8JKFyWgk/c2XmEdV9RnxGdK1AWcDvhGHrGY
n0xlz5uM08pmIs+mTFXwcm18h46mUYh/ylMS+5+AvQx0mpxq8kA6EvbeFWq51bdJRdc+HmEkDEbA
XGGt1pyiV98jqj0e3yPVsMy37R/Y41Jx5Myi5CgvsDMYkhO332Obmx95p8VNZuKeGWqDr0H6aIaA
RqFRZXtl0vDpixbjIJTlpEZc+YkGnazHuIfL+Fn3y8upppVBiV0yxOKZdqpbxbZGcglA2rBxBWMw
TJDmSMVDTKY8avGvQCrJl9xy73P78o2GHdbozr8l+1+qF014Y7Bi950vmMkYa/H65cVv9dhGQU8C
3DegEPvlt/YyozeiscZgCt+TbHnh2z96MWkM3Il4m6+4TXDx2UFGvgvyY6raM7W9akGAXFYEFkpn
q1zipbTvIlb0HlPJ9EAaqS3v1m3kXOo1km58akxgHrLHqJ5zRTfu245gb6rNFOBJPR1Lei+rgYtd
459ZvnohNigJiVDhF1yClIuny+uGqZssBOAWA0+qYTGmcXmsghfJgcHETnjBCRjoOl68wj4Me+tX
ympJ0CTEqtKgcBLINOY4aex6cJxN7Jo4Ig5LJXs7wYmAi3Y3lD7Xz8ReZcajOanEDU9tA5XdX56A
ynG18A3pRGhi1B0682rhVtLtQTsUjCGQ4Z5P3IFInOrJF9XZMiTMku6s3Sko5dC/T241gtHMPaNg
eFBSg1WtXC5t/NE6spqfj67ujcFOWr883RUmDD/AaLTgEaArhcvFWMRoNB2cZL7com25bvwp9ZVq
r9YO1I9b8o2/TNDMWdGrWg8vKaYsMeCL9ZTtKr15WPywTuNBr68PVAgvrzdoFjmH2LJM2Pl/Wz2I
ruxx1ciaTgZmr/lzzT+WR12tVP0qn9jttBfuhUeQotgj0tydfIpKKaHUWLHUGTzEEkoaQClpDIjC
jpgmaMg1irMJosJ8BiG+HFH5anYPw0+OrGOKXzjkKeCAzkDP/pLaMKC6QE0oyMw18ThG6TCJG4Op
BnFxnDSi4TntUR1cR8acCQChITXsPCZLZ/8Q+yXteBluncDT1fYFXdH4fosDyXsog7xvp97+O9Bi
NDHWvjqik/FpXmvERBv4xBUY5em6gF0QhvFlhoI0XGZkLe9CDi/g3Kdff6/UoL1x2KXeZKZDG0WY
LwhIT4//A/pZi00oRSFlU8UCldhRwEIlOA30kOVMsNcfPeX9DGbzbAldMMybOogwisxosI3J0bDy
KenNiejl5VEzsmvIzZclfXExu1DW71GT15qFjM4GOdMMK+jS2Yo3DHXULC6rT3R4ZU+n8PYxdNZX
b9CALZvfWm7hEHVsDt+lYl4TLPn4HHnbdB1t14iCpl+AfNqD740vnm9Bxm7w2uWFbYMjCzVvO+dX
jS9wlkfUeWKPTDG+2WzY8xnteV7hssFlgLtfqufVnSCShMIwDxZyZswJrMD3edlkHk2VMgaI5Nii
wvyIkr9zC3A7yeynV7LqjSjj490rMGKG1g3FRLYvuL71nb6ke+DwpOlrk2cpZhsydB09j7vSaT/d
36JgREMJi0sia80XvO1tH0VMXqTG5Ub1oyRyqlvP08si7XSaJX10RtIr9v377EM6Q7z3+1gc/CiB
/3Q5rIuJJtkY6k/LCY3WWh8bL1Kt4MmC6yDe+Nc3YcMUsV5poNxutjm3T3sH0HfLs/XLfK7yEPsT
oh6Qx1TJYxdvh84OqzyxSFoyQUmb72RxtUOuUfY4Ir6BGwY5JZEFq6DI0e+F+xV1krfSRQ/FlLq+
W/5YFPvyhRb6iwm79hAND1MCleq6ihgaDgEK54kksaye6opPWQyKIOs2D9qA7B8j0dPym3uANNM7
IrelcsosrNK/weE8QV3yrNu2Dyd3gSrbjBsAzIqfqnZ8pvhSVHzj0YTgdiSHTWEO7nUK5TCbGd/G
XxVk4SgO9/KuH+kmh0aNYV12Fg6A/7yZ6HPwAoH5dBBA4RiVJ58mqmz2HJlSQR/nYH9iYEN+4o3q
MIbMGRexycOb84mQ0Znc0dn+NA1nVBYRvOXcqNSpP5pjBrVpdbXacxEQsAIK7IkeeLPQZboqdVKN
rYpcg4bqb7v97m0bSHKCqMnV9KK1hQ9t1dFDbXa2AJ8dVPRFjejoZzDzpJvEdA7TXg4MwaeijcVP
2ZV23aiY6jlA6/RoSQBOpClAtWC9ubX/9IRs7oMexxvP4RmE3GUkmbuj0FeuIE4/tGudpndMwMcV
0RwJM0YDHV8TfrNgQwW4NxZ1KJviZ6838OEaQTtNIjOxZD9eoIrnt+jv7GBFd2nh3KFE0q4taLLq
mdKOh6LUWPD9IiCXHlTCGqt9DheePas1K+fHe8C7nBzImNMDzYLk79zdTwXRWYnhAmDfXfNmgHXv
HF5rIX4U+Sc/sgdGxlMZQh048jSEZYQ43DPVTNiIkMNabTr9Da9kIO3/EWw5TywbXQtyxL/xlmVj
fWBys+mJDUvRj52iT7ST5HyG7TeaH7Im8+quVPXsd3Tf+PxaojrzeVx2hQRf4FQTokvbgjv0MD5H
i4m/79hd7DWxJRqvM6jcOOlLeem7kjIvT116Iyb6ug9bX8llJIe7Sp8A8WalKAQiSI2Kt0MmYx2o
WzPRkD17UCxrtXrvVjIVvt9C7nbshDUkwoquZgldti4ovFuoZMt31deGdklQi+P09DvJA/MqTpkd
TEKxekLVd9A+t3Iy550wBObB4sNITniPoSzyntCeyNPsWwOMe1A214U5GmwhJZ4a81ycwrlxDUt0
KWXTeFUFqebwcdy2+v9iDg3jw3jL3YK18+DleEf/g1s4drINQg9NNebUEfXBu3As5cjD+CqfH8/I
ii00RLtFmBDydN+vAUlCFth80z3lu+5BD3SqqKnD/WpBm9+giNltTuLi7v4jsjSsusyaCbF4EPHt
Ah+Iv+PfDdse58IVURXPI0taX+sQ19692qay3ZsqU/4R4YkEUnXr0sOu6P8c9OaiEaG9wnP1sT/8
69YBOKsDdUZ33b/oWX31UPF7o136ISRa3A4rnpSVPmvoVkZ7td7RLGrd2FTOkyrf6f1cMUxlSbNy
0AGQivp2ZE41IVMtxcsGxU79lFfoer4O30WrnluNmGWv2Wj9Anz1Y+0ZKQWAxu+a5pBC2EWFhSnC
0sr319DksZpMZ/EjqkQulId2gMwgj4+1hnfeCT+Mk9npCpOiJ5O+37PsLZ+HZdfO/xwvrx1D6wDY
Ha1X/Z2wEfCZSdXOuA4G+aHeD1LfyA7cbslgMFbK+ZA4KWBeEr6k5kfPam/ADUUK7ihVd59eRKyi
ivahdEtY+oS0AUKXEKgSnC8jzJjJBpY6vSjArHAUKcaVSDYokGirvS2ADaJoFRNo7IHxD0mu7bxU
vGrVfcFclFLaOfmdFX4bCiRsstaD0BgM84Sfzbv5qod4KCORTSBjDEgCJBWa3+GxmfEDebmXCROH
I+po5kjjvX0/T4/Bt14wJRzYK1nFQ30LXE0XZogjdBLeoRTP9abI9+0A7KV8GA9CHqOBSw9PMemw
KXnbJRBYdUFZuVsme6I2PiZdgvXAmCmYF3YypZrHLt676uJVn152MHEzdMQmt9j+fHWjikUzs+dC
2eByKnnJTFwKKmM7l5jzH6wwrOZ7R5lqm+8Uwg7jPHbMkOM6l1vsb0fTm2Y0we9G6zu+uU2GGB1E
CMricPjFUspI3jgD5GT9EKhtRassesoLFG+oagGzc5G9aloyxnvcvAftbz7qFSxicCHUhwPNov/7
ymqMpNLlt+JLgo2C+UTNdIesJWWYUP5FGFfXXs5F3bnAH0VcwqrqtKRmC8sDHv2Wo4svIOQeaV9v
kTJkcx4z5iAsO0kY2yfs3leMopbYTdz0P9lwbNsEwj9uE8Jr7HNXdQZmr8shDNKA7hegzOGUDDav
lCBfLOVXmvptoZH/BtlOF6hphlY0z5DYCmfRi/oY5hWdEXGfrdlJ95dI41BPYnoO6A4aIwn0GUiQ
ZevJDMHesuZDjF/84udxkZWBcNnWXNPYdRZIlLJ2QD/LEDrvubQWLLOoDB/1Hj28V7//bZXQQKT1
vTMBgzMRGq2/7OzQdh++R4qsNzEzbwhn8qEliQW3W/Eq5GVke+I766yFNiNQgoCpRugyoLElmFlG
e2ZSCvtXqUFoMCIAbMJSjJIidMOzB/GB05418qRjzjc2Iab3js9RvrX3ycaoKLQsSK3f74ZeiU4B
bTWSnR/9liphlZDtGZNspqoGKZAWM0rj5UsbOciuWSQZnj1OUXij/92OxN6CWCeo1M6TkyQ5HGZK
JeKdO/FNeza1V5PCaCVvAaIgnkUVmzEcdReE7FLmX4tK5bNsF5bYByrO38uavg1PtPMQVsV/94fR
oVu8rwUI9XioPXL+DoTiLTffLpbRU+gQwvzcSLXRLyfhFyqLoMrtbOraTu1QhOIqWELYgRLbT+xc
gCdIuH+XpXKlXHpr8uanfJZJdbOsX5igYPlT0uKxlJl0XyehrsBny7haPTlheqsW17R+ZWHojxAF
rfDK38383Yr+AcuM40MuFnr+ycCGb220Xef+wdbDUL9z67D6QFh3PC30/TK0uk1nFsFx++1LsmB1
YIGNRkEPhBPnHillrFyC4U/Lp69mSm5F6cd6qyS/mLnT9TgIUULWPgPQF7SlRbOmLSlBTj38zl/Q
HUDX2dNtDTvIPfI60CsYn1hG2IMBiYOZKDF8CKYTT2uaPvCCfHlvwDBh0wTxCvfMVMCUUwjkjCvn
wq7/z27jMsIqelpg7/PefvO7dWWH2JGatkZwNVVayXb8uu6HfX7LDbtfzVYsKQ5oKGuOlKRuCKnS
HBYtOZ4EeBWJYehGexyy44MDLj1QeuC+Jk+rV2sdOsxmoMa/+GDVpOjR2HY+3/ARDjzkbbToueBA
tCMdhNLvtczB3iJGLDOmzgc54hzYOtiVOSw7drRaHxskLvjIc5sPyPd8EY/erguqs12Uykh8bGZH
2N0+qygW4uibutbG2dPI8wJuLQgZSe7fEwckZD/bG+AO6s/my2nQyr/Nf//QrA2Wlk/gtxtigYbX
isX7pLkgIeFHyA4HwxQl46wE0H2v84ggl35ubCCfka0cQh2BEIY538jwb66tl8YeoZoi/YF7EBZN
K0jfU2eF1v34VodoYjxUxUefJKZLPj4rzI4d4A5RxyeSrdt96MlEqgeOQlJ7UAxNNlLJ+Tx3+eSS
wP8Myg+bk+il2+kW3IcktyW1zvYspwc59/DIq3KlUzZbe/dWKJYu+69yigSYx2GS29Nityethjhq
pIrZvo/p58grGngyDqYG+p6QOdv0FiVh/5X6GD3NCYpF7vG3LKoy5cZkfOIYtHjrKWBGT2VH56op
cnoGrBQuXJmO3wulxAy469oNkBd7dtNRGVGmfBbAqUIxbDowle7hsmsHI/T+eTCaAk7rjO5yUbPP
2JdxsPRHXTcILNNpubiTvyAeqMs24DZGkYVwBD3YaIhHflwZqLDXYkkxoEs8+pJ0HjoL5VEtI8+e
Kla0AzuNhd1L5CTHccWGJyRAq8Fm/Yv2oqZVjtwoqYLh0aaXl87K2DO+lxf+vfJeCBV7AxWQZSvz
vpksUCr/Lc3792SEsR6XvVQfqPjr/zrmTZGq85vEDloHXIY9V14cPkW9M8+L0RtpqddIIYrIEaBw
crQPqvL5735HfzQqsyBmbH00WykzFVw9EvKIbJcn7aJb1IoUAeSY6sWrELg6gmZwYeK2YIiPMl3b
P5XmDFuTyh5SZaaoEfAZ6vo4WDjg+iuWgT4FHuuwHGnmuT6tcPVtL2SUrtFApHxXxfyhwNQxHHmN
PpCGktaL4T8y3aa+CECODjyGoQQbBVKB1kZLr2l1bOaTnaZBj/9tZwwEVHp8xMYkHW0hmn0TBAhV
ngwJKws6kGyQhlpnmdCJhNYpY62aLmQKJZBUWRsw2mFjcJNfvJc1csAYdMqygz6rzK+P7vI89Sno
nf11IVFOnfqSI8+ltr8RDWZfJqhHpjtiSgR/GP5JrhP9HCtNGKNGtJTW4x6mkHhLcvZrXjyT40Im
HcqS8j7qXehB31R+D9tsRXYqmf59qXFDa5wSH3+9hPmc9mB98QLgPDqFaEY02OeeojcpV4Vl7WTi
SXOcCKYtnzHBj+jwKcVzxZ6ft7DpczwUY4IBg9SecIaftiOZgq6besD81Pt3boE+zvFnAoTleulV
alzE1sRDeQik9G+Nf2wyqWUJ/3nMiNTafh0IKyA++doekJ3JK1dDedykWN17XSmHuJhdTGmDiS3H
UsmxuUZsnbfTk6VSwUWvU8ejA4TYK/v+eyo92ud3ZM33R9DfIusruo1pGBBz6hTivSY0Ld1RX+Fs
Tii63PYHk0aUcyvWQCbilYiipAmknORYTPDImRqVBpIyJrovs/nmOMKR+PBul+EVK/sWHzkkahTR
lfIfVkX2thgx23ftzqxA3OzJ9VPm4+2ilneyVMBGY45bb1jlZJDk2SfVdt2DfkL9n7tptEegNLnl
2ZG2HpCbzer26/zxvT5cWwOW3ZgVhHTtzuLHRiw2h1+T8fZEUAJKGgsUrOaapfGQzXivCkHcz+x4
gCaVS1KTu0r2mynWUOJygZwHGbu2qDvBtJBICjnwuxGRA2OZvVEmdZTO6UrwE9XPVqKEt2wcyvxy
nGxY8qDE3wiZC3zplC7wIVNBKeMd7vTwGgW1nCs5R0Cq3V06ycqyjvTleKX+FlVH4SngJD/VviQx
GV6RaB7Ryz1quHf+cfFCswFb0LvZseuBaIotG3WzTQrpgTJlHdhzzgZ0f+NFYoJC0Dflw5VKeE+j
IjAJtCe1k9TLUyZyxm5aAQ3xma/IQE8dYY9vscwUqaWOaK/8O1hdjmE7TuFDBrkrNE9iF7g7zh98
8LvS97psxpP9ZqqG1gnPrYjUpKllygG8tZjO7TRmoZgiFK6m3MmtVl0U9g2CEVC15zfwCJ6xKa+j
y5PZyI9RMAbaAXIx20kdTL3NwGdMic098lCWvmXM+Dxk+0RWqRylaAQdalWxobs9x+wI1HufX202
uKsTgMDcoApdRf3SHhNVx1ucETBD+EGqVbLJXbZ1l2+Xgf96ViBO0rB5KzpVzXmagaEsH0niPx1Y
YHjEF7T8KZABdzeCdqKNgnnvI6TZE6doFliXolVIpq/HuUAyMHp2cZd/Y/oagsX0CBXuE/7iWB2f
5CusJyvJOCSaaoqMfDcModEyoirrRfzEyneDTIRBKBGz5ar5CHCYqbQtcQLpQuiH/fvnc402xaSU
4ScGbOHoA4jyqPmeF/XwWRKScw3lJzzU5p6px2e6AFcTby0CUs17fgLUTSzeOr5+udkoPM+1qUcZ
tAP4J70wbjLRP2M7F8C3uI3vOpoE/XG5XGMH7HcjDE2aPELJ4CDo425WFnJ4lpgDgz6t6Cn4J0+y
F0F+7XdAKRCV4LOs1sT8n/SH1fimMJG7YBjhhjfzkDxfLYG9hIZ+4B0sAlUmObEj/UOwKofG+PUs
mSbigLs0nnW9BlSbTxyoLFtiZRRd7GVKC10YsYtUfWiMZBHh1XG4FYVayKVguHXeMMowQapKm9Fl
nwCRe+gypHAznVFEFHH6u2uRJIveSQ5pqUyQ5C63DD2tGA5H8NUI0Zu+fOj4VeTnBtKYLi5C2yWm
Z4bBT1j+4MolCR8KzrrJ9J3GN6lKmisfd2GgALTulWVgLvAAZw7uVCyqkIcAWbBhSmUuwLkbvNb1
k9dDZ97rl3ZusZ3mcGUMdjpEp7+h8GFy01eYUBRJDpmg5+iyzj3A0+ClI1eB2DJV4yGD2pQ9s0Vq
iyAhWWjEQj6of7mr1wzjGZLQAE5G2SK+NpH7Xw5gVbgOGIhl/p84GurJGkpmaIwhn6gMkkNDRAmZ
0ENHRWkwgA3z2B7RFY+/6T6d4YJWkovZb4Q3bdjr0czxLJcyTQt5fqCFTRPk+/JMY6HgFhLuneDI
SEqd/UMYBi4+O7VBst9d6AlftIZUjsbo9LfALzjdjfAQ5GF65YBtK7FAgaVlN/rRtC2uBgslPzjf
aynwlSX059PY5JWc/d+3kOjXwkBHE1wjbw==
`protect end_protected
