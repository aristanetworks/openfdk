--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Llc3FpGN52v0h00b+yMi0rIJaGJnaHbj/9W0hXDzTroKuSWrNC5rros7+upUJe67/uMJQQhKOqTN
aohHtRsEqyUt1jrZ6KtnKKtXPhJnTKTlBsXeEoU4CON47rXyG+qiJl9sE1tZ8+BOaRgHVSk4NWGw
QTzVx4b9213loqL6uS2zrmxfvva1wArHsDjlMJC3NE3YPuBoNYU7oeqMUY6T47+FG00YQOSQYejP
qnBDb+yLF5zaUG7eicLBx6QdujUddbukE637BCr2063w4I83jZDEO/R6MKD6LMl2ks3nq9KrCDex
Vwe+iICi7WS97XlevltxRfeQQBUcLpwrWsPW/w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="XekaSxz4q2CAs7dnOUKG37ssyK9Jntxg719/2cN9Qts="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
P1DjFQDewI+zq+JdvZiIovXE/SCu7+mcXv5pv43NlZrhlTsfe32CJLTZf9QLSUtEOwQ4XJs+mxg7
YV8+YLaYy5Tcs1Mfc94CHKzS4v4NBEofIMUoPdV9e7LSrDmg4b8TC3UiQi7kURckJSXFxOAFGcHd
vKJ+smV4dHD6Ja7KMOOewGB6s0tNi1Di+9WIkQRh5RMrwmM2SfbAGf6JZoTJB5H3ZztMzFMSGa63
xO46rVMdcFvuhW/b7uanHJmmoR8f8IfUoj+Kl+UcqrVeavgS2PR1Cx9yn15bAx6e4RqyQaps/T6V
68zbr7v3F37e8702LyWadS0+bsc7pN5a9lqmWg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="i3JguQ35kqa3l1Q7nvihJtwE3PO+QDaG7zC7y/3wusU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10048)
`protect data_block
cw0FHLwCJuZnb+U3wLmedeJz0keklIsFA8mxh1FS4BM0yZy+aMo6yT7Xu4PYVEU8gkj3setCouZQ
cEk899CQvjAoxmIodzBG5AoxXYvNuXvGJWOsoiTocq47O4Be5JKySRvkeCQ9hOmPpoU/5MjSyuEb
AkzblNHRmGGdhQp4OD93WLHQqJ0DWYDszG/77Mqss/5rZdmdXLbvPy5t7ZbhS5/6An1MkJ0Zad2R
W7mgYfUObucPEXKKfVcGlM3iqS29QV9pzBAqHu1nl15a5Nt7igc9Ch1OWJiaixgFnMJgJVMzLVD9
cOzEZkK21XZv2IiIjLrVPKX0i2a++4pY7JSF2tHH83z1flEwFMTdsY8U9XktdW8XVVBKyEWGO+qI
Xs4VpwvjirAulCUIu0yN+d3AhAYV/0D5IC+8tj7NgZWDKkczoihoyT41FsUob4n2jVPiLypfkgVL
CNn2QBSVvsIfbg1mgy+KUmvVFL8UgYpgxh/YtHmXaP28kfIjhztn1fHhaNHc5712UTzf/W5VW5iF
TgHqCLMh749yIlug0wQfTr5020Ysvb/PBoyTKFZpZFtQAdKIRGdAdV1xRSfBQIMkkzmAp3URkB74
itfTA1lgkmm76Jj6GzZtCjAf3zTpUSgnvu5fnDVZU60fP4Onyks5ccoVmZbakrCZH7xv6wOkLbw8
rG+wOzQkfqtrTbVkq6uJyB79zqbvaPp0CKkMbby6U7C91iGFSb1owxHnvyGR2/mc/O8Sq/x8T+PH
1iDw68WKpDTdxBlUe4FikL4t7U4GdasiyBt4pQ0hBl+KeFDt8AJUDXTqYxBo96zOWRv4llmXk/+d
saLs7qU6dxBFeJ2aTfLdoAeh2ew3VPngxMEkUbejKxNJm8cBWD7WbBk3r0kkBOXvYi/g6AjF5xMo
A2R5nW0/D3Chj5hC57Yz9r+ZzR4coGVcdhTOjpZmfmV7QPicaQMFF35mtWYDqC2NYt8R3u73RzrN
D2ZxCvSJV+x76mvKOTmJZFFkTJqRWxE9GwL4IyHT2NLSbVdNQcI5w/+I0PJhJuZVYq5v7XuBbCHW
8xsi3olF0SDfYblaNaUhM//Wygt8gwvm5HxBpEAk8pl7Bt0jB2quA2nax98SAWZAC4/AqEp2Uoyt
Y4iPoyrcWub8IEvB/tsnjMtu9Q54sp7IlD8LrAqCcobqYLZwBi8/qpRpoCsYy0eLE7QJdhLErnjl
YPS9q9c+9fL8nylKJvxN1zDbHhy+mN/dizB3ikDcTb35K48PrEdVorbzIdj08780wBDJXRFWKFrw
zJxLaBFEksO3aT0TwTZ5Mk2QN1xSNhGPO6IETXxh5wMY41wqqemWejbf/wAri/YFm++WGlZgbzoO
cMtFTE9BCStqTLWn1GoAsq8fEZOKKcNiSK3f/u7cSezKXUtceUVqPD7e1HSX0MObxaTBHTgYvKY2
fzHXRdDZbOsmB0temnJUILWRHvdhgAEeKU6NCizqIpjs7o4JCmNo9053OoqlJ/MlkbWSQUE9k8Le
x1yhV5DImBNsV2Ip/rofoyYMs0Esy6+Zpd6GshhKcoIt4c8uOid5llO64cfU16MNhz505ZBmGOaE
AdKKz5aPeHVHbBzQh1uxkQwR3SJ/rUChAGPSMB4g9mEWS7j7gwC/OSQcAe/rN5cVLBkggE2J/foi
iYHrpsv5lREimhT0DLOKUA+BuSMwg3uKGrmwVtE73NJ7RVYVoQp08gybipmEvz7g43ZDDU75cazm
+85U5lU8NN2+WCtQfU3XRw9Sqh7ZJl9AtAEttn0lo7vQOlR1sXNiQk79a6fzVJbcVx2UeIE+OkGw
SfcfrMmtwIA8mHWOeHu7NfB6K6+WFcdopPW4PSb5e1Wv7jF/zuyN6S37VSUFw/TfLhk0JPqALxjo
vrOgmHDm6+ynrQTNDwXqiXo+zC3MU6uOjRlhqenTFVTnlO+Oul0aBgngv1pJMQxtmi0oxmCG9QbU
WsT17xluErTnfncTBZfZHI3fXYMmzegWHv3b9FVp2euPGjRiCUQABGqxkJuPACaH37VH4cCOAgw8
nKSQ4Kjw4uZDu0WVXe0Dgwhzoe7o1BW3ntz8+ifYi4xbIyK9rptTObxf2JDRXRgeJAO39mbW++8Y
5TAiTPUdu46IIYlkF+yjZu1gLVNVA4+dQVi5b3Ud1+D073bGCBQ/Mwqsh9uiCN6CUEhR5hnaXR/Y
4BWXT6BvZe2ZPt+pXLslJ610U9NwiNsIiNiuVTLb6lh0OgOz3xZHXSFhc+Ao9RMjKvzOXW5PZeqH
n7XN0X17/YC3vqp6AMKqOZ0olq8VemlmtgJqOHsmExdO4AaUsofrj3z6JV/c5uPMBD8FJHBd8Ssd
c5T2mJGiaQqo8FO5AT7JewKLxic0nPvfuoEzqLB4pCCnoDU/K8sgZrhyNADLexxe9YVC+jrnfBFl
dPR7aE8MkiLGWdyW4ObV3B5KohdoiGGMBZ5aFteKrnW7hrNr6nbx2MngoIqB01I0Nl3sc5mryG42
LaxDiYngkwbb/UgQcr/3O8m7pANZJ2AokKPb4oibcB6MO/siqcINYV1HHC+raD2i7UR5JPgZejKX
vbY9gdRcETPiNSd5ZmyDREOx2WbVWY/NureukUYg/3KleVaRWTgCy9EjX2wsOtNZFwfVdi+eTNCP
EE+dapIlGoPDXltJz3s93UOtgjX9h+9dhnYMBr/pvhDs9yOHSyO6PcQqW3JSRhtE0QFsglCJJ+YA
lhFob+F5GRCX97PYDOp7FHa5JJIHbG01VVZ+ITWowtBIgke42P8YhRELZem9e0koePqcER2obijC
HwxVxErd1F3uxPEUIy3EYr0cGSMqth1Oobe/0ppILKnNJEk1hfAe35VrvpF5N3Vbf8GnC6sll75e
h60wnjosRxKf8bjoUG3x6HPZwCJSpU1envEjyJSc+8gfQkczgXHQLsuzBudKAHAbQ5Ao9HIKACx+
QstFp0KmZwmqtEvnS4HASWcltZ+OQcAs6KG1R0sPOc12y0T9cKpT5n0FV7DV1knENncToWaNaiWg
mA+h8vbapgje37i+ZCnbTm2X28EywfEA1h+1Rt2wfKm2IPrICZq9bALOz99lSAKBlneq2dBfA1a5
L1LHDznA3YO31PFFnKshMbUu8dNvHVP/kLoPetxRrQ3SzKZNQ2mIUDG/WaWmS+rHD/oF3P/CvzI5
uD0mPK2E8vOpplKpJoiOIg1B2+VwdskATkpCO+rkaHpnX1g/CCapTKj6QXTkC6oIAxBjQ6eo7oO6
x5lkuedOYPh3+dt8CwtO0qgdlifl+HWw8Q9BnL8GKOmEDKHcQSBO9ivf0oNdj1fnIHiyqrDfE31x
TTHGfhNgIdspEcAg4Ziu2gaKLCglgPkR/7Y0kd69N5I+tioCPBiTdSQpNS8PQucevCAmsTJxglyD
EeQFfy6k7q2f7bFUqH9W2TqjQC/RJInOmGY0r8QA8Ow+FzQhntRtf0ESQ4M7G+8M8KUwD2Lqwhpx
p5lBjJq8aYgnNasEOBjr32uvpf4kGK8Z61o7XwynxVBshxf9QxsmaBscckiAxkimzaA7awOLiJiK
Bb9bivezJj7Zq7/Rv7ei5TsNY7Grr/EfHVQmfFokrSaMM5YTmEyIMdl+xXAiDjwbJIg59pokseLL
UxQTLfB3SvlpkrWqAvVKq1/e/qRzKKuICKDVAIiZk5j1QqWoRtyRkAAScFEu/J/X4Y1ZpITF2gGQ
nbNBNG1QABDqASnNWIdSk9GTnkVu2lGTq6lEmV3m72YVtsqVPVCqiufyH/xlzdUF7ALA2SLAy/Fb
aUdqfUlyF8TBI/zBGJ3vQceFBOsJuS2E0O8HOLCoImKcgk+1rIGgXToj8o2DkGNon4wz46ocoL2m
qLDLzPfojeyh9l4nf1E9u7+AEvh1dEVwANKffZI6zovUsfSD+jqjtxLn1BqbJyw+iM+SAfu/vClK
NwbIRJEcXQPaodsol1SW/APRzbAl4KwAJENgy39yZ84zThv/1IpLIxI8TjKYq2kGdbYi1zqKKSe/
aLGOX7T69tLqkM0wAUfw5bayRQ4i78LLKozUvJuQDxxHp12qLu73++sLp43Wv6zy1HWKIDNxDB6t
exzAIELtFYqKDr5nRy5jp2M6C27/7hyujlFcdllCjO7GPhhnQponYUDmSux+pf4Ng9OQj1ZBqmgR
4xhXNaQ7BKCmK8kyYVHJvos9AlA43QmFi96KGhilrW7Qo7WdAuWv5okkPJqNodxCCVitFaOYVdAj
GMQ09iZW22Gdjan+SUm/aQUqZffQySMWYxhghkXN58ymLxzbey3Y8WfCrxXoFmzIOcfUn39HhsFq
gxn644l5yIp2cBIyqLje3wN5Xp7KSmkGEQb1p+RkOd5h3C9AKKhuIcsSlguntut8xhw39aTR6fRJ
jmqORDjzLnBWaIja1QXp+ijtUCMSKmSJtg2+XMEgitRnlqo8G+R0JiO83N5RDWL6vXhPUlCjtW49
OzX8tT36gKDUufdCxvdWrs5TNnPPm7AH4G2Bfqfzlw2B6Ju8bHHXB9RZrWGGx94Ky2qkkJgl6qzg
J0foc7bHvsb8zTl3Vy/QN4qDO/pdgn0XdaYH9m5+SeHwGGTSvX6/HZ84Gu/2rjVYu+VaFyGIT0S+
kgekbYl8gi/5VKih3grn1mrAGxJTpb9aiiZVmaug8RasC6UQWg5UkuvQKciLsrU4R9z9AKbOrZfp
d9sh/Xgj8+ZApb6JXeET0c5tUKB82K6/BlRJCMvXVJXB+0wCjJrNHzfxvBIAy9GBuPcyC2jrwMgE
sBhr9ljOZeihmiqIwzgveVTD5D+djyVKBOWWaWcRa6s8/mz91CWPi5ac/Nlt0t1mDbsCbN2EVidv
5waP7+20RH4SA3i+T4QaBDcfpWYRcCsd6EQOOcOxmIIc7oRTjz2LM8ztzBaWw5/D7sYXqsAS9Co5
yo2iV49zbhcDQLsWzV2juxqH9IahAJODUjylJeool/79Quy/NAe8BrqIs0iguyhE3l6Ri3YTJ5BZ
jtIHtytPtpaw7+hL8C/SubFxXPLxZx+l00C+JUzI9BZqQEuieNLlRfAJ/cbgKfFBQkK06F09fezJ
h/ly+ZqUoKGpOhXHCZRqEwOqxArTQBrwonFcysKJXHvV+y7Ggnb4SXbXkRLbjgKdah5mGYyplV4b
kvuT4ZnOwI9aV5jmykwm8TBVal06yw9I7drwUmVr4d9WmscT4K85hI/H7g4BQ5I235qE4AexXQWF
vxZV1j+YlcRWIncUaMqWiivzIhFzzPivRNd7RyZSOd0A05Q7QAwoHLlOEIFOno6Bi6CrIz1j8cX2
zl4dJyHJU/x2kZgJvZKY9mGpumKW1Luyq7kd5uiIvKgr51VofHAjCKHeI0voPr+qwKA84liD1jWZ
SqQZgK3u9tHjjKKI8iPcR32u74xC8h+0pkE7VU9YME7+3bFy9zXpUEsQvvje+oyV0IewCGKW1aHv
YVfQNN+aXTu3xcOgqrG7J9K9RNvkjT+Oku/wiEmzDZ9R1zAwycRQLEcA7L4uNtTtOIKwoYG2wNsQ
vg3p5thpjWe22B11kzhsaOQjPQvwm4FTfw+52K7TGYf0e06/WBc1ROHS7qnqmaRdFzVgOUxs+Vno
p+QwFUFMAfUsyL8fNUNSKq46u6x9At7N56JlwR9BdyxBehba6lIxnE4J3H9bHDJPzWJvIZ9rNgez
+xZL+Sz/soFNbwVpveNwVwFlO9F9ry3xJEuNM1HGMDZ/oKDhxwTv6WdDsDwC8HwmVL7hEtU8uafM
m7qFSF7OCa8jfDVVYjGmBMhXcWaO/96906aVfzi7UcJDFlK+hfIvr/XH8XsyRHUyEEr2purhaG0b
nCpHoNX/OB1z6Y9MYcHkzYPhXPUupUqpLCamAup1U2fxpyQ9qD4FVJP7npuSgD810OUxRZlUeiVf
I1plblCjkwVr1+HeLpo3D5zpp1laxZZDa4z8rmv9SS+wXo4VJ85HwTITdG+I09QYWzF/z7/PG5+e
7Z3cyY+fRnKa24MD8GrKZl8rb7VDUa3Owjj6Wq1WGZm+WI6wmQtrC9ensIR/EbMXdmq+5KrLM2Zc
exMTxLpF1TwiAPlnotA0LS5afwmGxWbZJt7uxaC1Ll9+hF2mXxZAmYAsifPzwhZ503lCeO+xL/Pi
240Rpr1Le6N0YfVBc91ovJLxJvPkhMR+jjRFniumVqxgVfKloVvEKAVZRBJtMmeoyGZ4kfE3LBQh
f0YbkdS2/6L4syhsncOZMGpHlURoG3NiG8XQ6bOSHYRqork8zbAS6mbwAd/QX8WBP6Z+TID9b8FV
QAboBb12Ug4uu7J9CKmqi6vSltuA7Cu2XZReHEvXPFvmPS8wDXM12rC8KHynjMT6TD/LGlYkHZwS
p/013RAxSM5uTdDNQWNgtRB2y4R/S+ZokZ8/x+P4sjR07C6d/tNVC8/UiOjsnGy1iaUntNpEpC4m
RQ3uh9qwIeCRGp+vPjR84KwiBmjaS3wC4fDjvFcvENflyW//05oS1195wISsVFSWqw7GK/usK/5+
UZp0ZuiY1vxeXVAFX5tACA4VLqv1hpBXUSRjaO9RMvhoW1IqS2AE+8xlx8NjQYbls51AZt617nU3
oVioSqjFncKptH00DLDWObo9D/BM/SYgPClZCr9QAjA4ARYwTEnJBptrzAwqBmfCOeYl983JI1JN
/VkCEL3o8y0Ab9doIA8D+CZBu9r//HTD3JBiQYdkd/DsS117zN49ONYWFGwXVhkZXWS2u9QznfVG
bmPft1eX5kS5SRFlPpQ3YqXXyuSLhAAGezC+V8f1ZIds766FPQb8LG9c6iYV+1h1P1VZv3+7FzrE
g8xVPp4Bw6gp0FsTJNxpoYk0rNwlvRL8EZ8gCrHU9oWy3oiOWcWiZJX0DgErNilv9OR4LXnB+p89
LiBdTVk7gkcVM+VTe/taY/XAu2M+9T9eYuU4Gw6+RUYwSEYPy2kV12FiARB6ORZReDv4xNoolFLG
3dffYrovowtFPOXhtoRoiJfVs6+oojz65kZh8lCquVl1xvIEUxfFhzfv86SfCiJjrciuuXAYkvnz
rl6lENQ5NqO2sE+HCmlYEAFbDw2KC+soeydY7QrFJIkLOiSFZBfFL1opClThLdCTZsNq+zx1L538
y4wV3ihJxLd/6eaoTzl7V+Z9lqq3fT8aWPrxFIJfCgKyTNBJioAQYXlwFZZXyPreKB3/8XcXqX7+
knrYKusWH0VWM/mRNq6VrmbTvFMH+p1LQOkok+VeFv8XTWFNL9ukF2lmxnnFrswbB2xa3J6MjkY7
7TDSMQoDfIbCSSMegUMJaTVicsYPPqnbaf8heJz9g2nLFqO515nSShOmYQfVETTVzPO/DIEFfWgm
Gg+k5lrOmWhXZWStIDol3VT31BxFdNDZOt5rZAc71FMmGrR40kU9iNyyVjfIjW/krsORi7pSjoF4
oM86Vx7IzYUNm0Xh4F6F8j9xbZyv3qLTf4F5T7pduF7Wj3VW7Ru19A5PoSCZBPl09aTi2Z50xVAc
5vTIoUEpCS5sGadNvF2RT+CVZODRhCwsJSPA3MrV2mQjvpdSfkooY7d6dmBcdKem2MzET+Pbm+65
S5ElqbCMNFNTKot6cW1OLHemmc1dhCz7kcD+WDDIVNRxV8LpnezExPPSpLJp6gYfavlHal2/kicZ
mj9XJ+YFretY8NFoSXvSf+2p1L9gSB3mkn4bK4HmX6Or+Gw/7H7iw9Nle5Dji4N8WiEdw14vueZD
kriq0u6kT6n06mH4qAszfDoXDbw+pPem9mwgvTx3MohNCnojezWqV/e6zy03XdfZQv/GE82PeSJZ
OP15R7ybjjRA1l38QJkjxv3dfWBWZJDEh58aZXQ0kN6Fm+M0eORmmb1Jtv5gTD2KQtr+4p6IlOBU
iNMSZ6pvW+zUCQfh7at1Mof7JvbhS0/+gpQCxT9YkFsLU2HfN5KG6ikTvlc6PLBkqug6NlBAgbGF
uMxpi1fIuowlRwUwy17C6ue+vgVx2nSzVQvKHmIHevpS/tUnTy66fXvpa3diJNQq/ig5wsrDGdVW
Q/puwOm1Lq2WUx+JbEVkREmDHa+WKhkSng0K1IMm6gNUnme+nbreLPhTiIYQaDMQSlIm+3+x+gq5
sWGsxqpk+sGEZfJRpllAws/6hInULQ+Cjzn9hI5wP2IPvItpYWBR8kwYUpz62mvlfY1KdlqCFfTW
XV1dkVzgHGvKUEaCLmeKwICw6XMSHUto4S3Q4IKYZoijxbjJl+jWHbVFbb9VTGx14qAZFBQGhe7E
ILgs8p7ico5gMetUq0TzhA7y6HqMVgRL+/UaBd7m4IJHvbAJR4sGCN/j9cQq2yCQegAXie9iDZ4H
ME7+mg3pMwo1Af52u5YcFsNCQzD6pJ0WfbAs4L3L/AdBtmj86CgnuBsu1pmljjnnbwNjts03/VKk
V5MyxauKouO6GR9zFCsYzJN2zy9VnWY9dlF05CVbslfEKUHbM9VUKQ75RtEQrY2dNoLtHmmEroSk
93MpUOulWakDDIZ6Omw8sjq2VF095RrpwasbQR4bjbdhMQXPMRXX0SKnE2mUQpZt2NX88gQYkYAV
vWnzt8HJbOof0W7ZEc2rnqLWJ2ndCtZpbPUZ9aqGJDF3BOhuOf1bW0IG/2Y0gigRi1tO5FlszwNo
i5WqaynVd98UHEC6+iuT17PmurXeWW8rE5hR9/08C2Od4K6YqSZdWA7xiam8hqMk7mxTn3rzx4mv
jDzRI6HDx7dDfoRcX1bl5V77ghLNmFghFDUcQ1h0CNOouuB9Txxk3ngbFBfHCphY+VRL2QE39doX
ishWvg78imZa55jwYRyirqNgitL5XPCuyzfWlX6QbUcnVReiAPhkgjlYp2VYbXSBfiaeY7rF8Zit
pJoTtHV7lQiirX8nPZ5DZRM0ieXzTe/whR6PGs6s2wVK1yWO+/ZSUuL/KgGZkAIpXVy/mRiiKON7
Dy5+D5phDTEcLwCUDpqxM7aKT4N9F4Bnz4VRvT23sXVmtpUEAXJV8CWJFlfBe4Ic0MrJK02/5Wrs
lLtew8An6z0TQQVDSYWvKlY/LcV64l21GLYyyvZOBNkIVwH0FXZeea8wVH5bSpjr+gRrXBGyIJHh
wdJYN9Sp6+KjrASi8ZhQJYSGnYVVlglDUrTYhU2E+ziYnKWipqbzbzvGcJLKTr0D4/Jt7+FB7ilh
aNPxeAzSL7taqiW62aY/RTw27ZBL8FAdySOeBjnY3fGc5r6PGcIQrJYX4m8hAaCA4sPshM4ACafy
4laAuQFaPIMFhLp6EaiuROhfayjVkuAndLH6R7A14K2TwsJk+eyAqeMY4t7mhClmR6DmImWhRQUQ
fSS6dFBzSVpI6Htttdbw3wkfQiVA0YMz5PLE0k4l58tKxFyAHulaEcWrOc3rZutC43d+0jz1ZoI8
l1RIp97gqfRotuzKJL6UMpa8BCHbX7rAxd/QlDfug7B98Em/Pt8ZgrT68wBFyp6dvFW1hazEGrxk
jCxlm7EU35JgNmxfQhH8jPXikTHX0oTz+G9JNXpYCRIBktnwLKwuxTlG293MY9xiBzU25gTlZEM2
En9fT/Xkgh8vmRuyNJcmrsEPAnXY6heWQGVU11RowYsITDVgio62uXCjvfJoqDi4yvP+DRcuS3kJ
oZ2RsyJNUHdgvpvlRRVML/gv3aMZA/SFeC4MVxjic28lheqZRSiDUjcC6BTooK3ytMKOYqP8h68F
U/wr34yCL8FuRD5Kl1mJPnI69ng/0g8Lh6q78njcGRHxkfE1VLpLzuDMn9dCsk41QthW8l7oSWRe
8sAkwHNdKrh8X4xNclVv34d0+2SDDKmWawAcCANmBOyugHiKpv9lTyn23KnPzYXrmfG9CvlJh3So
yoZBI0dszxPkvw3TJz+xNDG0lScqes8+EJ8/6KZq9jQ8wHHouIC6uPQWDuOAYFIHWMap7+9vXcF5
WqUe+P5d45hG28Mi/3Q14TrEn6eo3Zg1TYWE5PlQjdzKKg+ziRidIVpt4eoxbvMKy3TEhzun+e2I
BbpuiPUXCLfW+tH4HHPDKAscy0mpfadvFBZKyLqVhRhU5NAVfNl/7wR5gdkIe6qHWg1Lrp/cJslS
I0okuqVxkWcVGC3fXhOy2STgGx/2VmjqKK+qboL9DON4fcQX58o1DRa2TIACvs2psGYjMiJpT1uf
FOuXdJj3vtiw/Ujzls17SUWw8FqY62n5KiyiqH+3f5CRAD5gUTah95K0F/DMF/1csqqNbCX1Q2WY
YPjWNmHpFwhZAhwMicFl+HXqCIyBMNcFHPrUkGETojVsrylfhrzRY/7l3s/8EbJSwV+m4i9x387H
GqDBDJIzYhn56tffgs95O7dpUKnydjZOyZn1NdYMr0Ntr+1FpKboLQP3Ivp8PMYTKEo/rlkttl5u
F9bTe3An+nj/rcWofaajNXI77/ikfXU7bNV1rQk8UurkklHRbNhlzqbC7akE1BINxiEVZYjZACfQ
n3qc93Y+XRljt0eeQED4NW7Gf1blSKs+hqerB0jDJGStL520iHINyYaKUZr4RWuNJy4YMB2c+Azy
kyY3JLXvN1Zt1PiFPqWfuiBAndK1QIHX3SYt2F13mfRq7j7Yq/SbyvwrFXT01MX5X+2R00XK/30q
uQXbbdX3kKi4ndOb3CAeacT3PKS/wioORPuUUbLKLjJkDFV1dEs+GvPayQf6gAI4UHysF9puUjd2
j1yagJYrqDl8VHo94/H1WmUSCOC+sGGic84VxNljDDE2iDkKJj9JaYsNhBzlDDTMtsbXLFymo1Bs
FS7d3JKFCdNLLGn9J5lfoUO6AssqmfjbHRyBowy7CIyaoXzex0jY3dPA140PSsvm1gOJmTXDCAPK
/QEn7pXB75hEbIP2BBjvn3iu9RQOMXr1nDGG1Sg/w9qVVPxMR1mU7uPKo0upyVUMK52BeLVVefds
lhWUhFmDtY+PIvl31uoW3elxHFoXqJpASu6wT23aw5rO20tc3oHKYFVHqkVpI2HibKH6Y4vv0/bE
P1J0btF7pSNhnYRkbfr5iMhH3CpQ+tswr+Xe6hvTowkLbfuRCVxgpx2nw8SmRzoc+KtM7SecBqa9
NOZ1lWB4HUD78iDiZ4RBdBuof9KEt/G0AABD5OjMFw7cyYnQAnbvUNoPqcrTIffVPyJVcVhdj+x8
nXnu1J+KS7sWLVRjByfBSrXO+JtdLSVUOlQ0M47PTvDX3zs3oOl90VgHqHD4p1kQ2wIF1JFJqbdQ
RrrjYJ6lyL5yfg8IEWEM/q9Dzhp+W4Lu1Yqr0WHQHNi9cl2mq6uSsKTSZ2vGXgyY8aH88ILX2hYs
vk9hxxxVVzg7nidb2HVx5xZzjmLroBfma/OL3h1OmKwz2Ku31bmcdDSxYggQQl2OzYxNM4Ydq1Y1
iaf/IFWVlZpdPLXPrOzXuxTz8rBqBWcndAjIbvShPo6taM1/nG/hpZPPNkiMqI8RCorUsRZHu1Cz
ZpjNyPP95lyFKPt456SP/0e1z27wNi0Q6jduMxM6t6+jcBgF2DoV0e7Z39saUwi2GwQu3p+uhXc2
O57kO444sXJgt8vJmqlAHUAEXM5z/zQzpWcusfVI21FC+IYy9v62afs7OhQlc3rLzcd0dj4VdWT/
3DvBC2lQ7wTZ9GHruJPQF/1hU0jPQly+d4+N8RbjJarPP5ZXzNdKgJ+xqNYOCL9YfwYdM8xJ5ax+
8kPQbtHu3nWbJcNHsCsFGc/kzPJ+ci7vjPcdzvq3K5VSI1ZCr6Q15auS747NHutY7s0e/oY63uY6
8taRxcY0Ye2rIIS23AqPvPgEasPPVCbim8u2vQqDX5WFOV2mNjoYjNoUKvq8EqQjFwach8FbleD9
b5sj8Y5CpoRUyoV2hG/RwU1IMVhsH8CwNm6GNsko1TqQ2TSGESreN9KqY+FIGPEqzkNaIVDvWaDE
Oqk+P2JJYJzVG1gb21CQ47PhlFbOjQ7s5/xahyt8jvh+FnDPoMajGYavsuX1axkR/q2Qg45B+Ag1
P/zpOnRME4N20v4doMfohR0/Wbo3iXQMUK7CKhoFak3s2tiG8MAvnwqbES+xX3nU3BEYGMWLe5VJ
kfYhWIe+MTcczDYrD6A9An70cDSd0e69G3iHXO0Hq6eUR22XqZeX8gPcUkFJK5mX5HhnUBCVatJj
QnUPojkeuTFpI2x89x8n5zSTSfVPmeOSTQM2ZBIKSVr7+7MkIrOiB0fbOU+wlvST1mIlgQk574YP
5sTDNd6w6D9VyJroQSfk3VJkl+mmsQDRyiDdz0LuMyo3PdyrAgvPucpWjOgJMtDbwghT2BeFS7Aj
N39V+/Ydx0J5W13edC0fDdwZPQGZpMCk8Li3vkRg2hg2jPAiApkMlJNVgRzC9SuBhDge7vhR7qKR
1P4pik1YjumzaiRnMMgSgzuyy/icWCSCVEXAT/hiSgLKXkbP+46AxJbFIYJiRmBMerqZyGmc5Hxx
QR1LuJeKlahrJR7RYTXlnOrILV/n5CckIP0MxailbnR+iT41Hwm8FkXvBxMv229SqIoaowNCpToX
O2suN5w2s3TdQOyJk3yJWpB4rmnXbz/oXXYRF0HyIgDt/xvrFYqV5/snvKPUdiex9Ie1PLvzGYgz
DCZWsH9mY62N8MX/BmAOqN6j/zEj5kLx6tUlmgI2Au0Vt2gdtdhci7T3xqyk/lwceid/jNQ1t3r0
4PE5f2hNlnC12wHJyIbiwGD0dMeg4sOQAIGLm7jZn2Yt0wA06tYko7zMRxCZrnGR6rv/ciQwZJdb
YZSBoUjQiV2d25T3phEdXaJjD215OBG20TD87YLDSGQQAHb2iTe7WTrUHc1lxyovHmfLw2453YIw
DHEDZS/xJzt0FSv1x46cz+FJ3E6MqwspbECkPpfRdQ3Q3XjcpXLN7iCcX9o56QDXZdTKfo4PLGVN
noY+eKf6Xn28z9lIOQ4Y0oi3izmeCq69dXReuZc6neys/u6iy8idmNeZuvVMkl6LYJW0ztVIM2sw
0ekdGMvS7EtfEhMyKZBXgShct3k8s66rE/iKM3YPtdSfcf6QcfaFQ3L4mP39UELpkeataX5BN3PV
1aMdYGjpVwNtwqeBZwUzHWIBXijQx3YvOksVSRTLDfZWAMk/QGW9CX+xpxJOgVgWA0T4VVqPmj2r
HUbSmEbVsqjNS7LEZoa83a6PvnvzHEJO3uDkJcxcbzamkqC8oWzlYAwdz10noXlW2uS363amgUly
FIsBq+s+WfLfsetGwEKPoS6sdHfbB7w7chdT8WWR7QkpR4/ZptV7hWuF4EitnQ0DCajIwQzErObS
fx4y6opehcgJSxntxbr3zyZRuv5tu2Z7d0v9GFmrEdXvnLQR65oqk+hX44viaQpxtvYw/d3eAg+c
Lrj+QyOlEnEc52ALcRTxCA==
`protect end_protected
