--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Z1mRQ6lMgPxu8qw/E0ObSZBWpgq0+fQfUux5cfmcjnEsVt9QXYMZkKUXgUx1sPehXFt1tGFEkxY3
OWietoTUmyRFl2FakNoOmO1z8+KdaovOnXwa2sl8EUwnEbdmfLfjDiXJ3ELK5FAkMVYs41nP8eyB
wQ7y4UvGIxOXTOHymC+aDQsdCI8KaolBMGMI1PURySRjHX1KeDwgJsS+nGHhIVonpginA9icF3SF
w9xdw+D9N/Gmiq67C84KiO1FOj4cGjZsgp3r2jiQaWBA1twuw/deUv0l1pCmcb5z4Q2AvbJ396F0
IoEhw/Az5u49wKcQqbj30eWlZPOl/HbtSubbsg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="j3lynIy4MMQkTbYN4KUxasIBnBuV840r8KHvYNwyWiY="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
CNlPcdVA+Z3Ar+jA35pQW1WpCq+4EwJjbXUz4S4uZVcMFbW2caKpIW7Cow8Z3wxoGHh+aQ+TbCe5
0VOzZ9l9+lMUJH4a4PdSRv6RY4mnA7Ugnt48tXXCLmPJtcMI4PjHB9TtxvJSeJNxUae9CuF+mUPC
TYCgabRxUrw6F4kmuBmK1hdKy2PB/uVejIHfSASWq8D0VqjboOA9bupygdDrVqEhPrYJ1KCv53tR
uV1LPmHPTX5Zd6CVpsNadl9P8N0gS9XUgtnr7jEvJKrQy8/PmYhE6YFfARW8EVDoaT8GqGMH5YGq
+VtPN5zNK0MWV75CGRvdL0URpUCDRGjdcbwimQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="YG4f7HAZ47JnduNnFF1iPusWxyTHMWqssPRafxmSNWM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40016)
`protect data_block
Aa48ikoOoo/JbsjUCdOpuIWkLJjfjkBUO4MG6iQ4ZmVAuiCLQtSQr2OdxUyBWo3FoUZGVNNABQVk
AowaipwCLP6CvMKKQkN8e2LWLPIHCsc6jH0PtGH+ooxiaM+wIKPWPKZxWnQyda3lOdEn99pi8165
aAnQdvuauguzknZS5N1sm3jSTID8+B6DBF8V+W5XWqm7+mqKsIxK7Qlf99PQuynmvFgVgNRqJjvT
2cf05oXyFheLbKFQHCj1+4uoM0Ru/zweSSK/WDe8alqZ0EePiAo9fUuP+JcaUcB+7pfFWWNB1pY6
CvRhR3OsI87807bmhfbzjyH19UJsKBtmI3hUVAzlVzCAQR+IzyI5ZBaejA0tTBT42okky71gkzp0
OynBFhoUBC5q66kzvG8E3IkGHMU3rxRsfv0j2yDZxC2aclTdKox/PGhTnx3YCMaNj7MebQ1DrLdB
Ky+/oftr4YKlojXnojwkaWuA4RgK6WZ9KwDgR7OkgOcfydx1yyrcOXfoRMsXOHqNWmzBp+Iu6zrz
2sWf551bveiGmbZluVJLmrpkHw3KtiuDnWBSXlGTJ6/GvsiaO257VHhJD4XksfKP7OLLBaEiD6JH
iwFGkBgumIdGj2yIVQC8TLrX8Dk/6ouzpqCVRAEHb+VtmnW4/Vu7pDfq4mw7vCBMNXT/p4NLwtce
cZkkBsGgN8b/by0lTvQfmQyGJPjTcVnEVNBSOY/emsWv7pD+YGjfZ2+V13ejEVeh24EsMRsujfJT
ubFOowGnTwdw+0dV+m6AygUEf/f6wShodRYFuSIBS4frIpCAwoGD7glAPzWyq2poGAjHBKKBRTlX
LAuv1g0A/HMYwMYUQqN315BkJcgOQi6tudR/88c+0ffX0a/yzXghgblo6X+xKVJL6x25npxrvV1I
hyZZ+xLBg+3OAY0+Tej3U+SvpMxsu/x2i5P7DXV5gJ06wmpOVl8UFmfPcCdZhVpTmm0SiTvTuYwg
xa/h0EorZTPECx4h0/OY/FnEykkPy+07uddug9ju1Q17HE0uah/cLknwPaXYUOfMy080cUnnZ0BB
LnyJg8RSiRfhfYLRCf1HOyr+J6zT4szd7OXCabvSzXKtYucpKkZlugwyHYkO8HgzmFJtajKfVND/
kVS1/NHTATnqxDxmijqWWTtKH9bj3YzFgPTvlTYxCv22vIT8LM2MxGQxyiZRtqb9kDM7aFwnmT7e
WjmjAFxbS9JPxI1hf1sICpveVcQkL6JFk5PsgRS87eX3SUtZryRBkzJPXLnn6TaLr0coqvJfgIs+
ipPGS062zVRGBBzolRvjt6uqd4nwQmRgOW/pOZKw4NUbSERsQrZTlAXKIqHmBK8/5/j1fjFZGaYf
8Ydr2Fj5VBqct1icROoAtOCcZTIwtCnvTYOm5wZTtvTl5+6FMnuQq8L+k/eEuUAaYKNCcQJdOXtZ
Z8IUSnUlDw/L4nypiXhKq9UX/zXdFlOXSyAHklegoVI0Jy2spCmFVwITbUJqhWeEUoa7pwv/C4Cb
KxCP1OVMxOUinmFmr1/ZdZoUgGY6MP3KmUKLndzRfDTzs1IKVzIPWfStuzkESDL9dYEdS6mFwt5M
vmQGdyieLBByhlGHeJLW2PeYMMp5/WhrQj698+TWrY8p9EhgKdCf8ksxLLP5i3f5IQ5ypQL57VuO
70bn6/xO1BIWEqIOyoL5ZFqIDNrAcYjkj60q6dU++Ox07Zqi+ZzJsU41cWqV00NZbQzHFVOE+G0D
acCVk+uVyWiymfLIdHHlMSqr9nPZl1/dX3il1YdqIiyshkGeiyrM64pRleYqWraYfF85KjfSbc46
uDEwUodjDaH7D7WzNeyNGhk7Um/mN8vb7wehAuIvS+GGrofzdvKkzEzdqMXcmwgcjXvsnsW0zYRY
wfgVJIt4TvVrPDOaeKuozIqiOvyyzzhYHTaPbV68sS9iDPYbNmfTYVjyxHci3iWWoPTMRINrou0p
/6yU8PWfM6FWX5WQzMeYIy0WssIWkiG+s2Hth8NSNI2elsvoSwwkHvYGHwVw2uYYcASpff8luYnI
XEBAWin2BfPysYMF9dThNAoEb5YmqenIyQWsW4/1vdrbYXYCOZkbNTUYJQjgCndc1QZ/R8D0uehf
w1bLHaIHelJQspL429wvLwpT+qALTYjDHCZDzeQcQ7dwHbsXNXXT/j8xjHZyRgGhskND2BZsLmCf
a6oVWFGvyVlndXSv/uUnhg3nUVBrTjWWF2mNXgxVcnGlIK74bf0owkCgZ8m88BF87nnWzCTiVCle
2f/VGNMeotNWfJBcUEMSAdkVTY4MrmfTcCQAtisCwBk4IawA9MuBkv7pMS+EW59e4ICDY/H0+TJV
HNlSe+h1g6kb9bS8seEJe6FWmsjSYT0iKlYFVTm5rxP2LKU4Z0XSP7KamzIRoEjCl5dHIb6fJM7V
JwZ1dyrU13ahOyC8XhP7jZvfaeYRMNxlptv2MP4VMCEkA/7/ib0lIwO9iYuy0UaDhxdFFkKozjCm
b46fu77rep770+/Km3x84IkV9cdWFsCKxT7DpuTJEdT56LH58h+vCSBar+0HKZH9MvJwY2cYPMo/
qV60EFIE4ckw3w6mATR6IJc07HijIfDmFIntDNfQDfFV1n7MAdOFbwH72UkJvE8l7gNL1iV5p0wU
BsKbtgb8NUVv0KAdJMDd6Ni4/5yqXqO3Stz79g8CBBahs4ZRAmmCPgbnA11GYQ0h0IpUhDZsTJ/Y
KYokJlwY50zLmyYAK/LO+xgSM35TM7misbq9KXmakMLZC5zV4KBHydE8SM7wUcqeuZuD8bNVRNEO
WO9BLsuAZjs161jZ13LUaBq5JoVCpmJEkNjDyVxswUk2f03SofIsB1C2wFsExE+zpPgSPihRBnyD
UbH1HzZc1goL4Ka6U/DU8SCqT6a6HcOSv3y08kzAK9HvmTE9X1d1vGUgvAxNKy56iKWZeLgcNyPN
4+u7SBVaTSeUT425paRM1m6HH4xRtoHB5Dx6WQkT94Z4MBnuMKtPh0zrNhYB+OIL92BWvmURDHtm
BnyZJBC9Wr6xja4oj0tIYJTGIV8W7UOGPWFtHCNAFXPOG8rITR56Du4eQYvNMqVZzmr9QmjhJYZl
kxR/8xmtJtVGYOq0nVcPOsnPp8q5wz5IaKfz4wjXj9L0Mhql6OCMz93I5mfe3VamDPOjtlLTDiYb
c/fAL5cd/lPAcFHtCOyFf5Ngw2QVMi1UhlnQh+mFRsAY3mSqRoSHsiqyrcEo1ouR7zNvvCHGfcuu
mMbxZyVhRBC5p+dlVeyjFo/GY2540YgsvpAeQo5N/ZPZa+ohP2tbDMQpd1FQVJ0frnN/x5HQWazE
FFYWuMtCI960v1bjAvk88y0xflpk5hOG4hRaOKGyfs6AZOjqlu7aIgpskUg5GRSfGKa7ojs11aLq
bQhuSboWw8NMWAD3prOCA1TiwYT5bZV4G/lsN6k0bNO2boC5M2ojrw4yX3U3R2G8teLNjO4tZtyI
6bYKKIccVce8Fl/ZFrRKgC1GrugkQhZZGicrlU/eSON7FGnO1HHZQMW1TSmWk/KxSerRFOz0tCCO
+XtOuDPQyILSMUbcHO+KDivoanSUtKZ0ZroC0Du5yO8CwTA3vgjjylDcIjYNzoVTo51/wffRh+eh
p/XpB06TdLBD1+EADrySsBHH+8YZQOd8l7S46ao9+/c2N5brOd+++AI+k/+ZSiCXD/Z2Z/XOLpD3
Dd11K6OqkhYnqPWTyQZ4hwULOAMQco1y3sx70VPnWYZQrFNEqwwLRhvEMSb5x6S5K9XYLploMZcD
yU6TRp1ihJZfaD9gRaH/Eei2OHJsw2yEQtZBnyeu7dhuVV/TRDGx46Ol5JzA11anIjieS0Ni/HcP
6L3LEzuai0MckExSNlVQynI3fz1eQY2SLJ/MOOS6unjQCpWtstt65U4k1KNjweeSB/1mnQPXmYMt
s/R+xiUmH9ZcyIBaA2fkQd70ps1GY6UsxaYG/z4M00+lCQb0UOV8NpWL1rYQMpk2ZUykBYF8FEzg
zvrCI1cR7j+pZxf98HrxW9BfRJmJWkyWS0gq3HrEU2mJxOQ9IO9U060uk2IXKYO+Q0UjlM5CDFC9
0/lnRxgcO63xG8jyB4e+bGKhR7P7YmpSTaaROmYtg33TPvLaDiuJsFgx9dUQ+WUkN3P6wD9/v5pS
/+Vh7y4rShfF0G37dY/HLimpCD7+QY2LAoDKwOrw7IAwkIUOqIHe8CdXfNEc+9K839dB9ewnH+3U
tdb+gP4LlQxUZRDCLEcNTAjpTvnuqfNBjr07quIY4fgfMNfQyb0+MOmi1/zNtexGakzEEGDrOZLS
Hv+/todLEocOMNApQFUrPCVZidRCgpwSO/oOqfGDRtB+lWR1vKNaZ5QGPcmfKYs91gu0Zjc19Kp7
xUkuuB2F8GdKwOKVPT1d9CFTmOzveLpmSOPH44tv4DBMW8seG4mY/fEljQ/SmBjFJ0wiVGL2OAci
kmugUUEYaO7FipHBthBqNxU0fDtIqg2j+XRCSTYaUBATMEGn/ThUi/xCGJvBm6EyhUxieVNxxGhk
+LVb83CIZVHdds5u1eo6X/t2Zp/wYWbMT80JwtarVd+2hiJxvZSyYd57f5AaslAE/T/9nv/uRALS
eHT/+Jwi+UFF0AE5DCgPmMRIz61SAtELGKaxUkzCHp2FL+9pmsW4X9rDXbKSb5Uh2+V0C7GMFMqz
TX7nNlbAoVQVBBVUEDD1wpDoZRiM4r13T/7CzULo4ftLWC5bclXrEmWmj0eBvF+MehkL9jcBTXLS
7h8c05SoJC3jfc4louBefyHZavvc9tElupvTyOugFt+1eehnTG/U6U66PNVltwQBmO4ApwJkVAGk
8zSfvbW8NjLKRPMFs8P9FLDMRk2ra9NnZwUPPjPmTrDxl24TdRslgZuaVnvwfdhP6sj0QBKIDK28
h4hIjZop+i0q1Nym5kacn6+TL5z5cUMAkvxpWdX1hViyvwxQJCgXmeTbpU6WX02q6tfGIvphDsUx
wLVK9yt6E+eU5HcCa/sNHFLxBJW1rBiDDSHuC2GZV4P0NVpN0Qp5MYto/0DkuIJH66uitDpS887D
UaykP6ZMfLu0sFBXHxWEDTSjRhwI8rsxBOJN05a2yF9Dp+CRPT8TU2GLJJVYeUhhKZcVytrUKA9g
IfpI0e106viBC1ruJ47jrOZaOJ9Fcib288rUybaXLwcSJZ2O2fRwDNr7Gowbc5m6UDZ25tmg7lDh
YFquvmmdkT4QlUXAsr8PIUaIoV1EioKgUpIeY3mxKWf2jK5mn6/wgTquClD1M0Ka+qEN4ReKaKAl
wCBEjfejUigDg2BLy1G3ecp3uFOLtuDSdrUxD0Kmjwhg3P9OgJZ0exvktkhX5fKHv1F98AtDyv5I
qXD6bMqwjIwqSyq/kubN6nhA6t0NdN8iW4eY1HEQlnEd2fMeGFEwtgCXsTO9gb4EhcYHTm+VwbvT
9dXfXxTAU4Gl7EUmbzE4Y2iOx0xTuB0Z+FdcARFg+1NLRyCn8YJpCLPg1CHhEX6tMmmM5JqLskt2
cE1dyBfANKOKGhq2Ocj3QHUU/0zruNo0zttun9AD3J5AmmTLZ41sRaUJIfBisl9GKsWGCn341F2Q
WchuMHjy8lijEfkuTr6i7IzH/hzPRO3toBqvKA6rRXknRaWr+Hf4fQlGA10PK4qr9PdAho2LtM4T
GQZADGJCaNOalQIUokNVZfNmspMl8D7yRDdxD3iQ2gJVzzI0vf1Xrgbzbn2n081dCydyJK0B0bTW
VWIcT6NqaWBj4ruikx+4JYStFD0RQSaKMUS7Kp36GIJvPD33YbUbPIj6Jl2nvP3FGFRQrfU0MSBs
eTA7gsX+iY9L78xg6KJYEJr0HiGCSRfNndfFaaQrK+sHBikIj//w1FCGNcKXM03129hxf9R1JXj+
CgJ7xjTos+mRyAT3NvGR/TclGaU4TOlsC/Sx4xfruqTT+ViN+XR64stKBWNthbjxyib0n1mahCM2
FZd5yR9I1ZR98/vL9fL8lhH8BnsgG5c1h/PoW+asXzI7D7faW58xS46hHS+l3Slr21H9AmBBp1AQ
k+3SFZA7JOpPBirgSJwKvR8+R6mz7sSN9ZZ6f3qQblRfadbZ5c+W2f1vkLybMdzx15gBKKiWaPvj
wNemTooc2sCtxHoot6uzikT2398fmRudHlbqhXNS5GIvn1MEp676qQPS86f7921SxzmdU27gulXL
GuuxTvap5jIScuXoNbE8uTcwq43TVgUSLnm/9jtkY+IIaDqDFs2HlBYo6QhAr8zci3taEAuDJoom
6xyjFfIpKATzK2AJOG0kETLrfDOIEq16AgfSiSPStedvns4vvEpLfGbUWRAOeaclVJmgc6DOkSIe
4KwbHvopI5oGyBfJ3g4ijfHWnO7c8XGbWee0L08wVHe1P5VaHaTdaXlXBFH1m/BTE/amdDn2xDD+
i/lZsjav0O+JXpbnRoe3Z00lFpbsjldUCN9SXB1ThOI4qw5NSxW+ZvY9hyfFgKzQp4mBtO0dXhtl
5X2cJtNz1n3QiiNQsXYupvwuO0mnYMh0W92kvglYvjTi2BTLQ+e6J3QoOS36uCc/2VOrE0qu8kbY
SF715FQ2uPY+Kj8RwLtfY5ze0Im/a/73PzkAwGjPWBjfydclnkvUCXHoTAB3b+/yEW5eGMoq7FIf
AfBu8V1KS37KUzdZ2a09KSu6y1labHPd64DgemlmiYsaHAuaIAIBnVskHcXT0y4BcwblzDY5tPZv
swjz0vaKuxf0Eb1v8JwAh+0JcUyQ4/+K+6lzhnmTEg3Jyqz0Zk4wuuPGGxCgvVMKruASYVIu+WMf
K44NlKM2ScD6U0FnnXTelAOPV//JDtVnZYKtWVyDLVG/4hH0YuQilXoggHNKXYCyEgqrzs2dC834
vajMWCcrprvYoI7Wxykf0jpd7oVy/E1g1zdcUFrV9GvKdRAgdOCj1Oux+Zv5pRtYwrRNCq+Z06ac
aRCz3FRRvS+bgBRVeRKaTCqLmYiLnCFoTGH6MflxPjiWsfOlje4ND7xYJRFIiusAXkD2YCt6/v01
LuyYKcbr3+EJOUpJVu3iijBIF3eKt5jt9/bYB2adAjn664+y7q2R2BBjvnmccQh49Z8jUEyV/pPu
LIsp1kzyNvSHMWTG1CZX9ULYbh9C6yDozp8vEmqMOug6/OTw9nF8w8s8/ihIutNcFrE79xMdsS95
Pr1m1IBLp064sTvO2uq0fv4ftXrSCeokYPC3INzWPoq8JVPilFKtTQx8JzOzMyovM1FWGgzvv3PP
ViN8Uw4YVeElQAF9axhSIqGIRLtRb78qmeMm5cLgEoOAlRz6I1mtDcemr/KMGWvbttKW2aebD9FR
aQUvNB0t7WDxtzbGo3w7IvkKGSQ/GBNwrKXQae1OXkABfCHrYOlC/xzRZqOuqfJx9egECn90XPiJ
XYI1hIEgd0aeWdiT2uJhw8jR8DcD9EUq1qPg+foURvvKvjJp5CmI9+0HE9aEKTygvjK3tOs4PSqW
YdKtzbFM2HQ9SweXL5XYZl/E/OgYcKykfwNeMuM2ZSUkj6/JyAevw2aE5C47Wd1bd4Vr1c2rzR4A
rVrFowNZnhK/jcj8QcgLiZvGNk/USjox4jZ9S2SWBPWLen8CqErCmG7vrlg9rmTo/VooeXN3SQxV
JvTRg7NHG8pGbbXGPIvuo1jLP0zGYJtdgxK4lWrXr0NGvoq9cYmWWKRUnwhNPkJb3q0Hmy6x7aL8
yqZ6cPoXszB/Z44BLtzpSEuEhIbbttuNk1eMMvEcih3o8pohrAtCOeCLz89mtihKrs38Xl/6NAT3
n9x9DgwTPjGPgbDnF5+zkM9zMZEOZ0/f+AoKhmPRsbjFDKHyDAQPND5AWSWnG1OWkJWYMn595LIc
022s57iXJ84XL63wMjOQ6b8vzvGqLRRQTaC8frK8/h9S9sV3AIncpwLPGDWsKE7pV5GbuXW7wdDJ
blyTiuAgXKdsa9qQ/SJ5MGmXYzz9QpmfLgkUT3Tkg+I3tmRb+9SbRLOjEWpVHYf0UMmLhfiZj1vL
4rENKONDfEYIIHFw34pOX9GJ4DeSgGTmpQJdfJp/ns+pTM3R7eznUa5PMs6TSmK1Psbtexyt/QId
Wd7qaUtiyKK/nb+T8Ou+EhZNsxRtrOwItbM6G010+vhn5jOkS5ghd6qMXy1OIRYV4pGWxtPpDOn7
DD7hQ3rP3bBPTSQYy2UVbC7lDknQ5a+wwVCvLZPKkcQaKcCiN1izU2MAbZ39q9QjsI2ibxEFXAV4
CydMfPsrdOIPQKocBuDasKg1L3T8b58mK+2TXUuD/gaF690UJcyJoatXvUkmRCG8vKvaZY0QMImZ
e7hGp64W7U+zaY/NgkM9YMwrY8o/s9bEEL6RPGlK077U0bH5VMCAD6u9Cm5I0MQVyioZPfUJEr5h
LhHjesW3L6wgIsTcyp8NKoCAYZ1liQv4pUUby7dCO+qlqHSXTGEBntEpUAsI0uIj4dstvsRoXVfY
SYuU46E4phDH05kTQenx0Ci4WHcIUhpWTw/IaO901iMoBOXG7i6CUmpxx+ttV4nL5f77D0qpaYDT
R9aJLtyKd02JZp58Sf4erDak4okQa8CiN/Uu8xu5v0ZMr9qsMqXD2M9gAOszmQuJC7FdD4lwqekt
XpIqE/F5PUrllsFeFO0LXWT/3Rsz3Yh6l4xdczFESJAyo1fBnwrIavA3QmiYRpjJ4OZyZ7Czuh2x
LZM8R/haE444TtySMG+4H/SJapQh+9Sn/x3LlEeWtMLWbmoq/uLFt9UO+uJ2JIIXRW6M7lp8Jp+L
FZThfF7YGDOXeg10qohJelGmEflIp5dTBfDlvU0Fe4D62jCgb2TgCDKUCCnHO7RQbmKVMx2IoOtB
dX0IhBCQbx4/PlA/sNGh3GVU5NJbkLDF6NbxbmEhnoEfnMP7fm6C8jsLr+xOtwCV4kaLeHuRYXwy
urLzxGXYcaSkdYTIu7qJEv/KvYSjqhMmweFUMPogaI8EtjWwABos9pKtiPdclzaXANJ2y2Sq+N98
w12SBdXUP23AtpUDxnisVIu9zFVflb4YZ3ZGkjkt9eVQkicnse62bWP3cXXlZ3yWcKi00SV4Fi4w
2R8RbLS9YfO+FQKukwMQ85ZLWzm/QLtpNlJssL0fkyccBPPWw0kaS9jK7hlYCZ3BvTgPuTitORtv
Y794wwV73xXToZkhARF8JnSOhh6b8xJXaLaicZPkUko3xgPVHM06Njg0lM9Oc3nNWZkAdNVlK5lT
0lK9UPYy/B5aCUeCOApthX+r6GaTJfh+E3bWY8ScgoerNmqVabbRsjW+uIG64oRJrtLWkZoF5b8u
0E5b0IyWDXPlqp6aMjjNJRCvbcpU/3UlGC8XdOTYAbanpemKMGHFfuPw+3T/IlHWVLeOBtHmwVPG
zyv44vpa8J4X+AdWB+39T+LoPVm2fAMqjNDCvyzHvCn+7QFL1IMdjuyGeJt5jesuhW7JhQ2YYFSo
1IFg2jNG++TP5NZwcOufmb8nL1l9FsfrYqKXLP1Az0rz5PoTrEkl5eW5TfKkfUCjku7ILsCbODMS
5zaU/Mx+7wBJ8PGWxtu3jF2qHGKg4bijHb6E77mSZm573I3XLvOXDKc/Yufx3SAmLCIgw8s5qH6G
IFlfzzh2JilLk01WHYtIgNbqdYVYmEA/8mttliA6yhr3s63McaEJVmKDolrNvACkcumCeT8Aa471
1uUvRF3IlnoqDPQuxEMe0wzT5nbMclaJS8nHp7okM/90zt7TeAaaSqw0jpPCX49gZljMojlN6foE
YbzPcvjXlbZuOlesSsvcLqu56XmcnO/LJ2V+nHFBXGYgZgnVv5OYCWhPeiRMXcfq60P+2WqSp/or
Y/0X9+4DdOEns6+kTaBgOCN/P64IuXy7dXxT8loir9h1sXlaTHh9drDDLbQaR4JvlYWB0LrtlOef
LsN6bvnA9WWsT1Eh5Nrmi7kMzdPNOMv2trUS6dPwd8gZN91Nfvj06bh3snxALWYyCSEvSF7KBAus
OzPKpvbC5eBir5vCddZLBY8SrOFJ917BJ8ICuXEj2FUmRF6n5OQmt48vPotL9c1cawOsEO3QYmXJ
ftjVYbJmTyNgw8RcitpCTsdobi8/fcG+5x5qiLV22MYhJkO6/pNmNAfFFAVOH6p5bQ09Jtrh2Hs+
yGrgowHDw0szd+S5p+oyCH5jkGgYR9pGiFCSNthoV31NEncCAwK1FcBsbyvAv0AsxJ/Mgie8IetS
y1Gkj4KB4MYWoqAkB7HzrPCJVc8XP3KjPsCmDaG//crru1ilY2qtq1ObDCCmCv/iMRqUcXSbBsBh
uw8Ligl01izqOfYrdDC86sPT8jM1aD7hJfv0U+PUuIFF6IpU7hRdaDPNebUE5R3LxFceBChp/Nxg
BComsTWZPkJaxkewUlBSNTcYwGiaPjd2txYOX1wT59Qv3XukEQeOGkLo8Auf2OqSLzTbTW1iKSzL
rPOcRZxpeb6uZQFYUaGvG4iqn4BwYPxcthnv5wsNmtA5f5YBIkH3INFpvwVa8Jb4KxWh1Oe/HQzi
Fs4BvIFXdcnDOHaJv3Bfa+0RLk/mLmtg1x19mWinmYFnJl+KnrQXTDvzVJ3bmghHHn3lebXTnlGq
GEwl56ezbGd69FQyDKKQhF5uMfAEBHOaOoeVp+jXKDim5Rsni7SWtip3zDV8WaaYk5Z0YX+tmEh9
5rLd7U9xP/Ekj60/EkYD709UDI7oknFQbjOpgEffTwhMQK074G1I1AiNEJPBBeFuCCbvBHcwL8Ha
01QTGZgp0GqAskPfPJA7oKMyHqYCyCAw2nV+P7tcl0RawaWL9flSRAvXD3sWdTzPKM/LOsM1IolU
NONU38soy0CwhtSyvT58RuJbFiie7Yg+NUzI57zpYzFKynNnDdNrbA5WRCddgrKiQsUO4RHRd3ri
zvKJham6IkWLfpGHicNQgj+OpLxlLUYsZFIMVYi81t8NpVNuN1RFgmiu2CgjxsEgkPPLopRuHH6q
TAjWz0jXnLJVB93z9yWwKXnboJTY55FnxZEaPUj3UkXyEYcPXyqzn6uqsayAhWWjbrM8OhU1U0UC
EpnkjdpXmJ0KcB1peTGGYzN+UhU/SRvomMWDSVp6PK5Vhf+5PBtxr9/ls63vwR8UUsYCJKFbpl+F
CcAW+ct9NfqxCF7g7YmiWM5Tf2mwJgCiUknr2nult/U5TL95FXjPdzL4lx4PmBuMhigUYHZSuNZZ
PXmfElwrCryOZpsM5aV5JGhiuH2+BDbQ5wxSQHxmo3hPBygKCnrCT4kB+Yn+mKqVIxULhrvznnjr
Am148QVcoCz9PJeu/fIc313OYlgZSuaDvPD95MztuKGK35E8HQP7yFStTh0PpBTpI52xRZKNNIWN
hTPsh4LW9DWvdjaX1bo/vSU61xcr5/lWnhlUzB0892d+rsEcrHQ7+5JVKz7iip10ofmc5z+RJwB4
/TuOdMRimR7trVDpnbAZRKA1PF6QmnItCd6d3n+tPy1/q7amelSXB/sLk1++4yJ3HB2qyll494L6
i1wzM8EeqLF4NklOzYrAJNR+AFAcFqM5ub7ytkRnOcaPaPC7aDbo7sNGB2pxXni5oHykHSJqD7WI
Ul9xLBYzrXQ2G+LokwwefXb/fJpuJmc5pUAaxK0ZRV3M5XHDTYpM185g3BGX/kkfCucH90PyFUkx
rnXym9EMUX1Lh3fjlxFawoPLuF+9tlhBf76momxllh09ClFd0WkMatcWq81fd1O8QNOIkNzVcxnL
+zm03mDN/SaIzdnXW+eMgNNRaUXDb6IYXrySx57f1Cj8na8saVFyEHiRNflzp76mbrTEUtPHdZzQ
txA4MVPiZKFxoVbQgOLp7xcDLLPBo0bEFxeJxppBUyK6JC3tgTe8NGeM+5H+RR0ckat4x8Eoou6U
XkVLDdVX8zj3H6ZlU9Ri601PY4b63TD72DKbK45EOeZu5JExfRnkGiwvmZbAufrtGQ2lPHL5iVTA
h890UmR73e/aKbec2B2ZXCTjCYkpDycycSoTP3zToICqs1+D9jKImKv7ECztep2TlgDhZ1quiOPE
c/osfl4VEGOa2bLRKh++StUJy2ssnWEfHJx+q4ev7V0PZgTPbaNxqCg3ucnI0z81OFlWWlkwy8xQ
iXAUY3W+azv3rIR02oZwyJZtEpsAM2oBa16/pWlYxJrcyPJx8rcyVsFJ9hhE4FcfswbHeWuiaH94
aqXU+u1Rgk40QFgF+hC9+Dw1ywF/YvNKlUc8semtASsEeroMDZjzexXdM9iRTRlUWZj5xfTq5uTb
TmxPiagdQpohFX89r5MEJ92lso+O/tRdTjeMoNWs+9gW4Kptkb+0QTphcwVgYKopU9nQUZ2ItBlT
xx5Wu2tPhY5V4bukYECVW9l4FV/wXg5jQhPUL2sLvEinAjazgm3yT2HZhLUwyS+twrcGpyByC/74
q+Li0YzJMcekrXzya8tbeWI0xX4eLZ3uT8SRYBd5GQPcVz6hBIJiIrmStkrK7RWGNpEsbuJRWrtC
Stc0IkRAbuEnLRM55Yk/3u2GCkX6k8AbAmx11b61x40lFyTpnbV9k6GRNXYuO0lNFSfIr6d/yddL
7atxqEvzfbTFWXRQCP1ciSJqXTlxDr/XlsBzcKRizPQ7cLfI+RZ7D5MR33T7YQjKlJDThV0vxSE2
ky9Vq8TdT9EmOUxX3RZ9oADaQJl0gz/VhVlxAHfJp52SZUogYarF8H64F/rPzjn7hP8Chh5D7hik
6T+JHpXXxDO8UA8CSDpxWzYLniA050FgpQk4EObpxMXxWV8shhJH9v1GG5UrUzMNMVvx0rLW5OTI
W4WJC3Lsu1V8IZmzbni2op/D1i6RUX4b7uiau7ygVlZXB3I9qJTtm/8OvggVeOjIMZd1n6rOnnDT
I3PBmc2BEZXu++zcHzS5Lmf1B2g5EbClQroQ3DKBx7ZQq/DcFjJfz4QsV/vAxWmqjHNO6F1mXvP4
RVsUY/4vK+s/Nf/Cx+uMuKDsolUl2a5lVXR+mU39iX2JHhDiORNhL6NTQ9XvGJaaa85hMgeeXzSw
9LKt/daXX0b7l6MTgDp7/B/ghn20Cc0I8DpHE+YhtU9RdSxh/lmkDph8SbEPd+kFwb9okJVdx9ry
4PfapSPkRek7Nn4rnet8EDvv+DzxHn4XuRMpvTau/xeDGIwjUjrM/a9Jw9hZsD59KsYdvqKfsLrj
tzbS2Yp3tOXBLo9OhDVFMFM0elexu1EBqyBTGHTy4lB69emPqq245zmMt35hScr4TIKi5CNfmUqa
rdDXGio9tQoABqHg3AMzBsC4kWB6pXYb1tJq3VOdxF+PQbVVso3Y61rtVr9gpzD9+VKWMY9idH9c
SJptTJG9lN+n7PPgut5x7DNJcTT0k5S+s9IZIt+If6jeD0sneSRgSfIBF77qReq9anpdgtndthS9
0LiaZ8fQUjrWXdW7Hq1idpaaKhn0ijykXDYQ2W+bl+ntfuHbM4v0Zt2rSl2MZBtqdRSR8m1gGMaw
UlUg7MJ29hyawoNF7lkF6UVGdatNkZxIHVSe4fpSbV4iO4ESW2wGVFvLiNgrUC2grZjoEFSK5v3j
vJ0gBpycvs+BEbAT9WiE+idCKnFNmCasA93mC2fnjSYXvtEk9xjd0fTDPCnDXGZgV3Fn1WgSf3gy
6/nyZjTfB6VzhCZ3mfdcNTZwWpsrGbQq8YddeMAn4P/TxuyzVXIjaTj1DRSgRBdHkdlx5JCIqRKC
z33Ve/NK1i/YC45HBeQxlQYTAFKhMFCWTF3pKyrtXjR27fLxcfePZB91Z3B9heSYwL1J5pGzHv6L
1pPvs3kFHMVaOZvffl0SvJF6J3tTzoQg8Me4SaKEfMQjm3dDcOo71pqqLzj+1XawlgHwW0slst0K
Ozm9UZ9M8gyOhn2+o+XIURlKtCBfL0UTqbdwyfc1xKdUlvGZ529Ij4MIe3ZcXlWmucSnhT8fOvT5
kb6miwhr+h5W3UhJzRP2QxABTJkoWKZx30ldDUXbNY84LIB3CTUaoGsZJwQsVspzM8gEysVRaDgv
J61gY0pas5o77JFuyXuAdmMPJTDfZs6uvVU0sCWVmPnNUevZ16hwMQ15H3uaNC9pnqrpVIPUkIMb
fRdvum1Nv0dAhUDeNniYhcY15ndixC2jrRWtijU1vAL/8dtXSCNRqJ22z6SRRmkAqSnChRBAKMFN
rw5npBsE9Q1ffyqjCqe4T16HbBFdo9UY+6hNg5l3McnRTk8A6ugGdKOWBB55X1fSiFRxOSjf+uJF
nWaGC7AwnUaoadA0DW1ckLj/rRxYmD3sCmyEiA9GRDShe63pQCnx3pEuXXUqgrCVX1wUZFT9Hdhd
9v2a/tQnYxaNMpgshiDjWpXAu176UfylpaZPWDOgTtwlS5sStUp1NfcvB0aVMQy9YuogXIuJGesX
yT6ukRKEmXshU6uzHehOyXuINcphOf6R/kbgDnXhal6JA8OJL0kk9kuppBu4SWr9q+D6ez0O0+Yc
7LUk6QBtVCrjC48roQP1bgn9wBryLn0PiVicDeu1XoEfXJ1+9Xp+geo2j0aqMkh11Ejb/mK4jL+v
POBHSiZDoewCeuDHqRTjcx+29ar6gHxVEOKeuICaDTYnyOL0egIlFwBWR3ks5VnXw65MHrw3FBKE
TLVgsk/lY568RnDz8ntIC5lKhYh0IiLRC8ak+M5zRyxIK39ArZOiWEvBx9XIILc72qvRg2vcVOTE
7zK1IAvuWqt8epIWGJ9k2MUSD59H/SpEf3lBv/qnSRmj40VRTL8KFJiHrT8jTxornhlip3nippsI
lhXl+dOTtsrqYr24XxbwXBmmXSZQb5k0pOPKP5LPJgodAon9++rWf2mwE9RAIFT3CqiFJfWbTmF2
EXUf1ss0FQJGeBAdlJcrpTsgcH/PWot71cja7ZNCAYHEGZZJJAfl4jcm8QYIBOOxB/Bse7jU2A8T
LMtqpzNOZrC01Ft1z/o3n5r7lDMpjY/z7qZTUZTxesMPUpNy/ddMcKH3iIr8NXeHaXnJdp4DUhN9
lcsRCpYuGh05WRVIuE3c2IJNwAf6/fpauAZPlLl9P9od3lfJW8M1EzkAweeZ8o8jH1FwOvcifx1R
mtyxpAYJsY928bIJMPEFMS0+6GudeYcqtDesBFi/OKngcxHCbOgYTs6JEXSA43BxJKg4D5qm8K0F
Nbzsy/WKzN3k0pe7CDoyePdlL5SFMARBq2viw3EKgYMIPGqJvSwvzdaeXMDeHtJvRUkFyadjY5aN
jNgRbMnfATc8yifSrttx92dbkAlkkPoM6NoRu7daf6l3Ce3iRucp+cyoCGTz/FdCdKk6zg93lDcv
5E+ZI2o7VZLTkMb9jaVAqLbv+G9SKJd2J/vTqWzKn6TGa/tH8Tpn8AFfr50curb7RGHpLu7Cjsov
Yd8PUhKT/dAz2n1sksQT2RC7i68iZXlclIgHyQRbz/8WHhNSL7Jb207pzBwbTTZN/bzrnvwWNSHX
5Py+Et/h35nh2jEXPTu0G6i+Gr08ptmyrDO+sdMoIcKqan7wHgOfG01VFLh4JwBudv8mzh2kj11z
CAPJclne0Y9CIbX57bXOwzvBhBg1o+aUYXxgdwYlSTCgLPMhtYtg1bRQZbZ9UbdXnVXieqstuUx9
2tiVaVOLMF2Ekh+NTbtSlhMD3eRrZQu+q14Gk5AJkrHDiiVFd8x9ayesF//a2KnLof0zwkBuYyku
UYwUMiZpJdoSjTlxBWErXLm1CEFWtJo0JRMnWorgmW52Rv6DkxCm4GpCzYnsIPFpSknS9PDpb/6F
TI6H8RaA7zGf4gk0DiT7flPirSsfwvkuGnWabaMMToWHZB/qcpJ/KMbQ/4LUt5DTF+DPeWdeOSeW
8BhyNWlCtQErvUGXWOnAf7pmSxyMjKNZOFNT0XKvTA5N16izV4X+NkRoihI+ACOpKYvXopmeZIFl
xWTkehQQuFd7OY43Nq8e+V92ASUTmUjxCCmiwG+59TjxdG75tl6g+D08aVkW3IV6b3nf61Cr0TCM
ph5YJp0Lgk3CgbHD+VkmKGD7H2wcnXC0sSJIsyWkl7BVYO/2R8/DPd3WNch6RSK0bjjNyhexOE+g
2ofWsjiOip66/Ujzeq9CWbcX3DBn6SXYtOwDOF+G2OGaaxYZfLUkVZUTcUllaJZv1SFo6vtXgwHX
AHKnj49CL9MddZiIl8HWBPNOAhS4i1O+651FDNFpMuSowteXl+ITa6XTonpkTBhSH5YAIfVPYoY9
Ilr9kuwJp3CYcaOrCN0deqOXjt25tP9+MLtl/3B6m3gEI9Ftkyvxcp99IBdyYuH5Qv2WrWD0/uGE
CK1MpFiKuEGbHSKmQ5o7Xo1KLLSp9pWKnyLEuEhW+wP0Ck+E6lfiCADJyQkEie8CVpEVcH8gS2CL
1fnoipgK4v54sMUuq61nvMFiYx1/l4rTQW/9MyzyYNIj4TySHW+/vZqlMxqtrEGJJWuW7W+DoDRO
N7PxDwR6ecUDii6L8+Xp5ntGyqecRG5vNNTXdZcJdJR3FGvmeVS8T6bYHEKeoRFo/coux9wPv8WG
GF269mNizSI4YqO6eP5rx3+R3qAGxx9CEtPXG8jPq2h/BZxWuymLdUhn9SJWCIJXzluzfpHYLJrd
LBBV4JAmfJYrWmJPPwveXD94xirDje78spdS7lF9ZNxtyQZHiegL4RNFzCAO3zBgBCrYnyiMANup
VkkRd10bOzDtv/xVcnPZz30d+Bo7PVGJCaLUAHVAVTMidA7ScbaAJV0/ig2l7YLY2HNzH7NHXVGA
BHIMAO2ZW2TdRLk2F5a7soMgi+GoWkMWSvMw19iKd6+GfBvQWfv+8JbDB5E1LS0F5XegDkM28yWx
9M4LRfom/Xi3VmEmFZ2d7p82rYn0UfwUBUirHFPAIwI0/9OMmddwTpweCRH63aL7mjv9nTilYV1m
C8oh8Cr/jBdFFKz8tgryyLz8rscVmgzP1QzJaoUZ2Y04lIi7VY6PXCdY13aVu2UeEw/+RyI3loMb
Hpat+c9u4mrHjszkYNDSGlKZhM8WwwddGTTVsEbK0m736ZLt4s1xHQf6Le9b2jCzgvTK9USxgE1x
fPdjyPzdOBJxJPA9FTdcpBB1znB9pX6S2jMufQlLz+70leQQ77oG98YFmUsObsOn9eS77tbwlAww
PTIl4XWcfkGkunSg6BX7lhnwWfQ2Xc0iVy9ZCnnRFiM4J3Nkl+TKAB+zl2AxX4Nz6T23BCLL0hXw
YEWqWkJGJEsaUGv+x80lYLB8UAGjNuB2GF3KTUz7Xzfhw0FUUNkDEIGYKw8b+HnOqeCxavh5oQsM
f3iYHd9QlZpMg5HHykzzVSOKBIqO2boOP2RXwwqzsX61fnyznyf2NPP0e+T9Alj32EVUEZzOS42V
U3JIJ14iFdRbLQ8fbdY9fK36UGN0M65AzRRQxUuxaeORVFzKyV4XRB7IWXKl52wTW71oRQJpCb1R
QtEflrKypkxELDLEDu9buYb3o4xMelURw0uMk1DZqvi/kmzo7g/Iyb1DXcvjiFOrFan4H0sn0osQ
WcLFhKAsCQnhh+cEMpMV0oZal5iYoIjW/SZnKfpgVMjQ47n674d5pHPoMN22e0qSs2aai+4Aa9fm
SbXcS/X3Lp0KMb7JfMLYAgvtmGUV06kPbNbMvTsPb7gFAwsmY0mTUxaBd7VNw/XzFqedMa2rUCb6
VY0PMYKx5yJu6U9paB6SpG4tcCTyRH0pYQUTik/m437zKvNNXhArUzfdmBMUF+m30I8hYTUxFb72
c5ZtfKXMwRzh9DfDBsormNlclXizLpW4X374yK4elVZB5Sobe+9Dc3QhIis4haiGDqMgw4e2w4cD
zD1TfztMKouDe5fy+2XAYrb2+WrbNbxIyO5DgKKpkz8ucyuj8PUiD9YSLgd1/NvLQmAx73ZaslAN
nnxAywZBJfy29NXATd5CRM2DNdpeua0x59V3V2kYWNGtNhUBfMKnpZQrC8/ppZ0mD/LLzfyGbJWq
WtaQyISr+4ZCTt2l/JB1h++FFq596GRXF+QHVbdkQFiF7nv8rzaUlzaj4Rr0yOIvNc8HzfYeX7U8
uKrHEuJtgELmfKkgPY6Gb0vuSI+advQP3nPgSTHySXw7w6T+TThK/DX7tV8U7nzApuoqhpi+DAlH
vEvoVSHMBpidXGwQf3pLcKqFs+TWrfDP2WaBSLTiUNyU9c7AfQX2soKp0qhHKzjqqUwlF0YyWCHI
2woL+k9/dCA0Kef1kCHc0DQBl6BG7kpg3aDed2UevnXAdqw7Y9STV/G00TEgRk1MXpp8bXOEPX5b
EfQ+6uTnno/3VgeC9xwdPMs6AEOgolpu2u7UF02VRYgWdYRPCVAe0x4LtimDuQx5PO0/hdo3h5kN
Z7r5IcpBQBpimCIJvgFHPBHCRjT/d2qhhU8oVxRe60k86yGLfrzTTOlrCd9oZLWz1SNqafg/jQdZ
pmWKueGSWP06NgKfvkB9r1+kHpH9vVGli//gtsEDxDohEmbI3ytjsqRzPsPMUCRev05HEe2gYghJ
cNvHoUX0zawSxHlJByPZT8kJkkTL10Z3iIqN0UGACKGhzRrlre3SOuvjcrpX7H1cwl3TxBnQRczd
APPkNjEzRTyHn23YYg0XZklGQJWq9hnMSruaiwVoPvlycAYvcYEKjq3x3o1fX/rTwOrErCPcjWRJ
mmxcyUHvZrE7GsrHnwQxk33fn+Sz600AP4eYthw8kjrzNMv3ayRC76kwrWDP2w4S0+DUNX743HvY
qxpV1glKFf45aT+xChRqMII8PDBPQ/v5fmu7k9Q9G8t65r/DlRCCqZgXIXjZxfq5QT9yGAFGvGtQ
v3XWfpT2lgNArsXxiFZdz4Qr5MXDjVO6aK1/3S2TB4q4baYuuNftlKNPP9HNX5PH5OWqcwnF6s+4
+qztWj3SHAKoQZI3rh/UiPp1Tds3JeAOYKHO4WnnQKVpyfdtilrQJ0xZX7Od9q4jBjzjirBqjCym
9oelk2528oABiwGcNTgKYRUQrm+55RAxX3sWm0YV+56VauvxVCimp2OJx13BphPvUgBZ73qLZsZq
72YGdn24j0sVG7BB0f5Bwa+drjby4OREVi/A3x44DgLlOzLLS0Sw7JZ0+Er+DfaqqY001zZLN1aR
TU1soJFyt9OaTZVjcQIfHYP1doAFUMYUc8hQRRe+rypbJUvQeTu34Qdj8rMSvKOpiqgh8A1MuAih
5/pHnqDRuPqRfZqLxT0M4LXEGm3+SWzP2KsqxiKPwj0xLz1t1/Qn0I6nqQguDAaqKM7XWPZ/kP/t
hLWIhII+jlvuXDGOPm0vutbft/HnM5EpHobPsvXUybK8UUnNfViohoRmdjKL16OUF+tFxPV4G2NN
8mjWXzoSlWZJxo0TOLuaCJOEulOv+rRs33k9yA5f9ZA0+vMfgmMdGlu9o5EHcDibwLgNNMc4CHyy
o7uVOmMR5MMdNUZRGeAOij7RA/oYrwTQTwUq15KXpkdJOu/NUS39RCDJSqNA0VfnzIu4EV2UbQTe
5qRzbzFAbMmuil7pTJbx+qS75walePke/3whOPPOqOrYQ3h+mCCQWA5jfAI4kVkqLt3z4AJXvkg8
Qu+C5wubIpx+WLLka3uh/ICD02LpimRgd89+vfABnGuyxQMB/+ppwTHtJZ7GFYCEKPeU3F7vU5E7
KzTF4+T8EmmkOKWyt3vmdQdY5KWJ54N3p9OwG1DfkYYTESv14sPXZcqmX3HwnCBPpAQ6CJ8qGyR1
xlym6sc2b3lThpC9MHrXa2LRmD2Kymicq29JNYpFMOGdvKlrBeh1Gjf6DBkb0g9BzLHZ4jg5eK29
pgXjNTWTJsb5+492RMoWls9ouPCtP7HFE7jWAf5Wfj7FeLWPvAds73XFZJY3aDr2pijEU5T8RMJP
FncrLup2fW6bjfcZ4uhb2VDdw/+UwT9JsHlCLrX9CeTDmg8cRw75qwxoYsJyGvGh7Ta1b+AHfmBO
RQD1NcSQSfQWQH/H9P9I3sAQ7PXJGF3WKUXjJWHQVd3xj+TyXGZxti9bPboObwWL2SQwGm46R/F9
V/+0sgiK3myiWFTK/9Joznl5Eh3mtY8Avg5N1LmhI0Gwv/05tm9YDLEweNGArrNFoKMTP7HwNo/b
sMhB4aXH0RwlRM1X7s0o0uXYtJHYwdq4xrTyX8RbvQpHgRqq4j1nsRNWu3jA/kbAT/0XCGbvp17H
FYhQ0hxS7wVCbsip7wAYuJ6OnavKk7uoPo+OADjovlAow/IHAz4BsjyKm6Nvg6DdyisoS/nv+BS1
B1mbt5PdcJZKZJh/YDdLYK3jXHYzvzDxyxcnRpyWEkyAsTYySHStiUKNfc+39DgxH8vhRfJZtt4t
Ta+ZqIaXpZN9nbk06EzYJ/AlT/0O+6a+XjlTJ9eMa3UgvC1r0i2ddMHQqL7ejROmQgolb0J51DII
aaVfZtQn27aKYi/vKvbbel45GVaPdI2gWY/W0ZHXv4KOXY/IVZJQbtOtlI2DMz42Guanyhfw5U9O
QjVjjazjtBj/LtbHXzcT1iMeCW6RNRo8ChoxfrfZaTg3lPt7GaRcyNXUtgnIeB3qy/nl5Ru+2DgT
mhwydHc61sqf701kSEIdCWAqXxvhsTYNjux3jBQ4L30yYtU80GoRCncteTwVsaiCmFH5n3Y3HkJO
Np9WZNJyCO3I4CnQ1eAMyUwTMoPYcx+gP0axKVU0+lskN8ltqF7ZwD5PBQkSKi1XdVZtnZJd23gq
tInuURFxC+Der8nYJ2KNVEYV/m43naDtpraGjEAztw3MZGxI0A7V0TzmkgU//yXKmETtrIBKB2qQ
qsxfz/zeBMozoqJAZ589Cd3EW2yALg2ynfi8SMibXyKs3hwNbJgGDwspxrTw3zpWbgxloeTrep9U
BD5pq6eh2aDTlPorYJMwJupvgnGafKpQwqqGKVBFZM1L/QRSmVhysdgbQ6Hlwv5gFpBMaeDGufan
yk7TUH1AjpoIdcNNokOaOdWzaPL7AWP9syyIxJ9k34JcRMEP6i2b8AmjEt0NPyNDo9GvgUEnoIQ5
IrG+E9yZyllN2sIGAyxCt2S9bjPoCwiKQkP1g85ZXtOMjsPdpMPUhWRFCWJw1fkXyinu5ADgvbpt
2DqYcB7chKCceeW8f8OpBRcTQvURGdaVetr1ViiDWGJmNUxg9MIKihxIpXe5OTrE04QTi70JNnJN
zoWNo5k1U3aS1z0eW7kwK+8DoxBWuO5AthytqNaky35jAzGEv+EFNJxNdEADDJSfFd7njcsG77TA
ntOuJvu25GpHwiFKpa53sVoIm+/UXbe6Xx4XLXB87jiv/cnCSSyi1w81WMda0pUQRAWtndf/4QJ8
rzt9gcUTPZGndodMwaZlpZOVtPm32wz/md18nDGUus+bYJNEmLb3ZblJKVacSeWYmofgIpQge2aU
FAikk50dTPDo4ETA3U4/mWSr2iubmbMCvA9iq130kvvGdW94oApo4R9j9AUGPffSAsf1fRLbhFq9
Tbjq4LSaMMUU6rx4WKZbp8FAuGeffvKVotxE+vzlO1QbbIffOwvgBTAtsAMxpk6sZa7GChplBo8B
RvrC3WIiCXFEUaDuLg9LJNpS/4NfsfHF+5Ykguek0HTlzsLV/7Vy2vO90PS/T6qEbX3WXbLs9DP+
iCtS4nwj8DVTtoWuUH0/l+ZIa+eNOg6SzP3UoluKqq92T9Ph6MI0K33fmhT4fq86p3CpYzn1QmMb
ca8M09KOf0OysDNkq0IMP5SqnAbIA7S/kjlBOYUO4wJa9OthY7dgThXuvwTFyyyy7dKEgSjpat6J
4vHL+vV+ucWGfEdjvPzTMYZ7T+s5ZabQgWni87UD9q38JWL1/FxrJUGt24EgBzhprfoLQHtsAWzf
K0e+dwalfh9h9OI72WJujphhqgvxLhiEMrZJ4e7fo6mjdSwEcdOd3OAy8fF+4E4WdPKOSPmYeJF9
nAEa+rq8R1c1pOM4SDLl7ReLjjtqY8VakDmnHYB79AwWS+1+XKvMdJ7AnMP9XkuDFNfrkC0mxo35
UCCd3Bb4yuDpUpqg0v2TsSrwZb5PZzN0KgZVmeIhQxozXcSMcElRns1nbWBghf+DLzkaybnI/ZWI
PP2yI9xxQUtfqlQIjqFGTBM3tBrhpIWyA/MECaQSKnSRgLStFTcmUjVN0KVsQJrth7BxgqQnGklO
cVpZz36AmvziWYR5mCjnLaexszSb6vBSTO/Xmb71xEUTqv1ip1Zl6IOtmt+NmBsWebuv896t/0Nt
cglv3pHjL+/VddJmUgnc4qSV/+j/LbuCLnhHwmoVIjZqhyzEhBv29qWt1TQVW+A8sGrN+1eSIVIW
3Qc6eEUKp1u+bUkBa02xVfdDi/+KqsWu2JV+Igt7dQ6edP/6lIVbGPjA+zTbEa62jAC4pHNyR2YT
DXeLQQbyjQvOWxo4DOet5rOlN5lQaZm/Ru3uz5dUuK0KFa6LmDxuCIvZUmOlvDHRlkUOQ9ey9qZ1
gepKDUvjuGhkt5Dzk5wT++BxTh1zDZn640DlWucya7sZjgCgN/opMPk6K4WOfwtRyOW3U7X5jYtb
n1YpPtOYBiDVpJ5dm2oFLfqbGhBk/f9XZoWqqLqAz4f/qYzCq3Nbj0D43mdFHNJa1o2zu8Del86L
jd5VH1H3PEQBxFql5LaRJ7vo4lAmp8NFXShC1l3AjZAnXpGRziii+EksURK3qA4mZKJpYyr6Ebp8
5wOqqii8a5j9oV/KY9B1sh+MM/P4bUdAD+Q2vaD4cQQJUS1BJhGlyofkysxiuGu9NWU+ovIPFke9
hgidSZGk9QVcoA3/YKm2HDZEkXCV5kBoMYQ1o0dvhcsDmixJd4Y6AvRbMh8qqVUaBMFE0F4Tf9QH
FxS56zyC3lLksu1AIf247wMIWd7MsPTRlxDRwk5b6dOU/KhxB3u9qdPAT1f1rVzWvRffm5iJsrUg
LGrIbvbIR07bGrYnhg9FEiwGGfgRQ7FnSLF2adSbWf8R8oSidN5/zHpUgugwyLLD3kkQl9mzFf/A
V9TFi0jsB1ePIYZElnzzb3ikusKxfmH2TfzoMsNXBcwoHBl5LuPNkT7zkBELHPcWm2vOgNAe+Vdv
+M8n4McwbGORozcI0WVH0Rhyc3U8iOHR/cmW/0DufwMEUGXBDUp5E1xFdP7Zhi5bySq6O7/Ch6JA
fkis+yFP9SrWI6+quCEx3iaUoEeJN3KqjxhaHiVpbP7HcrY56B5zzAs95MZuGH+gjyvq5sA50S6I
fGuOyUPa25i4twpo1+X/v59K80IHJR1NhbuaJRL6aeziU6oMUeWVPhBz6ghUPwXOfSHWU3bdimvV
HRdIhTgDYwUab5jCJYIa6BeXMP9tMqIPGkAQHYULNmJREn1oW/+x3/L50sA1BTbmM/h+XfRg/rmH
iPXZUI6dBGv+yA9lUGzUPQKRVD+Tom1J1kMPsDYIR7QuyoWrE67U5+ams43WoeMZHjbA/j10dRdi
08jAPZ/qsoblaGDtXNxVxnXqLSs7sdyEfrYeVuhqNAkvvVq5Md555BsceeQD/JGTFg4GPKqDi2ff
JShbxPgij899S9f2TJHXNDGBpKKywLDTXA3aojs1iAvHupSsU8y3TPMKwcCm12ijD2Hx2ETC1BjC
NY/qtIvWF3yR0eXSwJLdeYNmQ127JwF9RAj8PZYXMoSDUct73NKV40mSfMxEMS0/tbPrV6yiL5tN
PF6Le/LWC5Bk3H2olqFhPgtc+XW5ukDMR/A4mDKNNVHwbgWxRCkoIjqFWueN76z8XggkWBnZ0GM7
bddQZCNaEr3aMgWnTunvcsNm8z0CWgbiu0eyOE8HzxehYgxCPYI5m/tNokf/mVCWVg/4J2mAXq+X
mOnhBi7QWtBgbXcGCb7K50/K7UYecBKkd9DKvYYw3akK60MVB8o76bYW/Odx5GLCSyz3/3S3QC6k
AH8AXz3/UQRhPzFKKf0nu95rmSzTKEGG2J74yNORZ8DLUyACyFhUUdQYnURr7dGKz0+sHCZdETq4
h7k8sjqGfkHwTRsEDpkLka8QqlNmvnfoKQuwK9leArV+V/dI4B9qeOsTwtNLQGPKyyKkZc3pt8DD
3uhcEE3WMtN1W4AKbgFm6RIWfl/vRapLEFoPffCg445KAfQosuPJ47I/z+Fvvvs8ugCZ5kd/QEeY
fx6sql8KHD/uCd5M2+3sV7rugLr6WVL6wYX7Lgwno6MMLLAKs0utMeKVasmowCiJYL6vHpIdbA7P
QQHr3inNYupnj1L6h6rBU7MqolRLVtj8ow8rBXlkLe/AI9vbRFVcu5UbFjS5AGWLz+/m/+2ao9Q2
97ld1w7fWNFMkfnkYW77Gaizg3B8vbQUD2hocWTHqkbTaZQZiO/hJGV5IL3Vx0nRnr+DofwdAzco
zjVnJ83cS/MWq1eyAH2oZcjQh+1piooPqdUyTQqZkk7SUSgYztUJlFDmsJm+r4dJPT7ImpaOOzfx
eKmdzCBTqyLBykdkRGgoEABmMgKdIyZRCCO7GjN/a8MMlHLkY42pO7H9rVu1yfx4HDY49DJhRJqJ
lwHjcareM86rctKGsdy9dD26rW6oCmCYZM/nJ9rno/sI2ICrx0iGwrHADqRWDldHB5fGvOrptuIo
F41863pHmxfmuXnsY6PpLqY4FwAVsCPU4vgufVuUbS13wf401hxsM/dIJv7AjoaNSmjn+a+6ArN8
0qLOgsgf4Kt4/j9HrnKVWUd5mjAGySvJGetaoUNqcwoWWwfU32AOfbqBR9DISb+cVC2QKmenYjr/
kDrij5ZVzziBBQIx1fL8aFfF6hYBhxs85Hlwfj8FgpAs60gF6xbmvLUW0NQgGTNcC4w+3EOdL/mq
Bk8Gh65iDjj0+MZsFkpC9jireZ294i7Q99WZvCZ8JybpzGaCHZvxjL9zstX/4Jnr2bRcyGxncUEP
LmtZsM9jWOFjbMqJ/LU4uLzMvTiIgf6iMKQDebR2G6xfTmf9TGdpJ94h0+sR7auTdDJB8etXlGy/
DSBZh9wLCtumHF9EHj/if99CL5toIBLr8E24HyASMgSpEy1YQUK7fh9iGYf8WU96KH7gXdShr4Sx
7dzWitMzbE1TgIxt3oGZZCBqh8nK4tBgbOh3R7hP7CSKd4L04nbw9n83Tuz6CnEglOf8rxvBbKDZ
RGADUumhpR//quPn/vJaZS92WBFMUIpBRBN9yA5nKue2qXyScf4uwx9A/bL/PQD0EoNl/TDT7Tcx
Fd5QvLCEYgLO4eVhZmuJ60n7pIzsVH7HWlvMgtlS1PMOcE/fEZLa7I8joL8PZ3LSVLuIuw6Zm8ji
qMswls131zLXgQi2XD+i97dhXrphdRrYd8gXGTJn1yMmFQgS2sqzZEb08EadB88dcSzDqz3KIuBh
tCeI+SqDQ6RjrDBFYlDYGZmC30+zDPBEL4+h/hP0vO7sCrr9EFkk4IvRpDCgUCjV1BRNU9hD4Xua
LxRCfOAz6YZIQphbBFXLcLT/gAFmqWrxgCkRUpEQcKbL/mAdR9myvQxnkPaJNKMN9eqpoBwSvHeC
2u7GZfXBlDi4wIxtxqWCLqcOnRgWRQ/6VrfrQxWufRoarbD8OpuT4n1PmIcqYcWgWq+KNcsRkMki
EKtjM4KolZWlxpm3hh2/nr7TBzOuak/S/r6qw/abwUisA//vrpO3Imj14CKTbaEbGR5J9OCWknA9
kPA1B3GVUH2RIXhh7N4QToy8ncDMuz0/wfaIHMDrpoD+RUoe4PkDsdiPF9ioriE+J29I/AqwZeoG
A37uXZUyTs4cjQToO0QnlvDYf8QhJ9+mnWkFvwfJAnKkpQrc430xEymum10cmCXNxCETAcCIq3gK
FVt4CFeNx4Cp2XCRrwjmYZuSjXr1fPFGIJBQh8dizrL5aw2obQdmCd77tZG+UVLTSlvQqtpktGFz
7P5o83bElQT46VksHHffWPIMk/LAgjkEWhsauZLsUwdv4MNdzeTk7YDZNTem0MsFgmeeoy+SO8bl
Y91l6D04cgQyRa/3qTmktMURDf9CoY6/3o8acvPSHEeVRC9kmjiiuwfue2h0VxlOOWl6O2pYDbOL
RRRdTdhRolbmgkfo/09p1/h7scUZVpuJmLdRN2b+j9rbyYtjNScrlhdg9vAOH5tvnNubqnlhLMaJ
Clsy1oRpZdICU8ZeQEoJytuExvA+0MTZQEYl4g0sfvZsIoH7k5+ZTUFlsPt5b0swctSVEcUxrJtJ
UDJprW9KrVacuTrZ6kp8kmf0Zd6JTKtP+MpkXNwLLYdDbuuh2V6ZCxKQ8EA62SH+oKr384eQVl5m
2vZsxhOdL6eQfEEduECOdbPNe59X+xLNVc75KEOUjSon+pIfZT9m0BDZctvP6FUzjLrESovtMmwQ
7sm6qQOJ8t0lerddGxp7i2Cb5dmy/SjqNdEAKhPIASzXzMUyH47oN4oZHkF/UNRtAwJi3GDsMsdO
I76RbYYFAm4lBEvjKJiReRNC13ibNiB2MS6i8pjVL9vUgT7xIs/iiZGkoP9MC2xsi2LLh4Klgj+h
rKmNQ3BpCeiCGYYA34rNYtiU5RoeBzrOAawEGHpAPuflJkHD/HL5298J3fHiZgJEysZmDgozHpwO
1SEH1tKepmeLBYEv3eNz5u7+rvQRHGxlUPcwqWd43QxUx5Yl+cbhx7FyPYE3Cs1C3ArIWLIMGEWz
o3BiLlXw66+BwXMJzFDZTiYUz+c9iafajBel1PUWD1E2+XBRWl7CMiTQT8XmW5bCBx4j4OtUzaqM
TXCWxvnbJtQzWYmeEu/UMtjFskEfMRp0j4BN1iHtxDTv9pUGm9qzBvp3eRCWblmFUDN0URQ38HKF
36SoKiY68s5buyXjGLF/SG6gz+uo9J8VRCO93p9aXq941JE3OEcttx7ceZxC7ofd0xezS8Dq5D/V
ctytZgc/yMa0Ujg+2aJqfXtBCIVLTAPHzAmqS3K3E3TN7oexPhiH0p2up87PoFlyeQpgi6gp80a7
TxcOD0nRHAKGEnF2mYDFOQt5H54PrVnLDZ882iERWRD9noP77BmMHL0odnH995z0WYEtEcjbKZNL
YV/iSl+yXXyVq2cCfbF1vRNdcPVEqb8RAAWjTkH/ApjZPGZfmZu5l//znaJhVSIPJokpgR+EpWW0
jZw1f/E2ZoQ3OFfE+aRzwI4+nTVQBKXTTW+p4Gpfe2MXHECvqf9h75AZoT5SMhMdHdE8DCxj8ZPC
yps1mJXJF8+G2oejxNzOLjJJuMCs5Eu4k8V7yI4DNJWR9hTHTi6eRuTIg5MlH8Arw9+VjK79tbSg
Haz3Dut+5DnHwJ9PRk92oeQUcZ3sqsPWNX64WLzhRqzxhuvqYU4daykUB7WdItool82JNVqVDU4f
tlEwwieqbQ7T7xEFbEc0X5DWnxlcyJNlAa1uKQFGpH29RHwB6tRSWWbNWqcDxxJkokJjMu+ounsg
R8PSa38tW6jDpwbe6jsMZPn4DUUeNlh/uM+mo3byvhTCom35LEWgOsfCCkgBC9Oo85qR3Uy6kDhG
j08kxoUNKCZrjQNKJEIJIQrW6UI2tTCTMg7TOQR47OPyrBbbOWs0hzFMNHzZ4DXcll/ffINwAkdT
BKm1QtkPfDwy7Ufgo1XMbHexu+X9ueWQ8bUd7UekbXxZZzQSXg2E7AkIgW1luA31fEJwqkaw87H5
2DFo3sevjJ504DAXDDQ2lIs+0HDx3/XHA151GOfFbliQH9dNAtvR8xPRQEI8C0yVagFMF1eYLI8v
HIdl0JvJillgw6L5gMIJHz7om5DH0ojxnsC2ggr1C2ws7M5GT+gZeA4JEb8Z2FnkXZmsi0Kf0i7M
WCis/WzQcylnKUcLmUHa6x8FRNudQhKxlxbbObeClKNG8YxWeBIR/V8OmzpLDR8Ffrtf4h7KZqN9
g1rqzJnfEApdhne2edq/T0SE8QppQArzdGU3WJa8e8R2B1Q7JhvSL/5apbeadK9khF7Sa59II01w
/MI9gvr/pdXRJBLTNVt51FcQtP43joFs5DybO92/eTre5fLY1me0gcQOjGkfp2fa2RLgXPDc0cAe
tUYfq03eWx2EwsWc5KUGx1AREPhyr46ZEBgcpuMstFDzrESt2IznPk0kXS3FNO2sTAU3GrKuaOkN
KqFkYc5vlPrH/vrRm2tXkf8Gc5Mto3jBcLjC8TanT7FzeHtY2n1kgnDQJhwFjwB9k2wwMXmzCKNX
iKlIaHtnjQ+HHy78lEHjprLr6RegmHKh9CAGealUXYkfSYkmPCWLl5fj6ZpUVyeFOn0yDerlEDOM
CjMgnwyI6xVrLlTM6yb9XpvNQUHT2Oz8rp8OtpghrvTYCXetuhfzabvAPTs09lQ13eH1NatMvs1v
L5x3kZVIOviA8QODDXvy3E6Y8eaP8LaODoUB3Lup2K1HDDOiOZY2g3/yM5nbQbIHJMlO4uLBkgje
osChurrU9x96MTCQUwTQc9fSDEjcfhYBP4O9c0BljjenIUkq39YaXA00DLg264LQb6lly2EV3VL+
VuAPK+oPlupTSS4rI88mEEU2JQFSO7KzZ9qek8hfe0aasrVgrlDLdQC6Ila0ezaUAXSA2qaBBgkl
rp3g4oE16qgbCM7Dk6iWjCMNJW0ZqsFSDAPz6oPV19osOsD/3fRV+ggxxq0iRgnqJ5cjpUku5Ku7
5N1rMg1RSKPMpC2l4WH+qZsmJppi+3FVl5PvtiNFJYooBVy+MRIqWgnwBC0lUz+xf61BTShRUt+E
JEfEwGbxCYTzbcHEoUxCoayiV+QWzV0la1mBXBVm7uun/ql+0HUz5MetIa7bGgXyzdNj1uzjRsxX
6T3yDYEst/UX5mEvjsrF13cmwludhX6Bd1otAS66Lnc/V+Soujb1ZlLbmJ0P7BHSMO7TDoQTz12c
P5icwv+Fjfg2RjWHXjEuXCIX98AsMlZHsg8aNT+BOBhN8ddBxr42BolpjqWCWH/ttJbHqaYUMThO
9vAS3zT9eTHN3N1d37enV+5gtBY4GDigDXREgSzhZC1GWiWfPTj4FqX3RvD2g0mGFT7AZlOeEbH0
ESL8GVNn04Zs680dh1qtt4SpPtuWfoVk66WihHK1PMHYPw9JU9iCZMO55g+udVFwnapc2ZhD7vm8
9N+I1PXsfXyObi0oeEKwKxaXAuGFopcnHYZ6YEyn6f/++xTQkVXWyt5DYHK7bqEnaMx1lGjobCdS
RP9XSd20gP2eYUj39y188Or774ilGwhWEmQ3GE36Tz2ce4YRcf+SDZldcrk+hagwyRlH7CVnagYp
CQfCymsCqmxTLmvkW9Z8CSbKc38Eg3rkjD00r/rZLDroUJTWa8aohWCD7GOpRxM4r8g4DxKTBMQV
317NsvX4Ksn5l+NkPtfBudWKTVDaXMfJ+TFGsDl3VOPN9YFHuWLfQ98dPOYATL+2WMK9WDv4jNVE
lD8wNkw3VLbbo7OZtsROrNsY8rjr+W56QmEuXwK4TdCDv3pNGdUhWxOeSy/H9R7Kc4dp8IbocLes
gbUnGOiE7v1Psu4QzKngeKhOBQKfAmgZWVV1EnPi7x/XnV6kp5kS8U1uefMLAFx3Hb1jBCGDApHi
bH+WlJWzqUG2vD7QlBqBRIURNYYRBPiJkW+uzC4X+9hf8DGLXStT6kgunkpE10YmomkPbV5e8hcw
l3f86u36wVXWe/jf/qITzFERVjM+A8dBvSn2L7cxCesd0PS6CVqZe+OxUc1jja4KSvPdcqr87x+5
hDLm5fhELZ59VHjFp1oujd3uj6aJBW9OESx35zhKSklihhSJ5o7AshNvkEAOtSvz+Zno55JeuDXY
dKi6rGQVBZuJQI2zn3kVNvacnpB7htUGoiyXD0TCze102934O6O9hJ2pf6p2DyqlGJCqyZbqHutc
BrO0r+Z88iVn8OK3yJNvXN/3QBuxBAUPNbuS4X/60UmlmLKQ5rgZFaV90jUluy/K2tpoP91T1KXY
kxtlQ0kZGMW0Ep3zV0TdmOHY9Ok8T4tbcFM333ofBUShuCku5jlNf4cSRXWPQWB/6E1WKCnND27b
u2/0BmYn1PBILE86Zac4oU9j2gbw87DCaRk2Dk9xeaGwxU973M/VpOEWtZXgy7bYZ1Mf02Knvdpx
C81mrOgN8p3kbEHbnkrXmdGaD1zbPhJ4rtkeNVgRtcWQNfwsoFZAxv1LiG8Cfy3oQogK1p7gaW+M
buLOk63wqovRk21lPO/dvUs+jDXHtQISKRZqm4xzAJsa4f54vjJdVD6L4bynkqXrbfTytYja+mEb
AkfKHqOV40KHWXomV4l6N3KWvKpkXsXRj4NnBM0eOTqhd0ef9c4lrsXvxdUdY60kRgLI5/YSracc
+7XpZWEQJYFAqHiAYAttxwoJp2MLQYQhVgMovaG9f+3XYSy0Ri1+YqOSkZNVj3R9Jpt+5pBq4jgd
yuxqF/nsiVmrgsPzKJyEy18NVmJ6wbp/oY6Hg1HW2yMfPap9hA5IjKntE8KwmG8d6oYYFwhAgsbV
7PezZ6W8G5sHN9k4RmehMrvGvgGOi6gIkIKne28LHwIwcNjL2Fnl9kC2sVqQT0cWrQf4F4hV7bsv
YRQzhrIyzsMPnrpZS/iOQYpy+nnjmO1+ym+OG96Tnz20kxYJ9nrWIm1UvKXPc9DEKIS/xJmUFo72
B4I/chTXErsEZu1tlP0cvfLWzzIidVyIQ1BiU6zjju42G+ks6+VUJgBx5uJvMUM68Zhq61xu8dUi
HGv5kb6sP+p0rQt6k80PZ2jtxhz/UqSdN/abz+whpCXccTMOQlEC5/2PaMzZKnNkkxjkEDmh1p5F
5IVdni+MgsVEotdNhbKuJiN53/HRh/UkHfURcQ9CDsH1CvgGG+DJ+3uhUnblDyrya4kS3WjJoxWQ
qjzYCq45t0P2o9P1uRTFcC4vpc2r3DRvDmMPfjwSz7gWy4I30xRg+9vKKXrDa5fPUxdVK6LP/Vki
3Bhb3nAz/Hk9S1ttwO++CFMiWfU9NE6Ss0+ZPaOc8dL0ArRUpZeHlZ3eTQ3Y9CfNN6AIOWbzVjGB
ew2lfZhmtfBE9Mmlj8Di8JgJ4fFHsSXBgx/Fw30VMudnuCYMibL+smmTtueYKISgtztWAt6atss2
hjSk/XlyW/Zgo3z5rIPvjGV2ovlgNOhfTwzG35VvfP6jMS44JZsC68hXeTWlCjdj5K4T6tzL/E0I
UnEbOxiC3GDhnEfrri0eAa1h77ONza98V+OwUal0Qd/FfdquHaFIqkg9hYeEleU2DHWMNFzqpKEL
ZR5C0fLf7+IWSM7alDO5AFXRLvflNWfPPK7P7qrcIWujVSBLbA6UxZSZGEzJvNmqYPhEAA5MbNun
HVRi6pFODXJvEjzyzQhp+HacjOBUR0K+tdFNFPEujnEo3PV6AE8JqWbypmhWxJ/ca9/tmM4OLydg
D+67ZwloDS3E09Lpy7h4+9g1PYe8WAe+LoNAJ+q44McLxeiNPBiDfid/O1mOMcYSrWeAjO+kfB2/
KFPeGKJw+wDsJzp8NE6N+S1Cp2VTqn32k6kzo2XFNDyAY+IgbN9k2JMmThJJOiNagbbQoDmJwH90
X2APCeOc1ImxsRVEtmoWBdkaej/ze5BObZF9kemSH4E7FMKjAyzge5RFdNG4rzwgcKGzwwi3RvnW
Ywy88vYBcZvcpYi0dmvGLUbTxWXlyf8nOXe4IEP6YcVqh+d71YJzQ8NRljICzN60whrU3G48sBWO
DFNSGWjJitXffMTB1pw15jfAY+b+6neNNcH3+79ERxJ4o1prH7kaFxro3AyUiI72HayEbWrlXbIc
aZ1kJX81H9slU2FNGGEOxZfkuiVtvpZ40jZdlJM/atsdcWo7bPFTHIlSoGNeaVBmAHbBigELhjqr
bgzVsC5ZJeb8zMNqFtk1cU2MB6FE602TTTbg4aYfsIrpWno9D5vcLwETQEtr9NJMoAoclCOIbquq
TuqIRVhpTi80yoNUZAM2SOaXwAnwprs+GcjRAcB0jxAhRp6PRkADq+/AY0sU0uQzH70rWxc6n7I1
oy3Ufq7Qkr3sNahz1BACny5lJ4Aq3kXbxEt2YGJNxZpVHxGLnl2+9r/fPry8XSXLOUxclFFmV+Su
ClfEBKrx13oW/+wOw96ZfSCc+8qsLNKG4jFGWsZTmrxQpUKGX46YphGbDZpd5TeDZU/rme4uOSlS
Fy+5czml2vKHQkybV2HOKnn2IVwICQiR7vnRVBWH3l7bCrLcpaZFZg4FDnuPBKTBGDKt1BHPIp/a
Pbs3RE1IHUrdUgTI4z+HljeWUxVzKUK04PkbF49Z/ALWdN67pB13rbnWz1KXfeIkU9gBYv98wLsz
lyTM9FAGJRaKMJwISWLTlsaVCV9FdzaiZDEVldaX4LlwkHYzZn5qP5cePvH3vPfdVFwgSnMPB41D
F1atjFxebqbX0gy1dpqyuSCCQCtvD8zzVqecv36mZFyGsV2IeSGKoMeecO+DrFrLpJQKH8Bt0Nbs
K/gysztVF8NlYvlFhsGnqXpXGMoaVPkLGOp4LJ5eE1mmFclUSX8IHflmImn5Bhn0Z2twH/psv+9z
6QVDkqFVop3P4Y8g8G7N9qu8ok1t7rGlST7GMrCyNLaw8yp1U6KOqP/qQ0xp3qyi30Mo8rzU8c9S
Z9WQvPha4STDg9VH7lI4Rzwda/EgCDimM2S5DHxcGqnIvTs/7gRPZa6oL3OrxNzlklusWAnsSw04
KV6rXRDPWR9yh3nYhpnPn828y4E5YgdxJCLVqJufVs4MawMuGgXMKdmscjgx0oDUcOgbPc6zyp/s
qWioPiEnqwHaZGoWBRqfXsW/Y6M9vonMX9epAOgzzNeMi850iqjB6sulOAK4c4MQK+2+5DTEM9fg
9PWisYRFvajxFq5CHcDum7QbyI4yDZpO9ilMY5nDMPQdxtI5nIc0RgdGJ48EruAzyfmYAVFUm4mP
z/4SfGmI9liO41/d6bKgxF79CFVa5aCXbaCeyhYI62ZbtPRYZpsQ0EW3/8vk5BxVi9X2KckZXu1K
vdO7B1JZcU5GjgDzgVJpPwLd1rLvm1Aj1I40ht1Bmt6fR9pY7QvckGLRk3yzXEta2j3UE8LV/HJz
135u/T5v0f0kuqeq+nNvdEYyfADfyXiCmYoDQ99BRL3cuiYdVCo3dhCv1Lm+9FCy3nOmN8ufb8NZ
EuKZSSoRkkU9/K9564NsvnQ6yEN4ibDURq315RCc3mPL/NTMfd2DdTttXO+Docmq0KI9XcS5sRTE
7BOn76hQd6FkHgOh8zub+g+iq95gG3eMUt5W0g1c2DmaE7/yrlRzsxpoA+tQ6yFuYz3s48b6azWv
DassG7W2UE1ISLdlf0IWT6FdtmfW1yDRyFn1WmuJPXdlFdxbP43omSMJ2jCRoJrXvLBDdgJmeVS7
g6GCF3F+tggO3J9YmCsMUDgK/2Oh2jc7LtvnZ0CpfWpXuZBTL5W3GJsl5+ovXX8Ra3k5oOt8g9uG
h9UC7bA8Np9hU2bClftC1FY7GHU85V+feM87OEWI4o8CweKBz2gB5S1MOvDCKjajExWwDtZSpjiz
XoYsW/jSWDc/WuWRfNSpLxw2YeTPi0aYgnq21+ukD1zLIUR87bpMFEA0H8tHk7r9ZUrNOOGac95e
mYDxj8M/rOOPKR9YANcZ9GNcHCMELw4xBe9QbSxmHxlfN1nTdMn3NveAu5YBisB8/oDxPTJVy3dB
t1WFS8OnbzpI3qhC/t/FtReY4B9ZU481eWPmaUPMsoW2zLtbRRUS5QahBENzr7Wk0UkFpTjnGNv6
ghAjSect5HOR1Rs1S7npOQcwgA0yuCP6lAIhUDd/gQc7+riap+4HW3xllGksB1RO0iO5GzHw0/wq
ZtvBBK2uUy40IjQp3OwA+OsWIWfHq+0uXdJTPz4H3rIxkD3IYNpAwh6uY2866YVkKLLxW1zXlx/x
A90+0JpvThqoN3EU6u15fAc2uDk5ChSjOckqhSq3LsLfPCVzTjTXaM0/FDakNXXsI3Zr+P9gPhsL
ewJDEbpe+Lf6oRPRxH3xGhDjM6isbd6w9Uh6jhILCMYxRjlwQu9lcDVElHwDfqD/PfA+cOw5xeEr
DRn6RwI84G7XUVVgwjxtY1KxNoTyZ87hJ/KhEX3FyQWaWUCXzbi5SyykV8Ztl7mGMyMpDdZtXBff
GHEGGPKo8Tvzo/5AXNJxcVraUj1yOuAMDdkdctXG6e0h3IrF9Ks4VJGFiQeqeLKfKpJnFiD51wfi
GMmbWpQYKM7cy5MHOYPaMk6z17JqnFS02iwlMwpdfLFO6hIvN87KD0nNTOTMwnUYFinefTSor6Ug
vHuVqO113sqHZyzbnPS4kUqAFOwbEQT75WjI+IzeHT1nbdK+9xGLfyNraFHd+v5NN/g8cYjvu+2Q
/FIP+J8BSeR2pgetkCQ8I7wBJsQiTQj6hz2RsTUiORg7j103tFv16wYR9REdIuD1bCMjhcWzoENM
tHJe9X214sZFn8K7CadI2RQ4i+UG2p1Gn0gXOf9K+O1gSAmwByDmyMgOiFFSpwvcuE8y1J2yI68Z
5nScVT/7QWi2x6c0nNjZFbo9y7UUbpP4N1tXVEnlyNvXhucFOVmTNOLdd/1m9Wk51MMvb3aGfP73
xd029YENVWZHf+Xez4iclAv5tJoc/UvyD8E4sKuP2HkMk19hX2FOUSbuwB4F1dJc0ogJ/0itmbnf
hmSksM0TGXM/CvHW0txl3INbbthnc1j6qzzbksoC4xbwQyV2erdYd2KLUYd14nngi0rhj0k3ViFS
wMS6OBwlBU3UnQCCJmf8l0wAuUrBhke39f0t5FK+WCc3xYHHOgQ+d/2Q462HMRguGbfFu6MzpXyq
EC/6n9qXJx7oOMPs1ZQGCInQHEa/xEi0NTW/MRNvHOq0H3G4kZwytZZNrTEjR6lw956ZGEO22wnj
1wA59PlIAO32aeO2zl02oCVQVEqh0nFxgQ3ODe9qYuDFcphK8ybluhEX5vd/Qck59k596U7gjJpk
BP7Fkql1b5sH8XrfzPWmQhkAojQeQNfS2Dd17dcyRt2kQEYEC0X9+dIvJTg4dXAcvsKY5PifuSLy
nJ7c6KnIgs1WW8N1gx34XQgKzOrMRsaQhsPizYngDMAQBeC+fDeqROQTWjfa6c6JmqUVP6zCsIdH
rWgJ+CLmkZzsgRtumAjfhPdKmdfdYj5dZbNtECOzAFuwS6Qby1RdR44Wx7vSQw+K+h84m/vRrMWq
22+j41upsOQr7cMLtd7L31NFaH6TA5hxc7QWtuwBPUAAgmv79MVwAD84pDR7sbMKnebFSHLzIIm2
tjhSA5xeJXbFt4g/IxUMZJVBfwUS6PYb/VGIcmmboEhM/s8Kkal6zBSNQs9oiKEwDMNqxMrd5qYF
UksUXf6DOeFPgBwQR2E8ELwuIkM6M26tI5IGLjZtnF0vRyjNHGGDK1N+DFpOSZKFrPIaeqj33qvb
x3PCs1YU9j3efJeDV6cdA8zvRFNkLaivWFhaFwZgxUT3035sQozS9sTKFkCnanVWtds67W0CeSJ2
dhhOBYB83p/P+Nqv9ZtjSyn7ES7shSAfSVsx++DNvhjq9aQ9l9d2eQK1VAeTMlofg5ldjfs+Fx8l
PnfKj4e1syw1aceV3FitULcMsN5iFsUlHCw8OR48JTteVF7G4el25SDqaYGrHWGqcqrxl5WrFd+M
ksS4ge0CKjKQ0o1pCMJiusOU5ja06ZgwShUlepJOAzjpWzoDh07guxf6U+y6VVtGIjBU/kl7RMFw
A6qnottb5C0pckaMKCmdLKhfrq5qYVhQaYBjXVrVSxB2yEZ51Oc0yMVVBOgZSCRG8bN1pCI62LtT
7/9fTXelXXgJ44xxHIlg8OA8wlRsczR5J1qM3awMhXqLjmvKaQmekVdU6de39sgSWqKBrkfV4i+D
etCLkZE5T01EXe5w6gfYEwVD2Cr/uZTlvCaWC68vr5VGyXK5AVWb/J9/ieQdsrTJ3qtEnHTHoOTZ
mvHt49nNBdwuha1eKhLJ0DsZq6wZ3pxeOLPNaLPEMrGRpYFk6KoM8czCY+V9hYJyTig9wrgtV63p
sN9hUE23CN3inqrc+qNso75f39yGWgwukIMVi2NZ24nw2zEBbPNqIsKBjLCkpOXFGgVA7Yk7y7ua
HQlE/dMYCjw0wvPg3WJlJ+YxezlB97X8aZfvsr/QmP0+X5FItV9fZdz69UKct5hNWj+aCLSiiMT6
sAKjnZfmh8CN+7N/bXHrcdLPJibQWxUUyB6znWcEvf5OB2TsYu/MIMnqCGP6uidjG6Me5/5MyLQ6
BV5uAvUcCsGoaUdYSIokJZfrWWrA4oGNY7I9snXvZBlxA1/CrPqRHWNN/TAC6HkQy+6F6eQ7oK8O
eYh6Vpb1aizkU1IwFmfjeSP0ZpGIEbYMHLz8GPJGTbmc6bSVeDCMr3qPsHrY6ULJB7byvVW6gefI
l2DTo0Oc+4HVen6ink2WRr411YOC1nw/AJNf+BrldIoK25b53RcIQtVlvCkIpNmUUQaLjB2Ot67X
M31kHxkt0DjwcnboE17cXvrqfutLxCXGbsf3t+zg70HYG6qwm6B9ajAXeyuQ2fPwaEzgeH4ovTt1
ZyEaGFuU6bCB8hvoqMD68LmcGitrTdZvchTG/iRkuB7eKMHA0ZRppWP7q+ihbXWPSHBfb4kOTQ40
abMLhCy/Q5KKyz9YPUfXrOZsG3ib+gQoVpwaO6Uk5zcrmJcd5ipRGm0mGWUdT+M0dhK2NVHrUdbB
HfEv5e1/lXYDC+GPIqEHk8aAzap6gwJ25CiwABSfjROZm87T+t91WbexaheMXYk63T4HJ1ROhbba
29tC2iKhYhETqFUterSmCNq8Ctccc7RaeRiMlNPdzpXUJIsqOx8o7/wMx8PGeec28HaYojmK6b3F
ovcv8S1Cl+W76bTT5n2jz53fsPp6csfISu4g8olaqigRtUJEt3kB23mpTnx5ZDrnMiZ7fohtxG7R
+SU4GL6vP5oPM/CTayXkEcV09LCHX2EUEK6V9sm4Af+Q+bN4d6diCkXaAIn/xW+iysvXcCvq6bF8
OzxriyT+1BoIpj/z95tue4j0+XdPv6LeEvLR0zRT1H7NWJ576pabflPnkwyE+oxq9WQdRVOPdAnq
f0VnlSPDX1jCO2+gnPlu1vISKfhwi6sG8H1Woz9vrzJDmYNpnmKvJOww85Pjkzvo2hT9NHQPiF0/
f397haUFiACMuyLOE2/3JN4GQrGf0n5TEd2fVQyC3oTnXU+aHxdonNMmAD2dm0Iu9QfV8aa0vvAi
R6RMr0NP9t2A9/4u5rWVfVadNaPBP2vfGdWj4BrsHMa4HQkjyAFCzI1ya4q1rjlaN4i1S5WdyRQ2
0kA8HjBSBlj64U9mnge4Vn8AoCqFJaRGLjg7aLG6d7qHOSca67FSxXE5Q5ydPoIAVrfO6WqkmQE2
kqEjsn9SZXoDErIRYfbEnoqqdoSr72hDGuPVR7rKQzzlTABNJn4n2PGKE4Wgm7i3VvdURMI6zr1t
83EA9sE4W1heA2wh8vkD8tL7TIO8n+8wZnBjW4+qR+Nil82hlBDYcgLXxWfyEbBx9CTvw/0eUnpj
OgUhrMMz/FjVLCtQibhK7AVKgr4OasPeiBwXImaOHM3EW1XuOtFkWr1jrNBjCHAa/pXTHfRj0Gaq
jQY0dnX9a9I9kVYDyWi5aHQSTym6poXILElp7Hw35cUyKE3kYdRHkTlNWwXFh1kD4/QE/xD9I43q
TZE4qCOGXUlUlTk+cE9KTan13wskdxRfSNo6vJBBj7xd5vsD9N1evpIVbRrxIuqYzSO0mWhIevCc
l8uxUxoCRSYw4bwTv7ik4uDixAXqVYmhjcw87rANpLaVkQlpTATolb+9QlSTkhK/suVB3L6Sofn/
Gc2Grex6nGZtiO0fQdLsICSYPMQm5G9nND2RT6zBZIu1R2qbEsFBYFZPqocl3+eCpuYjgChsAiWD
TFKUWr6bfYSMBQm2I22kB9enMl2B//R48e6t2tmt/YTYZ8NtgBhgXO/O3Aw7tQhxmLhv6ZvQTwAf
Mxw8h7YcH+JqHACorkrdGmz5whcB3q2spL3j0xo4DhiVHTDfg2HKDrJDcJn/69SiIuaMgKkCwn+g
tKQ940ZL56G//S9RyC7gbpqffaMjRXOH0SFP5CW2nRjqp4kl76pOJy6FnkZagZkWmXeB0K8vyY7v
qrzcwCCP631PaMkUB9PBIt5roAO+mm1CPS0IF3jJYr7yQtlpcESdDp17rGXFKpnHPJHDIF3fGD0t
xiBovuOzCsroid+lzOJdortXlo9IPSY/qvgjVXEu5kaPgiMG0CPQMi/zQbbUqlPhNCHitjnjrwWT
TizZTVAVnPXCiQH49D3ySfEbEG5pForA9IuiCLH1YXNqQwei4cuDfGjyPz1tWt9I70Jc0jvrCFcv
e4eY9EwRAwB12UZIqJlt9PlO/5ZInMEj2+M/7Lv8OaKeL38fIPTpkyeh4DBs8ukIARSumcnT4o/u
WbpeYa9Vv9CFzN1P3K662DBwGcnJYcRFyQ7H89dGpkljbYbLJ60vZy9ihBfHNaY11ySBmdUsZ40F
01z4I1SEABiIom+sabgBpaBPR6COzgJ+ha1CptSLyFKvLvwfyeg3eVBA2O4r8iJzMvdXkq0sxt0p
XEk7eyn9cVR63FTRyzyQTbm7TVM0LlU8E6nErLWgvBlREyxaCROVrBiYRiSOnqOQKey6iq5D8e9R
rqKOQique7VZ5eTn8RTKrtEbMuEfvsgoOcTqOSpM+Jl2C7eYlqbXxeSINzPk+lRhkfcZOCq9Q6ZP
UME3k1FygjK2YGs+Xv6ZjnTVqV1p/VsqZgsfX9Qs3Xn2Tgm+yoihoZN6jcpeTmouS5Sh43tatP8I
wfimKfRCk2U2HYYzMssjkLIudhdDe7+2Hb6Q2BGLz2bcb9ZuiDZQPEJEw012BRpM/sir8Ccus29v
sYIm+KFcGzGj1cZiIjPNafrhZE2fEiI5Um9xTsRjsTeDPzICoo3SqnqxrfnLRBpcnqDxM573cAAg
4PuqXyXZq4aBLhcXjBhL/XCN73ahUJ34/m9rJiN45o3oMspDrykUL430oHbTpjxAqSOl3u9hd9ZH
dVHzHeaPWKALiBEqqFJ4cfQv1nBQu1MP7P9ejB/GjjuGCCXJ2yI1Zj3kSnZsHUPsMB2c5f5FwkKM
w3BWQULobONCNpnaussI6+Y67x54Cq35xuqmLjna0z/qwTi6pPOSGWMLLs1l8hJnyK4+MB2eUpIW
/r3zJwNkfPVA4q7yiRR+Y5bx7i4DRwRQJUxqktgWPtRGGclNuGTLwYCu3/BxkbEeFEGOdh7+zAgs
dmvxS/kWM20javSlzofY1mA1fCm5JemktYpcQ89dLECoYIlwvZRvMz00K+eDeUmnjiLXsbg/q7eo
lMEvcOg2NdC3BNia7+SUEOir0O5U5cHjj0CoJK/eAPVqd3DJX4HNPY36ybEabz5+C/KtoJLaJd+T
G8ghNqcrCnziGEm5/k/1RYsitJz1qRPIYco79bqDoMzufXP/mtbImFCWvxJ5ACciutPqVUCcLNEU
bTF60a2sc7zNVzI/V3L9fYCWUoTCLMAMJhkfRi5JJ2V6ZXe8rWLGqlF0GaHjna7YUjvAgMxy35hY
JLXaCLi3J12Kk2jWiV6/wvK0swufsICrQkuHhKXO8Wd4KIj99KznulR3U6oFwVY8weP0M4sGnpVM
shwPOZVCgueiqXu+sCYHqnHAQZdqtOUR5soWF/X3/JVrIG4GP1dg2TcdBtZSgqb9a5rRsBxsTuMh
EU5B6aq4oJ6qbflOd37qxK6+PjShLbbOff7E2OOdOMc7KJnrt1NfQfoQ+ctRZ95MIquv/5eID0Mp
8KQiAyoarRvHxAM/b2OMd78eBnjY3gPvEgzE7Z/qDtVllYjD/Kt1Z7GgwkIFO7u3tN5PrUs8ZUby
etIaNBz19ADnBySffCcUnzmF4j7OcVIzlttj2wlpLnDzLTuYaX63B9o2MLlCQunIs4BDVnI6ZTjz
xlBeSUuTZbZ6FMR7plssOQk/PUvw0p/EJGnS/A9exfq+7yh4zGNx2KffsD4pbFxbhpB2ZJDukK1f
XTkTIE8JJncVA2dTfUcLmi2p7XaBGl1yz/Hz73GboRglTc92MFNLqzdeG+tltc1vCdtg0jSNzPuc
GQlIB2L0HzlRWB6+Myp8J+WqvlWDNqkaHJXyQoo4mtwrUYuysKjfRnyEDPn8/TdXCYc6SEMz2z2n
8k3WWBJv3Cvxpiu7cFm0zSiwjLdss6UHMP4Q7qL6P8faGG3YhfYNBEjvH0gDusirCswi99HYEU+Y
SWLJPiCfUA73LbDqhwWvReAVc6lV7gGTnHEpw0N6AxL5+HVQ5Z3BCu/C8kKd8LJhq0A4cWyVkou4
D7dNbQgPskzub84PdGHWhMR8TOO4JCbD58ULBPeIKqc/DjQbCs57xGnXQAegJYS91kWDA0M2H05r
rXqKhm5z3RfvKUAPZAfgHUGcFoKZoMATgECZCE96kmIhU7YwPrKo8OvTbEqbV1g3IgOC22y6ToIL
SEtmzaCkNv7sFZTbpZ23dJ8tcCv5hMd1YEvGD2Qo5uUCQLveBl8thfO0Ci8gpGc6WkARi7Hxp4yf
n5mybWsMbNvI+0sdqjZA+PP4IiueIhF2eSzkMtBD9wRCouQyggD5WFk3EOptlkRGlOmfVSb5quPP
TuZc+Cg3dZiMKc/GoR14itO9yj5bmtY/1NaL9aasBBw5kftV4UXrVasNWvoOMV/XxwjLYUN64ZkU
9FkMfugC3fDKkUU1YpYLWDa/wmA47TkiNle2MHgyFc/bEV30cWQ6utc/xdoKcnlG7bNJOqRJN0T4
1TFzRH3yMHBfPAbXoBk7QFTxzmtYDAJKSNEQXbHO72RE+Vazo9M1cUouHeSzIK7ZmAZkbgWMk7xS
4F6k4s4cOwJYFOpfJmsV8w21mh3shOgJ1oAQYxRKifQmBSL875YCdzOcYUYVZdSOWo6juGHWbYGh
VFzsecBnsoOi6BXs7PlurelEo1OqgLwUFDhtnETc5JBAgSPdHZefr2toVM/SOU3yx7yXmq3DJCNY
eDdGNtJZKcg9tS7XIbG0BhwVAc6faeFKopKmlgYH4BhE3GVEYvWFklOJZTzvXhDd8cqbmin2KJqQ
nsJ/4iUkHO9q2lewz0NPF3yavkAo8vQ2+LhYfLJINjVjgRB4JjfOmosF8l635SyXn0dAM5mt3lzn
55y2A1vIu9oHOAcEopt93dLVZaZ3exUbFuMmxarAGBMifJERFI35bz0Jrd6D1mTGki/U0DQPr1AW
KXujif63ddXwy8yE+MZwW0CdrMrU+vGsxhdUzRCSaWtq6TQQhIezJw3MV+E02XqMBvCgRjdXEOP2
o0C68dhywlAQOiPSfR8g4ZaJ0parxdXM7/MulxnWu4FGQcQf6DLjl641qSd9tWepFQrnO766H1qG
kCPdsk6B4L0F1mNdtI0DHLWoZyopTssAXqSpbh8Mx74o0cCJyVaufMXMgyqekt7hsP36jhg6WFuy
jw2OXj66YEnC5ISNGNuyiFeEpxhc3zHmdsIVkYD/vmAJ3ehOHUCqNZ/iMw2KfjpXjSCcFkg64D+m
MJceEuH/zntGGKuKNpc8VegC2Hxs/dMbr+UB8PekQhdrB/rfglaJXUcP4bU2n3cBZ1nO1ArWaEb0
Jyh1v7OgXfohdjSy01ez1L2TeOW3Z7o9cD+JVwa4fRZuOAMxwW63+QRAJ5KL0+N6OcqDigDeqJiM
u0OTcQoPomUU5mIX+DQcr3ziHEycj+O8vPX9Do4LF0MNvacgQzqCB/SaEylZHBINxfTf5nK9q7rd
NkDhjCx1E8nemHZTpRpadkixHboegJ08DedfPc2nNt8U91SUi/QfNB/Rqjx6btbmPpij8/8Bivb4
L4HW4rUjEYJXhQ2oHEPR68gHkXJZjSz1TB+Pu7O37CAkQitV2CVqOft/dgUHzKVhthQPFV93QcaK
yxDuuoPJJEv7hAg41Qf8J3P5tdsdNhkp9H61sc6mo5KpIvMt/tdqBeoGUwdAXSKtBVWt98Oc3eME
LBpUa/Gn9cIDJ1AschgbVWKT6fg0T+z92T4ceDOAYhVrUc/QbNX5ilg+sAg+RkVYlixEU+EI6I9g
S5i153mE311mYzjt49vsp0plDff2Qh5tYtOFifTbzvWtp4dBJK315+ox5J3ROTmOmx8upi1LXALy
tKd7+0jnx+vLQ2yKwKS7guTp3XjC+vn7to97zhlW9IkMokeT6Bt7K9BUNyG7jg6zp8b89qA+NIYm
nvnlbadxIwE+de97D6rUT/+Au8hTeB4/n91NHLmorrIilsSa384y7FiNXSq1lEZFykffbU2eZfrF
sbLCidtcd1GL85FGGrpPHy6znrAAEmM/vQrjVRbRkj7nY6cQjREOotOiCYATGN0M3FHNCGzZdisc
vMCwHKV1FJgopQ/P2rdJS/ELOdFm386zfW5uM6kFVYjdLb+GD2CXTJQJFvXR2dAfaTLzXZd1CAYc
CHZ5qhykRhAyRzt5G1dlUvajOc5fwhRqpvdP8iRb/u5pJnVzL7119oH6lP7DWrEJ4U+YOrHw+dik
hpQCWV6c9rHnQsnBtbu6xbtXegLgf6rYysgnegJbzCdEoygYS1hMB/rQ1JeemqR4GxujMPft5GyD
1lAdkndYWTPxr4cN6gWxVTjq9pA5tkp5KJ1cEnJr4pY2XmlwuCAIiZDqzqoaNlP12Q/rOGFI3fOb
7zRo2VUmSllqn5bUF1lxZ30RDfa04kzpM5KAD65TRihDYmhmUfWx9DiODQ2hQuM83ygDzvXQd0K7
HnxSdkOPQ2w6qvUGij5Vmi96ql5bqCTuF9pvfNcvVaOTbPJVKv95ue+wwuv4XTT5HFylmth6EQz/
6y2lKT0nCXv1SWCEjsj9F6+yTmXWmrygluqDioTaRVXPhJa2STlTl2pmCrQcRtw6M4uW1nPBPfYa
3DNozGqHYCPvHnLp0GBN3PXmRwO8cIcE3H9c5gNJKg2H3pOfhd9PaFE4EKlmU26HnE6gyQHNpeHQ
iHNcbik6jpE4Q2HtbM/ea9vQHI2zo0IMDSmHwUbJaB9hqO+yw3OQy4Zo3D8HZ5zBSypx5ed1UcjC
Hl97uEsgYHnwPnyuOfc9nfud5v+SuGNEcefJl+5sw2YFTovCEwmRAghkh3jYyGKpgPOT7hl2Mn2V
TRXXM1WOAzzukX5TCCHVGRTI5apWSBhhhiZv3Uvzw5sMZSgsh2bYLVABo8YQcSknOTYTMyXMqfuc
W4BmUqHdnAaeXIuHCoErJTwdc4P0V+hsxDc9FuSF6mLKMKnpr/ncS/0ztet5YUm94qe7FZsCrefr
3sA297DYbZlQAjGyq0Xt5tLp1iCHoRK54MPbWnL0PpVcorTJVu1250+xx+2iQTzke1c9+mt2wTGp
Ew9yrut3yXp1aBbgJqBVkEiHlGzDYxWi+m/z7Hgh8hgLqWkkX+1ZH4sC2Z94/aveyWQY1xkQbVb+
kSGf5lyB5vVi2mFShk9Cf0KyuAbvcSykERWyi9E2umIEQebzUPREJFMXgpRmQkBooZCbPLGd3C05
77WuYbnKerN8yYiDumQDJDkjv6NsIkNj67FQAAzQ05cBjldws/2dJXB4Fa9qqFXOcipzqlk6eQDV
iPjvoXezfyKVPGxwhbZQSCOCz2mNrDZmmOdES4ypRk09OddMOpi+Xy+vdAPUhTrurdJWl9lM7loM
4YMO+F4jk3UepPKut5/Mdnr75QcakQbVw+6/CAZwxolHLEXNMYcv8QW/GJ3MVwYRlpxEbOARh63h
ApQPE8/e0vD3rWIVD2lXwNINaUlyB4D253wQfY1+FKNAJCzOfsMDInpoh+Cb8JuwpNXWueutK1ky
12dSUe8UfhKoY2koUM7byk6HwUejb0xSv0Cy0wHMe5QhGlowpizjkzNiyAQBwWgFNG2eJ8f3SFFV
aDhv+GUFTaAd6AqMPW7einDDhYZHdgxEfc9TYeqDtyrH0BJkLc9erzVwxiFE/+0cPjO0W8QbqKho
+WeYwGpIHa/JNJqVeDIV0xI5q3vajBYH1zgQb5Wfh6mez2s6OQWl8d6NEJNmxhx3RSFNEk0wfnvS
iUTG15m1FiMd34GAZ9gdpsXJ6v+9PhHhHIN1KeGYBYBI74o5WenD1LyhlIZRo9ThFkJBW/tCOLWN
pb6wXxzJeyGJ3UxZUmXxSNX6/ZnTpU/hZN6PbZtGs5jR5r5w06ZXpRJKkcJIYVUNm2qa8nn1gLMU
Yt4tUy5NPkzQLG1W3TO0/h13TWz5VPnqZ8anikrXNo5+QTZPLLp0mQyddi9WC15+2XwL2VRcmgJp
pekpJUEO2bFs4wzhtoz7YEfeEaQdWeo0H1XoDp0epfpny1g89JSgEDbq2Da4wPcGnv8E04qygiTX
eigZM8/r4u08rPzrNhA1ZyRs7lZs4PO9U4lFmAtAU21DP+4YIJRx14ZAmA9iR8Cp5QeimReYvTIQ
qbxkVb8gCaPtZqYjAAWcJ/teP3kXrzwMK8v+so+epHaPTZfnUxEErhH4tr3CBWLNUruln77V3Uvv
w8Wf6crIA0TkxRKIzsFMS9S1K3x2vnRRKKH5AcaXp71A9dNA2kbBUAt/hxs2hG82a+3vpQj8Dtis
9j63QoO9yAwAw4izkQYgAqoMA7sz//Jia+gIkTPPY9/r5i4GMaTBEa969ls/csikWjn1ij03Hnc6
qsIjEYtBQ1rJWkjwgyZPkmKMubbIl6WeZsNT7X7xurn8dCMEcpvWQBph9z4yVMLFCmYXmapn7LSN
yzJwMHybznJL9a1ERmas/RyoxSteSLszuT3r/7WXX+JNWLv2POXVEEmwRqSToeyKPDH74bqxlRqg
cPyJCFtSRAcPl3+k8GT0KXb3/1RJ1iRaryafcu0ckUhxm9AQVl9w/gEfvyQNM3uW2y6lsM48JNMa
2FGPhCe4ywM1pi+Ec1IxaIq/9izUMVItNbPAW/hMM0C6yiFr5fSQAgJ6PTAi+i/OxCnmzS8x7dEr
m4hRfixE6bUOp1UfVgpKCShkWXKpmGa9i/jx33+ys4EyAZ3MvGYpvYliJwLUtbRALDz7LbwdG7t7
WeeH95A7KVDi+VIzqAD+oqbi120+xSLbQWllu87oSBWigIa03nmDD3nZbSroAdRy7DrfMX5VUrl4
0NeCLXEWAR0xEiBjNlxUz1LJ+EChYXnoGCKMXThP3UFEZZx2jlEEnCpKoNX3QrNACtm8qYj+8mUH
kao6v9s1VBGicAnjLG5GMfoSsKKsaXTExF7V9DDh55iqFhblh2EVrlEUPsfI3l34kUb7FSfdMGjf
MQR1XNh7rj62+RHljzbyJQHfgArHGrx1muG65gFs5UApZfa5oPOuMoAKv51vdkXPbYi2BCUo98gc
kpz87RWNDi9zvneRsW7IdQz8Q3mNniYt4Uy+a5czaSu5RkD0jSeY+Zq9QK4Ca/OaVa1+gsVADbhG
NbdtmPT9vyZM529v+7057AqWvjfWIAEQgf3Tb3TUdRVRJDJq7gErgqnBSM/vHVUD4nkjZR73WVl6
9cP39a9z0BAjQvAj1x2sHToRpDuNReyTcTO6CUFZk/qv+S6SdU/qMzd9Z9sgl2d1umtTIguhjKhC
IDWrcrtnQc3t5ecnEF87aOu8XRjAFNi321cZP1VQ5jWPPg37+/w9AE43aonGzm5jdo+zqaLUshJt
1Njed37PHz8x+CCaMgtFYUogUwgRCNYR+sfyfqmE2a3WywMnhm1YerTooumhu82qhF2iQCgwnc7j
KiGi+LBqUrm0VJW27+VmWIvDtobyg+sl/k0etZJTq92vt5mpJsh0+LrIV/wirXd3Kzkx9e35yK0B
H5VPYmibm1K3ZBUT4yV/dq2NSLqAOmnSQBiNTJtrYya+CX83E/omP4dmTT7YQkX65Uj9Ag6nHVCM
649Cc12aqNtZthRiSQ1L1FcQnTZ0uCNyB5eL1JG85z59USDk38JAYC6jQ4CauGlcOOGki9zd7ElC
yMJhwDDFXqjd5UqSmalk+zE4vpGst3nq+TcOuZCslVQ1a3igfOvcYJvnYQez6x2hwEfiVna3jUSx
UeBKY02mgTzFt2EzeX5EX0XtTRTsrWNHovftHrjcwIfPsT0fm3OQCMGEq0IIZv5Aswv7BSM9BsvW
9lib5W5y6i1fkHaylzis6bFZB5ChPFPHOXmb0wr8IOuii6BZwxyT2fVmFYzCmHQ+yIfcNhX6X1Bj
zn9uvSuVt9cy+uuljPoLHxCiVxS0M+iZ2kkZR1TKq1PKETyVGQJ80S48Z1f851nx5CGvBpxnVoOP
7mKHEaamcAFfeZycBFWSXAp88S0Nnnwf51TppK2dd7kgIBuEED1NmMeFXfWQk6kLX04aYfh14/2g
Q4cNsxaCNVQdj2njJwkCKGFmtkmGLxeomVRQ3fHZ8xJwSbJ5zFcjxZFilD9qYUf3MD4yZ541sC9D
bil83rSPzXa8d5otQRD+YMm/+XiU5z6/vmd8sMv2XCoSdssFQ55ehozMYtJcNKYpKu8SyCZ2k+T4
p0Xd9f/kIem89uJzgjyWweKAnMBjLgNz+7QMNo/sLPzdPwwi/XKOu2bpJd58ZHIr7Ul+mrRYLiuL
Q0SqtK0nTBfdpF+CCNtSiiGxo4bHlhnNcHEkOIpP2Z2r5PDrIqCSjUQQyCHGNLXSgS3MkHmafmXZ
0SZHV+0hKeiIZMLAUW4QIW0iFkV2rh6u3ESzB9E6MDoCgDcb50KylMM4HCpR0VqW3v5G39IWoHLb
WMZePzyc6SDCglnrJDCxgcUccwZbFtaaSHOXztsEHVGAkHCc0pqKBB1PhuzKumK0/7v2En8Om6w2
DgoeHqvx1BVfsNd883bA/bHto940jA9kPb6ROsm5+C1P6wAh1FkXPY5VDFwKoT5+6CcAEQP8+jel
ssDON3nbX3kznPaze5kgefPVYnluzb0wxSskz7crTQaidLtCXadqeheB9Q0D/b+ODs0L/7QeByDy
CizaSFbVNm1RpBJaP+szDi5xqrsVXtmXfW/Po1M+Yz3kwlXgtSM5y5jiP1+nyy2mjS/zeDtfM2Hn
71ePsI8OeMlPhMxP8vIdyFaA2c+zIsgIIW/rALiepk+ShvMum68k6jPQBeEPitVb6eK3lr+3a48N
BpEpmVJmQDGTRdt8jesym6EN3BCZiFkkmJx9yibXK8c7lZF5GnzCQIvSzaDo8fdYqX91U3bAPgX9
V/Xl1oFJR9IZAfGWTPGtmq9FY7YAnVZhscN6jJudymuZx+R7qeif/V9CuA4KmEl/0dYjimFj01rW
zZQ14EdW8S/eiAR6LK9jP7wWWrARQ0CfwaNR2ICs/ubMDvI1LceFZu03r5+KKUPM6/cQg8xltnnw
sxiaZE+NmZPYdQ/vmaGOzRUJUZR/7kD6CFPJ/YPQJj5UjSLTbPPlYN8NKZCTx2CYmedudqZXlCOz
sgZoQnFytGeWfL/2PjpEQQH8aAh2NcvUB4o/Lj5YqyY1tBkqGaKHCVz6tEozyhutLKXkPhQ43Tke
5tiIDtCInD2o28BxnTyigR/7qBwa+tl8XkrZPBW3JVvPwOq2eWJpxjlA0lqTyu4BJ5mrlPUE0RDZ
ak765Iz0JaBeXaGp1TNWUaD4PmgWOY56mV2m0gzjFXsz+XjYMS2/9QmXkL/sI4/kQF1wjMV4GWbe
ZTXXDyqPn6g+/6vycEF+icxn2fsqLWEpR7bKHoTlwC5oWX3BcruTM8ol12qhTaefLC/+2t70Cnjt
nrbQ8YD+6Fg2SayZEDure/zrB3hA75F3d7MzVm6E/UUnZZIbSdkfSpIhQujrg8OIfSzVY2+IODu/
qhJsIZRVTLUTW89DPtnRy5iG761lJz/BPnaqk39R+6KtEHbTZ+OMmWYAmP8FGEBF33L9NtHwBv7F
xtfMt6vtTeH+K3LpPsSElodCgNxi1sWnDGMI0O5nRdIe0nb4z/R/8axBFDj6ko/psvnHd+OVDFVL
Dkz/H0G+dXkXu7kmNOWkBPidhElhzHawRWnSlgUb1yvMqYYa1R8jawWqNsgEcdlvDuLZFbpPPzbT
F1IisbD06pG1ghXbNHvLfV1Hj/3Wtil60XtVwpT08MhrTlXF4PV3FEU4qL0lPni44clX8QxQ456Q
zyZGRhKWVsXn94V4ZYRRrizEW/cEORWXdsqd+GZsXDHwFyz+LSrJz/9bM7qlK23PLGOlvHGvHWgs
DR2WkW3S0jmYZ5ZYjBsIDYUTW6XkAN3EEpYkuF61g6lzUGUA4DLv+9H4KnEMm2HWhmPX460ud6jv
MKrPIeKAdUf77gAc97WqvTzOZM+YYvWsVZu+YUxJy2MT+7g9eEnU/MzJvWE/QaMu/Se2IAGtgjDf
54gihbnWpEDdm9wmFsdyW0XXVaVX0k8KSm/t1KZht/gphdaqtYpd7BySRHnx5v87B5AYY2wKteab
N85e6sUnisj00uz6wciBSG8UasTmXmvACIeldRhTcaPCG/ERSFlLsqalG1V4hL4k7En1b3xQ/oSi
jaeH330KsKtaJNXg6o7AXGM/RJ/Pf1HFTy10M62wu6PKXCOkkj3VJ8f8PnGM4GfwRc5Bhq0xO1eL
GW/rK5bB7oXPHGi939Ca0PghFzEnwTO0T8GLmKF+u9na3OtGfXgj3kEpM3UXyXDhs5UhqqGECkxs
dFAaVGtnXNl+56LW6mp8Y7YtNJ3vv9K6lvo7Af2VLjEHGx3iDwxb3YiV+TPbaFuyGDPKYLJpsczE
4iQtZCkZWSeGoZnIXymxsE7SThYNBhZ/ZCO64f6EGm9pYeyM2U4NuzMLM8XZlF6lC5KRXeGo9f4H
jFMWFfV/w1wKef8yvY7O2s86K8UGt2g9vDEzEnpMS3KdYgBnrtX6Y4JOgpEzYR1Dttno6cZzeYnr
QDS1aQv0bGWZExLDvxxJVtsorzY4upJY2t0RTjxdTx5KH19M/zWvFcaFU1Gbxs4nVlEG3qo2Xj2A
iFbjrzlUOCt1eDb6/VpYHaokTqiVIwHKqLNNIri+3RJzwQPtsRnq+AgwvrpyOp5xr70vHLmve/Sg
Of1TRGT6RM5GyAgffjSqAOd/3oRz7kJOZoM/cNoF9kVqfddWm4tyuVCiLGSWuaEKZ+zGeT6MTa0I
4/1pYzk3M9IikQdoo7gqEzPJ8VABOSlf0TvZKZqarcVUB+ZRALKtZBhuj1e+f0Ev2t5Y95AVOW7V
9xzIZJXeWxPyw8bQDrArfk3Rk/39uQmcglXH/i0mgGYwy95rnZvW+uM9QltEqZVBCvVZ3DXQpRfG
aatcJgQdKDAHsLMSZuz5JT4+SptQwIv3XyVNn/iuMWTNesl3/BB4U+CFB5RMQueBG3s/VgP2tJ44
o5ZMn6POvGM3exgMHO/uX5SOq1RAZ3Wx6RqrefVLL5bt+R7O8U/luQDY3dWy4UOgyqYNt30/RnVH
NIBfabd3NPCvdyJviD2tlnklvKYPGprqFkc5p8OMpLsATI6amfhcAK53kgrcm/YYF4aqreB8Ccb5
PcwVumpKxaFeB5NFEnF+JhcQ+KM2/zwpEunHgWTOQmG3SxPYdAJgSsqYGnLSkganaNF4QkxXJqF2
QDv5LDDS9UBWNnAGwGHyc9KdeXk8K8lebwhN6LbzSi7TVRqK3lWOL2xbw+7vGTIimk/6BLk1A22Y
MdPsCJA1+A1U2DQMHtId4k0P3xDRwm67YoTRhXQ2qXlDPpKS4TBWogJq4TEJHs1211BZ+KEQBU+d
1CRngF2a4Q0Vy3ejHUMrIsOpSejZ0ZW9Y/IwIM/dalhf6knTX1/u7eixvto3wQOpQtzn2Tgy3M+v
pBSlPTTAzGxPjNtdF/LufxJLyS7WSyHAOCKEfZiDtMwgmEtNXq8iWU6YERt2H0ekNycFn06FRcfD
mKgXjn1g9MgZqTRbl90Z/pKR0kb+8yYGdz2+pA6BPK/QU2mZmSULkxA7ST+WsHDLuOoV/nKrAScC
/SC2O5bKgHOIcUCgnMP469RemSSwnVCrYdhtSnX1uwvpSFSYxgamQCdpxVjdBmlsc2qjPXL7vSnU
3Vd/tngB5vpBfFA+wLfGYsxQqtHsGvyPGLZZpiR8/2zB0MlHoJGg3iLpainjXNmpfDZqziRYqi+z
W29W6NMcXNaMl3SNj0wNln/zVTXMQBgwz7GYc+PYaS0tbDaTJdJoEiiww2t/gn8AFNQSYT5fE4wl
6zCy+hyhMjcNIaNEGYFh1qJprGpfZu3/8FMmal/rdGHqXT9odOx3wabQIV3kvA6S+Khs95gIBwNI
pYjhGzSqCPRpr41Hpt2gMLAZKF+gDFETp9LuEAKB5JTYAE5geOVTJoCnjbHXDPzGpYQjFT1M4RQl
0pHKxgxgSQpzZUNaX/y7O266/8Bh4dQDP5B74nLr4H2BvS69+1UzywXrsyyTirY5XuFPjF+eiEkA
EUudj3fIXXQgGLBAfng8oyT4yR2CpK0KhQVWEWMBjZhVAc1NBGrxCGnmN+8fzpwdetlThhDFIo97
TpRrVF9HvJlSAIa0KdMN7v/h4DQZBbPRCIcpj4+bCEM4NxrDXDCtj5y3bcDIUksC5qnblxjSrvfQ
tM+hImO7nBJ9LYWCOgFaceXJXthE8ypRAeFhX0+x8spoqfAVUFLsT4Az2wpkaftThlctK9c2S+p+
Hds4buOp0hdOCZy7CWFNCqZlLDx/1igg+DW56AvLRC3rGANI8r1ekqWBOGw40XhQVreEPGhrpf2v
i5lGZSJVVSBmRAu0gxXG4TeQTS2X8FyzejacufJKgwmg+QbL/o3PROUPCofzoF1r8rEesYzNjvmY
ynpOd37apxp3IfBz5UYwNSWmggRQwP9PnF9joYcUZ3pG7B4va/gbirCf7qR26Z7cJXu3dFwQOStP
A+HR9iCXFDZU4jQXt4y87vW39zbijTqBY6VWSqCF5feZTNao9U4WRcTUO5YjvlqrIAnCyg/YpkJ5
PtOJsUOsJAyVlyHD/AvEtUzo43OLfmmQK7XocomttICyNiibexexgO5xjHZ8QdrYJRAyNIW+y69i
cv+5Na3bSH7Dl8Kr5u56OsHfgh1CeO/7zyeSZQjOoILF4Zz9iD+/5oDaupMxHYC+nNwlNSxIic3j
xxPQfUqNwjHTDxPIFCHqQycTcP6jSpVc/vvmghAkngVoiK2hV4YGiFI1CXmR6hIcuDHORPhtKm0c
WdyGpqLg0NQI0wiWwXHKuwYkCvT8WdKJtYIQRrRiQ7P89dwtmQ5AkDiXr+9znBfyAXnVJqeYIfCj
jAkUXLK4e4MzJkFApdIxZMfl+kAV3Izm8As9/HcBfwGY5zWycaKDPqzW3eC6x1xdnxetEk3xaY7p
bAXH8aogYwyY05E9fSIVNoMv+xjV+dyoJVZ9/Xfr/k9A43Ca+V8fIztapsrwFY24aGszsvZAC8TK
jCB/Qq3IR17AtIJkGM1k8hqJB0ZyyjLQrRssT7jnZK1Mnay+jYdFkYmnjrNjtgcS+ba36q1pb230
0BRIeaxQGS5J2bD5ubgZnLSoUagUKofRYvopOoD4GPlVZnUR2mjftoggw2B8qO+81Sqh1sA09OaG
MW8lrbdsTYccw6H+ShLBxgCt1LMTdypynBrK/ddzzTY7XLf8/TVBdi5s/BcXjyiWuLoqrWBet9+e
yt3G7p10zpYDneNS5faQMzH6wKMlBYhVqPU7NTchHfrMNTjulcNv0dzBTGuUCex5uZjQLUMw2pMC
lDWU7fU4M/BhYieC/czrSlIMvjHFe5TQXtS5YrnypKHV/WIK1n6zsPrEhrSdtuO0AqSbQ85XVmQB
+B68yK4IP7vmlTKob+kLjukEUnMmfPXZ+lHQT1BxUF7Q/hpSPFiChqF/kAG6XThPW5v8HaFbfr8o
K8tMvqZDIRaNrM8anWRNhIIfcOE7GL8MfE13VALwTKJYA2bynGkiKg+8KMU5il0r8k3qRwIvu+N9
MzedWyTF/H+iYf7RpilBESlApBM93Wkw+N7PmvZAMutY8PGf2o0jgr6Mom9tNn+Sfwh5Uaxccxko
U8DJCYjim43EgdMp1uei+VON4Y03gZGDvYsx24w/85GYjIXovs151OqFRRIGv/OzAjzShXL3bY0N
uc7oRVO6niKNlqxHOj6euZvqO33Bzkbxns3d3fkRNCAlN7tgso/C7xwGFmhuNV12ZOk25gSHCz/Z
iOBnTuHyVO/GxI5eydSl5jouwMyHLe3VWPcQyw0vfwfZGfL/POgdnUMcHQ2XdT5dipdNJdOR9YPw
5cRUTDGc0YcA9SWrpjVmfWH41UNG5DYCwDLTaeqEE9KG/nRjUZj33NiAvxAmmEvBwzqHKv8zf4mJ
ln5tLds9vKdn52Cxj9xWVdJ429josZJyFE5b/Y/l8uXSnbdNgZUdmXUrta+T0AUgwWghEuSrdFSQ
3LIZyk7/RIJi4rfrY+YL5XXflxHTNzVDNJQnMyNAk96GELzKM9HJPX5N5LLqyNU8ROIzIQI/jEjC
6lkyYmoOq0XQaLTnylnHpSACzGYBJY7G4gSQeUsNvrLRnU68xfidTqjw7TCyqZLp7nug+e0kZmJw
eJrRDBkvOTyL9Ll7wpmldLpZqujbWQjQoUIdOr36fQy1u6Ec8xwiX22cPcvOwJsO/YoLQ4VqD0Sl
xOcvlfKPd9YaZ2GVCoY5znV+HARySVdwDcFQ9MijO1ZzvoPfvk1Qd0UqVOpmlAViCmwygZ1uMyuY
zE6ZOKQ0XD7rVd7/JAKbL5EEKFVwK6+XpDRPIL4Oe/JmN5BZq1/ItVxc6dl1TG0gt55lyGyOMEWr
msfdb4gId7Senj6JIOT/bDRWePU8ApIIM9kzc/VxSsMiIEzXZWK+0FzygTAGJoaq36WQPijXRUEp
KSFoZ3QcO/SLAq43AZB6rTEAJ9FhjACCRE2tpla4ZLyLN1Ih6YPDxOaczaYJq7qkmX4E1Gvqr3g1
H+3b43EUxuDDH+Z4T3CE+DzKzWsC0O+7rlJbkwDlZKQzUjLDOVyU2ojkeUuJQFE3KFnWKhxeMccj
2f6AhHTrqQBpm523owccRv0eYmLj9n2Rl3kk4eewmYb94kNz+4NLL4DQ1uk2MhjMIAGW4TAimhSr
mHqHseK/7OyvZPxPVhCYs7GRyWQXdjhgjhBpU6gjUNWpsfFPUwZlbUpUgDlZ/a+E4imvVHC21BSF
tUTlPyz5qbj/+iIofcDc9hdFYzbWD262FgTe9PEJkx55W4w9DTJ1+IbI/3zl+bMVCpjeTTLtKtjp
3QJPtppQM9TUlLv4VTHYSM3iTE5ucR+vZ2z5Js8qe+TXECyQiMeSSgawsDrog7Enh4S+BUhHlj8w
o2tFNEX4tcAlD9jcrQ52z13iYzrPv3im6yVYqChbtg9L3XeUbRxpqEB0LuInLmsB0rcD4PwDVrap
/wI=
`protect end_protected
