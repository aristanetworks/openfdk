--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
cMfVX2OasTpSS2n0qFpdQ/v/1spgZfKTyWDNkbahEVbGqPU7Z+fqMFOMxXwXT7VfRBFw70nPzikv
SJ9qcW/g1YrmlecIRUY37/z6RZw7RarB/0bzFkb4oLcymW1pNKJE+5tx2+XE7teYCfEFYQ9mH0t2
Hb0COhPMEllSdXUCCqvyFNalgxo6y6kiuvfb2XeTTUxeaJ73IcJh6jyoeFhEpH63ZI4rRlNnDD9R
ApVvcl5P7JMl6OOABba9PkeHPWWeEBZ5dcMnxJdUxFEf619XhMe3OjXR4bt7fsVnL+MGNy/nMy4+
BLSTkV/jjRXwSQpqCp1Lec5LrpcU+7CdBNfoJA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="7FUuC5CBk6PdaqQGwm6LBALnaeIkpunYemGy4LSuTU4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
rnDegK2/DG/nKrpzAIfAzQTBYZfX5RDPJdHxhOPaWn/TaJ2+ywqhbDDcoOJqYAR8GHFrq9lZ6jWT
msThFxREjje/GjF8ho6OM2w6yomYSGDTVC2zPagFCkFNU7At2BqYp2h1HOurPcGLIwT4R+rqMwwh
1gghV+5EbPRDgwnHXckTII8sIYgHT5wiKlmt1eCHVT1qa86dFKxTEBC7I8ppsFlYU9PenmKJGWlx
CJ602XHmplZbe8mcq2WRJ6ywLRcOc6fMikqBwVyTasKqshasi0L0gmKLyfWLkshXCB7Fp26JjBCf
vuEDatk/Kz2zxH5xj2TA+h3iGdnOKm71ikY8/Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="3vWqXT6NzN1yIZW1nwZALl3vqoiX13eTpEVcxR7Xixg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9440)
`protect data_block
8dSYVQOohysBuN5iwSZ9LyNVJlJ0GqSN2JgpZ++55KXdLJIm8pnSl2jjie6zqUGVsYe8V1zW0Dii
pAjm/XDFbmmnsU7IlL2EP1HzO4cplPievq8w7E9C87+lsfG7cNbyjAW75XgOD+BrRqyktq9iqrRC
JjgMoqnmi/d9UhBCZnW5Xcqf03eulQr/h20vdZzKhDiPMZ+UoHs3oTfYZ0grRh+gveVBUr9ctDGs
T8yHozUZc6Ex8jw8v2hTCa9FMmf0yuvd5uFkR4vk8m/nkwqmZZ2kK/rttvNP3AaCCLnBDsQjAzQL
FHDjkCqMHrm+BxIvVUbRjMzPzdC0J/CxjEvCL9ySRvqxShg1Z4++yYMRxO8j9iB4iLbhSOCozI28
pyvAHBAj9IlRy9CNUpruvuM8iCYNwJ/i/meIqIGohwVc6Fp/TXJanv0BzsIjEg/XM7JyKciBXZcR
LftBAorPzquaR3KcRy06j9UOgRX38GbKbloZlVMhZagH1X+V4J+u6rxAZw2Yl5xttpB80ubcCd5X
6yrAbRQaJRE08/ffnyCsI7xndlibCmujWuBDynoLGXQfgdEeF9sc2xNEQDrf/e2BBHLrR3vfVYoB
F2kuTd9gG9N2dw5nth8YuC/9DMNVpMD4Ju//XlA15LRDLTjoReEFu0vNOdZ1RWw7ZZjqXHcc4M7T
kDpTctsJ3niAwBMPInDpRRVokuBgNzGpXnVL4SyWQErbo/lH2V/D7Al4XFwIRi6lVlMq4o8aSAfE
M1Q5khGxfBDoO9sQGcxiRMN0Q8ZNbi24uuiyzZBMHDnu8yItjNO8SIOeBYgFwyC6IB16mAgc9uyN
uXZ1hPUX268GExzCx4J1haKca0gNLivA/VOgXouPodUw3zI/zh3MVVxqDKhmHMYm64cVwKFxLUtD
DpglUnGNyEe5rlHYHV6J0foW/1fMb6Ywtwe3rXpMNBXrCG+IYE1caxyKwjJ7jdT2UwN25kjmYxjf
dJwFrlhEr218y6qbTuCFddpOTiCYh5vZFLH5Ap7G/VRDb7NpjQbiSg2XNvPNQsUyz0lzwUpN8BKh
iz1miCzQ9o9z1P8xFHmUWS6Fb03K1vRlI3nf97psVxS7dXActHn+AYjKZl/+Q6klex57DG8KZPNc
XT3vUliWaPWZYhdRRKsXfmwoq/Zx5AtF6ApeyrDqN1f4Iwsp8DdqWlKLoOOPpyvXzQOXvxuLVkoF
HNx/GCSLmpuGDs6M8Bs4rpvAyxlhflO97eEMkHMgtpCQamAyKeVUPYQIjlgE0kHdObaB1Dng0qOC
bsxg0YAkbtcvATHgZTE+I3vfRuSScZ8Oav2prO5VBSldOoVcLI2H/r31wvAV8iR/0Qu2eAQApOyA
GrHaBUysA/bVE4D5w/DMWJ0/hGcEV2y08xuxl4tyTe2rn/1kCidJHwQxXhMiPRxe1k4lUSI8uBXO
fujvF/PSgYo57URGGRQy+xhmOixPzWn+RrSHqn2AaGLOK6lEfz3GrF/wJ8VuFSw/OxKtBHVfsMzb
SDbIIveFjMSH4lZO2KVZ/pDdD8oFi1i5F1lFUtuHP6ys6pOU+i7NMLZg4E7YADzv6Gkz/Zc09ctT
koTphYYZ30q3qACnOj6yeGO3HXDuhAU62vz6v8jdIKyq7vKi6W6nW+QEBwOlsT6GjDutr+CCBwcz
Su4w7NArn4r460bOuRBlJ8AK9+sRIPgwO+9UHvynKMFhMN4X01h5AE8DRDA3rGQYIgNE6DGKy8I8
aOgq6cf/nMy7IfjDKk00qntMghwq9zgpBjmvq9AhqufEzi2yBqQZKYyoI1Aib2y0gVK7dhHJy4J8
rxwkOPAT3JAMaJIrCZkvztMzTra6E1b6LJJtsKBWf5txrIl5N+jVqR9OMTPhyr7T28t1+2WEcqXK
Ib3UFCCsRc2oCapqIkZnJdVWdgt5+Yh9Fyxf82HBmrFmnJO6SXgGwgFjJ0txIdm4zrRr2iGeTz0W
eUUlIbT7tjIvXn0YxfgupBvJ/Md78PMexbpnzVJnlI6XFCnlem6xdJQnGiw1b6OZJLFUxJHk2pif
QIl3GXq1KeXC7wZ4hCl/6QMswzRjpx6kfQzQLbaefeEX/dr/xSYe2HKIYMjERmHr9EwgO+0Zykz9
Qe4zuCd07eVH1xJ6cWCpse4QEAE+7lMETZK4zb4Ws3mRn46zoM+et961Ir9mdXXbA8M1/b9ZcPVB
NfM8Lam5ntqLsL4ZkBGbB7v0AIKKRFlBMHLapyRnoOo/+N1EMf6T8VTaQvisL1FrAX1QEZJG3dUB
w/mp8mU7F6yGVN9UBKk+Xs25WAaOwbTS8lvhw/ooIaNkutbAdpwbLqzQg+hXa7/WE+pWA1S8jFiP
oQD/gBCppDDplgBnAdOF6L1Edkids6aZ22Q6VNtR2R9bw919HRZew9T8Yk26mqLRXPsN2zVH1Z2X
xp/APmf6B6HB2TDxtjFkMMaNJ2tX9MH1NsvGP4hsEzFTXOmxfH1mLcysAWUghja3Ja8rXIvpSR4x
mGrb5fcvBj/Kv1+Q+kRnkdK46bPVrK3tq+qqd/qKTUMdCfk1/jUnTVK4by11p2aSj0naVv2a4mKV
5lDJ5MxLcHGq5HhETs4GW6eTWnv5STpRIi1IXrDN42Mml2Jqn4hI1c1JMX6MjR88gxVW/USnppzV
fyDBBNwYQf5q/PTf7QMGbU/4CP5GdSEjI7duOq4d0HEippcacSTeBhTuSJUyHR3VdfTmqcr6yLQk
ZytpbevVvksT+cG+sxPDHHDjqUb9kDM4iBzzM167fvY70wKiQZNCWUdZYhxiR5kJ/JuGGW4YPRMM
aVpcmvE8ZLeihUCmeti4HDTmLbGDOiiN2B0eQkJX22aIU3oXiUbPGVYDPm0LDd95MRQiEpgJQnQv
XXTjz5FQwmiW38ZtfnyaWeH2T2Ee59bMSOb3G/yjsrdGEQgaqvIp2G0hDIFHIn21NB9F6x/27Qvc
U2gO/PTFoecxG10kb3IPumVMoZCcoQZMt85WM9OshUzGB9rrOfeoO/URQnyBdzy6i4Cz/nqJHAlV
vICO+s2GMffJNSYCxoId5ASil5gne6YlfqPWIBvS1UP0C0Np8RSuV68O5xva1p9cxNaA+Bt1GAho
tzUHaCoEaD/lFCFqVVwLe98tFKnx0s5WVCTbR+xYyqkVNxN2PoT8yfu1PIxY0ypo7CYnLHpkq2Nc
PhGkPe35a1zSCmrJ/oFuKJd9UZ2has+m162FR/XGg15P1G/4OV4ytXsJsaACgMXyi1V5Rd7FXtBK
r/B/0kileU5GahTBpdzAmxyCOnNsjTzLJUnoD4YTyDNEuBsp4kgGiLL59RwrPkUcSctYppl7bDoA
5DyO+kWPhi5hmrQGoyJetUNE2abKk5/9Na9/MoLjp2/pgVdkpml9P+vwuejzdG/E77c9XqD2WIFM
Y2OgxcM5UBfV6VMBRmJzjomJdFh3S9qFnjH81in3tbD5zwGYgwubllIsSPIgEpTuv6e6awL3HaXC
WgcthRtPV0tdiITZu+G62143NvEhcBJ7jp3fG/gIK8XVRIOOOxXavyD42OArhF1529bYTBOEgZL/
qXXUhrntssvyWPPRpyL++QR89uG+Ka7RM66e/XsmB6WO/kvqa0x89T1Au6D9a0OZ/ok076T9K+hd
CySUYqcug90r5HCNAcCsbFeAP0+jH0EX5/f13naRP/4unG+uxQCMkHquTfIEie14fQzfaD3Qe0jd
Lb9Pkjpw2zSJduVnavGNlwL3FWc2vDsGWmZNxav8yJekw6lcrGOn6hZOmbL4oXcOgAErb6yagUal
H6wCsDvxSg820fwkVRsbQVfoN7zt/9hqfnOAyHWqm9mHeelr4cULbMraxJfNMcl9cuGr2Q1QlpKA
wGDTFVgyeMZ26633M3lBFflWRuodP8BhhF34HFpif2g4BT2QON8Rlfs6OQPwJS8nWpYVJz/79btm
lF3wY9bBoS8dk9PHj5FsoNRP16fQ/MY+AJQZVKtdPH8PO3m1aFbIUMQvwnuUY9t7mb3HEgqOEu7V
WK8FtsV96uP+Ga98lecUVFP976K1ThUWwYolv5GIDENxdf0fmUbPUh1CpzqwIy+FVd8pg9hrYACa
HB/KjwUGMfXrfxeljYFe2lNvTGe1RVGQyazuLCam37k+MuqPEgZ0hCuQosMbyTm33sbKZex2JUt5
J+P/vrHuZEoWxSTpDnuKYwJdiLKG+C7GSqfShQ7SbJMaD+3qcA1JhVkmjJ9Nl2KeQzyUCq47QZDO
66YYW/7yFkMrUmhQpEBtcGMnR+QoNWp9JPQB6FT+Gb8rk4F3eyv8wHui/u6/K7rrT85KsYByXB4g
vW6F3GX8SeSGT/aQr+QLIL6wMivXAFJkHaJaaNP40E0+ZPp/lnQCAN33erUQG5GxIrAxNGvJUQTJ
qAosU6AOGhMOsfqERR3kNoGzVk0dVfCmU2NvqZU+Z0DtMJfvpaiTk5MF/R35sYkDDaMxE6OC6sxE
AHQJdFQBWanaDQdRObzvX/eGevIWOHwJoCQf1mjeqrnLqalc73LnOOLV36gmzgJo2AM5ivtcH0mh
IAJfBEarla3A/Eib3GIUccxI+3M/iEhQX2bdnck+qVlQdmibeUyksbdyr6tcyXteALEpYmLTZt7s
SnibHLmjBkGxT2YU1fyjzpQhHbX7SuBQWg1XjqjGE6TMJIWeR3JsiviZR96snHNM/DzeOyoFSLh4
xy36plnPaD2jPUVJqyHpnsfbAJ8K7l2IB4NytM/enkg/ZXgLLUkns4PywA2E50RwBJVkryormX7V
RysUDqdfVRDv//SsQMM15+M9O4xQcYYBAlJWFvqRcKI+oCHsQHDYl1ppCkmXZ+k0sid8iSejfG51
Hsikdvgv1ugFiG1Aov4eTmbqnK/DpIr6hQ+HzYcgFVHK+OE3e1pnV55DtvYpmkk0SWPVVgr9D4aQ
7Vv7dHzs1JBOCgbuqJsvpJSJo4scrbmnNYdzIphJIlnP7fNL1PNP+RQHakJb2DKZufzR9y+Ta6A7
t2wLnYLPwzcM8wHIZCUtvaLvYDRbtpW9VFAsnBsVRZnirr0sCAJZxlhQGiNJe+oWZ0nnyEDnyyj8
G+aZMIlx4+xzWPpdyy5YuhPmOV5hB2zGLfLhLsLvhk9iOHFdh6QhDflIzyOx0JNpkgS0h8AUMzzT
zmIG5gwWJRgunrBv+g1PFyL7Z7i8Vm2iJ7KWk4nGXEBafQJI6pJuje3kAB1p/+uT+5aNQwrj6Z0U
oeWApiPDHyfy1YGwZgA/RsWPHBSoJNDnQhR5Wx8YvIo5D3RpHtDzc1bD+wFXPsmazE3vM2Jfcdde
tO/xjUsuWeyZddGsOIrFiOEhLeJhK5omqBUWzfr2vZ8u8mciEcBld38ryiqwHd47uI9hcDZr7r5R
W/CB0E9FQtkcU6l5/n/LEiTCRwlApg9B+EtPK+DWOG0bhh5mMs8yTEx32Ou1UhUMM0MSKG4yZ3KG
OxA5Y+Bu7+oyKwJzGlEEJ6yvFAf33zvNxF+ix8cfV/QZNCywl4ZhPHN+KcQrSLENKAZF9rRD9COI
E5HOOWfjEIraa7laMkHGPQmb4ncqqIi5o+zqg+QrDCar0nq06im9fy/ln5F6RZjc0SMQsGIe9AD3
EAapMTC4wJFJWU0Ks4lZfmH1lodqh9+zcS1XmmowaLYtR1NK/2YWoPEL8/K4bzr6EA0zYEFZ5f10
UAQTb1naSWdywsVozZ0EMENljB7NzumW2zN70era8Cke2bsDxIBC1K/B8vfjYvWvbJ1GA2OQanXB
8rvNBmEqqO9R3LGflHwksPeJ9LAJ5YyUekw4p59Hv/Edfw3kFOKcfxLJ4u1E9QMvhesFJMubocEz
hxskV+Az6KUMBeva19zKu+dZam86E2PlWGegXJdfoPKJVap9wGCCpN8xqGzuhnPwW8hILlcBDsRJ
a+ZJVjakBkXTR94V/nWd/n4rBIU+kb6W66GqYoCFkYKj4eE7MYZgh16MEfzhWkGbk6bPY1mRUfdu
LFTGIbuLjjSWMYLNSeKv+bASsw1NtqF/qxlIYN77gJqM1YTJ8VirsB6b2l5KAyACd3nXwxNpFz/o
XBMEuHOjH6KdLSwHRz5QsHhByGpdpuAK4PyYXb2Z5A1jyfZXQwgAsJe0pUcc5NJadB8BBFcyCjYp
8ucvulX/4QeoI18VqSuq5PxbNQjrHIyHn8PcMjoODhxSYPr9EyYhMMm+wJju9deSziSx5PqTNWES
RWgkQU+LRRXlRjdTFsBKeFF+44D7ssT6oP0PIbeuKWptK/GqrdmSUm9VUnI2TUwAxHJUReYmT6SP
Z26eNwvYQH59a6lNf4fE+BjRv8Cxf8yOZ3nGZnBAA3r8ZH2cwCU92KJLnOEvuBFvhM3uq7C/8MyC
hBhQGE/IW5VIBcBGBvgWECpJUPzDuWrsCvNeL9l14g4pU9eQR4qzlSsye1VoCSWGMVMrBofVBesP
DdYPll6nOLlHtiFdbyKCZv7NsdGHRAcBZ7ivm+vxPFB+9I8qQfA9tTnD8ItstWK5E/A5TcXvSgU6
TGzTyN3KfzNtUgMvUEcsKrBwzNKo6smtDqBLU3Y/xQpM3s1BRFL70/sQas1YzEDzcYciDkIlATBb
JsSjZRhIdC1kHlk6V9/6tjj/PBSpcXR/QjAGd1SFd1fnInXX9wykCWbOHsdPRqaPopLDoxy/pOfi
qTzzsJpnK6pUf2dCZT1qXnv7ZxO08nH8e9B7qgRkzxG56CTlC/I79QEOAWyP9z/UJSZaOJwbP8ws
x9RJqEyjN9wUm4J87PF9smEdEt7EfUA1yG4CS8nKnKT7bFkYJ+g1zoxqkdDtHzGM+dkfjPz40bi2
7KFLQ1oRwocvfFiXQyskKCVapougFq+t1H9WsEQYC5yMPi4FqsmtzPo3bJa7t3on4PW9i7ismcFz
Voz3qN9sTn3TwPD1C8JXytuu7oeKeccbf0npSzr6drtGjj7kFRDE6gcjPDpY9iSxaFK7BD835frV
d2Grh2F+N3u5sw77pZTtpOINYIplCTtbMu3RMr8s/vQslzCIAgkjpHJEsHODsbPPdXpCjQN7Fy4v
+M0tNQtaqVtSeHACVAdM8RvZq+0jwm48q5evndiQh6X8WXaGXz59wE/cOmg0wIsYwHBYBHyYP9Xs
PMZrJ10zqnbGc3VYlvQAiCtm+jdfj29wcfsnDlwOaf+/eI1mMeRRv9XcfNnT+8EpnwMqFbEEnqi+
izi1o3L6KmlS/rT0jy+186OPHrMu+hxy01ej+KLSnN+l8C+m3ZJkHKSF9MfFMFmgcwxcTXN/5uFX
uFdGfQ2E4LCDaHuV/3MXJGOvUBb0kW5pAOiWcCnqiCq8EJTUCpmHBaDADjGI/UHcAcSiEdzvqhNe
p7jeijKI6mDVg0sYyvlYX84TZp26Kib4K+YkZGlveRbPByJ7sBcotf7acbiD8Nb7QBLQxND/mVbC
1SGumKVH3xXcNx7FQjaJhvoIuLx0de/JrCdG+juFaozy3ZhKpr6LnMQXKlD1JJSCtH/JV8T4Rer0
+53FyvmX5FKvS9pTCE41D7pb5tfkt2Z4a6E7J9pplXiB0cRiVGTk8toFldE1XwJwQFBnAmTuCCY2
l8B571hhD8P0N99cO6y6URzdFut84OIRS33XaW1hRvI7IIc9NKhuA9XAJkAH/9cWHFMQ1XgfxoWW
34+ySJOQAM97RPOAYu4HNq0q3G/UJPzu31jGhuYRnYQzPemjChvh6sOXDQY3kq8ifx6rgpfOuAva
UtSOhgNDNhCmb9dZSRY5iuDEZE2zwLn0GbqWLZWlOoEJP/r7ZD1TBMbL4IYYfoPtcY0WIoERGnX0
5qwEv6/GRt79IvGlkwXYGueWKqQmX5LqLFAU1QY7QAtHXCs95/MbeUy2VnFz1schtse+ynSybRgd
R0UKcWXllkIUS8KEpBtUcV6uD2V7jAV6JE7b2Q75gyQaWksoJj+zUFFI0x62lcMrzZ0JO7d/Jseq
eTJiX2iMLDTm/Iolnc+BILP2Car8nXAZ1ZvEiiLpkrfLZgFimATf+Ei8rVvAyVpUSVyMPn9riPfX
SDztD40+QIznfHjPIvoZwwvL3HDCMS44d9QmDy6/5OZJw63yn63kMNU2nppJrqekV8xS5orBKkdK
W8HLDSq8zVOCxFpPwSTZcffhQyIFji+uXyKwJRwuc9d2YNVDulyHplheGWbNxH/Dmavqig8dA0oU
MJWZOez7kHEyvmHhIAP8FjHqvzkozCGnw47/ibiRaN73xX6GdzlJoVhre72upfM2lrJodK8WMHvJ
sufVJ84Re2INr7nC4teg3ZMTLGiSfqy7SNJ4l4OdAG66y//CPPk2JEvKU8c8ko5JOEN7MYxSP6Ti
CotG3B1ryFRg0f/oM8miIu8GVAnCfvK0qwmBW4N1frktudo259Ca3nZfA65g1nxH9JEPPwk71oK9
DIYnoKKdw/r2hf2vfCJ62XgB20XWvSUc0hXpy2X+WD76wAZK2ZMV5BW2q0RLE19A1eakogpgCIIJ
raFtC3MMI2HdytpFfNtNl4g1XmcOnKnSIg2sElrBVJHtaAoD8AtKzfNru5AG/csCv79MMcunOA4v
vBwY0GgCn6JPi6sgJrsf+4oktuL/lm6aAothh8nwBfSl7JwBJskjSRoDbLKFyEn+GyGCJqArL/0A
R2GoD7pXJDDKqC1ewKmP1v4PeF04815vePVZ1UNzX5rokDbHluqbf9wjr1Yw+jgZGxzV8BdzCkCz
kgWHG7aQXqiQScKnXasSccbYLTcpMc0nhULpQdTKnVfYeQjZkqNFHrt3R3p1O+N1ACkWcwkBtwlS
ttu6lOSQQDI6si9BzAmRGm7OLdU6fwlW9lEdI/Is4sq6aLFFmqD0/k6gJi0PYpqHkEYZmke/EwSd
/dXtDPOEHBw6IIUSkC+Vz40iiTfGPGbFNdukpALDpWMMni4TXSXf6RLskbFLV0dHIR5Ko2iqWUKn
gmdDzkBPdhr3t7iALCK6VrgPCAsdyjLUqBzJcTMHpaLhoEKdDHSY0wmCelJTBVcw6pblnWc+jjmI
vxoyXBziyMXvIYbzYP/t/gWFg67jq//nC6+/IOcnAfzOgKtPmyrkQ2uERlTfxMZClFn0TKb7Y6i9
W/vDL325FMCsl420qVXWgw8k212zOTylryC5ZNsVFjVmpE0VDQAVnxkvDckl9F3rKoKZ38kxctI/
T5j9Q1ThhVpJ/B6RuWlRWEI48nam+jLA4HG96+BAOUzUFNy60I7gs8E+LRurkQ61OzXSKOrD3f+W
zkaSAV7z8XGrLZi7z9GfmPRVBxYsbflZ2WDZqj8KKh/ympXb9AJkNQiII3A2GaFmTqzgvVKhjEnS
e36zbAqvkJwkO6/+1Q7fXhQTyTZ5gCR2gHK8gbgORK+tPxIMvklO6VlX2ISTCvCIoXto0dpYwUIu
U9P8f163sp/xtrJBj6ltNnUDtZBbhiqUYJidC5IVfpkGyzYI6JUVojWBEdh5xZrPpyUw1j0KHugd
fD5u5kgWqdqYQ0PLAKhN/qUFWDow0tIKp5rtClvANvoMcjsi26uQPRsgeUW+QYaZviN8yW2D/TVM
vvbAg1PxWSbyEJD9iqgAkojDnwK0m47RUN0+AkrsRorTzPnbGf3LgE5QAGqDyte0OXWFYFn86+fc
Df4N0YrpWXGtRYfzp+Q6cHWDPqfUVCWhglhRM3Gc2AdTAOhhJD017W3tYFRIWTQoLt+Xbc5/vI8X
dYmMvnev86rdXKN8/IUh4Kemslg1LTLzoDgYDDxpOFnu3BuTWf5caq9LOMDYbx5oxXT9EpZkBIc3
LFHy0LuPCtVHMKvxz9pVQ7hKuX9/kPtWqEE9Z6z99eegsB3PoOwpkhV2sksOJw7KGyuATt+2G/SC
hfY8E0s2z0g0M3A1tslJ6VIzGy8jgRtdLxinfVkzHPyfJSjyMVDu3tkGKG81tCPTjzOXFBNLGDDr
8xWKxbZT+RMIXBLx25NiBiLo6PMoxEaP18NvwIDjwMLl363V0+InOzXl3YpZZR/uzY4QAFJkOLTu
78mD32czRNivG9J3mBUwv6GlFcUCACyCX1JW+W9+EmOrg9tRIX/g97zqgymKLqJbwaEBQ6TwaB3E
IgREUew2GT/vY10QM921p2jo9VyP3Ee/TmyN0I+TSDL8lXo9rIqzYThHsOmLTKVx1vj6S342LmJq
5a3WnYzUupv0BLeEElz8TVzLTcYrpoAZQr4dbVur2NcGX3DcvPZHdREmtOkpqPaLAmIs9VnOLkVL
tfC4c5/DZkZbykUEIKI8/XyywsCRfr9ZF7Nhe1LbVfvFx8p7Cc1MB87xUQSLfbcG5buTZ7vv9Qza
HOYzLkqnX43kMGoZeo5tHcecQUm9LUxvoJWKGssHmZJBfklFntUmDmDBrqF06O4eH9XBY2tqmxqC
BBqS2iqPbvaAHZ10HlGiHJbuouTZIwvU88nv9B7/MxNceTpQEQpBcAvzDyDyu70b7vUwhZDyMiyj
qL0BX1oADl0AyV1uAXYq7not0MMleCw2IbhHMBJXurOFUCFzUypQ2loMrFIwvfQ4TWYCkCtA1ule
uz4Bq7HMEIb5YHt2PmBB3Tc6gJEUX/v8uxlfkhvXMTp04rGvfspJoExzZbdB2Jv4fdveAY9Fa+cK
EDvCOx0lK6HupXG7sMPLYy/q2ZVKDVHVI4mIh2Ne2MJ9fk4EtNLRxwOIP28wjrnngAA9thQlAdTw
n0WKaJQyv3/1E/q2L66DQTtx0PRTnt9PaOnOGVMvTj0QHJO/E4xDyTy2rSrU5cPg/YjbShbG3imk
WAD98CVZ7IW418ZO0rrzqPA1qffjDdoNCal+z4kQ//pHDHLXL8G3001nx2RGda7F+ChGBB9SsDF3
LxsOCZ3JXZ9SZsVNvH2QcgGcsLannn9iCN7GYiirMnz8UuCgHh09mVWlOodn3BFx95gdR5c6rNwx
F0BS4P5c+dYoSLdSbUhVigwviNt1D5lAir4I0zHuRHp2pQDqTf2xSW87Hh3AqFfIEwZ3jPKyCndC
EcIkO9gzgIBZVM5OGivTYhnH54lrtE4ZYG+N3NCtp6gWJDDEHK/aofNflcFT2HPUG2ARkBhtVCig
UH57H1XTBlcPTFFuR03EchAmeAKecSuibAREb0/gItxS9ewdmwKw3tAeiUDN4CZxTMdqLM6kPkfe
wcvpH8/i3FYzuQDEJdDighuwm07othk0lhYab/VaWU3fHOrHv7Ug8QWV6Eexd00lW5olEhUOSLDM
XGThLX3HCoDnSEnC5J4CU2f62f/zpgmIbxTtCd++H0OgypW9jdRNuZCPXZ+fITDzSnQJIHW5TQG2
Nqkmra32bRl9Fr0l1z8QpVZN3wowWIM+ah+ci6Rgy7Gte+m17dus1San+MpCF8BJEytRfHPVeYOj
5xGNRoRVduTDRwF/7ByYeor8XZB+FcaWFSmtFxjvfzVIghz+Z3IjC6uMooj1rbiPdqRaOGCIPD3/
AMH0BcjxL9ED+Ui1xLdgeu+kt5dDM/e/4C0XT+zDCuDhNWFn9yHQbbCEjFlziDQd19b1qKp3rtf3
uKsRw92vIjXeDdMqwNfRMDlLD6QVvMySotTK2+cvoEqawDZR9gxMOUpWsdICt9tKHk4GYZSRY7vZ
mvphTO2szC89inmPIZl2b9ljhxgG+GhGLDQX3h4NCwv1w5q9Z3Xyli66p1JL33liMbmc5I4RCQVX
ZTEggpyAkIgmQnezuk7mFAMoECv/Flk6VEDL7Xf8tdC/JkMvbRJ3tHdU39QER9jGotJ9wF3arEUI
7Nm0ND3h5ohmZAe78kpTE1uBMgYjgIJQ6H0Danz3eNbbj74b2ffzRBB18wiYYLfN7Wf/K4sB+ggm
IAh6kaZ6EvwId1r5e2MEnqqQd8VKbZLbAvxIuTbv3lVjiGF2kfjzCOMq03vZeG0ogstfaU13VGck
hY2RQXf3kD9yMASeZaU0zAAoPOhHncRX/ld+E/wQ7ZiFdSdBClpPpofecKIl64r5jfbp26/lHjLV
5LfCGkBbIXjCHl5zUZJcYpYPwhQfdWJi8Mt4FJaTKU0TquGBv81Qie0IAHNv+Z0o4Y8y6/bw4MtL
uEG067bYz3U/+jzNgIuQ35R8Qr2EUIRUS1xDVidhcOUQTVaRNqnW90XHsF1YRLkfX1Vnnn8JpHkQ
w6Z5um8m8pjgxQJ3FwpsvxweKM8OgxuXd3VykthxuWpYLGY/FohRQQlvR5ZxTrZ0Ue1ry3rwaBmI
ST+ZUFEN2TPvxeGM8E4CZ4YxwIDG7lds443AaRi/w3lVPRgHJMOON9h8AqOk6wDqpAhZeJQOkBtH
3MEMfRfq6swTU8tJqzm3TsGTqgSyKco56imxl7Ag0UlEKKptHHUSs1vC2Jzq6TSTno79SYS9eXNo
ofP76lNGkM9ZIka2GvhZg4Kr8nfqd+qdjU88n4XEwZQG/wKZYc5GDKl2NmFuViDKPDTxOt96v1MS
Ol9JpeLP6vbJRHZdLuJB2f1y5bALJPKE+3HXifHJnFrjypPYxmfO5Ahilr4xlr+xv5z2gBKxI4Xz
RkOxmppe5PqXzSd/fsXhy99UGy8rGgtM/acqnVRdgS4PVBU=
`protect end_protected
