--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
gtvEEK70MgHJXXCo57ysNwMoCeS8VxXUsQfgcSgbC2+sp/kRRDYBPUvcsnxw2lxVBBL+Uf54bi8j
lmt9G1rXw/xBNC+dhhokZBke8WYlMLSwj0lpJsvTRADvKFterfckqA+4mfOzkNsdU+54GteOhnpK
yweGdwJgaYZXieQ5NfS40eYntTcz6AxNCZL8fEtGEr/cRUWX31kmEBZ76t2rNj1S9Bd1jYabWoH1
bXERvqGBmPe4w8zFFhfRMPPtexSbmSgcKJcqpXMiC7RBDEYVPdjtqHMgzYnITMwycrUY3/HErWoM
6+jAI6cE7YTed7WpjpCsKRdPzrBrHW/n5FUTsQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="70Svn16qJ4ZFsYtku/IqOiVdot0gZw6PHAeS+6se21M="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
BKQtZIVhxsGryoLDQ5O5i9DAsyufJWViVydEdIKejvqHBR9j70FMhcINQIVfsuX8czjBGDj8sEab
FyQxcINKZSr2FcZ1IGuIjzJ7CyCwap+toW8EXH05wZDHh4lOdjiY/8wJeJ/uyRyZ5VNwUFIyuSzP
ni5cVqZIsb0CwZJtyuYqROXsX1+1Q8BuXpIyk/oAU99ojE+qgpuRQv397UmLri7EwluYnNdlvY58
ar9EYyiVP2kaj+kqaLe2/GNTIqGTy3TwT8T/mtPEbHz3qerOBhiQyePiboZQ/SY9SFoyZzlFbaVe
671I6+fWyA6sM/mcsFaBE8IVXAC2Kt5L2x896Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="4bBxXqSaLW4Kukdc14AHbirLSovyH3E8a/n0sw/E0rY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2464)
`protect data_block
Eog1I4YaeGuQwH49iWWSWimjBhQT8a+td1ajTXJWsz2jJ/y8nT7FafVHprgV+ww7qX+UeIHGxxIo
SuHRoytMeXYP/ApePz1yktNKm7kG3xKiPbSjLI3Rsv2ikdbnzjDLTKV449oxARIJmGrsPnRFV07g
qxtp4c2nHzMp4iKPIiT8K0iAWTJHsQtmo0pgIq7kNy1SbiAbQr8ZK329OGjiqepaVlAav2T8/BpX
o4CYeQYI2lWgo7ndrnPhpnyWI9V39k6NknXPrg8OYIldLPnQ+0aHUAP3+Nlb+pjolofOR+780NWM
PxGQItbOJO06qxV9hhDXCqMMmW/9INwMpFe+We8hyG61btoZYtsDARO1J8yrky3OICBKGkGStDlz
15llfXpnZ9UpTAc/KjX69RnzI7+S5PIPQ84odVWjwOvbkB5QTM4R8N5yN6U3sDBUCoTNO4sb5hWx
WXgeJJNeu8KCw8N52iPZZNRS6ie9iR5szEVwV05bDEyJRYdW2jUIdks0JEH0wg88MXBC7uood3rn
IDQMBaVmWjbH6VSTqXlweM6ifEKeBHXGigI1l6NDjHzpFCAh9ij7Z3srTgIb4/Zm6YJupikswUIk
fZ+oBmh2eOJzTiZpQ/m+pLDYS9A0Yp2UrBB6HbBupmJczxfBB7xHN/5dOF7Q7tCP2lldzcxQa8Sm
vG6lP0DQ9ZUAe+oSV4pGtRTYYYGAzxHq22FXIdz7xvyB/JEGIlKhE8KWbsX0lVb1oIXDqXjegECW
c4HrihTAGJKLvAmZmDF9Efre4u7LE3TLu7j8OS2ueeStSnEMn7W6I/22+tVuXsrJdstfhn/P2EXv
eq+gycruj/sZVcpG+LZdDdwxr8DPkX6x9/tZXd/8uY9FW3mKtvAUL3eOOGKs5sxyxzqcAib39Pbr
+isBS0r3g+y0EtGp51H0Mp/7pVd1lLlKQqPe/PqN9ngqPmEUT2JPlH6e5ui4R/X43ftO9gXx01gd
pXT8gkpVv6iYhmfxPCX26Ts+ogrm92CYI2lWl9inqTmWvADJLKwBHW8SRanyVwSjsvqVQS6np5kk
IPcNwLT7O3bI+GbRYZHR9YsnBbaw3cX5AQAj0EF3XmACDPaAEFvXQyaQruRUwa1oxcSKk2Ljt4FI
kXFKpCK6yxILSC9Uk0WLnewEZ3ixC98QhMAuDp/xvLTjjv6sPfU0Xz7wWT1DuB9xEkCOY2CIun6i
EtL2aDxdN77Rn+4wNhgEL4rOi1TQ5PVQflwBPC6JYJQpyPMkXaGrmrItAYbATJ+GTvdmVwGShMka
RMZD375Q5VEq6vohykUuvYrXdYyUehfMQr62/mkikgt9Viv7uhG9uf3f6ucAcVC5W0NYPPLDyRse
LlEOicuX7Sp1jezuhj9lXjztE9sH8zAS2Tf9A7etswwVumBa9QequEFyLYSknu1MUbW1MEVblMUa
QEInXQwvWELkTWi6DWQBFdxcTjlEB9e0ZZ/b53g91cqtR7z69e41S78bvL7aNIWStgFpPuPQiy+k
//0NElhghfqDNjdt9/fSYAVSfAV+sE5gwMUwqUa6EYcCWgabUORT+tFBdX/pS1gG5tYNIQHQT39a
I4oDf5XCuLKf9afpXWqPdc0/pnIXVqQzE0jOCbNjc0ls1l5hgiI+60vaIMtjtX7IwR9ijJiBXh7p
LyeAqcT0qKFEG7Y/xWfddiQDxhbtBti8gbMfVAQMfM2PoYzMmchppinAKNbcukZlxk2NuUlSPSjx
A4PZnMP4RTq8MGP4j1s+gsXTVqylIcjmmURtlVIs5YRghABBzPCNMacIOos/q2k+grGZvtb1KDBR
rcgpx8TUg+NKAJqf/oZlYc5naf6UdonFivLKXBuJNxLd5mHkha29Yl6gpYkaCK4CJQWBoOIBYRJ9
oaW6b0yQ2fFnVQC8x3uomp3hsO4F4rAS7uRjCXYpE4iOfIiAZDZMo0Rd3UxwPCowXMXeT5elJFtE
RzCRSgfTug79NZHzunPxN8WRS8bH8vlus0WxNNn+rzIyDED7SlcfQI6MDKPe1TDTEdo6qf7VYAsl
mhXb2f5AENmLNkfxSa+4TFbulBLnCsybIlVBuKOtOcVwJhWxZfCQKjr165911O3MD1qI+ZjKqNqc
TCNHU4fYnSpsvCftl+yjTg/hJamHK0cRuYMa5l0xUewCD0Sy73aBU2Pec9Z06P844dsEIr1vYxFu
hnHyIqQwOF1Xm65QO6BvVJJdWTVDxWOqRDqMo3/QH42eM/g1fl7sOPOSnJrnhzSnfaAsw1UsiGUK
83yMnqlB7kOSaiAaJ17uLn7AaGOKGgre2jX0Hp9XfJdBA0wR91RiNf74oul5Fe+z87aW724H6B0J
gL8CChnPKBz+1idLp0feKsQkw8N4+GUBaGXAZE02NgNgwJuE99JN5Xrp1WedO2YSlJVM/u0g4P6v
8h8Qnbrz36uo9M7e0y20fZca8dfvwNKi3PCmrGs7hUX8xeBX37D+xEhK/WXFAVnrD95AT1py9TkA
f7o5gZ2EdTMn7B0HUnXarsSaoMjpUmGT5DsYcJeScrKFXnJvn7e3xjNtQS6W6LYdDlWS0CAw/Sk/
j9p3d8ZUOXcClRLhYQJ72TJUPwIxmG41Z24fnmYqIoiXMrlSCFcTw106KbQCxccBAXacuB67mKE0
yKtgbpSjZ6rWLedglS/N534QV0StEFOARzhgIeQL1Z99mwA+4FUxkxXbulmALBSAyfJgp9cw48Ri
GIEn3ftfGSNqZ/evWVR/gZ6seOjNDV3puZ64pXN/y+3W7bsvgIlAlXkQqX5E8F1APFA4ymqKxJV0
mOK8cKXiXQFL84r9ZuM4kTGilyB1SHZYB8qRAjdwGN+2c5IFnZScnUKljI9NC/4cpCwnrBLzhMuu
1NfV0i2xITi6FjO31g6wyNezUS0Bs8L8XRowJhHEfxIIuKPa4t2QOMFIop3QOjBokt5dsKPftquO
XS2Twc7sImoDz2sDVulbgQUfuCGoX09H5fwExuGyP0/amvByG5RIAGVGHihJ81g3vOC3NirbxXpY
BTKBFhsm856kOXle87VZeBc/HKsBJ2yavsVYSZErsmNg4Q4fHvSbQsk+3XPYWmHS7hXHECaM0ShT
OZIN1EEazDaTGOTtSfwk0p/0rgfmTAXCHp3KvhrtiNyRKxjthbCJ1M/9EeaE5JupG6gbgb+Ef/Ui
SaSBu05Aj/K4P3CNKsOuzOFJPwxzibh+YZq7CalwnE3/FEDWhUngA6QVAkZIiXBhMQzA2ZF4kdyh
SRzPs5nn2O+1f126Ow==
`protect end_protected
