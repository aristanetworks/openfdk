--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
XMyfYR9C2ItkSsG9Pdi4vDtf//wHPwAiQvnhLDJlk4NjqyyToI3EqKqHhw6eORUrCgWLdBTQs/nT
DW8+BKW2VNV5IIJ9wFX5n4uk6LEAgl90QkNnr2bHxFQ892iahlT90VtCrDW1HwJFCO6Ya1sInJxU
gUnynEr0t7V1yaiTPAfRPG5HWYrdNuUr1k9JGMSv+jxQhCzi9Sl+c6iM9odqBgfywaH+N081W2eF
p0Gd12U2XFlgdKZQcRiYtlV4w1muR0bPcAW1OaiGASagCOx7kGvK5EBW9x0tGu0mygy+TupdZB3O
QhJHoZaRYRwgpagEay7kIq46kSEgt1CwLJ7QDQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="dXatfWaUFogeCk90Bz2xYWfQbYVegqlvwG22qszq0xc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
jf3OluBMZJXTvE6d3TjzcaDWpVfkgH4pd7fDDLo/ZtB0lKHXBp37dwv4EDJBwFDwGAb9s3/78M+3
jlapfSFzIKU6RfqTUijLiX0XEcMCm6rMuSPjObX12xn1ZCMtAmEcDwAKe1hROqMQZQW15zvEzO5x
8hUbYJYPSUpEd+z4uCbPffsJLrI4gXnWhkH/dvCwUWk65pJGhIqASaH+4mDAQPZHls5NhxOAhfU9
jST9RcNLNUOZf6kN9TvOZJh7X5zYvOwmAlX8HgSb4ZGw3NzCpqgnt+1QtlTcmoNsdBX97L3wmWvF
3Qdnf1JvhZfGH1QRhc71I1V9V0/jDqNd3S5MGA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="aaw1BzJEe8LunHsoeI4VezbYEbgdCIxlWFhzt8lv/7s="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14320)
`protect data_block
njRZmcZCJwtqznASR4dt6pu9n8o/supLBCgDMu9hcFaQS1zNq6czMD/Yj23oi8AH8Bl0Ufy+1wNW
83zZHFMvL3UiQlKj7DQZE+wsXtwOhDxxtFGCMszJI0ffYD6WodMeaDeLqdXNkTGZwBXEkn/mmfqi
ctS8TG2qhHEdiX3pjg2DoYqkGMDE0RuBI3KzDzB6yVdCygRz6uLu6fEdtwcqPuKDRnMZgFwZK3XT
ZgOxJUkX9x/5Hgl6FAMGD5gqcwqILbaqNL2I3GFzrStFKGpWMN9UPe6AAjqw2BtB3WLM+t17IJPS
G94lAYFDmjM+fBZ5oX9FZk1q4hRDHbR+pwm3OCCn6a7d4TbnGJ6R80Dty1fif5jAbe4VKk0q+tJ1
ekdQ+mdk+1Ack2+5/EzJsOgLTWFt6f4gMvy6D45uM3+xg+/7DveusSL2GbClYmGkpm2ywgC0XOQN
4LWYt6WmT7k8Zf7b22olwZ6MBeXX6kqeNJsCIEFBY9TGgcXc5HWohPAj24vQKiItYJXe6xE0CZos
g4sW8YH+G3/RaE+E0tCeJLdfVFPX+GMKJE7OB7yA6TZbvIja0jgFR3MACbqmghc7xtPi4D54R6W2
ELc44sdBgMnqap4EOxu3QP2lOOPe1a5esTbx4vk9KseyRN+Y9FE6Tu85zSRSuE+wpBUDlvm/uo7o
9dK/w9CW6Jkp6G4yP1DKMeOsWWQydGUaxQrfghHEwauVkKNINqXst4FJhaBPzlS2+aSbVtR+8WqF
kYEmw8yXv7vB7QXlQSFLxsMc4L0viLnsX6XpKAaYUfeKRn+Wyr/IoeaPYyJiZCAS7Tz537P8eVKD
pGkp2CAiO4/64Ih3BJt+vIE8NhkxlKSceyuRGVqnkwHitvJCTPJivl0WWUsRVynEWIS6Dvm5RPVV
dG/nbqWw4W4UkiNZE6CJvs/T7JegEiYXilwxd8RIkZAdKCN4CIUGPc6YMcY2UZJEctgznQbyH2Dx
64aR4jL9cZjfm7HJApOq6KK2B1MXh9y1zRoXS6E2ojKl8oFbRWSoMbJW2RPgzBQCNPU8erqvxaxV
LLvA4SUzq18ViwXcw9NjgXTuPEhrE5EiOnvuRTKSvfD8mgrM/DTHoGE2QOYj0Xo2bcOQ+xxKOAj6
mnOczUOFjGucHYVwqem1V5xMexW1svmnuhQ1m1csD5bukaEFMhn75P9QVbuHLqGSw+Mulod2WUMk
geQFtOil4o2N9xC6K3F7lSc4CO1Snze3OSp4/rH/1slqWXhmrgbJPwH5Ul29GRE+MTEBU7OZAkr+
/G4ttu6k1WZMODPfGZ//8GPwaMBHiPyqDaubWE6p1rWQ5BOQTUmMltYUGNT3nfsW6VnVVs6LjPXF
MFYwHJnBc8dw+Lsrc8ZTMPnzEKqHlEza1ysdNrILKtQ4BhUsZN9darZ627pNQ+PahyspbyExnzgr
/UqhDOsGecuWfX1x+kZtnjLW+tFyrZSJMd6+lPBMSZjtg/thBsq8rnINkjV4uDNPEEl9Fy47FUDb
iE8l//nvqq9ECorYKVhjzZlnp44Fw684CRWxl4Hu44hRCGoZByu2mMsMuP6aovQWtAAOS0s+fuBr
+KCGZgZRuSCTc86/3M0b5dpcN8+uucE3FN9VLJoMXCPb/UE7Hk6IG7Mu6fNOkCUISTuzEDHJ3J0e
WzqmF+rf922ahnYs/lsI33GNxcZElkpTlK0c3RZQ5Rrol2u4UNTZp2hsbydcRYltll4NoTdZV0dg
XPHT4x5klsYjtbre++NCUb7Kz9xsA00nBfq8YyjrdD4gZm3zA9c1D7lWk7xcHEUWVsw5XwL3k++L
vMcqKUQaxpG5i97Ql1wriF/DYEaqqisYic2mKqxqIiJmgUpH4FwK9Aul2tKOK/BnCOG2GoWlspgV
LgDGI+wxYtgYpWq/kNr5OYu/4EXYacEwPnRGzPJF5z7rSTgGunbnDBmJFm7t/UXLwA5y96Go6/d/
WPogLzAvm1tOCvFLz8X5BX0RXNfwXzsJqxYDAOgM2bEcv9r0sLdc0VZEsjYkumYEBDkKftOZ6b5Y
5/8U3W1Iz1jkBWGmvfBDGqcE77Bdamr9T/p06hEs32f+rtDffnweMaFcgg1hWTG3MkMr/patI4Sn
j4flfBaN+FeksZJbfcA5uUP8vG4hMj3rOq1gSkDobrDBrmXz/fYORnWzQmiHXCYKjk+dzMSMfp2e
x1/h+C39IzUtAo6Y2r6ksJCCR8Sz2DqrCeRpXET1TsyRnpx3p7anfG2E9+8lTXUGZ4TQTZvce0lW
J1m5LMliVaDtMNMMmVq24kliewzw86FfAivfxIwmwa3OeJV56B2U/4KivVPwY15PcVXtRfjFRh1o
1WzefsFOdfkmxU3Ck7yIIkPCwd5c17B3vp10PfkTNy8/7m+PoTgleRNh734m3JSDlG5X2AxQboe9
7Xo/ykCxtj8CWlHsiJ0uCVlNRzcj10hjyIIeq3rEstTVnGwMPu6Y9p2ZxStkNLK3wRU4wghtlm+7
qj80lpxAV/azQmcBS9I+LJDCpqWpmcJSYk0ndwvChnFHk33D+UiPb2rb5EYlWi5vemDz53xrBAru
nCDfoZ29mCV5qx2qk4x/iDrAiQDcDJqrMZ1d1uD8MSngH5yaiPHVCiMNhwtGNrW7vGFM9r++GWUI
v3noJp+OY6HkSj4+92kvj749yCKXLfpzYw/KNN+bVMjh2iUneDENaYpf7+bxzsjLUeUQgxfkjFo3
wSeGE7LRtYreW2e1+wMKYa/nS7azgnct42h1IiOdWni0NBO3R5v1V7iHyNcsEktpmFmC7Ao5W/ca
e8RgvINZubIlcX7ZtLdBAty61zQrmrsY2L5d4cZRJaiTya94GDRRDc/c21kcKyOqQ+Q1RlVmnZoZ
Za2xbkC+kTkKR3Ty2wHa3Ktt0wjsyH4FVtej9tz85/G8Tjbmrwq4k6jpPP7sy0BZSVD2URJpBBd+
tlxvL/lTSUD20EkFZTYj5c5R4/hsGPCNU3AtA3BgpsxmzwbBorrkpLGSqFMuEUDc3ziuKyIE9DOp
EOfGZh42vGZ0DtiZEtuA0vPJ3qzGLsDvhKCq9dmQKfbz6EPc6H1SIVBjUQErBIdRU7lTGuqG8U0k
xLcQ4KuCfTE2xwL/y6vnI2G9In5NrtnYEbmvoqD6oa54b1blGMoFwat4He+nvLWCLxa424JYB7fP
qLdh4EdsJuVm9+bfJYAlGbNlGtA6k/mRCmX7WfEqNxPJmZEkWYhd9QTxfg2eky2KM2iuub5tB+Fo
oaGLva/XOOgvsCi5ITRPcpv6BvrXKWXxKOxA1LSPld7Y/e+S3/gbxnUYFD2ouXNXHZCwwQ37PvpG
aZ8Tbfi3B3UB8CSH44XX2xLOGC8TZ4gpiLWyOqBRSqAFZtdXgRhe1HRlmcCXIFQm2Q297nKTm6uT
gtGBlpZTzHU9PsUkn0BurPHxTDfvo5t6gZhqqp8jxniChF94wmtdbVK5DDcL74dAUPWVqpNXbxA4
MA1J9nDO/xRJ1y36P1SMxfi0Oikd+78H2fq/nmz8OkhPzv+UGyQxrUWQXtk7ywb549wxvFolqTUJ
Ol1d9h8yAcWAFAxF16610FyA1kaze4UwYmS3XZQRD2fvqpmxurlY9cYi7t02XX6Kl/41ps5kzeAV
j7L6aXdM5w/f0gYRZxO4tQh+r1D50CaWOj6iOBVmopTqbVDkfSkuAuJ9oYnkZB1PNO1UWPMogfDQ
dH8S9IXJQagbTMXXcpyUkQt4vp5Q24pM2Z7Gf/g+o71hF96gIpZ4+V/8RWd7jfEtLsXUmIqTqYOc
aXULIIzQFTwi9Knkw7cpwfzTwv7a9UpF0FiXxVfdM4QoT2hVGCglOnGipcYTzWo9U7yrs1c2EjRx
8BHM2wSQqcCtGwNe1IMNPPW4h41u3+4jBWhq1ZAc/G2q1nWtdX94+P8mZZjM1R26BkVD84Bnu1Oy
figmMCrz6P/y0GGIHT0eog34lEHmm2YRMXIg6MlSonmZAKD74O/cCh4iPALumJlm+yDz/a8q1xAo
GYJ8H5363kXm+qGCJm079eRrmCpK5/KLnn++dkAR5dIWjqszUr4o+xmAdT1xoGI0D+CS/tRRRmJW
GNrhX5oXnetMFn/zXUQP173wkBCNWl+hbJFpa/5e9b1fTn0chhhLS9mzHrbLrs+8BcuW4R/6o6eb
DICoAHI+JiPchv4P5RyMX3A3hIu5IsG638uAjrG5Ozp1L+b1nk+WxhrGqzjPNxEXczDwR3iKCtqM
qxfFGkVvwlHSt9/i0mtGbudqT7P1cC6LdKOwTu1BrrQLJlBsgrtKdv8gAv2cGjJPqwf+WyLTaB0U
0UYlMYK3zJD8wRmUu2WRoOIhXHhhT+Ks9sSPuaoFn+P7XEs7U1V7Dl74AmCdX2te2FIEZdm7AjUc
uPGgYerYwkmKdhfMvPNzMnevoTdB8nTClHsS+PXNFZiKN0owDA/9B10fasW5FQKlFle+P5tzg8OS
mlO8UevCqKFajWCuWeVMXQzHc2Dy1UrkjIzwQuafQqGaBWLMPvZpJA0uP77UwOR8aHhhGvtioxVw
k6VwzufFOkNZiFQWVQhFwhEza0EvJL/4LDv5Lub+sTRt9AE/7jaRwWqcrIDx1HzutulfVzXStD9b
ZjLwy3S9vtXAZD2NEs0tosGUKmcMY/FyHaz8zd/gxppeKDug4JttnzOruz55ZITmNrZ1wdjrq/la
W7mNSlVmkaUF0pnujoUFn1HxhzGNFwZM9z/tdlEaxJUOH6qMGh17LRpZdEUzGOePmI++WbZ+/Gft
uAqq7jtiW6qVLW8ruLiYs5jgNCdQvrd9tm8PODyW+a3NddoDnSHQ8piBk2/v37WsSO1DAnzVibpW
USBWsfuBFBt85QctQEI7daNf92uGJLOb/t77bpPWsNNUEkZn2NE32pQl6WX0SoDKeFiSwVx5nlMM
Hki0H8jFuHVqADuFZZFKKTiVCfcRDJHEQsz6D2OgmDv+4466I0R6wvn7RJV3JGfbZ5bl7WeGt4Km
Kdc3u5AVcJTjFsR+WDFEFaO7ITZU8CkdSUl9b8HHCateYjt9yQIi8VyIxAbSZbL8KWcjazDmVU4O
FymT8kboBmz3OBJ21xroNwCZytpTA4JTRwXyHJYlxbeVYwl9PjHQFzPFwupWdeUQhd+Azx83JmyO
JZnQJXD8Yx6cVw/d9jlL0LF8X14GkOC6Q18/RLdCE4vfq7+BWYh1jjL7CGhM70EtAaLfYkIRiUlH
mGDIYKUCynK84cRicAqZOhpxQW7bAhLgcf4cqCSb6D3Rt9jE5ZV6mehL4v0jBjeMWi8lGBBeQy5v
bQZuu3K1rDq2RkeKhNBjxyHxCs6uYEeHl8+LeiKE+EKa21P/fSpaNT2FBK1WSrQvY0MezXXwJjsG
Cbk0sStQuBQBhPdAWfelXEByCJTaOx7hbYECT4gQSEdaYLJsXj+Ivq3DRqa/cTslDB66LVcOcvQW
0qg6X2e7/R7XBp+tel+eV1YfTCbXmoEE1KieXMPtwXBo9AkVZraSeqQ/rd8p8HeW/YorYrUz47ZD
TGm5xP7rMynNwYvZV9bxaKmUhsT5EiWWDUWrAfbJTgGARJoqMOgYl5dLQW9DGpL5vmRSoM/mkC8t
SZ6+V8wZbBBZaJ12CmdwA8/Gvn3e/il6rdvI/i1aCcDgSFHZj7t6+uW0RgT9fDa9dXXn6oFjCZaE
/ZPMReATzck8DfE3SCuPtwtqz5UHCbU10XK5wl8YP2sTsdRSzL8/UkeMtA3XEw1OUMjq/TFSkYrL
DytTsV1HJIS/15pOZPabARpcea8Um4sa2vGz6N7NW+mrrdObhp/r9tFv0MKgPbUb0dXq20iUVmJE
5mlLyi1gGQ7+/iQXA2rYyPO5Hao+QuJq7ooY3uUZ9cDNBwE9XOgSuHf5YMHkygWFoQkjp6bJcrKC
0ojuONIGR28kn9LMIyS5XKRofuN5XEDO53oVVroMYI0jCwQmhNJnwsv4UxZ23wboB3j4KujE/R7t
WOu8ZlTm4HIkMIYbGgVmdmAqj/SsFqiKNk6gV1d20U5zBhkJdcZzxyZWkg0NWHAhGjBSANuh4KBN
mlf7CYvQ27ynYki7fUP6FJPhyLS4Q5Ymnh17MsACopIU47zfKpx36ygyncpoBgCtCAJ+3oRkwL2I
incdRDSOt1D2j6NQOibrMGSbXGmhOzumZ/OinbTbKXM/Xl3l4/aI5i+fF7MLxf18muzcV4gWOYiH
S8OR+K4wrqIjjalUY8wvpDB8ynxk4Aars7b3FrdPaTPrERxAk7n6YiLFsZcUfbjNxkSTzHD7UpMZ
n7GyW3wBQ5JXxz81sDqahgpE+629Z6iJIGJVimoPe8W2D+PgqY/DlSx5vS4Zu3LlRBbNUu4dkeYr
lENTFIg4hERiLc9KzXT3zhZLaSUq1qyETxVfK5ZvN87LgttCLH0ei4HXRFu7LnGV0M9+RT1wYY+h
EnbgtwoZnIdixOtB8K4x8dBc328H01y2uT55MjHJzCvEQDG5dvIC6DnkpXdrNNh2xXRwSFVHaTle
Evx1v4vYD/ME6ZBkSEJiw1J25Tco+idMFdDI02d3N5HUIbZb3xGEdLCM0T1nIp43ANvgFvVA6Uyr
OVnyzD1z+/jhScEDgHNPXXMr2Upr/MfSYPqxLqYzdny6hWq2TT9JXAKZ+nERH/sP9A8p7O7f8q6r
feNN0KpvR8nI2VTro5K0O0sFiaAurLRDDugNxALQcfEr4cZiqWuSujm+0wl2AjCcatGjYD4ecc22
O/HbhLPRwS2Ey7qSNxxBnq01YQ17EGpiwQFjLEK5p7eTK7WNQr/wdgOsslBgJrBlv7tnTrq/GTZa
qqlHrF8BMqvETOgIW9haEUSsasRMPmvrSNPRv8RIwccWNTyn4GPO4OQQE3NcukOl/hNOYSAcDh42
ps9dYYhvdFA7DtSnYA/+BXyyQxCiYCg51/Xr/qpWU9CuflxulzVit8qIyS/dqSh2r2s2a2dIJD+1
k98mxqqq6ymz7yQCXdQDNGudM9XsQ/RRCbUrrziwZ2l/X99gEYG9kVZCLUXwVteYrOb6mdnOtWD5
bg6v3QedIFzJIKJPhx0DxEY9dzSQlle/ZrI7/DuXLTBy1KZDse0sXHEZLosubW0cSvrIsWEWdjpY
91DxE/IvPiz1IoFM/lZj7ACHhRjC8gLlevkNn+7Y7kp+IpI5+E8Ok8k9VhSbsugyzN2I/gRdf6Aw
WwWRhMgVAEzcwTCAScH8F6LQ3KtVjSkT/Qnlvcx+nV1M5B4opxQAaP3t7YPYZsH5x2DAiz1H+nDh
z7lU3rldRb5Q/D77Qpn7UO3JC5RdmXv3cegQU6f030Cg7bcmpJpx31s6ubIl3AxPgC73RgIcKeWv
YTySmNrEPtglRHf6DrQ4pgsZaDz1rdu1tYLWz6ptBuhVUsxYgmA3g5BDYwUTu01UMLBRClvT7XSy
APzg1p83Ym80WMnA0qPoq0Gfzu6qI5iN74p7AWPVLf0y2B+EU1DMjsJwO62RxqDquRQl+LA8Ltkk
jbJPZuANehT6MR0x2T+WmidJY4MOyY4eE5qleKWWe2KOMGBN3OKwdi/TFrd5ZQFBJQg/P6LLGXAP
H92GgGH137vSEz4bRLzzrZ3rXlWc3BiboUnHfu/C2Qzc6XBRtjVlOjKBzmjSXhIGtvZdSZPf0uqG
nfWnbZ3gOwY6FgLhL2v9Jsjcqsg8Q1ijLI1uDvMwKpD7OsdcQiLtZ+OY+xHwa/S1d7vnNPm0FYWb
MffoqjB0+CjXxWuYAt7V/5fHQCfMlfsLmFbp8EWpD7Bn0/pXofsl1vIobDPFZQKs+pZ+DzArfqmg
+CJRAyyNjbkVfgAvbemcX3w7YIXu4uwsUSYd/A5elWfIYw3PY4wb4tpLV4uAwBx3BUMzrFW3hmCl
48UnGB3RTa6j2dI9/jPFQpLSRbU9NMqyNODCeZ7mPLCGVCum3GDcsD1pD8AbtoaxY8UKF4OxOqWR
Yv//5w34JzAXucMEmXJ+mTDj5pjbI1GN7MvRJLvA/dkXJWHWepQe9Jo7zfvxk18Fn+VXBdkFzuep
AOJknv6hHmq7Z57U1FhpwXvGfDsl1xsS+ZMZTG4JGM3k2g674JlAu1pnM1p0yUQEgcPLrUfLvWEm
O2QV9fbqwxgGNY9hyDtkNKyQW1hqNhuytnoFnS4pEpIzcE6/xfEyvJ2ZFtkbzVjSm7NeVsLE/JCC
0UufszFk9is9usF5tNddL3sl+QnR1zzTBkiJNnLVtYdVCqipTbTA4OO3eZtj2iKJ/LdB51JgrBsZ
/Vke+1CK1JdL7Mvij+fmAmRfJPfiRK7APvp65UW1pRH62gpcXvTSobUWQ5OFd6TJyyb8rNVusMpF
L8jOwxGTb7bzOX/+bjtvblfKp0epYTyCnASKn9+Zww2nLHznZITtmAYsZKuhtS1dpHqS4krgLcNO
4MEZCA4ojjsJi4nUJ9/dp/f34ZvIcx4lFveQfwQJZ8/b0ogW/qQuvW8E/9CyPxEhToEPB1zEFsn+
jGUc3htV08KRJimHh5umjDyvQ8AS2KvVvUM7eybQj2oYh4Zh/DZrjA3LUqzrKpyzUMn7wxDAbNzS
o+YkrIOfzcSJXZuc7GnV/UYWKuy8NVWnmIU2Ak3xFCL7ola6sBS3qUqlX4bsVxaVa2Fvbkbz8BlE
L7Gu6y22gwunbt8AF9seHbL/HBNkpVSlMpJMO3AHdGQxgU4fdg6uNfJW81uZUZvUG3IIBWMKnWgd
fUF6PLr2lO5WWfB7kmfSQcPA19oBszt41JmNe8SSVw8h775okAgHTMUpiHSyFua49hyDJfoMaGFv
hkG6AIbOsWXBXVce9qKIcbsWZAfi62kDHCXWYujDKIi8bxowVImJwSFcRcMMsEwJn0uC6f5KBL8/
8k0fEv6waIza69T2CTP2dQWmAQtWcZvDXOIKHfPYoms1zekW8M/c69ayTxZaCX+jsLnzSmxzL9dT
aZ3dGIeQao8HrCvjQSnMdFywjuirHWMs75qUQqBaICSEruo3aKicELwdtzEZeSNUjb34sP1Wi2mh
ZB5lKa+g7+QfGdHJTfJOutUjeW9La8juPQAfvmiVzhbYD+Z8IC6SvDZWjEL26FNuYwXuGKsdnF/L
A5myFc0xInFxKlA3pzTlNKkAC/ZNlFr2cIxFTHU2sZcs1KP1WbtNzw7KSrB0zHg+bBCAAaAqc2KJ
xMZ/7ZQXSvIqE5xJ1XJbxPJEL5lOK7r05l2GpbxnchDB/86+MjTOsJISTsj9sAhRCJyg0rVIyo+a
09gL7V98LdmZBEZM7mWm8f9gVjw0pq4JZT2pw2cLeyVhbp4PrErcXRJioXiu5efyIO/KLot62Erc
7CUr9WkxHAuS8BKJXVbus8d4W+aMaFzJSk5QwRnqrmvSNB4XQ4v8H3NSrM3qCrPU/ox/wJ4iXOSl
Z36GBcs7E5w7hzmWLOAeG3w3QLuMqLR7HeniGnoUnL0qs3mXDfj0G2T53hpGT12UxZv3sYOn+CfO
ezsQAfBP7ZTtbppOwvoqc1Yw1ZYgvaUKjfYoXgqEFT/VCe8w/AEjlDj3V1NlD96bad2JUJQuTTel
7OQ1CC9/mYT4jOIjurk+6z5QCh8clYYI0zd2Elg6lNSqY7O0eeSP7SAiCtXYt4sSaxLderahpsvB
4cxFDV9RiMchMK+KmxLKFDb/Axx+tCRcKy4bG3a76h7thcpuL/rs46eIRk9Pn0r+6plZfInpItQu
0dCMdT+4nxerpWatJMU5n/uWG/hoEWNKPwqNfrdfJUmWFvKDHzW3ZJnU+kYNxvuDZW1G3A5l+DUk
KqBaE6vfppHh/RLySwA/4J7vKpc0QXBRFNOcyhU54UgNvP/f8saBSiXOmERuqZ4AP1S8o+febQGF
ai/BGgKsjRHt49NFIfOSkRi8d+LJPvh8VYJ6IwzK5sgH83zv4WH22YnqPW1P0PFTYZYFNmonTYbS
Ue8fYKDHV0TkrtUwjxYUr4uX59/o1BpgaWEyvpeso+/LfCqspTue2EuXA8CMTcxVqaS91dCVYHQA
Jq99TBjQDWMel+qTmff1zDvVHG3EdyEP+ctSRxyq1bSFPQ1z21tPUDyHnCyHzciqTbY7XhSkBHlj
MtPdmHHJ8RbM1vTA2uQ6y6Hj5YDDaygDD54Bv6QE9yPN3BiYFMjhgPOMFhF8oYPGv9RRY/VZ+pM8
Pk+aLMDNyZ55ejn4M/TUZ2ch2mwaU3aTNzYv6JjfKSO4ymHnjbY5Tc0Pi+Ek7eMd3BrlcF91iQym
LOYmasBheFEUv+3KA9SAamYZly58MXPchoyW8gLht/eS4YFijAUqxUD15p23WRWsiDxLsfu+N6t2
LmtYP9u/A+5Pv4runNo3JWjRWZmCSYpcGUiDgE1mkr+QqGJ9V267QfbSch1A4jCWHPe0hWjP7jyY
6Y4JLts6f1agAxz4l/KK2ZHPruEuxyWW4lBsHNmVcUvlAAz9YOw1KHh0W58hH+9D+/Xxks4PAXEM
3ux7Rn9tQI2PyorxKUEhC8r05opct4/RiONf/LYQPl5PZ9qv7K2aMwikN4eH+L0+5Ku/VeYypvfB
cKInFbNBSDnHUDVj/6fdWktwyclFt8WE0DQTefkzamVEfeqoyM6aJeDVTuvj+wO4BpST1e3I9GGg
fGt/O7g3EuFrIWZJY9ELHElmKQgSG2jsDjIDnh57vUVFw3C4O3oi574L4UmMaxgWWqMKJZ2zgBNo
2/DimYRvpgV70xLG7ysQz6aqRfJDEU4lNIMlxaKtryFJsSasDrNL0ZxC0qloKfZRCU8lseItmz/i
fUZ/UYaxOzQZ30xGJX8sZPmEqBKkvZFKPO1bvoHUH1g2Rw81zpicaXFiOF9CYihmHEi5XCvrt/yM
f7xWn3b5EcojrHjoCy03aiWSxCHSqlvcogSehjhAnF8ZM/boeGHz7N8YtXWLXT4A1/eb0iy/TptR
tk3Lcv8FLyeocJ6ASOOV9HZdiwC/2WjbfVMFQu9vVyI+sJd0WDJpuByj6ap66MpJB4SDFBMRXG8S
F7xk/iuObtwpXX4+EWurgYRskifVpVkz4bUxl3AIuGT51UxPXzfldFZKpjDjWeRQhPOuZ+T1d52i
8tfgyrOns9I0wmOnsc7YWubk0XmZp5v7wdTOVq8tThHfB1/hoKOtBhMW+xm1u72de/bClVViYBv+
5rHUMpLjpc1RfUKQz1gwjpFCpk5vYwboiLbbHalWpLdXeoJnZmixOkirrCkiAnW3CWm12LpPAMaj
esbWRbn0mexBdeCfbRkda5EQ0Rbgvjcc/RdDJLB2MnbX9rB5DQ74rMpC10a66ErgCN1UV2omXst4
Wg0MwY64mezqC1o60C73cUpZoHsGILMtJgs7j+NbrcplqVvz2RetSNmKra+Q2csJfvrW4tutmAar
aVI9o74O1o+aymFLi/feZ+c6QN1wV6744Mjo4AQTSu4dtUHTy3dN1dqSyAak88Fno/JCHSwkxDIi
aUA0r+l7p+9UlcmvlDo0R6KBeaXLnU3OQfm1BKorEXgeduJF2YfMw1dMiT8EmmHWZJTVT8aLL9VB
Hn9xdjKZpbOdsvHppb/ZZI9q+AvEt2/oC+oXdj4Sy5AfJPvQUvHlNzJmvmWz6yoUQccmArVCdXb2
MNwdBambsd5yZIyYGfTqr9syTpZfHXvP1MPpMHLRYEO98xknHPurRdluGnJtibN1eVLhBqKkKz9Z
ICAVzscJ4islE518eV4pb0bpKy+KEMQ0+Ngn9qo/4cGLT8RzD2xG1kyGa0n2O8N1qVJ/oUeMTfeH
APk0emT0eFBYOf4wns85JWJq3sbQHXgHctWlLwZ+bTTtdX6URa2FHxypf3drUNtpl6AbVgqlIqF/
ZAdaxZ8ldoeismdgpbUHbZH+PkEySYQACKrnzh1zdtJ+9nCTOvIUTEQR04BrOBhA2NoSThYQZqoi
vCFvS6j9hHU3T75kEf/++oQ3KhXLrCKPWbrAJe8dp/6F3RMNhUakZYL9Y38SmEw4F4cbVd+Lr8ho
GXqOa8LoK1eBeEjosIbcgtbgHXsZBRaV4zR+7mCJdqHsdY67LvJ8qobV2ENitDHL9MqSdGJx8Ios
etYd6H7ovHENL2VePIlwDgaTUmtnLqxpLf9uP/Jmu9jDgVgiUAIornTfpZ9Lf3s8NYLOXWQ8lcMv
4O7F42kLPzgv+Ob69x+M7KMUA1x7YMkMsTBtxNw7NANCl/++lDLtUzH1U2llpOkb/9c6z4QjcpGw
4RwcXRERzhuKxm7+ccHY1oZBLRvzcYQFOWGHvQ75tnplx8lNQWy6EH5FVhxRuFoWElUWMUgBBmvZ
PEDlnBTdwCCGOCg/tHq41Gk7/Xo0O5GF7h8+9lM7tC9a05ui1IFlI+bPmzPKWy2STYFKgPeedNIe
SohMWZltnNwdw67fM2Zkx3OkxNGbG2UPqbMPSljvAR+tDk/P74Y1vJcgLUlszOqHl4lVUn9Byo4V
O0Vzp0hvD3uYPOhzAdEWlWlv/0mOAh9Ehb8+6e8dqDmSvjgSgcgn8myn4Fu7uVWrffkSEpj6h/hi
UHRjqCytj3nkA6wa4KSWPsGm887Q+povVAqv+UCbsQKLoqsqlNtG2wkFt3CoqjQTqIG7XZVEPIrZ
crkipIrZkzY13fIlg/Jmk0rduAysvA/wbW5nEz3VsWwweA7rXb0D9zsvetC+aRw25ih/49rWwPgl
WtACNBPa62obR6WLjH88pnwrBpPvDEB+JP8Pyn0DUA8WXAeASW2yDBCvkQU/WYE43WXeDU0WMW98
1+3jEsIjJfCLN0BIGKoG4m0dpir8z9fJnI2EDTuAdkSaBNf5HIehmYTMJmTaMBvRgxKbRyNeixw9
D0N2FkF+iBMqximRZs9jVojEBs2051snAGHSLEXK6OoupSR88Nf60zkcGGegyNtbOuEzQ/LtJ8oe
EhldaXsa0rI8V4bZ3cU3ZqVaThbMKYuHqIOeqH7joMf2xP5jQroi/kdOlb2wDgqBWCQXczLYLW1T
iKg0uVFQUm8wqn5G+iTV8Hhe9Vo/JrvGCPYYnmBCSzXVEbaOxVPjrk16RTr1yB554uQq8AYMqSq+
QRaI6njxfHEhSguYSSa+loukEmf31zpV3L3Icuxbl8VtI3SXxMzm2Om9kuXzoQEolINq88p8RMjr
u3XypUTGebYn2dUmBKDHQJyc7CFBYLB5kzHUVeUwN2Knc7VBgGnz06iE83HDsSM4zk7Us/msBEzn
b7MHJL+6a/6nrUlhM95jERiNEI855U7EVkziDfk8EInS8P6bDbeejbqSa/O62K6/gm5D7WLZ/MZZ
yYWX1t41S62WMi2MMEaftW4aw6RVpb+EdhPjbDqYeYYOVTfZY7aGspfYyoFM6sFUggS+iAgx5hzU
pmzBQ3gPGVQ4LJV5oNy7aWDprkHMycLL6AMRNZGHJk3setAMuDMdP6RBOzRNMZjHIQvy8PYvpMzR
5VRRGCPMGZKlMUzMzap9Y+hFdJs5+/fUPLnBF7RafMkHeI4B8OB0uys2lLII/f3MCz2T0ICLZfuw
NLl5rJ4Ao7qUHa/LqcbhzVv4GbP4nJPNSHmz3UzN1//znY+L0FXGb17W8dKrq88v1MlVMVhC/sHO
zg679eY+A9droYoUQsugMggZaCIXMa1JPD05g8X4PHWBZUlK1WhZbcPLg4LNsBg0UaPZxSaIR2xV
EXnAZ1eAj0kvSPMrM9xDk78RSqBKgmih7to/+AmY6Xh4AQWG7cL6r3FC1iLA/NwcYbzrvdX7P1gA
ulsQzNe68HGGU2/JPgf1QzBdKMNFlzqZVEsJRYIx1Mcdb3+7/hbjsmZZ8pyw7pIYVv8mn4yqEGpp
lYb8XfGmsp/QLB7evmxh05jfh5CaE/LvnujHL3W3ztYCdgS9YOc8BMBaQTdQZ35lprhajGONZOxd
QHdifFicFyvcc+pgHEB21mw/anH5kzBWAFVZrCgSTzORJFbMJufd5aiN9ufut0akXu6tFDST1pcY
c8bJdVkvrdy9Pt+s9K9dMywVVv0DiRyUoO6pz7LR3nnBxQvIfPy0qzTpSuKT33vtt285YYLmfLbm
HMj+cxXlI+3pAAp1sVkke+8Ld4mJAbCxKsovKjzUeS3W179mrzcZcCEP2OX5BkloGdvOGKekQi39
XbXxO5lP1hr2r/hdKQpjvUyD5KVYJ5QQdBvcpaaYv+N5jH1loeKuPtj28K6pxLCR34AStUf5sTvW
DysT3X7jfyfhcEwOb+Lg9zcLVEeHfgdkHN7AxGLl9gNdziaolB1OxctpY7EiEi5bgaura3Xfbouv
iQT/UrfWB/xgQ5v9kDgCNERyOMbrzqCkASUCGLR9Osv0O8ojaudMFd/hnUGG9AtiY6sDKX5ROyut
dmSUu3AEAuq3xNN7gkBIS8wYW+UPNTr5A3nC5Xfcl7I5zDm2RWAHm+4Eenaq3Bu8WxHNSGjNPgQq
rbFm4J0vaI6kIKMuAqXOTSu2NpiwvZcOs2I7mO6gDmSPwY3oOfnYMqJSD2zY8BqZ8PzyeMkSDUJZ
F50xIyRJDsatQ/a77QyAaHE0fIatbmynel0jxVOFPtZTj59pKiX0Na8cwQZQDW1inLe5pqfPP038
ayjuYEExg++/nQVi4QZaXr/6ypS+iXbHpD82bPYOInGRVP87Yet9+bR+N0ReI2qm5e0eqlb9Tp3D
n/iBw6nVs/yZke4hgTFgKiTI0OeO8mTGSdXRZ9Q55ks01YTGK4FN5naB+RB1ONCmNsFWohT3YdV5
xRD/KRRmkqlrekblJGRklNl/qrHu+8ROss2gjYTYrCRDHupJbnhhKd6J5rxvLyNSHJtJ64KUd+Cc
Lp2+eTPawDOIngd73w64i68sy8Otaj3ti/76ReXQSrOxTyQmvPTbo+JuCiuDtrDS2AajLqZEXKpR
EesDQMNwGtLFysqHFI4BrbUtq/KCtLa+O/fPeI+Xp0Z2fqU00qaZ0iKvYz3FQZXt19ggsE9w3u6o
hiDIToCuWToQYCWesb0Ugg/HHxItMy5lqTjTXfh5OaltMekrg3T+arwN1B0130ciZj9UHKnkuGUt
Wk1W5tmkrrhafIQQI1XI6YQvfnwJwrXs/MsAhkZYyvckQIarxGF2HQi1i9Utzyt1D3FvxPOv0Uxc
KMyv2Wir3yl5WbjTZ//TySWOUFkSMFwORYAqYspRoWotjmffTGvgrAZxRyx89T57Fgt454MScrCm
QPp85rV/2GrcXpoK40UnhYo/tCsP7UP5rwSgROiMy+gWWw2jpSmLEEIii3Sr4yLRsrlGdynZS98d
Lvrhj5Rg4wpbX5/V2QRYMQx/PfrtaZLvQ4oGVSmsAog2XaRfHCHLj1J4EHLOT4moFfYjR+F5xnU+
DNdqGMSLy4tpEOF5BMyNyBhORX2cN0w5V1ufxAm0Y2/+iVAqFobKjwhlhnpIqgQUgkmXdoiYo7eD
gO9U0L3yUcHoipu4QrdH50aTEr+pRoIXMXrgngysQfe4foZTkxtuVlzMgSjhTkefTHXklCg192+b
6cmaxVyQvCpfLzYRfhVYbU19rU1lC42UzLAUmQ/zCwEMg0gsaoXj2KT/Hl+8j63xkQI6i/2TuVyY
kh8P2oy0n/5Ix0zmWNMkUkAS4AjK48gjxiIqGXSgmUvyIf6Zcptwj5I912GzO/jdyYPlkKQkXGt7
TAil7+5LtQ3f25DEMooD88EMJlOrdme4BfBml4vn5k1QYb7+p2+ISVCE5QO9120toX905tbqpg8E
iArj9kQDIAYDTB3m3sXdvR66fh0JDX0QZXKixDe5cuCy4lRBi/Efmo7tYpJiW6DFOQM1etvwjeLB
1hnCIdwSmcLplicvbT9GSra/DgCxzUCEqkwuBiqnKrsT7BD98AJq9t7IYkWRLUqlsqk+gnCPIiWx
4NgktLzvv+Mu1VOomnoaRwau8wfOjAUwf6fCsvhoXtHj51tpdhoxQ2IVLhd2e+gZQZnAQ/yk6xVd
iUuuwjH+UuaFnFExTubeJMVrr5iSNiaLsX45Ui94f+idyYhMoXKpy8gOsXpNEG6KLiz9XtxMzu7v
O9zRMoEK9DabYdWovikXMKRKwRC2ZgXscZ9gwvDw0fnMR9jQxTAsdfvOORDx5crB880SioOazUD/
CcyP2VbIj70XoknXwqK5ExmDfUCXya9W4YBe3MWzmjs0U99DIbd6h2/bbLEiMUjZaoukOJ6InShq
0NQxWMGSaXjL+MKm89XVgL7AG0a1Sr1BAE7lWCP3ADUkxzXZc3HxUgtDwr0yD1z/oX/JjXKGQ1bD
nJtb6VTKHFsqQ1KldnVVUfpYOGU3bNUIlVBimzr54vS7LSKnx7e8NKAkPH739DaWN7w47m0gMHEV
iLVcD5/cMbNechuISFNt40P34HAeKjYtp2JtY2zkOSB/X9uE5AlMKXJu9QvRQtiJSTC8a2ej4mHX
r0bGwLh982kRa0D32XJTTHDVKPCMfmqJ4tzgb8hFFDMvL5vSo5VPz4WTZGdEhxHanD7wItq8zwjh
38+4TcV3DRA5WOoP572Xu2KrFj4G5iMx/LkqTA3qVi8AEipJW21r1hu0Oh5ofmSld3PWEeDcN6fY
4Ny94uEq6Du+BA50NdWZQSFMugCI5Few8xcEDtxeyWJP3KSaghjNIurTl3E65jO6/Qf6SByjzfwD
4QWmaneeqo6qJDok+PsFDlm/w9iExfUEW8hL6puCABGO6fU44yI0zBesot0BOxJaQzFLhnummnxd
9XUSYxWU5LD+SPIkcW0NUK4SpK9z6s3pwF+uutOK24w0Nhjcs1v0Ujr+3qJmHACAGnn9rksuwtqK
6mwAMHH9+Z3+PDzyr4DjDrni0qzVl38VoRWIU/88XGJ7DK9PY6Maqf6Xiz5t6AF4JOWLgynqUbfI
tXEYxrrDxE+MxaboFinmprmDUevkYmp/ZadEm8LjNHPi0+YEAkCT5zGw87chFpfOpSsWNgBreVU2
L0M6w/WptyAXUbxj4xVoAcX9ZAsQ1MIJ66f2es3/fGDlygN1SeF+TDpuWcBCIKCJT67gwPXM17Z2
KDlO/xflSUV3u23OyZwcmxuEHU0K8cgzA64jIdtL0pMWLte/s08TOlAenzx+fpMb+uuMwziZY+AJ
4v+qwo7oh3LZ7Qx7MZmprb6HM/oNA6F9ypjQVhFIhXmxSoAGuBeqp3NKaXf12CdOzSE49uinuSD7
TotQpzGvfY1S5eEhYgKAIfnh1Vp8r45nLjtJSuCsZhu7VwztJ8lBjurvbRHk1noAgzTb9oeg1buQ
2YjFB+Ivxe3hqyb3RNL66W8uM4vhsINCoucidrejnrn1yWQbPqO2dRNXLrG36eZEsRMrNDsE5Jub
g/q2BBhPfDut2cANFppjivYgqnmwfLOoieFkVrGwqkYorI+LDzOaPCYHqlwi6Zx4ER35kTT36gJp
yGhYBL0tnABE3vddqyIglmcmJeEGr9/gjr7GXc8ZENM2OCfynIjy0WxBfhX4uVcrWafYn+VS953P
USGKmfa4Kic4dzsglMGm8oyz6CCzDCwHJhy6J8ZJW+29WXlAK8bDjWYtvTzDDBWIb59cg+ZlEUYN
d6328Qr+PH7x+kKI78rzkMnF0GIbdMGLo7N+nBXCQIe/isSNgOCM25cKP0s5QAuj5rgrn2gpM3GL
JHBrBizZBkSO2GGJ6cLDekwsyScTix5sFG53s0fWzGqyYjbGMmmmrMHHN4TPWKl5JsIyma6dAJxl
hlnWvd0lqYk9HnMbTbm/BKVmOCCc8RY26i3xB9KsVq/5P4hthyx3osM8aNkjbxqE+xvT6oKqCB3J
LnueB+0Nv3HbeHXh2MDROLWxSsCbhNuBL8gs9Mk3Rsv4E1Q0HQ4WNIjlP3hA/MP2ShydPApCEuuJ
blDPh+dxPe5jiiMGd1B37Xn6kW2l+w9nNQHsFWgA1bXpE8AvsWsS46DJkP5yyc3QwklNxaSYdzit
CPcx4PqlaCxE7R4UAtRFQtDHInnheGjseyLHkNO59QnXSxMDih8K9VcJdQQOaUkShC/y6gQfBbW+
a6tSJnGJAUx/5g6MwGDWQYGZbamvnTQpKSUo5bmuB8mHs4vX1eFp7oodcwFpG4pas4Vum1syvpFw
YAOnJz8ppw+c6oHktX+kePMSG+rOrgQsPhyrDUUozH/PoOMuHhUUcaD8DbGNYMlT00FtnG+h94jL
6X8Ji7FwOFYF8QcwXMHSEcjRi3+HVM4xzq0O+/CmLU2LV+eIZ0P+7Q4B6yV47dc/KmRqPoFaXq21
STgSCYx3iDljTmatfGpQApDvEm8dtV7tOX+JGTiesfAa8UTLq9tqELTeQQox6cY/2DLzn6t007T+
1wwXWpeDsTOrcXrt8VSwiGS8/7us8wsbj08cB+JSvompQ5drXXHX2O8E9AR/Lig8gP6ottf+knso
72m8h1Z/bOBf2VhxPfESmxvZx41SMceB3i1Nv55I7K3Oa63Kp1X157+2Jt3GIh+ObHA81NQwj8ub
YaPxZ8x8XvH22bUvKSTLgoIBoBzMKUM3QZ0hPQLMQajwF4R8RWcZOSY0CMOhr+uQGXclbyeyv5ub
rDJ/DTfcQof6iy0eBI80bHtEfek2TNUYsaIlIiA3xIkKZkq+fPy2j50vNFufWwhyyj96oodpRfS9
iYWkJvhXY9Th1GcRg45AOQbl4D9tQgzx+g/555rh2OGhP62B5uWKAHPffNtRlVt/aZosrlBiNSVX
pCLqViCKe3nLWe3onI2/dQFYUGUgCU37mT1k2bwpLHf0tpQGFj9jCSUIjM5kVxNbJFEmlX9SMuHx
wi1f3B7n/1nFFXYYxggZglMec8JfYXt3/UW1Gj2K0iK4F7RZbe+P1UusME+NcfCYhraoYRtcBSDz
OOT3I+VeS8+oGKv7EaV16AASBMjKnB7CCREFUd4svBhXK+ThJ3iPj/hmXxhkN5gVy/U3s8e8UAq/
pV9Cy3LBDPvOBCltQbAMbj8czqKnIu0uglqHJ4LeC0DJRGCsYLzCXLB9GQk/tPPBsbCgUCxOnG41
p7KMIYgdbniXWZXkUsfbxf/TwQPpv80ilUAszXAGQXvZgBnaLSfWTvgHPl1nHemLlT3FuaOYPL3y
w2/wqdnST3DJQkcpyg==
`protect end_protected
