--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
SAxtzGvOOuAAVWOZXsUiCReyBBiG/7V2CnBbmUiqTfMQ6gA8ttSekqn/DsU8POwO+MwV3KCthG7l
DIlzb81x4NhXfmb7j/C0rnSfijUOsOj3G+3AOuIXLPdViEP8Z5ug0gU3pYGhp/3S5P2dVzvuwgyz
48mWQRVfPPPmL1YCvCYMcPWK0w+k4SGOX4Dl5KbBzesKBgqrrDeA/oRhMYLXk9loSCpvjuLDYTfN
zpGvSYTykq8eFFXJ3z+mMMM6j/7lXG/a6Hs7iGT4IDcBK3Vd9Z7yYff+by7ftY9J3WLh3MDxo+7F
zKGoPyALULU+l7xf7EVpoLhtQjWnjAnqFriLDw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="YptZ3PLo4ckPD9pjczScLpXdeUK/Vku699mAA/z6TZU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
QYuUsVzBZOgxy1xpQeVCD0S5ijQz06sJ/ZnHwldagg3VpNKtTBNsvWtkRgW1wRoaJIasWp5pqqYc
DXc5pKSQi79leT56QGvpXk4Rwvq6iHRujkeksTLpYDEr3fByNMrkwI9iwCcYZxJMSEBz8FL/KJpQ
hFcQjvriFbZ59wkqk7/PyI9emWoq9QvmNt9SHmzBOseezG4OnuEI1FW4dTMPAXsdDWuCucfXNLWv
+Lvbp+aVKYkSIQduOmqMhTkSswYGVHcqRmAZNz4zq/l9vuWeMpY2CoU3c4cwhpN7rxs/UaJnvMK4
lQE47rIxFVWgyDv6qtP0O6njcOuVpDrTlowsjw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="wyFMKJV9G6H5GcPDIRdcuNnRYGp+ZxhTcDzEfDlAjlQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19584)
`protect data_block
oX6b1lzbPPgXocD8tHWSa6ZZ9Ve3ZeX4kBiqnS9ZkzjU8uLGN2/bjQeWmJ/xs1CgBW8B5qwGl+3y
sDAA9vnSFvrUWznqiEQhg2wMMEjXS+0Rut5Ws/raa+FCxAMWpUeYhBfTE+AxIdzNFmuSZterYu+5
ucPjNLxzim3DUpZnGOF98h2yuU7DDDKp9+UZhhy4W/LoTVmrVzjM0NH6wbg4/iu/GEgBlauetrsT
f0E9nPKpsz1mlEc7Xi+jQSg/AgSzr+AZRRp4R0NNfiANtAZb78O20+VRiwBxf0m+kx02mVurjmEK
LOe4CvG0POBpRNHA1UwC5UPyo8Qs69SQUm3xcHx/b+5dWmRDgmPuXj0+hUgz/87UflpD03fsBPGs
+7D7/SBITDQHl/oxTVzb4X6zYON15C2mPF2MV6KysF7ob2/XEYGHrQ6HyfNgz01KXATX8cXoKF7u
+hIYoFLQWtCXuxrwukZF/uJhabl+z8B3H2C+r3vvg6WeBT7+X/i2AojaT9fxEeR4UKLkOlCuPLH3
WBWAWc0x5e7x41XBSMvRueJB4xFBfd9QXUbdka4gTJ96Vvz/u+GiggttLueAwFEcCcYZ+/3mqxaz
WiwM10AACkVhWp8U8pu6rbzbmFz0Hn+cQNSfczMl+z9aEki0qWFR4GuIk2HuxQNoCs/2BET5PL8J
etYD67j1bZ5joT4rz9Y6s23yIqr2pp3cwpjeUhVBcKCpTq5uehrAWFy1TA92yzPLWq4MWKXJhKhh
t6Z6O1tH4/KRdhXGBMETMiFItFYg9Mo4ZkRZ9S4Pd3utF4JtP5cn8B4dE7vcBtHPps7fSShyegN4
+aKS7dDhTX8osIfGrt6htD5F6N4RvhujJJQbP8l9ffgylSZV4qQ2wa6Fp/d0l+BWksas3XufcQv8
pH+iMRQHxuzO24j9fuicbcisj8TBDw5idXXBiTJhU1vpW5y3Bn4PlSQU9ckFRxT14K2xvkV8F6tT
GC/268V+FsdW8rkjpCYeK4+GCqIB0nD59xBuC0RMGlbEBemGsVBMM4VkJqJEEFFbF+YJQB/xTwhL
PB8SQc3Bx3YHej5PwykRLEiDN6sk/mtLnArDR9u8bMIRuQGPlYBjMHSt0YiAgCp7kF5FlDRC2AMg
Ivv6IPwuCQ6sCXX5NWooeiXU+DErXG9UnnfLYLv+x3jhkCu3PBCseRCyH92Y34Zz07eQ+BqwVFTu
5Uj6P5HFppEwPpiMKRuX3UVPPcewI2b+IFrRLLnmUqezbLJn6egpfhep96GDXQePFoXW4CrqYWGw
dLcps7Z8HUJU2+JnHVgPaaJ3E9RBoxffsPgBpX8hd0S/O+5pS1srNXR+W1IjjdRECK6/MdoF4eHl
tZ5S0gKc4ygWQrl1FM68ejOMI1HnOc4n47Se4r6mUeshepzl3Tths0OtnC2qw5tAQZ+gjm2HrGll
VNgwhMwEsnIIVYeu0/8XIzZIB4Trk41coU01OH3yZEJx/CFbztAu6in/CsQXwubCCSxedRqvaewi
u2y+K9/bJROkQ5p1NRYro4BX8+A/9r9I+8D3FValBQy6YGbTzlH+E7lEHHLwaMILSP3ce1wWfgp5
CD0wZX9YXBMl7hE/xJMmwAetUQByTT9W+HCS7mZd26nNpgz4GDXIX8+dTTzXrzGLl9awX4XYGRSq
/fDyqPZJ0aKLmnyXm5C/L5aTb7Y9o6K3haibBsxtgm/lPZoz5IzCll8xlB8cOE2cIRRjcRJa67TD
Dlsnl/nIG0lDALFpYCOGiVy6H3KpWWcTFa2jKs+IEDJ87t+HgRoEyrlh0Yu02euCDP8d6aJrQ544
v/P+6Cpwtpj3z1vDkTTGBktiWpoNhimSOxT3Gi1h3Gq9hBdOuJ64lh3kZdjRNnWcW3S5sbDYriu1
wZ9tCNw/X6vTIWEN8dwGTwD77m/zH6hvJ0JbzdhaYxPVbGOGDFnTzrM4Adr4mug7ApuHmhW2fsBI
HSbPondpPW02HD5EF7czhmmay4WlkA7tD7GYLy6wQu5TrQUb4/SBmBiVB+lBx1rmKx2nTyr6Q9/g
MxrDOSTkdDcOG71oJgBAq+KJZssAQ9mGlnZH6p+zhBmbFwt1lsgesLYXbpWKucF268QWGa+oJjRu
hdWux/drXkGSwGcCe5MRC80JNPDOW1iKykKSZE3RwqDfDARZ/0XGyBgdMrwg2k9bchojbs+WljOK
smfAkvzQvqGGOioTZ/xPWOlOI9hNWqzrN1LqKn6uqLPTeuT6Q/ZWspN+wAX3T+WGyTrjvzw/jk0g
5pAtgOmbWgbwF2V93ugC6Et9OtL5jWVS+3vu2Y20PP3CXc/u8mQtz5jXalw2mqSMEwCv08Z0cHR9
4CbS9VPHPKr0Tu5a36XOyEjgINW8Oi3TWKTnAn/5eyuhyufqvGQK6dNL1aYMHKj/4dQjZIRvD+N3
fwup3J2FIl9Q20vY4mKOwFCBmXvl0Dq3CxiL4RgpfGR4nRQqlQins7fIRP2esd9w3Xbo3TSoJglA
euoQd8BdNblK289/dhhWbq88MTJr0qk3U1qa/eNoB4Pij44WLjSeouI0RNg32VV6+8lgRqIjLVbW
o98DOnE58WZnieVgun7S1NtsnNu6iceI1xXjzoQvaTE0ZAbo/wOnORm5Lg48SuugS4lUokPiByrq
OqhJP3UTHgMDGTlKVGIw0fgfhQNyjF3UHQNnUnRKheE0inFGtURW7PbmHUbUL/0JwmJqeYAIvROk
SgPZXbv07T87n3pkp8Z0DdEij4O3OpjtcRvdlpmFgPA5IhlETp+ar6TiTZGYUa9fzQOCiIjocysp
vNx1IfesSkripV7peyfdb2YFb1tYdKcagX045bAJOgKwWW56u5o9LvYw60qOXz+I+Dgz5pDBOI3g
sISX7Wasmro1cVDq5OZk3KhGMhMBugkrPYd0GEiT9SirTqodC/BnMEgofT9/xZmwtU0IqROjIwjc
Z+WkgB/P4rct7vrWX01r6f5EZ1IJ/u0ShuOGUoRGleKZwdSgtOd5OlfiU5+gIM8PHREYR+Xvg3o/
nhQ/hDXunJHanNB0MRv8BmbTbwo7e9fYffcaMeTNC/nAxlm5cAAfMx8f3wriLdst4eXeqJVWIvRu
QuY1Q+JaLbvDrYLT69tvlivfFC4MlSduaRV+aidOwjnC8DtQ/v3O6iXhrTGqWb87NOhmYlomfEDQ
MYrmDH3vEes9/aUWmziFNGgKWZJgv0ekzZx5ofzJrOUdCKcdOTT6icbWGlBS0l0+OUBtLmHYDwpA
7hv4X9ZS+OXYfQPrqfZXWliOXAFOcfQYla8xvJoDS4RgDGME1oeep8Z6OUMAsecnNitEvDC0O1sC
QGLZU8YVdXiKYQxhLOv/fs2YYVdZo9EgPvU0jlreKqA8fVH1ttGd9t0zg9KCjSmZWaxfcIQDffU0
9lOUlnLsyIxhg3WNTID82/GFjsX29LzM5JrejEd+023QkROpzVGx+RTDdeyvc3aHVEMcIB0cltRp
3BWx1M70ndaMjaYS1qzO1WhdzVjSe1Igv8v3hSxL46h1Cqf6bhqnxauQczHePDr4QIiSw8Zpx7hx
iWPjmKEdN++6seRcUGaltw819PvXil2YCTmpMTzTSrNqRjvssR+aeFKdAiISA0BwuHF9MZQ3oSL1
eMpjgCqg9+fnCDPwMxkucYq06WoysyEMM/3ozw7ApzuRuE6QrcRsFFxIfCVHFL/nblyn8VWVx/wK
cVH5f1xcs5fYkMAtTtI2fGbxxo7KUdBzmmYyXicucwxK2A5qTu0lxuQckUM3NX+bUdBcFWs9ZwsD
+zzF+YmH1164NNLKqKbhsltkb2cHKIf5Pd8Q/6WiHlceKt3s1q+/dL+u2ft4SLuvq8M9htoRaIsx
AAXD2BVqiASkFtisRIUNpTeyFB+FZ9h05zcNUKyMkwILmUVJqNpmeHpZnYf16iuYwsoLHzDKbIoC
eMSVCesbHIuD4UfLRWkCDoOwoVtUZor5hZpOFEyk5wXR2VL3clPjmC6BiHiYfB64zXvzodZE0Xmn
Mi0ns1mGs23b3MIunLxZg1CbHOL1wID+0ht55Z2mxmP8O23NSN85V4z0nNuxu0bw1jLoenXQfKBq
VZDQVKYsZFvejZozAtLNGzHbt7Q3fVsyd8JrtSKaHwrENNpObmK4Ne9xnEvrzPH6UO7onbafo7Wh
QkDj9W/GyoKmS3tcYgD4s1KwQzrjiYdgZhXXcgquhOb7cuCIaWk7rpfjyOt7wsoo2TRji9YgXXgR
OzVC8+g9V6L2VDFEhjwHce1BzK9uUOa3O9GYiBdb5sIa4b6KrNyCsOgwjmWuFR3A3DyFBrUHfSmR
1zleOKD4tQPSzS1n0M/hOu8Pvvr4iL53AJLILIDr818tJAyHLgaGx+ipISmxpkcLmExWzkkCVOW/
ZwATH9LxttL4oY7JToKe4nnAt36geB58L27MbC3w3Ut1118GKgBN25wEjU+WWSWgXt+qEsDf5qR6
OszaC5RoQhQdAZB8JUhdB89kFPHJzgVhZl8XBwT6ff08DX0NnR2PEkkWgXSKHyGqaoWT28NQ66Y+
m9MW/G7tlcQYgjL35/O/mZxHcSaFd3zk3PN2Zs56gw6jUKdOPjREVwvx9WCfPsLvvDvixdstFYdi
wmmEFyopf1bhXpQjEzBFEAuRePCy9G1B8DD/MbjbshEyw+v72ZC42CyYHSYyNvyDc62A2IC9qchb
zAP26aku70FDILJXFwQZNNK8ePqR5hmKQCkYMVTUfSS4y1mfTN+wxIVxhof9+te+baiP4JmoO4jS
uPofyfSnUWKojIQMsIkFTP2tvAD09dLMmR+er3pI8HHo9qAPvDQ0KPs5IYy/qZmUI16ig76fu741
MO6GhgusVWOF/xL20v/zjSV7Ho/gLW1H6PVwcqqzBtFb5mjGW4B9F9d+UoZFu6h8YYsExl0eksne
LfWCUNPQfNML1+p3VAZhXCMufci/dCx8quaBUrli8jl9kPvCQii0d5RiIQyAD4odO7Q9WlSQhdV4
GqD+kFryPHogC/RRlDyIERWdJ/EMBKBtdUh2AiOTGGm+DXShwgvGfVCjvIASDIw4gJw+DlbcuwBh
VSuTHu3sTyUlhsu7gKm669W4TWVfJo8MFIgv8PSyKu9pzN7CkxpsAX/DUhWjyFID0CweFb+hO5hN
A0FcrZ7fDjCYoqN/uVx9kCGCC1eHzaaBva1EEFWhXhyT2Pdvfzsa0vxItW5hT3bEE33ZmK5qFSCM
gjchUjRBJwFHtrQWycpU4oPAE4UO8nr4OFpZJ54umlnJWpl4R0psMII/ZJh9DmihhAtTHIdZI3Kj
a9tFpe15Xh3TUyTgMOnZVLHG9p3wLXPJjG5Uir3U8pySfPi5XBVSy3IEqi5ZDJs0oHeF8+l39jO6
68pco2bcP7eYEob/MDOTIzKQNs4xDXwVaHhUns6w6J+j7wfYKOPQgZpvWwWUkGhus4ttXjt0wo+J
zbBQvGA8SbfEVaEwfvNuEp0sitXZX+O962FTxmqeiYO5v3MhPSQYiKzalMtnSxzViHZUqYh/926U
gZoCduB7K41f2wvFJVCAVSUKdoAd+ohJoc8PI+aAQkyIM+N0Tz3eKBqoSlntNU/fEBo8RA74ZqyE
yMzRtSG4NqrpbTX7saUdvXAf7Oo4TK2eaUVL8mqt6eWluZdNQAOj6v8faiKDSOpPtpU8BKowYM2R
ak66QEjQb0Yt5Cxzp884bZIQn2/X8ofBSxi8AElZsft3AqtF/w5tFcTBu8fRYOzxrA1Et6GAZ2Ht
x6W/LpjYwfi6W3DM9CkPoiGpbWw5p8cUP7kfVN+9MuArnrm3+gswy3IRY4CNROEuTqTxmrx3NXRI
YjbXTzScXeXrciwoxEmtFlL43KGyNQpNq+WDGt0cKiMNFWRJPq9RiVn1d6ofnD+xX3M9KBDg3+PB
Kuu2opkhvFZB6zZ8yfPk01rpxE7Tw4wGexHzFoSeCJqq+kXP66M6jwrFBPXmrnZ3h3I2zX5xSM2v
ugfsv35OyZGw+wceM5hZcwkOK5eHwURt1dqedKUyk9NIDQ3dBJbqOyAcbm0N9yBvhYmQiTOMek1d
2EG94a4GO1q0uTvNYxHpQ5ublpfjwzmpmVg7av7BMxQWmEtpbhQu6KGOb/OYLvFRBuYG9qo1CNxV
8uOp+eeWtbQq1kemfkGw45E1R6j2np9I/ymNwmedTzCYlhRnqcZzykQwYd4gqVHjcApC3LpOefk7
9N9XWXKy+yrb6o6K2bshhnDuHs/C5RxX7S9UHfj6/0iLB01QrKOAJjDmrTeSXylWNYQkc2KTyW+/
P65dzvEQBhdSB3qBGd2XStGF32QMTtS54LwBdRa2LFrFF1TawkVlJnmXoNBVowGTLmCtDgeNymbf
8t4ikq6ofAYocp18l2+qGmhEwpfiPyYIhvx6jxOwJ73Z62tzT+NOCPBKB6IU/RgymJbkL4QEZ4VB
zjDD/tVoNSqzcjamrCRsZ4W7x8XvnmpRwxUEwPD5zKLKpZZBUicv04/MIxUnledrVgkpAojyC4BE
y7r0cAQvgcd9GYsGZbtEFuztTNIXxRG9AKIFPp9/5U58YHBEIZMjgWE1WZbE8D4eDM81R3rkYlvr
YLFgVoQAxk/l2TTneZvh1hbG5EQ32/NK023YhmOa406AJiyoxtJ8ywt3twgkR2XJbhenAeFA8nP3
KJC4Zhq3Ze19OrwJq4DjqtIgLb9z2/RA5SpHHP8aIKdW7NwNmk/WWDeBBwcc4Eb62gL4qan6kQdk
18haMkV0Zq5mH/QQTb3KrgafCAiyobjXPUtMx2BQGkCZRUDX4QMU5RsAHhpwV2F+ofu2pCeinX0J
wZb06e8EcCGDXT3KmvXJBSS2ecRmqEE620lvc8PD2NfHbCcVyZXGndXVh6Km55fTTShzWo9Yocgy
ghXlxZC4E9lVOwxCJV3y7yEgs2omNAW8v+zFEPQv+0+A9iVnX8t7v0GfXjXDFBYik+3M1jSDqCYW
wlsR40O1kwPhh3kLIt7/dvVBbVN3nOL7NrtqeRMc8xmCIrkG8d1/eGw41dOI4W8XPO62zpMgYT+A
XnX9tWgO/dZrPe+TsKF5BGt6z7jXnEiPWsheOB36ysXaNvErALBcBzvr9HP7gfvq/hwLOj016pp3
/ed2hh1zg3JxLwvKDqFnww6p9gJSW9KvslxLTQGuImNzlpqw879tjqvDFRksFVmv7ZMJo4ZWmxU+
fnthqpKj+lYQYs29feEP1vd+eBPR92PptzdTE9sy5wUYoLURdSDX54F0NPsqiANKpc3KTjWrJ5Db
o/52dDPh+YzHMocGZiZEnaIju7IQRJyvfT+hWBoJVzF+OLIO1K6KwbskezA5IOzNZWQ3nmMiy3Af
mqyyeGIa+3W0WIkBwG4FK0YSiRvSTVKGerWbfadLoSJQjLG4ArPdR8GrrNFaIX0xf08mLdSe1w60
Ojjw1gVffv8C7JC3PKyxzbPLRfLuY8ZUpPMSMJqjVgYs53w7XzfYZIgD0+lTh/bhDLE4Y32kjb19
yA+LtlO7UlW2f+7/DD0r+LnovOp37exb7m6dgkMLwvaUlSmCCKoz865bGersyWfxXaLnjfBFe7DI
4hw4LxFmKZMIf1wNUdgHLo90Ad+cWcb4I4/s88BvW975C5bCTeeNtjm/smI0K4HH4/JmdyEi+Yxg
jtsOPxap9xD3zgFfh2vgVo8EIYqmoRuWgMApzK2stOb5HIeCU8gEwf1IDx71BcnL74WmG3GBaCuT
Sadm46LaiOkPJldQJvBaVZoT7CY4nzHkdOsPxdPLnB1Hf5OBywNyPa4NsOWlHUKmz99MIIuN+0A9
/mxZqK/uBVr3UWaN6I9U7uQ9IaGwTwea0lv1at9LNaH2bJZLuXrutejH7o15xHXnLqRa5hR9PzFi
kP3UTS3o30S5ubEf0XOzEJvY2b7EkwMM5gsjmd4Qzxc8aFyYgKyW0gMFIR/Nk2BIfWuPyyPF9pie
mt/QeE+vHR8X0ykxeXVt8NmXxe7J7F8FYrLtbAzoJBhG85HGtOYbpJFEPS5KCQjUcgCBZNBVofXU
O/LCOTks7DQHRR/N9lE4dCcClSiHCJfnI4UTBxds9kN6k+OzY2stkgVzFA755rhf1yKGylVPBIqD
S3ZIiwMn6Y+KnUkEUNSdv/DweHnucworapXqyr5CJZorbJiWsZpOYBiCQpyPe2yLJSzfDh9MdnMj
nJ4t34XQqsLuxavwlqX4V3yYBWF/NrpVwjuJOtAhhfeoTmPg8uTujOHMe12d4SFVDscIc/YUw6qE
dmgVALgbIBE4LX/fgisxrN5rLlaTcSvo5bbc955IOvb1C+Q3QqGKSdAPQVmTX0aO5t1n8p/6dPw+
N/lFkrsPhEzgIuyFD9/ncbvrwQ4mndULr0Mm0GnciJf4r/sVnG5NkouFD5aRwtaUIW4B/PSVugwn
yEFoO16XqAEz/B4GnL779ljbIaMwvv/fFC2sRlrZ7ANntXOm+ECdu3Ab3VU0wTAGsrSMPAIBjfWh
NUOSZuPwWY6xELFwvAqiCfJ8G+UB3RGGSdkATXqtCMV4ZGh4eVrDWTd/b/BqvljNBMUi7jW5xUcY
MOxvqoC9FzeARK2UT3JQEIYmDSaBqVomS6Dx9yGzcP798cjWwPeFqCjF1rTAi98TaIu73CH2h36R
hJujlwxQfmt6tEYeKgjaz6hERTX/y9JhCg1T7LUeyCXrV/jQcGQzMMAnpPaBLsiQh33wzQNdljti
KaW4NGhms2bwoqnw10qf7oh8lUI9AxmQkVvE7kHbZFo/qBaUIxJvgp78rXBmABuOMg9BzSKkMZoB
ZOVE4oy53ghHUQUj1OW4dG6khDrZbkkpQWigpGA8f9XEO4XxWyEFpKflCM9OUiwpIHQ7IAW395DS
29R68L9u/d1wjpm1ULO3R7Pqcz91Hi+xucGTr/z7gsYK5rBNomq5yIre+aMXcdlySQZQGoeapWy1
xHRqVJ9IhcociBJv/PNv3v+H56rS6rPlRVQYSD+SUy+5fI7XLjdP9ghYkIr1LI0bXtaat4JaLXBQ
pXiKj/y/5yd1ZUyCIN+HdS3zQn5JDHuDPg+iVLkwask1TvkiMd023Dqos10rxye0vD5uQl2M9lXo
d114PWBkhWM5ZRluaRR8jRc2z1gmspGCE1ryfDfcFdsorpe2OmHh78MU4HOQKKtxkfYnWRGp7VD5
qjQ5/l44Ghj50fAB+UWUYMQveVmf5n+8ShqvPIeJolcNz49+eYDCJ4z2k+lqgqH7VrucLUIMPF/v
IZ8m6M/fz3hHio1B3hX36/VI6YUdGD2M7Yh7lXt1QNkZFCzp9ERMk7PTfu9mdPN6OkN+yhHQNVUj
QfKj+TzcPRAN7DEW9m5RxW6447n9YYQ3L6wcBW+njcY651RSzmWVY3JAM6OIWh5JN4PHj9m4BLOU
szxS7grsMfqHseN7geRkVXDB78zeTM+54jXDZ63iB9RbsSo6YJyb2YNC1r7cvRM3/iBP05M1HOs+
zDE4jugFwtinPNrXyBvj+pCfuO+1CMOoGT/oxmUjAIIqcvJ04tVNpUY5am7zmXB1NV+IcvH06XWb
Ia9ufT+J+ZxAsO2+x5F0jxFTmqjMsGz7mbW5CYHEI8KG7vwF1HNgAwXl96H6R5LLGbB0vFVrvd6P
wSo6wmlc4XbE9WGGy6HCL53RdSAMp7j7pxcnBSKgNRLm/nL40VvVgKqzERfCZWUolaDGTeISSfYa
1I6c5VAZRgyPMokY4DJawuWeaQPSW8vr1rRYLa9Gy6E33PprM0s6mFV5UCzlxSasSVJt+5er/VHL
lOFxdLnt+TvXoJijGxffGTbFYeNi1A7QvxR3fPxQC7I/L0N92HjZpg4WA7E0WUkplmvNWRDW4DXO
FmDdUCSPdxvPBbin2PEY0pUSF2n8idqatyhWWh/4Nd1GQnCfnlAUGCdGLb+MDErK+V/LNDiNknTG
pWs2Sa8CP+gBdDSfo2lBnAhZ8awXFUGPAB0zsBPmBg1npGvHUXo/SR0f4O2fjOU43fAowRZCjdCA
xiiP0QAZSQoHX9klWI2evYt+FDkkWlIAPk4blBALseZwL9ZPf9rTmAU3hEotXlBmTGOgXwd4gEtr
DY4dyZMKDcJDw1EFwbNhdPg2oMx/zCB5QDs2IMXIUTe1LywT+rSDUs+vAjNVhZWPIG/Sgr/Iqf3O
ziffquMiZLFk0bDA8tGMlz8VSD2eZSh4Nx8dVJd8EZIg0mbMOmFAwPXliQ//jck3+YS1vLQfmHtW
sYFjXTou1R2UoIxecTapOjNgl5tLqa8m3Lgs/Da3KjDTLzoXYacJFUSPblFdlpn2Z9ld5tcOVvbI
niTHWienvuLuN2me3ka0QARPFe7HYwQ56ACHEx3qRit/qOytySOeR626TOkEjPZ0imCe9eXPlpzI
UxXTuJtWxzuQrEw0GHwhHT0mhxURAaP0QkORFOcjlw4PdC8q/dkMznA+2toweWRgHdYQxtzwdOr5
hjqxCd1yTgfRGOKyIbcRmS6KEWOzYdyoCOgJAW1cukfnsxuQE1ocCG0hFwMnc/FyZsUVbom8T/QI
6ku0HdsKAerDgBDYgm1FqXC34eRWJIskzT/zvHBvXLR4S/vYFigcjR6oi99CsdJ+reqfy8GtQSqy
U3zue2QPlkmFfrYu50czNZy+A8OylL8Fv0pM32LWUH9i6pvAhphiZa3AAxoLLNBAwas6HZPcH+xq
FnWGL+zYS0ozAhaaMRXncwrqFWXr8SxD0U1lU4Qgvx3HwmkESp2pIwKQU3lbpFdW+iOIYnnTa2Jp
i+LTmQeXx2ySoGa1srPQSq3kgu2gJWg/o+Wy58PfDfjsHvLP0uBY3Uyi1foB4T6KJgP5o3qbjbZG
QQP9ygtP7PiawXT/SBCZZd9lEdQRsLpgyHu90ROlA8fFO2HLWtXVvNZIe/+ePfBAwMY1Tvc7gjg3
6vRlEDrEIomlrtqUkjLKdyquCuOiZLEdEJ6G74H6xaG1Rofx9qGDl/2e78WLkovJ1QhW+57Ukvl8
3VWIlACGktjosxiK5uAt2Z1tX0vDpH5ed4l7vdWCA/wi+JKzxyiZVUGlS8OgkH5W6qcwdr4/YxE1
TddmZCL0xQK0jaDI3CeoQeB8o2aY/1KzbnurvxrzA4HiI+pswTbJsfQ4mNmH4XvhKwQv6ffd8SY0
jjy4esg8CfzBo9oYD5SeyH5txfrQmUJOU6ePxDu7IK4IsDcNheQQD5e/uu8GVLHhTqRVtu7YaLv3
q8rVc4MUKTBLo7NrKxgy/7gVbFcchJsF8FDWLhoE+hMyzweTMlDa+YyX9dFuNF65RDDbLYukk2fp
Rb0RPwwXmSWAdY82zR/FN+5a26xaX/G66rgd+JpT5NZ3oTOVmjknNojZkk+swyufMGYzuAZSS6mP
zihYGj1E/qQB6nG806/oJoVocdlZdqa56G+rQ/gR3x88zq1haB1QcHu/2tGr1Ivsj4vgWGCJ5swg
9Lhs6uVPH1LO+5H505znPtm26VjW4WtxHwiFMHw2jQvmlVZ7vRDjekCkYCu7AGcdfMirjANeCVpm
SC3CUcykZVyWSiPS0+Jg51qJgtqHHsSzDasdroGByUKMLHfzzYO0HBzn2q1QDfWkCdigHBQ8z8vu
RmMX6jBNJi5+ZAEvrnnlKFJzPC1m9EZ/O1qroykWdv/kGjlJFccnik7+r/8+bouZtqeHDJz/N9h5
uuH8thJQMVa6trHWM3kPY7M+YFR52saIngRDjniZLvG9xsByAdqnOzufJZ8JQQo0XovPb5oOIdC0
7nW/u+ewApFUWYRt55bSGlP/ysl2SDBVQ7VbJOkuVHKhg9wysxPRJm1jjxIEboKRBw1EuRZcdBhV
VBT3l6HsD91MZOQXqRR+cYEhEHWekP1N4p+XzkPa9r9Eoggzg0TOofBpblK9seFSbG1tCKfM/sbc
aVukLEFuJLK4msnWA6BrA5n5rKThDOBZBNQL1YZUx343n6fnz512g4BkxaReS6kIKsBnWOH08Qb4
aajdZ9Qh05HYEI8qa3I9GjwD4bFjeOTjXUMI6905ZgFXUvNeGzFqM8yOsr23Y3slhB5iLJ/+EG72
xPfSDJI+nNjVbd9ZiGvkuF/EFsCX1Duc9vQO+dK/WyndItz1XIX5907LnJYt0iV2hVqFX/iIjXsn
0TYFQGrbdfJQm3C9MwwmlK0MQCxOitlmdNSZ7+3ySJbTVffSHSvOycv0bPVoApPGuVeFTVvq+ojI
L5TI/d5Es1PXWBMPpl791EQIjfT+EEM/USe5WMv1I5IVkgFl/51ud8TMwe+nVRbm5XGAWTWNfGKy
TUEHFV6v69Kldcb4QeVpY8oJuyOwPR9sMEa+bRH/X/EMKAJAM7K4O6nQHTLKoB7wb6uFLEH8NrLc
r1i9yp/Ffdiix9pDDCbHfp86FJk2XNwOggfigXZz4qL0saVXxKOpji5FEovj5lqf49FDifs1zyo8
HwRxH2rfyxzZSp+M4QKxq3BOTL6vIaC7XOAfKUt/ffhOYWXQFjtJ32GBFSF6CppkhmNRPHkEAa9F
gBK9ExT+2hHXVVSBBrYGamaBwLG99WtzEPhGXyFnK3JeUSvPPMGJk+2A5QQlOoWRvl72IaYh6gP3
NdKvsWys7dJMW0U8JIJmIi3/Tih4OuuKk5L7Ua21XaktNqdnQf96rQGDL4D4PMbU1V/6n/z/3FAU
YvpmiTnpS0Vv2SpD8fI/jN87Hr0SZCcDfrTzWhZo6JbummojweEFwU6Q8+7ADSM8jSntT2lfnjCT
JFkOaQYwKzSDKszCRBQcd7xfSYTdIWfm6Qa4xn4Lm1326Bg7DljGHGlqhOt1AwkZKxLPpfcnUueW
xqxHd3s8D9mmzGj8+ZFB7titvoptNN3pl2b5rotOIZvJz+lUfKPJc/kM5yAbvZ76WF6JSp3Vf+XR
wYIPcCH5LohTcAJApiGDE4pomCdaB6CkRt4zmvXt90jmJYlp93R7OWzLccx4WFJjvOfwRNSuDjqh
i1LjxwT/KwQGdMQb8FhO7Qyln6Mhfpgv4pwJujuOmG2xtodX6YbA0FsC+3nZhbl05RqoJoUwYpr3
WIIa8hVgBT9NSEWbCHpGW9sGqbFgrmt/am/ki41ov0UaUUV7ct49uN+XlQdbbcPZLp5UDy1pjX7k
PDassOe2vcYRqwWCWUJsFQory4OsnYnAHvssRFpMkCoWHWSPrPYIeeAt7Kzjvm9bKI0m6Zq2WSrf
8yyC+N4mfbjyTP+2e+8IlL+6bbGJLfosWJjRf1KvxLrC+SMOd3YgdgkYpj4arhEaHAJttb8m4dFI
tAQtzEZaZ7TQ3tlFAHlopINTfmMeQxqZmGJUduV+rfC0nfhPQ8NBiqpsaknWzuijpYsHMeiiuLwC
EZuwx3biEkJcVVonqj93+a3b+zM+luMjRPEpnGd68XcCoNWBNrZoa5OI3F+3/OJDsVruCyJZvepd
EGOBzv1kAH5NBEqvIrLFRnFuvjX3ihen4SaGd/1Mu1IFFk4MRIhbVoj/W5v7CrU7W+4Jh14tfG5i
y4QTyvzaB1lE6yCeUEXYaDLJNPqcWMNbcW7IYMRZMGKHdwuPm0O61fuiPVykdjkT8+bBVDV0gEvW
SlpuFXq5x/XqAaE973mafmNNUfcjwwXMOo8bEB22f4KcigBI3rar0OzwPPTGRD+pcMhqGcJaz4RF
bK6WaxtqnmpTWECscsU1j+ggeAThdYVgvKPBGflmW2u14S/FnYIsjiBZVh4bRqus8Ncn1MeCobd+
8FxqAJgXGeUyqTcJFXlVrfOAQ6Z6iIQp0UDbH16CTQ+HyF33nijxTnq/olAKCCXMau0nXDoYFz4K
ygsxW93WbEr+HI8sDyEWnR3u3+Vw+2DC7ZbKYlsJvfmgcIO9d64IC+v/FlNOkL6dNqs3tN9xCvCT
YrBGxgI4r3///2kL8rKE5YpQ058+T9Psmvi0Z21RUs+VymBteXGp8U0TfjTdXipsBoH/KtMo8vGv
44FFMFyLyVEvhcLc2p8JlvXqgqE6p4yj66ZbbdwS9zT2f9nv9HBPvNdWMVuFdvxyXV54ul07yFJq
3bqVm79GB0WcQ/7l3aFIZlfksSRxpsT1tuUpK4oYJOpK56CHXo34ULnoCw29sdnjz1cI7cjIIqDH
QvdZzANRin5ASEQX7q9yhO3Etpy1fi69b4TT7NBaDetVCL1opIyjGHinpoWJOx6S+14+8gJq56Wg
BcvMbaJmtjTzz9n/i/b9y4B3W3y6PODEp0xpswGxusAlHRw4RyGNAVqSIDSVQQbRhR3r1roFRgAu
ChnwcRPhdO3Q7+TswvPiaUw9oGuSQsYNpfhnZBkqn3dOQHtGF0lSrEYLFeUExE4NbS+QPThfWcDB
/42H0WdhyHRIqtWwm24tdr/N1AlHA9ossCUrH2ToFFf2spy8ZQMgnucJvLAmVRXl2DY5o3a1/Y9y
miVMgVWGoi8/LrCOziIxIGxbJoCw1sE1Q+YiDZswnBzTwXTUgrCOg39EPaCpW9lephZddxrBt8WY
eTTN1gPI0IU3V2xoTTJI7c46otYXJl7umMCahfRqclogqcSUiq0ogHlErTcSGUzetzYaWL7ShCRX
dBNJTiYsGAz+tzVYEvGoYQZeILHGvPEKkhHIDl95qMv0w/MfXCuU8rgjsYMIjMQ17+0bSE41btg5
VFpiXyI5D9eUyIKTdssuf2f7Z0P4lsvTqblJrJHrs9au2M2UAQlX/d53/qVSH+fD9do9N+z9Jchf
QzFkemRubXovCTqel1hzdPXppIldYNgEozT7Zl2jWLHXLyem9xmryiXd4Td58LlrUECNseKDBqv5
lApve6x9k5BkZ+D1Abt2QOOOnw3xyWhXnGGOK2Acr89fYsThEco55gfnhSTqgGObTTtr0+5AKpZv
7nn0164ION0oEeg53cVQfHOEdVznW4/JTJrTx952+IxK5jdKPjCtB8Vau2XjS+ignh/z8sPnI7XP
OlvzZRyaxWhWhGz2nZPLvshg34QqDWpwxBdhzFo19oSh2vR/s78uouJg806uCbeC5MO4cDKU32Ap
BXSMXI3BSDKfdN4lm+HYrUUI6Tt30xOUIkCHONPRgSGUwZqjzaxto+YvA6mCcIz4mudvMceHhJj9
XVjpXOh27S9piXRNKcNsInES74w3/X9OkAELMkapjNdHKg4HP8E700YwJKuYj04gNgHep5TEfDau
DxAhUTw/sAjFldgmtUCdgPuf8fQLUBijijOLVRvyOo1u+hWAEjCAe+Ee5yH+xcBtEYGlHiPLEyBw
kL9WSsee/BQGoCMcqs+VI26fG0ziiKRvjHbyePIORUJLuRau52gKtMhD0VeOku04aHViT/1rTq3T
L/83KGcB1BsOrliJJ66fDjYb70vnELHYP/6zTJ1DctKHJPYG07atx0GrsUb3SU6Og8qgQsPppNUp
PXRYvZ7OqRVElZ4Mh7Jf8tGOsIyNo4gShkZ9/GSm4U6134f1rddYI3aBrtqmABwdvt6eSKWy0Vge
whHbnWuKC1zaK1OErQjEAVSQ3lID46jH8p2Td1EJNSUrsIszW6kT2+PHYiNrR6uKsSPKXu2G1yzO
53dYC/+lOAy44805xrlzSYQbjJ+DnbNPOE5DFsPbToGyDvo+BWHTjdpPO23GhrnMBcm/scd3DHMj
/u5gft51bERlgG5YT5oJDsaOUcG9VJovsl+JSHXitc7jeNsHyzCzRVDCNRee/c2WWbJK0ogj/EIH
YKuiy/2eR3osXu/Hcsrcosqie+uYTzgzls3YBqe5vAJ9i5CnVqQK/WtfC0SYj08c40I7J9ak/5hj
jAesxsfnRti8Qywx19LhDCma3caVh6E1ViVTml72J8pKaez17e7y9BOUjFevoZkL3hEWJbuygxdk
+5mPyC/LzrKvEaaFEAbYEZCmyR8Rmz0Ul9XJxQeNt9iocZLlUIHdkr7/PycWANSr1BhjDQAOS7q3
grUsRkkspGifme6cVydPgQiNpJf32p8WGsozBHMzeWuHGUxKf73nwXS+HA/4HI2CfBPARLqfsn1G
h399y81gN/QljEfZmYRBNg9iwJl6PsDlQXk/OdIt3HNQzfXAL9kQxBWuySAxZDtU/yJUd/BIM2p2
xqvCWfPrHgU8pZhrRkW2fdnLXPrbl62IeDRQGo5DGhFJPQtVIBy/7BR0qtwEumRJlT6PfvbseBOa
ljsYcxRqaDuFS0zI4+XYSlGuxQWIoD2u18Wx/C/Kz13ccOWGXAiu7mT4VF6FYOHDQ58bn9DgtrQm
kaBw03yKVOUTyPR/JygvV2lZktuxBuzgL3M0QFVk8xb60dBpRU6YFa1EbfQdd8CN7YtSymcL/2zs
6ekB566Ovh1H1BbMj0fbxpB9gyoXYYxNn+UxCKIfJQW5+biABgSmCBtY2sfDcLPzURnH7SONEqHC
H3rvki3FEbACf+5bxAkMIZE/Fpx4E9rHe7SlwJlMUDBgK2YQBaT2a2xMPaaFjtP25jwPXI+2mJDD
nqnojd5fS3Yre4wDfFwIrTHmUKxLZhVBwptZ26y1i29dfx96IiRGUEKKPMN1fpjR+RbQCQkPmEF9
qIMCk9Rxm9QEWrwhFcemoPDjDDpBfGfseij8UizM/6+tnd9jRqiQAPZ3sj1nn0xl8GppjVYx3P7g
Ss+p6P46CEnhCqkKRvupE9HPppqmSeYNtoYolmVdJzoglTlMvGIHS7Io+n690lwGmtRnAgHxL30O
CXx5dMmS0OfFqcWOS5XXbfVIOuNj46HR1oYQxlJDPMWPT/avK9T/2SgaXxiXh/qMasfIpNtFesMK
fk59ea/SJAzYYp8kMcMkqvCrlulJ51m8Bdl64+tcUrslCAmogLzrm0tsqPXEg9sgQUvA88bN2rvV
ada6UcdnE49VKOR+K9uTzSaCoWD5SOo9XvcV2vzgq2UEliHFGzCcp4r8UgEprj5ZyIMZe924tkfs
RMTQOqacOC/hnuaC3WyeY6s51dJHIt4Cv2iXHZcc0bIJJu6sSlp71Kcjg92uB5uHR6CjurbzIUBw
dzvrroDxIwmPLl2UM0jkMitPStFGb/EuwiaeSUbi+Xkuyrl125U23vCBcBPFooRpAdG8f7XpNC6V
4GJIAuCiXcoNYLcIWpXgnY/V0SaCqucVO/Y1jtjv5zF3u5QGI/bfJp3Dm6/Cd6yA+movK0Wdgehr
/Q05h0u2W351pNo1dJ1VU5e7wEzozxZeiaY6H/SXq9i0lnCx18QG9fmUw3z2m2GX/OBoS9ZBCEkF
cQDpj17EuM0mAhk1K2ahk1sP2f0GJc1BLtlE49A2QbXRagavgbiDvQC8KUtKK1SVegd/DmchvM/P
6NPAaWc2ixy9O+s2iw0NZkPzDfKwkCYZr/BSz8KU4nBbFrdPtoKLrZ9bv2VTPXj7W45qV6gMvJPt
8EnJfjFSHQVjByjJQr0hceT7maYcEc2ixO9//ukdOVSQIVN0739N7TEzL9gUjhhNPFqagfAw2Cy0
qAoFph8XbMVvTCvCefCXwA6KGiNOTNmSJxo4lCC1iDldXS8TxAWmS6P+S6rwWfte/71CLC9Vdwwy
wsrEaxJ2GC9Mt+5T8Vymrc1p0RF3Y4Rf+BgcnPuQni2q2t/KK5GUG6lNbFTF83x+7ttgNS47A+h3
Z/nT78/bPT5TQGBlg0+DitfjGeSsbG4ubpw9t8c/qXbjUVXCzLqVPk+pZXQb0flfI+/+FUfNWMZg
Ag+hoCHIPYrwF/PUTkk4CxQhXFQ2kNdnxuRRS0wg0aZhku85M2NeMVM1XwGJzk2AV4W7/DfIutMM
6pZh0S4OsgyzPUNiETGXtnJ3q3FGVXTHgsgTnJOPHc2QqGafwMW4V0paKEA+5e6GsYBh3A9xsVu5
dcDaEAobTjSQBM2AE86BHc8wFqOszOSJLyNrcATzHfyp+3oAi9qBi7wpAnMDCpdrlHBn+Obeynpp
1l4dBN15l3WNVNNkuG1m4Cw1ZVFQgi50aWx+aAuyAj48rDEe8UfTiwOwrMPBuJQ6IjytdBMOuMUM
uq8f02tHEsMz+EkyxvQGzwFVj4ejoWyPPeXlUckykp6wDBX0YWjC1Z9j4PK+I+7LQT9nMFxA4khb
3fTbw5gKBWGsnf6qzHnmKfYIVN8kOcXxODbUzLPKatNSwTXv0RMapHImusXf3HqG+mpyAwOCyStb
JZmLF5N1OvsyWPHOJG9jH+br9NG69Cttzleu9vJ3OBACePCTm2KSp6kmxevB94KKmVa0BEhDHg2+
4SLU/N/tgruyKNhRuO9P018cxHik7cHTCszX12fhKYmNdgCjgNWfZQ6DhXzNc2BiOCPlJcWlEHQB
6y/mqwAe5sIJuIB4cKd5VT6l0M0YWutClLDNQEiCAM5DkGzO7l0c8h70jSXA1ZzmQsiMRGPM8ZYm
yV3zk6oJ5E7oiduh12p+z4CdNDsG7+cdiNvDeWOgfTaxz2P6Ik1zDkJoe9dryEoQ8Jm1/+sXqjos
4lvcZR50tTnRnwTbzn86DEoCwsFoZJfHp1L6qjyt1k3Gr0kW89JunXJKXNWPcg7Iq+ifBLPpXNzy
P/RybUE8tN7PhmiPkXXS5fXYUKVktuvbKpVXgUUuGBfot9nX+BQu8/h79RimOefjDaMfhyD4RGQ+
Bdh+ZFyK6N1Uo8eClPAK2BZmhSKx+IH84KlQsL2+W6ftkZfeS8WsXF3ZlWtxacOYbYRflzVem9/D
x7GAZcNeg9uoOTD735jEIESN6Zxy6zExypNPWLd9wHf2ksbEWFKZWpicaVQbuhhL7W7s85sUKUsn
zavY3UBXiD6+DwDfIda3uWCgToDFCpugJ9O4Qw4ZVe78jXjdqQ2L9O860gsg7YDyfouIUYqXnAEe
jbVYpM0IEgbCg8sZL50CMLnn4zkehcnCr64xb2NK1YrdSIV5xcZaVPaf9N48Ac/3w63nBcetKpfJ
f4jRqn3x5P/7O6lh7jeV88yMIadNvFOAHTIyPi5YCt3K8SyqHfjLTSByhwGSSi8rTML3qPCIstc/
fuxW0rMfGOGxMc8Qlw3iA914fG3ePseVpFozHXro3+8PT7oFJkEAH+1rF7AlWQ3bS5uP4+8YeXGj
exs811pvmpSeeqbK+NcA2P5VQS0obCwMc5CQ0WXJRE6ESZSZVr8nv7ekKgtKpLoDghO9yNHAQPkL
iOs1xFEdl5/oCJRsRNDw1+EjE94ZzDbDEs7Nx12gDpy8r05YzJriKddLtvErYHvosgf37HxqDP9Y
eoN2jIu7Q8k4nBaAEFRfu2SNPqz5K3O0USibmf4fqsb1wbaGnTSUBx+VFPUB4li0pSmYHjIdIs3E
4JNR2qs27tCce4cmCH3r5EYgZMe+NTWoxd3TFYsLlbwRB3S4BjcluccEbFGbtF6Nm1UuMIl6UEc/
Udu6dySezAyuwJhjoUCKwLMLRnKsl3J80TT9L/gIDqb/a0ab6G2hR9fyTlOZY5TkvzVkGXI95giA
9vhA73OdLyEGxibr7vdM6qa8mr16l6IR/b3laMh8b156UlXcihAqLdoeySZjpibzJJ4Kb+7Hy480
ey0mLgFx6LzFbmWe5eT5Is7yfvllymWbLJyfDPqyK6+8T9CJ8KKf3Ygo+UsUFlwcV1TAp//x3CUa
KyAfTXIE5OUnvfMl2JqwiQLaqWt9D8qu7VBELjgbr+FPjC8IuUvimfuDbJYz166NiPYLpMlIMlYY
VzWVJuH5cOegrIhjSioywqX6eeAvgNsPZK38f8uRJ6m8FtyGrJ20TJ2eZA4CSBCCrjtY0vuYcIrT
rpmhoBZ9O8BtXVh3XSx3a4koqSxVwpMcjyE12Tg64Zg22XcZ7SJsNW20s0UrMgtdRFglsWAsCE3H
BEMlzQi0GwEDrcGl8IKgqmYD392wYdb/f/3I4HGXUm+6NDqXF9YmhQiNOckRXcLTonUOQQs5kzs0
5QqOp/ztg70d0kkSYQkYWCCIkFN7y4cMZcBtuLDaqvJkqAwBiphg2ydCdUSP2lA1+lISCHVJO2AR
V+36yysc8r6wbjBrN39NAgLP/qJDjAR8Xg07eTfKBrNFa6+He6iWneiC0WrnjDRhFaIxFpTSpOmv
bgBE875zFDqz7AnBeg1hiJrdqlkuPaVR6rLFRQOujGxmYECzcB38K8kRIe5xeTGa4q/Quio68MO5
jTr0g27GB8tp8/2SYGyjvhQ0T8daC3g8peU7kD1SYAu7Za/LZT56GXYuf3cHkZhs5BEjkOOmgeD3
PuTONiObwSZLYLNYJveDVrRVfs2mfaC9M9/8btLlyr7r8UPQUeR5rUv8CnQ4rhotelr+5FmuIBV8
BPCUcESf9OY70BGb8sVg07WoCx2gjoR2W/FONYCO2y6tGJayDneyEqvhaKUMaUZbD1fiHezOIInD
uz3lHiwCE/qqVrvT/ENO+TmW9HiV5YMoyXtmxud3klpcI6cUWkWxMiymFr/ORodqoykJ5dEFZuJ5
ORgLU4y5wU3eHyMKGn6a6ERI73R/a29W9GLKZgPl3Z4TAf0llbn77HsJB2m8P6Kkxw2lu3zvmHZm
QTA7SnK8l8Ulx8VQjGHiR7WohwM/A8GX1Eyd4viTQxLIT5oeWFK9O+GzV3Nq/XZyxBDSSeK966a3
jHNnkxhspBEbHqg4GTx1jsQYi8QonDkOV2ffTmHFoXTmP0srZN6j3SzWHJivxIyl1aZtMkaSH/CC
a1XnsrtgGFS6RyWuA7QJDcB4RROFnUErig5o0WEPieA3HvxFhkkAi0L0nRsDrJC+R0ddFgkQvHsg
oOd03jAl7AGlng8XzuZwC+Wj0VsjydwL5bnvDMiKnyL8bvoSF8TtI5dV9fa7Esud97GLQrTUL7Uh
CU+nFa+KweeF4uOQ5vr+wF4JSdqpc29NJWINae3hu2nLEwQ324bBSmK+A2fNF39qvc2SkF4As+RK
iv9RhuHX2bZMH3C95DJZ7/62wD2D5YDweXcj+icTRkgSx40+BT4YGGPQNNfwS/n3atjdcgncRxEQ
Vjnva27bGANOW1wPET2mq29kznsm5phs8TkwwCllzsSVJHHpA3LC5RC8oP4hs5pBzE+f0fEykrBU
PooavAxFE527B9sHdwM8CObsfIThkivpP3V3saafAdvNSrWI12K46PCSWEhVcgZj1GLDJSeVqiMH
w83gVStLBCGCc7HTLqCzCbEspW2KPHdtjEUZtX/afhU6ShA0A3jzk4Y8/aZwvrjFt4Lj0waUUHLb
kNG2kERlioDTD6+MUFh9iMUPrmoP8/yvdw93T847JK8K25TPGjhCPYJPQnhFalFfiL9aEEigMHLc
DFgRnsAUmxZcUKSXIlAZw97SPy073b47A5SUYzyluVcK0IdCDBdmqMtm+ylhJY6AnrYtg5xPSBSW
pJZOKsW2+ASz1BZETFq02hsSrk5f83jnAFsnRzLgTL11qmC93eCmz9/N6etErhNNuR6RW4NYjKau
IZxTcp7Qi9ohUjE5o7SPRzb4Z0dUrk8EFDlYxIZ7N3WExRJXq0H3782TXvT59jWvuXXgDC0JpD0/
thhZGyFxDWdQUfVJ8B7r4iDEJE8PazcYBJ2vawt9tcXyrmmWzetF0xNst0amsvZ0ZB8NrumtW5AZ
ml2DzmqncAX6ZindZzIk/6RcvTB0n+Jhe0yOKmRQBKcarPftnR85dAojHTYqzM7crxHuRqqbzv7Q
Cs1Um4ZyNnDKd+qzCkzhLEyw2mZU5mZwHIziDHK+x9pcB9MuIKd58+JnTGCYDFdVKCx90I466YWY
5JS4SqWb99Dlw2OLhsb6SqRpJbtgwrKzIAI12gukVMl/d9GzBuhkYH8quHd97SHgu1cIrFjqTWmR
quV+CVhzImAXGM1NyAWpFqbkkggoI3iN38u6ftfe4EyCdPddRZC1E+u/GudpNVE75ooGKoQlqDhr
TMYPuGSx2B3Xq8kPnVa1ORv2oVj6vjJSrXZaFRTO+HKPnhZSe2LmWSbPbaFLiNsKPtY+dPZQfp2X
g4TlmNMRAxXQnvo1BdgTxv1NLtd/Nj+R+M12fTWlmtrmoBsDx7+ER9TIwUXLQ7ubzcU/5/D6Qk1B
33snNvGRZx9N2NaaU73t1Cweg2eUpzoP3ajcZafvbploh8/vghgQyanvByVRlC6ue4myR3h62/XZ
duLijZIVxhY9SEvSqsfyf/CkLBOizcD3VbD2JC1zawf653OPEjHSeH70YCW3Dx4R+hQYl7i1Jeyo
OthBJzg/cXXRE6+2JlZxQ6nFsOHbr1pCrE7KoYu6xXmgVWi2HotTWRPArpROI2HhtVXT3ygLFkB0
y7AgRiTvvNHOU/jbndEO4N0usscKqH+eJ/VyPBVIyfAx0vSEfS2jiPYuC7CyhtX5XFSrt926LuMW
zsxdTlgAPWF5YM3isjMnoKCfecKe9hqMu86egKAUFYq22fvYzXWCxkwhHW9ccFVV2ZlK4puq+Was
M0E9Z+ofY7L2k1fCMERWK+gGQwFsiS26YZ9XSj2QXG1ZrOtlOjRvVI4+h2uphWcHBEzCaiPZXJvR
T2VlgKqzzmw/3eFkcAK9vxao/5zcHpqiW6zuYBPZjpWVotvHvchwnRpPolacY+jnxQ8uA8DW5tXS
1eJ+PyXx8lwHq84Hoe76KlUrQFT2bOO6A5yVx3Ai+6YTywsEJUMrpdWzQRNnlSexch+J+lIJql7z
ZdVn0GAIUQATN0x0IXr/HKY4yiv2nuyjOwWGdLSeQROwpbjSrjvB0UYc6d4TLPcsBnx4FIhyKN0Z
DflidY71rhRxMSuQITPGnFtL+nVDWm4Xb9Hyb1JgEjCLBqDHhj4UjcjmPZfO912QuKksRfkGhPVC
gZud93ro5yI64ilIfzpD8Fa2Flduu2Z+PMW7f1vFcjwTGPWNdP6MP9CtMWR0DUblQbu1ym3pRLde
pMIKsV6RTFFZ/caaPHyLDC5K6lUd9PloobprUAV3eDaoIoNywh3pKfePea+7ipTmozWzaWG4L24q
tb4bLMH0hPtjH2l/H6wn2/wrlT7u1B+2PfO/W9YI84wHq2Ke6JAS2cjZgWfl6a730rUzifwD85QE
WR4ZHCdNChFwxQRS4ze1tDggcq3DSX/7ulcOB59m6RwDpnrsYLEzg1E924JRdcXwr+VYH/ETau4z
ruSNo/kl7L007Gtp/19t4LFdFIVPpZFZgHaicUuQHhg7hcZCQP1/ElIk8891pv4IgvM6twQOUqJ1
JoxHik72TrUVUFJvkU4uCopbRT9PRyc9sqvQLxhI9KzWm7545AXxlY72SHvTIx+7NxocCb0SbG+/
1ZtovlrmgBOKgwGh6+9IKSZDF8K38Z17B6DiWhjFxygR0ij6GELbiENMnlw259k1aDhGVpHGgRMw
5UNDj08l+ZZTwZo637yrnfP1FMAyEjurNdAlMhoC1c9id00jGLaMNgq1xwAsjeiEw/AVYTGyQOBN
we3nwTmqO2IJVKEoLDRsae1xINprc+IMRCWWqOddEnNYh9XxW9pmAtBRkk7+h20yy0ixMmfeuqci
Z7GvjQm7+1NzpmpUbPb9jyspejjJ8m13Do/HJBejlVy4qTaagg1LtQMKJozm/0cRotPom+8UczXx
Iv0oevRusSkEQ8UHUqm7EP5XguuFejQlUh/BDy5D/6prhzyaTqWnKA1HXHUYxB8Ds00LjmdxJYXI
UiJcjpkMBC8tSyaRTUjjwbEnJS20UmU/QSO8MvBy4jqGbmzA+8Zxwn2qhXgelDBhDpOqE41D3WCn
l3tvPYgdfRr3Efmfd6PC6WWVZby7gHFPAaPkZ+KzAiPXAyIvzowmVFDd6piVgW/BAHBsgT/XUrS1
w2jiyixzSl7Noi1wFcRICISn5vlEiMUOFNHIQDwUyKTrwOieK15XJct+kvlcrg9XBLbAHhBmqoy8
MiNt7drXo4Pnz58rfXj52d8wsl8Vmo1SpHgo9flzSMQU74fc5gr6e63c/abdulKt8jpHWXLOlmCa
/5ODnjh/a3Mg41KTOfJ9EY/Urrcnz38Kgx5o672r5BWOYSeC0iHSYPQmEF73OzrDfEigb/VGTknI
NExhDkEwLwgxsAE5/v/Th8JvpKsUerH3O+wRTmQhIG36UiYvpoOe2GHiss0tkdN+w42vHcp3YkRl
qFZdDjfYRB74Xbi51h0xEdBw6C6LYHhotk7HLLtZ5QnkiOPMUT4qOEg50tUrw1Y6sbOwIMVU6Nos
8Sjzb+SLNn7KbwugnEZovp4rL7oH7KptEo7T1TzYdBots5UMhc8itWm6Cut729OdaROU5bR+6fdS
3xSARoxFwA3l8b1/KAGc3gk1757X2f0lUwt01guZ8MsYfXSyPAO7tFbrTbU+kR97CAEFaCESwHa1
WwXCbgIylC/hnyM+ZUC6UrsIWP2aKJwiUQYirqOs4Sqjljmcm+H+dlqE4s4mu+A28glxdYstigKP
+lu/1GNdIlZffkh7rONXjBEvh5rXABPrMBY1HG0dOyGi73YRhXnmUyQJHgXfqKNnTbXam/6mV6lh
HEmCrLpMFLoozH5W5JIO6vHdkNl+loYYTWmTjbrYHReHOzojg+GAqIE4wQ8Myn3HXi1/vG/FT14Q
vvzg5oVcwxPrNOsuOVYlYw6aQqcdf15+TxitTthQST91IfiO5RlkLtT3AwiQQhkQhlWSOfWV0VZZ
wxp8WRMdEHyTOaZjE0aZlUXl2hhzcLL7XSQ/f73sNUrtEEc0E69X3snbqNdVdVFXGgvwevTVRvHP
SbwO3RPgOpkSZJ57XdUV5OHWtjZ4Jx+HCQJBYIk2G4wGlQHijcJPK7ZAMSvoynbZH2Nsd/Fh5FSv
E5akqPjiUdIoh5BQEsUkGxlhkq46x0YEFJijnCIVJz00jEXz9fIF+9k1mBiVHtgi7or9VhgfhbWO
DkBsUJP7ozD+xswYCZgpe7KMxL+YuNsz4w/b3oWYRthcWzkFjhbVcy6ibIm083yAe7yrLqakyP/E
OQ+9UjX4YpyG3crAxmfCYMiMpON3YFm706WMRnQa1AtePb7ZvoGhuf7z0g6Jp1yvfAK5tpta2Sgh
j3IvphLPtZGOtR0RcCJ7qHMk6ASmnqOx/p6BDmjChvfYaymS/x5z7Rqi6lWPXdXx+HpyIJKxAOVs
YTaIKnXtxklcgqhunBwmNhbo1FpFnPoot50VLGHRufR5zA0Qj5IkVfY96udYvEjsG/nQ2wRUNxhr
+kjtbKIHCNBNdLp9dVTG9LniE3LoNgcknyZLSaze6R+aLXjO3h9/slZEEn5C941MaiU0O994Prb7
IP1vFPVE1gq8rmuZrolzUwi2Z4sgG9uY8H216tJr5riwHoyAKiKHgKU3ZKjXpUL4+/wrBcTAFCHo
7ZDfe8Ko1nUxXQqT1wgBTMd+Mhvp7vYEtwEOf8jB4wqPXXbXiKhPNB4qSZ2JmHXXPXtOA92Q2xoZ
nLW1hgHbBYEo/Iy4UFhkfN9zPT3hLov+699RdqncDdvOvNSyCNlRVJ6VBAn8kIsbgftLJA/9wgk2
9VrhdyXCRYhFrL8GXri3z8uovA417Ne8rCDaPJIlpTCqfYKYQXF8fjUlTyoqzO16/1Fy2wb3akch
FotcCS8ys7Oi+yoNkMOZ/phOAi+7Q0o9/6HDyg1hq9mK7clDPgcoMoShk/KE0hZORyg3WCg2SZh3
xZjMEB7XnNt7mgcYqbM+comGrKi/+iN9mEeFfANUN1ED0vYvudD+73bY7LsY2j7gGYVpY7yK1fBT
C6zw4pn3Yb04c3lErUJn6ZvMaqdwh4BJIyHntCZDCz8RUQvcNey32USFcuyP8e1tOB3bBnU1keQE
BarrookIGCL+ulkmH19PfTXAsz8rZDgdot6me636VJ2CjFO0Fe/oE9SG6/GnBDlLSfJmuGBfVp7D
Tekw4YJ5SFO7zaRdCgVE6X7+z6b185qtjCYxVQt0pdjt5OsWKqpTCzwtKVaTSgcCrnWRNwV4FD//
uKK5bpsFlipzFUkd+LF/FtWTS7ELYo6bW7nu+kLuqvDoEIZICQHx4rhuLkJWS2f1DzOutL+6IjUc
yrdRvxJrzl6Kuzl1PvvqtQ9zDsoNobJLDT37oOHTdi+PE4cZw4XA1mV0y1Y26Tn6ls+Doj9Ura6s
KGhrH9pd5+mVP7zJGhYSHNOtasIdJ7C7+hTwRs1lOOqR
`protect end_protected
