--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
lguK6UkW0F2TjT744btiW7HjJxX4lnSS7uFDLDHyv9EO+a/JsyN9NaZlrxiKg5Q0ui+/52SXpQZX
aH9hbmTk/wznuNmhqwRNhzYh2SekIHIHGcd8yX0XXJMcm3FmiR5CIdMZGU2i/vDbAuy8AYSfgFo1
19c/rpESyYxpSrKqFvcLO/Zph8rMGgu+IvP+ZvlxWb7Rk8PHgdIGUrv80ijO18orRalSQKMblIO4
2r6pz5cf4yFq0f9/w4ferkeYrN2RgxDRun930DCdp8F+UPAj4Pjj/Lyu0sXBLkFma6MNEYg3OnCp
DP6b7CXlfe8yVbMRE0gShvP7gaco7f6jTb+lig==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="8E6brNnkLeqwfibAk59dL7adVHbeA8htOtszBRbePXo="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
sWB0m1lMhDeH5iNw2yfJyDwHpvpRis9mKY5+LHiXFL8tbVwaOiirXPur+QuPNovJ5+UbRn7h3kzm
YB2ZeDZU5xdK2NYsxH1y3tJ2Zu05rtIP5sSjoZdjQoobLNESTeToyOgkWyNMpPiwEDbYH9K4Fzjg
0gBBQqx1njLxhoMElabLBY6QIv1R656EBsGpvCWXKv47TY8GLXb55sXgqSIwIii+8boVQ625qUfa
gDUJ38NLmwRvLSBRSU28wfhQ/kCTGm+RP0nhU9ww/Jbaz19iz5VawF4HHK67iGlz1Vwm6xo+irBJ
HfowjbDDxSQ6H86mAO/47aP9h0Vea6Gufjo8Cg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="QdLinXTWuHGrW2QmV+rmwxcQDWByGFf6QeeRnm3HG48="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3824)
`protect data_block
BcL4+piRKZ4Ndoe05Qv+jFs+IZutD1CLXiXHO5d2jIiAdoQ42lgFur96jlOPvfdMVn3ph9zlFrU/
oSUYp5zRgDFAmBhOmXFNjtFgCrVLx/fo5iUS7C6AW9d9lKZp8zgZytgmpedJkmI/trJKd6jtAMkK
eLHJYx4vNGWm7n5BdxuD/Jno5byhF+5Ra30f24wqdE4/q5Pi/8kunGaYj9MqKhmyIMOZT5M8/lEp
xK5bKHHxyMZ8yV4jk3/2Z0jT0pCh161ii/92Z2XQE2ihCZkK2uyx76SL/CBZAOayOzmsTf6Is97c
dfqCNuE8grrJaxnBLFo5eAhpI2QVucoEZGeuwdeaiQef7q10LvaRW6DhlVp46JIYJAgrrnAfcolt
F+/TZoo6oUMUnbZU7QGIn+EycsNSB/Hkh27ATFDs8mBsOAfD8rmvl6ywZwye2CP4dRuDgFGK2hFM
G6m2w/gzrchBt28pXf+eqRPURW9sEyBZROIveSM/i9gCSZpzM3MB6iiDlcFUNBwknb8nORS1fgVF
Yj/q+i4h+GiLQxG8n4zURrRlAauDrElD6Mb9FqI//hp8oWXroc4GbDCkkIZXpq+aHI0Y2L4ZkJPa
hZlENAVRsXZ4FuRF0kuVjW01Nrx+PHfV86N6RlmaZvJ6nwqH06xdfDFh7XZOBwJvvYniqPXChNOQ
rtJTBunYvUQZA3F5L5EUjUa77kgKgpxg4HAI4+lJVVx6CrTi2IbpNhD5UqNCh/T9diI9rSlc1d+s
M4rZSCkIeSrI3tYfVYhju4z0qbTxi+4TrQcmJ5LO5hnxoxdjGiu3EpvmUrxI4BjbIbzb+JboPWSR
Qc3JfyAt3LDl6oYsxsd/n/u0KOK3qDK9Ms1FqFYNBk1sD+vGnPSvFFxVsyCTiyvHZKyBpPx0SmtP
fM9QHloPzA99KorCxGiLEXAw7yi7YX6kKqEwoKLsXJflf9dXCn/8BQiiEnDqWjZXTctu8OHVy4wJ
t5jePeAa5/3VEPWDaV3QLL2YqsWdkOaTzJCpOZifhx9Ivc6PCLdA51HoBsdARXjhdM5hPte67wwW
V35bhSTZ8H+WcpAM2iDLI+X3lwJ2fFOrAIWKwA05nBfgJ8HrUF/5rWbhGV6Fmyaraf7MRTzz4Y76
kfd5D9qV5Bs9nA4dq5oRam9TUf7SXhXoJC8SzI6mpahPJsST92f/aZsZu+oq8pFmYsrUysQ0SLj2
PFSfJHoQ0p5x9h1lUJdHTq0QeNnJ3IArpBYDw2zIVpFE2P/Py5u0JMv+Ct15XkKMjwdL99wzAl5B
WgN90gek0DJCPOX3tBgamaLZvf3BXYvUm0Wz7NIVkqM4fWMHDCKuayouua2Adqv6+KTbHW4TuEbZ
aXA0Tjbw/n9XF2aieUmfgm0MRXBP2Fnm1dD0yi35Xm6oXvXM6n67KtJG2AxjXOyC6M4seWmJ9DFG
7FjesTazqFEYtcodUZrVins7jqmiIeJAhl+IICVCNb8keNHw/b8zO9rJkdbtZ/i9pAllPhFkfZNF
gHItr2B5Lx5fcu5L91zxzsVPAsu/qjxND9nkGFZVcWTzyOmKmaYWQ7jE4+BISX4+KX4tUxtYCWS3
iXx+J8/1MBsNFd43Ig/XFJ0mR9Zt86qBsNr2QmHTUB1s7rLsUNWcB/OoY0YAXlBtEPlflKSFmPfh
PtQmIA5ROsjGcp8oSG6hkMUy66tj7ettqDErm7URMzirgnm1+8fXKMbp7qz2B/OigRtCNFjJmN6F
em9s1Ua4W/mrwSpT5vaZgrj0f7CvXjRHLu+xOneTbonzXd1QOjWGzA/BowWfmckgjfvZAEQvVwW5
sCY7PiXA7cjdbznz4MlrLcAMkv39NIbANMWhWO+vrai3zp5710Gy+pCZXOe4U5yDtuXZfWAzlhSZ
cCIcaAAxB6XVbDZHOlC3vzmOhkaO14Eu8ceoCO/lt9UBU1jtu4OHJ+RnjRyvKz6DNPAqfSwff7xd
LFyXC9JTbyXryfoSIzSrRZj0P07whkyxpbQuPjoymXRZ9mT9mylCX6T1ymQ5u/XY/kUKFVfCUgkm
5gKoAwXiL9J5r477pK9z8791HMjaaSzM3TrwgmjPDnZZXlB7bbwAGwB3wxJuE4OqV/aGJQqeQBs4
0FjhJR6HY/77eltS5l50DRURPjT3BOLpP1thnAli5tLCt4YeSVCwC+Cgz4x0Cs3aQllmBJpWmgjl
UHDiy2Ohx6uldxLzQxvLB88ha47aB/XzqhTxUpfKKzCBRYfOx+ZGSkKzyuNfUx6g5TKneKQOs1b2
MLNhoqQXyyqymrvugvzz+JNgLZ8lKWvTrx+s6KfHtG53rGxMEpzYPOSHMph81yfQURXQO8xdhERx
IRbvk/FPwl8+EgfgcICa+mfvrHfVzibSBYGRddVJuLDXH1+eBxR3Mk9V9kbxK6udcE0CJGQqEa3d
Y840tqkTErMOfFzDFCc/G7pS4DSURF0/3uY3rfwYYdCVe21Ffu4eTdM0DEYUa4Nt25dKDIZ0Y//Z
VK2fpxFVlKi7O42gtRatlwcP7HQvZKJdUEvoPwypIdparkYV62LwX3pE8fnkK1a9amQXfLrtFOF1
NmwZJ+6MIFtcchUz6ssgATsvPN1sA3Gdy3kFczVpf5Py6uvYoyJTEBqbv0GykQLhvMbO2vzaynXI
TEuptZkQ+RvRCogNpOA9EUY8EUnVozmyeA++7uQ3qR8S2Vqnd6V10+aUcQ/ROhidmtjlVHhfRMQF
ZzYHNeeRRXHMQ8AoWqic41QHsLtiJM//jLetyYpH08JYrg27QfWLe0qPFmqxfN9YyJfe0iwJwtfH
5U/atf9aWkHynFL1Jz6H+xewfNZKfhnwVQqIgBKvjdvk+fBbRf59nfwPBfFL36HYwQHjj5pMw7h/
LuXSlLLjiiB/pV0yfuHJjLfL1Hk35Gro/EGjEgonIami2VIkc3uwGtXn6fvqwysFhi2U/GPYvXtv
pVP4WKSmqjsxOacXcd4YWCzIOhZUupb27P+VsbQZvAyJk5CWhkzCEq1A9ssq96LLUubMwZRSQ078
WOtmyQdMAM0cgCJRJbLZZWDocrV/1BT82WEujYvrUFYoTPRb6oHdQ8IyIE4RKfFiOQuZD9dKSuJ5
d9xtVHIFFlS7g6y91WHEmH1Z12rLDMnhXNIEQiRl0ZXdqwwQ6DUsIpQxDSj0OJMq6KRBPQ5FviIi
nrHBoc2lEP4bfr1uslnaUFoTk5iZ8eWgKqiS2RHagE1x2ie7QcU7jihnkljRX5teP8V6iC5fq6ku
A2rm20KcvHTQfhaxWn2omvGotNuiCm2IlQxm8jIYigy74MZat/ZBx+b/V/VzCaC3+oSd825glOeb
VBJu0bEWYeAgjJfNMYDHno3dgfdOuVYEUiofla9qSUDVaNdmkVoYdK8bM2Ri4hi1FqTzjZW2vJM9
/3CHC3H1oNs21xRoZFWWdA8I3k9aQopijMwcMUaxsz1GgHvGYbGIZG75Ju9M1ljH7CE1pbhtkuy/
BaEYSf4YC7eKDtfIt9H+uBWb21OpgvZzG55CSxjW7qGPjGhtuBmh6dfyu9PZnS4P3cu7zRmzDxRS
avpdiKesU1jhmopCpaqnoDoVWyATlzE3YtQ/ltt+81+AUc6RVLgaHJxVZ7R5vNCm4wfFzbOhn088
EOKgDcD9kPTK5KR1e3ge82W0RMmtuKN28FonD6jVFy1Soq8yXTGaRdEb77FSdCVqMZkF+4pgPGBb
JcB+orYMRkPgo5FkuAY6xIZAxu0mSY1I6y0w5XSL3qASwFBeyu269ZAJ7ANL1DjbN3tKDYE7lzcw
dXNriE0ocGqUkB04Vl5bxrTrZD3E3/nPFQuG9OpzX0idtBnvSG7o/fbtE7gF61OTERgezwxEGSNP
1iTXcm3uWrTeW5EMiNH6dcowIz2FiVzG7pY5xKBmO+Yq0mkLPlGhCcFAL16A6oSLvS7ilaFf4phj
ugppoK4RDWOBQUHUGFj64Aj51/TuAMN7ymJ2kNEx17shq4t+nkWSgjEvoFXu2iZG8lyIzFaIFl3+
iKXMEInrHpSPmsUvtmVPOQ3nRl/YvoETQdkOJfOtf775GcMeo6TehqMfDe6lzDkLG4A5DUV4G0HS
CEu57pvaLOc6SWwTtI9byN1nXOG4/jKGkjlyig7lrUfsq9K0R0jqJlE3jppH4jxTFaUlGQxRVOet
Q2WtBZoQ280I6a3Jd9dPEcoKAB/p6mikAmRcXxXAALt5qt54di8UJ1Wz7+yuMtya8FWTS0MFU0/u
8E0gbJo0RVhdxDzFErRmObln7SCNXD71TBnfio3FnO+NJZUhWDW01TqEAW5RVLb8vM8mmdCisKAQ
cI6chI7gytn6IWgqu5cOGVTZ18FN/0WT4LJFrWokM0lALLEPxGHaV68qUqn/JhuAqjEPSrVcRPW7
VT0hBfS/kKeGeJpoiK40qQnaadIvT4UXpiUWRQ0DArHWUaOewPaJfGtL3F8HkaSEME3ZNHoSvTCg
tjxHQxbSj+VHFbgDIl8V58/Zqs+yjYPSgRQTpt+XcRGTJZgbqUxQuyrey50EBZTC5Hb2U1HFoBER
215VNh2wIdp+X4sWq0uM/L8+RVkias0/HRMM4ikh9miCp8h4wfaM1S8jGEZaaYne9At1/YYhPkFo
HvGv0e9WFWaw0LIxJsYZY8nHdkbD1dgQGsBa9lmUuaSL15fg0iN6jzBbWQBC6VStPkPrTI+H5LQ4
Mcz/N1L6+/9YckwcJm2XTKEqBA1/teRQLVIwWF62HLi5CPxWxHVSAsFJ9gsjkgPgcjepl2yeJVKW
o5BaAu4nRt0kgY96HKSMBySNA1JYXA98kGoIC4q1snr9M41b/ySHF8+4gP2Dr7XpkQo9Y3UBuoUO
qylrJk3nVr/Z4JHwneLRN5p8pwfB7UVcPA3WjSmvgLZHdjco3lNzeiU0BquCb5+tZ/mZwgdipDkt
xD43JOZ7lZWtJBVl07X+KQdNIz9xpmDLaJl6pfVdsi7zvSHQmfeAGaQh+ZAX2prcs+GWQywM/2hH
vUUWTMHj+7OFbI4hE5QvvYCDm7uKtn2Cws5N8arCDGDWxp8NUsiTmDbMRtGZDK8/M8buS9unGjfW
HzLxy6Q=
`protect end_protected
