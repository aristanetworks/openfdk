--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
RvgB/t4y4fVkPzoTRrM22x1KQqeVBTYuM00/6GBC8Fb8WrFq0N2w5J+jRi+OcQAzY2Hh973CmtN/
b9lAT/6I6WvDMm0Y94Fh6Z5EqmIBD1Wsdl1meO3HLnb0IEz0P0ieDaqoH2zF5T/U6BNMBdw/Qe9w
dxEdZMUr8xwzHMOyITtnjXhqjAchBmw1QjgGv5POj67y+eElP7a8EhQpho3UeaHTnP7MhbM1QHhr
ffVngh9Cv/Lc/sgLNmHdx31f6giBQVmKPzTHwym+DANmFyPUJ5wcSoaHnuMTXG89gGkew2erbyI5
5VnpytBHUgr73H4Ec8ZosZF6R4u+TnchalgP/g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="+EMFR15Jf3yA1IvF87CQ1IkPh3mast602F1/yHM6bhM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
KgNGkj11jy6EMkq9eyDMZBqZeUDhB3pBMkhdo3CtWzW1i062HBcYRebdQpHlvhjRMRgRsWk+waIn
Fnho/HJS3/h2RCchiQCKr7klt6AGVztyQzJrCbKDjIsL0c5cM9MEABmhxznXVD4LFlITGMMIteIr
sjawTQB8pT7cMojUGsljsKEYK8h87wjU8E5kd9OGEg1zEyaxyAzfjYGKHUW7UThnLrnz4O0U/RWg
Frur+OEJbC5Vn66WPZ1spbBSeXMLkyzRd06NHXTJRauXMdj/0KA4RV7cb+FlWfIdJIoFm93TX2+5
JsUQdUINCokiSQ13prcmV9LJxzTVkC/U7uKQdQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="LzTOfmIL8j2eYNaVGdI6+jjquwN4qvMr0oNxteaDP6M="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4480)
`protect data_block
cpzkOvJ/dFIGYYCVauuIstirydwHPL97kaUZgFq4lWMgsiNcB2Gt5L6bgeeEgiD/s0qP6YOmLL7u
1BNZwp9wfKuIfLA4/jrBiDb5nsADdGH58FWzgpT7D4jVdyttCuKKMcXWvs30lnPorK+3lw4PIute
b8Zu3dvPmUuqj/jNRbQJA6cVZOoefgFU8X021CeAAqrgId6Ku3OTYgeTi8NfysJ2Yfhsq6xKZGv4
b8/rSBV44IGxZGYjHZ60qqoLDYh6NzYQRV4nKSafKOloPBw/+Mvlbiv1B+ubkfbHWJcZ81UY0eja
koZZOMefaNOPCuLq/G00J6rwqawD/Fbq4AZK2SYPK4dpEU/vh+D8wvrImchvOIFeqVEGjyqGH4tF
AuvaJckzv7VxqCrjQkpw4FSDwKwW2zDKc0iMYLCANos3tRT9LbErs+VB5EWp1K4plRwl7ijc+cj4
rtujcZIm97bySSYAyVt5BvWG5fpuSrmnV30KQjfrP4EUw1ghMID4aBMkuIeOzlGdY54ETKKfIAet
idzIj1yCLSQedHgrLCqBjur56U1LJl9fI6wKOleo3q7DbnZeXtQ6DjdiPZBj/sGOBXY6L5Q+xeUM
/ZFjtzNuaaGMko+lDdNWC1XxJexGw9qjAQJ//CKJcJqX6w5jFwHANQ2i7DHofatblEdgHJseKHk1
qwjAtc5dic/gv/7DYbZBkKl9EQM6GvWoOAMxr73BpTUhE5UhuLTL92dD9iwAyVGy8vYTnRvtqQiq
uLI7fpUdT5lvsEB1v+hHswqcq6nso3u7WeWHpkizPgisLZ8vmN1E31kA4ujIL0ibIb7LUtXj1tov
KjEVG6QCa08mJ+CHYi2zOr88lbaU6vwt2ukd/wKU1S4jEL40ou8K9e4Ed2RcrOo3Z3M0NeWasO2x
GEFVw/iuKubiG2L+DZ4CUhcvPK+DGk0jbLxElelcXyE2ZeCls60RdhC2RERqdoSUJCQk/eW/PILb
Uy0E6OWYZSS1EfYcXfg+C90EsTBkPhM12l7vnylQMbUlGbMIsbYRq18Fa+0xae+TawQgFxdq5J6E
f+XjefGxJ6CpqRIPRJ/tcbnz02i/aZe+VmdUm18a7Ox8sLRLeWY/PtgKi9Bjt9V97ViQ7+K6KQfc
CHCZMP+iq2bhfbHy3sws6cxWpUNn87pEqcbQRPPaGWWgyOMaFr8i5EIJYKP0g0YHa7EGsoanLhjO
I2aDpdmwYACdVeXyJYTd9dWl0wCYBBMpxS3eIdaN0iIEF55GpzGvEMuwl7Mkh/a06K72mMoBZrqf
j4kx0Pj7jhGvJ+U63hyxY+JCqg7/ypvWGXye0Rc50338zsieLnLf3ynBNZpAPg5C87nuahCfzvAF
0Mae0IJZspqjaJ9dUL1OMIWWOC7CU7P13/2aO8b3Fie6rKOVKpHYq2sxw5vZZBJ/EzPjkWslxp1P
qt4vYrGvL9JQ/s7u6aowWJZOKN+l5Dwk8G7A/LXiJNZaYQ5JnAkSCIB9Zc2/9ruIRxKwq4wZhCtz
a578jFi00XC4QqYZS0lzqM6m9l85hx1k+DFFk+U8EKyi39YbmtIsRdKI8PS4vizTNFLg3Nnwnl7M
+8CjFtfOlPXXG1B84PZ/h6P8l5BBsuGKBveRw9BzzHj5IaOYgAYswkVPAFYC9P6oOmYccZ+kk98f
Aqt875nix/TXqQEmaitySqFQdQJKXbMKt7dMpyvA2rVKv4Y7QbQaX4h0XXdcS+gS6W4Da/gQBTia
l6nL9C8PuyOl/F2IvI+pXC1IcfO0d6gB/46Evmoel4bXTwrBk8HnB4/mhPwjl0lIHwbAAZ0zh20J
tlnqdHQN85OSWzDafXcSsLyBRTXyMFLR/KrnqRrXNCDcQQSnDjZZSNZ/Rinv3yLs7CbO4jFhEI1v
+t4TRvdj+G/+uGKhGcG3WAuDVg5DMLBdf0ttjuwbFS9Bn9+ESHLmaT+Euy3/fMn+tSkhv5YwA8Lm
gW9ZlYfwEnbX8nzjzv7vC/7DX8o617T5EeCjMqrC+Ov2/LknNMH02etAeRUPPDrrFy17CyPHMxsI
BKTEFl4/RCrUuhGWwyHAeMPqMwj7M21gYOCURByMwLd1aPAfwOYyXn6IQvzo3b7LgFoCwzzzAMcd
4E65gkjgmZb755N0k9YTZHN4PzWhRPObJY3VADwdYxL8c9llFm9qAXTjCE3AWxd2UX29+7WiHgFA
lNZ4seyc6kB5UeXQ9bNAbmgUONDh6iTZ6bwMf4MgWATlSx56h0RXBizuC4maUG6q9KdfXHrkq/hm
T1pIEcDMlXHG65uL0fxlYpl12WXwjB0plJ4kfV+j0FzR3ZWKoxMKqsX3XrDrXwHxwXxv4Md5j1t1
mrAorplf0kTPF+DvBOhBc1mRFkpqvkSbWzE/ORDxnTue1cdDmbx1IotQ4y8PYqhOMSqLD5ke+tE9
s+ngyfBbAChb3JDNx4wtYM7zb5Muy2w4D5T+sWaK08NyvtoTtWzHkZwlVzd6l++uJSG2hT7Ybi+P
KtFFjZKSBWuYc9lyN1ojyqXDRU+jc356Zmqd1Y9Vm3PoOp7nc0bMYKh8yB0AhFM07LhfsYnMHplj
r9bbA14UuggS+QndwZ48EUBZY2KoPlKb5yJ3wXq+GWBfb5bxSv9tmiZdS5ysL6sou2g6rT6wWUCR
Pp2ON+Zc2gXjBXnWrrI2RhRK9qyERFUClq9oh+CeG44aLcF6jfXcPX2hPXVSX2U4ulNm3BnLiPpx
cJ1fXwTNFiUoEcv85PL14WkBCQ2wz5dtKE6WTAmYLzlJ5dkMPCPwQNZsxf+p4SZqwgZZ2s4PzUjk
7aBnBWKt/9R2PY+ZP8juJ8mjvNeSIfueSJU89ojO4ZgdaD1Te+UDVT5uYYMAK19Vzpm0lzpbmX3+
P5btPA8GyUhh0yqF5H0Un70U0c7Wr9JxqgduvGxb6JF8jO6sAyTvu0lsY+KvkgKxOgd6og2RJO2h
rGe7kpAe4xTQkdANsJQWd0NL9wC7AHSUKIKbLiRIJHXAjGPUZtB2xhxA6RG2qCc6IxP9Ryo8Txz/
vEoso41EEtGa56kSaTpPeLkEUaEHIlzlHQ9yGJjZs0qyZaULxY9XHClZM/tpDVv7DjWtLhURKhHs
By9Kt04S1Vu6VTnb8HvuKgEe2FeLqu6a6eMwz0S/LF9z7ASlg6nChgAM6huRQgd2mWhCDztlbsoB
bIsDngCOWB0n4m65ZrAdEN7e48qQosWiZ52rGnoCKiRKaYVSXSetwRLlkQebnB4Iz+g8RkJWXOAb
W/095HE+vu7DVkSQdlhu3Sd5QSSk4zjYLSOwpZ6I1bQ7n0CJqV5DyEo5Uz+uYXpMm+Ab4rlOWzuO
t+q4fY4Eqtxu/p8UPdIjh/uGHLxxandSIKUni8G9cQoPsRYfQi4xe9m/42tSz+9HZZu0CRqxFZGE
nKFfDp5ykevhnrKzuX5Pme63Ipku9Oem1DTFC5mY9r1e+vxn3+R5/jMIa7+7MWiy0R1K6fZLMFdK
xK/EyFCB14zV3WgKCs15aT8rJRB3oYEISV0hT/vXbsuEaTIHXfEHL8xhvoRygWNYiCVW0DmitOf6
b0HFW33ABXLDLtaXop+326nW71CnE79ZeXdKZ7S6gk9ta72yCQqVEz39BeV48jTaUFTf26VRnUqg
xriSVYaognT1nbqq687RxMNAnXYbvBj8T6ATEv5dqaNUFy+g2X4wL9+bTLJ8J/YCWYcVzhGX5HDA
tq+SXbcU4Cesbu3D+RNRx9Yib/D4JxcOD6tUDeSnuck3auglDd91uzqnIXsPidkGUrRwraUm39+f
RWHhlFV6Bf5CTf+6flzQiMYxjcYZVuOsl1YcQmV7Twk88sZ1tqYc4GVEekWIhz5eA7/H7mJfbRUq
GSun1pZZYR3HA6NsYlYYHegZZXrwSAOReMJ5taTBY6l7t8HYVDhodOrtXSXgZ9c9AIeoZMBjhR+d
xzrL8nDF3qWtMGyVRCOhlBIofbn1ymV3799Et7o0LKxGseLzKakb+ANyPAu2BRgNOI44n8rpupU9
GoV7FaLNgNMZRb0JhPUau9SX63HlknHJb0Z2sYTjcpatQlHbMvncMYoTNxBW9os52lZY6jAj/D1E
P/5gjTWOROx38ky/A9RAI0VReMvv3VpT0DiFcD6g00bDtmtFAGvM47JGgmUBXgMDnx3LyDjPZiFf
zYjTZUuN+TJc6VsSkgyqo5hbN+oW7yHrvEtvMjTe+/gGLQyHAI04ulN0KxQXZtn4seVsWOmbtFdk
AnqurHGXr2vNo3SY6JeFrez1GlDR18PmZS9K9f0EhMWT3Kqz8U3tHL7jsE9iEb6JUWj5qbO0kegh
56774EJiZ+XrkCNLfLKBapX7wkDbJW+5iBJ36RF2BWB98E8tB9rl4uCFtuKZ5IUwsXIk33ZpYYhf
AmO4zq08ZHEg0kqSi7YgAK8/mstVtY0ROXRuifCR0ozLiFi/LSNml3vRjrGRXgqOINesz87QAk3m
Wsekvh7FMbURdyrds4B9wdJzcxE1aEwKNEGqGKca8H80xGuFiwvV9Cvh5XIa5Sr6piT+pgNGRwsE
kieISCAHh2ArNqLH43gAfmFlECisYvQx0t2Ng/03N5GpRLGOFZxA6ka/eZUtXjaHhse6Safb5gpD
newisanG2dnaAp2XwwenmEg5WF/VBfGuG8NybCyHIs5aRKRsQw5dwXRlVvJgVLph75L7r/2a/0Vk
6VR79Tm0n35+h9LozIeIPjekdWXNn/j0XZxKZhrKqWjvA6WyQEuYM6JfqYeuGK1I7tIXWZfnVsX2
zJjPx7JjKrc/x7iYXSgMb1FVQlAr/ngEdHL0XSqLIdHvaryXFSzaPNBqlmY0wDuyVSJTLUvWFMt9
63U6EeYgFAzbOy3FAhSy+TyVeNmIX0gxtKzAsAkqKHWIy+A6DmVUndZ9ayMMLd1MFIDBfu4/cpMB
0GU2e6wTCyo71JzMPQB/VARGLfA4Kuho6kw7vu1BU3lLQqHDqshDQAk+CyouGc8knWXLnBu/UpmD
k3YxiTrMYYTdRMrSxf5jFBRuuFxi20D2aJulTBqt4vnuzLW5K1KDi3cDoSqYXAxNEz1SKeSvGMBE
batv7qpgrWLgXdOo8ljR+Q8dLT8bG8RCt3LT+waQUaSyvWOk1VYNjV8jHKsYTyp8SQHHGl0FWdcw
e+w9Gp4ofOQCS101m48yRCnuoffpaJNZqWM7Kg/T8RwiwoWjj25CXvhwuW8xfLsbhQujwOvpCoSR
tV0AohXDkJNSnHQ01rxCICVUcZjhB0wjZZky+G5OIjY9J1KSB1WAGxAcnzfAHtCDh4cRryg4RKT9
iVu4SoefED6ewXWlINliX2cGcHgUE9yoo5qupYHNpHBJU3eiaZ9OD2jdDQi2si4ODlWV5JnOmVOv
WJkYXN3U9jdtXQ7XyEa5/s5Y0TIJ2JCTcVjNck/eZ0u98ffC3TycRjGFCVePh8gI6pk9Sn4dvI6N
AXf+XNiOBqE6fxnZEp/AIWXe/TsxoHOdfUMtZK8rNOHRIMK/yOBgJQSuoNa1ZuoiJbKQjLPE0RJ7
WXteCyq3+BuRPaNobPdYn6mUEQd68O6JeI61wugT8/Miv8GRHDdPmPn5sjnR34+BQks0kYSVbXqi
ipB6fRcg0zVZ/yRFXjwBzNHqHV3imx/iZtyPXPte1pit9DAX9pfOE3GrNqEn2Oa1sWysW98O1mWa
yZi9voRz2qiSoPoVWsNj7tU/kDJB5RczG2r+wdRbOJNnxUD/QiOjBBOR7qVUn+W4mQk5NasGLYXT
RFFLgysavzn2Q5DlzRTu4sTMG5PTJAUP1K/IlMgOm26rkHvhqYzoMrcE7ltXoChKJNp51ADdrgdT
LAKFcGWDkk3zpygbJwGThhdwI9HHxxeJT0wtK1p1siILjAOxHnnu4aVWDhmxyr358htB81TsZhzf
5Mqo71A+Lrc9QKRgScxquPpwDRQJdk/CTkKcLj3N3cggyA==
`protect end_protected
