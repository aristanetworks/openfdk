--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
BUoL4ccYaMO4bsYq4WkJouRFdl5gDzRhLKp/jHl5TQ44S+jeDDf01a2kAkmbqB+GxyRFlhhZ1+Fg
Onu/RzB8DDGZgU9o24anqniOmh4pszgbfTZarsh9/eFye3qodkCDKj7TFLWVCYiZQtXC196LEokX
V5p1s0oLfGb2fegDFMUi8z+xp4g3mtHA0zt7/u5HWVYQF6C2qY8/9SSNzHGlYcLsDa9ICEX0o/tt
NfkFNt1Lg8Q6Fopz341R1tb4d+GdA4RaaBjhUZ3TfQcGHhZDLIOtJBqLi6W+RYNdQxuWz5dW4dQZ
klxRGZctZMUZpEYc5yOZ1W1NuWF1iaCujGKpSA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="0gVUmUsAhZfmjmHw3iQSuFYOP1VPdkg849rX6P1G7Pk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
pF7XylsAlfNxJ1AlIO5GS5sGRpPDKvLo3EE1Guw5PNwROZwmWWU9GjSJsbAKW5ZxoYvbNjzBqwUz
z11B8B1vT8SsPJdagvH4Eb75XuQwqbYBcg7omjd9wBHToKYsgJczzoNCCnGhKkv7j33VE1W3teFR
+gAhy+xy7tdj5pXd4k1XzifRcMEd0FQBxkGFmC9WNgFeKPfpUpNc/Nczisazl0lBTH129yenLU7P
DwyJfD2wSypNbSufCmh0M4tMAXDR7gKRMBUvD3713leVlU47Se385dzNTzkElevpuzTCLaauchAf
3P+hb8LFgphlQ5oqaHk7pB9WTtqcqusGiLMuxw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="4cwU/iHXrIfYdi7srtzp+SA8YL83fcGajCvA7KwTofQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6640)
`protect data_block
5qBTcRhykY+TzCTjn7/lHD0MmcaOuWCVqwnkAPQQ7iI8c9OV9Tb95E/mQODNYH3CW2rNM+2PfqVp
GxqcvbPpc2/1ltwlUd6wFHV0l0MDNsixQhbrj44nfoTsBSFjUVqk0l6+ZqOzrKfs4YEj7/2xAilQ
5AnSaYkG0hzZWI0n9sLbECg9kIKdg3akKGAA3Ov70Jb7WBqAyfNJQoXsS4dSd3zdBy4eQ7opcaNl
setLOSfiVw4DydpgqJNGA3M06J+gB4d6ikr/uc3XnZCup2QkI1XVbyRUCdilcKza1ZCpSIUTW+qI
WB6J9PK3w1QMaiwvkFjd8dJ3d3l7osLgmsRks02tZsKufvIRnR9pG93Y7lnVGKZK5y9iY57UhSRw
xzBjFCHndszDaKFMyV/S1jHThNLAgFSj4iuQFS2j9ECw0uAL79GzNJ7MUj8D+WnBA750TeG8rDca
lWoAB3MUdY+jDDPbgYKgb/0mqqxsPKCRJXjnEUfTNsqeDLdJOrh/ZvHGABAdSOroc0VtcdhZL/Ar
Pv7vS4rOlnwj0IZko4iomux157Ee7/QVb4dkgVE+RFwRxVIa79yrlgALYPsWmJksv8mkyydKZOve
9ojiwgZ/jzsl83sV6Waur4GCQkHXRtr8+CPL//qckMZPXLLcEBKF8NCyl1Pt50MqTDV5vUgG7EI5
Z3ZMZJGb0LNXxMY8UImuvF/rC7ksvGQ2zLsNP8QzZiCyxm2PAFejxBpt7LM3leW8YmUfN0nb6/zy
nqQX4RyN5r98SzbUFHl5RjWXdm2HvG1TuUUSELWE3Uh9cITVcYdL+ORdoVNxuxLdM3rDRjaJuXYp
vfQejQlVEOYs0U1mr4vc2iTVgmWuxk2Lsj/POGLH395YLeIuQ7VI4sJA7JIWTB71a8GjlXYkYiL+
qxqcAxWoD//mcNJrUddRtc0e9kjVIZMeO5t0O+UZd5urrblkS0KFHJP2016lj4l/WHuCoXT/iNoc
b6Zo2ySiopn8LQYdocB/mlQNdAj7/nLkQUjELVXxOJmdgXomILtIrfZsUK1wfJ7nPNKG3pXAiP6n
SYNIciD4o6nskfJhZsKJN7Pt4ogb/9otmw26iDKqieTUOvaxceuZ1hrTCW8FBSjgeNtVL+SS7XSq
9/g/gC16F5462XA74e0t+JyyCUKjgPBYKTtoOzDuAUcO5NlYzszs8qcAFciU3Tt5ghJq4Ey0IyGw
rs5mbhRBQC0vL9F4D+dFtKty0mtq1DEsJk9wuPzwFnr2RhKsSMqBbovMa04+EccGpNLs5p7mTbFt
8OEEvhH9f86qKayalETGHJ+cniFCyViIjgTrLewiNJ5/9vgC7mPMDVQCVzMqySfEnVlqRWIs334H
uGbnOyW3VizmOTiBvckhkpCcqF5sqxj3k6nhrbfgPYzoJGlV+gLow0XfkOw4lhJOWzXfeEQ/xlWr
tfJv8P6pe72gcsczGTjNWYKRe2zPGTexJf4+uevRqwC71yDE7Ulc7rwaonk7Pjzt5NuFIdss2264
XXYKrOWtvXENk4fPKI7pm+dYAbbbYtiTRoJMbIXbQqdxW0GadNjDC30jU4KJHSZg9HbLyGcVM3xc
Zp2sxH1+JuJ0HClmbOyoDORyaW6+f81iWqXGWAjxtSEf6X+LAXIunOtWpbWb6SopufIsfpL4RLGU
faEeWLFNODPaNlUsAsrqdqVmXM/rzVJ9Ack5Z0TRIDbTs2y1ypNuK5LpYx4sI8cDL+HToKBKTOCr
hDB3123aRcC467zQbM5A1pzGdr7pO5BjcoI4Zy1UYbhbCn1+KwiDXvnPZQfFt+4xYobszM/3kbFI
B3/4t0QHLgFdZrh9KcgSe9gu4dMahHiLuHQ+qy/mlsUn7NwbjQc/Nl5K1p4XS0ZITrMTK+/DbZyj
Uwz4fQKzdFbmKjHHfVWQ3l5uYDdw9GGB6+e+2GMyZwcUnG8gIGc9j4njQPNsMiuxx4406PnLL2vy
em02EuhHoIp2NzjxShp8GL1KfZYWmMxbLOvVlmKfIcDwUR67LrmGIkFheGLNToFxNRYsjWDTemlv
dwzNchO8qu+i69smjx4/M+9A+qlibWU8SgwiJEjpg91E6QT4mi6aWKwdhG8i2O5tIbo423jCiRcu
cVj1xIiwyzzyToL54IzIM/9DEZVVx49efX08Mq//sp20UBG8RJCk7ABS2sd7Ke6+AAAfa4HBUcbB
w3DIPx0z+oMpAJmryI3aMlaWoa0a80rjP5jXuwg3t/8ynpJAexI3KySXXeooRmd40IUexgJqOQWu
cCgqFB9dPJtLsfawHm5xbgDIw4Dx0BqmJTM31quHggXQeoxxRMy87hobHLPv34HYUr8stVAY26eE
emNlojpk7hhxufbN6FzaQVn0cG3RzSMGTg0gpDYXn2DKZq5vaujWXKspiUntIu5+zyEw8eOnDnSc
drRn0dox+V7cumGksfFbBG/OGh0mDYttlVyB+TWNUZqpAktBp4C7WPgpggEHZKMvPEzHNQkJlNLx
+hfC0Gv8O53bQTGss3CLWBSoVhM/X8TQdmgp/81+7xG5O1yYHwtAXJcQrsqQa6+GImXdkOcEoulW
+02BonYOMRyuqRawTMo5EsPbbD4FFM6h0f0pr6SJHyPQ9t4WFrmKIqIocBSx2kCPcZ161Gn73gPS
vNgwFTVgilTH06m3HV9Sa1wG3kWQQsuSvjPl5epM3dDoGmA3K+yPu6dGkk/Mlc2YcLqDlysqVdZJ
Tdj8h3iY3Uxp38aeJ8qMt8rpYhFsyNmfm14Gi9vHsij2rjMY5TlOUEuvNXdSJKN3BEyM+p0j7G3q
WSxjgreuLr/TGrVZrLIyR+zhy/+pTN5Wq4CE6zVHgLjAcgo8suDFHrl//9dcqrRFtfML1oYDCN4+
uhmiugHPA74NN1xGL30BNWt2CjnYFG7X2s5B4/ow3Zdw4Im9bQ4eIudud/wMbjL7xihBeqnjuwfb
qybWWDY8pC/XXSpc76r8ze2dwzeCG4dLSjAxJBIWqoRub+uXaMatFHT589wGK2FeyBcZ5DGMd8n0
3de/FKxTRgmUQrg9Y52oXCNIUgULvhiLFx59VzvNrixxqbV3GxZgNIt5BSkhB6Z5sLkgS6Xr+uXs
erz7gH4/hnmfG95ImwLbaei7JX4T7MHCo3l9W/wZs9r2lEgQY4/WbsPuIyfq46WTai1sZuTdgnkt
NYNjPrlRDPbSTPwVQWLjanAZQUDWUtNor1ygaUARXIWwqrlYniUt8NZfwq6UIlIuTCppb7ouCTzT
Q/WLdpJCST1PHj6fyiGEgivedaUwXBkxpZPfZoeE90glnkd8lVo9iqcxTjSDdOm0G+3eaxGwMf84
OWJn8DYFIpGj2WCP86lG/5mqdWKfTjdXM2vDY84hGr09RDtR/GDSZXFzziyNjtdntR/StQOq4vEY
6LNpE1BttfXMxkBc0ImdHYb+87XYD55lEvZOpXM8GGs/OL4/6+k/E177wOTtOuxHnA5R9Rpp4EZN
yFe11Ak0im2duC8iDwOWef+hg9kk9kNIqphZh/swSnPhtCUd6ZLv+efLtf8Xlmuv5TfSXE0sjuPL
82T476dNxckZJK4OGTPnPzXwr4YalffDVbDL5WtFpUlgKH7RyEvaBnjriLbr9Jf2yUGwaeABYsjD
eeRuCJt3aW4HAdRF8y5PuyMa2NPRdKnhKngvJAYKTJS0UIx8K795Ua7iQlfeUch6vLnF3QkIfdPW
CmfEcLO/Oq+6eeDsoCFcjvVkIKmoWd3wFIBPvWU9gr2KuNLguqdM3wQUaCN79UKZL8A+a2H/vSAW
m+QTrvrmR4pkKNaT+tfyoHKxYGWVj6bdSBA+iMqAEFirgJwW0YmDAOsvCYFe54FmwsWbup7voedd
aVBjuI1y7Aa4pU14yPPNRQ44Mrggsg8g/US/XIoc8zv25l330ihJSbchNVqHxUxomVOocJ4B3CCS
/2Tmo9U1FdSBGeVpce8B/WMEv8cBEEsOXJIJ+5CXhM0B84M57VT9JO5ebnhGLcpEeBFOe4pESgYR
HXEVX7cXAur2cQ+wLxdrgUhpV+ILVi6dvJZ8U4+0hLX7Tn/wv2pv4lcebxYQJwpBJcuoCdpcYn//
8R/cNnMD7v8IcFI+CctXen1ni+jVSTylZXlac2RCv4BAr++0+GbDhGBtmDlOhTRt3SFaK5cnBcMb
LHL3HOZfJEpjBsm+PRXzEzx0niZ9WAFN5HpQMGaW3z0nBlr4LPvGXu0jI6XxoUaHGoeBF6dyjivD
66A7Ox3jQyhTLd/XiTDHePID3Jl3bUysSmy6FcSHGKs4QwvqbPtlIL+ZnGgmDLXO43tQ73/h4KmP
0XGiOqdWQ4c7onjIuxO2ncuArb17YYMbgAXxzVEj0DCGqYzdTKtnToHe89G6V20AJKTxaV7gKpM8
GmKFl9OSuJyZLyqo8SYlCEErQ+FvofpS3gaIAGg98Pr0AtQp2iSBFErR43S8S/9IpmI9QCzR20gn
pNnbQmG6T+aQIsJNIlhzWJxp2erKyIHUMjCTOGqaoyzWx3tXH3lAE592WjqwR3JO4krV1jxDyQfE
w4yvYHne8xzCdaTQ0KuovNL1DOBglqIkmfXfIZxt0V06wE5/R9vJguRtJBBTDKbK1cBCbnkmUsnE
iVS+OOhRMpvIT5X813sJXPaSUo6S8QaFF8qVpkdSn+JY9+j6zmwwgOtEHK0FJAS7pj1c0YKzY3A9
k2h5bR3K5Hk4Go/NJWJpwJDVVZ5VSmPeDlNXJDHGbT9SwCTQNOpJFssz4xANPosQ8vh18xY3pYeF
6II//M5+ZwPJBBMPadBqs26hm6Im15fpQ9BXEUooxcELP3506fc9rgs/sU/WFQ8yH0q+pAEk5r+C
Lev2aSuIgMJqSHpmSpKsMu31olLleHKCqYGnD+qO4XGBj4E6Nrfh0Tbw7XIeo8g8YNpoiFvHOvL7
LtDFxv5qg3D/EUR7drIDYjAcUJMDeMCXlfBmOfp3fnSBbGHtWuqhI3dpJwSOrCYx3ue7RKtkBgJc
oIPklj0zoO1pITdFXK+77lWlcgtY9lCD3aPMQ4GJu4xqUjGAnAWBif7fbN0ZHe8uCc9XwdBEdrBo
dwlICZSurADyX5gABnXYuEGYbM+Lyezq43LpxHbtuh7NEDDiT68bE/2pDCihyOuADuc0IlsM+w0M
WVa9fc/nehc/hgDm7dbx8JoKhrKpekWuSBEMAHqvt6gAoYFWTyeejmmDLWWrGEwOYWXQddTwbwXZ
fEdBdKKaOXwxnYVco7UAox7ooXgmCiAQfP6paJqNBlKv2qQ5BOMrbCLNfYO/bJBHXhBEfhllKfGi
NY3x0nOgi/fyq0m1D703hYazMoIWUM+/9uqdtHwOXMSK2xUZDkPcTrM90JzanAKt6naluxjrCW5j
fxCBlV651uREJoykFAfJ+LrDWMXH6hxan5lwmQIhhmihZVHzZwyivSbCNAVOD07Iyq9jPVGfgUn3
cwCGuCwiGVnbt4ciY1FBjWNw7IIxRAZKnadE4stFJ04Osh1utEXYGSXxheqEsj8/wulVML2TotGG
wMCWaNen05SQghjXHNkmU/Wa/7eQnQjEY27tmLUFB5w5scmXBYPRW/58qLjLzbXvxuWV+DsDVAiL
+nB2bXV0UdKg8AZjDMoqVmqXOBdp5ueQca/yqPXMdbsHwjmwW5vcNjfeI8JiNMnK45V4AqMv192B
ZQFRMktfOk1BuIfu0H+m3LJxlhg/HjvbJP1QRH2SszpYCSVNU1bCqwFTrH++Ly2j2n7vE7sAVQgx
ieAnYxPYJFoYfC4V70GGirqlDCdNB6N08XKqBBJ93yYIPL7dSiJ+1gQuH4wbzRReRWC0AecRy2ei
ruI7mWGUF5wx/CMjO+/zXvYoaeGgkQ+MAsBlyyqT1WDh68I7J7PWlK1wz6fjPslvGUEBK21biAZL
FCZGHC67nNd/upzFZwX/Fdroh/DM+PuROsvkvhc4cW7SiibH0H+AwyGqwK7DiWzb9aWYuilNh2gp
n0Ntg0wKpz5MK5byaIFLZWbhTE+aDxvV9ROwdBMhKgPD8jdqCGRSF24JLCH8nDUrEEBWDMpNIwx2
OLrlT24kXN9+gcc/PTT8sLjVRGJWmAyeZbP+iN0fK7V0SB44+Fs+yIKxDBh1OetMaUj3Ul7A7UnF
b/yJAzlyR6c4oEHN5B4j5E5uOGycC/x8uabiAJ7RMR52HnAm1Swbcjxx+Upp7d12qK18WYOEkMEN
ZKZO/SwZ6qTrqLs7h68326AEBiVuOoUIM9VyoLparDeuIJOy8HCS53dlRjYiFCnkBvSp/hFScLFH
1D5NA9vRjjYGUnyC0CEkVD4zKGT3W8kgRpu5zZW/QvwU5qjhFR/IIkRzBAKr9AmPgnd4gZrlhExL
AVujFk94lPgJAQEgmxNid2TpvHp2uF7y+ooLCnjphcKnanDPhPHrXsEhc7BTHxNU2qfbejj8Ae9V
N32X4H5LIVdFjIHtOb4tCQqYOZln4Xs3t70QSB+mE2oQoKMv3EG9fm7AaklBnVy9WNpSJ14FPr08
3koG9Syigkgp7/R5bGEa4Qxn12AehSjr+q6GxP1/X8RxsmZiM3hEnUwNfJCIuRafxp2OFY4EnAWE
VUap+8oSXPX+o9cPYQSKtHy8Sx1YS5PdmKb19gicepqymy1AvuTiWHY8YEqqwdpHwJllwV8xGKrF
NU2fpUDR6GPTUJ20KF8bid4mqmv1k1iJeiL4dPPyLt6U2DeBtjNlMH4qFQ487KutWtagpnQv9p/O
Pxcyffjbw/XNC99dvwXBduD0ug23SenSmpCSdCGEDosCW6MDHAQaC2NpWoWMlIHCoij+67IYTVot
LdyKyZlUYF6fZ9GFFnl0IHS1xMhoqvXp1mZiAWeM14VP18v+UZMU07Bj2cRVYdLfjAJujRvM3Prd
L4LKO08xeMYQDrJiID5oVBFZoR7gSAprs6bAWosb3C7bcNvfB6rg0eWHc5ib0aqeOMNQ1fNrMARs
DTQU9OiqqJ9+v07c9Pa7LjBfX7s5igKqTQVnU+OOb3V6ksdPnFzAqiaXZdwQ1z5liMzFGP6lSkv7
zDqf8+p+9ijO1YlZBSPN0zvQ381ITSOUclaeUy09Ly6iotvG5DaPVkZ4EuoOa7LYVa0VqkEEUwf1
22eXBhkZE11kVWVA5AdGPlJ0PooIHazDfjoCuft1hxSptP1Y9GsLIQdJrL7097koww20f3FgT2vR
ToSwEOOROxSRPPfLVxIEJEI9kgAvai6LEQv6YLNowy+q9ie2dnCORmavq7EZehL606JQizF+j8PK
K4xQz6Bqas+gfrTPugHzadaH2bmQCEKNPgUO/VqFRv63EZd5Tlggwetz2bkic+VxkbJCbd452evy
4rSdSLbPlxoUjIDBYadT1TWpN94p5jP3u5wT7nDc96UssG2NMqAKVzG3ISEDBIRX3IHFW5Cgx2Cv
6BG1I2vl+Z8LrCu7RKdXj68yvpgROHAPm4tu3EU4zAGLBkSJsF5TxktwBg7bjtyh65hZTsAxWvAW
FcRdhZs8xj8BdnyZ9G9a+k8E8UVH57DBP6szvYGaYlrTYP2TfHjAcgHfEifPaNUuZq2HhPTgrtZG
x3vqkMy2QjhDY8EqBoOB/M5AjWAHC5gQU1pBOLdJzm9GLICxHBVivdd9VYRr1W6p6hQXpsdc7ZwL
f2oTvlW8hyh0bLuwsw50DlyHLWayzgJubJ4y8Bf88vae8jLc1wAkE3NMjkTw1BtlkCenThyYQVKm
eCUJb8M0azxqeqJgm1vdM9kWM7FHv3hMHIde8GGgyJjixxjewX6+T3lzOiUt3EHHJqg94mN2cVVL
atsxFJ2a+gOiMtQuDiAGonzXb/Jg6TERRRatmEp8JYD2cA9ohC9LxCld4t/zbh+Pj5aPy0uvG9TK
U1Rm08LD4ElSOt18ehbo/mPk4x0o7dtYtZKs4cwKRUN/dL5Fcrb34bzMio7vg5BJ7Q4cOAxcIStQ
m1MnqK/3v32Iv4uyUuKDSqshg/sVUcZ85VfUslpwRGxaSb9jyL9KoZw5AgyVbcD9LYOyvnnY0oz0
WyY+BypAsrZPP0WQydAQ8opVjU0m4yRL8LP/wHzU18ljkErngkfUsXot712ia7mi7NoZtzUPBFT+
ltqQfa9+bWo/dh++hnt/rOW/Ox3ee7kSi1LPuoOF7SryBXOfEAqCXXm4zSnKfefQ36tYZThYQXA/
ySeYngwkZzFgVC/gf6mJKF/7LDz4faR6Bnqfyqx7pDi4Y9OZI51gR9hwIy8Y+bJOkS/eDg/sHc1D
UQwfrdPP3rCepbtFyQiK7NY8LtZEWlZn+UfbU3Vt+iiuyKPt9SNWiyEcis1Z5pKEk1eUE/Y//Tdf
N2ECeRM1Cs/Uw5z8hgfiAzcZYccTxq4pXTHyVi0xHuE8jR6tB/0jQ5T6eSva91NzhR8kM5WmyOp6
ww5MBOjd5euzmHbBoJvKNfYWx9HCwudfkZkQYNnUk3J9PGSgTRCbwr4BjdN9sm5UptQUyI50jwMf
biM8d/dnBoJeV+PqX5znucBe991om3k+/paKOh9PYe3g3SzEvgCMSmltwvd6DXLSKKKXVszh4sUg
H25V18t8oNQQFiAHBcVkH0aB3dfK69vIdrG8zEzZlJbuDjEu6ZuiAmm/6fgyhb8NqOlRs9H0tsL6
80ZGgnsjVBPODOTUZAGU7CGXoTD6Xx/zodCHLHZUhjLn/x3dt1TM/Y0yb9UxnUEtz+FdhKzMhMD4
oWVFWzI7zdxnjCiyLFPGERSnsYW9PRhDbRlyCMH7LbHkbiD+SGsz+KCFLJHq7w3ujVg9Wpz32jvT
wvJEkkRySvDKPfpaAvncsRVo9KBYtTxz9IHsPA==
`protect end_protected
