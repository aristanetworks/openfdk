--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
hLLe2byvq8CfN17iKVdvuLdd4K1pdlUj122OQZ9K5uRHDHxtNVLTdLOozNgNKwIl2iF7UfiF6FT/
CxznRr2U7pEO5aMIOnFzkTekNWHZSBK8Bf4aNoeNxAhPHdIA4Dg7Cv7OcVPellwIcBJMYXhY/LmK
qTtZrG8YrSeAcTQjRRWZOZfMrwhkOXF2DhTNbTB+uKR7OInBNvqEDEUXJ9aZYNubRGRaoFB8woTR
GZuI7mejjhMsk0+LaRqcoOMWog/keeUrwaFUBqB/Xb/ww2VDlPwX9jtl51f/o/AlgyqXaj0Q/liu
uH3GUvk0vPzUDI0UbTJ/g0kNeZ9hXa/2qnJQCw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="JjRcEllJVOjmk67RXL5Z1/C0RyUmIXGZ1d07yWD+Ygs="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
VyshzAl51fMzJb4FbCv9TyfTqzuHXaJIva73JYvimHp9vsHkFO/Ovk0O87s6XnpAcjRidxXfQgUI
N1LOBFSHZckkKzrCM9WW5gZFr0YUN3+s4yaAmebA3OwKtZ/35RQ/7Y8m5BpzG3FtlVh9/LteOwc0
7UupwyLxXQClruf3i/tQCe7KYe0DjYRTtiMoZoUCgGrwfNGVDHVR4wLrLyJrAaadKjJagXbxt/fh
o2C4qpKgWLYbqL+aV/ir3l0lZb97aUgxFwzeZcY+HshF/3xD0DYosz4FE4x55HDe6sCKbhnka50s
AoX0c0Zh1BcUH4s/veyunQKc5knopM8od9HEIQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="3aAfy9YUJUbtLZpJD/LPkRVZAIU2Qi778zw+PM8/MfU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 38816)
`protect data_block
lbj7f8rwVbd4CHyXApxetA54DR6eKGgRWKM1O+ZtFrLGIDrfO46OkZ2LbMBXCx47s+0tL9Ka4loj
avAbJzMUZTwZr/LklkO9Ylg4b/y2m6tsLGKmdrpx3Sy/ntKmrl/SLm72idtIr/A7wmPSoaQxD4N+
Z+CYO4EcdzmXYeqig1oJNBOyqF7lguyPNDsQssplOThR/0w8Pdds+7XbMlpTWSZx+bqqGGvQ2PEe
VgBdR4H+0l6MNTeFRNd65lX/ekxbHElbBhbmrtA9aHsbkdpLJhmBbKp43rCHvVibZea+NxNLbuoJ
QjtzhJSXMwjMEbZwID7P+gYbIwvCRwt/C8eMAFBe6iU2ZXhu5vl9qucZMY9N6r/RQ0Hza0qhFQS6
zNJJJxnbjAn0yOyfE94kCMNY4U+nLH+32EYfWkEyerFtE9E6xGLMrw6HKQJ6QmcjojqLUwoxJTdd
IuMgG9ntyhVNkQH+oA5JeHjQ4u0GgU/maRUl/zRds1I7PeuDptaDdzejQ7MK7ajGg/DIiwx59vLY
Hgrke4OcNZUIqYBrftTljLCDwTAGdYFVoi1zvrUHAQTyaI7oGJhClRVQFEnRcFDnh5h9Lx1d1nl7
wAytuVdKtxDKvquNF18gBpxI52OdiLE2xkMaJgAP9M+tmPBVP+lYa8aYWZDi9sQQPkQCYvbbqH/g
EKJjk1nBhWULEEEUf7RqB9Z9ZTRCD4n8wRXOV+JoZ04k4wvtLVBtGNUBkNDzWdZCJxcdrHrAeikq
pG8O9zKI6W9X7un92WsRkGI1uKYolQ25UCTLk8slu+mdhOCr8ffHpJbxhdGI4nxtWOWkWr3bFxby
DgUNMJ1o8wTj6BPScyvjZOAuXp+wlEwy1k3rL7q0zyLJuPe1MGdghtnxFNtNG9IMrXIqgMF3Qvb/
73htch8ox84KD36mJsnzWJzPIfm3X+eC80puEvRu4M8cTm6czfDrjKZmX5YeD+WaFFgqwdm6kHmH
EUkGQATkI67xVggxpnlmU2qBRTNyIv0L54SHjhMdUw662SnbgD2rMnh2bQ3/vM8JTyHqdJlH8mVK
pNnZmkIY/vc4R4QbmMfQMaZnRsZp9iwCbj2SYxc8A0QoZsfioL8WbcAP6QBnIPW3RsuAdhDVUQup
UVLX97G14a0FAlS6eqZF6IwOsR3Ta8AD5kXVU+SJlGEjBzu2B08hoaUPRI40MOrEhT9J9ccPUOu/
s41qL3j93jKu83RO1fxNpIOzbE2YugOFMU+Hi3ofgj+z8NjsuM45am+E5b8LXWSvR0CAC2AtOtdK
QR8bB+4CBEP9s4bdSxutaXGd5LjQosfMN4mV9I1iAJCSrjZQ1AR+ekyXiCOY6bL44kOefwl/TG+m
hCBSB3q6++AJV2//vY8H2jxnsjZ0+z170pixL9kSzGnnt6kYaGC6jMRJyBPqzN1mG6lIiskn4608
E5wZ7Q2n9TEqTHvjoYRc/3IZvwUci208gjRRhplf2iHJSyAyUJVsF90+3huYAbPKKsBTgeTrsjRo
rmXnxOHob9QihMnqDzQGtjAcknomcvEQ9pD+9/pc93J/e9DHYJdDQJOQsiWS+YRZV3V5nNi+4SDM
mbkRRuu3G6hvVTarvPZ84tK9b9szy56AK6r14JTFjYSA3ezBUTIdzwpKzRx9p4w2iqpKT68wLmHk
QDij6mrmnUVHUvgTdfcOFfVV4nx9Ch6kAsRC1W+aGWoNBsc5r2zC12s19nWGn/Eyf2GAsCdbEcAr
OlnkcMj035vzr68+Lk0gy3BpE7pYGTwNsBl0F9I6bY2ZRfGU4j6XpgTEeT28Tx1s05pELRZN+KnF
osSx4yEy3sJ9SMItITqvDFS+hMErjOyk0tbgjwvKkNuN/7YC+rj4EdNIMBSbBFnlWr0kaNaT6Db8
cmJ9WPiG/2GMkrHsEcCwvz7ogspZOnIPyDOawTnuHfYc6T4psLWff/9/9XDnX7ZIQ+sF4iSZH2bu
MwQq2iM1WbKo60U1IfwG87lZCoRCOHY9P4sZa97GRKw+vSFSX6GUk8BFnofHHzrVa7y8Iy/I0W87
bLMo9zd20hlet1ISh+022Gk3Cn/7YXI5sWvj7LxA/PNuWdqaeBoEg3hrdeGRLReyekX0k3dNchDK
Ts6/BAXYM8xXg4oDckYUHOGx+APuthgwEJQZUb/4nn3uW9hrIaRBLvUkQvBLCfG984kQ0jaCjH/V
FqawIsyFZq7Dzm4hpXM2kKTLZpNluanGSQJXdJU8PqrPIlG0xj7lReVYUVRKmjh+YIFJ8I4jGMLe
6PNwkTQv1XZn9jr/N758tgl/lmg367xPjMZ5kCTgaeLgk/iTHWy5UXoAOMGdYJpFvgbbS7+Arg6J
HhfmBeTtJIQ8hYXcZi8AGXqP0etOIO+svQiqmDaRUb9WGDQpMr4tG01z3iVN8//j7uF+EiSTOoTG
HZ6YVe9i5KAoQgFNzmLzPw5swBsZ1cbDO000VwhS3YeRflOdlMmXO4IC/cXn/j0LAQsiFIifHEsE
md8fDKWh7iqLeU2LOMaA63XUmNfLni7UvyIJTAQlMwe5UfYOQ1pd2UoK0SWmTz8VF3RjEt7hhqX/
oXjJAc7Sq75V92gLvoWuYkDXOt9LTvNZUgqCE8CyFVGIDwogH9avW2nUmR5xsOhvW2MIBjb79bQS
hr37UO/UzmxS5XIDxPvivfsPGHkqbAOJCN/g+4CZM9c9iYM/PX8eFaI8a5f0GWJ9cScjj/iKRwZI
FwUutnA9k5g1rzFGvQuJ1XhOh+rRWy5FvFodx6WxBevK57a4gQrYFWRu+Cg0fI2EhD0gQtWKLTBP
wf9WRnEI7LBdg6asDewm3BsZwJ8F92E1+uCUqDtDQuM1G3M3kbcdUfk4DM5qH4OwS1FcZwQ4vfIm
lch/sfmGRMOXn9gG77U5J7lt/uFyfEh7kX5M0c5jiM5cwxiqu21hf82cL/UNIp53Qta40i9HQIBl
J5Wq/vtAamM7nsWfFBRlbK4gP87jHkzNCFiCyD3gZR0x96GxhCNU7PQ9UVJCNtgsO2peVJ1rvRMG
K22erSZAoKkFYZ0/UAY3vWiusuyp0n+YnTApcQyr2kPMTOMVcZWcELF3gUrpTGEU0QWgVcuMZuTI
m3LU2JdRU+/6TX4iehMqxWX431XcPMB9ll5c4PdxlPQRBsWmDNYPr7iuquE7kOG4xPayYbTwd/QU
tJQ1FDrlWbgHF74fX2cIjnp9n+zBXx1PyOUOU/D8V9nKsLGD3BYhnD4pH+lbZhtcipNt8qGWM+V4
juSM1OUhToIo+2JG0qllAPkV3lSseYP29BvuE/iv//RlUBAc9rY8V8Il9BntEvyHIY0fvXXVPqGf
Lc20yjCxQJ6mUKaoXUaclWdE7VqhdZF27RSibLx+7c1dZwsX7hdrRYKRe7qJHRyeoeO00bJkQeoP
WFe7Lrnj/Dukw8PZwzaRywnT1Bf3bDPLSXEkQCaYBmT5rakueeQJBGNeAuinvbE+I1kBE5XxSGyk
6zt8JIb5xTnvuhSZp3yfalllvPOhrYVSwk2n58hpsmuQtZ6DOtF6uYOuqANmV3H1cIFFVuUfAeuz
UNfpE43HS/K4RadfrysYktNgklaB2d6kTqOxj2JQ4ZlTh35tiPLt+NUzf8PeyNWBXsaqYOUW/33+
y7iNLvOLdKTxSWYUKtxmaswEr1FcNUQvoI2tq6N1KMCkH3ApQw0GGnxX6ygP5igwSiQ2WtBp4+If
4eFhCBL/+R2gOwosrct2US9/Lpmr9bgelaF5QbnzsG0utVKu9Drh8tfUkawvvd/DfURH0JettB+s
iJYOuXzmhbAPOhfoCaOOPA7OUIQ4Igne4ZoF0qW09n3wk1B38wSztIU7TwuXkXsab7+EjMGVAkgI
runw6V2Dst9B/ckggzKDkLO2lxKO2VERWjAZ68fjAk2IQsyxT5FyQyQyXIikBB4S8nX/lTaTQHBI
qfk9FfvvNPc1uetjNoA7gUi5z/j0jifFvfZhJ6yc0/S2HGn14eXjAsCeuq/N0em39Rq7FVDUICod
7yiWLMIjBuEUu1mRh9+dyrVo1akNKSWwSoTxVvUu9VnqZsqgUgXniajtrGiD5KcgBemUBBc6wkY+
y1PnyU+bOGGUJTc40EfyG4ZmDHmIRRBX97rBJUJAiZm7KikcIwJN4nxAECFlRO3J7KjzOxI4DZiz
OFtAIqUsoSYVB5/ikGRlA7z5TMnRghWTI8HG4aQoYUx4h40T+Y1e+XdLc4LF9nuSb21nT2ghVNgf
sNiI9wt5BJ3xp3KAhHaiM/I4xF4iGVhsGDwFn3+wqYRaZKMWD+Mn3NV2t9Lfhy35xD6XMfbDXzT6
OWCDMZsH8C1p5AIGe1m4I2GJcOeJIZxeErpi/9TOP9fClWW9M37SUVIHx9z4PAPryUX1JFfFsEpv
wXpnfpoV9TB33bT+ZczY+0aPnluV4S7H1uhmrIUscMmBJVfezRlN4MiITMHnhkkzP3zx1fOs5G1g
dK44CWIJcU3780ETK4uGJ6/1I28tE/52g4wYgyOp47O2r0X3zdu+XnFII8jY/7ID5+PG3/SmfwD9
DtM119BLesP0L0zXmAbfA0rYuDuH5IrMin4PL1VTDIpmtma/xt+MyPxLht+7xwn6oeLatTU1UioJ
1HxxzAaC7p0yAHPaM0Tt2EusgoXvs568O+xGXPBcCisIgTTJLHAtbxHiKJ3tKm7NctB9ijot2Gpg
c14+BtBqnqNlwVGPzwOt1bFzPycSIVRQyiFqMOBwI6UC+hzMWpEMrC3i+i9MxgCEmH4P5Ol9NEoj
vm+dwX5UO29kxR6Ssbvcz5TNToSSoTPJ0lA9KvmxH5vOmUFNbkNqRbyVtx1XyOvlU3Hgxd/TBSwk
DqQo2r9p+nxFTVsM4yodccCbFDHQ5nPAnVA5Y1iHBBCcueQj2zLmFnH+P3H714wLfsWY0Yo2SjKW
bGvko0yAN1lYoYfsYR/vZG54O8lp9ZTL5/9En5qNXlyzpR/a7DzXwUpkeqvNVhrxXyvodNyIs9jg
1bGJSUiGsOqXC7drX+cx/ZoAxh2+5I0A+GfH/ZRF3ZjGcG9lXKvG2un8PRuGBgMXyHVqYckz+64Z
sALqokRBrj84NE6Mhb4E/fVAB+Oy+J2fCFfW+WrF7EW2aFaP+Afg0ByV+BALwP2RKbtqJuvEN29+
boTrduEHwBAWLepZaYsQ+0cmeLTeQTIWK8e2iJH3DJwiqEyir4JGTuWMUynDGlHQlKbfQjuymJph
PTU6N04YVm6ZFCKPGD4vmtSo0jElJVuZc1alSjPu96cSMBlv3TWEYAVwJ7hrO2AZo+2Mhc+Y3Hj1
I/QUMS9vBTKdZ2pl7wafNdP0RR/PQvlS8cGYEXN3DL5PZk041BWqjJ8REtmIKDNw/FIuXdTqqAR1
YNaqscLLqNpHJNeNUy9fAAmrIpTMGglvLn9vXW2UkrsCiltX/gv5C04B1crM1cIuAFpc/RJfBLhY
ZM3pNe2G+H13uFBpv2thKKLLLtRgyLIH8T/sE7z89ZAx+1ey2UtPEDngsWPWlmLi4gIe1sKMjhDG
pnV0n7nLQMstFcf0fx028VlbQdidOVMI6mFnyW11MNlNZsx1qq/9/Y951CSryXOhgL7oPzI06lLi
1XEvRrlXCZr5TrRaai3VzBl5DM9m98DNpEhGYioOy8zwqdoOM7JbbL5UEsSIGM3fBnZ/40Jh6ny4
QHcjaZR35B6dKFiAEStUBzzY0yg2C5zlASHs5jtGQ2YLs4HRNURypO4oCpc1riJM28oq3Kh4iMXG
7F7nLAd1dggsjK1EVEieeRyoMPW8RYXa+knwbwJcaHR7b60eUT3bJB/LoTH0EV1n0kGMojtNmKfJ
KSGApzVW1mh4vupcQ99O4avmOyEnjygl+5fN099s6wdiYw8iPRWAZKxedHJH1wCVOfe8D0rsGQ9W
FEoUCuRWnDG7QDf4pYJKRZW0ggBnkh4v+5FAWQ8sIUY7wC3LJV78LTV7YUQn2VJ5gnjVBvIRP9W3
19LnNdskXdZyP1Ohcc75wmCY9wEBv3qDA8uuSf6DsZ0bWbf1LAaNWu4e0Pcx1qOCjwWI+gUTUQft
f3/iiUXg/pu6JBrRPZ19oyUPw+JPA6pJ+fyi0d/QunUJ+rBDF4UnZmxtZZzui+ll0uoHfL3EHHKn
jX6ShiBAK1U9B8x4IF7JbYUWBywr/YgByDX8GQbNZfk6MP6USBo67nYebtjB5zQPHSAVm0iVvEzF
M/YZx7fG2xFUIwU3PWUE74plsjR3tzlMDL1CG9PJxjckRLpl73tOMR+hyoCCfpDKdIzBDjgTvns3
s0oqfzN8ur27SnL6IRpiFdEvo2cjbDdjtqPOhopuagkZd/ZnFti13Zx/zfGnaNp3TYiCvWcOMmil
A2e0uOJvy9EVTZ6JTOmk5ychbl5x6TmauoZN/k1cOzvIzBQTKVdVnJwJkPbT9GK30RO0RpqKUDEY
WNlgzFJ4qIkZH33M8OGf77HFzwa7O+qqlUldD7pz9FA8fhUOn3rcy5cIrA3oxh34XS1+oqZE3oq6
8WQNSf8NrZ9msI0CvUTrUhcu4x716X+r1qToa3uxxaI6hbUExAqE5p49nomYwYKXIf06SSXXmzo2
EX9dDnmwHz9+yn08mMco3iaPeTqlbVOM5P3BXyuVCKhM2MHI+Z0InQ3Za9s97/yVD7bxJOMbhAzA
cbdudd/07fU21o27yflaP/0+ttxJNEm9RzPsac/3U3xqdcWN0t7Y2cZ1wK6OkuXIldSQYyzcanAD
tMZrbUBcqJKBGJqzs3FA7bYPVQcW9QlY5xDPKtOCweSsc1d6YBsLPIh4glP+yMjRCk87uoWTSS9U
vWud+x4XVBBQKZFrB66qgaCnNYi4/nwRisWND4cGijVu8QxugZEagfYakY2rhsZ1yWhTjU8hIXZh
XRKV/orcgtipVskKK9W9o6TafMEYV3PaBnbtxyfYcf/kmVWDiO33LQ+lYRzGIuG28vtGx8s2XBUl
N4Ek7SRA/8aZScTyG5Dg/2XU0JNPFw0yhtFhD69WsvnO/kHw9GypiOZ+dhNZRNmpVoRGSS4z+/xR
bkUMzyCa1LT7IQMSdK6BTqgC9NaGZnn69nvyQ2gMl2yN6ZvXxRX6iQSGT5UrQ4v4rD1517bbFG2f
JAtcLamiBKDWktahNEugs0t79M1JmcLc2ua1VNn0QXPTb30WMDqapCDWrBJCJTH5w5gNGMpHqCTj
3hI2PkyK1ejQdI1fPYDbxYJlCN9JYSJgvpUxPgKVg89eglZUGMTX9MyLDbtmjuO/DqUtWRTUxurY
TCa8i+akKUZPztKPgce3OxR/moIZWJW2ZleSwqldR3biy1kojwf3pfpwACcSwC+tl8K+uHCSrOMj
LvTkDRBWofswFuvIRqxy4iw14XWKh9VT863Ol5iRQtIK0DxaaU0vAof+HfIbpl+banw+NIj56U+u
vEqd6tweKT1PcV7J7RIXv0bgxXzukHRt7rYmo5pvHWjBHsbdXrViTAhsUs+1SBwOOfGjI7jCNRqK
H80jMWt6NBl3xGZh3rs3S7yVBTNW8XjIS48O0w7ELKmLrutXR5CVmoCDrQkMzXFfDC3U+JEpC8LP
SM2+b3E2JEfFeQs4WKx2ktJTvjf2YaEEwt9b/FEa5BIdV4OWkZV5bRjyVkaM9IbVqIUokjD7kHN1
uIKhkeUcVejhCGw+5tr1EcpuXQ/i8fTWxxA2nZSmPjLhu2y6OUR6A+qx1MoRwWK8xrknbxWpi/8M
WD/F8UfTYgHz3aJSwCHQz68jHuWJUbTZozFFZ5gRGm6tZmLMhbVYziakEj1ztTht318o0BaZrmeO
w0gGE/t9fLfIxAotT15bxra+4U/0ince7qRWFJGuypupGKZ2Rf0JuqQnz+Roy5ggCRFe07m/lxU+
ZQpBONONViAi24P5iRnpT90CX0d0duMk0qDSum7KHWJOzHoG6LcPetv0VfBjPF/6ty7xhPRViTM3
H7JBy3Nrcw7r1gud0MOtSsRTh8xflbLItpgNOuVKJaLRC9gOg0/ZyULIlL2AVw+BfhqficYnsM8u
1F4fFbS5v+bnOgRDctguVEiBY0zrp5rVtt/xNQ4Rcq7iuQBdzg4HDnzq5Tm60MoQnLBlsTHJFOup
GB3knvBJLFLtI/D58xoL6yfN8299i8PcT0Ra7QVwEuTAYFTrk7e5nCHjjTfoOLsBWjHOpmJ6CHES
WH/5gYlAB8Qb51z6sSh+WJPfHEBhUpVgdW1wUehYy9hsljqJKojPDKmyXGnTGut24WXnb76mcRJj
4ZalP9WA5sT10bZcfsHO5cOx88zzX6iP+dP/c90IzTMQ2un/fdt57SBApG47ztN+CLHf65Tz1TD6
WEiBDLZEPwB8iMe/lYPqcyOgeGFHpjKZiudeD5JQ5/SaF5J04WBavrGt5XI4OpZMK7DriejCUjoq
hLdlfnMNJrhiFanIrjpuOn8D2Y4eQykCx8HQiuBwWMV1iQCvODz4MOpFtlLC192R7R/NFApsqKdM
bkinKjB6Kg4yAtQcIVOVo1QHl+eeEwd5Hal/SU5FzOaU/hoiZtYawqrEH/m3XCJP5nUlubmgp+nv
WPYwUNvvE2pqdXYdW4aeEhFK7rAs59VuwE5fuToimLpCe1D9nUcjSpptyYAg+NQWLai5WSqQigKq
4fSmvneIsA9JZ/SsS7Tb3RO4Si8zOAqPDaHIIOVID3F6f+6nLFBTc0WjLhrOWoroBm4nSXV43exF
DKJIlc2IRhh4lCUpfzL6nQlDS538bSnuFhi1pm5hLSM5q6h0gWe9/RW6ANYdbNMQmS3px0p6quGn
cDqs7lVNNgUdcHP70u3g+Rsaq6dAo5XPQlklqpqH0bK0UoKWi0JGeKMTB65e6OOn0gVUAQ4tjL1t
D3HncPmGOVDbqn0sYdVzGZj5RQ4CZyMdjYcjYeySC9so0EGzSTXt3wdOOSvcS0tKYjrutzdOZ48k
YGuF/vL7zmWlT5OAEDuhw9amerOQ1Yjdu7NQcHFAA4duOD9MZ3yrX+JWGsjvzrB+rgaPCsk/nC2C
9GvCDfjeCGy/gZm92/KTe4Q9+hAQKumU8L1n3fcasSQytJT4oKSVzv4VmXrVqLqeR1bA9USpHz/F
/XbvbO9OAw0UGc/1ONLviLpGbIJhIGCq10paAFVL1qq1uymLw1Zp7XG1T9lPsMn1E1LWR4oBXcHV
uwcOBQcwR8kHuK7T1lfW/D85aIlWZX4pcGZHJOKQEscL8Tlb6lm/ormcf8VDJHTcIdPrqZrLK5W5
cv55WWKY518kRuAXedjSPntCB24NkKqkyalhMY2mL32nhrSBfdRGkZyBYKsrHfOHLjPMbhnLOQts
tEnJgZv9iH0MR4OfHckeVdbk8g962WdCCfl+/xiI97/LRj+dKYKFQVt8Gorm6qznbMavOIulaYCn
iz9X2DZcd05eEMryZnvdJ/8UTnJ1KCo/lYtIrL8YeSl+elwv/gVYDnSjX5ycNuBLEeqwYlJTV809
a57p4eLvQVPFGe6wIeHYACRefVMtf2q133VmQLS9l4fLfD9NGmp0nnDAI2lZCavA683rrWf4emLr
kpmd0THzbsDTKi0ty3zURi9Rw2XhYRZJJWfDtAYiE0/ptYt1pN7L4JJqwdG7Y/f7Qsr0suFaxIFt
IplEgZoyzBwOfBd6Bfvo+oB84rxmrzOAO8fBkELWenghHsVj5Q1GMTI0HlN0ZlM0/pcbWjfwq512
QVD6cVOzrtPPmBDYOH7NLpFXn0aE3MCM/3h6ao5koOyXyIqFD9ATOkOwQ7NB4NTdo6+2xa/uMZfY
+WG6RxBa8yvsy6c1+9Cs6lELlvQJfFz62x5RYX4f75Ljiu+7nzVIpXOXb6iZbAIvqIeNaaYogPjI
9HkcTKSewtvIubNpS9sSjJ28zTBtpX7Yjm9U3pX7KGTFmxAVi/MpNN7MHbpQOes/uZqqRsLRb8dH
QYajmSjWIVULfEcah9ySQuKM8/cg/Q8bLQ7tfnvxMi/Cly7qf+g7uD9nKcET0Rqy0XkedcHCG4Oo
ym3+qEgSaJbrYI6iz6w1XMkCiVhYuuBuvefcqjmTgH8r2Nkyr0bFnp6f5M0fEY+uPNKSexM99wdf
nmrufOzxCidsxViKTHy1IAS+SpvIv/7CTdelXs+3Z1O3JevEKWooJRcnFiPsYL0Jnx7r+L4XXUhw
xVAWDwb+Hpob7+gtx/680peCBSQDr7by/3bBEcT02iXInwaS5K+rlCgCQyvW9lrQ4GNVO2DW9oi7
H4QxsOBtz4AZr0N27f+UrsOtOWR/rhekYWCu1+DM/fs+RkVZWRAvisMohxRUAyk95sM0lDctP7rq
Ti7YsLk8M9+e63th7EqgGs4S+tTh8VA2H2Asi0Rdy9KxPQDxe/9tYGL/MJc4T9P/MHcZa7fBdK8X
R9+m4J18ce9F5q5YfH9e4F0DwM2F9fxY3uBABSpHG9nu7BNqGw+ep/LwrqhZC9jH7t3hf+iEltJN
Ra5gZ9zcU4/QyCbacoat8nw6hRbkmxXk7qMK4iJ3Yxt5oOsncjg28PLu1ODzHF/irmyhsteRXthr
pkC9U7vS7F8JSIa39+OdaHDlme/X+kewhxyqb7lhOa6b3pavy2z2eAMw59ai9gdaNZIk3fzbTuUX
DL1rWnavZCux1cvrzb+fh1n+/2ExGdEuC9gssaZNdW0PqWTDUMiOQxndjaFXTxaySrQcuzyJMo7P
NJj1YfJmhXb6R7SkXRvx7P2upsgWrTN+WB8/HY06djqAFiv/WiQai4MeURQ5cL/UL11piEtaS1d/
Yc+HM+YXoZBYDl4JEtfRuemXQ8WeQ+G0WMGRFjVcg2t4+azlNx7UPzc2U+oqhE7Z3BiJCedHx3lC
GYe/Hdd8M48qFM4GYTu2n5hCTzUpDzPu7x74axH5+Qo9zpf4orCgvsYu3STqecDbUNe1ZDrZZDm3
Q3fu76Ww/75aHpWqlkB6uMCPYF5AuQ+ruzpWAJ0kUQMnMx7BD03N1RJt1HZamUnViEgldgg3ejyT
sWyZDCEUx9HjQdHU/wWydi6nGrwtNATwytmw6SRf17W9pMx8AHqDxXujNfdpWnbnL8iPxPiqIf51
rb/piGlpkN7maCN5hi0Nrn8Njl/v4qZlR2g0VAXNhCvPVLr9Iz0iKvnrjsCSsmekax0bLtrNs3l3
EEVRkdj1sJw0cEER8KMoubduJAmZJy+3jdYb97spPAa4080Mft2gmCxxv4ZimHphXQFuyZvizLIj
En08jf0tqkL+twf4iKwF48G8ZjYs1m+KLTVXUoUckGVmr7BKzwmEcrPEPU0ygJYYAqOl86jm16eU
YZhjm8DJncgPisIvh5AShFFpossREqA1wv8ccBs4EmbUYYYHFhF3qTdtxdUkA7RrDDH9cl7FGCF1
ZV2g42l9QnCH3YMwhBHZI0Kxc3aBlDGzYhG4S+M7CzdMlVW4Z7GZPWBj44QUuJFc6V1Aj2h8s5ZW
Z0a4UEiUvGRx2/MVNvC11lbbxaUfAiFI8X3ZmGMbRsYqL2kCJKr76oh13LQnPyI/2BVTEcDFysXv
KEpz5UUstijstz+q4WwzD7ksqb1G3vk6PBnN/TxnX11Y3x/oL4dydAgS3JNzW0F5WvhhcI9cjmmf
QbrfoyuWtqXWqGn7M+4Oz3vMeYeg7TxkAPHs+8W1YzJCcqfg083kKbAQYaG9Ob17POJH1D4pwglh
EiVPzRJB/U1kd727QMFoNDdWtMlHKt/ZLOgbj5/So0fWiua/1rAVCr3eYlqnYU9PzUyaNUbIETqh
H3KKGiYjj8kpZUjD9b2jR/IdZ6Rzj9b0+TOwDETk7IP1S+k/+0lOVQ5VIodOYxrEcRTblvRdPT5X
3nVlR6q21mNdPxcZ8/48HzrUIBkzLSuP6BoimZCEW1W29V4iPVv5J6Mc6sP6AtpVBr6lDOQlZHKE
n2RdvAbqzkzmdLlQ10lyT1OVJ/fmyrgJGL8HrgbF6v9wtqn/S0v+n1YYrVRBhXZ3LCPraCraRxgM
vOkX2XTDbB0XOBJ2Vden16/5GnW6gvUtmsLg/MaXUeN7fV0hdamnDnnNUY91ZUREsuhlLIWiZOsn
qmtDWFpW5RY2QjhK+3E1S5fG50m1tGfzQtZsjGkMOkIkiORthTYp9SGa9Rm+u01kjPtl5FOOcOaO
ggHRgVFJVplRIyJGbIYtHHqrqiWDF5k1lI39qqU/65TXTrNXqfGPaCzd9Sh+F8qb6Bq6hoZvQCCy
U69cb1z7O1vOH5xnzyRJgtLzDPtz8nZaXn/oEnYE9bC85qtpfF1tTGPoEm8J8tjzGKDKIJc8u30U
CE2RlUk4LUZNuj6vQTq6gTBeo+QvT31IOJ4IDNcSFmmokJPASphFuyhkdkYFpXRD2d5T8VJySl0c
i4ldRPjhWL8r1wZijC26wTKmx/HziH5aST39QFAPIxGSirDox3eRfalpWuWlgSLXwS4AAe00lFRT
b0NB9xrJu450W1T0SRNtXfHIXgmnhgAEjAXzBjjzGW1LRPwY5gkAzeeoDDY9jv8wZ28/RxV1FwQf
c2m0tOnhZ05taM/xUcc7thmmgsUlhhSd2WGocwtIUEZUJvMHZgYtd2Pc2kjzEBTzi5zY/fFe8GdB
vVFb1f964Q0A4SS3+h3xFyl+DBu/MsOAldDsCKxQFUhvbomCAhkNZxPhPdqBhOoL/44oBYEN53Hb
LZKnAAvjJFVkCfui6ksG/nnNSH7m4CzEd43XXoESI4m/uj1cm6DETVMvjeBTjiGJFREQ/KK7/k19
XJLbGZfa1BDKMCBtJyrunVwsrbGUUmFqJg6nmS5blqPuWNiUVk/rLrsvMD55yuHYN8+yTas60K9F
7HIGEfzXy4W0T3swK5etbb4NOolfLP0kWNMiahLHufkW6RnNWhVb99UztK/E0zSA/3r0THPl6Tom
fr87NQfRc1ZlZoPbMWVeTPjh+vJlDVCw/mc6uBfo0SY0zs4yhpUJ4xNR8fOlGQy2goLPTS5N7RXD
o5MmDSRtMI5P1L6kLJZoSNBMz89O+68acgb5SLcqXpaBcBSdIxLJ4g8p2eXRuFRvQfiLpvw02GrE
K/b9NTAHSZHjk2MLWeGD1Gn/dtiP/KcOTvbSBAquBI8lWOoIvH564aMb/XzNq+kbJ4Lc1gu7nxsI
Gd54vLumw/C8e2MISk46jhEzhbpHSX01pvGlqmk+fIY9R1x5pjI4XqYbd1dvX72qXfppDPdA2vZ7
2X4K1mOWRIGhDZ6V4xbwSPDJorP4Md8HIULu+qhb8a4cvRR9S+KlbhN5cfoFtmjxI+b8ehOypS9k
MYTnAVRiK/WcoLF0UrbSIAhRJriroaTcridYnv5MevFg5CtdY7ACvjuT9WhS1g1lUmBqDwL6Hjlz
FwE5z1giC0OdqstkqeuFgXkTyHB5i6dnOafeeDEb+zYomA6P6kPZHmPyE/D/V6jdut/cXbUGnfwb
Z/ThS1uqw+i6rMXogbr7IJBr2E8w4swx2Wj43hwW/stDMWO+bYx13Qyq/b+C402xUS5Xq88nHtJ5
Lg0WIPfpSlymYho8AJK2zVTMIPxuy+aNLMUC0NLmyDPZyUTO1tke9pjsteDVl2ZDGdGj1dyL3iHv
/zeSOjv+dJXRUpbAbyHfGGcasN2UZJY7mYN0/Q/X5pT7CqyXa33fD55xblwTHVvfSVyNiIo8b4nQ
1tHVuXGWgbfJLqofyd0Lk5oM6NGi0ES1ohAP11Ao1DcgtVccehtNGCkdtN1EFT0UFqo/tZGC2A7i
CPF4uMDRe7t+9WrJrZSgBHscTPZ6becpelp12m87ZEFU5QOg9/rcREUtgwdODI+2lf6Zrm3xF7gj
mTmHPtQhn5O7L2akfEzIamixzzcqO9N3FxE55qIGcA5E4qM+wWM0dV/HZQ/zqpJgBF28t4ha5htO
gu2PPJThLTBTa85PgHGpKXYkgn3BcywXYqprrP/CE3sbNpsVG3qsAWVY+ISZHL2+v5jaC0EpVnOz
sRirhh2N5h4ap17BmdhHMFn3yz79teHvJMEanKTxh+t936X62GIJapUvrogSYebehr5iTKcKZ7F4
R/JVzzN2zEiTHzaN3z1lxQDARldcry7a8k98q9TWN9MnkbJaVJVpFOm2YfW8httClQP3D3UrSTCC
zhQ6BT4iuvfbvewRg8Iw7pX+gEK+wujue7d89MidM6BEppbhFScn3jbDN3O05hKldmVvlsYRjnc5
CQkp7aQwuxOTohPmpQLa8B1elYpxElPDxfO2hBVbSxa3l0PTWbmkIoKZEexFZdfGTu1cgK1GNoT1
kV6kOoNPzjxYzIoEAxkcj5bRcdDHLVbitMpRzMtUe+U6kDRhIS7CH+2NQko2mtmrFpcX0ps+xKRM
m/hb9Shz9chVBX0vCzQcZgBfXQAITEpq/wXONgKyUHo7vK7X2Oj/pYlXw7CEgBimVX7tUWKUT/2l
u13xtYSF+CN+AyLOvkMqEmJDm/pySlc+eY4ppm6YGrvtPJZ279d+Tcri/HQvVOtXvUT3HOniLcXn
P4pzylTuUumLGH9BrwDzGEKi3hhhpdWDgayBlsS5wb3YHn670DupEag4zY/t/MrPXV4JcefKNPzw
ems3gWoJkU1D6fBNOG57buAfaoMhEvd2ao9AK+vLuHoIIKOmK6LMK85fMbpmVvXufVZyTzuaJA7H
IPz55qhkVctUKfLc5jRDNE0MZfoaX0AYuEZ0vrGEEPug015C5UvJBK5fdLjUdyke1oDab44UbzFv
5BE/pAu9++/Iozd7n9IUW9DLNs42+z85zmwDkAhMANV90sKVlcLfw6jLjTdWiUPjxFp9Swp+JIer
7j0khT0jPN9EYw3S7SWy6uuZULSVgIo19Hg+ugqXBr5lRzqwi9kXqkNIMpM39iLVlwH8R9xCVs9w
qkwl7aeV0zWFw5+JFkZ0L1SwW+LrvtkNmWBvPMiue4+n9rB1Per6dYsYkUUxNUZmEJd3z4XUfB5M
vtOmD2dSCGSC1oWWRmwAsFO3VwfL8suQG/qzzFnkRy+mnmh9LBqDwTHoin6kJ/cuErUB7e5OcJSC
+weMG3VRTJbZTuGI79WrocN4UuSgec3Qa71FUEYFPDwMrEMbsiWn0klJ2llACC+st2EY3DmWCVH+
V83sIhC8jkMnpPNMYX7AysFM0x/u0rr9T+zla/SepUxB0TdT5aEP+etNeOrKRc2XZ2CDt+t50UgF
FvFmxPxXitRGVtatG0cXbVjKiriWTxjwwDYqFM5atcO3XLpErmICV6M48074dwXDnU4e9ad8KB0S
vrqRKTB59b5FgildxVIg5mxkF0NHU2lHN/gd2MjYCnfIrctNe3XzRmWtf+ybaPpgAeyg2VD44bj/
nGq6/ETjgit2HFkFoVJum3bAtqPEr16dDgSAoal2cAgVeP/AG1nIClv+rAtsqOuPwUcfvKexuLmJ
YZKoyQI4yzvHVvLq9mAF8FioyDJg1k2grGZTlOs17OLRk8E+e47cQsdtDLZN/Kh/Hwa8f82k4wGk
NsNdRryUebr3fER0wmi5OBPQ5xEzBUPFNx6+ZpUbFuXwJum0nHtUy8HRyj4WZ2CzTgw4tvn5kjaB
RidD0hZbx2Qx06vmwNXP/oQ2ChyNRjnKIBJSzdbw/+2WcL7b3qsIPqe7oauLaa0SzykY3gXu5md1
V/HWWeTnivMzFDRc8PW3SLA6WPkd4iN9cQd1VWNTF7WbzLGRKLizpN4CdD+NeHBMwFcG2xjuZ6xn
gErklA53xRLJO70+u2Wgz9VlJFpQDoMaNp1Fx04nVUb9TubK8VbmaN4kGKNVlIBFzyq8Jb4vB08R
DXH2n49TqnoDaK802/UDfPwdhj8B6tarvstcJzwGTvyA6Mms/OybeU6GG5gfnC97xz/6Uhagkdgh
OGHh4EvkhbqkJ9V1LXtITo5hMNg+owBoeys7Axtr2uZvwIKdanjwYMsP7J5t0zDPz+HTD+ejOgO7
If75ZCiklIPGxy/l0WmSXBDqUd3Ad7Ics166kVq2d6ZWA1SXUXixjktdqHYJD9AkcMkmYm8nG3GH
QAAtX4R49i2mL/v2xuWORn/gch1wju0439pbl4OGENwW+FgaTbPBq16iM8a2b+cva7cMCAFNu8DO
ike9wPaZKI/Yw70eVHtPEnOdDHujvI+EDcv8JAn+DR0CpJoMaLnSQPi48Sc1Aha8VwRWg7Lfc3+L
ZuBp9LhFtXjzp92cC4GLQKCKP6ZcCTCJCZhxRDCn32aB3IEsGTlZjF+yKFI5Hd0Cc/lQ3xjwBjeM
EC3TxdNCVaQZFc5pdnejzUVW8zbfRRF5XsjdpSgTq609xR4vh/uJSq80yLy6N7K279u4aXkF2k8T
d1jShsi/Wj4IiB9qBBNJHcaOK5dn2UsBHrg4xiYGlXyBSslmUfU6r+OUaNhNuJIqj9m026KWlFZN
KLjd3/lqchlV8GdfPkP8/KVJnfNnijlNfF4/Bcvmz0Hu3EhoQuQyRao6h/Zt/07euuwQvdHkPeXD
X0n5I1Yf2Z6NIcIuwJkH30i9Ql5HjPjUmkuq13vFyNaE7mSuIoF92hDWAwp510OOzpFJtbk9aW3P
C+zyd94jkoMnjiqQIIYcxgETwzKCAYaDbYuF5uEbHc/MNXmDVR23s2+LmYvumLVVyYNaoZhGE9Gv
Lqui8HOw1bv3YBwPwwokkPEiK/jEqClrtIP7pEAPZtERgCGxkdONKLPplfcV1cWX/b4CgyebivdZ
YKARrGZzTVNDzjGLKvrpkL/qKrg53unVL6NvfXDH6kX5NUOJBvirMDRQ+XfvwgAsAr8dXjp8pS5S
EH4ROCgZloXYpI0hsQkJMuG4nW+Bsu7PyC7piN0ayLm1GEu+J216Hal09P76KsjdRvwso1CrQfXH
fL07DruxKGUP4kcL16AvF10zfzrNQjVhvVyLKrRvGaoERZHFJn0Ji+0Y1xoBWCA94+5B7tg9FA1Z
AIb99jx1DGoMzFjG+P08B9BLpkyB6p4qZomYYuhrmgSXbQcuUmONbzNm5hR6fbdkBpVSUqCIACo5
Cpjw3MSisrz8/ZdLALvaliunbnh7NdPyzUQo+wnL1re5hZVg6Wuvimv4YgR6UFRxtm9SSfTdokPv
lys/wllQ/gZp+nfoUZ9HB4NrYG3QRt+kL7iq+0gsUdFhU0WWx0oB1jtBzwWzyI3vgGOIHIU4MI+1
lJayzNilcq4ftOXgcddxfSVwCPeTse5r2t2Pf/GJrezpPJkaALSuRYhAakqAnQ15WcZRXyQXabiS
QJ8TxPt3YHdJ+l2TcC0w+lM1/vRZkfWwwRob+uT3fGic+mWGGBv8kQae/Rnho9EHwD+1EHYwliGk
jZGJAKioruhqgkg4R7CU6XxXTQySOejQ6wqCEWHObMgKdVA5eg24KY6Z3P8JRm2gGuRYGQC6dXdM
KKcBA6KZ1YB1m9xvqDjEwmoeWi/QqBNL9x3G0pur7Zr19X/tsPVek/bGL2p/E+9++exvzTVUv4IM
YsI6guVHeNwLr+oQ+a3K2xPetI3t6pSA+xqsqa9Ead70xrEDTNdCcunlqSttnzDqicDA0j8qbRQW
OXD7cjtXkCsZ2K4V5BtAUJO64tYGduqQ6ZZjlC6dsS9D6sFyIL4uGOVjsQ7YN8zN91e1+AyDxO3X
KqzMr4eGZlzMfO8y0eRHZt6Q/1WLrL/HEFnMO4HTletQ1FFo709BXSDB5Ob17+f0yQBZ/35KdJC+
DNv5ibkTTt4/Nkd1OvN1Pcti63Tblj7EGL05GgkKqwwQl7qmxD+4+pllLTscOXLrOZfhPM3chCzL
uiLlRLj9PzczIOAdhyIeYHUjhGrkeYePVVKxLWliyT83rv2jaKNiUubHYwQjPis9jcZbK3MZK9oP
sCdj7ixd2ikFftVqp1n72Ie1ibTYRaOc7y7lTZ+WxxVxR7i5Eh8KSuv4A0138PjeGOqgJR7Q+0LK
t7drE8HBJIkfUVxcpI1EIhrD8yLNDv1C9nPwWZifHvnNQTnA4/HPmTO0m/2XyvOA7Lfhs3s2wJ+o
qoXW6yjRLz0KcqWJCBH/Pg9h4qCfAPrLkSwiRsvtECsxYD+LuaBmfO9RP9RdLgxbcv76xbDDNNkV
D8rUh9Bl6VALbcXBlBExtsQaymDG5SMrL/nT5oB4ZUqtpo99RpiEeAjBUw2mv7wPeF01L3fyvNfA
4gGTRfcvMQXrM6X/txed+CzgGXe/7A1IBfkANRXPDJrxN9RySKNoRvL89px7PQDKhwNve1iIvKer
QW9yULJaGG4KpLF4IzLhVc3CUdbRelZ0GmMz8gnmXycYH4JR7ne1+E5nzB62qczMuwDIkIqykGu/
YoIGSvcwPGJ8rrRvUq+wYKzEFRX28tb1yAXEYStqqvjYT0SE81wabGP+kVggMqWpoBLxebyntTVK
f7fhNBk1jESgFcHJYW7XlzAdzgDFi+tr9Eb2pTLVzLelpTLWwX9ZFfxGLsJvLD6/UXLgR+GY4Bbm
peamxToUuQjN3YoPSWQztzEOnX8DCD8JQJPZZpdtPbLq0PKb2HDBkDO7aB21VFSAAXXWgb8ZPMNY
Qvhwuy49KRmmCPInpX9onZscLdH2kNTMFT01nwmvsoCOyuUVicDDM4tRLc2X85kEnrtyw9a5D/h3
6gJosoOYu6ycY3nOEWzx//ZVy7ipNaTFxPD2+1X8tCaYE5bq3ib0k+tynKWF7dak4f0A60EgZfUR
hD9/EiEu96TOPtddsw9lJoZ9QfOJjrw68jAACoRT39TG7yG9cQt3KzVLvdMUXoApDi2uBlWkSgdF
iQGPE+Dkbo3m5wvwylbBFXCfJShhCURm+jyCKxsJG5hwutbJEBcqbghPYuOvLLtGcdtu0eZiNqhQ
ticHA4Tde1CDHsBhX1rpxJVo/gAdtq1tM0OXHLr1Yhi5bQV4EU/ZW85z00zDCwGLbW9T4tyuLpvo
1uafECztJCYg6N/+A6QgokSp5FBP46bG8Bj9LzdGT9JPSIBPuUmZOZYxhuJtJwtCjUFVnFW7ZR3/
+QlTulUNog9Rqetc/8dqVC4VbBa7sgZ8hBexeNsuPsvY4DE8Hd87dV/rqW3TEP8sY3UWShfoVYYU
d80m1fcFi5QWcv9fa7QwE9IoDf7q7WtBS1dR8Ig6CFDFxwQvONReA0ne0UVQ7fSVf0P643/wmyZF
u32p5ycQY3QByNzNaVttU9hknbFBBpqQzLaLnaKM5qdN6vBJAnBaxzS9VuO6B/DWxm4XSDtXN/jT
xpIwRg851PWnipI45B5CyHqZ9vbaT/66aGFYgzhCuFqXz7eZepQjYBcFz0SncXXZ2HbzYZbPFfjX
Zo+/QihJl0TGpdz1Df6axynT+vIeC3wIwn6jRDD8rPgmr9rpz8bwf3kUckJM0JRHJOvMro6911TV
kW65gSZR4nsiuo+HnKwZQlFGdIoq59isrswbHDFdchLLs9CzDIelsdTKpz/91VBhdRuBSMHsagy/
kP74HewyWHUmM0zZy6Db5vbxWjyCNKqZvZ8OnQbl4Wvvb/DUBxL3mkasTwgZ3Nuz6FDUxmauceYS
oQ7yRogXEmerWAGek8IPPDFy+j19NQ6VlWr3By5romSFRE3f7bwCEepfFiBSYWku150kOpM+F99J
6DUeUKjIRJI1DBnUVIK3cJz4L8+W8I8ys613TQTfZyrChzRWeorOuBks+BbuzdYUPq58IT6peDEk
96QFpZ4FgtkTxax5HEy+vdTPlQ498vfVyOF5/4g9Lw0OSe5l5e5h99wSSREjFqppvSB9eEBCZO7f
AU9MHxnrUIIzEb4NXD2dPmTRo19LfQa6fR845ZIqXoaSiaRhHVpWvXSt7szlBbeDHKWkWJlJfQYs
AI9Pd9WK1JiDQIgoR8Hqzifa8KoqlReru4++sVg9fpLLIk6Fxqpl2WGAcHcuZIuJEXcVTRGDwAOU
+ju4urApF6SWLokH/qGjPEJEZSEWL45R6fPprGC3QtrA0My86JBhsmaYtWAkShHVuqaMBrMK5Mdh
TanU7p6RIPAHTeGNyZoPjmmwAv9MHDY+7TN59uJVK8trhhqwhhBekqWQhBK81PWZigm3oZ+RGfM1
WIztLbOIL1Og9LGNnrdFIvZUA8cv6xY4reanGDn2E7Cc/aopVGSvIkKka1/EWhNQX0hOQXdJBDz+
wL1ex20SwQm/cNElT1sx2ICr3qnHCM7DwSQU/7G5suq2gRuYqTdKnwdfoalO+PaNwWn2Eafm3nJj
m5FudXAlaLt/YCvILToJy55aSAwsB5bLDHadEmhv4XIYeW4D7N0x3E0ziwmg6sDt1M/vqQr3LXH1
XYT8PxKRxE2KiV9J2hMYIxCIuTpQ4AAylmljI3ulEyl5w09KwRI/uu2+nQf7UEsb4MYX/248YTiD
m3tjjbxJqsEnA1E4UgkV3TlbSAVOkpQMm5ZlocNjQMj/bORQOReEVUSac1t28l+nIwhMMHsyjvOV
2fkrhM1pVKtDHq+ZIokupdSyWsfnfcdealqhdQ0YhsU2fzxbBOplUd/0VwMTkZmykpVBdrsUrO/O
xATJNx1ekY4XvPS6xQ9D0A5FhnZsdvHXc5Oc1Znf534f4xldQh/iMx629gfXFQ9TDL12JRKdwiWH
DhSdyhQJ9DhxgqxDS0QObbQQq8w10Ke8kdKKIYw+QvgqalhcTdp0Tnrt1zAaHIOiSiGnP6I4/sdM
ESMYfEWIv0Krmow0/AHvGq2ttFqSQjSsAAnk089mBCr9VGVXYuvktDk7/Qe6zIQ0Q4ZMgPIa32i+
xYx14bA8rp1qOgJRz4BVwYteg88I7YD6MJYMGBfE9wKKJWOj4Gug62b/R/Jkb2SLYq+1AX9F8HhT
qrUsT8TA9UxDd7pVD2009HTCU8GLdj73PW9sGxm0JZaY0ve0oUmbO054ChRR6Lw6N7GRbIgZ8K/P
faT1L0dOGS/FGtct2UMaiUFWMeieoIO3c7n5fThFh7BlWIzyGj00PkY2got3IGRXEjFYFJn1Lm/Q
fhNN7xxXfkZOGEcoNtNsSLCae9YBaSIlKVk5NT5MIzdl1wmNU4j7oyh92u0Ah3e806z8m+ibj711
9xgXUWDDNyvBFBfmbSnV8BNMEUjhZKuWp/kecIBu4Sf5p93w1Hy5HKLe1N6PPk97pE1R2fY7z12v
epexzD1RDqfRj9yL7xwy7vyGpWV4PL89mEeH+CZs8+XfAbpqWeiDdlnXZYmueeKCDZhQn3kG8juj
tduEkSn/EVeSTuD8UCPnVXTfuIwc2M/HM35iE2WxYeM1S5FLKT2IPiT3F3LcwIQkmC/4ut5dsbqB
Kp/LoSHPXaQAPIO5PAsmPfMBgKv65JTdwYsSvIrpAiIkQHMOVChN/KD1llG+Iu8nvJcJghFJ6kcw
x9jurIm9f0z5a/r02w3wyIuLb6G6T0nLs9dMlKHYRxrL0SrnwYMLbSENuMU9EoWG0HV7UNOe2yxA
rvN7BkYVvmVQS4WWya7NSa4VJTS6yrOCcRdlvW1Qfhgw9DarIYZgvpaDhcxBlGdhhZ8SRCKVchWc
+mNCLAXa2K1GYi0hBagm7G1sKxxMDF0f/8NKu7ZVG+IXPgxLfSgowz8E/rpZlsok9FjjGpQNdj+q
Lii8S7Y9jB8nlUNyp3irgPuPrREqh9/OEDkGmEtaF3Hz7P5j+DSLjHwPL7aXglDTZtqizcsnt4Au
GiMCzCSI+kofAnffOEE8HDL3IwlbavSAY6eMlAgxCLe6WI/JUm5Lm8na2mke+pLdgc0LUy0cr1S0
k5SQWqdmez1KPvVqjPmiAoVgyO23Bz3T/6PbZaa8T03ZEN1nOix4Fx/7Bn8vbIFcU7P/saj90QaO
0emkq4t/iv1XcX1+PBvHyUC5TRub9SzgZQolcApqg8Iccs5pCpHWcl/ERXp1RVkzlg66QOFlzWwq
bCjMmDvkUoqDyhV1F4VngFmlFdeVvc1FUOjPEtRVrb4OrQoV3XuqQvOGDEGJ+/qSlu12+CXOiuAP
2k74x3n+uHPeinuhSfeAwYcWFMFJz4Y3ZugV/3tK8mEoNoXvTGdIuZegewW4mI59oOxEUu25gDZu
6pwkqTwcb+3GLceAPWE7r0B/SKZRw3s4m3Kcrqxu3MQdh/8h9Xt2FDAuLBbTHyhQgFLteJ9Ku8xJ
4mHyVvIyRAtDhFgZVjWrj9ewe2tCgusUO8S8+bWFMdH/uS3YaKY3tH0N6raJCoHIJkvMNnAWgQ+L
clLeALpv/fgRRWJXuvRVxXqBiduF+sGlmStaPNyOk67xolqGlJi921TeuK88u8uW32eqEwen8uqL
QGmWyKhaZ/OIcjYamQXm6KHLvAVWYWDIexrMJuZPpqLvnTmee9H4zGhLK2ynk38ylcHgRO6fWKUo
+6xxKRSUnhFPSXFf7l9EUpSV3y98BUV2gt0x3rDosCIAz40TejYRQMBdcr8V4AY1abzcdm4cFoDT
a6C7NT2cFZYYHwHBibGWuTke7glKyEh86AHdeKHmJw7fwy/p9xW08V4V4LTs0btAZ6ZIaTyJgAow
fvcXPzzO1vIG92PjEp6Xy8rJpwYj5IT/v26a1dXHq++EUB9/dqGKJD4iMsALMS2MNGrBy17lrgre
3koQCDMNgoKAKUMpv3z965vztV2OCaQnwVROGIIr5PDvLkKKJJZPvmBVSlHJNUNf+llviVBSpC0i
G40Z7C8k3eyYuKhAwjJxKoqEOiX7Dp94L7qnGV0WDfpVO44rFIGpOt+bt2cXZBY4TZZJgHn3NBqD
bOCM8VlOLURB3FVhMgHNw+6iJZ+sz+12LtgkFw9neRlKQdJ4H3RUjP6gZZCLhqnSa0tZeOdk1b4v
RhxwViwsRu0uzsXOSpy4KvTBb9XkjJJnSXyB5hNoAu9cynMdtAQa+KGX8NEqgFJ1Ar6DMJkYXjE7
F/lyv4mMjXAoUj0IiPdyiHqqGVYUrpeW4VX0n9zY3tb90QnN9Hh4Lz0z1VDkH/RlEwyyyqyNCd99
tl5Hj8RoDwmKTjBnI+uARAYDM88MyMS0ZOsqHndjZQ3ZemASur7f2dH7eUzeI8Kc1e3G139A5jMV
SCEKm0HgKiiUMv2d674DpM1LusFpse3v2fMuAlHqoZ+pxFuYcb9wvQ4IHS4Kn/5VGvgCrT4YNb8X
dz9Z574oX1+XfJTLS218YHQbPMdJGBnz5F29xm51BLych75ot3kDmAfrAjhR8A4WKuVopgirXvBH
nmYzfkiFujXJMjBf38DzhDODIKYysajG8zJSOfR0biiqgVQs4wBgjHjDCSPXYoMg7pBlAS4oeAwu
9//mNnz6lctq54b1XKpqkisQBv+xjM/GffmFOunM8A8fx1i/5TCGx+MkJXxuKrd53tHgPeF8X0f2
1AVx+6LWjfsswwVK6TXMsvz6NMqopchhpGWPeNRQqsmtjjhmU3eNuk8MMxM1vTthTuqM8c3BHokW
TiFdKeCRhcja9Zg4rkWWZTbxQTRaK9ES3jkNWCQff1/SfTPvsoSQAzTs8N7kRLMndts2Lc29s2/V
ZIZDHCxJd1LNjV9iWg0dLsJTEWsVFUTrBxbsaOiP9o++HH2EPpaxHDpQjqxJU1LKf+dZCHVpSQnE
uuXCej+BRHG6UOUyyxkqDGHE4RATBlqDdMaZOMyJNZFtL8zdas7LGbilScydKh/gb6kpX1fRrJO9
eU6J/lJht5geDpaPAKlGIm/yr50Do/FhAMDUACLcCmVbFm1/kVYVBz5SZIPOFsNfzhMOFXBiDVv8
FRX4Lvqj1FSO3urnwRFnpXOjOw6mL3cRxIazaH5cLTj92z9Sy0VsfVW1nmiUPGEDshgvqc0g+6TH
zDGbwx5xCx2O2qM7WZ+sj5j5gmemZWNyy7w0KylK9Lm1DLKMSSBmXVhGVfDu/bT5d8KqVPVZnW5i
1lqD6sraKzuakOdAp/4fX3GJxA5Wu+62wDy7UKb32e1jBeoAYbrpwWz78z1dMfq31m70hFvHuE2I
lfyuUwgI/YCBRMO1auuEX8iut71Qs1rzryAnKtB0NWD29JJTB4+8BbLhMoFfIlJvIhDT/SlhuzLZ
agob9M4GlbIFnP5FchlMWKB8X5fDERHZaUCGqRLUjxOzJIKPQF9BWkvOm3WkFMHnOURP9sOT+pc7
iK9wL6LLZH/u1jW+Uub/hhDMuL+6E27JGlXQ/rt6XUE9xOk8Ikfv/yHGjqfpapPVLsu+PIwU9hey
5DPJUc9LFQEB81dsE6fy2nMF0ZudMURKxMv1uOhmDsJ7c7ta/i4swDft4zSBDV68sBPbmz9aZYtY
jgTSBcog6dmRfuoe3369ctP/rYtgk6z4CEZCxdH/sqYDlQla87q5RIQsy17APge0zRkQcisSq2Pk
DFlM3qkVfzslIsm0bjUurErHzMP/Pdn/PuT5J9Y+rcPsndFFT7ObxxgO6UNscTHh+bg6nsAg1zJS
LIP/Mh5WJZmx1l4mp3W6kc53+k5kmIVP/z8bYgoTSyLNRJix4bfmXAMJuxcLYdTCiITrWuk/nqji
71cmStE/67/I9EJrj/yGS82k7LeOu8Ig/UK3adsT6TbpitFc/Dvq4GjytC3EbW9lg6hyy+rugasn
wpHT8m6yYsK9LjqSt4Z4298Gg6Jy8t74V3nlxDTjgeCM+bEUntz4w5G8kjvSSNyF6tnQjg5Afwyt
MGoe23Z2DeagiVwYfhZKjKxhRof6Yuy4UU91SxCHmYQiMbQyyATXaXp8C2lYHGqFGzEDKUG2Rcx3
zJuWcT/8IIdxCQYV+fWE/evBTGzZ7jLjCYCGiiqp9T9nKfiXSoKmEybGzEVc1YTWplsMJtvh4Zlj
VCTG/u8wMMjGbFMKdyMrCFlFOz6CUmf6ugNSHagWiFKcZjwlnXvEKycP1Tk+gprGKkgHIx0CdFnr
GHU5Gt1nBGXs5mvmnjs1L6fZkUmMAN57hrCoHg/5i8j4HvdaenhBUN5VAPW9aqrurkPsh2GiYJka
fiuMOhq2LtSmqK6jt3RzbKSxaPy+lmdou+Eb6zkl+ZxR+8h1vgok/RS9LtowCKxXhi9JfWmbZgOa
3eOvIQWinfWPUpnL9CpoFM03//FdE8BBdpKm0dlj37Ovls3/C44LFdr0Xu2acNCMpfAkkVbT5pDv
ofN+fpRAdZ6jVLoORKeaEW6eKMcrDZWjMYqkrm0RyGK3UUrTHWAmhT27DBdTWq9BE4W44IUhHCaN
lxYUwm9/XJmwXIoYh+vVDok9rG0ru/HDs6bemNbOA0VZ1DwX4jsM07Z39fbC+mUVl3eezyvIlftj
VExnlkraT7c9niOFMnzwsQMq67fhm42qV5tBx7dJTByEZHGbX8f/5qh3rWT8aj/xIx2LQnRoWFtO
DZPwE0v6vsTi5QE5Sba41EgHjJu8rDEIpZhE8ZutbZ9FYEGBsM/NuNndbWLGRDsr7pvskNQJyQyB
29bYS5ql1Q8graBva6tDfLP79BICzmzrY64mCHw2w8f/81wo9xnsrRARYXDFbV3Pn9EYeFWhpdpn
jNVgpLvz3bfHYRauciA/SNIA2/hUPqtU9KaF7/gkqr4mNidcQxZGR9MRT7YtnBnXia4xZBhQFTbY
vy8LZbcyKCRTcrr+wPzJFj11xkXIs4QAV1Q0Nqo7KSrzkCpzOiHfCwTh3UjSWK5aTAHSD2Hi+6IQ
z6gKu8r81TfNDv5HYTuS1xMC5HiNaIvT2ZKc4ON+Gu5SobLMgZh722O3csdEN6wZdJGZgRH1rIy4
9EA8MyWShjaXN8/P0RcigafavT8P7riBesJi/ih+Pckf+3MviQIbfbDjI/WaQ9vSzIuLCTEtr69b
X7+SjWFBOPATX4Y0suKeTPdBQU2awQrN3DlCc523JcJX3EZJwacE9GUsP3U/FV7AZ/yDVfh1bqqR
jCJM4Jb1/iWMgakR5MOzq5liMLuMdc6LmZRlOqzX+W0BdU/tuEbxRYpvHWDXBZwVGfO8idrZRNor
JY5HqBmPyu8ZkBhyKrWJoiIYxz0kWzTDj6x8gsbsXuaZq1OpXqzaFC/V4EmfTklm2BQYoXFTmzu1
Hmk6wiOWyvQzGU1yf372P5C9ByGVZWhmQenFx0a8b5RZvWxiorIyXGGdCVhp3tOsZ7ehzBOpEHx7
MHOQj3GOzuU4deg6JHfYw2rfdyR9eKzfeaZOtSI+5hMHXsOEBZmrdYTLkFptXSrwXMQo85sSfLb+
P/XqU7AGFlCEC1Q8J7DWBn2dWzCU2ZFD9ooJtC0nXGRj9VB7hqcuf1pusboaXu7OVCD1Nb33tUTJ
xackChebXj8E8wV6GxYB+42a4kTF73X2vzb5AvB4PYjMoxC6XHzRTyCszGMBy32WILk7rCWprmIE
kwozb1AV7dWj86O6v6CFj7P7lNCPuFlEw3lUe7TuvqhmeskilTokyvWaf50TPOyzy1HosC2P/Vnu
ScBd6OG/3DCKQIrMFFCSNzJD/7fCoiINUkE9wL+5EQ8GlqbS38QSea4IsutDyRfIF+5ZUubDAKxC
2N0NDO6WgYjFP2CazpHj7zMZaII+VDMUnyQtP0o10suoaV015Gp54XguQ4pT+JJrh0aDwONg0S/r
Cr1d7XuCNKqEfYr1/f+6qAw1EgoS2J6G+w/mVEV1jek8tKWNlSEbB6sjBISmSyiOZ5H+uAhQEn5D
2eIJbe+F1HGqMYphrC8LgOqzYyBe3dV1tNfNtNckqLpKtycKutdNsCUAAR5S/OqQukfcSkqQVVoh
94lHoThWQUb7u5iWzJ2Zgi1A658A/P3TZnJbdfR3Q8Tt7ePfbQwaIRIDnz7s7LqPoGKzjuZq9bSu
1jXsejE653J5DxP799Quej8fki2dzLBMog5f6lB/sNMyqP0wCUlu2qiYmtKhBiEyAHxCUI7MoLUd
+LGtBHd21cVSHIWRtjM2ONfI654cRF691FZOkDuJljHjGOTARHKd/FquYY+b3DFjAJoZQVZbbJBb
M16DkbmmK2eTC7cNRbu3S02VWH8MC1VAzxpvPs5c02dO3RSjeCh0IW7dutyweK4HNG/2QtCNSori
aNKHE5dM3osVkjXhdH1jdukoF3s1EEm1d5LAzZOOrpP9xQW4e4V4TyDnMb+Xm9ANz6zCDfu/QCA4
G2hKPOhZg5VQuSKRhu2ifdZR9W+BqNW1amwFejajWsLsWqfKgDp3/HyUQIXonFfcr6kMH+L7jCTZ
eehLETvI3Y3CGFQykDm+RreKBH6ROTceuokK/Y3EZn9vvVOsPAOht9qSWv9Rl4bYaDmXkeZoMdvN
rUFbnDZcbYK7mxUrsNz2JNm5Kpa83KBxwInAN/VwI6IYBSLP88gz4CMPpLw3uuqvANoG+BVLO6qF
qjpOvc0QTStTVpOFg102xQw+pk2Swdv2fGH9U1ZfghKLHnHkLcr3K/aNZUEKgKihjRL2oWiZK0ye
WMUnVWFP6eGcjyOiNXOP/vBqe+Bo/puGztYYYuiVQ9QFPKvhKu1yQyD96X4xkzmW34gZaLTuOh/x
uR4EQkNPQMSJmwflQDJNcR8OdScB8H+IjO4oCJ28TJCLWKyuSBTxLM8490VS6ED0JManonhRS4Ka
ZMyUMUAz5HUWiCaKc6xuroADKaxNQU+AokDZp/3iJU7pEUex4PWOOwlj+F3qAPICDqEUHhte98OX
n/gAe5Y310B040E6eiuHjLMhq9dHONJVudBqMopTPKE+II3n/zZQ6TeXDa/n3uCDblqLqslA7Z3I
+RBWi/3eZw7aN+X8r4ENOFLI/1/9Gnc0RBDa8tlsLBN6PJmF0gy0QEf/3BNJ60wdWnDQ+ZVfij8A
mkpne4vv2kCaelLdu866tmLBez1iPUOWVPxpYjWAUfsncA1+c6lXWtPTFmQLePmpiXVO/8sWFmdW
8GVAh97fkhJCmImZpvzcchUpXHRdbiIGhvT+rRPeKL55nhfENp+B4mXBnARSmLZBSPUCMPWlx2/s
4rLZfISVCmLqZ5vZ287ySIox2OSJPI252xHWPvY+ZkEvaEdQf3TLVXc8R7Z9Upt1PpUyq47mA5as
S4nnXlHbwireeUpBq4DUu4ScHNIq58obDjelxrwpBQLUXX3JdebE3Buu7ZmY8n4QFyrcrnHXqDci
WECD4fduoFXd5IutsbmKFND0Xz71XCuqz7MraFc0oIveWLEskAImJQWOpHkw/fi5IDqeVTNuKLXs
xywI1NfYx0SD12v+KMxst89dgDl855DiVyrs3GAnZji0CNL1QQQThGqT32VENTKQyDlOLhygrz8Y
T+6/P46IIUl/dwwgoLHW+n2nNk5+SQJXxpevhS9jdKMXeUL+C93BSmXO1sa/uoKWgWvVMN2xbN5F
wt0PYtjosgpGEY2tRrHgCs8F/Q2oSMBRwvLTFR4HBepkWlR7H053YuIXYS71HoS9owuONi0z2HPR
BwCjrUDjUe4rBQi9LdL1Pa1Tuainsxu+i6VKXhs1JBqp/jzJNUhOpOh/IdHLastu7b2Vi/YkfAGA
xHum4pNhu1KfLRzeLXdOhlDD4SaSApouhYtW0o85Yg7CKufqt5Iwfedlpg/9GE4pZ6y4Ah23baNw
3MMICBcXqSY7PP/qVfykwE5lrxE+dlYL7G6uixMcjc8ZkayQ1KNvlxkCJPhobsAAjZfVRunItJRO
Qd0hyo9dm1qzPlDbgAZbJrgXEds2N/aT69nnhgHmHRMVNOasxcyaaoZpox0ujK6mv4U3W4h594DE
XWkhwTrFwTP6voJuHwnSnjXFjmpqOk0XokHkbuMTWiGwiG1JBBtUJMs0r6tcSNA4ppnuGjb0oqxT
5PuKO1gnd52XJtk20uuD8ilEAbZdCKZ8LhwbcP03KW6CGpsEVzy5KeiSdRc8wV0H6uzRe+YH7IhU
Nu2RGbnaYV1vZACzULQVuUsUQl8UzkR8e7PTFpzUeOANYje9PHS8L9KdY324bAvIEDc8ZcoXxfuR
xvOxGFKF+iux6MmyDwkGe+Z1stiLsVzLJ0fb8/eNZSHlgEsAgTwX4pkj6sBPWeROsLxs2EBw0+DD
hzcrjciSLR1b9+ql+R/6CQ+IQIbMvQudpw4rDqtAl/SWWvAzCNQIiBtQ4EFP7MhqchS+JJTz9BKF
BHXN42y5u78MK41KGFL3CV9JJPg22yugMIp0rIYZ6qUH+94Obn4AsH0/umpuaUDsYE6ztzhcGSHZ
aCUxgUwa7ovbU/hIY9naBZwRv3UMvWZvd9WU3i5c3wo0R63xEFLUO1ms+S8NybOWNEcFivq/2Y7O
z7YRAIV0t9FK51tzlpEFJeqAO3H9jaEpmNsMCs4IbI8z6lQJrpJkz1oS2l/vLy0nAZrcC69dAEsC
VvI/VmxpkjzaTa4ih4kNkmk/hJiZMfesbYCJTyaNpPQ4BWnHTIrwrC8jYyc/EvbeUoTXOE2osoG1
6plDw4vXVWNA3VeLkkwQ5IMyZj+0dHUFm4psDKZ05HhrfNeuJ+qZ0EeZpG5SaacFz4JWRBsv0wSs
lDA16t4HaNOJmUMQV8+/qLa0H52WGiMkY/bjVezfiPUYwmsgp2rj7nRrfsw2dPXFKYHJyWoUL4bM
Xr8FGB2crAO8r/vxnHIfXfV1bqKgsQO/7VkFWrOuTXLlKe3OcCtHmB7JQdNyCsOY5GANySMvGvhk
xEXBPsjg1EYrbja0V8mxQ3SSjQ15J24w7ruePTSunRcK3OzunDhb5f2Sw6CWg7UIGVIQGMEfqhPB
0TKFV1gg0vwGolLMgLhrPr3p3cLEHf8yV72PEXLWHqVFWibhljr9xpb50IWNaDotvfZW3ApP1E1M
Zj/j76X54kc8IRHF+IwGBMVIfb+Ymsb83FB8l7y5jVnDEiiH+Vt66fRYeCJNOMp+o5F0E9ttwoQT
XFMLOTqJraQhWiTSzaPmS00njT3rfR7U76oEwH0vjcVtnH3N25y4m7/r8sCqmLWPhfU1nk8uO4oE
G1RDGiA/rKnZWjhIj26U1xG2jtaZO/g+I1seuH7OglgLt+8BYwd3lHUph1fD5wc2FCxt+iD1I0Q2
rV5wMMkfY8+M2bKISx0hn0jYsYlvkmWpzwqYx9l2rkpEgacpvW+E7jlhh61Uj5Is9JO8j35k/c5s
GsRB/wWX2L+NpqUix4355BEkwvooz9R9EfSM+mSvIcL33aHyjV+fhZQOVH0sv1pgpkUTbGntxpzR
F56NovRxbN6gHaEY+hkQbhntfZtHluO3ri+4+tkDachCtHBaMcRw5adMwCOk5q9pye/5zgJtCyD0
5RFx6RRroC+BxnjL0PR6QNGtQIwfATBsBzy5HuWo/SRN3ImMrR3RxHHGuqTY05db7KvGQUequUpI
YXQ4CmJHfDE9y7cHi7CvV+lk7WLl6q1TZ6DSofDGLNaTLSEHkEThfdzPe78x/GgIhr31Unbg9R3N
PSPyhqO3D7nk662KxFl4fO31bYa3TZGh/KsrlWIT6L2kagjNNEB0NyOeeULypNa0aNjU8PhX/7f3
W9KocaoMEBv1BpeFP6BZVrJ79LXZbc4IqZabgRSfV6k4xEtXCYdv5d3QaDVEMnqUnNO7jehbsRp2
7IZTDt+/+L+WImUBhbpNbzGOrY7lmJ9hwU8t9aKnDAuV8KISKeqhmorNxtfJZPySi9UaT+RP8LY5
ucmU2FPz5/wnnI83WrDpW7MDDvxwyEbgV0AqVheQK8wiL+M9Nb+Sol6QHLQRtlUqyFYwqRWiqcmq
ZroT7qo+q/k7vEkbpGcCdwznCMwB/hMXxNw8+5th4+0n0fuSX6qPRhGMKSDZsfV8kvtFyf8a5IhW
+BouONNI9RgY4uUC6JHCJxLniA9JR62+U8IP8tGuXCK5K/flr6F87XMghXP8PF8AlSrTi7cVB9mA
ZRBEFE3c6/lcdEYvW69taBL9gqkboOd+lBnpd91dPuyNnR6s2FXSQIVxmkEWbkCn8AX3JwHd0bPI
SMFaedis71Lz5f8RCyQVrh6YT35Mwa+9ZqroQSp7Z2NXIw3ytEPceYDqPhfexFXQYR4YXLzh/1et
zeH8vVLZDaHkYWBbtn9xWefUtY6CsYG6fJYNij+nAL3tNZf9yYaQT/5oWXF4qmYVqHZMjFuEw8ut
7rscflH7BRb0pE0u38gl6SAjc43tLxjor4CgSK0TowniQjfFKwqAHNyz195Xl9p22/Z+E5ppdi+u
ardLQ9irc+ZFjXBTbhGjYiXs+oWBC+99ZzpjJA89QpX+NxTbLPZazwk6vUKcY+W6MHxPlMo47wPj
fK9VJdfP6bvc3XKc1ElHpObUs1W9H4TEhbYjeLfseXm2EkpfY1cWtImA73ZYsoGWDvp+H8aagtND
IRd/y1AciPVhtNNKVZFTv/ya0VefzxqV9Fgt1N5HWdPQamhLilrMig4FLslcpWRR2ju+0f3U9QuY
/XovHGH9ja2WwOIddS2K8/xLbXqGUsH8wTO4ZQJMNzd910w8NqJAPzXWblj4EGY5jWF3VvPRtE0G
QuWeoE8QKwMEGU2Ix5QmICkDEwHjmWEPFW8rGirA9gZIszzYQrULowZSuehuuqR3rrNjC2oHlg8m
5NLfrYpnx0bZ4edL1jYkPZSfsc6hplCREzVMlOpwepjlbxdpQNS98YBK9FEPExuAxKlfNaoXfhzl
Wtf85IovBWYKhojwkQRT+7lh2UJmO6pnTp0uUzPQ0rNXo93S9lOkOVpXR6hdpRw4DoUTMLYCBUdE
Vn6ar1MiVCsFfZnLpUenwooBQk4EN8be8Yjns9WTTvi4QhMkQFwz8teCZvUbfIopy/D+o+sHDBmi
D73xN5PHimJU037sjhffn4K/fJNYL7yNkScJs97rMZL2iiRWhCib+iI2JwhN3hP6KGOfosFpovRv
jA1uENRDYHXxSOSPzngMmfmfCQz42vo2nHfOHHCxn1vEX2dxHeGeS/XJYJa+x0Snn4WtvRZhj5XQ
xhp+Muj+tSrZyEYMDL4CV+OkNiL94sL6VCSYytYToEMnOE8IMBBW13dhAImeXpNCJsEN3uCDHpy3
9jQkxMbDashh8tT248389XWqPO7zFho9HKofGCWvivBLzUglcUFKYV5UVNgS9YKB4ZwNRFyhNiDp
cizmgr8xAbjfJOL5iAAWJqfZpdxkQsgWblZteyvgVnhna5yvnTRwZzJEc+uommeTxWFERgnETnQL
BfvW07+O5AcO2DwMbMRgXomoCU9C2m9OFyvnES8wiOAZ+5XhkrtuB2bp7qgbBCnmDtJVRd+FOG3W
lObDAJuDokkA202oe5Er14U2I3MwXYiLrlAfAYLPU0FMyh4rGLL/Q9AZw6X4qzwNpmp77Fj97tZj
uy5cOyqQa5RVkvQakzoNKgj+5zO4fU8Wkryn4xga2ITyMIOWcrjSFAHn5nMgcvaIPibBd0ph8BnL
TOuMRjAFbSt0VuJqW3oRZ/eceTpFIIwpAH13U7q/hf+XqnQLgfDhutScck0sezBbAnpAoTD1NuxM
cq4kjTgqexYVP8PA79YWdG3BBwImtMtLRxPnZ049+Sl57YuWK7GRMqrexTXWdoUzQAWDohQ4ABBd
xDhlzxOXnluFjUUcq4oE+l0SwWxbhJ7Dw3y5LQ174czAqZIOk7kGS70ysMQirc4X0l9ACdafDvFl
qvtNYRw1PXZx0Ly49WDkU0lkBDSCR2BKiNJ8P/khM3DtkJJO3uzIBgVE3Rusz7pfEYx9f7Qjq0Iu
sHUE7Mh5lyyux/v1o3qqlgV7v9poKJQG64jGUyfP28cp+0zymj1TZxjJGjTnKDvEIWgSWdDYZ7I5
vi2XN6FQkS3PV/MH0jFi+j9mGUVqbZyjICJxz2W3Yf7sxhaveZvOmLE84vk0uZyq/e3Q8RQ2rLoC
e3rRP+Hvihgfd/Zn307jMa/LM4s6j4On+hbu9m15ZhlZuN3MPvUkgBppFaLrekCBh1hE3tJqGKzx
lvEfr9npzSsCqAQ3EBSLp78wZ7oXfaO9YaVAETPKZ6MTbBgYHy3VHr03D18UzMCxstjP4xtexm61
gSCYkFhqQKB7xfspomGa2WjTcAJvdnrNjJ7P89t8hmh8Oimg33OqDQSIwATmgjGjDviW28XOFQfI
9wBzI1rgN23ZqmGg1SzVMcdFHXy8CrPO08mt7n6EUlDGT6lFxeZbJo9NkUoOk6KB3UCwLCfUqiWe
3JWp8UtcEZhlIwD5/qDW4y0yqctJtonB20zb58w+SCczDHg3Iu2SAA/H3x/ql1o01CSbkk9XwmQg
1bM9pa1gWWgV2AAx3oquFtS/2sozt2GvbaZfSdxLF1OKenEv/UssgsH0yWz4v8Os8GOP8bqDfMZ2
QFn333IQ2mBDo1RnMsERAOOjUAEkHc6oKX4DCNYYvdTH3WL/93q9ykM5ybbYiIWI43F4wRZPjgY3
/u1PznXS9xRwLSRkXbd90FWHGhfgrjkVDnZCNjXzMNIrUJbeGmcna2pZSKVQfIwO7tL7K5Op0wUx
vyshFY75o/hF+VWOKDQ7MwJIzhmqJntpeSFK1+FFVYBP6eqBBFl2a8GIzftJRtHyjsqaEQv28EiS
rV6cBbmJ96Tqn98c1pCuV+rpo/HM9Ilu/CcyCLzjljRDCv/74AE5y/LPOMq5TYhXXQlsnNGdaC5N
7pChCjZkznPFPthqg2jqWt/jV0xyqaON4VyG8RHsNv39W78G/ucM2HKtbtfak4t+aVCfVfCUR6oZ
86BfDai+nQPsP3kLckq/w6Sk+K4WOMaIwKbDN3LRwgwR4tVdWe220TB5/JMCPA8WXmfByHt/bfBs
fyyfwv6E4MrsGI65hhqZZqI80wsMTfm7loc7NR5/82WcxPjPODEuGVyAizwQ8hlgwkU8j+W/ZtKC
Xe3S7DSqmF/KtbK//oPCf1FjVBQv3rBcYe7JKmUS2mb9uQNP4gJsw0tyhpw8gvfWEqoZM4FYiav7
URU5uJKR14iqpzzj+gL45smZlrNzVCowY4ULBDW9v/mgzvc5EmWYWCVrPJLzNh+VHtIRf9/6xar/
bjACMlZuUpdGtNQqGJ3zNWwfZw+Wf0P/9WRatSrX+9XwZw8B06tkyTcrJqHzSAkUSF2G+CxhhaNL
DEOdG0nzvfqw1yv3jM6sLHNAoh6jmsd0eLRTHgr+oaH9EfeU6gosk+Z08qNLuQIpvNeo0z3qo8FV
FYLiPb002bxORyfUc5OOtOEGflVDOm1CDLgjv1fjxy406yw+9FWQS7dmTb17Sj8r8B7vCMOcgCAm
41C/JqIKjpa7N7cnWecLIxnBq6LZV6R3bdvsU5k6z3reua1H/lxcf4c1bpKnIRxg31/oWQFZTMjo
Ayrb2xmud57l9DTB83VobhBPLq4uWjxytMbc7f+J1hVvhx+d+LhZ734ocpxQediX7TRTu44XkhtL
zA+zRrSSgA5H82y77s5u+Vs/v/02b/1wCACqrKxLtJ4YgQAY+Vfu2m45hKrSyfxGYHUPZPQQgNe6
H3TDUVb6fCKttXV8ASI/5yWGe/UD/gbX+8Nf0DVVYJB09O/kPxjkFYCyrg8p5IAMQQU5kQFOCd+d
CixBVuw4WthwrWnwYR5zzGLPvXPZlGwQxXucHtAcZhaIWOzRDkbwf4HHlxaE3MK6fImGjjM39M6S
DVJCKEDsAATVGcbeNfbqvQCUA3lbskKVUH9KCqdx0ECiWa4FP76FFgce9Iok0PJ52om3Deo+vp8q
M1N3E4abTgFJmt/pXNcB5uwREYH6MNASEKD78Nd5ktd4hmHioGSqqInCsccCnGXL6O6ghuX+NOV7
riIvIuUNYCD8Pu2CV0OEw6wjKe6ts6sV0eL9jdNTSZ/UifIFDs/pnOX6ZfS5AmPZW6fMrbyMlfQj
FNmWrqVQg4YxZZAopW4La4qjjCIkZ5P1Hcq5DS7VeX9S6naun4CmyQGbhmOaU50wU34unsDblPpP
zQuHDNSZsJVLykEbSRZDlv8awaKZ+2pNevOepcXuRJpUPPB93JURB22OFE0IpaocBGxW93fFzs7T
Sg7Sj9icmBLwAIgQ+vTyUUT6ON31Tpwm8Q5Ny1lJazR8D7iaqOHlAsik6u3dzLlgqvjETBH4wHL3
CiHyBISsZ5e0iI2Z5xR3AdBV+IWP/WF6kThr7ySK7VJ/QF7211HJf/njZPA2zuc0SStpFlpSXDm+
wnf9zfuCqCdSIKBwPX6rUh6mizNTTKSiE+aehldwtmc6D8mNkKOC0AB/h0zvQp//LZNBwdneA/e0
4z8Jf+6kTlEe6bx+U7OE+OMglrUUSyzeHmt7/xhuigF4gR8Rbwt5zeAk/enOycmzetFUahTZRpcS
tIIUa8u1xJEaay3/8I9oNGRNORjM8w/q/IPttpgbACrpZAtX43ynp3bACgB0DkTZrS+E9gZgSBvV
yM/8VFVUkIMjtfhpLfCqjrBV8n9tVP2tuM9P9EHZekiicdCqPaz5v2GYrI1KTV6Yawp76MCvPfYN
SHZPadmLriyYTX9i8s40jMuK6NEzWvSXgceafwwu0A3P516ST+vgdrMFfMVsB5n5rZOIpGCJ7nLV
kf1Z4CP6r+/Jp0VKL/OCC5c+JrXWogMqLmthKDy6D2AVsKLW0DvJgFtHwn9ESUVn3Eo5R6NMC4Bz
VG2n66dy1Ds5uXK1hKOXkG5X53RPnLRunvibpQ+6nm2GFUe69FhhRZpvkzwmD8DIOArfK44YU3wM
l8W7XY9SZ5SVSKwxQEEh4IvtqjAkOuo24jrmNQ53y4LLMTINStnfMWdlUEQL/oIPVjP+tGD0F9Tn
/WejRYgm3q8HfPIehqipk3sMCc79AObKDnTR1ZldGV18yOXrYw35zaevAZEmbr21+/yM4mcu3ia6
kY5E8aw7p9pTVXM/0xxgPbmh2sZ/KtX9IkcuO3Kxo8JNnE3R5gXWxsh+HOswzd/xSJ5MnSEQNCAV
CE2xdd7yi8OY4GLR4SGWqtgMYBMeZwjWS5fTpx0FPnhVfsx/qBXOXhpMdYmZH7NLPyd+R2UE82Yq
76hg/FC9OjE3Nz4PsZZ121bizYlhD9jmwZSYeTPWubtHQnCb6xGjt2iXp8BtBWnNAlpacw5r5Y3I
GM5JjMQppGsqM8aB6DBukSUm99mZNXz8Jr41zAeQBiPgeXVYtMLB+b1P+uu0TS0dE+0JfkBKtbIw
dVhjKszwIiB8zAOzAAGdh96Dk0cVmXC/1vjzwqX1MFX9xBOs+ViJoDV0ukwZaGYGzhlPPNXX2uz4
0B3AEuhMpGR9fJD3lje5qiy+9mNm7s1E3LK01+17bqvkV7iBDa/5/jeSLhoCgtIiiuXoqpEbtfHk
eKCBcB3kOLZ85yaqfAQc+fM34f1T3qKt/FrAyd/oe7IkgokgfXjp8Fzkxd5BrA1aZOvzPGTiKjS4
vg/PRgbNW7UnIHaIJh/+FG1tCco2RWbo49fJ7btuh/6Puu2z8tQfk917IujDvB0nCu2GnySA885i
CYU1pa8Eb3NlLCs54qqp7HbvRevroznsXcK3HGd3/5GWv1K6zSQlGaJ279Ck4byIKHRSotj8mYQI
TYwL7t8wlm2y7HaHOJusqhpyjEFhACIZKkG02TfaaY+gbqHbZcxQj3VFqdzRw+xzvKZmd/hCnfXB
WZfMM1OX5zciQgwH0aIYxAai8ZcbOYIF2qHEsEEitI8DlsnMM68Xz+pFbFNL47Ula/xVas/5cJN0
peu0YrtpMtVQ7tk3X2ej80f/lZ35vCRun+E+GCCt5ywyl6GCgQzxPT7/1iaplhJ0SnsODtEkM3Cp
qBx1s/JKQIYYa8jEOyAM26GognVqtA8g6nydJLHU/5WXndIUu6Js+ImczVTpptLBurEutSUfEB7E
/tQ3ZGzzcfDLmxEAEu2nafiIAhqzxOuYEwIa8v4vsLldPDV9ziZN0Wmc/AsyVsdiw0FVElCUjXLp
MuV+IuPYb/AJ7yjtSqD98Z07MM2pJjgsA4B+wFH51COtnYQnwwyC81hN4mudEAaP8/l8YptAGEH+
MfIf7ik//L1osTaC5VmccUG/Tb4JwqFHAKwfmDtOWP9wqeyHM7OSR5vIqKuSbPjST1gsASkePzoF
TJmd/BUJ/w8mUmM5GOlY/fzIMPSlrsSAii/Dfd8YVaoOxOk9gG2g+QFHTkpq1bOQqQx7LvMVXYKc
mtKxFDlZXO52Kckoe/h8oCQJiU6RDSEOPCA9nV6WLWnFkhtuU72saIgtFXXeCptNUocmH8+n1qdY
7eVkKfjy7aCMg+jBeGle94Kju7b6eonXRZger/Xy0/H9LQtF1V38LLaaOi4RVOgOdBH9jJqh8Nam
uJvome/gumpcoECd8vAIafplH4RxR6e6s8d0qTscwPpCrNgBP5cA9hevyMWviq6LlZ1jgnaS0s6+
aJ7xKjTWSbjXa5uqQefahwE7A1JBwY2SmtPgt52AncF35f0WK/7m+L8ajl40k7g01Ebq0eSYTt84
UArbGn301WAW8hSAAjzlmr7jVBJ2caCM89HMXzdMtgIFcW4mdm1jFICJW5sdk6hBOxeN14UJbj2j
GcUO3brQ7uf6p7mGFuEYQk3pD+8Qnm1Y8lKy+zB0Ir4HwCQYETrBBxt782CQRtW/MKcHj+g1dW8t
E41XdcOlsxG/MUgRz8Q21TtfDhBkU1QWrkZdkeGQhgrndnPGbtMcaCCDh21si/p9oyUEV9oWqYt3
Uxot30WcdZw0ZIGW1L+ViMl/HfwgXevt+Y1QwbCBj3D2LPSmIZaszeEOsKswSqNrWk5/qBXGsRMG
Et38IkZtv8bVvOZXazPpAyp+ZG1XQW4/20ERrtKuAVeYiJPGnq/cKAR6sgkz8IbOBt66e9xtgc0F
YVichlFw7sT7o/5PwM7Ad6NyKTWslzFR6YwAqmFai8LDd4tMmC6zKh0lcapYzBAYBULO8bEqmv3X
/4v2wIivFuSLueobN+sYRK9mWmc4VfIv/fHrrMCe9IkUZvzeFNeXiEaUelyEtOdMmMzzEqT36Ktd
Wv05E3idqM7JbOzIUN5pNWHMCp0yvQ0S/ywcTs1s2S2K5tJsrHIqymOAM30x0Y2XxgctxE5qh2kc
DUPjt7sqPVYXxS0yCUAMHkkzPR1D3QfhR6msAqZRzZKIGfiXsbE7RDYfNL25AgjOTwI2lqTxsMBf
fiaUtwlJwRw48N+0hlKO8k3RUEHm2d/qel2wmLyEBfTzbie9Y/jwTHVqka5pism+NFZjDwWSVywl
O8C0lokIuEXdeaZw005qF/JS9p8uuHs6xlsYk0QW7KZIgpTaCd4cOz5Ok6poKJd3CUHWaqJ0wjR2
KlqG/4ADEvlTlWFfbGMvo9ReZm96VrtEomVKa37FTnoPxIa5TE8U7uSTL1HUbv/ghNO9tNvthkQH
LicQbUZyrA7N+oM8JhvduMzHLGNO3RInNwvdi0pM33NcWTQ9KhzB74Jg0QA8wuIrYgK/xEPCYBU7
bgVoz8gKEcFxJ/iyjfH4STYvfFmNWBPk4UZSVpgniyaToiHA5ZhPPJFGhlBIn+TSWt5p3tL8+5b3
RpLMBzW6af9kgIGd3OAUxJrrU0CjECNf0sLWOJpoS2ZMWvHYZrx/b5mUl4ZPYoWroei3rvqMGM1B
LtXG2ZObEFA61J2dwrhNciZQt/QLoFaEkOQtPagHIhvX1r95CPDr0mELsPumEihJDJ6Tj3ed+Ued
tp1fAY2Pl0rDZrTIo+Lv43gNwulN/RdiLSpTEvN6huN2kYRF7CqC/9KvZIekgPVKJip5D1DKc2CI
vmEaGFqmH7pF5WwGC0m6JICL4G/ufmwLCV1/KwlZfJDoD1Vyw2ZbqKE0wb1LDRFKYkfuo573QAp/
nCPck1J8kveyFCfK/vy07mJDKhsQiKDwSbcuGLaEBZYhxu4CNntmU6Mp3h7cPfL9m+cnR6j8zQ9Z
VSPhK4gMWvJOGmQWIW8fljuME0YRu4QHPE3I8qkph5PUE8tyhvDyxU6FX3o7E7lr08lzrpx8760h
iAI0eb1qQwxVJ1BARI+Qnm0ArvnaPVEbkhSHpc3kbYHGs0XOOoma6/dIdgFD/9OFBfkCYKltfObc
mvVrgrD09B6uOm1cIFTyMHk6TGlwVOFFg19+I0UhZ8bJCgK9He9GGgXJLhHbd6b24giDnS8FdOWs
9fsGR+mskHNdypDcKyERPSGj9ochD37BbRGhvC0DZPavq3wH9qUIBH86xcNyMqUeDX3Pm/nUSmKb
yEikWMZKWi7ackCMYS94VCatzYoIdVbbUcB5Zi47IFtVR2ZVDVxR8vysdWFGk6QUn28IaiyyI7yX
F6QjqTuqSaMG7R/yAdt33bggXOAkXwVHXVJ0YTlWAt15EnnsEZYYwNZ0mLB6Mu8wkd6J/22gjYNO
ycIfxQR57MZEe+fq8/DXuS3/edgGSE0TmUdtmrFGE5fzJYTXDj1WBaJGs4YO0mMm2Zdj0MGWbVOj
EYn3QF1j5h1yaOzayemiJxVv3zRJZsrCbrZf8jtq6rhSLY4ctdVQuiCg0HhRLcvnBXhSqVO5GmKm
fMiszrq65Qm/ESiIbURCndy7FXn+MpSi06G6wX8/arZAWIAsjyQ9VG4P0uulJ2WhB+5voFdHPj+h
13yHxesDCoLybBL3I8fgMUc2HFm6G2euEpGGpRdgCheOAw+8a94bzGTgV+d/eAedHXVGRvu6H3kf
qQTPmfop+e9WYp5d+/IqZWe7jY4PeVAeW4MN7kuv5VfFs8ST9RbEWK8kcfRxJ/dRT7TlfvEpnS3T
mBqGjEjEGsQ5v0/QT7y7MyLTfBc2RLf8ePB7d14YuVZttnN0Ca+pNAznsga7BUfYZEvI2yFTCGEr
LQD0nkx5Xq1BVpZL0GTardSS50B9uNLnwKkmkqRb056icBC/f5tRdrNLsUmck48Q2YMt6esgsxWo
Mwa2+OZ/+QyQ5HqItBHSsrv0EmxHC2Cb3Ihg5ETJoc2vYL3ADUVx3DjGs+Sb8oArA9tlRRU4J+Ib
c+tcHpHi4qVk8t2YiG5uHWyEF343bYiiA0BtGeUzvObKUfyTSrJtmvOzNDINhS2jzolSU5BH7z19
MG69awECoaCg+PfKe76dTscg5FMiSSHEtQHR2jpBoc8wOxNUw1BGnka/IaVcJS9TaAxJxqbH68up
6YfvKR1GJLKU1JidssmXSqXvA4H5R/iXQuqd9sKAhsO/NZbwYqp92AA2xbVHTQ0X4PUNNYAsYIaI
iVx9m2VLICG5lf/fgO6awhTWoEiD30rjBZ8nO5vgxYaiBF7nuEkIQfBsyHluVgdkuyvFGOoM2sDy
kZVPBsD/h+3ZLl/imlwbviOXYR6yAHmeUYCiq8EqkdnOTEhGUUoB1r/9fgSUBpqYPl9AZggXCAA+
+zr9dV4MaqRlwuYntQKcL3pAHf3tw+gUtdbCZS9+64betWoyu8qtfnVhjPInwqADZUKncMV8LGKB
ZZ/ANIu0ZJ9sqLTAxvq0NaXHzVkiitOHMaWSPnK0hjSEEmolQMFRmdzaIjCub3YTmR7xTV3go1Ql
4Tra23xi+WFNUIhCd2nfXI/OlvQ9M+rQdfdpeKUjIyMc6wYm/e81NyqeNjrC2zJu8TYOfJGMbXz5
fXNOqP2G1OrYBWdfKFeC/Lqs+d5beem/w4yCKj11DKNVjqHpV1AGy1Vh/NUoS7iRzsgCq0ch+3dL
Oja6r7sK0Hzz/DYWciotOJ8qEbgyc7mb5Ebakf/9x8LZdAJPuFgIA5QwOh2prGVE5fPTBWLKoDKz
nWIxIAnYJF9cN0cjFu7Ru4Xx6wpLJOXjRXrlslyxUTRrgXHg3VQK2Z1927A1Qc98qPAFN8edfe+3
HYlHONg1y4JwslAwy3Jqb/qCbktpxMN3iuEz7LU9lrd33ukAc8lVm/t2VR4pwCjIkFyLsTD8Ty/U
oHbhbcUVtGCjvtH1hIGMpFeWM70lM9+PH+Oa9vrK8xfgu1m2X8lxEMmnr4HgBHd72nO+bFtpdq/i
IL7TJFPZKwrWNU/zPIkWhwGfZ0lAgai/rKbxSeXbEQgPbaGqaSpT1d95euMiwQSLbZc2tVFwfuNh
jGuMs0jYFEdJ4b4f3v2gP0S0gUGzdua5wNUOR4XGXqS923XIR8yWCIq03mMVInvSuxpfdq7UYu16
N2bXsPn4FtGzsI6m7Srzc8NCyLaz7hTh+T6+PjFpFHolKN8Jb5I6xYkLZX0plZ2x3eC2Pm5FnJR2
DJELSKg8hIPVmc78KSvOugFkZj8v1B9vfU+TGBNUwPqK3Jt1aO+1IiibLmzTJ9XvAEhx/3tuIZdL
psPwgjHpaG8iqdCZ1cypKWfY6gDE69Wh8xk+Ap/sJxaxMnetKGyuWhG8IPkZyeC0PT0NSO1tiH0V
gyqKbKGPDUPuYbEio+06TcltS40hIzr4BLS5hYsdt5AepgwdaFnJyX4yvGWxdhXJ+a8r4x8SSBbX
g50aOt6D9iSFtbTI3EjhlQklE6Ri8aPvjAbJC/uFhqr16DyfiAb/Pn1ZrxeRZ1nTAedweLWpFNsc
rjzTfTM0WDrOtJbeDr218QvtAkBRHEQ6mH3K5iG5lKkyFzSW5SnDsd9VmS9xJHeu1b89PpaFpB0d
4QgVEbcKwBKXrzUsnFOInMqoOtXMThKX3ZdlbchipCmQ99J0/U7HLSskwCflQA42LOJrvBcaoChW
/1UR8SbOxLKIGKgtGEc9Ha1qLFW97+nCG9cRHWDrjXWHzCm/Knf6nW5zFOgSlMrB2nh6pEJr1bDl
sAQJgAGEBRNQXz9Px190gbHOS7UNjoj///DPd0YaYn++zCjqmYl6zPpngGYyudc/+oTxYpcRqV7M
0MgKaQkAA0zuVEIPhUieYzCUwo30RYb4WCWUbTe/StRJzu6MN9auqEK3IOY9TUAj57C6ffsDkPsQ
pROXBM3YaJMxctUBfd/LgyjQQxjucrpOVaxdQ896XNBOHBvYAMEVD/xNReCJF9D0tFZk2ss8YiMi
8gnb52xtM4QaIKlg23ew1zXpmYcq5C+3BdSRrgDCT9sOvGHAjVBqc28kPm5/m9SnEtPCMvCKU0GQ
8KRoBNt2aEJuZpjoskg1UT4z5Cn8M1/FG4utwb0tJ2AyPozk2jl8qQrI4waOq9vECKJjdlN5z+JU
opFbjnkCw3nQOsIf7SeMudOd9g/itfLE83xHTSjuyXZ8m/WAb9c5pEgh4e5V8SZImrLfzMP7eReq
1MgdFlymLB1Z4o4yVFaFdna7uhmnwfXFAnyg1X+AHtbbvaLc2VHH8bJiNfcenk1VImmC9sxyngw3
bFt+4hlrkbdH6oK2qyEa/NNJ/oDlhaKBQPR0PlPoeWSDoTipqKpdpCv0wKSvVFkq+8BjhaFRN+cc
2uBS/zsrIlLrF0/hIEW2W0LbS+Q6Q7e+a57+LJ+/OlVDPAcuecvqRP3i27cJTsIvzJPl4NiouU2X
m1D6pkmgKlJ0iZPZNwt5xg9oRW+tiiKQY6VGFlNMNsc25supzQiUskpid9Qyipo2A2NZIdDP+4UW
cJP9qgXoknrQUKO7e+CQR1zG2y93FAW29nk2nkE5mkdNVkE03Waa6GRPGHx52WTvRBFSVzx1atkE
ym9BLeBXGH8WMLIiyKNdS5DdngbQwc68WtNyFIGwfTNidM2NhUIJD+oZYconHcApSkY6xbN8dHfG
UvlcZrcVP5WcCEBHxEfvCQ8Vqob6KToHBnNMHHkHtpW66Ynyb1A4+krz05Nur7r3xx4CE2rjEij1
H86UwHQ4nFJsMwh+R28mYqi2wTwEBEJZQz/OHL13IhuneWS41T4wTojEv6zaDx8W/2cf87dxzRYC
QgCMV/qI8+yEpdt4qs70cUUL6kAU1PnITiLsca0UYZntbL+g9HG0fLSpuKyJACUhRhRR6HVxjls6
YXQRaj/mpjdO5noZ6OEsPqWnM+drqSbXdtSJjwGsu0WDA3wFqRBfRE/GZoRlqcGX6fGy3Ttfee/q
TtS9X3mGYl9i2QQsQjTwLl5/ZIuE4m8oQqgZ3p/kCOlJ5KQe9H2UHAl8OJmfpMXyXRuxK6wp7YO1
Z8hK4Pe4oIDZfZZUX2TyyltkXwwhH0vOQbiJSv+7wF7Y8o9z8dMCxgvYoe3F2KcRgfOo7VNlELEI
k9mCy3myoW1s9s1bCM5Vtt4CGWRPIlJKt3amaEqEnZ150u8tisn21fC/nPDbwEHee6nYjewrJBDd
ulXGlHDLpCfjcFXPi3oQ21QpgP/36bA8HvrSAA+PTjGV2pMeR8/I0sXqDIrhCKyoHfgJSEM6O7pG
E74NmFIXiRtEmXyA3+oQqQ98NW49KtgTmURZybkbpLoc8ukE2ZHuIGoOqXOCIoH5P1arUEyeqmcM
XDqYZXz4yoPNZPXnEpKBy67SnCwGzJ9F3vj5U9s5YHJoSLFiQ2sEpZg5qs0CgGGpqZzmPDHmFwkO
w5/eMt3wAw41j9jeU3S98xoE389CGVovzeidyQCObSM6DCyfoQUmzwJnv4NPKRKVokoUfBQBzI/2
OJA0kIXkutVQv0nZm/W3XBzmqLK9WxX5LF8SpYbNQQNyAon4TXkFzLkS8dKAKfotHGk9Y85zQW6u
BcBmTWaMSaIBulup8DvWm5gsCyderqbksozmg1KETAW5XEDjWqJR6hfb3ViswZWD4e8E/yrxRqoE
7NbEzqJ6QkLzr5iuvCsBc5d6xeRZQZ6Se4oTo89SkmvwuFFRoZmGkCzi8fQNA24GYTrdnJKobNCT
ZzLAqj8DCqLNqro1u3O8iRybEBPFMrqxBGBFqn5kBpQnc5ANQ0B1EhLaRJju7JBnwSyLHFekZoOX
qXbmHrbxASKz4GEvB8EyykqQp3MM/rQH54cFvvEVtNtTrYryPO68tc1xSbODdTXw7ig749azpNq+
GswSSIs7y9NTEcGUAl/skJlPq+he3BFf+XM/EdoeveQo2jg3GvDnTfmqCeAzRY/NHDwfOY/hr1ju
UlMaPrhjyqWwu16PJmHwg7LV07TvsN3Ove5zDXaVSqAqKlm/HffiUtDr6E9GsFSPdOViXNIr+9yg
9oU4Xn3XA2Lelrl25aKrxpmmqEivNE6tPWBdJCHtefOq3c0NSG+g46MVbaWKi1NNJmivzwxYvKhG
LE9KdIo6pjFvabCOI8521PDjiaKJNTxELVXkc5ivCWNxjpw1xvWxwx5tlP7NQugTt7Ft5EpY2Pko
4Cqq4Og2kYfTJIpk6iDcR2nW5qq2IuaCe/yHGog5GLqs/5x6UsFrKsWDkkk3SCJZ8PP/MYWrx2OB
NlJDLZ9AkEPUQSgsUemCFqFReVcvLg86/TcdSSVSMSAAtPuFtqSfSIKJJVbYY+KFUe1socVApJBd
cGLGjXxGomKrH0oEUFyMGgtDyGXEMmo3ri0ia9MFaRL+V7DsOKSK7XjmbOGR69zDM1xGA464yNxY
Zj23leyYXDo7deDz/tBaYONr5a+LRQKl92K/dEZC1DXpILtuKcyPLethsOMLZZUrfob6lJQfZ+Jg
/TH64vjtctFD6T+irKQQ1C9RGWJ4WnSFQSvn0e8FmvCEaCiu86sL8o/xbYLAqCwLsmswCJqHNEas
z0p8WRsWSTV/r+Qa32qDP83RG6LZFbV7fwvZPn7W1ASwxcgmMTodikizU4Wt+DWQW0gqP3d26X3i
ViVa8rpgYWKN+/aLkh3KUE1Z4Io38Dcbj7sIc1jL9NsZXZnoYspqhkzHtCC7nk4ND3GgBZbZqEjD
nDPNK/e2/GMaD4GMa28pYtIr9Hc8EQkVmzb2QCGcyoCcry4PWpVyYcQRg46Skejtj5z/rVD3MPcM
n9aMboWsrAtVFPGDwBtOrbX9VbmCfdRkQsmoP23OJklp6T5irKHgNuLzx83DlpV8tl+dCw/wfERH
0OQwPULerrTlzNOKORAqsxuAicaliblS2WfhrdWfWahoHV/1+llL/e2MNTQcPRAMW/9Xjn7U2DbP
2L1uhN66B//fm0dUGmYxvTtLi6fsha/t/gdTZCr0GL1HrQsYSg3JxCtIhQFefq8O3wsdV0Olbw9k
/2R3EiaDNubx1rj2/cIm4LeWKcHTUqStc6h3Z7s8pXPDUmZA/x19WVUvDPcH+gtoMq9WluStUNx2
0dhRlog0xL+BPMRzn6jSyAhQ6vituBNIq5JPlqc2bVdG+RaljqnsxHKbkP9mrSw/p8V0RXXGdQZ6
N+lfCAhU3SY8sludPmgGsOMHysXwYYSs3zXoziXw5Oq4maSDHex6Y0+lUfh9R9hrY6UCsqBK2rVn
My7QyQEhhEHK61rybdhIbUfdzDG0s3iGwHygf5euspnIQdUcg5508n55mrDyS9Sx48zErws2MiUt
eqzpotTtD8icMUGFayqgLTLGLL0NvFfZMbuGWBAyTu0hvEViBTGrvvv5K6gYkKrLTCmwXa4LnDqr
ejntdyIew9FitRkyeeBasuYCnqfX1SqSZW3WEQ4u9jBKqbcdDOvuYWeR/UY9E36j14k4kDuKlSRx
qYvmW1wRiXGjCYz2KLz+YdNqOk9xHejaGBU/KaAbSeYq72cuKPlcvmSVDMWIBSs5ORQuRmjuZYmR
Y9JSTKK1j1pkQaiVPUngiZa2gcD1UJBU4Vv3+j9hwAVxWVI51YiZJ/T7uyM74Z9LRaPE5qJissyq
h1dh7gxUOPhgrzzP9xDIiaWW0LHG9qN74lITFiEwtVYnGmXFmhDRnVOq6xfnGGZd6nDkZrc0IT5C
XLAd2PPtJpSEcf2yvR6p+D00ITsdTUXHpVAdNY6qfkM3nRVDK6eKBfvKpzfgxPN1heA7mOXg0pT5
4RutfjWu9W+9dzRXLwQ8K/ViwMVGiIVCgdas8UaCkG+wmdmanXkRb1KIKA+jzoSJEqdkzM5lBnRO
qziK6r8BaRmGt7mEpfGcFzWAgTFhLbpVL/xiwg3do5Ppbgt47JbGpKKnj/h8DopJkjFGqc1L+H0a
vhNKROoY5MYrcRxSDM57laM6VAkvy5frpytOehFU+pVlizDJLVT4o2H0+XoFS/F/X2TT4mS7XVEc
FIuTw1tfUbZicE9RunHXIB79xnsZpcpVW0hPYsxxmVpzaXV522CrHP80rrw/XATHXwrShR5knonv
mU77lw4ekKXps9eBlzUStuaXauy1O/gVUSidORHYSgBHSXB4ROc5+JgaoHf5Q20G9nUWdFMO6uDY
TrfVTHtkcigI8btMmb2M5rBUvS728qcH/Lt7fZ2IQ+XaQt2P7zSmZeHhQigqHYuGYNtm2JPqh/Zo
OXLLM03xh4wWJfQKtCXiIAmEf40CWcj+n9LRlsiIycMDlup93MGsa4QhSmH8Az/haV1hKDy7k7r7
+zJdYz14/oVvgRsTeak7EXJp5MWsXxYvlNp/wEFsHtVujF0/p+vZGo+E1HWtVzPdyd1s8BJtMHjf
XqXea3GlpHTndSpO8sXkQez4wNxptTSXR0RQXpmz3VfU7iLrKCWfueV3h5V6fsnya1uiduwgivoj
pWPMduMKdSuiIVLGPN1C7GnpFJztq8ZF3/G5qP40tI00EeEBkE5N71j61Xji9D/Ku1Wblk4XJ1Du
xXYALOcYSJ1+JDtyCDpoL7geZEz4qE0zYRv/vKK500HjbV4eZdjndmfvVCOD5pkVJUMdy6YBnfB5
CJ9bdanL+hObgNBwu8YIYVYdY8hVemmSdZ32S45pHH7CUffqgHCPFmNNK1585s3QXZhc3AYOYQ3n
rexELfQaz6eMTvIA6JGQEZqlW43wwSe25T/jJ0jgV6utwGcKqU2e4bzHdY8qoUs9+G4CmRTwvmX2
GwgnQUdU++GWVoKDKpqFJe8mt3qfzXbKsxL0NydNRBdsHhWWx6zog7BplrDrGtR3xSeSGIy5cH44
I9KmVuZbG2gFeMaPaBNBXWVTq2tSn/uTCF8Zwm/CQFhXq83FEy9oJWZ1b9BvRXM/V1iUr8vKqmSb
BL0nEa9Pagh907Nm+X0Gldi0QG7y7Dba8gnvZN38/HthnrqS4BLa7X/lEd4DCPC+7yy9uyPDsjZO
cIPNEpiNoNKGizA7pOWDb+3OrP4paEV2pVj4MRlvPVuT+a8gXy2yit8ZoDrqBZvq8LryUFEE6D/C
UeR9gYC0ACWcgKIHqE9O0T147vI4QdQ7UpO1GCp0yLvA6tr78cRnk3NboYT1iZrEoU5NQsOlzQDx
1okA0oE1jNR71OChM3lFpg5I1fB9CJMi50L9VS0OIIY/9hSb9kdWz535e8egsI59HMDXZJJ8iRNi
bDbKfr1Mfu/F4jVNStj0SuEuxzWGyyR9Xgkxz6ILOfke0kQTGRhnM/ZlNcYp2jDDIDz4BsjMeYhJ
6QWahaQlMKirs0qgK4WVhGwLCqsEiRaE7qX/2cbvl/Y/N7BG+jnVZ38tANydYYrDh5P0KXH6DaNm
nsyWf0up2BiM4ikxD3YLmIJ/8mNskznBqAz987IgqIHzthuIhS7wnTjcfzPq3Hjz6VL1UxjgotMI
WZaafsvSLscnyXnRQM+KZxI6EmMPpb0hd3WWDLJmbiyh0Qc2MMHXYS5qMUE117zVe7Bu4MvkTZzE
w7AF51W1nhnuWy93xTHirIoLLYAUcx7Ho5mEo/AEp/zd8v6kVd/EQuen3lWdl4qJqD5UulZrPAAi
8gvZsg6HTpfDb+Gls9AiHaUw27xLJxwXTDQ3zw47zvLdjFvVdZ9unUJlYi4mouuCOCTi/+XeolRd
ETG0f5aDhT/CVvOfi9UpXDyzbUdfbwJt13zu6kesyzKjQdZOQECLqsht/At0gUZXBWwmahCzssg9
5tCMaw75O597o7/YT8AavQtiNR5cqPN7nNXVkOHYBsBuaojfg9B8lp7//x+4s0XiuuCo0upu2Pzc
Zvt0hYpUGXe+S+C4O4h9TI7YkZfHlsaJBT4vqjFKjnvKEOw7010r3Lefd5CISyup5ZwFPqMffkAu
+7oa9ih0GpNJvpA5Z37DhnwzsFc9miA47nF6KtClmGY3ZtGROYEJDSCqTx2QuKdvVZK9/P47Zs2a
nPF1IwPh385pHCadcEPPZeTGbQyZBUBk+Po2TgoBkIzA6/dr87EO4R80++s/pr5Z4/koIXQ92WlK
HtDZlC/aG7Jhh7o2Odphl/1nar1LOo7eZnX2XK7k2QmpJXXDPpImbzmgC84DI5Vs4SVkkJoWHS9R
HWmVlIoL7Kp3CivfEIgqvWAhjvPEE+OymP6Dn2yW4w4yUZgWt/wdIFFQUE8GJ6Zv2K+EPhfNG7nd
xQbD+5eWVZamy+nWA7rE7DKxX7dVxZxh9+GUviSn8xTnjzy7dErx4g5M6PN77TAn0E5jzvXmW97U
++l8dd6CWYB3sUHpec3a+6JGUPaU84k6XmIsDK+bpmVJUjeUiWCoJSx8rEj4s/hpyOuOE31+QQsu
fQtr2zHuI3f7MDKKj45Dl2/D8AOQLmAG7xHDIUKOLNXGqSN5usF5bx0NX0eVj+cRng/VZiHH0Cxc
sKCARXgnZRtWwuuw8eU1fH/mCBC0ZM2+LAAY5ubjH/xfFXrT5QVTnv81LU8XqQvpEfPhr1zgrUNm
PLNirOlem3VgccPcEC/2jyUdHPYcX4jjIki68/wWdZqwLhUWqWklxSeIvFxoyvQmI1vpYYJclw2P
DKSe7NujV74ueWfHg105qo5NzRMOUEw4GdNcceh7g27y5NcCBkrl5HhqXTn9q9Zt/0pMgh5ems4m
wcxLXM48CVf2OPaKWxEHI4GQM5Xmq8aLL9J/g1F/n++iPcm4xidokg4XQYF9sE3LU+GU5oIxt8Pg
ZIQS+yaHKoUg5agDuP9+V1urUzUDuDp455onjABokksO2NFD36MxWfhNgi1pSS52UzhUbtiqb0cH
vVKZGxCYrj4PFj5/MlxpTJtr41sew7x2tXO+Pvswcw3BK+oY+J0gbvs9yZtPgRcevD243/C3Z6bQ
3RMiFa3V0uH2VyHBUGI/bYqwb0qtir1j6y3tkVvV0sok2zPqqVPpObwmq4oApMBkxdAo6Vz/Vv9p
bFuRBjpikU5xJAuJlUAo1e5pfy2YAQby0WfkEHwFIL75Xoik7LSrQCPBUHFEmjwZMzJSZYvpMJcz
XFVioq7qF1nlXqJePf491bQWpVNQeJjIyE1LHsWZ7VdyWc1tyAmj/7mXfLcmMjcn3QqE2/E/+LGH
2U85qGWY+c5Iut3L2HH72twgySvL8i0TtCoDtM33KIY6hKixc4v5Py36LKpnUAaveP8SMVIgw++N
3sbs+0+p0Jm5f5aFjO3shtlqgscK2uAgwRnlBTQtrd8kCLX4v7FcNbVZk1kUawVBigiQJer7H8nx
JKoU2wfEVy/CQ3cxuMFtGba3y+Z9trLc5wl38vrTb4MwldALZQKkULhZB98OhgKGeeYOX7SToTEc
pgzzKFKYwB8n7acwKhMZzKbyRXtnxHZd+691+SvmesVpw8y5TsQPe/677xv5FJlNW8i57abVXuLz
EzHTsRwNfWA9fzUblBXSNvm5b1Q3c4IA5QJ9YjidYxgX5ZkpUZ1frmNdta84mN3eLmd15rJ7ATaD
ikzvriXhALnLwqUEGim8K5kZ56b4Uv3hN4KF3ZUZVZuBpgeK8PSqFHC9O881wNTplE//oHRo6QmY
SLlZBUfDvm+CxEYUIlSgDS2S38DprbMDGSkUDROO8thKFXO7WKHL6pEYK7H3zUnET+W5RqqNMTGE
GHnY66qiQqHlqWAaEfN/wf4pXCZ2L1oKT2VFSrOKHXdBinp0nZ8I/wMwd4Zyaag9uWwrlfpEtKQd
pvqzKwXIJEQ0NApfqQZfy7PY9mTYqc0JnvujeDrxrecc1YMkQmuuWZq0SBcPEV7tQJA7XSxnorzl
VskPD5vaZD3faCubG7s+NNYxJ5VLoPy7gwUkj9NXYqLz4PKWR8E1KEFeEJFpYfUG+BSkLb0Nlhvp
Gqs8ja+k9TDrhpt3l5HkG98RDJt0nXo6IIcusRMhqctauLIMH/pcjxavZH2I/Qiw7Ei35RslgqF+
bivJsOYLiuMNLM+sV3OnqyCex/rw8Oe1v/fOznTVF2Dx9TMtO1ZEascDNX//9krcyUlba4Tyonnt
xzZcwKImgh8pmZb4/1en8UzNgOTWLIPMIF8IqYg1f0SO+3E/RhlAHan+9Wr1Jrs2uMzQpdmOsfyB
PA30WmcCfcqnR7/J12NjfNjjxUtYCXvfRT2nwx37o3/r4q3g0638IzyA62nHlBcFdzLkR61GgW5y
gspCjsjQO52TeXlihAIoaXAHIQtE/HftSUkI4abn0NQgTOI60F0s+dS1nrQygI9Phhfh0cW6sXdB
Hf3bd9uNkgZvo5iM/8NuMlR2mzIqIRZaMrKOAsBa3zPBBiJkNVZn/t3LFiH8eT8edIDgXeYOGd4O
vNRI1GDGw1ZyVqrTsnzYcFIds0iE4LBKkk/UJ0o4W7YRouwB2+T8ZR5r4j3of0DKhItvnu4wOmwO
wEVL17c7r4JeXNg6YP9Lv93buNH3q+isfH2gPrsYddpFyAozPE/ze5IFa3WbNgdE0WJsIdXKOqjQ
z8lNp/hVOR3x8IgCTJyN4b7G53U5eq3NAI/e6VP7Pta8Y9a/m87WO/BY9hcotM9C5Uma2ushlG1B
StRzdgfRtPz5nEbc/9aiHeOoUylnAyDqIJGfb+WeidAz3Rv/iS+l/5NIJ0/8WOrEaeKUu8n0Ed/r
37T7LN5zWhGWH3cWsjZQC/broPNRj00dJw8DX3RRkszh7yISxoOhpr78JTYR3pge8PRHkb+d1605
0oOgljg3WNZRdjD4TFFu35Jz6j9RGPxdt5OhRFnZvK6g044zz+ynjPdkoCi/XRodxjX5q/wxc10k
Uzxc/J3mB8pOG1UOCxGhy9IACrZbaiJNAtiIt34Ct0YdfeKwUVDpme2E0UYwDJ60v/gIH5yrxvuL
1/fHD7j60QtO1BiVU9gIyWPwD1+g41CNieH8WCkYUslq8IM2KTxhlVv/ybArzR+Ib/shzuOhzc+/
+4POnV3rViZ1mH986riGJwTHBqDERAmP/r23cLMWD0wK14DRDw1BEOmOJq/X8KTGdzk5hOk5P4em
gLCE4rJ7LTOTJMe4DhqWVYyAWgEPG1L/+TzQ1nISgkL5CEL6K8T72YScWI+4nQPQ/fEzBvHGWgyc
ur9S0qhmyKASJrI25v0NoE9SPHu/jcn1/oVedUgHpEqTCn1FpTWkdOChT7mJ7hYFtonyodSmdjaE
/lu7gyuVoP8VMKv4C6H0GjDzxvXYoNdbdDbQWMp9p+06zaeSs+UGe3qhL7CSl+jPFIzvDhu3Dj5E
jD2rwsl7ndQis5K4tfi1JxvFg36mdZ/J0UlIFjHWz77R3TczHOfn0ygg2OFx56tlO71yngl9X7Rl
wKn+g2abHXqRP/GWwEYw1JA4/w2dHHlcIG2ZZzov+n/SGmD3JD4urubgkXbP/Fh1yIx3lubwW0YT
FNrbMMRi+RC0PBmCpcvo9aLbzeW0na+/cr4SQnIDWmabLkp+bABr+V5SgCi1PqifSqBrsiz6iZIG
O0loD9qzWEN0fi1QnCJaUQNRPebIlun3Wn+8bnBcPXIuq0uZkHoinxjE6NMg6Swh8UaxXEEzJF17
dva/53v4Z5dg/5GfsLu+dNARSzI27guP15GyIsk0+ai/6cGjdLoGyMhiPIqO/+VPefJJetbRcJhJ
XE4cfI7rip+9+DN3TqmpQVjcOmGH65dsnSoMy50ZM91akGX5MSSCrNTsVPBLkab29HeFdB8nRLsN
pVcUz9FfHf6ZM3Tgp+LxLRu/AJayxvKQDJECSQ141ESkJtOGsIqA1dF+fc3Na4wygZ0Ravr/zH+o
b6EW/X3Aj5yPn49vcMdsH+pplA93gSp0HJnSZdld+8nMklhYaOYuxyWKnnR8GIG/mtZPxnAwKN6n
E8488692T7zDlZ0UjCSLIufVue3gkOvLkpUpV8Nsrx2vkgpbh7gkhtH4TIOisrkKYx9gBpQ0pFg=
`protect end_protected
