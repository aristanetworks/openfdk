--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
aZJEvX6rdd3I1DZFb8fu40S8kKH/3j5aCqQldR7Kn64Q0mVKY9pYhgpS/5GSbqx5yQSKXCFsDH1j
Wx/h/OaiKXiz2qVNrSZLG5DajHiV5VVRmGsCkAw7R/vCzsCrmNvEhJjz5qUzHdF7NYke/m+ozQxz
DK5GyUsJ1zUCPbrndZ3psZg1BwVtw/9PTPDTdqr8zAl0fHwWwC80SBfwTW/IqHx9Isb0Fw20lOtF
h//R3jMYuJ0TBvH4ZxrRh+k9Z7bfeR4Y/zKzIFs7l+ufGm6MtMZ0zH+1iRcQWL7/yIerPCjZrmrA
C248C26r1uCScnZutXTCHfLiTYQC0CL4cUsafQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="mX61BCqrnvZSlUB2sI1Bo9mkE98S+XCFTZ/5eTblo9s="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
kBQXkiMpShARLo/MvN4LX0W1h3g+dACoC2q7NY3PM9EYUPb8rJ+WUDZb1IwbNJT17HHjt6KCIukW
MUR7ISf3Fs9va1e7jKaiJ5VNlbcN3esQS7LR2aWUs/gYIPDicA2SIlLdqY4ECRcHyVAgPLk41ytN
luxMHnYEGqTkmsH8ataSUcGYdTDZz4Uemakoe67myalaIj/Nh+r58whS2VpJwBcd6SBZAObncM04
lYo/+mnbFfk9Klw+9YCAIAbaiGV73GFtLxFSVP02NPaguyhtiWWg9Lef+d/8ZKKVGlM2idnTQ0r8
TPrSoVjoUuuYQiNsaxhlWBW9y3wmpd9Cn4vfsg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="AMmjQjiWMZRYWG+D9/AxfZZ1yrGg1l6FP6Owijrrhh4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10576)
`protect data_block
pmXDRn71yuvEX42mR9xUmkCzTbHAcsMFMACmn6NKhDYWzRKrvfxyWK6Eou83Z1ALFbY2ZmlVDqzN
K6ZpTSNTPAQrdop8lrVN8wYCjm4yD67vgcOR0u4rZvsu/EruLqejmHRLzBMSBm+hIyRZmDvyWCMR
pYGNHGjbjVgKiSNyU+HpPtbq/4QF0nSXPKe6QkuAIrhYpFJ5hzke2vkG9NwIim9m1Z1rOIm4+ptt
mOFxNN7r5m0qVx4JryuI8v35j/yzUhRMqAxghFELbYfJo2bD5wG33wNuGWRRheD7vrO4WKIaLKAn
XOuqg5On+rorfULY5mupXIZQ1cvge40klT8KWLfacSP/KI1P06NG2O4vdS7d6KjVRi/40DwmXjoQ
mOpXXsRX8XO2nDUX4WXkUT3TmU/8WJsRbzH8zGcs0XEDBCsMecZNSKBmXr5ORv/C44ZCX9EFlY3H
mHXOc6DvyW1WVABZIKsWkWxT0jU45VHJwYp9aQdu7uBHWcFFd8PiiV5hvp18m43eZYWc7fFZ+7Lb
uIoyMchIZ0HZ3rRi+a5BLP9h+OkaXXALd/hq/1e8rXelLOQp+Eo2f73T35KWWKPFRbFNz71QeODN
mkCtY5meKC1NMPg9c/ln4VXTCjwEcHlW2TVpr+wjlYhMWsfscq8Pj4aet7cZplnnMNJi6atSI+ns
6MhKBM/8B4V9Z5O9Ryraugzp3UeZFhmEbsqRPu1+4IS7wBe2Ir2EorU8B7dXPo/u7F8ulIjrK6ao
X+lAiBXGCBryO11gY6IxFAr8uqG4AJPtATFoF2GA0E/lE6xawlz6cx5ZWlfa0k/IKBwXjyy633pv
1UQ7YJ6MaGzKCR7AimkrDVdQ/c/PV67ylM4w6qbBasc0QvxmUGbMg59yGZZ2hCbtAYz8IxXZVPbA
JWZBGwZQ0TIJXHQKopT+3MBxK7stJNqZu0GPWnsMuQV31X7hXch1Wq1OVx7x741eOy4x4l9xq2bD
L5m5AWSs0+tNEAjadz5si+7ICABaIPUL5D0smKB0gblQLVzWQscsMCifovnUKB2/eYG553zFhafC
uFalbL87wxO5xQ/CA6Wv8H7/oAYRMJonbbBB3/3kxb6dKb/sclLkb9TQOIRZaGS+MZtZE18Ulz99
j25MOIxJgYJIMqCyd/X1tDOvU4P5urdsl5Q+n0rFJfDu7u2LXznah41UyBFtM+nIrQFRzz1RanYg
Zz/CKYKHe/LtdzW4Z2VsipAE5Sj8+4bM59Qu8K1Y1qWK6Ne2zXqpMyEN1HcF+dVws9AsauaogIQE
6VMNGeyflzwoumA/OIvXdq4mKjrvQ0tNi9q8XjtKuwN1LdtGkoLnUXukKwf6p+a4z0gAyuECnZkD
6wOuzcx+rzr6dEtUrozzm72HiDKzIg0aLJtfwREHiPnTX3UVLMYceffH/zOWKtWWr1cYNlTlTEtP
cWizQ5Md7x3vH6qJJbKiYZf5if4+jVZzllHIULAcB3D/9bGY5EY++aOSR6Z/XYVtN6qnf+rrQhvF
bZ7YR/vIVLgW+ZjJZPZKG6Yqk/xuK7l+88Kz60Bq1burTj3hlipFAroWg/HEpmLFRjNDFhoBJ6EV
DAD10A6Rv+T378dLr5giBscV2Ee7+SLuZceBkID/83uhfMI/ckeFEPOr6I+2u/1cWS3wM3FNEhzo
uqLB8QIO/sH3mBrT/9m7iynyP4sp/ddnqoyj7PbGeqrRHn/nzChT5DP0Ji8xxx+74HlFS0vW7onH
KkVhbKPSVCnUuGxC0gzeWgI2YFidnpMw+55Ng5NLCwk+OaWN7pYfBapLaxHvE+GqM+5QRl8t/Y6z
gAw5d5aKFRqUu1Kk+vg+JuRZu3B5+WZYMwMfBHwO+WewMPrvkCycVagoBecE16YE9xlwtJfudoeY
Kxym7Q3bSxtJUUzzx1Kwo7qQqhTiOrCTgS6Bos32X2gaZLlrD8hP+K4ZO+pMrEgiaowm1Tlhni5+
Ji8GLpw6U+L3JrMRD0iXRDjtwhCOuNQ6Jp2pVTub/z0jpyCbeacipKlkROlUK0YPMK32sNo1BtEk
8ItuHjszu8JztBJfBEEIWwEniVI95TlDpIZaLWHypJXlOs7jqg2qv/r8jdI4Q+6y24Ecu0ntdjO+
+XIak7X6sAhWJWesromR6lHSkuQJt8XN4wjMRxBIBxeehb6nAhytOOXzfXGLao9h4Scq3I5D9fFw
Biq6EpPrmg1iIS5TsGFKpPFS5U4e+kvDviZf2YXsjHQ7VJvB0AM5iL4ojga6DwugMTRL3rWEp/Jb
9ICjdOp8PJwEyw2WZreE7oaDc4WjY/RxGv1rCz+IMOMooR/VTPU+e9HI8G/Cc/xtM4AejGLb0zVJ
+lQTUV3rBVzB6H1NmxZDmPWA5CHuGqZxTpBajjUFzQ5V41sg/yOOKCAo1t+NpUx2tpYSsqkR6XRE
ItYfVu9vqvqogk+yZO0ppWxfCLv102OfgGGvEwGHZ8t1UIMVHGflJLHeFsZDIZeIYuoe71cTshQN
aONgEwBkDURiLkhlTABX3sh1SnF9HTHvzUZnvAkz/ueZS5a1LcQ5l24lTkkynfc/Uafb0BxQZsMG
bbF7pkc6sJ5nfY8DzLWQ8AxzEncOo+1mg4PxtGbCrwPfhHChSNC7vfJLNcE5KN8cnz1rATXExOIO
+Ayk3WVIMX2lcntjIL+pZaCoCZrvvhouvK3buHat+uxL3spRaPTde0YBYimlSbRo14jOM+6SS3oy
QfmTgJra+OI92qWpZSKRG2Z4vJV5LK3Uhf7/ePJ4Nz/t0WAnkH7BXt0LX2SImFwrpoe9n2EeGBGO
FudTHaVe299iMxVlvC3rjenYuuT8kgqcnGg4U6QAfSzhZqmVDZ35lxhnPzfeUoG0UhENcXyn8Pj5
9+S6oGnIbD1vRZx3bi0FCbghoKaXos9ZOU5mPlKRWYgyXkFeixywlBVAkLrQe4hKW7rs5nC7jkT0
Ahk+jMxFIalqUxGGSgMMryExMT0yQqyzuPuHsS4e/x+ZSlLtHm5bydhPIDIcGETrvVRWdOnceqoQ
IZkWutYweFMR2bSyOD0tsAc7/UcVhmNk+wXr/XfVJAtEa4I6A02ZDJwp6a+MfimQ7Kq3MgJhZpDz
4eIJ5r1UR7FpQkhDecGtQ0NmQ/CvneT4eD8DhFADawQQUou+GY6gSbU37AdXOcNrsrK7YxcigJx8
05ud1ffFfFr4QLzg5SOf3H5u0rcFenlxxi4a9dB3ICu37SreRWeJQKUaChD3zPIAHTFwzUzNSfI/
qOIj+PirslO+Y1EptGrTUWgMq9JOuxkhK+gUzacArVYbCGZONbXRrsMu8ajCYjdhEYCO/NE5eVLX
G9nkZhZDZrVkGN3ABf24bV8sIb5gd4MTYeFqCzGqNpm0pRrwvQSwRnLNQfNy0nyObyAYGWztinxW
ntPUkK6UmHQ55k4+GBk98jkrQHf1fcyFU4vZX8lpq20UedINSVxN/UxuICx1k5ZfL8171kl6K1uM
NQ1nQhZREcNQFgHAb0W1q6M7bWTgb7zfafJcHXYvmW/mrcRxI3XJeDylPVqhVHv3XFYUBGk1q+86
nkrEpeaohnnZeEAtUel2wDIsQLg03Lep/yYu3GRfa5soE4i7zKDtkivxR0qmwHMujtQKhgE9Evg1
5OEQpwpPkq0IlLmLx8rPkcTNiBJwoBsC5Blf8Cwd8MbxuFdze9tBHDXs+D1SQkEAUQ6qXC/ZLPAa
hOZ+j1FcGcDTO9cHR+MPMlZ8Tl/3Ful1HcQtdd3pT1I1CP9szoN05Hlo714/fJRJ+Q6jurotSv4h
ug/3uv/M95mKvvYv6DiqzyReaEmOYAP0vd7xRKgCIYy3C4DhG0Qt2UYlTcapxfnmtstrT4nAryVt
UfQ3qYZ6o0awrP7bHwxDpeKt09uW0NgZOh23/fX5BKJ/f19DaOgD6YPyfBjiCBWg5vikC9Gy9o1R
qBvTj/bP9vkK0CwpIWvvkoe8Kb2l/qTLNxrsnoDwbSlUk1oow6oHc3q4/mF3E8hFb959alvI9Qti
uls6E710eAYHIHRTmV+3KTZPYTLq3DhW/CrbEs6+q4to8nAC2pQLCMoMiesvgdAMP9k3R7aYKd8D
0eI3gyt6o5mLuEkw/EhF2x13R36gs2fhubakv3Z918x31GhMB/KUXQkWbGAQA79LdnDNZHZtwi5k
++O1fgJAFU59Iz/r6QNgKzXXGPgr1Ayxj9GdnNfRy9bfjJgb+W+iokQZ0fa9HKS8JUwDC0na3SJx
n7IJPwiCSmVRpVq9Pkb2p7uB4qR5Froqo2x1jZRTYgHg0QF41MF2+RR4AXfEwrkhBgYKq8txi+pM
76d3ZYm5tiRrt3p+XY1RF1kylkZpVOQtzeMK4nNjA7QNNFbfcZOAmvMfFh1ju8sJZSWFxcOEbCef
XGkWm/37v1xAfVWfdgedxnMhsuvDy/fMrNzhTANeYwebSYAvBKs+s6dLnNJ7cpdJco2d6RXN+oPy
4Y+yZEMQHEFBx2VRTMZhBMLWIu/v2tkm+vdXwgr3SHgxSdyVb6Az22uC/PLQo8Z6Qkwi32K5lKYR
Ddkzw9sKC1KedjA8pAW8p09QnCfS0MWNRSY+R0v0i7FRejwvSC13TzxPORY/1FMtlmqOX0v3k8YT
ZBsHpp7FaKaiF78igJSnOmckAauFBzoxqkj/+SSl1ZAEUfxp8hkkmAC1Zr3nRpqSc6shjIsjmtLN
PCe9gqkFi0AfX2sgnPAXDZGMJCsZ0DhGSJkOPX6sucSvERG+QC1cyydl2iOZTAqY1Zx3B7KT9d1p
J4aR2KLgh2KjjBTMKsKCpe7kuOKe4ndqJIiXXJlbZRFrVWMDRf/FaAnGXnfUipeFCwRV5rzGAOyp
uwHCl8jkt6gzKybfEJQ5159SHLc5asI9QixKojnSugmoVBNzgRa5pZKCr1ZsIDumTwL6SZrPV96p
vMU1m5cpA5YG0t8qZvCngEqSTeF71LxBLO+K9tzQh8SBH3gJhSgCcK7dyDgi/camL7FkVoBcF08G
5Mk+pYSZJ7NnP2q0FELTeVgCI4q1F55TJ7tFQWqKrs/nEVgs78x1QpmEymmlpEH1cvkdOx0TaJ+S
fkiv77a36tjWJyLYWBaECeyyGOux8tyoGdo67YnnAXl1HZvDQnhm1PWxH+F+DWmb0EwpASGKphzD
Fjk+LBVi9I/gwpJbK739sLlE9X/q1V1sIswh1Nqrci3LLeoZQTMDWCHz03PQPkzFBtEP3gv/IlhI
ENcIWOBvNqlVxu9xml0TJWC+aBwd8OpDEr32/9v6z53OSvC+lZdknELLKoTRH8uVibng3y+pHVrO
PaDCgJCc73OFPkNl6m6W18kKIVAps1JhxNLcosDiu1+mkDoYq1WEvGRPEik0GJM9yAUGVDMUDHT1
N3yVWAzb3ZTpN57eP0HtllFkDYOBVqXCgVZ/+Ri6su9dIwPqy14UdI9gTgwgdJvdnJbcz5hx33zC
1zcqjyUTDOTqIPA6hmdYXiirqTqPFNOwUwXgaPx1U3K1lQxf3oPUhbEokS3Fy+cUwjQfDY2Vgt7i
DVELeLfoiFZ+S4Kv7kTlGnDvP7qvBTqHPi6fVd+hhZWlzVmVBj8NJ1t+AM8Mdi2QPInefY3uQz1L
yl9e3p7FNWbH3BZZykIBPMs9C630h5JnPtMDNpFCQJ7eCcPxXe7HZInZeSy0DmFdO+v1Ku7JOhbU
A5dt5BYuubnPyszi4EKO0FShLFzJOqoKDnqtvZbTH0NQEZc2XSe4AIk87M2TGI1qykZPOcYNsrfL
K5E/d+dYBO4d8FdpGNp6QuSyRF5m6s17aOOBb1NmVSRn5w0H0GjVoNTGVIBYZXEIcWhFKE5dd/Vr
e4dK2WHRAfqyingI7s3Sp3TyDXFukS3Hc75UyKGUOxnb2IQw9YNenyhzJPzZo23roSFQXUz66+cR
WEYZkCgkzXXEPfqdVOGc4RaB/UNu2unvN1M4ZgdqPs3gtWqpBpDd8F/jNiWvJOF+UXfrnVr2ZgoV
gf0PffEgTWJAKgx8CVALUEM4U6JW8C5WxOdbXycfuqXC5O/7sq47KiP3Egaar0eI8I7miPc8Z/Ng
U7hciIpy5eq1wbBh484tiL9m2FUNIXGWcyJGV0RZjHLTfK+dlj577f5ycmT505r/WwcpGl5nY0p3
FCNrPjI61jLkvB/o6eIXLryxh1GSQT0wuIWGTqNCTLJEHTc0U4kft8ymjBNNChZ41pf/UClFgk2w
0LX8WwrjlwvF4wumvL7DQYrioNg1Y1M8IV7Gxn07qXd0In+oB/yUPQ4zytxhw4hlTz5OQHRDMfC/
gh9HE+38dDMUkzE+bMYXbDQFvITjGwz2Lx9vdJpjFpx4IZUtgnY4YNFZ8gYXKNYql+n8PGfUHqzi
62WpNZDyMqKU0Ff9m93qhGL5WlwZfOTdB08GhMB62NYYmtWgAbP/9wyFWfMLWaBXr/yXgb+/9iV4
v4o4mjvP0L3uBP6kK9PabZmKQgKipC8BmJC/P8CmbZt7P723ZnCda6wplKj+w4w+jZZ2SIWuWeBd
Qk5a3o0NbRuEf08hJOu3rcJZNXLHGoj7ikK1AQjsHnbdIRGE9Mm6ucXPYWz43b0LNie2eG3aNvGR
M5OTEYtyZtzOr8bxeNjp1nSCmq3usFvvKiYbmuuBk6YGFwHY9lwFCbHvvugtmc1KlC1ppBONoh5w
TsiSwEoddV9iq5EwI3OPDP8Olk2gjpJR9se5wlPBKsO6yTWvvvGtkG1ifmaBUgNkMrOHiTcTpOJi
iO6yIqdnSADHbZVXdOlfh2ENIv+7SkqlFt9x6Fdb0+m303gst90h8axtylmOXrnoTIIRNKhy10Oj
0Up+ZEkHnf/MnOdOwotVBXgyXvhTNAD6D/ECPHn8EEWjZ/Hgq/PbFsiXF/EhxN27dfp3Dv/oIL+Y
S60za1EMdabbQa3qhDXeuAqjkVg8O/f9PJOttOrziWBYdui8z+jyoeJ0f77vTczw+eqKsTw/aCVD
6NmUNsZ1Fxjfe+1CnDsoN2qXS9kR+M6QtwKPDZeK7TKM+Sjgc5caPedWF6SDWEwJtIlM5dlaanMq
klt28vuxCKADeXGTEPVnKGFrFvcaE/pybPKBSkiprWZOw0X5ASdkYtqvVyRLTQtiyLZklSbjcMr4
4JlEgiVF8bMCFIrYih5hjCk/9I0+rJuaMISmsnFxyS4zuZXq8A4/nV8CQ7M2cPJgPtM0tpo4wSd+
dwr1+5OBUj04R1c2jPVShNOwJFkkqGwFKHsFYfYlWUyhSeRwpAxIX5WY2fVhBPd+8JRGH9LRYAgP
5gCCY8Q0sdVaILUDflisgC6s006+I1TmTAt89aDDmoBK2+0AV0tdQBPwdG0zjEgWn/8sRep6cXS+
I2rUZ40s95vg/XTyi67FyrFLKw8oho5kAfAbgvFvsCWXVK7vE00MnsdcSbEGy82wS+yov6Sfu8e9
o7pNEEMTNQY7xsf8byafAyQ4fMYRoN0okcRQt/UvNuxWqpgO1fIhmVSay4olFnmoxo2UbL6VmxDa
yCfmH3GSE6RLPcKiYiz/XYBkbqsBAGtX9hXBCrcg9VpUBx4jw32vwEo9fNeVEH4/SgWFWqn6ktGx
7ilXE4wr3gbkWWgnc1zGjhkM7UqCwxHEFX/1GahEyRYi/pk3Lwt0w2IJ/zpKQvLJgeV5wYyGsszR
RC5tH9x0vfwlZp24EDefJimd4oJ1ddI5chNIsi1IM9Ce0pLSPrNvBO0FK00UHa7OilEmLNziY7vV
bxZvtLplmgR80Pqg1Tua5h5Cap8NNxE+USk0Pq7z13Dp4wzAFhBh46Uj25ZNqfTRa/gnDzi6XJ27
xjESqB/nxAdPSBopYEDbGtyvaqr1xk44z2E4uBMWul58UDvfVwqntELb1fwUBouwm5xkgHGbN0tV
Anr5E7AgjmzCPVtSRyZfgWEj+J+jwVOaItovyes8Euj8tMgSxEH+gtx+wXbT9452A9cZM7kDCS/X
SPYrz8jDQ/9YrK7I90uiJMPI335V7SecLQSrKE1W2xSJ52hjz7gs/7pQUdDviV5GIQOFgy0QYUyB
xy42TGM425XheSsuM6a+kvaDmvHYud7m0E21CStyR5lGivnBJFl5sosZS9jIJvNzkoQ2IUtYtfDH
n7f43pE0ggwvxs/MCPe7LOvja7XPLxV/0fpFMthNw/2LfuYRjxQb5GSkxQ1m7qOmSyHiIcoQZHaR
nFP5Rea5I9QCzFWXRlm1OTs87MJOtJGwySBgHi6qAwsrAkrX7JtC55BE4kh+FD8v8J6kOVpsPEh1
4abdHEnt/z9GNL62fgyjAB/Yq7sZkpDlQaZ9FhoAd4Rxq3Qlpby9fQm9ZjV4Nw/xO5lYCaT5yHLX
miSzHffESTRxbpZ93eisVI245L0o4CJgjMjcSY4lsBtp4TiZ72BecGaaS/WKyOtSo6og/SScSLYc
aTXBepf+xXEzWcOAJsfY3EOErlIdI6ANnJEvK/q/9giW5Keh1qkFHVjqNEVwxJXmd+WK4FCqnLUK
fKjhcVD1YSolZGJO5Kuib7d4tPJoBSoRBN6KMGlCpc4wEJQrjedq1VugsQlTTcdhR1U1/S0SZNmA
y/X1TmiFVK7bOlwKBHk36OZPlW7Q0Pkpmfi+Lo7TOOyncZ859rH5de+ZN/Q5LIv9vPWSds0DFBUl
dAWJEcE0W+dMUJVUyKah38RoBm2yqtDosEWn9vTnTusj1nc3vIFUAUMGEGRFNqbg87pe+Ly5/dXx
XFyvvW2VY22RLhe66ila/ke+4nqqHTW0vRCPwZ7pvfD95d86kuHu+pae15rKCvBatab3bvd14aZQ
WumM435DiCv/IrKQv7z5qoTpxUwfBNsNSx056wS+wgFGnFyTrD+txrayK7JbrEbLmEISuu6ex582
WfFTE1PzpkfWyGjGRxmnMycdvB0dhd9tNHwdRKhz0lRTio30yxnOKjlZfVyyIrhs3vgQtBXCnBwS
XKa5yNEq1aBQYg3N+cd97CBIZo/wGieoKhpLn/xjgquvlg2xnsCCoShO8JJxWHg1VcuRLmmr1Cn7
/6uHDehn/Jsm82fRT1Rbz4DfGmxwPt62hJRZcJmYjQR0gpPD6Lr78B6K0WorckNM3pkW5NxEwscB
25UGYYubkV83pdhm1whlFNFyJNs055KrqkdG5af351U0SB73gweFsH+Eow1nNqyoSg9K2xeNBGv7
3WLhCoo3URg3uuQxP1ByCMaFQKN/t8rAG28j1B5GoMgIY8z6nmT2DhaFs0y5I7qwqv8rxCbvfYbO
a3VFjDvVbFjAalQ9iEq61elEV4mj4iYgVmK0w7xLzEyqax0IGMPGgV0Non8LIk8DIjUaxg2RCxWv
b67F6VoWFJXoZ2Rns6JUolxiet8YoJSL+LVt6sAf8OdllVbgjEHlE8GVPTZTHwrNjAI4zPVU8ekp
9G4QonnZJSWipnGkUR0dYpL3c64SvSOOGR5Om4W1LcTPNNyOs19xVPlzOBM2un7bDPJ8BmNgfs2d
GYBDezmpRHNeGtEvRE7EKIW4a6QnJs6j/l1bLE6AK/v/56aCQPWX8S4MrA28KkZQk5kA/skdyiYF
l8vWkoAEaQeaP91P7yxdzj1VBgIx7zh9ztCZ9GHYOb0xBbevW6sywFa3KwEGigX/EDEgtjq7KCjQ
HusD3776rpOT2689/wX0p3+GM0pCIk7TzAK+y1Ra9pS9svd9bhaGDrQ/6CflINq3FdZUV35+R4QL
NMfk8Z5wiZnz5Y6LLrLBB7MTBuzyLs06HOYNpCCLrNeWWfGzUFxB40qoj+MuO3ywxXHyMi1Q+SPg
0aSAfT04YUyKH35+sTxXQStoVQieB4iuaQAkG4La695Vu2eP43EDtbfcavaNUk+ACq6uHpzu5xjy
/tvBpSvymoIKyv9g6eMsJ510lv1JlIrmtGPGtiz62uIFeCEY4fepgakzKWLvmhvmFjW+2NQyE2kc
f1JzqUFpvV8uPx2PlAwlYka/A3UIXPlf84G0Z9gMvYXuplcFGRkGhVHO1fIrzSUFuu9pnm52brQe
HvI/Umvy+A8IseCSTmt9zjksK/wq3+XBlWmq7CtJcVSDEg9tTevDGok8at0QuOiuHPoGk9j4Eb17
7iYrdXWi2D2ovOkGTebgcb0FcrX+vZzXJMih+qKRW/fkJTTalyJK/iYgFw2tCcXoADTq+Awejr0O
/7jcV5ASvKmqjxMjYHKNZDPGPxriNVdezbNH3OOZJDYyOvE9QWxcvtof7SzT2x1vjKj7/BJLkrKV
iEDCuTRjoSoPcUeK03Umj8/DSj7MATo0ZT2uYPZSMcXya9nQWCxFPwItBNxsK+qt7VOa2YEWPg0P
v4MznLwUJGsUUk1R/C6AjvA5yNrg00G9RkpHPA68RKlESMWnLfjpn0GcC3nkgoLNCmD2OWhHHmhf
ELddJz3UDRZgYEwmn8scIvL+NU0jy+7fNLuOUgSRQZIdNfstZEKa03YcmkH6zW14pVhaTRTaSZsx
OS5xIXem0BZy5jDJaCdn3uxy2V1UVLfE+8Muso0/558HB6V46qxWHSU5TtOJ64S2BfKA3VPpJa/Z
zWmZYUegSf9PXaKeAEKulFB3QQLd0gr0Iade7KWLYZZLKSoAueNy7PQCvsctOzwnTEZBld79yrf0
eJC9D9zqiXCaCsrcFBs2OzeZccvMGfxCE9o03+H4eip2G/x6ax/OEn2rA5XxHN1bvlvo0VE8K0qO
6jfNAthpZfnQkBh0sD1/ZA/ssV62nU2sUE6zK0zkg3t+n38yanVuRPyCtYN2+Aoy/9cgWM0v0dm8
sECu9IibLt+OSpVyCy21ne4WqI+jSzGq7L3H6bbPvsOnkos/Ec2xZMhxGPPlBRBrUCqcPgRXK1cr
Djn091FjMZ/dD1S9zcyfNFj8bAy3Y1JkO2kr8GxpTXNTAFb+H/+3srNqJeZypljvrztcHCy1X4W6
Hfa/+oSZaBxOyg7sXonb31FMuhKgK993+CIvyj77h8Ac4nhfczrOrgNL4hsp+1BnZRntNtTKM1Fq
WL4Tmg4KBDiDxkMDe35xNCew4yzchsl7jrqy3K56PwdZFKsNboccqtxfOXA945JbjEYrfKy2K/Xd
iU8UEP7/S50t28iSbLJhvKhBinUEGrqgCqzugjxWGWq3EW18tJjGbIIy+xlqg6XebNPitmqK4ZBg
4vEt3j5mgyXTukVHDQFiUTWzBYHF4yhm/6ak2788V0S2WwhtSdpk0Wh5pynd/7ubFqK4SgOclXkp
3p8qcp52Go+639jM1Iy+g9qgbEEw32MxBSrSnpsCQhtY7pm+wDeqRvBlXV28yK+yZ2VdFWfEEY0s
xvSxrPEYVH+VBajC+7Ea/Z1lJxaS6kYNTFMCd91pDR8un3t3wGfgABQlizSPf+mPZJPdMGcbX4Dj
NBkQoa4kYGb3psB2ZcvzxYLbH+j4MM/wN6qVbaOKjbTUhB3Mnjgx3k5l1os/G/ZR4P9+FyUI7fIm
DUDifX9zmoIBUL4YqLa6MSEt6x3A7dT/eVHq8/Pagrx1zSYBWyRHKnZSPnT/7kk+55Qa/wrFB3vb
ra8RsOxF6Kb3RNZHPaD+ZubBAovTZzZStjiqKEGpYiaf0/MHf55nLIxXvVzBN5k1FxP/BVVTXm8o
XdeQZInAhfXl36G0UNYfj46kw+vrrPvRtdWLh8rBQBdHpqQFI57DrEi0ZeUrpHeGAlvwfzKTN9dk
WjacPIq8Gz3Hli5D7f6mfhjzQFoS81ChMlegWEDhgoCwnRzj69R7y7KvrVKpSZkchNIMJNgUjezy
frulxPSrteEQnysE7mtoimdzv0awMpH1Wv4VrV16SokeYsMS7m9Vvx5tBWDbr7xkef0xrLEBGE/T
uN8V3gZfcl1rAcAEsF8jFAK44SOMza4n/VeNLMRWRPuEr8TdwnAHnTfMR4h+PdM354n9vwRzR6H+
4JGA+OxCggtFc/ksLjAtHTIuNhLTHfcY8nT+7jmJGibEO4Mj4j/MCPJKjqrS5Po2aeQxEeOuZzrC
HCe9R2rytsx2PoHqgJEq7ciA9PMaTwVumi1is19VUqMY2WLtMJtPDTY6YOBr49GU1A2riasXMshm
fft/hj8Cauna5GQ0ac/rNHliK2GaiJEn2alktZ5UUYhWl1xtil7olmfx3TPm+1IBLgKZBriy+bss
4NOpszLYutdR2ml7/j+z9anAnNDDEPTKDaMaLuYOMDr343dZQxkHQz8EV3sKM5TSwyPWd4hASLVB
ID1FDNZMhmwJGGkxHF5ve0B3eFiWkbcVlb1hvjGauwruTrenahalrnsVYgvtY/dZGL1fgFUf4too
qSHSHdJaOR1ELvqTyBADbOs5ohc8faONBqVV8pLaenuRa5viWZgUmbu+aNqLcCIS4Po6+B+vWuIB
1Hl3IoySj9yuMvY5ADS20L0k4nNff2rrehl2+Xq+NKyVyVmGTisPKw75Fl5Lc94943Q1GX5M2DM/
QeN7W4iO/JLMP5mk7h2zdjD43k6USCApVuxL8jdWKK9GyUavFbrz7sx+ijgax/Y80oYxS1OoRyz8
OG+NMbGQvYph3CfcofI0/S4E9HNeaKg2I9LJOjly7BUdQ/M6RMLi7Y4yzQ0ou6JkTT/r/dNZ4rV+
K3ZIB15a4adCh59Gzy3yVjyQG4rVm0EPHTpRJ6oaKufgrY5rRWu86qSPNAWa4XwMOXPeA/hbVdlG
JOq/nqbM1OQXcmE1ZkO6A4x2cdbnlWiSqAmmAeRGZ01zHp5Wcq659e+J1jEyAx3u+sd9NGvximXP
QzTUo28DMrPMZBm0rhWGlpSW+uJkgKN/yWQFRtQMlboQzwFOofNvK6l1qiENp7qH1LalNyIqVQhw
dlJaHlN0TVuSMFuHdQccb9FBzrHFQIcAy8AObPcO1cWe8fvm0GCDKcARJRQKCKvfTdP/3scy+4Kz
F21eCX8ZAgVoyG6u3neIWk98FZyL6HwdwAy8QaS8IsDfJ5FtvLJfCLLNdS4gmDZS6MWX1N1VXuMX
KDKFBZ82Zpg2DIhJz8+B+w2liC5vo0IkP2Y0yYE1dLQ7IwjyhqNr7IEaQRYTkNHZQGvVUiq7vvni
PwlJK93LYG+OZVrA2FS925FkprcWnQ5BNdGVlqD4I2UDRwn47vycrZmrcu+BSNTmuIREWLJNFuwp
gYkFeUQE0UEnqLv/6GSyUUEw+HcaRE4rpxI5SXeBrWnWJapk9TxZo6N8CUL8cJotYIQWFD5WsASt
BMV6Skrxewqn3iQBRQzPHcMHApYs7W+GTxa0L0IVW/yfjeRxAGO0GyrXVy7CtNPv/twW/cBj1eDv
nEvqsHhGxesZw6WLXHn7lINdg1gjoMDbwQ7+tQ3929/qr5SLL99UczOX/iTfx8OF61BtHvIXr5xr
lIe+fAk8nfjaijMs03kUp9z8At3Ea2gmJy1V0LHk7t+JP1rD7YR6BAYnrdT2YoYUR9Th1YFFuNO1
hJnwiI21c6P+oHXfZgoWsI66QfbphGhp9Shimmqlvufp7gJO64/ba6OtA4FrGXj9WgnwSN8bDy0/
1Z0Ax05rrTJGsWJZvojSDr+QjdEKhokN+yxYSz4B5ERq+NQ+/oMuGoIfDgMy/C9G7a4JwYIFTGj7
/wYjkN2XNTEDO4g127B0swxpfmdklf9iZmHcEFamXaNGdwhYeNqk4nqRGSf8TuzaqWZJXv0g04L1
XpU/ksF4b9jgXa78BnuVGYUbO+C876W+sCFR4lTglbhMpyQBljc3ClSzZ7xvAdnNcWV+qkP9R7iI
fSRVAWdNUOyU+AWT9QnvO1ldMlomC1zVQ6D6tv/VmQIWM1qX74EV03NwtMFOOnUtkFehxF2LEX4b
ZFfa4RyB87ZqP3Z4v0Ijhl6naRtFG9+YdyDAi0b3grOnYdFXLVYh/vyWoi3m39B90E3eCGx4Nsv+
ogKbo0UDBA2LGax1zIeCg6yhsSBETY/rgwwKFMbXjUkIiPN9T3Olii8QByA8MTvzSh4r31kiyLgl
vr3F5oBeNBPgcAr6gstwZRrWKDn/53cwAzwCvv23dbh77+Czkus4razDyXMpUNwH0ro4yPtsv65b
YEbHKI6LYoEfBQSbT7sDJ8MJGkWVriYS8015l3KP0A==
`protect end_protected
