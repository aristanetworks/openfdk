--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
J3SZ6K3zKCKWwzsg7IfryXNiVt06SvJCBwNI57XZsorqgjGYt3zIqTQmXl03o8HlzxULjTbQtSPc
or6GbDD3JUNNh6fLs6F7nCx1HRA0WZRiYJZKh6kpB8WlejIKr67yOK44o/uPlB+ezfzeaJ4pM7YQ
mRd8OjlA44uI8fGUm3fk/i+IXpb883sO0F/p11UnublAMsrRj2dRRuqDE5ol5/dR8CXVCY/4ZJaf
k/ce8ZCiNWvRwFbnolZB0B5+mdIwMUKJFciFKPbO1de5/tPZhzEB0p/n1LD2cezq1O5GY1mP3qgJ
KmqlCFVHpMN0fZFCHgaI1t0KDJ1wYTynyRycqQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="LMV9adB3qMeKC1Kp4653n8xH/AZemgFTFElPl7pHarY="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
Be/nUKxuLZyxDEXWnf6xWFO8eLrkpdur/4m7hvhRfFQYu1w2D0pIufr9vFB5kSYen4vIMg4QWAA5
5vw+f3HKVrlB7P2dr1E8T/xyRVQCGXNJzf9CVtpCuHfw72iuSjVDHOiPWjsJcLuRaKXLfQ0iS1h6
b8vwdkU7d2ME/R/qT44V5uXddNu7YOdD1Rl9ZRrp1g/xlwr0zRERBde6FUmaRnOqN27nbLVVNku4
wXLpAu1mvKdafksAHC9VpSUt9f4ln6dfg6OX0+vtg4bcgcBqobs4t4Z0KXbu0KT5vYmGNRKcXKY/
HuMqQDrEznk5OyMzymsQ8cSyL7xLipiYfOE76w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="6XBw3cYdQfNQesjnt/qWH6so9AsQL0P8zcqXGxzyTc8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2784)
`protect data_block
y+VyZWAnLGpqOqe1fkLQMimroTedHrMl6ToW+Ano5UCZhD3XoddVAVW8D0N6qzQeskuPX5AC1NKt
fAGPSQ77z7tZbgBaS6vkxfhdscPd8ji91ZjHKfV9JDvgFUW5zAgqTMjGWgJHcEeXYMcM0FNtguS3
h/CCQkWYMH5qx/fDGFtFOYAHndSNR9bO744D54MdPVmJxNAmX0WpXASXinmDEdLGM1k2e6lETtqt
qoZ9GdUt8TztS9QAxOGXalBD0Y/mWZaxn8lfUdtN3ShNWhbtCupZ8mH7HH6eDi84MRxaHgv8AKka
NToGIvNbyCmqLL5/b7zWImCcZiooyRbXfdIgYPbTLXoSRY5wTVoXY5tXy1VwuI8CP7VaYbyc/dIf
zXo/+nJ9augngHY1mjy3Elc9LW9ioNnIkUJEo17SEQq6zK39fU9JkfqT1Kq/ZoFSQo91gjble1Yf
LjJWcAV2crpvYsySV2aNem1hGPF+HqX0AhT1or9UWk8yjMIov0f4er5VXF5pe++oO2ocEjB8a036
ZMNiXkzJ0DrpuE/T0QV1a2KQw+iDdKuO0pQpTbionx85S4ofb0m3Ng19USZlXYRZktfKgyvtv+7G
GyVw+0Zn1fAuvbVxZ9Sdongtwc68cbHooOisOoSQZFiVAZ3o8TSnQ9XpSdcDhrC08cEShhqRy3FB
isEjXvc83Fsj/5DGoV1zmXFkYMFZ0me0YfKEwdDqMLXFEP6p27Pj4Y3mckBPfSXFIPyfsm+LcPzI
asj6SVCUMECmktIr5JHxrrAKL+vfJHp9yAkwbBPbJTnf8ymmqPp6fpl+fsIn/tDpzl/i7xR/+Bwy
SeFYpW/0j8mTDGYWSIPZ337vwSr02Wd3NJBJMfZwKUNB1DsyhZQiHYs8Q1oZiL8VmeDlDRM3FzkS
UokhZgf3kVJG1Ee+dMsYiNIxKkD/IFTuyqpdTer6LTT1E3s1wAD/08Xx6uIh3G5d7CdyN67zcM/T
KoCMtos0SU79xsIDSjs5iw6oUykEtaRJeZVQikNd4ijTMMyOuX6ucuTY3QWZ10ATVoDaCuYYmqfi
Ku7MygXbbCmTjkiYVDmbHSptMXOB/ccHBOIwtafCBYxDGUR8wDyLvo1A/YgAfBfHYtfTKjQKC+Xy
dxp2btqaWvDltFYnttRKRsoPGqB2wkcMuldsTtt5LxzBsHy4Ty5NrQpPST3u9cyK459ljgJPy8ms
MSrwUKfxwEFxtC/cpt88QON3WpvBNzDBvm1v95pLNfExnZ6fYsrQrrYHtrx6J/k8A68STE8sNFOD
mTztjefhyFdZK+7bq301Im7AyJSFK3mICezIm+DQORRAj+JOkmNIWmdwpCWQ9BeCid7By0iIDFGL
LsZNsuL6gFH02dgiriqfKh3g4ixtv3OR1ChLT/6ffUFXu4gIq3/WoFikG6fMtMQ45RvnZMj11w2G
C/eUmtlQfOYI6vVj6o1stL6JfcuAZWxznMt4Zv1+9GsepuZVmfkvk+30yQ797elTtHgbniCPcxzy
IdExKrmxe3JF0fRSj+sgwAnQhTNX3h1AF6WoLL/sPtgofqIKmbxY/VmCjm3lSujPcqsxyUTz7Owj
BeZxcdFmjI7bxZmUjCyDky9GYM8ynshYQJz9veFaRnLV4L6x0TUqO2DkT2MTPIR1N1Qud8cSkkD6
54VaIICAiAkVVoLgWrW1qKm0H9i1blzkg7Ne9qpxtmqTl09yTFij0UmIooRskXbLa0SrvS7/uHld
guuChzo+qHrrkydPncq7lQU0GSGNg2gkXv5VkPVMg5zkhI/wef8gW9MjxvDAO0E1VKjJ40DWOWWI
8JChE56p+D1/D3NWtKNr/Cm5Hl3CZONK1vsK/S8xYskJ8VMcCDYU0MSYremSQlqb4+wY18DLXhXm
WUwLuc2Vghqk198S1ytHIp7bs2+nlZ2qVKP41CbVa85R0kFVb4P+w0mKT5rtNl/veItYpgYWm7JK
yNUHDX9HhypTOqex6KoqOEjod/GM58XiYxhzjwR7ujOgAfWIXGdWO4eEZsN44hflb7UGYwA3z/bX
Wa7M2c0/S55aMTaxFGBYe8uHKjXElpSWxnZpbRK/FeFodnN8UPbVZksYawz4P0D02UmOrbdSu5C/
R1IHb+k6U1n8M6Wv6h1myujgPzlKaueMojx+1ASQ+K7hainTKieVzzDBGGQO8vXFmaiZnUXfHaBq
JwJxzvjXkgaTrH6iZ2lleNNSqiUFxfFzsYo8whod3a6Qg48n0HZ5ay5MVGlrSxyOe9CtALzYNiQ8
BXzALrobu5v7Mfx5lshjcgmkClMg4PH6VUj5F0N+v/W9aZkK6RcEPuMDGTJ/6P1HjyH871j28dbz
23rhYHRrbgg7faWmAL/0KDhBFQIiqWqDMfh105NkotQaC25gXciSG0KYyoKxaNE80hUCLoy80LBO
R2VrnZoZkVlVzxPF5ogQc9tutxZGASViFbEPBulcoJPXjKQG8OhBAJwzQrudKlvxuv0LDr/ZtM7J
mzjpXwkI72CtgCrbl3KNW+eIWIbNMgVY4rxKan2Wo4DriDRahKX1DFvsRsDeZAbxGXkSP1N/cEeD
DcqY/1ET+Lyh1LMP8IEI3Uo4/s+qllnu0VQ8BjwFOLHGd9c/8J0xWZqMgd2OQjdZ8E9jPArPJUYQ
oCVJxKCWW/l9Z2bNkj3joZhbItohnTShCmVnoXyQ7qLUTA+qldk0Mj6Dju4QclRXDkYzXW7kgleZ
cIHfzZe84taoOZKbCO1cLl93nXcfEnvaQQWDmE838Rb9ilRsuHqqTsjCLhyL3JY6aL12bZdRVodG
T4hu8bwzP6yN8s0/U3YZSbb37lG1kFXAk0KU5AImpj7eaDEsixAPIJjI10Lc01vuHbBcHTR6tMC8
zex5vrZjG8+WwVXNFW7Rf0UUsEmg/AYNVSrn/6Ke01eenoKCIZzem3w3zcVEk04TMjGnDy9dNBId
KqhQRHqENyyrcSNk6m63aTlEC3OGzkT+bSqJDLD5qkwPsX3cq3jvWdG2GgyvC1/5uMDOEGasUvPu
lHHkhPClAjc2f2nz9YpA1xb0y7OMXJkptdWt7sB0+7ST8pWs0mzqXy7GztT032fsGLNGrdusF97J
+xUGn4yF65xyk+Jkbaw8qErS0ZvX0gJ0nvwN/++CDUQPyUlu11daELb/xCWb/3TI81u7QB9mCjvz
8E0vXmZMFulVsinSQ9d1J9HU90J4hmTrn18ZQCmnotNmnE8XPzZVH2OZesLuEfHy5sBMb6Xvbyr/
fuCr7tFtmkMkUHkphgiU6QPYaVopzpQHcYLss1pPWyNbQmsxobqFmFC0RMgp5z2pZCMatFbatGUX
nTYoqBUPDALXsDzrIaPwgmnRlTZdcVYINDGL8Vfw4n8qDue3yxLtWOSbmfwjm7f28wtiJS3LOBX1
rvOkYIf2tjjXBzyKDVu77ngvzuesh7HuubSrlSEze040gFJ1u0o1NhUXrEe2L39uY7NHdUrSM29V
ao2nCQkBgpmvZUr8Iijv5BSJCZtIEdrGfoipq/+VNGto8P/gOG9YPJ++eSlvKX6nYzBzeEEHHrWQ
BOVx4728ps+/nUxivka/8VbqRq61Yu56lHhjsrf1kf3dGTmahbB/rLVlzmt9GG239kEc5/05zAjP
T20pA6fTK1UlWReElbtyYLlgtO1iJj8RiD1I0hROAOEtfAIhALVfHi0XNLPivUG7
`protect end_protected
