--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
DumbRp3DEnPXoFlusCJRTOBv6xjO4z7CMgW48hyuEuNfkQVUYXtBRyxMawj6vMgS+0+AlkN9NJ1z
+7oKw7pEcf9eBP/7rRAqk/xaN1qQ1pxnRLH3sV+sd61/t4TX8hyJIZdOx5VepgVc4xsCOoSXmbx+
6eVOvGy6fmd7SXQFtTi0HARdkROyRkWR73NneTFLeKOuXHwqqxef9NSleRFw4WVIs8iZIwt6L7YH
KthWZ32GPxQqS3+0TY5fp2yXQIxTf7ftejVEpc2PkiE8qIqHyi/MEHtc3xL1AfA75r2nLZ97W7qN
8IheniMnLInelXDXHXe9fNbBNmvD1Zhe+/NV4A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="qZ7F98Mv8gziookTyAnBDNACV5ITNCQGo+kqX3qMLuQ="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
fb93F+gQlJVnnuQx1C5pUCBFau2EI2ufF1+nV6ixp92fe6UZTXO33J/2mVU8nsmGAy0FD/b8kFU0
54IwDzAKTo1J8YkPSoKRr6xnMJbfc+sK1UGdsV1erohiNbzMEMrPi4D2YYkJRUeST3h2nXNeJdmR
T5Lv9qbSSvWlfmn0tK7R7x+/6uXycoJisNJuPCo0m4DRstcW2uN56rvarW3MS1EtAdsgvkvVPKXY
E31hisLwmDniLNym+ePnME4KWaEnXqHrPCvRHLQltnfVC4And8AFIo7BvMujiBs28ZxaHBLakh3Y
ZYuOO9Kw0RJMa1l4XhGQVWBxNYAjadCTmV3X8w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="52WNoO51FebwGHxOUYBP4Ntmqt1XER2/GIpZN0GMdNU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15760)
`protect data_block
Zhq0KAyuVwEVQ5nGlMi9JNXHc+wEdZ1dMVCS7GltSYnvfjQQe5a2iv0+BplpeJCJpjh80v6SWbUW
kqEY8wA4Pj90Hag8LDNvfAc1yOi1ikiaLdgRmaFGvWnQ02ExECZawzI9CBV9D/VhB02NLX50utO+
IEA1FHkZZkd6j2/9KI+qcXXBUeqT8GTPUR95mIJ5KrF7W6f4A2Yy8T41Q44QDhSbkV6oqEpdhXN8
dH79/YlNSrhC63hu1i9DmSXzrmSv+lCM0SHYdO6UAtyvOFO3btYiXealksnOuS2ptJ8kZwe9ghli
Vb68k22F0GDZqT0fOGPBnr8WFEbQ5Yf9gjLHicRnvBzM2HyyYMHjFzMP07MZn48Spah94XUpDFtu
b7MfxI+0VyEh/izUyKCjdZKB6I6WdOOL+skeSf8XgxgBSGLShyaWElmSrHvc3RhuuAqfSrq7oKBn
GKJCgNYZZRsRLghfX+mTPpCm/GsR1Mrps97hen1cW/r6BkJhlWZhWAXV2E44Q5eBaAQ+KmOKcywF
r4gT9M8wJOCEf0TGJcoEBjdxYjmU2YJI8FRpniqQNG18l2dHcoZ98jFdZHj5fOSMPWO8YkLX0Cqy
BAOW/15Sy3gKcZRdsRiE4yFgqvt8VzUExK/k/HCYlsV8XvhOeb6CeRlTIZ0ZJQ7926RX7kLyvTOn
x2efv5AeYQOIQcIx2nIPuNOs5tZoym28ZZxmCtsTo+DyAhJatamkod+j1dmFuMDGBD78ZTV3uPq6
RO3hltM0t9dln4y8ad9lw9sHurwcNOdyMmGKEzh22sNsEaBmtAYPoK/erABpYiPud/IVaKIFd1+C
ppK5dbNdrmXxnlQZAo9AdJ3GOZHyUfHcZfHE67t3ggWlap5I+vvAPQ+/cOw4v6LSLPBZI1IT5m2D
NQ5ZV/VVpdCURXjnLXL5uDmOR8zwXGBaDNCiBT+kr6AvpUbgMxeZH/5xkcd4Wnm3msZKQg4RYpCO
ZiLGnbKUwS6mhIICECphHQAbd5OM23FBaQBH35cAuVynhIMvUk/s4s1Q9jK5b4pLzy4TehOo4OHw
IA/0JDLJSFy6at08phGtCpnQ19U6amZdOA0yqBeq+/b/6rd5jvQ4QCJga3to7N4kUUjacelbl16y
pNELSWw1w6F5LJ+WvwPGYxj9IUT6FB9OUjbed7fy/jkzxIBE63UVjsgUvfF0dZj/lebUaEmE906y
5O9XHZf6cCF3ae8ErGllLorZ34OdgjiQH1Wey8lDF98TPckRR/CaOc5mhTPv8E0W9+XoSY64OHtY
dGLlB0xEwZh7/eEQbmdhSbB8c1DfRNeJlObZeAZXhvPqB9p50vuYTbR0Xtu8P1pISTGt6qKdapux
hwN4JQlr7VfYSvyv0mGsTm2W0FF1SOcxT050/UO/B9ew+By5qnIqQwKxnycQi8qJjOxBPSM7dV7l
Q5uO1eqthLZa2P8MT0asd+ZoTCADZMN59o3GMZVRKr8RrAbTTvepN8CyVa9i3FMdPbHY/HVn/tJ2
Brnim2XZLLXbX/UmCrWmr1gb4K7IzbS4fcVwU2EXBBmFCO6PuwNFRLuNPuDZYz0S7hxxHyz7QhLe
Ck5g/kaMhEzp6rsMq2n3fMLsYxF3EcSRhK8iSCS1v3BAoqHMlBGjwGiruaUcYxCgV9GFM/wBf5Cw
zlmb3C/oEim5tke38jPm+UC8YjOKQclkdwZP7IlK81PtZrZ+LlGiDrVih23EnA2dczPQBHmMEZp4
KPDx8UV1CqbvrR50K0Ja1bFnDV2hX/aNoNG/QhiJ0C7eA6RNOqv4dRozgisqEJVrBuEdpeEFEXM2
aHQ2wUxG7X6OqLC3ATVPMLCdFNFDWT+eHP5qKlQFBCnt3oV5rgmtdpQZVohJqk5HmHMo/uBA14IL
fbza2cccg0JIFVV196IRAISZoyZ0qSTqnuIrecn++dXtjPqdHH4GBCyKHZajGIxIAQ4VygIxZdzi
lYKRQsjAuamksxkMVJWm0NC4fHaqISTY3lGYzMErcMKjGUNg4F83xRaGIQ6KFOi0dcASnW99E31H
wIp6J17QHYj56aG7KuKj2Odc8I6e1rGZqkmUYisVRoMLqtlKhT8g7qqpJnbTYEOKpYjMgvW8vAS/
aV29BMywUv9eBk2mEPARQoESq+5QOZp1FD0Drc76Ul73bDD6deDJkYe/fhyXyIXW95Ou6gf+H98k
YRHLDsJE108Z0gb4HGV8/aIah3TMBckPQ0myU7ASCmG0pkRG8XNHTBtOIggqdzLMNJ1rUwBY05M0
eranExkpdVVnqMylm460+f3DpzCzURoa4oxb4Kcicg1J58xcTVxpgMSy9V0ficfKyZld85vc31m7
bjA/z9iTp5DtcW4h2fN/pcgYJ4CVQOQIb71lmBY14PzUFuhjQMcngOuIj98WXRnrYumFaccuNKIN
Z4B/tMQHgRhLz/ZYcn94Lj/t+UkZ4pqySBOtpX1ElIIqASY2W0SoofGx7FaPPm/YuKxpMfi9Kd7R
eQoJYtIdvbPM6PDzvRnuH5NyszqQT6haMXXyQbdHFNAy01ZBVEdVCwL3yNw8n3fMVUyhJdp046ps
kxWJb+KPsU9tlq4ANNFscu93pEhvhakPD61B8/0RFH/GHpUWITohjBnKQUzO4S6PiknB+cjlDMe/
+IYW8pyfpafes/KQEJPDttNgDaVduOt0mMQ/rFOKBREW3KRfvirX42vFAifk1nwDSzQsPOl9Mtf/
nN/7y1dHHXTOsg9aUTYaX70cYrtPL/z0Oa531mLyFXe1H+Z2zsgHKEp+K0uRLobEwqcLs38HOxrW
mwnmf6xKVVvF864LTSL4gWOgdL89vkLFkDGl2tYOPfIl7glDUi3YknIa3tbOmjinO1WgkVgEggtL
eFGsRk2QXcgy6WfjIs4rKpzCcDLKD1aqgD5dC5EHaehglBxoEW9GDd5bWM6y3CVe7Xm/8KFNT+4U
hm/f7Xxnhl5kqzjICo18wIkf6ve+ikl4I9NZCvxs+NDIetMwU7EpAsCgpV4KxUFJOAkEzHV7Eb+5
XJZe17nqPJdKc8tlu4BYgoiT6Nh+chq3vC0G/H3dI4gIWYbLcfLgpL/ukwyBCepOg87PR6CKeuGY
T1p/aEoODsPA9XH0cttXL1g3bghTT2IE3/zie83C+O6qKHkwm5J3Ii4bdZy5YyE+v+U9L2S4Mueb
OluxtuTqj2Fu6ullbwyOj7OrGkefC+X3HG0h61aWJ3mHSGZRBujLd06txjPxYqZWyHgKfRy15HMp
MWl8KvZZ7ufrIMUqyN3pc3IRoHMEXrRNqpXwJLJwPTNamAZ7lPiyJVgxFVTBHp+CxifPjVqakt0N
jfwyYmrDvTXaLjn1vq3qzOi1PEyd49jmQpTXh8hi4eGRBhpCSVPoZs4/NRrD7RmKvLFVhPBzrHvV
NcSU8bxGWlDMf0s+HuUgMgFZZr/ve/8XKceAzha5cWAXR2221I+1gDZDV52+dhOhf1TvBcQwv1MD
FmeLC2VKdRn2+cr17P3Kpo360rstH2xW2UP8MJuiDKGLr+OpA09ics0joqvIyZO3RHJ9UYglXlVP
ZP/nDaPU1hYu+OqqINsKwgUqRSTfJ2G1VDUTV934t0XORIs7RHWP3okO+vNN2TXG9a780CgJmOBL
DFH114zca96EJcJgzPqF8MjAmT223oFyzmxEDP/ShdvIOAiaq1OJW2nH8wZYFaqX5gi3SzgFyuR8
VdyhzLK0Cbn9wc9EkOotRbgSHs5r+o8mNXkglQcCKHNh30IrLTob9iSt07nPRxVK3LzxQAWLBZ/y
WzSXu/GjmhkbalN6Qc6w5bqB28ppz5vLJMgvF8kNzspX9JtX4iv4WSJCGg/7aDP4NYZY7p5Jkfld
vHkWC4s/bMee1w1Tceo+y9uv5DNNJ4ucwLFj/TJxT/FxRgiTPhJmnqbX7+QruIJZBaQEOI8RQ8Te
ImQv4ty+NcQyHzFNoawVLyjpa5OJ5Um9J+jgIAof8DTCbY94H8C4DLva9f1orl+Si/fXvog3Xv4b
q59bnEh2T6osFdQv+hIjEG+AyjMHW7v4KW6LHGaInTrWCQGYP1qoOuhkO2Sd3YCMuhZtBI84wQXq
mxEMntLBa5KlKfKH7/RNqar6mLy72ME9VsK/85PQYpZRyJxf59Pww0Y49bZvZ8bFMpkmcjpVQDmC
zRWVi8/JJ4cfy/xIcGK/yhDivZCdaZhcDJoWqB2ClFrW1UBWDjdejwZiLcMRDNpQCReCwAmjJWok
aJqbPqjwYUmMk1t63HOdMPOawN2HnSWEDHGivqpLHQJFT45z/Pv5nlVFSxWxceqdutGRkqgaA+Ol
0eoocykNNzKOFyIcIIKFRB8piaiCtWT376ndvEKaQ9WzwijAvfmu3r+95OMhX+IsTDXNlY7qhTBA
wCRgPNnn/Y/EKIfjRNaQLHmqvPoSGg3Ccur96xONYNkx7D1Mf8O+HaoIdiIGImGnEbvcmsELnBRV
x6+vqkByOcf6klbqKRVFqO1xjaAyq7LqzzZWTZyKEGGbRPJfSamNiCe61ZW9GA48NuXcmhMYVRoi
+CjQDH9Z8tsLLf7Q5YssvBvOkW0EoaaGNpKmbIrzpd804fRJQzr66QR8yQL4fgZFkLEWwlp8IzYR
F4uUeO9AvRS913ZT2DEa5DS4KIs9+FVRAT3UKjtcLIMkQFsOrJ4Adv6jxg1ZluPk25oo6Lobb1Aw
sMQyG3987rsReOXhZcAo0SrdFO184Qr4f0WrPzX6zeDczAD+pS24ANcYZpZQA0M7urqYiufUjs6P
0GxVsdshbew0rK4tK7fWHcQnZmAdi68MJnqVeqyHsEAoXOoHYO1vCxFvaghBMYu36g65Gc/P2iPr
2rTYXrAR7c2JmvLOcqwmOc0/TpsK6HhR1zMWcNfLnlS3HTstd4SPmNKibK/qB5h9S6OL884qL/rl
2W1irzKzSFBbmxhwNzoYZu0WHuRxhYbhwHjpucEs9RbhqppRhrv10UEKboeeCeM+kYBEXf2vvxKV
Rl2dd+cyJF3+0z1RDcpewxUv4owRLS/7jrKPxD9dZ/vByoiE5irrr9nVNtmd2BVgsNrhWnuMdkzn
CSyIINULdzjVUjXeSN1Uld8PNxobVzwJfiZIiVuaKSjmUgOyN0y8JGlHlurR/zMiakGho3CACeQw
hPCoaXN5C/+bTGHM+aIVBWf4Iwd3HAJQvho3cpfcFI+tzWxZW60RlUg59x3smaPrzicijEx8+nmw
tDn9V0aQVpHT+nEW2zagPnaEbZ9OUFxcZNaHoFFz1aPR1gO22GN3XmlyIjcugHB99kOMCiUVyYs7
z73WqVP7CV2DSgyTuY9+Vlqhm0JgtF3SVcc/mEfveLKh+nzHw8QDT8E1AeR2AtKDNrPiYwz94SIn
FV9BjDCfVBvpL2LVIB/KrqoupTqkpiLgCtRfQPikShFBlT0HDPlXXoJy4ktaY0MK9xc7+VQ4NhtG
2r77/YBhnUxcriUJ5RBOtOMWOEvHRYosF0P7jwWUA8LLoJyE3qRerrjDEwOlRJ9+q29LPSLCIGDP
p1+4FKMB+kAifFTnIYOdS7ahnLcaMeh/cWDW+TAUJQ8y6pikA39wpF4qPiIKKpvEypcTs93mH4VE
bpLbs3RdxBetzznNfKHLnh26YYHYo5iSczOWNVQJFE0s/ejfwvfNlOrqyHW0mtAnis+KUpfz4oyQ
0BYB8XLBSpTA45NSqA+4TA/J+4hwyVnIEnl2kn8Zxg0XJm5G232a2PflNrm+WYuVMXXILfF4VzuG
VAOrGAdW9+uqJOFpTxbO602bgY5qzKGB9sSsKLUjq7bLXWo0TRL0DpDKuOjpqxE5BMQYvBYcBqXo
s5E0CNQLYEpoGYes7oDv+E1Fg535Yd4svuny6Y9oXA+rmRFHMfCefrg7qWS474X/D76nxpSYjngk
TSbR0mhDlJuhuyS1E0RuD2/unXIazqHkPLQ9riXQO4jXPQ4AlAJ4KS/lIcik3bUUjb7ZdGLvs0RM
BZ4NTjfzijBphdDch48rhvo9HHffk/6SY3H0UAQBnA3KjiOY0c7XOyTaDUDDsLdoeQV+6/5dMdGc
vvYpmaRkQ6rhoW33JcqINRjsWM4pNXc1bvzynLToPZ0OXRD2TLfeF7x5AIOy/Z9kNvXPqxsg5WSO
lnSL37rNvQ1Y70U1jBMwJTyKFVpUhh7qcgzWTRWca6yPD0ujgKoMsQ4MQV/hvkf7Xu60sK6Z8klO
f/z1vmzTigLLGrQUbk3qZwPNzrbzS2tzIJzMxlKiPRHOeULQtVlFk8XuwDcy4/TZucfkQ9cTi4h2
jnKgA59CW8OVwjsNNyEu3MLlzxxjjEzmwn3vfRnc4E7zH2FkkSvqU630+PF/UI4ajV2Fb6+I6CL6
krI5FiRs51Nqgg0WaGdQYzhHzRAKcz6ZY7IijSIEoFIJckHqJDeJnwWPV6gCmI99AZfj+TzX91t6
Xfvb1cnHab/PslOExLeZfZNcfzORBfJL8+vtGIl+Z6xzO0RQ+4yymt0yXjgFnQfFsvUWMZTk0yuV
2USCHA4H1tUVAYt6EF0xmMSlxXOxoNIklOt1jUrQ297s2MDTrkNDkxvJKeI1waumMCmNsLORROy9
aMoInZ2YQ047WS/VJECVUtlRXM1+pRvjjeE/WfvIuW3nyVtH8DHx5otp9LDHwHjWjvFzm4OrVMNp
muT0dIZu0NIdhjf+Cbg27+4vd59Vr/KA0+0lPErL6wxyWOEpx2ltu/pohSFtmUeaQ2bgEnut6NKO
vH1pDJVJt41tnZHHieROSyyYMMGzwDrtoSWnMYnfRqRq87Kn7HWwobcpc3ZvcoolZlPBV7enP/D2
FmvqN6YfvhXMSonunh5EGydNDlMUpFLtmKed9UlslKgu6e8jS94c1U4fhXSZ0PMPqTD1lZ+dQUCA
r6yn9PYdp5WhECh4H2tKHO3U2rDKTxYZ/znEfBlHFHfTCxmwdza9dB9DzmrSWqRmZ+J0m34Vt9xJ
fykENp1LqduuLHjPRy2DvclvDN84VhiDusRtTb0JXneIWGJdg0tqSLW8Zx92LBzaWH3Q0v62k4Bn
pSlmrm9egwSIZEOt7h9/FDF2EbYap+Mwtmi6YO+Sw6Z+ooIl791H/mDY2suaQ1ba3f7TajjIuPFB
B5iwNd6ZrDiq/O0gjk28ziYu7Bnwpx905znJoVa1EY+jLNLh5Ss+XYFd2h3zetvCBE2yGn7WddPU
VW9y3Vd1wGgmOSzFJyYyHOhP0WQ00Z5hXKHtNp+Zsr/vZlFg/NxL1smMbSW0zcWRcKJRQrSrBYC1
XA8d8ToZZbSrfAdZrqaB9pE21cagOKLW2e3kkABdhTkQ3+xvccVAdimgXyoFm8Ufr58dgfk06tks
tu3t8zRdM3+9p+KJlnjsBajVqmhBYMcZ/6FfDH3CB/0QehfBZ6plweaqTjBhQbvuRoZAIpYDyXSe
BuxT9rpT4I5Fr0mAsuXZuMyH2gLmy1zckrsj0zRFwdVA4N8rpZI02EryNr4/XdcXpwB/diBZh7Ml
6f1Z/4EzTNm5utkYuZ8XbZMPQn3ER+5JOHrET2WGwaTEulBVlxFH9ir1m/IZm0uCDrwYfbWnqHHe
MBc6Z6PO5mZgTx5BWWKo4yGGsJwMNLlFVPhzn/gohg30fHmF+u+/wXYtwIOY3HoWuad+vJPC2mzf
dGmFxPAB1wJ/DRzX3RXxkdvcxRHL7G33wAJetSv72bA5t3Fr+L+l3ImIdpTwfroeNFP/3ZEeAbr7
3t9aMLySZniYKF3RswhJ+fAC1Cfj9lbMbo2kKnIzGQFB87U3iKhzKxrLOpvE1Alb7JBcvUOQHSTr
+Wppfa7uEsaRintKmFW2AK07Fdb8zbb1lGmw0dAaz+karGEZwWu3yJ5+x9KShCOhDwA1GCaxX04a
8GTAhFgHRbwgz6VJRsGZ2BUY9Ss5isfAUACalaL/WXhPyO3q8gQW/TaaM3SyBIB3+3qwV04Uyl1Z
WV/WkOjxjl3rGzGM3W7b5llmuVzyGIAd2944mRq6Dwg/l9kt208X9++hON8N+WsfQnArOnMIbjZi
jqZytw9+jVN5x1/WIwZ5iG3p42bTak5ZBp6W2W1GVcnRNjavsIrkmM6EEOs/c4pgdvRcNBDD1hkm
MtprfwcnDK103Dhw+6/Fm52j3upx/zfgiT/0aaFR0+yAdXLaGd8jgMqgVsElihyvrRpGyq8GtgC1
WsUaO8NmVOdA7MlhWR6eFgk49kbXmuNZWGH0hMMF5FiQyA76uBzsSyttEzLRBQsonAsJDUenSyGa
LhcoLrxqh/jZPXc/FZ22M9upttoYscrjFG6i2WsN3eNILC5cJfODH8F8uj7S6u6X5tECfw/EQd0Q
nZKjamyuQBpeRBOazdjUaU3bU6OX7omdh6aqDMHPK0DJ7Cdtau/kkrcK1HTlzZhHvbjxSPnfne2H
gw57ZG1VXm0MatTpC1IAEgvfN/237A9Bn9dAHuUL7nXZ1j5/RAJFuar+PUas0cxsiLrLdDjXnLTc
jbeEf9AbUxkTsumeoGnHcwpBaOfF9MYiDZ0G3kmHbtsuDgN0SzUdeIxSP6JKb5ZVq+8JsU7FN9bt
WrO1gAQuupgABKAAsO8TygCZ1/2p1RrK94NbQG94TmW8VAOzNxXb/+TyvMe4qz7M3CwO8ZdS28vZ
QMVtkC9INhrKe2zHeo88kU4QSVH/w1U2apAV4Kd1KdaBNN9h4TFJ05L4I3cSrARd9RdgXwhx+PZF
8Vb4scZ4WWrCBe4LyarxZnMTc/V3VqDeMbSgvP3kPgOwin4GCMqykDIwvvaV3BMgFZ6j9sN7z8VC
i1P+a4v8XZ0+THBwXWIDZLVgIorTvvKkKzu8GJC4SLVhv8C7KB+ZWQ6V44WSrTo9F0I1jfJyQAIQ
fLDQwZvWsHTDesaL3ovk2msflsLbJMtLV0/aQ+yDEEZ6TOSxtKZ1Z0jL8lu9C00JXh90N8ntZRMH
gh60Uyx8QRi8CKIJ0pYG9N28qnnyG02eIBhDRB4rR8vxogGSU8qxnGpRD5WWsqrB0CMlmQW7fXPD
n6v9Ntwktc3i06iPYdp9y16IHnomZPsMLENb45ML/ugtHbc4uqiZ9owRvARh235ie6QLQSn8s1Nj
dsnJ7QzWllhADyN8kNYI8+Ax2qQ3ZwvFVkQemIF/LEZbE6/f3nE0UY0pQH8+/7g3M/zDPhbfSLp6
urMjFJ22dVn8xQgMOXgOsKSPF7cUiEgZ9VrV720kpDI2U50xqiFqOgg/guHmxr/PfcihsK/YH147
OWFF5DYVDNKtDYyjALT2rSwJ4PeoBoHKXyUmVDZG+nklkFmveMiXs8N1DvlEKljKGBc92HeC7WW5
MLhpLKVDkaaIyOKl+O3yypo7LZK2rO7YuSMFaoHwbWZghgSbI2fa8xpfKo3YBD7PG6o81Fh/BpG2
sr0eTJdQBiu72yln7brfLE1Z6MHCc6oGqxVmBD8TRN2qO1Uu2ANvrBJlhKHRZghv+Yre6lej5R9T
ML6zitixHb5+Ej49mO49CwwCVgSuWlSgo+VONRGUSdBGnQWxP/OzndXpKo0mzpjI3x7diNMblwwN
Srvfv4toxT9pztZYDeKS/i0G/ADJBGrSJcCuPGetznM5nNGZWIeF7Tx6kiFAb46PyhedaN1EK5QY
3p+YpdZAIFgmoYiTmeUL82fDXCa7bfGGQiv7TfZjhljrtK/CO6M6LrE6ESZKFLNILd5s3qp1TvS6
yBIfZjZTwJkaLmA2ywE/YBmFpXV1sJvmM55MZMygVdbNh/m12TIpmXYDeTfDEX+PBz2AXCw0JAAH
a16jx6h4g3acxCI5La4T0DlLwJG4fS8wCADyXCY73k8FOic1ofUaauodFfg3FjW+3L1z+/2wCCnh
qT47FvEhvXw+pqYvwgFnKx6uj8BHr2LPGUZpuZVwZvNUxawqpI71laDD/YYmwSO0d+s0uGRbBOCk
s5/el+DjB7w+AixGTRmHA/hW/A8ss04y1gbej01IPKl5ZohaHMnrXb9U0sRCspIJSfAXxR7/4rNr
1Apuv9aEHyRIoD7jNsmjjw/EjK3wKD7ItMcVJGByfsVllIK6ZFuCxXgRRkctoTW/1o/Jn+WI2R2U
i94rB8f9uDvtECXqkO0zajvE+SZPVeHgBfyEhD8CObYavlbDOvwHpIBzrdTLw8pFMbLX62MiLmXo
gLKqU5xUVVEHsUP2gkQahdea8mNz2ZXVpuh8VDMqSkQ7xeXAeEOBDQZhJt8oPg2qOzuaV+BF5bx/
7khv8VznnTIyw7ySLwwpjuDn1k12S/S1yh3WIbnbKeH7/g23POoJFol7hnakdsmdk+fRKRv0WOry
tfRY0uOiTqIE83cH7/pMJzwsrIwDZW6iLTNhQfPgkk85AWTY5LKKDUJUNFmw3fUX7ggYBoIuLGu6
XadO1z8trq9IXbcvJTFZJ7P1FDYbS1aMKTzE9sZTkgdVh1O9oBB03Sw2e57iFHrTV7vTTjz6T8W5
eTVmhx2oS57ZQp1qhh5J+Jrd+q11PttYYsP7xxq9zyLcdoImSv2kCrcZGyJGKf9HUuuc1C3OmLGV
XoeF8MaW8Ed2SGFJTUHv/cnBRIj/mX1arr4RMV2h9ZUY+vr3qbY4R1vVJXK60tmS31i4v6SR5lAb
GWBniqg6gByJ9VzVcCMBwmuMvoiy8jU5ZKxxAZzBEP00CXGQ7IrR/lfrPnGBNgWXyo2DSr9/UDA5
h8vbZEc+1t6QrWJKJOmuyduBw3zs98mjQW8prGLI1GaDjTDIMEhdMBzeIa9YXNJjcfcD3TeuMuWw
9c6ahwUNeiTPMXehRFY83cZWmTQHPzj5bZv3puXTmq8mgs21rh4j0yxeJ63tH7JBFt0JZ23937vk
EnGkMagDcO/eI9lOX8sOz78tjs3TWyNJtAnqNa+YV3ok8PWmjN5EMXgYIpUssGmrMaJo+mrskvCH
dTWtitamkPW7Osds4eXUKnPClf/MHV2m4gXnBRi77sl3hY+1N1DHS58MWBH4MBh/WcZZk37PBSyx
kxbILjJUflzg7qIzwmpdyQWyB79gD+ApxDxSa4cN/1laxrwJAHlGj9HW2py5PtHtLKzrZzp2d8Kt
/QHVwDm0FgFqZPEZ4jN1JCNXOirCFM32FCchxh2OMKrYL5VrbO88M2APwFJ8QYbj0U/2cLBJ/xPJ
Xt5YHUh+lOp+bekRaYVFZ2ENwIcsvlMrv72BZk4672FITTG4FBwayc1VtuVvhGfK5/UrNU88EDaW
bjF6uh8ov2oXWIuAo+QqqYHeKB+jeacnaFE5z45cy2UgrRC6cYnvHiL0UPjD+HFReWMhx22jPJSa
4HNTyP3OlvNnZQmCVYPsSESTwd9kZlI+4Rvg90DlN66O4gZag1YxwoNaT+Vf9n61ZkR/ytLQdWQf
uK1bCNlJ9M5EEqZegzgx4WZ0Cn2FlEMeBEy1Z7Fzpv+Gn3sqn12oS95OBmMLmvna4LndxDvt+DSP
B/3WyWTSN1ZjeT/nPafn0f6SZviwpsvk54JSA16blhEww4DCWyBlXusfPnyvGLHkycCfP/ITRHei
3GIKc7m6UwMD225f9t6bP+BsDQULNeXczHFSz+unjNUiz+pmJ3aMCwv9rLtF6PBBkrDOI53Z5dfT
pdv1ZC1471y3HZ0dNJFcUkKf4tFRruX1uAb6IJzhb1jvU4BE/PIM8WUR3IW0SwBHvSu+KxTJT2mt
RqVo8xVvKe9EsVfZ1FEYV5P0Ii4TDeQeUZ+23Z9KU3pP1LG25aOG3LZZH/fMOhL3I7VYF5/p7NLr
r9+RC62zwUhbqFMRQuOx3KZIPD8dM4z55uLOFsAkpmm6jBVap7ObttT2T+BFXEQiWR6HIeUb30HM
YsQSyFvnwF6PpgE0NMKBD4BSARFcn4bqU5Xtk7xKQ/g0bjMz4/0+QDn6b4FhVymmXnRtdy7TA9TY
zcf2rbCrfmXDNT40BK9rCFnScFGqEJd0uOAwCFYXwKTe7k/Q6OqdgcXY/2HUehglGGWmOeQoppm/
LQyTrDdrAdxNvOgR6d6ZNpBS0xHed42CkOhdeGfarBhj9JXEeak3E3nu1n+EwDRxCbsSyXyNZ/ot
IZRdo3llMrkehT7aw0hNT2abSv562geKWgaCMMEwWbxlhJeGBTCPIGMiU88sR2+OjcRDESiuhKsa
D3DC3oeiaG4i8Qveo4EKU/ZP6Xtlq++uL4BYcTSDY3Wr0hV6O6OJOV1AjxCoy+n+hYluqm6n0n9o
J42tLe3J4tV3X8fLvlcV5hBpWdDY41HMQX4HKeNrlA72KyQWscbi/02JArdj9CN5GAtIfh/ry/Kh
xznorpLZiFm9UtCfPJFhVQzkOc+Xgt7tpR83UL5GjFs6d6geUaruFohLg9OIgHwHJzIvrvSAMKKO
cK9dy6nZl5Hh0EswtSUxqovtreHTgMAEGFZe17Pq7Nr8FJSGRi/2UiQd0hC6hsiIZDcKj1IDEN46
cPymmEIJYQUO6pyRUEtrgDfGrL9LSfYWnM4dzIHBCNMnu4zO6LV5B+9eMAMxz0B8vV5MEILmBiTJ
rJ7aUNRdn04JjVGQw4vREXev05RvZ5M2Ev29XJMICYVL9R3KsscNgYVoWQ+/mTwHZDHFLVr+SgTK
8NmmnznodohIMrUATJayNs08Gy8zZv12DvQlL0Ts+boB/HRYGbKXzMbbIp8FYyH79pgxpT8jVWdg
Hr1x6gnUwBKACXKZnG8AXXw+zXdlBnW07HGa+Z83DPLoXN+2EDKRrZA9LvYN8CXL+Ca22lX799aA
dP3zs+IvheNDadFpVZqbUEY9xdo/dSOaBfjl4QqunnYAOTvgpbVDyWuARQ/z9VikcVkUBoq8TB3T
TcgMfN/p/ttWky9xgDdpZ6WvbJBCQDmmkmuMCtgtIRsqjFqy/RRMDvp5bNuY72N6E85XEKzQULdY
L7tn1WUsF1Ks0v03BFJjWMA22sIT+aWNIzjUTJs+lm0GDWP4ZQU/+dc4gCUKw72WTkWhmP5eh/5M
HLak1kh7cTyY/XwyevfPtkHIKUrnfyapTV1ycQP7H0iQohkpWiDX6YJYmYQH7DNW7be7lbPOoShZ
OC3loFwh0VJ8iDCA7pfU6c5UzyzinPFmVOvsdHuUkzhFH/Qe6fErjWmn7z5UJ8/d5ST26xesWU8i
30U6iv8Ee6m3VhUKvm5XHwc0md/qBLRopdweX59fYgLlp3Eo7F/cwZxUmdMsc8K6rWT+wBO99FRy
7CyAD6D8bbEyG0OaSZTjpfbZR6YG61LA1/RaXxTH1DWLwCuMYUCxaJrBaf7F7IU0s7rQ+7curuzp
JcioEtmpk9U77dtweCDb4sUeYqRFLivkQrR9EkO/8aPXTUYWE5Rt4T3zubBIXEovLDGAEzC/Gt1O
L2cKDaDDgMBV4Qf4Ra5MLaEUMk7xptXo80v4IpvpuIjmaIIoc1QoUgQkAooT7hmWRU30VyLyWdSf
HWG9Ry2tkobx9lo0b6/Rb09reL2G1oCod7opFmu7eIe0SwRM0UM1dGxWyMQMT9S66oO4w2ht3rmc
Bp7MvWdSjZ5WXhBRhanpWUBrn8Mwcn3QdKSZFteWFXLS4o/WIZE3o98arrwA/mWyB6lz6UkvEDiH
+EdXp6oRhhDEuSnigMre1+EjqpU4ksDhjt4yRXLpHI2eRZwbvpx2hq10px15r7rT+PPssjDqPSFS
MrpQ6HwvQta+1yC7/jeDKDNMMPfhiut3L9DaryA7eokOachqNwhvy6wMJpK3+d0ndlEX2sHtUmta
XLnwTnv6MJbqZE+uO0XD0mxk5T7yIJOm23Mw2QgibZKZCrhvR7U76huLK1XI9fIAcwKEph2xArzV
OnrgZcKJAp/Lpd453gPTslu+s8q8Y0qpSMZ++a40RulCKpWbydz9JGL3DPceqeGb+0XgNCOJZDiS
fPNPfd7fsfu/wHqgspTA0MPa8Ix75r1A7L79evyXYzhLHWXZnEmt+4LvXhkzsMKyIim1oEmuEaGv
oS3BHSfjKkvS+iywsumGTFbuzIGFU8osOIkoUwv983e4/DG4S86FJrGTmWOalPHuQdQVL5qeNqAp
1lWsrioKEu+uyVVk7SAMSE6gnARKIBxa3pLTILlGoydylsDtFEBzct+UM2mVD2UBKKvUkWrfce4j
h2bPi8AHlKgXvqjSmD7ONUgkfyCQrKYAgjrhcKjjeuqjcVyRdwTcnk8vqracjxcPfglN5qcXtpZh
wB5ox9Igz6bT4CIArT6Xez3mX6EHPzphs18L9+0K48BTwKIrTZs75XnUhpKod5sdLCyb8c8S0zTv
+SkBJ8+6f2nOe+acSLluXRA1UUkSPBPMR4W651KfjIy1JPcueMgyjGAU/MalqHLTTLU2MYuYI4+H
cQx8dZO0FoycKSGVP/cFHODM+SjNpo+s35HSA0qFfwc86fjbxhuuYmG0PCtEk1B42lxOPlX1FVu2
g2yNGMNtGF3pM3UbvEZ2u0UHhG/qDbWvCOwr7xwvABtl+bjFT6WR8Q/UxTKZ5iV1N811WF25LEai
qKIwAT7aMTcnTkvxIgjsxW/dP8GgB5Cxu0BRh5LVCXB42jEuMLQwQiv2LLey9Kunw/+gjVszYk9D
x8LlVhWb0OckXXBFXJm8tILPdPxmeGiI/z5o1BsgtlKkuBFYlGuq2Yrs7zZuQF9aDhr0Tkw33s57
VFobKOxZifpuJk3zyGTuSC1f9lV7WxVuGFdROsnmJhM8CTFrGGfwsTvFxBz3crKVs/Mjxaf9h966
PfyBYciFlfQiZ/B030OsjrRmAIQ//Sb/6id7oRdmaPgzp316ft4UhfsElGIpBX6BIR9zfUOwPOSi
kFrXYzkw4ghodBETuJWmGCCv7iTuGpusXa8FEbhoC4E5jwgGmYki//eyh2HHIfT6YRknrt0itDKS
oXiKZhSi/r9ND374STMBbpQAwHigvYUV+Cu7NfGMxBvP/1Uq0H3FnsJM1V9GjZ3f/pPNso48STAH
XjBaGujXfEtyYe9k3JkEQSaDHOQptXeZBCTDHvX//Cn4wHD4MP1hkic5OMoGIwjdStBbh2sr8QgG
XwPGVXCXVjtB+tpm9nOfYe8OkEfvAHxqfustTLOlF3BtxFTqSvK6GyvQk5e/LnH88AA5Ege2y9Rd
NNWiTbTrgWBAGiYVcTlpnEhZUKHbPRuRcoeCSzWgAL1eua9M/8MENIB7fbzxHJ0aWWzAxucFNrqF
hnS9YKiOCi9vkOYOqY/1XFPAm5R/pMkZnrb2oCuqieVp4LQLl3czdj5ER+JUIp6vveqFqKRAanfz
aVRWW8S5mT8SHknIQPBWx+qqWUeVQYdtG0A3n8ivak+yeG1UyLMPUHfnS0TmlgzmhNTTRFUGOIAT
DWTWHvDZxjzmVKb1RdW1OUG/hOSjv74DY32wtxFMupkhsRpNdrD7hpVxK2xZtxwRZhdfvrQeVFhb
EKWKG24bBP7ecl1FMvZlH3DL7rkzyVJ/6bcBQwsh6c2SkLQVeiAL6HNZtZmUmC9toNvWpEjv55zv
kq6iu+3P7sRArgR2+R+/XYAegBq9QAs/KVCa8nI5JZ3laikcRo995KJ4IVVOon9nU9xSyDHD1aRp
bqjWKM+qwfHUaB41mZvWzGZ/lUrTh4D76DVkWVeQq9GdX9npb8xyTF+B1cRaNX3BRGAOyWA3NfYG
4itOS84/kis5Z0BRdoMrzDyoKIw8Wb6amlkgIniKUdTKhLeOjTrR22e6MWrVVh87HhMVBh+ap1o2
GIjJl+lxFVj6m3ydTjIT/ZEHREQCkwBpL7Hv1vUnYCiRTX4tTgP+qJ58U+XF32caBkE8XZJ7LR77
dzGcjZO0OF7P7d7fe5tMweYXU1/Ds1P/IQ8bDQ2h5L8xWlP1HDnoK+tnfHR61s0hymaQ4IVHF38u
Z7W2Vnw5bIphdXUFlKoIEsFFupYGeB0i0kPoBKU8OUkO0sGQ2QZkk5hvWftnzSto+GMBhKgtfkmt
2UkYkW9Y0zDQ1OZPjZo53eQWkNoJyNOILTRkE/yD2NXGYDK16w0zprP0VuZCvx5NXMbresjwsDhf
O1nkLeS8cZa3mS3elxkHYLGZFhsvf8r6M0CctVxIeECOX1OTAkMRDHj1vIyjSgIYDqwkMz/gcb4c
8pOdUjs14K+dAvTHZpHQPydStdg7kfU7rAH9cX9ZS6NBGwZOdrZEhGptaiYQ2vNauDWSw+Rcv/g8
8X4IrzuBbjzQUFySFMop3aoAq7n657rZubQWy3966OXEocGyg+veYcD/13XZi/hjFrXnEurz9mfO
+HiA8GJQYPQ81Urr9q0EiKqj+AsbEgL/0SiQotinsA/Ky1gNyXeXAM6B17WLuD+tk/wJZk9ikpfM
6pXfig53Fov7xf2ziFiK3QT4koXLbnbYcG6OAaqoaKec9xPbMH5X+l8PUli76+hlFV0jbFPl791z
5mdCNfDlz6mpnO/2r4VtMEJdaU9HeltN1EtgGY1Kdzd0+oJols9xb6OD794HDsuOMjmgjAL9TWsk
OatlXNromm9vN113gmDl62DJkUKdV6AO6AmYE2f98Wh7SWkrZ0xEo3O/ME8SG/fefHeq3sXg0EX8
mj236B4i1mkJTqfkJU5lyuxejrq+1ct76j2Hn9ZklrggJp8M4VTR4jN8Bt/SN6GR8fkOq8rAPz+L
veDspp0v/6f2aP88MUe8u5pV2Sp2gaQ3+ba3gZo13PL9QOMiA9wLGkc66cEvOsphPuS924q5+O28
dF/3E6S/8VrOO1FTyzrCcOOzQxAljPLoIQXJPuHeOvrsRr2htGobAIo8hbgsWTd2/ywT/kQA4sMR
+FLw9XuMXEFjWT2iakEQfYkDB8bS60B0wGUAVCASQAfmsbMH3LoGHBI9d/L9TAAE3EaoC/LBtYU2
UpiG53QYTvJDQFIMG47FgAi1dcbjZCgdsJ9JDzTuJhvnLYDhfuJg1BBuH4zueiiMBmE4JrxPlqEj
UOmuAYcTavB2E+WV00PJ7+W02kxc5jECBTnnUoBwGOjW+mDDDilbBuMogsjsbVezsui8ocCaykdu
WT1npjdamwY4LSKJdtQ2dQM2v4M8rqd9TA+SByYKfI+98+YSpUngAJD/mjHpdt5dqXe0pQqgR0+h
2hrXrwclT1GsixV6t4n1kbPzAgYqgHIp2ygFgrpEjAdioUrBy5Ukw6QNp75iBgJGnoMMbGOeG1vW
JdSWElmgmi50Q4WcxEYSndA+MCm4RrcBtvKI451wNY+bm8gigLNjwL5HzDwaBRdypTTBVBuSGIIQ
ZnT+0aLVFySXm1/d5vaEn6uuSZoN8RhW9inTGTF3eX5qSbQG/7RdkKx+iMviySArqu2np+3LUw0i
6z39Nr2Emg1icivodQSbcyHjMWJfOLadv9LeEFhsQQ4VMx+C2UyNwo3Y74EFRK0jEaEkJb1ZNGnc
WfMzAOlK1kAr7yUT9l9Ap73xEz3Kk99ipPHI9Hdk5GStHtotV6U+0j9QKx6m7m0lrfkIifaKzdC2
WpWTuWWb4e0NfEZSXuY2IaOy8dtVjMXgxJp9sGBSUc4UJQvopayPIH7IF8QEtxDHUfSErvKwqEMW
4rKSd7Wnx8NLeA4RhAAY8oktR+zEx8hFJQXJATuQJUjKPLJOGk8sTeXeYX3rZ4OO49B23KaUEHja
QIFagrQZ7P1xlyDi5L/XuGhjzDiUhd0g+tVdRCTvHRsVB776X/3EoWBc/IN+Xn/0Lm/TxMWlc4YV
gj94407KtsUBBjdUn1u3XMPQGInq2U1W98rv1eeCgY2VUH3DOidGdpggUZgjTR3eg8Rxxw0UluJy
ax2JenddrUjHssU90bO70VyeQQkdmGdKsc2B0xfauJ+X8EwoBTL7A/vUS3sbiLzgypbLu7+x0JhK
oROeA5ueomUS2PFf6Qg7zvI9U0HSf47dYWU6pHd7u7D4uesl9TciTwnq4rg2mJ0PC7ZCVStuob9w
S6+07V785uakekYuGFUIrHwW5dbvWKrVj4aKJO8oH/k17okBlWgjpFUiBBdfGYbvDfXBxFXYANAX
j+2xjZUhdbbFull/7rb99S+0gndR75ekD8Yh82UkhPn4EUXdKulaDZ3F9Gowvgop+gSPetUS2A6C
bJkSvLIsLOLwMFqwaluJya/xY6ByGeZYYvghGalEWHXciVAx3q+m0F+h8UXl61udPliCFc566Aye
BggZbmVMYRZ6ZANPJ1KyanZKMzXsh8rNcjOfVUTK8YI4X114VagFUtsFxEz2bm4/acsu5V8vQnH6
/Tx6Z9ohsJ+khd+LodMQ8/yHF+SNTSVT5g8U60Z88zfC4APPrVcywiL+zg9ylhCaAXJWdHJ4R0Yf
ZwynTEwWnaQcnGnf4r7Gs1qxswjd0iz2TiTbpiWIJUbX/Hnl6741Nwo/1sexVGs+UwOgWkct4hih
pt8f4shu3PtosLWIZ7ZKQRSXtsxH3rS52AJofH4rVgEK5DHAacZIftWOhG1STAbRQHRl7hEwsyik
e0PzDFpvdRAbYdHO7/LOfHJ+rovny/w/TXk+FWNQQ0L+KWq7HOg2gjREHPRpTRjMwWWcOHpoXtc6
YcllI5INzjpuNLawesTB2tk4oDUI+sIgW/iVIfg1lrh3rcYQjMVsWAFFadF026mfwINQPn1cwHUd
tXQRxGUJ02ixxGb++bNdx+kooQ05J+iHdQW8fWIpBUIxe9nPXLfdKHa7SjOpiuqTZyvIF80IBV11
B2uyY6hzrb4tFTiqRNm82+I4VFYLIqCoVjFcL4kSjIoyfUNNMDfjrD5XsE9S0MJ9qLC4d9uxGBUm
oCdrdHhmKoqUAr+Jw85ANe7adnjLC2WJkgGBLnw5YNsW9uFclWj2qDnsIsw5PmYgplRRz5eoAbAQ
GyMycawzVyy6QaawnEDcQDSI3veW3Hm3UE21u2wxNuQRDdFAlI6/LHJ32Xwv5PMZ0cNzG7aVmq+y
R56AlGK/aVvpClvhMoZKU6BP6znbHWFXol3Vf1G5ot8kmCshFzI6PQeWtN8LrR07fKjj3cwhrE8K
C98JF6Qdry0Rg+JwuWHCdIXeqYSRbiO9i8kZbZayqUT8w3LrKxFHTGXOIxU0xAbVYjTUAPqOWFjM
tSGMbWrMa4PKKXZIlTxv+Xm5qCEnIeKp+mSNMg56vu7Ley8Ky0GXd7NJXS5q+l0SwNNLu0NBWgWy
WFclYQkTcQf+Qkv4fDmtbns/AIMbtMgnUItnR9BnNE4eXOqP098PILLUd4krx/33eU9pf49QwOl0
Z3E3jC0dS4Ki/dEXzZXuwSORy2T4XYwWpUuOmG3LOJn+0GNC38+QflrjwZ8eGz+8OhzqFY45+zrj
G6n2kHU3s/2+7b2WIm3gHly4QMfxl2v1wRjIWEKOOEF/dDcd8uNN7Rpy0Pom8UkJsidhgnw4F6Su
PG+DyBl/N6PIlUbyqHJavY8SsMsZ8PIkuzUGu/n98wxUpAFE1frsrEQA90hjXJ7kyZcA3O6NLFAf
C0jnpOmgAiO326IALexpxNdMVoEeeBWAo738rQ2NRpL+2KC58SIRjvUr7EO8d4qf4uvbe7ncI2zI
vtRlzPY+UQuclztk8fjFdw5bWEmfkwUWFkJFzNqv72DZLzUFP+Y+/JdFIoIGGwi9yGJVtKoVaeev
bFhvBYJApIGsPBJLV5TYP2bMsLJy2yBqrUvAcpNFzg5ZffCHX2ZRUmbDgAJdNlrApWjxFggS0zYU
OLSYxHIS1zcmR/ZFAlT6VAGEX0jKPPuhTvkDGl/TEEWX/ZI6izp4WFo9dG8eOtuPzmm+Y4+Uwd+L
nGKwU5ggJB6T1vY1+gFl6wWHjZ1fpH9UQfaC0/XGbmrdd2znCTx1F/0KdcThXZ5DR2i3nG549Evc
ElZ8zHfK/9fg8weYurk4FwgM7wtBpXN2cw0Sfj8cCZK0Qln2nqjMRmJjtPfOWfWBsbIOINsNFKsD
9HVrXTRc/vg9V8Cnz8KrtpuytgCF5tx/LRkQSVJv96AnOjPLH8F6mqruQS4/23BLHTwqa0+aNGRt
HcRYr/7OCDlBrZ3cI8bTXpuO362tI7bBcZdrgl7UEc6BjEMwOP6WGpRfCu1frzDId3vXYP11SCqr
vrBMVjPb5C9os0a5/ZpKfmaIITNrfNszzlHUN7Tc4GkO3+EdbVZcF5r/6yqJOTnZal+vJZpI/AyE
IkXqbYI9g+ZKY5QQmyFBMSsOve3N9ucBvnAVwI4B7kWwzQ8CthJJfQkrJ7GZfmbjJbvRZzqC0zoT
nrhfMMGy/af99AG0n9BvH0zA+gLj3gv5DBSytS0bqTYlpp+O09noYggf4TbUprTe8cRak8CthaD7
SHGk1avyC6sYLJqwZg7yXlY9MVSpHBe3LG9RaywxkI1rj7CkKsaD9MxF+PqJr2Q7C2ALdBCNrfkO
lH3IFjYO+lUduSBeg4hPSfM11PvWJx3Ar7YytT4Z7O/8LewbZuZhTQlSqf4o0nEVGH+cEI9kmDbD
1epMAcfQllnNBjInU+lmdNCiObBopMt6tRycClLoOT/JemzYGhvNl/Jjy4CwXA9p5Lu9zec3ycwd
/FUbroBQdfGGzAM5vD7l+HmKQX0HKafXay6uhrKYJ7rkewecGAVSm4XcsjeJT6lVxE2VbHHa+ObK
/WfvZFL/NE6xt74fjWhHsh5Rj1+qFJ4sno3zR3NS+EFTAbPJuMFRGSvJYAUwux1+umCjcO3cFLP4
4BcF/5Fzh9dGYQS/0dEz9jDySfx7ANxt0BKWCVl2O+xbwFnslQDKStfHiL14vGmqmw9AaLOQSEI7
UE+HLNeNGCABsCIKxoCqDMtO4jKAxEXuWarHx6tsQKrQpkMMWDjyGG+YuGgtSPuwx6cTkkkyrdOB
vx13OwivxMETMTJM166AHQvQKO5kH0GogL4+AKtDBjXxeE7/24WBHmNU2/N4VL9pYShdbXPzcZwf
dexz5ISiUVXeL+cPl/8aNSpg9O6frwa0uL1gvrPPtWoJzRBAHqZBwQTqsTwzOQV1vj9pRRFGomnF
YcOatBLR8AtmIs9KH9lvuzKlo46ShYRD/6sRfw==
`protect end_protected
