--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Jd7/oMv0Okf9k4MLop3OwDIKI6nvyE5uC5IZ7JogEQWdhmy+VpQWbRpAc13jV6iBwP39OmB0bZiJ
Bm7YgW6Uzvij3U5fkB1i+RdzK8J6qXsHzFq6yn7lAhtCSOmXArVoNGwmh92ef8evY+9awlvx6Ztk
NAR9Q8PU6AQnDFxGZ0WFTdPzYSLpE+90QF5c38qpfl994CQxiSKPcyuBj8DYCKquy2+ONVl65Qpw
8NnsxcnupcHaq4B7/WaxTmBMlriHP40cTcLYvm0d9RTNC/RAdwANjScM5KQU7WlfIM09h6ujwDT7
HNGEbcLKt6RY2AUGguQbEIHRUiBkXSLApjBUMQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="4oehWNb0b0ZA6NmUd+QQ5DvaA0/4hYdytNNCQmtIoDw="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
cxs+/LepX1oZ52VIk5SQZWNcH49CMk7jCrNyusZ4qtyCjphAKkRUNY/H/dZoMYAZBDCOafn+VGRJ
yD1PmM/ERf4yNok97hgky8at+TEVc63Q4pATmD0Hkko5ia4S5/fHcPBFH9Axp9Hz0lLoEd8bDBL9
SlXyXgtuxVcjimqG76m6JYOIHGWPR/z3Ehc9bLorZU7EzN4qQDSMylcQCcjpG4VOkvsd6emTiXlk
CnJmRGNTn5I8de8Jlatym4tMgmw3Sy/NYL1UQg30h0Iys0sa1HYnCcO/3DPs3xcXtwe2yNfdVkH0
kMMCfPlBPepA3/I8clkg1zoq4PPKdNsTJjfUHw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="0GKfBYI0oPthM6XGyO2T3vC/82UE4hYGVkCY9mBIuTM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7280)
`protect data_block
uqXsFne+VLRQgvAH/XeE3QDnrU6Sxhz6n/94y6V/eUL7el1segIXBEexlU2Ct/sexf5jnVmNBygt
7qOrP7/FDdC7GWrkipW8e05r+oo+TdpT39byVkz93XTkoxjxS6zzczrdwis7g/NtMJkRSyfqtub1
RgkXkHC6sxXOiw9dJMBYBVS2BO8yun44Phd48Xs6VJYf8XkYY7100c98yxkxueqePO4CmNeB4pcn
9LlUDLjceee8fVp3ps11AgysXD6jqCoojagY3b/unR71eDk30SiJylU4F47/K8GbZHuKnYnT2t0A
LmJvInlYylIH6stThK/krT43weAD9g23NBf6Fqnbo8ifFaP17uN/z04fHz+fWECB34zUIo0APNCw
m3toOcRvaOc8v0dUsnqHXlD2wQVOtm2i+cwEWxa89vKDSM3IGoikvl57ucqUkdbYHNhsUxwr7b/9
XKN8PF4MbANFQAc9LutP0F1Ay2Oiqr3R4v+cbiW1/EGcbgrHunaMWIQ/LJNCNH0oYAyzSwXufGNy
Bau02zwPWWBQpp8mcXe7bM6TsuNFadQ+26BlgfcBGo0qg3HiQjZI7rGd8TY+3Ve5iPZJVr9310Xo
MsFPeCcZ5cobWpf9+H3vL2ekmWW1WCa/DDxL+ULKm/7xNf/drrLwMbaT/1pTEcwlprAPMwam7VT0
o/fTnNSsu4p5ZPrA8OVc8Apla9zGnc8KMJCx41u1hl5/1fxmcG9sfR4vVde8Zzt94D8c/WxrajUx
ecGqIe1Vm9mj+vYFZnvGJsQLqTxgqfQQj0zj5B8suMMpa1+NA1Ky7QCZ99qNU/Q/1gWSI4QPzogC
KS8QhD72qPGn7JlHfyrVOyyuEhlijZxqN7OlQbjgQZEoigSuqDPJDWLK65SwMGfVS+uhhmP8VSnV
ppRFXGHUy4M7u9F2opmDzFpEuhw2FwBQNdgL4Lvyf1o9Y2uUn1Dxoz8otp2y1Q8dmNGJdtSvQkkO
ZaW3B8IVzywZ38xIh17yoFmuhj5tsZC3Oog/F3dhGAap0RrGtE8jSRFa4R97HvnZhzreo/+2YJVZ
ZnaEipHfgLFBoO4i7EDzs2GliGFX6sVWUZ81CTYWBbwpj4Tv7wW4Jt4jgY9frmuxeQSDzUKpTUQu
q0KFkmfj2jpf/huf6owCw6ZKU/+JXxg8VRDKOq0C4cv99BpN5/BOimp1BIYN3u2sG5BrsGTWeigq
IuF46/WrAKS9w9WI3Ls+RRSrZZmu2vnIgVEge/hKJmx71L+DcR5vxbRy6q2Or6U+9K3jIyrSVdsA
UHu7XqGxlD+LBFsygnnuNH6kKpybP1VO2vagrt3KYTGm9W0V1niu7hwWnwPZ5UuOPiO/zNPyzvS2
QEUkysSCR1sDGQQJBE+pSZW5Cu858vRg+sq+TIp9dQBt8EpBoajW1lE6sIAQDFeCdEhjP1cDgabg
hTcExUXtfYvGWFs0p22ydv64FoXoloqacadBOe7oIXps0XXFm3YFmZMZAYKmm3WGEBadA6vLFrxd
eBibkgVtsrE2GS5VY2wGk9uoJJyvFDrslKEq4txziy81kRpld689Dc/QMWHIrWsXqLtI8Qx6corX
5YWuUaMFrI1FR+1wv/MvllPRZcz4t9i4kYYGZvz4qLI+qhshz2lHzQIWry3G0F0VYb7l+vfs495b
+ubWHGa2opfyr1pZ9bO9V8lyU68qL6Kt7adv9oIJA+U3HC0uyjk+HTiwwfAsN/Ic/vXIJ8rwQUya
8GNxy3eVJ6XwF6WL0zRIBicrHAddZFPuaodWxHe3+gL5VDyIRcXOQNprBp70QUhjkH5LKFuRyMgY
dy8N8o/FJX2xSW0rhW5k5NCWr7PAgXnaiUf9uOTQj4Vqjqr3S2j9Xk8NV+atsnjOLh6mhRdgsfRz
VLKjPCgyDlKfakUBM/1tGaMUVBKRd5UKwiDnQa9JVDk7zyMtgKjxMKTzcSsL2X7iO0vb3n6BuAfh
CG6/EOljN478h/NtX7YFsqGMr27lNCu+6xODJhReRapUYKAa92q7So1YWlpgdygBLr7LzpjRtMBV
cvUrCJrY6vp4Gue/0/LBnR17Pr7GUmk+xyFaAcrkSTmGFlpfTkIKoY+N4jamA3GUkTMBVkXJ/S6H
eHuk3DH5lcUXjXffpPyOmQKoIIDD3BTOI2hpAtXwGvrS+93AzRDN/5CWAiNuVvPBqko2vO2vp7iJ
ERRciBGkyvZ6RNp+AeLJmBXXY1QIcNGQtrW6+3RefkD2driFafZK16DKZ5VwOzciPlMcGV9ar/Nv
8+5PpNru4KUlZAY7ZNIUW2+9OivAQUJx9tp/USGhaHt8aIq/llDOU3iZHZzt6M1LUM+lWPmeZ1PW
6k+FjO7MzAw4pUmaMQZ9F0RsGMdED8cxk+BHth125z9rjJjzKXS+ZmMH7o8qIltaaWhMRqXqb1y+
OTQmHtydjVPhxl5ev3ipVnnb8TBSicdPdMuLWnMTXIOFTtllVadx32yrYtVnkqbb7sf2VJoBneJz
1sy76t0M1pCFBxfNSPqV6FQYjVj/uBA5IwTGUnyU6y32MurOLf2o2ArKusvsa0uq0k2+B4c2uPAC
q2kPyXt4uR8PPiuROrDQtwTq6iVuH0tWMjbIvbG5KDZxSUBm8HAgONw84yBcWPwDCeEnyux2Vcat
biTvtEZHgU5poHkHTuKpk7DQ29DuM3r8lTJVlb9ZQx9uW14zINWFs2uyllt5a8K2B91AnxAuPQHp
FMdIYkpBh0XNswALvTUBbol2ndORphiD4gnOXAYYe2A9+7QpRR+6y/S4qMQlTBbMK/5isBKFFrHA
ta7T7bLGCLD8pV7aT419KoqiqqwYva6mJ4IgTiU3KrqDhohF2K0/OtAOf1vnFPo+aCjsXo24WW/z
f+VLyv45zGfCZzCje2E2ykwHVHBNzbs8+3ref+JNHfoCRE8D2+B+9UvZDVsEmS/4D/C2eGth6cA4
U0HlXxZlxIIoP5dJW8F5A3hQnQwoPCkf5eJBECF0+NnFveNJcSeDI/W+J1Il5SJi1rm9X30JyRYP
uB8O7U9xZW5cMWA1XaRqZvtIiled1Omf5KYMFyOckBUCvYsEYDL7C4+ccmoq2buz/qnFytGcy4DJ
ftuulG5VTC50qhAjRKGo1xotp/le4DABx32JlBMWHu7hgfSFE9OHva7vFgxLV6v8sPV9+FirZ4iZ
QFu1IeRuPBf9ezp0OJyTA+olgVq8R7Qeddyb29Sw6uAk0Kj0ys2c/BDhFJGwQgcFKddGzpo3X4UQ
fNrYQ1bXkwi4adwuTK5IcBp3xuSglscI67hPxynC3escDnZTaHCLeqh2R3tdQR5x1AHyNEmOCblJ
EWnsC8YgE59hQn5yGXMuygTazaYrDtQ1HKa0TeTfyOUsPJVQaJan8L87URUKezBky5ZrRMNfA5hR
1D3b1ySAl+gap+hYvE8w4jRgmL3YhIldN623UHxUZXsFmxQFdiWZkQBHB9zDqd+mXSIRJIzwgWDC
l8OgEoWKmNByy/g91uENDDTRd/CpI8y/o2RZwxxfYA4kOSK5PlQriPlxCyyo1GOFLb4WM02vgwq0
zohCvcbIyuMu0zzR3htruvx2u57mO+YUfMdfW9JYdS8eG7IJ5Z/EMiF3aU4ratSlJtjXIxvWbtgu
ac5Tr3TzHnaxpbEiiBM/hRuA+F88/b10+ANhibl1OY/5syIYaqKYcc4c1XpSd7yzK3L1U+OCP9CQ
/ZyoYD1IZkRU5hlfpdmH3NoCv1cQikXfQskwX3KUn0gyqx/EV98mW5X3cBKhm2rUcFr8BAmzFkt0
SYJfsp/LWJmqcuv5IhSTzfLbtXRBJGYGKZe6zV52OUoILB+ZCDwOMBuJjen/QH4udlggrcXwAA8g
pnQ3YbE8O+puN8z7a9e+sp1qwCn7GjsoY5Lf3DK3RjwKsg19OvKad7lvRub6BxAVwzIYtiR0eNfU
cnGGCe06Bfg/nDDT1FyKHgUYj58afuGWwqtF6GdzjVfIdwcd5PZlHMxoFoIi8QGqP7AaAHT7SZRl
EmV8gRETqXG+7u9frzhnDxopX9B/a9oOyn3AP5Rd13tnb8i2MDgi7ogcrQZpHi1EPebTgv8o42Uh
mzLaXOMGvk9DIQWL7v2YoUsGA907yQ2J8wr0QurNjqc8oUCW/NjIe8y+jaNAA6B/6X8/2e7AerFU
tcQEMizeKx3n/NgkviF6C+4RU4Ys0pkvsTS1m4ga3rTST5ZwpNo8bGRMpaj2wldpNs3HxkqFIJR9
ulmw7ewyP7ex8zAAVuRaxjMqw4vDxQhWJrvtC1v1sK4UP2m6hlNOah1Znc6sWRINBLCVn+vbUM7Y
esnk58vYzt5FvbxaTbsJ4jftaGkCUK3c/uS9nIlEY+uG6XUD4KuF1nDP17nA3xOrZFLZqqPKJV4e
8ZL7GBF4LbrulFQsLiVGA3/zh1z0s2h3nzP+ZRHtaqW5TAgS8DmNJI2By+raFhUuIOO5qqtgpJ5b
nwBH0IMeeBDl6FzuWHVtEQIptT3Pht0ue0tS47FxQgou1feaOzABL2n8J+jandpv0SN/D5O+9G67
sIfQh6duvVabJ2WhZX2gpwpYevn4AmgN35a7I2cUz4rjHCg0Vj1nWauM1gMYpfQi7BTZwemSjH/i
S4dPaOrqn0h7s3Dld8B1jzNUqpJclEFg4PRzM/IAgvCJpMW2cOpgCQ1fLRkXdO6le/mEW4jByw/O
pcT9hum9HcSjVmwquBmBB2KogH/1gvHMxm836k4WV4NOiFKa/X5tO+x/Mbjtznhr4dLlRuktjkhC
gZ+UWsx0Mj3phARhLigbHgGUXnZmGEQND4Q8WvMUhqrusUR/B6qT6W1D0VXXIDcHo7G1V6TRQzbg
NhT8rfFvmLR2XK6Sljq3QtoSUBnD7SxnE940luMmXgI5uDVQlwvP1dEnTNYNtuIKM6rcYR/dCm2M
6b8WOA0Y590diqbamO4hZGFz7MFDHpQ+DCxNrIFMBSkTKWfyDOwVwlqKC5JtBS7aFIrMHxqtoYzq
dtrgKLHDe+0cKu489719ynRDCkRNNGiv3X53lTAqJT0d+bCocjwwEsJFfUzXKXSGME7h2Iwxfdjx
+/aElXFhRDfKrpTy+tewkTx90GklpCz0M5xfItjRbyJdlY59KVX6IzNgc36JdQwH+w0HixgP1mCs
Mz4degTy9wfughad5xMUHSW0Izf10M5alFREfj8TOuT6FI1SlnelmdX906SUI4uqpWMchvrTYXek
z2xdtB+bhysCXvK/OTSK/Fo/Vm72pT8cg7Tkw2xxBI4SgqFEW1j2c1Qe6/T5T3NBACihffOIeqhF
4oVKVySYT7acyPALAlGGapwIZlKsbT1P1S7BMtMdIAwFGDAUe4iSHGQlrf1UtSTndy2eSXkgF92g
KWw+9oHb0YNPxQqHRIBxRP5soWHCOaEux5NacKHwxNJUA0sCV7hH0Q/kDYbI28j+JwHOvtNQ2idh
Jbk98OoutcJED47svq0K5tGQDIhEFspFAdRdYG2ULPIO69VxlkogHdjMFyc3dgkBYRh85ilnRMSE
as+jVbW8d8FI+LGltyZLiuwsu20klUea9DvuUslU1Srjtj2a99ZkVCsSWv92cnCfQOUCwbZeeNwN
tg8uOkj5cR2n0S/ViATrITH8wRfWf9VQNVQVWfaCJ+s/8b96C6V9BLd/7sFEErbPSDbGBPAvI2XI
qPpAzlDuH9kZT1s3RHSZGdvs6ED1lsTjBscLhi+iPZDH0mUjF8C4fPS5LFkSR+RMJldb07DwTH7k
hnz+CjuRP/+HUa/UqYZZ6++wyyKD0MNjmp3ZAbK0BL7xwLQuqGY+h7Bt+jwR1D1HBd6rJDSyy/Gt
jHdI+/xrCr1QtTci0+Y8OINWVf/bq/sVhzs07+rQjJYyP00VlbPBYiTaBURNgcmbZmQqHm8cqeyO
WUdHyao9pzmIgxhIuJIu5GqF698rSuThAolL2nIKSMNnLYfx4yP3PP6H6StfY4h767PRfRlPptB/
Hdlwp+DJ4JxqV30yXdNKnrUeKCT5Z3qGsuTMOU/ZIIk+KKCLJWGW6edZxtjWQqw1aDKJQu+xa8Eb
KKBAOdHUS0VXF+adWjWZy5rwtZbP/V7eMBQ9ZgWuWijnj3WEZRZklJw9hewuJMIMVXHSie4vmabb
Qiz90ASKLDtTifhR6ViB95v+qUhQh/VYWYeORKNa2oa3NtjMNlIPkHwtz/SuugwwC24fIkZJfVXf
P4lM6+ywmuHzz0mfZSZ9yIBvSiyyztEUUqMil47rHvGmNoIkICKIehA87zonT1xcqhm+jeN1HbUA
2W93fCjPckyperU7l/IQuzufNyqHAzZY0xBYTD2gNJdmSTdprRnAdMX3wytFID68BcfS4j1D0p06
xp8RwYInJQ26pJC0JQBFvZiz4e/6iMVh+lMnJyuKKy1HPN+mpn0dfuYEW9DU8qymZOYgX8MCDOml
leUL/00MycjMjuVPWc8Gjt7rsUkU02LlKc6x0PtO5Zh50YJbjp4/Ptuji4EjMTJb1Ge78MTV+E2f
0Whff8k+a6eZGjHKQCJJsk9vvQ9Up663L3j4DO94/LG8srHmDwItj/DlYS/TIMr3j+TolkACQGks
yvmMsqRAxrunyApO+RFhxXcvdKEkc36ALFI0JIQy7SRd8h/tccdr5XU5U/Fc5fDy3yscGaFmdE5s
Xt5ckFkrkKkg+M/YGrLwFqh3v9Mj27fiNtDicahE+yo4gkiuVduiK3aO8tKxsJamj6JzXEvCoKpz
xBiWGnOuAgFcZ+OYLtrPTDbc5t02N1JQb4/EEwDFNBQwMm39a6FjMkoPZ2A0vJrSy8BGx07yl5Ou
MPqjW1LVAdiFgeCEpXE8kHOb9KLBmKaIVPqLnEPLM6qOtA+Xd1sF4lBq9PB6Dy8JvtrVLSPplSnF
D9bCESXO7bvKhipIJP0X9mI7cyJEDqQTYxPA7U83DemYNtk9ae8znmrsldrviDhPWYej3BZ3Ob4i
RpUyYD8ybgJWp0Ve0hE9rqejr7CtiglXOL5b15ySSC0OxkbpXRDandL8ffdjhjNXz37qYa1HRuWw
bGE2KQ6/jYzf6m4R1TQldQQNT/ouqiaMGGaHaBKNwP8FHSSNlyzUB3DQyc54mEhtC2tivkMgfsJN
O+rmW1YkRTJe4QzTBLqhnB9iMb0XUIunq0R5NYkpXHkvRuDLTPc+sv4od03FcQRYMtoKBX2Gci/q
SK3qdnzxzomJw3vnCpYyAHONXSlvuI0J2vMjRVULqwcROEwdI2+DYdKu15enVAGTDgIjyS1bjr3g
v5d6Qjfs7aRC3KBZDOeU7/SKnxYMOsmTv+5vYvXFxxtwbSS7guPZrGftnmTZb55OuZTtTqBlbv9S
LEC0csAZeKpJyOh02CC86JTT2Cd3emF7el1Wd6evB4NQFVneZrVZo3PJzxDM8HtWsU4iKRwniu11
vu6Pur93VUOr7O4BbUF1tMPTimLjiwng0uuxDRa+4//2tL+zmZ8YGgAYh+cdc6pZAVH9DnZx6hBb
eo/530jmeD0jHI/p0C13j+DTvVoes21AZzAKj1UxTtJ+qUG7cG3vuWkUsG+DGw/52TUGCruAfnFc
XcBpe/hwuRweyLGbuCaZ8vOOi98q1UQYH+5BFyf5vpq6TAvJeeeKg/VcSoLCb6irAl7qpTc7iBdC
p0ePteDQOULlVofJxab1ZPpoXxs+Mlerzir/gbQKjImd2w5o41PmHXIz6/hd8qVhGQKzPL8D9O/l
rhuKhTry18tz42cvWkvrhaTmxVGiusFWU5RioNvHFEAIbralBm7z85+rqM0fek57CIJ1mIsyf+sg
9SAS7j7rnArgbQ+1FtQHnfr1oe3fNAB6YYLj+ppLKVBgdpoIdbei1BxSeP1LdzPUUhXXI270BQgj
ypp6hqEZOZrYnpj9s2hWNCH9ugh3vuzHqboIBZvVxM9isXjUoYb508ircrWN1ErZ2SttpeaiGw/c
jA0a9TntBq1tR4MBOMw250MLXIy3feg5IRB05/oqWIw+MADDPBViG3PI5H4ctxIYm8S0bK5RkVV9
UYaDl9fcuyC9aKrE+P++aFWwKkd8hYB3plKu1Elip+coBHz5ihk1k2Dmz4hLNnvpskYoCCvgesyT
zLdto0DPFkCAlG9vYeRVFPCNvVLQGSa4/XwmtKHjPHZ5RVK+x0IW/moJQpOnbNKCDPEMHi5wYAcm
U7qk3v1E5EXum8rRIdaJYZsYfgGbvjAidoQmGYSrX01Gez7T30EVLo1b0/DPymsLqx/XRpQ/SA+O
TQumwt3mGmL3SjWTUGpKT8KqVwyYI+aB3VDfyWrPwDTjSBVIRV8RmHnfga3OSwAZrgDYfs3bD/if
Ir6LnV0mhmr4iffBr71K2Hq9Wx4cHdyjUw6+fx1Bx/R+IAgBcFLQ+nECnD9ISZCCoCC4+RBMsJma
Kv+4kYnlXqdlfiYCqH0mPGB9sNqsjYX+brNjhefkteC4kTGnM9sbBdwt/VC7GDTRvyJq1NZGQghA
xfhyUcVZbzx2Q+iSTDk8KhP2Pj22EFy8f7TX7DGAWd3lvna5wTFrk91/nYWKn5IdyZ/h5inmZ/b7
1rblq5KbAbz50jnerLprOC8P9MwQy/JBfVoacVRY6CONH+l/ZLkuyAc+aCbkfpfShHGM3iDnMwz8
yFBADfQjDjlqt6vSnR9eaFWhwT8aALrEDladZGASe9uCLewl5ZLw4LsHdUHGYr8o7GW/At+q7XIv
SpYvUWK9abcySkXKsJKJJVzesqb9boGJ5EIn3MFJJmNeVNTQ8bfM6xjwKnanYZH4FkpbCnTAj76d
J0GKfBj9lxT2rrqFTtdvci5VMW+givLQkWxUkHvcPfKYpNYCOHvvmB6GDruAZFsGvZt9m0m2TQfB
OCEZp9TbuCG9gfazv0qiGzDeQKAKIYkm5NYLfIEGJpZqOOxDiyAWhdH4Qx91Vf80gG3vdLSqtRzN
AkpobDIYHV27rFeoRC2fb2fxMxgXptIs4HmifG0DTXsJlnLTPqXj7XADqmgGe59kS9AfDdaL5Iyu
4wpJL9c7waVto5FbYmO8u3VCn9/Gj4uUQUZ5EyANo8BDtpXLMVNzg/T/AgIRCZpCH0855XcUSedg
jtCdj7prMj3XzjlRVXV2lSzsiKMHDVC5ctXjyc4BDry6mqfqyT/ldQPAcuwE7gOtITvkoDER1HSx
w4NJzsNnVJGx8c5j6DNXEcgES9WcUTllez6Lcn46gFOrsrF6nmIZLifb5iY1eT/6CCwCpLwwO1aZ
l2pYELxebAn3/3/9+AEfqh2+tSdN3iM5y8FkYxUShn0JTs71CkMUd5XmvMJF4fL/6+2XhuXpS7r9
GK94YqZW22NWLu2RXz7OdzEDDaxmGJ5XX99o/TsxYSaSPpt6Pf0Ocu1hlsGCAIzJaZ3l+bEkaDot
w95wSK6bgdle/YPYin75b4Kp2w08XpY1rm4pff9/V9tirWs5vVh3sR3BzGPNifzLmw29fMVxmHXb
+b6skvrHle5PGwad9iCqAlRTyaxh0prFnYcOZJj64nS62oM7eP1Rqh9f5tR4f7NXEAsjV/7flH6O
NFXSg1mbACzU2mxKAywWpMjdeEsjsk32LEWI9z5MGyctHxSW2N9RTVXfeR1AZBhrcVE6x3YUpBOu
hbYdmipHlFp0BM+Cm4CXWB2KYOMwBfUKkv6gWmItXODM46Iqb6vCygo=
`protect end_protected
