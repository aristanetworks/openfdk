--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
PmZm3VZq29B/5ohpK74FfWjsDdC9uGszrqQIoH01LD8xdRNavF+8eCzQJL7XmPsUteDeAcwuxZno
keCa/DGXLxGHY/wTNvmF14Rgqozp5lA2/S7airvNVS70ebi3Od+vlNXEHmgDL3zYPQnlObGa4CVL
9Ihym9TO5rW28zFd8vcoxbWsGdBzIrYLItL9QJHGa/tEU3dgk59CXUYeUjiwnd4iU5nDkeeYczV+
mYRH1wzlaXBWKmOznH8fhWr7TqvgbzNBxyN04TpQDLJVa/s+Ap/3f4aebc8YmQFer6NGcJWPRzAs
i/74eTX3Gnvvv3aWXoub8qrP6guLZYZNN9YsXg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="HMadYH3ku/doCEmaLq28i7tf/l5yY5GCqBb9KJwbUzM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
qyICwCmiN4b1aYwTx4+RUZ1KLjZ+Syz7Mj3oLSkjt5QP29PSBvSvxd80/l+265IeB+Fhg2UuHbXe
hEj2CK2dzI4y4fLHvDb+Tj2VWBt8r6+emVRMtmzX3l6+/3blZ8JZKiBb6Gf7g0gj48jQu8MIdjlc
Fdb0qyJmUAI4IqsyMrevKjkWcz5qCa+cRbfcCvGjYEv0Q6dVhLngXPHyv8GrJn7dNduLLELZPq2i
PEjvhEXMlktU77vaGvJorf47N92/IQu9H2tAqdMe/90yU/lGV0TAq8oCd6RbbvdwTfWcaRJ34GDE
pQVC0o9SJhNOkrHhAWAM/2LKxkaHz4zavHGFZw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="dJedko74dMPGpuM8XTbz6PH7wJa/55d45Kofwlv79m0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 68896)
`protect data_block
G4TJtItVLFMFvwcKe5eXuno42eHCmbOXp31fQ4PNkWwFohnp+Fv7K0Isp/kQ0iqhnExJFVwkv3YM
bmJ1+cheSkfoRj/cRhaFiqrlvLVpNzDNvQ3oFAxgFvemyybvQZRqmtZTK8tculjGV1e7GlK9+6YI
2vMc0I9sNBrhmmBIEvN7s9rtDN0nsjW9TrgVlGc1i/+hx9OpKLDob+COjBA9TKKa0RN6af7DUCXs
dCDLfbdI7tyNC2sQNA/Tq4KM2BJkcIIwz12fWR6e+gpFf1H7xP95XqHDovvNf9VmfFGXhmD5Gf7V
N+yZepoCdViTpRGlVo5iOGbgIu2OPGBZGgbLr0rRXRb/Z44jFIEklDJUUSqI+f9Wmxza/qzStAvo
K586U+a+5rzGBBSx8GWZ3H5CzlZsDqDLxrgteWHzStUk5qverIhivqqAis6gKgPtjEPFLY8kVvVq
+EzQygNPycKrKAdbgyX8/fMb3EuKGHPvQMMfhBfW5a3Z2GioLKb5eKn7MtHJAX/+3CFtwfJ71qHQ
e64KfMKRiEOK6NyNBdIl+vJHPPGJO9o18GTDpdUlE4F2MjVPu68fd60TbrqTFNFHGUDmhaQoPbtl
z8YPuRx5qb4PBNX+7Z2SMjog9dTesphk7KZ8fRYGvqnisUogFfgtq76I9XCSkzxNwfOBAizjWw7C
6hg6AHatjORq4HaGHjcPzGvYmHP11a+N8miEnDLbQ6MKZu4M1Mcc1JyEOmDDtMxyY68lO8fR9lW1
9gl5Me1by+xJYaAJQfC1/wqkGqcGzn+DK21DI8S28PJ1dUqk1wC+f/BdwRYf1t/J2DrJtRTaHHL0
0p2ZhlkQB+3EaMj31C2Ttr/X6B1aTc6GhUSHZ8xMwVwT2DPeKISSH6iVz2e9GHObKUpXHQ6/t7/A
NVTMG84jJ2ALFLd7JTfJgHfVn0Pc2COLCPP+3IGwahZibWuiteszrgsGelO/mmjjLHR4qUnICSO0
OAcm4+PhCjdZt0HcnmlxrP7Uij/xuwULKHlPugnKRdyD86eOGONZrgol5Lv9R90skrkuXjKG+ml0
diAJmNHWZyXxHauQtNFAodv08Usk3ITlMC8kHA8I1jEsH2Uf49VAed9TDqiE5Hva5luRhIyFY9QH
evC+NKEk2JBZJ5BVPDp0XH9SWXZ4mBebKeO03ULXKnpmKTVFumg8g0ELsAvdMaxCQ+ffnotsB5QD
P3E8bVtiitNs3WH3Ymixy6LNtUSyKrFxD7jcCorh8aQG/6+zq/1yPT7rF/PoQAyMrOJRwZ4D2p8J
lOL3EphrCbPgpMgL277DPdnzKLSPvDs7dml1x3P0q3Oyljt4uKmGOQZh0Xm/W/677uvyWaFm3hP5
CyTOrPqmkh2OBjHlB15OZDiwlqdS6hUa5ht4iBZMwjrW87FLGDBADkV61L+KiUgtmljZ7t3ae3fK
P9QSlL8XrMVLl+4coPgUa1Ax5uRgLubiIJMy4fmFQWDAcQl6W7oSU3+MoxmCsSpGrVBVtXe68YNk
UXQMe+rDqto2aBS3Ln5XhgOXxSADVUPwi33PA3Mi/UUIrORpzoSVAVTwMz/hvRLmGvpr7Ayj9siL
hSlniiwcQrCOpOvlLTLj0Cg/0r5jV1F6iSv+kJHV6E1K7fj+lY+fa0uYzwfxEToNf8rEhN66PTCs
NgBdq0hh4Yhf3xtsKaE0+Mjm7YJ7Ju0EisnpSo1mbSnKU1h85dh8wjXHWrrhUCZNn46Fo4w0NRq9
e37jCMzM0E9ROoPZLQgqTd0qLh7CV9jJz7QtBZzQ8ctOy342jCJaGT1qETjkgrZWtSTCIHxF9Sdm
82Sw1QY559NQUOlyGgGHVcKEH03ioeKc8FU8joRd0NAv1w9Vl/nX1c8uOMbJRS5hAsItPsx55LtZ
ZWxVoCMDUPF1jjnwfus4F9SAxLfavBFmpClnVkuCvJG1k1yLXoAamsSC83hbZYDlb8s81LyJBG1r
98Jgt+6g2szE/gmLxXbptqAIURgK2mxGFAwxIlYLqqtRwxbhaTg02vFTc/9JiFIomdg6pIyDllWB
LnH0pqNs8S8JzlwsA+ugfHUByDwc4dA13Yj7Q2kVDgmGD+eAWreeXMCUiQEPOZaPCIKVHQZQUclS
peQLGTEsKWrNvAgCZlZ1x5+XG8pkA9msi5C3iXaKix+ZqYoPaq7IjayQIOdg9f8v4SAJWVyRYAKJ
tzcB9ArLBJc+t0ms2QhTpwMh91dBr9BhTZh3Z8Wzd4m3Yt6grlmJlxTD/vVhqykig0/DOu5tLds2
K2TVLM+r9vEHVmO5UuBEw4BdLk7hI5KBm27e8u5kE/Jf71bN2fRgi9GCfZP2xJLILRieLdIw8CUf
YZnqW0wg2mAziGWD7pWVXUEuPc22KL5AuwpUFWZHLywgT6yM//uUJEYFE5Ova3RS+6BGv4NQmLOe
sUcel+6vtffaUqLAmSWx0pUWeK/Y37drx+djJ5MPz9T4K7K+PpV22fzklqoIPbhTJBskCTh4dujM
xDUbJt6UvcXAfjMf71Jpxaud+dwvk1woTF7BU4Elj8GxcqL1w7DCRyOSfAYT0IbsfS8p+giKWVEg
XTLBrWXOi56MKmTuBsBpqqYmk+mtJZnelJCEt8pGkU3nT1YDNoETCLotL1mbgMxNpWQ2n/nvrfEJ
/Y8WdgBM+P5bpUYvExDTPz9frxzluIcc0CfkbtmGZ8+YNfWuomSzvAWDvRODvhOqXmdbNViF9NbH
Et/IPxZ0OkA0QKUMRjkVncTNA0LDaXRH5xBN24o/mWW1q1AmcLFoqaR6jbAmoz8JPGhtbI0HpmLL
/oyujTu+VFPMZZPHrhiOlb0Z6tA3/mljOfgpOzCKZva/31xlV4XL4IDkOcT+wFdJdNmMXsHEMV2H
eZD/cjgWH8r30MQZdLm7UyXIBPaxBKuSSETstB26gjPVbOvD5sgW1i34qxBtHU19suPimZQDsvlu
M8avvmt6nfU3hswTDs+14U1Q0pELcs55Ff+R4iMz5FzK5+h9dG4Ltz5Agna9otOpgoxNuso7aCkv
6C6iJ9w+7uh9xGRttpyelEDX5RBcVEEdTt86DMo003l02KCRinxRO/s+6QU/B2xHH59Pc1/k2XDb
dehV7CZCKwl+Xy5Opx4+Nf1sDjL4tdQahQzpLGzw0JNMv51cSaD2Bu5tdBu6B0tzIn5dSf5uWsr+
ogsKV0o1nhaUiq2gYDbs545r62x6381RbddmljPb1hGFw32l71IR0KlGHcRXT4b4UHrU2jI9AVkX
RRgx92pXRJxga+WhTNcezDJBYgkBFyBXSrjjZ8BxTZ8/jDPqM3ENiUkJbQ7mxPvyjw4QPDF+q9T7
U56u9a+qkurUIyeS8HOEhtsYlE4eElCGj8rGEdpAwD+2+aoPRANjmPP0qCs5BD/TI7BFrA+UuHxM
ACGdAn1+IKdpG8m6CQQ9yQvk5sgpJJ1zz8tp6H/zFLGrvPVPTQRjUIcEHVmWskNtrMzzWyXvSKDl
XQcqSzg++2HLHP5Jjgr7fYt1ZMmJgRzxIpTE2kWHQ4LIPsnaR98ESQSemNOe/snKKDyLjKINBGle
nE1mg0i7XjnurXFKL6wy8BldfMU3YMdORfutM4iDP2OXTUJ1fI6+EOnGxp3/NQPM/GBAp7bU+Gw8
Jqx57USJPfntnj67bvmLl6BfLzJ77FZh3dyvB9TLXRwSlhDJVHJkNY66qSKSeapD8l1xTMTjd76v
cgMfPfIlg6FP4SX//WwhWV4H2zZE9gfNFCbFxcXBDcrRFNyrTPl/I4UJFVokJxMftF/iWLTu7MMm
ayB0OQSuF5A8CjEcndSix7wjXO7IO5KzdAoFxPVlyAhvKJnb97s7B+MdgBac4RsTGE5cJf9N8q51
gjyDhc/kYRwb+zaxzCR5v8HR4H71W0NzKMUD5DRqX9iPQRnsBS7k6oI/lZm0DwcvZ92hPrs24NlB
gCFPqLWahgqvtXt1yG4eRlQAl4oqj/pgppIyBEVdyCeDJeAcu+eiLMfAChhM7ZtTSVwKNhZe5GNO
I/BD6YTnObTXn9QKTa1GyfOpxG1fHvZuC9Dm2gGUZp3AtW56oEcem+0OKjB4QEyGy4RKpk9FUCW/
prf72Uqe4HDLJ2DcRgzXp/7/4xD9INU44EdL/kfwzblLI3qFDLxIcafyqnMXc5F+caCRU1Dd1xs8
bbRgRLVRJlmGDNQnWkyfzdErb+7j7PQ3+wynpO0mG1rL3NzQfCR1W3AVjY7H3kN5DAkDZNZTM8BB
EHd5Tgjbtr3V1D6EHeL5X9PURWmvTcQGwAWM1TQ27SqcXVzbwsR4mudtO1XAyeNiWAK4msajITMr
vwvAGRXSnuXjAM5IpcjrOpnPUlm+ADi1l47VskUFrIcnHhjSezt77kEY3B3IeTn6Nueq5W3X/Lms
9xWXiZeZeIMiQscep0OMhh/x0iR+mbt0++lhpFW89MhRve+QXHFjnOIoWZfo+4hsy2RWbEq+OpkU
nQbp79//7Cf7XaPE3PDLbGvwaRsp886uhNm8OEOk05InyEba1+F9fyJCLHa6qIOIxfcSDtfNr7qd
HzSvxTJh4EJZEe8g6cgNo/iSzkpWklxdL/GSoVtEwY/xlnNhbeXPFqA1+3tSyZj68FqTOKoHvHF2
fy6RdXRu82RhNd059KADeHhe69onrQjIs1QG4xC+V837E7OAhRtg48KLQF7wXjEunvHyTg8zZWQO
rIjXtoulw0ZHmb1k5zdxxCGxlqD29JnWtto4VlxVPUin9Ta7HDb/Oyym68uwLD/j4WAYueU688OP
Wjjhr0Zl1kzxn34dAyMaa+huqkPFmsoG3nY0IPDQaN+0lmIIfL7uJ966ZDrDicvp7JEo9rqXWMaT
RSLf97wUxVMrVGka82BZHwm8kj73j86fKnle+1sN07Ky9tnFOtvuo/XPtCkyezVw/pirAu8ikwaC
aOzXtZKjq26ljkdS/IjT709nw3ZoWSycYvpIymhC5LUEgR7vpcro+clXBGeIeURJm+mz1DOnCvpM
8z2/gkcpLHZWJI1gputXTkhnnFU9Zyx1SDpC7uxUvNCo9zSSeFPKP1qKqwK+XxOHWYe2Xbkqqor1
Wkxdoby43bGce+jHp6R9uiLYMFBgGbJiJzgncHH6V+H3HSVwlp3h84O3qIkwWcwNqU+ySoiIYbYH
7wGdvNq47YxfyNl/bj1iPFtUypXp7pB2G3MoALvsNnke73/YtVNEfmLGm+6DLBqb/6W/QnRxuQ6j
itkyfe7h+Y0LvuMM3tPMV535VNXeHb5Xk9uIdeIInjYiCG5x5YI21rZThI6H24uDZI8ZoFVGAEyA
i2AHMC3r89yrT6UL57Vy0unWWj65ihfpRLWT2DDIvZriuF0rRF6RRNl2inFcazrvDcufIucvz8pZ
04/LUKa+qsjKjyhKDqkojNXygQNqaKm2dJ1HWVTi7W41D5Hi5AaHzrwu4x0hvH0ZENct3y63wp04
Gby8+0Pt1tvSf13A4Weachh1FU49Z4svOdJfHQLxS7Z1uiTFGK8nYHUSHiKsUvO7YV54qZh4dnN5
r0TIj8rLEBT4IJ+LEXuGbwU9dbbfiucl6drAVCc145LgudWE6TVSxZBiylAF9DuqZmD6+CVjqSQw
hD6bFL835tGQSPmN0CSGkXQUaC9MYM+nll4af+CsXvF3Yr9EHtcbvRVwjbUR8IGCFI4S92pJysHc
S/AzjsaFh2cv3q7LyCo0QBBymWi9mkn4niz1q/SF0asJvFlcebLf1hKfrDdMK8KoO1IjQ8isYpZ0
mUvNFLNmSATbDRvLGlqC3POdObODZVc0mBhLlYTrM+XzcrEahXapnqqEGtYmsLLKHfLMpw+Ysniq
JxmJZkEG9ZqaepNYVIzLCECIgHVEB4hlqd8FRQ24NeuSt3rMKiS78sarbV+r+GIBujjGl7BWSbeX
NfwsQkus9gcdhLnziM2kPqCYyrBExLb2MHhhGy4q/Omsbz5fCPZ8ykqtsGj7fstcxdvayXBeYwVA
X/wBJ42yKapPb4G2raDxRCDytaa+YYJFYUPi7qTuWyEzxJNmgBePpe8FGSQPgg3TQF27ahCjMqri
0s0jST53rsZO1vqJEmKnDTvkTRz4Ah37yCH8uVhImq3c9mnc5Nh11Yxj6mG2qfKoGMfXGwP/wt13
gbd2MvWT4XQoh4qQGvxC9kQq/PSsw+gJMVSMHw2P24/xASHzaBVLQizF5tuQ4HjmgA+zygPAF6Ha
fnx9dho6egUEPqG7HZ4jvDE7lJzLVAtaGyhhQEB8P2RarWce5E2p946lMhouLl/pHO3S1nPhOf15
7aQFYTkimvScb4udNv0Z40mYn9kA/jUrKqGu3Uiw6D8JJuv8VmMWaqNdnG6GQNZL/YnHduJRkbz6
z9eHGzVAOsETmwHlShWJEn9U7pLjaLl78PJYgWWF7tA8K0NgD9ZKeta3FQ/A058tloexidW2DvzM
4V1q+r1kTCouKGBQ/jnq7gUGifnWT1cRCL55SImNNCaIa8ah23WHONwVN+az1mD7WCZpiL/w+VcK
AEgzAyk3KSjWa19a5LCUa6rVJOWsuma4vRnmEkE+pKFN6lDSTENrktPFuyDPfm8YyhI8MK0XRzQh
1JLPYAFbgYYYkba7bEpCHF1wVwDt7fYpk1Cfi4yTR2LXvhJUT+tmLVFQTr5JcFzWQ1f/06TkmBbh
BocfgHNUbHCh6suMsi9NeO5g9aGzucdCT5KAq+PANa2RmH68d4p3nj1j27fDb83ZAyB74ET3hcgc
2l1c8NnLI8nU2H7NVyZiAOXz/eaOMU91kqDhYxHcGrLQzWKO3Enskn/sTwwYnmqxzRQ9NuJ79tgR
SGNU0g2M824HjBM/ZZzPF4uH2F1WIjT3+WPisHgnNGPx4NGwoAZBqA0Et6Ca9rqx6qZRlhiseB51
V9mK0DlnDYtL4F8RWRDVnuriv9CKl9cfyQ/06AYQXRfPtowkpVi7CA/CpG7iaI51e63V8Mw7oGTi
7vy+D/25Z6rWWWx3fMRmwKfcL/uqh8wsCrZqwiwZv6hd2/gsOAi0Ow79StMOh4avs8jxxZAL8/+G
pUG4AKfgxTNLP3b7RZwU2ZCHJVSKkjrfAcH3g97rmw9HE1tXNJaDhZEj9zvJn1Kp2i5KexiK/dhl
WmXTMnxfY7MMhEtEhcXizDtzsKe3wUcY9wmxfnAY6Ponjc15+KFlfq8R9XQV6UpjGFUUggCX3Iwv
Q4k2vFHETCzqQ4sBBbLaE7xJFdAeR9M2MSgWtpXYFSpB7W5dMy9IF/wLWPnaInaR9yqI61cE6rFH
StnEV3Xil20Md0bZIiD+/orxUgFLgEmmFg6+tYQOeTTNGFY+R2IY6YpKEwodTCMURgG6rqsdCE4T
cHqblizN6GeJizeBCkzKkm9aquSukGLUbFrmvSD+xXxvZV5/49JG5io/ebOQixMnlDUFSNsXsyPz
A+rJHHDvqghHUZlI0Pe+uc/GEbrLoLJDTho59PTG9PIyb4ztTDuu8jrn05MTGIhiHCi189I2M4Ko
xrrRuTATjGvh9mQpf/cBysrUKAp7if0U/6tiodNnif9NksMxp2xSPCqRYeXgOe0IdYZaBq9lybdC
TMQAtSWm2mLSK4nZlCZ0KMTrKD3k7u9OyEyuh7ZSJZkyQEWtta226kmXgsSKilxdV7OR9YRD4dW/
6DJ1UmTqnzEuj7IKV37dNqg0cW/aNVlnmSYhWuXGO9FUfUySQ3sNPZAWnKj4JTZxinahr4XC0NzT
YZTOL0w7b3AURjkI56+AscLejmthJwDVAtAScGrisFoTuf1bLwnSf4lxUyv/s2K0KHxmzCsXohgT
5/8tlNQuUmcgNhIuVCzR9ff7vfLLvPlaNU2ZN1GSm9xhVEUNizcYD+VymPhOM39cwnyttlEwe3uc
8qRWEg3JoKTxyhyNtjWEmhEbdCFOy/ZvSmk6y3Kfwc4ouA7Eta0NR+ClWe6+RONEGBQB9wRAeene
P3SKqCOMpLzby017ijSbpWaRd0mhbbyWrBeTnmaot+0/0Znl/u3BYGzEUn9SaZt3i2Z6tgrVJXS5
D5b1vNQ/g3R4r4JiSxjctjLJBldVoYwActbpg+VxjzKWaoBuhVagZ2CE/z2OyOPOw7Fwnb2x6ZuH
8rZnIjYeICdzx9Ycpj6VRrdv5zsrcnTRBIHvsbsVpZ7TX9FyPUYPda9235Q/6ZA4M5Vk40Sc91o6
ciatFGd78RekDC/Gd1N0oShwJG56Mi3D54ylT33/v5412MKQ4CE+dBHnyTn0o87P6GB+FpiqjRzB
s4U8qkAln48WrEgrnl37tciBnEEUbWqfoht+FzIR+pOJkRu2xCAsh7WOCLIKcJWxVmpVRoDK7b6W
G0+u3xXVls4J+EGfFzBMyyhTGZDJMP1wZX9DpjGOS9BOEXG8oV3J6xcVQlGFqgxy/TEfThiS41ql
t8O++sQ0Um1wpd1lUbWR/LgAHPWmm6HiapXx5obY+3VIwM8v+OJXi/2jCU/gMO1850xhFTl5Xv6x
zRZqVm8S9w7Lz82bUrhxSX1DxsAg+HRHkppSM0AaZ6JGjaX7WVYNrXFPSRfahfiy57Zd4hZZTe6n
Mf/fSZyZv8nyKeZsawOQHBfYtDrW3j+dWZdMp/2oo+Riu1tAOS+7JKELfP/fLhilaElJem4l3JJq
NmLNf37cLE6MzRKPIuO9606L25vUqitPts4Pz+RHh6V4zlHOstqPuHsXWsPhj5rYpngPvUEMGPw4
1qWeCq8NPG5/vxv8yr5wdEUhgo3lFHZDwZPa3aCfOy7+rUk/chLtS5Hmx7HV97Sa897bWcQZRl9I
NKKaHTHMvfCYnE9e3VYuSoI+j2c5/vw3APX04WmnIua0p6mq98fV4bRHgHGT89YfhLNmlCS73rW1
u3nOIssdt94NLTi56INBLL6NU8BMFsOm8xRyd+L4WSqb4fIOtaffROOIj3g//b+Lzp1PW5ypRIfY
x2c9MU8K8c3WgaxrDk/IfWGZg/JYl+/AkGv5fXUiWWBTg7T3nlDHvaWY7OCe2BYqc9vNOKnd178B
f6Tuo84xgUvTdT66xqk00+AVCtYG9gbItQ28brAJu6xscOPrC9FheuWHvoq4FQbmyjdCUG9wgFWs
tyrMtGUgyxkY/Xm/yAn9tsKMIyYaEE8ansPDOLkk3qPUq7SDKu7Ue9BMoXUTjJODlu3HPDxxe9eY
xNHV/OPSUTqp/v1ngw3ZzRv6he41VC02iMdHIdNetZZ73CDYLXBSfWIdU6drfJYD2nkjo5xGxX94
VYp+rV8lmtqRz01a5FSKEJ7dD6+Z7GvgtZV0mzxJEyrZRMznob8ZHjAZhIqkPMY3JuT1Pmi7hkiT
3QC2Gi6ltJM5APUtdgQc0tp64Wm4HaOFJ5UqFLJqLPI79X5uhUO1itRaJFBCJtNcH7s72+CveijU
29JPNWiYFwJf5bpr1lbFWIhw6sA5PE/Emik51UtzVC+DdbUx8HpI14K68LcWDrTtUJMv51YyGAHn
gKkjx+jjqDk4a7nGOfAx7eEPIByYAhVUPm8Es69hbukkJwI/pANkuYtS2U0AsbJLPlNur/7c3zYy
TQ0/WPc97wuj45M/gu8fFI2PqC6+D9yASFZOUYzro1AAZrkEMrcP4Wme3HjGlYuExB8KG4M6gFOt
NP1Qz40jf7AehOYM8BWGMmLOWO/dcB6kpGdh4TQASdqDPDxcM6C7hg7ZTio1+EUFtHnCY4PIs8sQ
+BKN8ro39x9DDAMT1mIEH05NPSInUEfmmz2qKXatQXQgCUGE6b3uOTTVRRcG7KAYlqVdruDfKh/K
Vpuj9CpDrjtAceSkQ3+64df2xit0NMRsBOy8v6mt1FCE+swaG3iJ8CCx8aNVNVGkXCH/a1cD4ygB
K0zzuGVXN7bIhdbTs8Ao8U78SdtCCa3e32GYjFWrwjx2iRITtlFgxgQLAQx5Ghvrk7bSUb42KQcK
N/w5eT5gIAqLpngx5khwFZQJp9y+QW2fqDcb9sV2BmRGODhs6egFmbJiJRgnpTLmCEb074eFCTK7
CU7LWeWEQZHh2/Dc8zCn0DN7NhTH0krRPV7M5BAsSBkNQ2rUWiwFsr4HCkj707A1wjfn0AIyMum2
JXbwpTu7TEC41mPYk1SB00bWQrK5nBnaAHAFhRPTUIjrRe3KD4XQxVwMhd93KofU+MwY/mlNe5uq
uQfj5NjPqbsU3E8rNAwI7JBzIb2ho7M8XRk0OpjxG+tEqhRPxmEQaHTE2rNT7s6Q/39ufTFuZnHw
xQe4JryM+J9p53psTY3kUtpMSedHl2VeOwxUaQQB514bqIRZGnB/5G3tTPYgy8AcMYAdvMoiCgy0
1uNzwaodtxu2TYq4lBpbMTxJ7KyBXV7e3DWS6QibCf2T/bN93sVlTqRrqr6s70BvJUzqrgUNOoMV
SwfQabH0jW2U8Eut9byfvuN5N0lCUBL0yqKRXYiRWfVRvvQ/V3fW5Lo7jduW0Vy1Pj0/askPZgqv
otsLN82n8Dnu9EpVF8uPUb4663lfwgS4Toyd2RiFwap0KX3EpAd15o9O5mb99l8IuWWNRqFcBvoG
xHKlSX5Lj+PasNZhJbtUG4Fbsgh6KwLcvPHExVBr6TFKbD4mWzypURbzUIyRY5QRm2fvgTEI9lLt
RRLs0JRledGx1S/DbcaquNKst8sYqghMhpVPPsVOGLn9+GNOX+tXzX588lYuyOhlF95/Nx33y6tC
2GcJypwmj7I7ScuM9AzEVhBuYgMQC4OCT+kugdVtpOdAU89uaEjsXaPFxZ9I+G+c6x4SPUK/+9Go
YTEedVlY08Bhhix9qN/6THNEXVHDxy5hWqMm/WYzWJ0oGlSqicdBiIqtuAY1SP9SiJUZfrdXUxah
3rc5vHsqm/+i+NP0KooutdL74HaBAIkndg8AqqfTUqYetRdwS9rESSKcxgTQlEBRVTj2czqVFvoq
PfKopCScE+L6hzdi+iv6DI3qopXTK+Xf2aVC8BCh2JAqX+AbwhVpMJKs1B5642lOuhbiV/xoAtW3
2AKy9j4zGUJ6yc7pVrsQK8nYlVD09xdPkSpcwARDQTsFw456thX/VkqZ3ldO0jF19zXarA4ifq/8
UYlcR+EZFHFwnGZ3jpQfo14qt0Yga3TrmMdzFXJdbAusLyN4swndgWnSo2GR51DI2ozitrOf+L5K
2FIwnnEkWqcjP1JVq7wV/wX54naGTFyVhtCo2jXFMGhJCdYskHoRK/yXc45rn65Cyur4qEdVFDzd
pcMbZK2zj2sE9pMPnjyaCcCr4l3VENRp0/tQ/JxONivRAbupT5ECsgrNWZla7Ut9+HzGEkUwk6gs
kEfjmt9aIrDOL6BTqFmW/RYlRCsTceb7xUBX74oSeQvhuao+xZg97wb/3W29zb+U3+5DpuV8DFQH
TskXesR7DoVQcM/VtSBWaayYRJxwZGUb21DqcXS4w4ylXgnB5jqS9Ce9HhzSpA1pu+4gJ4gKA4NA
IcKLaKI7hNb+imi2uysPxLOPhUvbV0eudqGscHav+scFtNSBJn77YcAoNBvo6aTTpAc0lZO6F+h+
qEQ4BVHyXJkRTShXNoX4aDuU2uAXBAy1YE/aSQ6zlVE+/XBviPLG/FC8C6MbAp7EQ8XbbH5qF26p
C3J65DUqhwkDR4pZsqj/cVEaAta0ciCGXIVjYdmCOx0KrhXCrBoU0qG/sUoLyurclE9f+1o+ohXH
f72/dM0wTfO6mlX7zysoBc9qP+Su8Prx1si2o5oKsiJA/tT+29sBlAdQecVeer5F8GvyLc9n2M1T
HCKdES7pv1CV4HZWnGmsVpTTwEmq/OqaomwrJcBmB2/qqtzaJfHbQakdajhB76yt0U7RcisuT8os
R124Ei4svUnCQmncSUTyh0CcZ0zDWOyuboU0FR4hnVuydyiCupWI5EErI8NxyDkFQatrSfV1KcMl
DDcxNO9qbO4WntkxV/8ZCNty0iLw95UDVEwANjFUUZWMMPjias0ubPYPzV49wThD1kX0Pz4X+chr
J+eQXjwcGiehvcz8Bika+cBxgRN2Hx4lL2LZEPuFDPGvh/eLfQNzQkey6+r/jCfICHH8XeIUUcSy
hAsk6QG5vJ4Ym/PpuSPk06QSVUlc2ee3zLI2nKw7PzOqmQbNQUyghgYa68Old/stKGxPCU2ARcio
fzVetzGcbEyQXvZWR2himBqoy8dmAtWQ1XFvmeIF7iiT2WPugME0sCwumV84YheSlksfULjxNItE
bsNe9dCz5GmtvzAEHOpSWdOU7vtyagGGo1KWwJ3ZoWlbbpR/23U10TY9zBGFzFRSEVLwycTh7oTz
HnuqQ4Nn0k5BOJ5P1uOPdcom8JIqHZsQm9k2bDfnY4iRkSgXjQ8MU2RRz+uZ78JpN+3wIGcmmChX
h3FT1t5XL3k006I0Fcgjji1f4aeEgCOHRlDGY9pEIlYYXaiOLavVQ7qR+FPzMepVuDE/gCUd6ZqP
i59kgvtY6o+/1iYsc/Y3ltuScOg0mvsV3Axb1acrBCLtFetpFVonaoBb4fs6MqeKjlzkX1rKPBJV
0ExumC3/6n8Op5rTmlqhuuWkbyG1T6v4UarMNtmZUD+HKnfIxy2/tBAcCywqxhq6/76R9fMPypcV
MvTHjgArqKZ+C8QU4Z71CaVPoDmLRqc7gAluuGMIHKGHNp8U81UqUBD+pW0OefQuN0WxksOfi5qd
W2IIdn8fWDd82CvuJgu/Yshjad/DwdDv+yonVeaC1Bnrj/8aSoho8Gq/ENPU89ZGu5TUnctEwwXc
N9xtqdAX+GgO9IvUDfrGd4zgT4DYhUaHT61u7SToLzrT0SmzLhGqQWCMf5rEDS2MvZm4GuKUKaCu
irUNjH4Ld5fxoATlQ+88+uuMBehzU8S+nRRLaatqe6XInlK+rJ4qa7rhZKRZD9k51Osb56G7U6GG
GEk7UE3PrEgJPBwf/tSar0m37UqZeUeB0URRvvtyrqlS50MT2kTDJs+WjcuvhaqJV8++NwzwvslK
v8lf9tH2W5DwRwSuGN2OrTVtGZQFwOtkXb6agpAZwJyevLJa0g6X/1V4FkhTv34IffvuBijmy4jP
KGJMyp4S3x9a7g+PwcNeG7FB1Fd3xfNFuVPGiQBOwcVKtcNebgx/hbEjgbUy8WUZVu5OD1zT4VmQ
o4bhjCXXJLYiKswKket5sVGO2NpmCGFMpsoIgsIabQtqVjyAYU+We/zbpqyvf8QpBn9m+0RkHiZT
NEDR1nOASS/SwaqeQL+Ow5ysKlirJWyIbWAVbMqf0jqUEFpd5ADP7s8tKjLnScoONhZsIiPN+Z18
3LeI/EngnuN7kucYm4KAcnPk1sv68hTwTIqLPIPL9fvvAJc1CMNk+tGUjGkGh26x8SYsYeBPhawX
c9KNYonR6gBKSLQggI1q8VJn3zHRCHVeNa1jqXr9LVf89eIm3xvCudo8op4Gh5hHqXmCRVJ0fuLR
wa+fkUQSK53NnOjcfC/6MPW6dGVEFoLhhh8Si4h1wuLcscHNRPWAUnQ9i8hRgjxxs7hNrm49weVR
3snFMA4RsYI3frg1H7AMHmmWiPtRK5NOwRXjiuADUPO6HrtCqtywCuPFWMk1Ho7v4g7/mVfoPPko
ojRysTZPnzQmW/ORZm4u2BkCYVqv3x1tPbDLdZDnMwt2bIWIUnnlVEkKBdkqV3D0Xi6suEHjtdL4
7DkQiW/UoRJFpE0pjZrdmKGpyLAu/MiaYegy/pmsXh7B6JXfUFZBuu9R4rJeDhh8xlJ0CfbxpFPx
Q94wdgxV+3benazSU5CeXVBiqLKSrXVP0QwSH1BOZNVl2wm8c74eubzNJ3HKp97CNgy+rmkDkdub
5Ml4LGr272U8s/7I9PPqqpaq07nG4d7Dz5O12Sk7h1i/3ygI5d8pRsOibh6xaa13eEZQK1SuVe2u
OqNPOrFS1fEGd3piIqjN6B+Oos/nZO7XCleNBphJZAWX9c+pmfiNiVAgTNCMXF+l3NRNZMXGyrtd
uLDzG1NxEMc4pXSzasZ5Jw3ZmILCeW3GaqYXyuQCF/gyOONQY7BLLa9r4NVGnzHaUvyC1rASVtiX
1XfIycOYzHKr/AALrpaaYz5m0VnrfgcNG+TNzr6watzNXwzY+sk7ZRAHeojze5VsI5dcyuBgDUMo
gKDREU6zLQGHhx5U5fV7oaIF3UAxy7YVAGLg1FHyDMkdMaEQASRR6w0KKdzgRjNqnyjGx4Uw9PYu
fSfhMAmpXz/0KXl7oeq1nViN89kFqvHjaL9LpQhyhJlfJc2n0aynwDKLfuwaC6ioAs22tDiE5DuY
6r1RFSl7WJv7lziFEjDNzLX2C9kxAe9oQ2ejXauZghxdRMgCLALG3iVzGySqvOqz8fqEALU/cZqw
Z3+ykX4ZQzESCd6Nuf7K2bQydKG/MiyettXqSvgG34p3Rb9fvKNJ44fz2VN3uqYcmWa911Ou755r
3Ga4Ixm9JaaBt+x2wmitb4QJiizz3dgq0Ys2/LOzwUr8qdHa7B4fsYqKSo7hHwcWRlYV14BWZWB/
ryEiP0bvORmG8GCZlrlUx7futccfe30YSLut+ZWaFS5XNHQwau+hrCUtJxrHGQR9M4s27m/lDsl4
rTAnOuvECRW1Fg4ptrnC3zI3esvPuW5f3C77evl5znu41rIPFXcbXlddasCbpWpfRcyO6wp0npro
w/X2hu0YuYUlapxGPpRsS2SC+po98fTeynpInLX2azBVWX3bwnIHgEzof/KVb6oyIoxpYiWnQ5hN
UyWtWV9W9dR9QMmpThmEAbVGzFr+eMtIL8I3lQJ06e3QuPXclzNYyAtS0mQC/vz+gyhcPzpiZ0Bj
YV+g3om2T7HaBUmnXJ4MMLaor5Fl8pNWAcfYRGuElN716IVEPcLrHi2gKhhrNYEMHDVnjswjAHpy
Rfrn8nIdYhh8Spm6MKxRXyRKCXmRVl1TlgM46uHQZvTiCzp6o7s2U2o4KnMDBMk848WZ9XmWNCVX
t6EAwirvkPWQMFczXjsmMLpwy4bz2ifWnJ0mli50qL2/y+sqVY0ilPkY640DpT7CFjT/yiDgsd5K
8T3NOQj6gMhM35xVtUqDZhSRizQ/30nED6v7f9GBUcy3PEQk2zhqRptorCU5NOiTcqEo/EpsSkPl
ZPVdxD3JDnsJ1OcISQPssy8S1jqfJzz9P/1eRn9yrhaI4AtAx3dPsMe6/J3a6W9ZgutqUyjHpl8Q
shz9jRfyuLhf/iNrXoUzBacUIZKft5LacS9wy0PWI537TdQS/Hvh38LFzMYiyPhO7L/ntUIEuW/r
TPHmIlUhmYOKydhnRM3hT2A9HKcy73x7ijyMvGIsFdyZK04fBNIC/ZOzxsJmlagFa8VmNH9Li/+3
YWxOsaTObM8RIDsMMiayv7O8TZA04h/6LJTR0awULy9VJ2SKEgA168cr35fX8LdGK2+Apo8x5Ntp
X7hmOMBmKw8ar4UYwKUT7Lps66+FGkwzZQAr7EgBYM0raDg1kDbi7hc4gRmU/i6Wt1DjRcz8+5Hn
OJg8vD+mjRjlgKx/KSuROcGuvbY7/k0OGJkAATqI3dIezOBg8PlTkBbHRX7bVu/MLDAwg/MRpFwS
0p5rlADG1Va3I7lR3ZEFbBC3ul059lFUZhD9Tnf9yie8tMm7wJC5CWq3ZnvsE2tK1Z+VbD4GQ4Jn
o9u9BgDCPywMLY4yvQuXvYLrS601oERQNXzIpjb7qmFRFMogto9276kj5B6kTmlkfAZy4oUYkBws
OieAUTrK7SYlUXm/LB3OgWuXhiN7RVNt1GTYv1FpHnCM7X5BTkl1d2Ihl7UMlvGQGk2h0vISLSFf
XCrDkSm0j2oYjSFJEds+OcS3am8r3hrrnF4LTPDTF28mDTF98munFjF/kLlc7Y9F/I8gAlNPxfkL
mRkBCcJmm/dN7Jv0bEA0/ily8DCpA1alOYVHcCfpMuZCYYebb2VgulFBMId04JZ+z+d2Nr7vq0m9
TYfFegaFuh/KgcZP7lYIW4UeWatqJNisuEpGtVxuha4iYKcIjFeHkhN6QuFrV77lddsNVM5wrL9U
FPIR2gBrQ62c42MUo+hKR+3zMNiscAyIBrh1jpNqbRs7L/ZudhHHODx8FnBj5hYPl433YWW6jOC/
pcPz3M7YQkvsH7aApVtXEj4p7P6ibtQacsQFpCkiXtllUlK1XYX+FnNm0eso1NsyV74hNUMFOrv1
aUaCoXdo60uZkoI1jn8/x9UzEV0W0GVcpnBdQDz7DMpDWEcR3r1XwmF7AVY7ZQS+dZE1WvlJwviC
8+FiBq3ePouJH/qFdZ+ptKxKdFYJ2Q95bzW04zfGYFInvv98m6g2Z21DOtMLcbpDyPjit0/MCQCe
ITwMNaN2urNPdDrNXj9xo6qMttbLvBReH4j4aCoB5guGbqAyXnpuLzIcj/uxJ8egcoSZx93c0glY
kpHmHNv5ojb9AiiGpa5pxZGGhcS6EkGRY4kl9oX6/BjRfEYm2eloTbhD9V9nFcS/uUXzBQ7WojcI
ZK1gqquo/VV9hvoz4z7SkOOOxGHuOrLin8CosW+QEaNyrltwk56XDyLS2YMEDkLMUV8CCH8TH9iq
ukF90HRRqyxK9Ml8DOKiJx8qevynWYTz7agvcjfWlygTie+UUhF9Om9JYn2A+y8PkW1QpUwaCs1W
JnezC7Zl7wrJr49/jGSx2gHHY+XJzizImq3jND5FYaKfdzdGZhiU3DfIONhbyvDupdhRmXfcIGAj
pNQ/K2o00ivYQTxps8UToopEM85SyFFSoetA9Zamg98sFJWqZ837hDsO230dNSMYHKYD2Pom1KhH
LGmPxz+6TGvHY/SDjkbgatcObflywPcGGrZxQ6sttTPMrquzSTi/yQi8OaK6rxN72p3cT8SXjTOA
PJ86UD+eNMzZqhV81x5sY+WHAM/CReMN7xhQNdll8UL2HdyZgNrzaIReg9AzMD0hwYVDJkCGV92B
VBJRnAvVvR4W7jIN2l/wJ107EHdvu71ZDRx3Ad6ce0oIe6QGMDE5kj5wBSMeCGaaXrTISxGliZ/Q
mSpeenWQpW7zJ40psNi4pXc0vGot0Rl5NmUKgPwrATGLqSBeUANaHxk5QovVspifUrC80o3XBCKY
uRj2O7rh781vvNxnu5Vc/DTUfiOEPsgiibyaUmFubnWsp8iKHvKeLSGUjE3CvDYVRd81c4V2MnHr
DNBz4Xki9qFQcbG0QHODNq7PvRGL7TX+nqaEWLr6vI3KrbtNeRlpHMXvPqx1Du7pneZYuB8FIW2Z
ixMwha5vqDKsBLItl6/bCHuAmlEX+2fTTE4wd0IASilWmd9sidip0RkxcXnBbflbduy2rp9T5lW/
qTc6bxBiAHWDUazVvesVD5uyu64MJ4a3s6OFJ+Rk6f1fpQED84NSwLklzaAHC3Wz7/aQCEX5mp9O
NG3mWafKfv7jhkpFqYDyde/wkWDNyGKYmSpuBx69qgpwsgF7XDV/YtbOttk+tF58UMhUCvL96GRR
lMTCB/ZlUgOfI2iUgwi/8Xk7YNJ/B7cXgiuAjk7GIY4BytLlrgxDy1LsCgkrWmdweiOZQi4/xtLa
u5P8k3y2Zf9OZNt+qwmtCMD0DllmSQNb7VT0pbfpOTHmKBQZ1t4NXSZlBQsdaOSQ35Hc4gGbOV4e
djv3QokWb2PMCfKUfU7Xz/D/KjUavEujg566XkB67vGFPaC2NNEqbJQw65U3w9kCcmvqomaZU6TJ
h01s7pRB32esT2Rt1LyVv9CCGoR5p+v8aoMQmNPjWi+jCUP8UJpNyYVnYKTzarEUvOH9vjuSHtJ1
0cc/8WcuSDL4hpvwEqmhNjFG1QQy16CNfuVBWa6GAAiuaufyYG1huZ22bbA5Kcg/OadiCXdjOcVx
MXJ+S8wEtQmWPOD1nXBPGu4ul0v6BLEss0Z+m0fySS+tXgrIHpx/KhgqFX1kfT1PDDKbj30VuOQB
P4jg8EoEikislXii0jGfe5fCz8oS+vzsz6GoQjOYhB6D+0AGZOUZIGeKpkgsS0Yx01hAGBIsF3ka
30vW92M7gzs4lq30Ss/biyOS7UY8eCvBW/pKmRIbS0rC6r/X1U/vKs7iQ+S5Wy3HW8Bg6+vGOg3d
/6JF68A1m9PwMOtL+lXIwbDhkSnYgAOiqq3H+CWvd4laxZ33wvQtqT0xkveQQ+oXvR6VDlbTWx87
xc+tU5SL6KXV0UQz67iiMBOMT1OU10nD1lMY5YTTDprJyrdSozfaEPy35X0I2aiAP9G6oU7Lat30
ocCx3/cCEGBMsy91/v7eGVkh9Zs8A8b8Z6DgK00Be58CIQaNMlw3TTp4+9tu4Tec8jHcyguzjGTk
ZmnG8Uuxv09UzBLlq6Oq6EnPIzdPbsWFNqbZI9VG9AkNd6Z9rRs199yGR9hEmOx0WAojtzFEE2nq
QEVCj+VcYE9KLn4qwXGhTra/ojo5xc13uU38yeo1UcF3xaPIoQqwPlGDCOVT+usLVFsoaSTxulNO
7PCQtCZIt4LHGqLMBB+T2qo3RdCubN3YnG1LB7qaPkvFNcgu81GymD8fceUhid4Ju34elCSXNki0
tUv4/LuHDDU/ni/7g4BvTkarlIEctpzk7axF6LdKiTkm0jpfN2O0qLDYza9tOf95sR2g1/QS/TRD
JckYXba6BpmQH1XYMbCY55bLiHKcNUOM0Fj/CjRMzjzI9n1Bdidb1Z02Xq2a0AwtcnJiXhJtLqJ8
BVlgLW1P1rmc6oZjpRLjMsojfKvgHZ/N4W/f7J7hitL7Ctrl+QM3sHIlyYxl02npkyigZFBCzT0u
bq21SeUtOz/WFOssLCubVyxvQYwn7hBDsbXZDvrDvvaRzU/le36ZaW5og/XEN7juISSkh7g8q6Ex
olJYweXVbB2/Vfeti//IZXOXAixygo2EZXBswsqPe8CAViIHMZ4We1XGnU6qgGGNdhm1OxfvSzk7
ODjViNpk5bC1E6ht9RTANy9qndbiSavqiN73cCYDXiTIZEGgmf66qo1vEJjaBExyLAua/o7etMAB
mF1v+BIA1SqgHeevsNoZKp8iFSk1NpV2XcxtptBytm9kaqp9xYAMVoFNA7RH+pCzVH86ujiXjOl7
xSOaCl/VDRGvzaAD7XUOiNQSO+Pg5QCIfxzRk+H76TAotUVhvBq6FBRY7O+L4KH6gMbMM1IfXk9f
y1KPY4Ms29XvRCVEwCfWW2AbXqZjb2HxVmq3cXXHhAR45HRTjevxOIOlkIqxitH7LIhmplOofyzq
3OUZrjB6gXxdMd47hLkHUknDQXxkGkLI6KR3601FoHUIiWXXR2R1nDxpDMeBLDpZY2B5ckwZU8+q
Mije2ynLO43LdS9xV96AuNjTnc6ZDUUEOcvckc4ohRisc84aLSdMLGK1NrjrcsLSIbyx10rmYN1K
tFlpWJy4BJSJaZvlh5rYXjwHR+YY1i5coYLVCVxMOrRdErVZ4VMcALycmCal/iqKs9NitOscXe8H
sitXd0ss3+Sc0YxhQhXhTaqt5ss28RBrFIOr1uL1KQnsdFdcDPkh8X1vi6JerwUFOyMK7qP9NExT
EJtw92IGYkquOaqkwsdIzGgxI7lmV0EoeEl2xL9n52MWuIWj0410MFtIixIQ3GBVfclbNP2f3J0v
yOqo5F5HMbGIdmNhLZCnHP862RYqbj5hfVSIYKEYvdyvGzfFAMfhi2SFhq9T3U4IhMyf0vVWpWsw
QjbGDLO20JrQLxpQsv7el4uu/Zc9pQIXljeAOp7Nd9m3IgX673WSRBj3RWCkEwH7HPzSAgM7NSx6
fi9f0/zGvI3ickglawtJiJqSxoMuemGV+hgQAxd+QW1xE6b8kTZFKfbGWD3ElgoUp/6nzbnlnu/f
mO45nm2VfMQNLRtog744+q5aHgKOY72kbqHnGY0drVx2JKdDh6LXJgJLkyUMTgjWdD8CuVqsAwKK
GSSTDr+aq+5DrYtmAvbyNoL8jMcCqEiDDV9/621zxkLt1NXdqfN7hXyUh2IcyX2KLE7RnttBiJSR
/j7QMLKg6R9lJDlLUYGHYHzNOwK9Lj+ldZdU8wFC6DBFA1iT3JlvAmyQXyf6fgSxJoLnqNogO/du
WigFKlArM5ErJw5i7gZj+3r1M3/Y0LOEkjnhjg0K4Atxv2S/H5+2oFHbar+AXhdNL50JC9CgrnS3
qwMlJk4n7rLXDKRCTjHaqvVRp/d+vz/pA2AAvQIVCMrILNf4gaKZb9smmx0GMb//rmAAJyjHots7
O34/8/0MP7S1mWcMN7aUjIdXXWzsm5EMQEccXWRc2vMGAkgAnGVahZYxrBTLa4SRdCGD3Xx5f2F3
Ijyfsg4d9bRp4jjfl3MeedGxsEKKhR5K9LfVpuxjMs9G3T+4wfhI72kdmzBx4oMHIYT+WQs9FaYx
tPpovrdxGTSFH774gBn14rVbnmRuSPCv7gk+ea3b79OzydS7ZJQplSAJFuCiXvbnONEt4Fx7cU/9
5obdT6Ql+56a2Foq+aNoylqaoMysjmyxn9ON8QpEAyzgWreXJ79vyXlBYGl/oKfgzfnu/lm8rDLd
8YA+XQQ07YT8HWvmkk8wGw74mlLNb20a1d5dwInWtsgc5NmnvbzmFobt6CEVrOIeyOfs4Lf+eJ+7
AlBtkwxpWDoJcnE2fLpquJeZhMcFg2Dz01A5aLz5aPGxbJYBL9jbIJUfsBoUB0R5mQBWA6E2749U
kw68LL5aQ04ipUwb1oFyaWj6nwUiEvrOgC+Iun9Bvb7VZcubEDeKxyEMXRdwIbDKcK+H2EXRTW/n
ax2FreZqXIu1NOZqPJOsKgNZMebPJC2MFckFHl688X0oMvYSqeD2ow+2GtuSCWgdLYMmXmkK89BB
ARdywxJ6xVZTHxd3lPR9MQEKjpq1/gCQVWgb9JPgnTiFbQYqhSkgmr3mDQSlIOSzx7YHmTeIjaUu
fFlHUQSPCqKgmUxwU0hYMOo51j3Lib42hTb8MP30xiCm7F4nNjOlY7bEYNvgy7iY2nenEDjFEetF
1n9ugXdOyO0eK2fXw4XMa0j9tHjrv3TXo2QwkUpzHMgGON/nDhrL1BpYzgzvvcby0LEN70wxEDBX
gZwgiOsKAFxx3FqNsYVcM260n1QyQk2uD8bQvAKQ3LhOzOoMamtgR3PBRUC2LMTdE35p8qpWVcWr
kpeH4Psf9pBKOROadJcOwENassqe1XBULwarh+3YJ/OS/Xj2cspw2ZqqyZCS5dCHyeyLtkmKvOPy
BhlVfDnj/AAExAd5tgEPjQWxpN45XmHCGIRbCwdKeOvMlEQD00VhrZQMvlLsCO2E+Q3bJ/z28Htj
pX4jipSYp/DSpqjZTuRU781+rD10+GnXqlvMHj9GkiXJJyGk8d8YQqSnkqpbZsSq1e1282Be3mes
cq/9EetsderS74ekk0l7l6cEPIgMQWqoAKyFKWhpnxFWs4b0BrkXIckzGg1HT7Y63EgxtwXRjrfB
OikSkvRO3veT43/H1VrB4IjJGomKSUGA/5H2M3RSAF0iHO+THZ0BcllfTF9EZjfD3pJL5oiXRaOb
um9xc2lDYTzLTKW5D3Od+EOat1QgLlY4QhS7P6sugdu1XI/ZDy7rAuT5w1PcmAexX9Ytlw4Gs79F
8VNr36/dxe0HDU0ewxd1XVY5SZhKYc8NggZTlTkpDvEz8tRi1peW9cHqd1wxyu4/Itje+2Ki65MU
IW2BMgkgl0jIixSXW9c0dgBCNAIf+qRwRleQz2TSEI1gfDUyWGAtu7OhmjK5prrwy19S8BDVmx8y
smcNV/9+P4eTxGvGotJSe8QKMj1bew4o1MLOW1rrY0WTEaUZGe1CFRGRmj0T40VC8742mPqzlOML
Cw0WaFHgwdAsoC3cokckKVl4q+rXpW75nWlHv82IKtkeEQrXTPcWSmzyiSb3O+e+pbneQoI/RLHn
pJHq0ZlAG0EKItrrvB9MSeGLNouC3G3MWAcprgjL4QcDMVSGHhrRpckYTlRSt5q7XDu/694eeNfy
/+bWaL0jspTg8wjO8Rc7z2hFj36IVwo9HFBLJkYgj+a1om8DRfvD/hIAr2G1Xgsaf+FRfqQ65yqu
FqpcrAhoT1YoVjQ5NPmPnwBl27dq/pyuc0f0onvV5a99FX+gMbJtk6hleKgd2Fc1bt5Una66i7Py
aCq9Zg+H5TVlU/hQSCf/rErl0V5hJWsQvTVSr+dvkUuCLdvRr5LrYbIf0u81Zc0lJgBp7dTznQpi
M/O2uk6FVsNY8/ONEdwe2Ii0NBVdbmGRlcmeFtXTRpmf90FYmqCFASNAM61svKRwaG7RzCFLAgZe
8BfQ+hnpDI0YgVjBrMj75ZAwnG71lcppRg9F+tnPcRW3nJVFU8OM8DduF71vAOkIEo+7Pqwd7M/E
YShoS7Ag0mb5xW6YAHwqk5nwnx8uPka5mgUj43FnKEPOP1INEafCTzVbQ98W9CrgskEBPTePtjUq
ON7muxw9rkgZbCSWD2Vwm5UPyqruKwu6huR3XW8CPrDVY/chriz8KJtq2t7q/CF2N3N1HwwjMeZn
s6wQQ8LougboxAkXI+tPFsVQkZSNwvRY13ePs2aNKppBCnEjvzxMOSWRN2suLlhsleLF2YTcJ7Ot
rWFEMHmOD8V4QXVinAouDxtM/mJZghG7P1yxcZkGX62hBEJnL5i/f3PQPyqCS9zjCCK1x9B/X7Nu
afV4MTcPhOctP1rwh9oeofVZ2yZPAKNLwb7D/LQZ7zSHpUlsVXU5K0u4l2RFefV2m/vlQBv50xXU
fSQRWnUXrDbwZVs4LVpqres+MOGEG9je93hGZ/cal0Qr8pzrzVlEw0Uq1Gb9cOedPcU1kjC6J0HP
BA+hoKcmBLrEf+Sk7tJo+U7TbjIMw1PpVN8v5awUST0gHm6TWmFr78hXs1KtXQK+3ZGRuZTKLkWc
fB++2+pGrBj157cAG+ifxLr00CdlDUC8k31JZ1ayZXABfZFRFXetUrESOKXeaZ7Ytpxx80jZ/jt/
x0w+fTdkdU+yu5jLdBA+ygGEyW1GmRAR5HKEgqKhb+FPyApZWj2In3prhg2f3d689l3TeqJ/qg+p
MB+ppPZlWn+1mTj1SdmFLpeNCQas3wZ5OpJMUjbAs4PA7XsD288ghpZsceMpYno0SZdd5ssSSYEf
7etEMfwt/3Cvf286x5jnoxRyryOAtAlXhuuZks5HZRiPsMNb0zOPqHWxETcy0I/kUCnseuvUBogK
D+xNils/pEZR+8NbRduobl7M92j19AOoxGM6hX/QMm4erNfReFtsCBjkVbIJiWjuE8Iau+PSoPG0
CE7IEBN/0EcuN8rfctILUYyrjw5v5VPybzDRF5d0oYD5xAvtHZf6S3cnluCvlarpuQmXN8+/tSNo
qE8rh84XZXs9AggVYR3vy/SAiRgs+E1CgBuy8btihgS2G8goyO0xWbaadGP1pSbtBJSw58McWrqr
ZeCnOAbmJKMhE5BgADyModjhElE8zmLzFm4hkwv+/NNs8DMnsHQ4BG0e5m/PoMAX7vQu8QpvkYeK
rIjaccMeeqBPPYSMHCk0+kHAYoj+MNI7pumjInumvst8QGU73KCdM07XA4kRxfbTGmb6vN3mWwgR
mGpHKClAuKMwVrj6s87WYtlB+Cjoz86hU65yCgMg9yG3278Ghn2XfWi4ueXP5iDDl1oc3JeebrCm
fUITlJL4onw3e0PBZfVFO6HRmMw0dd90EyngTr/vtWOdWRoZoZ53zEtUvLoILKYVc/ObSKRZZuCu
p0ml3m3qYbUD/1hh1CqHAK3Fl5imLejlORAoWD4Sf7rLS0fHlYI7B/Lb9v/44so5CE2a/UUAKLC4
WdqTuO1Kj5NKkghYAzxbnZWDkMRpE8eBAxh8PoZXhq+iM+fRi6o3gJTw7ANoMFuzd29+Km8S1r6W
mPNX3Lr/djfcYRep65qwiJWlaGwW/8x3pTsgZQMn4Az0HOCqbB4JvRadBgljbzEbftdUIRZivZ8y
mGQE0/gGenDOXGq7RxuhWdDHRWkzUTqDQrdjAC8PbtD8/2pwlImjzfDzQ/vudt1ZNy1074Gn6O8w
MYrNquZ07hHsJTeDmEZCactrxYO5xYxH62e/cl3eijxM95V6kH2mlCt6z7PXpftLcvJRNPfTtgHz
Fwlunla+mUTDF+OWpiwMl3lxEBjLetfOVsh8fW2z38Quu4nVbmV500WaVW/70b/oRw10hQWAUKIv
BgW3ggwUWI8ff+bkYPevQRLPDu7Za/HaM64y0GbmCl6D/HI7YxkWLxMhOpPpWd1JvBfZ8CXP0tO8
0cn6m8qydPLeQ84FFepFom0C/ApvZZDo/Pl6Lh7JG5QKrD9vqsY01g1e++RFR4u4EqWQCXT33qAR
mW80fGGvjWLCyLFhSpsSCMN/uAmXrGgs+i6xywUi1Ej3gmFrizlaOMkEjYPpavetceV/GiQPsG45
LEy79vwFv5jvzGgh3+Y3P8Q2Hz+7ikSKDryd/9QGqxAiSw5E61W9UalFR7ZCb63G2VUbk7G65Ijj
vQF97wNdS3TkkspY35j21hPc28aqLXXREDZ3sRnnCm0W+f3TcN6kw1OblEW4jlsSahVAlm9NWraW
F1TRQtlrCM7mcbctv/s/vr11YA2xt5Haq+ImTYKzZ+YeS1fAofGYEynSKqtBrOZ7PpbifiUwpz0s
mzZzUbcLz8/KrXAZNsSxZUbUANuj0kcpp2E9PqYe5DzXkcn/6gCVUOXqm/TMV+AoIlfn4z8fJg10
aEfYKEdWGLzdKenbYkxlhq6cVLV7kwL4oidolpmDqn2gKfwwToFjhNTV1yuopINSfDanKRHaKu52
vfkAnhjjH/PRr1OZ7svwTLG8ohD47HMNk1ozq0R87WS+Me2IzjsZjwbpxS5TGzvlXzLe8IjeB0xg
FLUDlWosS4Z1o65eNUdS1j+1rtf7OeM5SyX+M8KlLwYHt2NJomPWTkXpwxPB+dalqGk/lukfQs3l
unlN6unXsIsLb/JdzslK2X4HG2aydPPZ+ZUYgKz9/GgNQ5iUOciKZgWhTvVoYfZCmqUEE5wxaFFx
RcCNaX+vWPOiCUPDXEGEeOePkcdar4JOQJPKlArfCTi4r5tAnnLxZL1pxqmV8y3JRGyv40SwIZVT
4PbVOMcZG36fGq2EMWdSqyG2va3C2KfobTI63Ij9lb3NfgQpm+L4s5btRxEQBP66YpoPmvSXtI3Y
/Y0s341qhGQzZrypTFCRux/7IvZ91lqo/x+45mmpBrqmNM/8zGyEuamXgqB9/hN37uJOhM3CmH2W
pgDrXK99AIo6M3lsMZ5+ru/TDvJL5nv3w5buptGHpEJ7CbjFE6miY4ZyDFmBUxniwc5LH7ziQqMT
xSERbvhJFAuY7+M4oD6pOji0zGHftlQXBEYPhcrNtPjLrBlvj2hYdhlbon0VLifnYmr1TFOwHFo5
EZs+e0cLtEuwGROF0i981dp4A0iaGpjlSLfVba2J9J3PBmafpcbziBB1Hum0Y7sO+jCKiU22fjGT
HcAUTK7Gp4Zd1TmGSh/FAN6QK4rkF4P3g3LO5n4SlMevD5nSJOFLmKL29Ein1+LCMRDOx1hlCpvB
z1MYETkQ6v7wzIegwPJA3sRhmlzII0yfor4gcaiREhbtIcRKFSOx09WV6ciCYhnifGsBcekiSWN9
hFqEvV/Gqt08VioPUTeLfJEWUCXVtEoK2YnSZlhaGaMGJumnj3dB++sm0QcQhMTDKpK5cF9vaMWn
gvzrkRWPV8AD7clRdRPFWjlAIdc6SGXeUTc79sEWHkBK2mZEkW9vpGWSe74eKMRalGZV6IIZ8WkN
9aemFSCaO94QimjPphJNq9ev+T2JxjCdl7EeaxCJUKkh3c+8tACiF8o6xeLvV6/sVF1jnA9bE5yC
iFHiGA1bQKbD/NewKNouz5KV7mynz8xphg2t5O9lu5zGPoI4AtjXeZOFzKMLAfuqxe/0A6pxonBY
/efPloyl/clZHHh64LlswBjaJRSwodmdI1ck647chxF2WS2DJCEYD1+lPozmjfAisNGTsLj9SpVU
vFzX9Vr2Eb8NO+i9oMM/ShbWFsi6WTi3whqIbgpk3YkWGiUzIKmyTNw9aJdN2btDJVWAVeXOzPKf
jMZBQhe5KsgKgA1AYSm0K3w4Kph9dJE0ky3ha6+UpI1rtWK1cAYh7rGJ16PBf4CZqkkLRhsmnxHA
5KBerefAtxgEoHBQATg5/t8FMg3jJgFiaCpa14Td2mItpG4JpXcMwBWx+VRyrEHwM8U0u2rSM6W4
Q7qs9xizTATKBbes8CwKARtePdpk4h4Uj8NFrui0bUsaYXCbUCxO6J8B5Wh8OJoE1TuQtQbJUqXE
nBr5Z4X6tB8qaiNBijQe+oolQZ4W7SV4HEBwd22cUEQAgJX8UXks5Dg/PEedjD0lkGcDFrsx6Ztf
OHRQqg2B6JbF0icG6NLYy8kbxwmvPtZq0kNVOopaDVCMNzIOhl7YwUEDYglPfiStW8Rchj/KlUIY
ccffU7i7nakfZyScb9nSkBh53ItnvLbK4UQCr1VPqrwtLsrbwwrbsjcyrTAQP4xYptTZtKsAZU0x
UlRZ4BDMYuIAwbureOgLt+Eyk06JBNHVOgHlvS0Qgrl5jll4I38Cl/Di2Z96b7/nZIBEDrDvzMpK
CXqUMYJ+snAu9Gp4tU6d5DgkvZ0yBvQev8CfxcIioVgOzFojDZHQJgHwfq243NEBOuSckyX6sDZ1
FpUorJ2NXOxb8uhyoLUkt56UQCZ9t/5Wh9dPMH3ErxtANomW2N7CE3KEbQxBz2w2USm51mqxWETs
iAOXXOtErPtVnsCSOqmLT00Wg9P+S09qdHgUtpTVMnDMp4XmqHdiigjNuUWr7ZRLynk4U61faqVm
e2rPF1BRFXfabh4URovhJX4hZZClEdD1aUtCaDx1s7sJHlvax1X0BNjRw/CLIK8wYytZxt41rn+t
AT2tpHd1v5YiiU+HmSdO3/lcuK0gW6eOLvcjzGHXrHEHJTJPCJqYmjIo0mt/j2AI/kMP2ozlH7jO
6kR7BGzrLQEYhBuVprYs08I7BjQa+rWPEl+vR0/F6Nzs2vl6SKNRSoKIH+w0k/fblGKLj10XzgOe
6jEUi/I3Pp12zllDFtyzv8igWNmbC8eEl+F0OadMfvMP2JeUMemshsT+Htrr265hE1ssKOmB86hQ
Mm9ORCCS68btbeOxo+o3e3JXchFWE4wrexIaMpHxKmNv/XLLa9tsYsxQqZsqG4YpH/zCoZpNQWiD
ciuPw2OunIGTUDz0v/YVGHsoi4puNI7v5aIfO2U/yASF8fvLCQ8rOFHMyTPpGzuHHRFjFM0ryWpP
AUM5IJ7IQvNxxtZgfTZ4VMYIVR+/sJ07ZTR9NKyOYKwGyt0xfec7qnSOvmPMWYtDLwLHOdEFoBC1
+sI8QUBkAyTUECsA3ULBXAX8fkgh1dGTdJ9ls00JpFFDGAXPBBuh6DBuT9BhLbErQk5rSADOmE2p
o2ZmAAyieYSXncBkXjN4aUKJXrbGEv0GuqHf0fYhVbNH9PQVhqmWecDncG5LcRNgxIjP8P/VU0hX
iBLjIAQqYuglElRBPRC4jN0SiDu4xDKQBlfWPqiKSPHk2mIxPHQvYt0yddwObd964GgMkaassTJ6
zaJHNiwRgrp3sL6iQMN4jehhFS8ejlVEGZzS+si77Gpe8rKC5O192QzrZVV1XVjzIhoIUBRWYyP5
OD0edMJHp42yegffMdmdiUY+Uk9Se+N1/HGAfkJZs7v7NVAVsDtyu6BnTVFQ8eZWgPz+hEG+dJFH
ALvjr3SU1+12cAWtT4KL8JKj/bkdTZiCYIsKeZ4XYRU1K0NrXJsj0Rm9zU2Rzf/Y62G9oQ9jdEhA
VusCX/xNyK8Q/XTdHtga6BmMZPr2PclmEDsWUdyHwV95J4gj+mPnRzoDbmB4AvdJGD2hic8vtqf9
ioefP26Qehu1P3K92YmBdDExdSI4oTXWQQC0v7HujdbyvwdJyX+uWwDGpZk2FarwrE50otYjCMuo
S3bMML6YlFUUfoVV0vVSWtZgsEOnFDzOsLD8grYm5gIFLuYG75rAD6HmhCNuIE9NjjhwmWNyuvU7
0X7Y3TLbNpTQ0IQBTB0L4KGzAmxlKVFMMa1pS0XKXMoi+wiekxAvVi6hlC9XWmT4a4exh8LUdUzb
sujcXrUnOn4vKcxY5nBbMrbgB82LlZS1Cn5OYQRIdUskzCEgCnEBDH1I0Ew6nZHgX9fF/WEkynuN
Xh98HbgaVUFZjJnW1BTIM8ghiUQpmZJk/4K4KoRVsKqc28YmU6+0NYuljSxr5cVstsJOo+XEp3Dn
0PEL/UrQCRseEFUXOltmqH1QUfNCjEdUJyfMWVWYbZr5SW9ueTkc4kEZoXu6+9/BCDkIfaGehfwo
qkbsWuZ9+YLwkGFO2aS12jvDLfeCj5UxfShpnZscQYnGsBhRntuUXIvJcxrENb+K0Q9xpUAQnG1b
6RXQSOH4BfMY//09N3P2RYlLlD5e3oLPcI1WITA/BQjKLtKrJ2Mcid7rqxpPD9TacSEOXr0yspie
0RNWDV+1NktNRCAW5gVsho3glVnXQjdH6LEYGK7WkK4V6FvjjZUxkadA+gGWijObxf3Oa/uywrM0
yAk9d1gzYt7L92/0C7wK1Z745Ut6WUZhI1Z1WKLxHCnw277iv1OZuxwAIfHbaDa4eAT6CKEcMo7H
qoelZeG3nxACVqsWB+cCatRzB4Ntjs6HSwqN12hs0DBP3rQAfR68J0i+pXGkURA6yvuyZAyp31U3
3kj0wnTqFxFWJYjOd4DTZQaY3dChRgC8no5H7/sflf6DvuyJEmSUTOHwnI6A0uA5sHFJFcFpFBuf
jaqNDD90aC8g0B2mxLmSVfakmyZGiVudU09fuhM6CWgnafCj57i/JiqZb7N1//wJcIDaW1IMBSzK
/ezRdziFj5PsGccxDbRvV1f6hnIJWQrb2ABEZ8aolfQs+BMBVl/pcJTHljX0N8z47W8WM0VACpMF
qVy+RPSG4MFUEET+zmm3JOPlJP2pYLEa6fyxTdxTcHZEKm6NkgYqf4D0viX5GpkGEtdJI1tzNa/2
MBtoItW24mvKti9iFA9qBd/h9v3JWjXXF0kcNpdlnREh5+fKn5LhLzXrsN8BIJwlic8+2Q3M9vbF
jsU5AJ9QIzFT8pHKiy0r7lHEwYSgvO6zF1cH+2EvrQGCB6fwjrxpt60sv/UrzNB+CuMJdYCVNYTn
7F13QW/B+ra5Vjk9QpW+YdpNqiSYnP33IEh/ZbYq+dTJD/7qXqDokqiCaoWGSqC8xRe7n9mkfoaW
dZxR8JcRqfIhRt6DRvdbgah9yT6nLq84yZb3T7AbwulSJ/OXQQ7wC4tetdfRhI4DaOPeJpiw1kZv
nltFhJNJe5m2HIuDc+toltKOh7gbdzjYbfqOZ1DRLrpeAkgLPUOMPYO2R+Yx5l2A7nS+LJUCOOjG
F4GGWcbmkpryTMM0cnPEhw4X3waUKJsRvknXYjoc5W0/Wo10YR8Ctv6S4c5LEvX+VB6O/u5TSKDx
ZHajreDuOGC5znZ2Wb/x6bs5ZpjfpVUp9qAcF3gsDrgdXfRMY0CD9ZI7UtQG8HvMRlxIG9VDxWuV
oH6UPYNAjoPSR25EQBG3CE5knOrWswTQN2RH5L4HnoRg9vaom5PtimilDzhM03UxiliWkxxuEYNm
LdSzF3PiCv2W82qX2iA/iSOXNV0xPIYYpr8kFlE6KUQHUfHD47CuXFQS5Oejoc7oXbrjAT3bEp+7
0bDwEOEYqpaPpyitOtlRRMF0i3TW/zE8Cf+Ey95QfQKToGbFGXeNn+60RTK6XCphcG1OMZdXYdAT
3u10rMzZJTe+TP8X2p6JNvGPtbWGOIQ/O/2LeDZ5hh6JuzX5tTdQ1zW2kTMMDFVoNgh0IWgz+qlT
Zo7xSZllu+v6JbJu4AgeOWoN6gGzrcvLjyUibb93l70eQrHDhZbftMllA55HCGzyfRYb16gCJ4/q
nOi7kLkkXOjQmOdplZPJFsdwxE3UZRunDOZWTaLijkWSbKJ8pAPl2qib59ezZiixpxbDzsVXzX5e
EdOjL1voIni8As1MxkTbKqz8dsMS/oxb0r3dxhvN+0OQIfRrwfAKJNaGCrzthYJXYPqKcArAax9+
6E1qTx54/ygisfWyubs2uiMFivfQ48WMj+7R2RPyaA3la3Xf1fXa0vkM/nPYnVbI4CCUndHVLmx2
xqwyxEVMUtvNGeE0l4OEisLdFTWojsYEZQoyzzLMFIB7d25oWRV1drMyiPtQKAyCyU0GXM1H7/m8
Fy10eFaqNrkb8iO42CV8SMNr6pQ/KIg2PLwkb0QOY/7sbjdM6tfTKe+ew88mRNFWIldhbUcK4gVb
/pbUzw11efxbLaemaosoZMnQ74N99msxaprtsb3QwSTX6338MUP27Ojp1rrvI+eKAvBawmWGO/9o
sd/CfxSl9zOT/kb4Qe5ZIpe2YVFNe4I1bXMfIRCKsX4LIBcH/JNkIS362c0BVL5hqkaN6ZD0vfnc
vTQUecuw66RHNpZVhSJJZOG2/YdL+HTMPXDl0UAyv3zeDzuuedMKVAx6hYcoVggtsgIkvxh4Smd3
8DACRNOmlGkZ+kpXswrAOtd1Atu01Mm30ORlkY7Sc10gCx+UKdq7av3U9Gm+SvtupVJB7+tjJivm
Da9A3rkpifdwYFyYVCnENQWuVwfHM3kcaSTGSncltwgruz8btiRbWKpUxHXDl3+JD80fSYVRLw5R
BEy8b//W0bpDa8PeM6lNZ09i9sArwZaq7MwYjflslEcKkdGo0K/CjjWZlXblbcV1KZ2N9BJHl5J2
ST7zatlVvHlwx30tAZz4/LfTkGKmtWfQejN8q2M9XThfrN344t8Pa/Lk1u1KLke+aOrM7HoE1OoX
8jW3TMSetUYYl0UBDXrg0Cm0rI3NS85X3BeL2Y1e0ifet0TCnkVW9G42JapBfVTUMHkc8z6JjNoS
+q9QCSAbllFAnolBQvVs+WJP7n61ZM9MzoZyaM8G+/lT2nMyp59AvSBSmOY6lozToRvzjsH2/8JM
59oPUymGY5bcLoeS79SPq/h7rB3LjJtBVUdrHvaB1LWZkfPNSUUzRarOrLivkTtLGR1qRokYwkmj
FoQLQbjL7RssEulkf0VL/Bhy6+r3LFdSdJvrop1le8V6i3DqFXUwsnjKn/9zuJ7x97oK1e/ZE1G9
D5iHmj7YCALtKlKQCHtyU6tziLPi7+GdLG1viEc6pbRWfpuc+znDRfwnc1l5IFYOUeCjSy1iGBrh
yKn2cO5HJJXh/oCfFCQkBKf35q+2AAHLHeog/R4gR8okHXhFEYmvwawTdr/WGllNKJYRdOCEBAHu
3a9zknY00yLfbHfCb3B7Shdv5rbCTWrnaXmbEJF2w8k31fO0yEJPU5HF36/uKU2uwYQK96nyB+ZJ
gArit3EPmCPSpQoOHZtHFMK+jQlVtLsGh4soTGU1j+6WbcroBE+ahHzKLhi254I9YWYqy1T5Zc9J
TuY/jQcA47m3SqYGb4eNfBstvSWRu0DsDnMQHauOshz311m82+PMHxOYJuKco6KOKms84xKGi3Ca
w2gbDrGxXPf1sjkniBvarHVjDAtHQNGzRA6grHZxNFgj+t9B7P9xKXG07Yykzl8X3IaR+UNUsQIW
1sDvKbFDgRZGQAlhZXtaM5be3/wLiQWzfoSCaN5wgRIfvzw8gisG0pLRx+OZznvUxLITm28hJFrF
5E11AHH3zTfSyJ4IAPyDkOwRyjfhO1Cgqi1N/+V3UIkQWX3HBl+LYlm/RW8ijF7hyGPcLuuhZSUA
xBkmWusafJWhk54pUkRqN7gYYdE9UM21kGCkMo56a5SFDmfNTyf/kVzagS/FWZayfIZn6e7t/y04
AZCzP6GO+0oWt2rekLP7ZZZMo9X4ccG9VlPpI8ed5Iym0AKgw+xX5d6NQj5Nor247jaq4kdPbSFL
HbX6MtscC2YJOQ+JkeayojdES2M93iK0FpsKsJFaHiGFj4qLwPNFnXQ7QufGX5Y+NI0YJs05gbuw
GnUzma1u07VtkLVPAdoG0keECn4urxdYyjDeXtS1VROIhK5PGW/rdzuaDFGIe+NQfl3GEv3tOCwk
WNCDPkoY2Ar3aZ3sxtFNZbsq0kALxb3q23xhfeO3q3h5Z/YCFXnDzjtDm7Smdpkx2s31OuV6ubgW
VBCgVPkhfEiJ6T+huaFoC3eYy9TcoLPCsr4Df1UWVD1l0F8u819NDBCf5aZ3Fxpj5NToAYmNoAvB
230Xl+UGewkFiv4sqGiAqhDZKkgFLB949L2Zm0cZyAwcNqbYRcJCnv45B3eiy8Pe+v5NA71pUHr8
f47tVkLT4sPH5yzShuXeWMH3bU5KtlXAupWNMRiXCXv7WnQwuKEAF7gDwP3qqUUAQcEfl843j4bZ
YpDM93QC3i8ZIq7Vc2cv9HTQPoTK8IgnA/flhYBaay5+pF7bZNVCfF3IWp3qtv2P7FY6e2w3R+tr
B9q6pyNwJpkStSNNJbC7Z+XWU1T+TiUEAQxY/5dvbzK4NxGdlrb1Sh9I3IH1NhjFC2vfTHkhEo9Y
viSLcJDx8tAC7vgx9T7NTHdbKZZNEjfzXTd9KSnBLRaQDiIUUooStxzDJzff7tcW++9CLA70DSmZ
wPcO7pnHaObOF5lTcewPVDirWPPg6EkbUakbINg2MhJsAjxg1An2CmHBr7cYhvvOQvEy26SKO78z
aWF602Jf0JkV60nirGDGxYQc6uOaNWP+JXOFA6VwWoCPc11URG3AKtRhni5nswwDE4JQ3N+Klvnj
FQx/NHnI9hgqA90/CXHjT/EEJhE5H1CYpvZwQmekR5HV5iAShZppd9ToN3J17AKGG6QBR31qEyW+
xY2KfUfZzhTQqsbB1SL8Wdrf0hD9+4aNjO9DkJcpAZErSp3E0RUMx/86sRW7nq3nAyvUDuYkSF8/
fbHz13t+Zxdq2HJ3q4dNx/f2++Xe4GKkCSTld+wjIMANsRG0YNud0Cj3E2kwAeXR6M959Qdem5hS
yentHIOjYs2fIZiYSCgm2hwQIBUhqpWyCpLpQFHId7CVNODqeLCYQqm+WrK9XweYyor7enTeu5G4
1/R2kRbwrr8CfQdYpF96AlE/zAxfp9vJWE6L5jqSA7kd7vyj91MQKRJMCLIxEQJ8KA3ydDW+XFWN
v8m6vkgs3d00GQcKn9IftYmNU4LhqXVL9ly/RObTySftcn6qTqR19X1CaMXdfGXAQjQG9ineCoTN
87QzIYoz+LL48dfRebF60e+rRK29quVbMZSOm4FrfJpYtCUE25iNix5rHJUwQwxouvxhTsjK8CjL
IIYmH5y1BOYNtMp7y9MvObNzAho73B61vkPiOjDuUSOKeyM037Nkd1KT49CGaNznQZzoPt2uM4es
0lfDeyeRhhOfp4BZOM8fGPC3qq5124xrIFcurUiS/Dr8glnv7FMpxmVlqqGRhEZ3/ziU0Sju1PI1
shUSH2fsTKBx/xF2IwG8yRpZ2FxF+wAsemSMkDaIAsyDgX/emXS5uOWiTzxQKX6xI7R6NRrD5RSV
v6BqkgIFK0kBazCsVkdhIRrLv0hlZrXd4hZl5+/VeLmJr8R6t1vi0SFXXZ23OT2vaZT2q5RY0zoa
JgMI3UdvzloohIsPkKtJav8pJ0AOuTBGEdfOBu9P1avSQXGCUktjDRP7eY8hUlv4A7IscbsG5bnQ
HkYJy3rsKHRqObUDQiv2wZtmUPNt7rnX49Sb9wDhMMhVPUB5k3BxCG2K3bnnU69i/mfSX5rsIRJm
MyhwxZj0AOFGV+b28V5wvcdNiiZPEYcLZO7bRVbWz7FeCY9GIaYleOUIBhmLksjYFLZvkesGYz6x
kykR6OUImMuQfWhzcoRIVVlabppM+Ue6QM4GHRBu0iVV5yIL8pwXHZrkmRWxpXX98oSBsZFno53R
Z4a+6tOgTCuAicl0SOqmvUjFwdbeWOoxvx/1RsTl1oLBnkI/+JMD/f8f4q3TQVIM3IVtfylExnC8
XC1rZ4WW7A5MiQ8B0uD0Dh6LAztuGFbRqrXbf04PcPFHLWmv8IOhO8Tm/GZQ57GcQOYNN1Kmq3L0
t0ZuMVL8bH+/O9rxwRqcfmzUHT6pxpIqpbsIdZ7VmdMJz8tX+zooRWKj9NAt8Md8I6NvG1j0nIPH
tZ3rylIj2zH/0O58uUI1RwAc+HEo/4r/sk79OL15EZym3c++1EMydN1c/TsDbVUhF3a54ObolgPh
fxwvjvtag3GVZU/Jo6mVXUozhV+zASZwbKwYImDsJ+CRTo6OhPf1uSmml2mIvHaGlmhI/plXFpoW
iM2O4GvcQrbGuRtdwzlSkSubHS+RpxpuC5epFqVwIpM9wHyBPQ3HduNgRGvcfaOcL2yKXx/MZr3b
O5eMTtkxCNJTeb+lPqjvw8TM4cLN15x7HjLDXlyiMnfCmor5MUhX5aMUAGS72hURF2BJ7B/2cLmA
g8/FGfjKET/8qGOT/tBjaM4j5jJ5dtAU50XtZvsN6m6R8IxyiLYSfpibbs1YyMWq+MprK/3Qdjli
JpKZTnVgoPS3kZIBX2E/F9jaYfYKBd5nUB3TocEZnuKB3JftIpoLAeCmY9ADfwO791KeuGFh+cId
m2wWeUAkXQoNJVE+16ujdR83ar+1UsLQCnuuPyIjDoPxIGsJ6ptwynMReKBqRPRTm0/rAhfFbxxq
1L/rtW77mPJvJCHSYMTBHNjBpxaE7FFnR4uh3rhh6V42/ETAbn/qBMoFOiXZfp6AWZcp5agNJvIX
+cIxfJZoV+/vYot4mcmGe9rhTdWIhWmpRok8jVXir2noAZ0PWJ4y8zZVWNoHhUVd12K8tiJjGa4j
fcW3JxcBixS6W3cE6hPK7zXfsxdtsVaqwWO/lcuJ7fJ05msKy2lP+AxJhm0ikLQrFVbxwuHuaCIY
zLJKBEhsYleq6Yndb4XEDBpRfJi6QzqAQrZe0nY6c7NllnQ0gtn3INUwo23EI3Y+t0XFSZlMg3DB
0YRQ/idIXSa8Lmr8KC3WVKKq0n+WoX7aU4d+uMdiLr9HGTFD7NbWXYW5Di0jvOD+JerNkewnhuYE
wdyI/zaILOUvzZyEAsz3kaxqnvKtcCCfn92GHlEEQO+FIaYStXq7iiu+h+OBt3hvplvZZzVsZebj
X4SRyGLjlJeZ9diQoeWRcCNRu4moJT1VYCHdrQmWD3QOpY4k7TSlGkQ/mfXCPT7/8+kkRo9pTfXS
llOKg+dv9hAxubueNZuXOGHG2a9JQrhfgcoETrrw6r2oEg4fbXJwzHFxx+OHIR9q+eBg3ERgEXOs
Wam2f8/BUI68AqZ/s/sVAyzvYQGb2v3vX6XX9qcI+0TGdDsK/GSPjoGG/qxO+kg/8Bl1hqk06yHt
eiUc8Em9LbuVoHvbOjwKrZ/Q9ycPnTo11Ba/DiE6m0CpaSLm+P26B1k0urt85zzheOOILmLGj6Hi
DlA4/buhimewQpz/qN5X7uh60K0wl4TqmdHhCrgJcxtxgHBtQu8AFsAM6P5x7IPTnMXZDKq6pNiS
yAbrhbuhrjy1tdZyF6Axy5bR2fj2ihlFl1LF4UavzlemhiQKM2XSv4K26Uy+YyJAsgAfzllbElel
v6I+mZqau40Q90l+0GBlE6FFweqo4cO+/Wv3TxIrVfXcHOfi+zMW7Wy+3fRdE8tY7Dn+oJqZOYsm
4MotiGu1dpncHePdr4UocFFpTehAQvBU8SvEfHzzHzQoCgtctDIh6hJa9r/Onq4z95nQtkn2pwhR
9/DMSgSkOxgC752Oa/N/mMYL4PjNr1X6f0IVq+LqFfl1G7NhNDMorlaVeOZRpCWOUnYBLaJNEpbq
b58RDoyRAgAiKmuOnYOdXqmQ7VqhrfGbwg4613UKlTchqGcqj7IE1p5G6/7M15CpOMs+Wfk7ODez
3Q5lWpqf3X9AF4HPkdRV9i0uRVrBKq+dlSXqISR5jwTFgpLTFUVe2HaLI5U/fQOa/qIakYDL13/J
MuAl/BHmlYnCJOM+Ss/O7GarAUwto0+RzdjeWC3CFBbRMQszrjuXhoHGsTQBvZ6tVvE+qO+GMThL
fyG4chrhPR23Zekv/Sq1X83aQlkHt3yvF19I4/wainosf57JIPcbVA/yku6KxAvSR08R/fu5Rnus
ST6cGX3bHaV21sycRCBcf3giB7YBbwZuKf7fHI/5e1Waur6O+GnnCtYBRByeQrOj7QsngwsZxIc7
D2XT+JZmLWnV3Te8+fr0+VfetpF3WZceUz5hhC5GwyQe1dkvDzq7PIOGnj+xe4pw7tc7mNA4bSz2
0gK7sBE/fS9POJtHjP8ObxENnm6DKPDsLutCxqCxwIgCt5pvXG5ZRNKubkLDT9zd/q9+H1h5I+KS
rgE+ux3rfMcWOP21txMJJVBItCJnZW1J/jEt+fEFtixTVJqrXnkXluf3hXq5k41PHW0q8yD2UilS
5SiShv9MR/1d5A0RpCgEg6XCG8Rvy9n8R/2C/1n1SA3pzLJQS9a43rlsxs+itmpwx86tNhEv7Mmb
DeIWVhs1A9yy5Z5eIAYF/H57GwdAFFd2wxO3GGxV8S/nsmkcKkSaBZk16okVp8lOPyuocykjisU6
gMXoE5Q1FSCzmIMEYjxedaQYkUd/3JSNDdMgl6ZOO2VMztMRMq0/u0qPmjIvh6MVBNCejYijEMDa
cbKA7yK6yi1Afr0V9rZf/Mg+knn6qXSeHdBSii88HquyI75xYcqH83HatD8LbnuFJVaQpVHCTHDm
zINF+EbjkFLBNFZbAzi5M/zmilmdmZRmxIM0+TlH5PgSKqHUMA9SyZ/DjJlH4m2OviPREBfhD6zc
PhjCvAGmLrQ9524h/PIa+RnaGsYHekzYB+1u83F7WxbSS7Z8XO3WDuwsH3Qqop3rGd2Mqbnae7qj
cc789P3QBJ6OGT2OxXCJ7bbZRVJUXEGIF6r6uNCG9ObQ+PCUKRBpzMAZjl1PIwkgSXlWmfmcD1/j
0Vd1zGWX1JYHTQhX9Ult28kdAFaKqOIH0qbuVS8W/AkQEhdpIH+vbu5PCyBSg6ITJmThCFpZjN86
3IcgtFIQHn1jg+ieaZGdc8HSAuvlT2e7VqdWxjmKdHbokMPdM2/TrVNs5lIiZdKIrmmAdSErvCBQ
nUBhjStPqXO+PiO/ibsyz+zSx2BeUzgU3onUSFnd/+oV9cfUD1uPcwUMWRiYv/Z6HrezDAPWMK2H
yilysdx8OOqs27qRYUsSRT5NeXLGgMzRmJpTjOjUB8SC0dG7YMr+UzTdtW9Ajgyo0HFXOK2RhK/b
Y4vIZDf3RT9DRMGNmGA60OSk82zWlC8SFZjmt8P8TXeDRXMGBX7DjD9JRojuP/lxvIdKEjZqQ7so
oIh8OC9zHNxowgOrcxfiXJD0VyRFEKB1JWCuCIcuDq34pIreXMfiwSXMJqH2tK2xgMJwn6vk34mQ
oBPnzEFugD2h1mJJeTCBDEakivO197cMgUbSLdDjl5NakoX8hDTNqAtTYsZyRnCUqwNCTmZDXsrC
m9k/oT+U478EosaF1UYykEw8pIfSkAvuH9SvlCwIDl0uljkj+rWLVWpsNj+MkM+xPJZcyIORAOFO
JhNwqA5Azg5vaS8857eVxJyTiGaGPLxIcjkbdrBBzam7CU/+W0UQ1hWGhmOu36OyKuq5IsXmjBY6
puyUnYaLICQ3b7F5dZ/5FIOTEgLfSsVmcyNg5DuirloYWoXLE8UsijI5ZL5jIpc1iTRFNpCx0z99
tiRh0Jl1ITJIwwv5KFhBFJAA2zmwkpgRRhXdTOCdKetQDlGau6T+5m46eWXHNno/7VPmaju8tyb4
o/TByQw8/cfl4oM6VXKs82ICyjnIiS16nHDiQRMz8F+6umi9IDx5/SGm2i66HMcKj5jk2W7kUnhl
5AtrcPMq0v2BRwWecXTThQGdO47HpLeR2Gh6MUMOQnbg3dtqAVAmrdnys+rA7uQ0ogk/fCYn00OL
R5UKmFYbNNkibjtWJjCZo9Vl2+tBaLjFiw6HOXjMGkuPf8kwJoVZpuKKAMI47HIdAj8hVLJ2FOmL
M40W8gc4vybpDni7yhHz6C33RiQbkMRX8pEsEuTlPwCPMKSKPeCdoM8F34fAn4LfwbZxRiFbnp9d
lCSJS+ez1qa5p9uH677oapmnnFuwwap38VUmxfLOUj5XBJ6f2WRI/02rjxHVF6bsNtnLy2jxXOG5
m0uZoUGS1X3qimM6toyJ2TSuqqk/S3Gr+CyiQjT3UMXajMNkzbQ8LKFGH8qY4fO3RqfjXiZSt8Db
24QuiRj4TIJwBPDE+x+5DdcgsQwKFc4QSmuQ1vN77/dzGZ4wZQG78/oorJb2QHZ11rEKM8B7b4Tu
ieXNhjodZWSTE9S83JdE/fWs1xlxIciIV1v8hVcccC8BvDOAZp9ZihZ4dsO7K/1USO7UIHtz5uq8
QjH9Y4GDWJK50LTsKT4TRyqyJJQe4gGqWINHvsa2SSgi6mTILbSqEfwuwCkItxGniJTi+spZsNqQ
oXE+XhL3ypKeGG8bH4cTjWlVGBFjh1V0fqHafHelbKgCogZIuoVixQ9KnYZPXZN10DxmYaJM62U7
OENrFbjUx3nXi/N8DjdBK8JF4PvvtJQ00R7PYgDY2UQgP6yI6O/PcAjbiuiYoyx9Y8xlxUhL7mpB
fdx9wM+kFH76HD0qu+8ZerQsZMnwDI82rAevWIvC6SBD8QLDxNDXzttoaMGHiTGVjheI2Zk87FHg
lC/rINA8Y6WCK9ExXU+ukNfbhlrJuiW971AlOGZzQMFOYV6fonz/d1qGmvCAogb7LJPMcBywQMGE
tYD+jblP+WcaNEZyG1eZp0HSW3YQoVDTfkR3nxgGFO9mZ47uip3pitg2GG+msMiFX7RGIPWdHQzb
e49OjNOXFrZ/xt37308wjIfCAV3G7If1ZrCV0aFYLrI5MMgellNEbMRytbNwPpwfTMszyYwyRI8d
sYmE2G/XdmO7XSf+fwsuEM0rbt6y7SSaJVV8rlEOtVKa9X3x2uY6uxF9ctWsWO1Mjfp/9TPfhKK8
VmkCpJx1KCe7QRY5g0w8l2ApZ3y8iI6Bk5M/iQWKy5oRe5zEcsOqlGTEgdD87QMlrxSNJUqTGMr8
GgpvsrgefvEBIJPKBGrs8KPlUg+lSt5v1nuDeCsJobH18yOQQK7ljng3OIEjDxrZb/5yCQJnOOB1
+dywKOXbvZ3pJMdqpXK2CGgIkU8AS8nzkZuGh+W1KjRSoseACBdrCgDx8KMh/F8tXNYU/XCYdUTi
BsG05GeBHvpZrlvFejzLWEuxsajvpB5COET+fGpNp9M9wEsl3Ba82fM41Ra5y/ODX0Iceog3GFxy
7fF/1B96YgN5pSNB1+XOeKdFxSYGcm+dFJF49XXSs8G5jVJWVgX/MOIozsM3ceLeRKYnUYrkkhJB
96H5chhXQqjDFUUyB2U05tsfLC/NIvVwffEI3tu7ZyyB/FiLq84vX3Z8BlUXQGaB4VtkRgijXZ2w
4O8q7xFmnSOcytgXTmO/8LyD/K8072FqtuazSIoZJBH2FeEXOm7jPbZZZNO2yizER1lr6+PQQeHu
0Ppfi1QpR0iuUMkCtvursy2lG1M1Px2/qkhVum6Igzbu7iXBbkW2MenlWMXZ30FDKJgk1ISxKPMa
AAkYR+3lJ7qdtgRuXgxD5PqEKGOndyBMq++PD4j9UIqjirbZil5dgrS0pEn5S22ycUJcSvGgJJEy
WqEBTLvX1u/4ob3nAZ0Of1yUsSb3TrnJl+A1oNAOlKcSr9D5S/PQzcjubqHVKeicvIcFbdR/WmYC
XXRSyLgTtU5165uE+Iz83rghvvvdlMcr/VABSmCfwUxSXVTgqLwV9Vfm6fIDuZShFn57+sjOcSvI
D3Roj2v8Jo8UiUqeCGQc1rIGZAHqmh7PPKmd9a3vgia0OYLO63TOZxhcCVGCFiYqoDsfTItyNntQ
RIQoC2/J+MelgswWSl9ikeqyWnF9yKjFd98/w9rFFnF4iys7gmHa3xbIh8v8aohEPnd3VRPLlS3j
vhTqvCQ7HyYAozEMkuyHADI88v5tyYIZoJqXldZ6er2f1KY44LcKdQPlExPz46eJoKQkl2fz1fWK
cR1VPSys95OgREx7z93Qr+f9pj+fa3E2Dk/FqC8rJS/Q4kRmbbbbkG+23bGpYVuTN+dRnProsLBc
TxFm82Z4dS9qgAR0yGoe17TFk+LXbyLqGRwVbaS2rB13pauerh0sZl++Unk7YNtU3Fod463epgWt
x3xzwVObydWzyefKjkvfe01dmjMDELTqAPWMsekhBvzOtR3koFLqmWIfFmfPkefRu58uNa7VK72L
/OencZl/MP97iPkNUp3hqRK0icqLTnb/Tk5Vq5fsuQgVIJgCtaTsNhtLyT4wrSfZdkbeA4Y8ZSbp
hRYylXS1XpjQvja8uEVmbcVrMbqlKYgZdBdPsi/d0Haf0PwiXv4XJ9ZcRMt7gu+6nd2sr5JOOqC5
17PNnjk7vOeEs/vl+Cd/nn3nu/2an0RCYfj4U52tE0N5eGwqIVHTbuIUhE52T021lKaVTNTMY7t2
5EFmBkgn479Ci4x6UJ+QFYwLQbgIulyD87ESnizPCJV9D8D16aYPwDIFuiRLFMumkF8pzUlwd8EU
r93yr/34np/mcnGxrEb94AGK9EAWpLOYBCmbmcGYlD+rIR8z3TXnQlSpnOYfdVam7pzSyjzsTYvO
4Bras7k1Wf8ImqgeXfRuxuLUf6XQM2+Q8TzafOG/xRwF/o8oj8DrzNhTl8OHelUm8cYZ8O1MReP8
HNdUpeIoVjvHCliIa/BeoZY16RTmogDGZSHsJAsG08mfcd/Pk5knsdGKM4ySipKhSy5bHb9cTDdz
ClWngOoOsqah3cQmYvmE7Dhs2keqHo3Ltowf/gfwm5f1OV9/RY12H2t0vsnD/dgBwnvFppproSNx
09UiEu9KRvdYKZqyeJ0uQTBIyWy7c5gdqEAFXUBdG4Q4Sk4iN19Ot6Tz3WC4YVe+TR6IQ3aqDErX
d55OACjZPCLDlFrO8XPzM0/N2ctMDWX8TWxQyZM9TX7B9dbElu6bxxj317s5+xRNMm383aZytaSd
JeIPvb290QV4K64lvtA9QqXzjxX81y+QMpW61PgjHpkaIUdlyOkuqR/VySF9egxY1SFbG7TLG8w0
viuBo5CP45fV38iF+L8trOfkOz/U+JtlAvyvLkLRY3vcwYwB5hwL5IYSMfDbgGPRdIA59vLdib1x
VWOI3EL5BtZurTGrrBCpkg59u5hctiFS/l0E1ITTyAEOPJUJjzq/GAKqTpPPdJNbsp1sdDFHrcM9
ou6xdbdVxlcZzUHc9cb9Cs5TX0JlrfdE5h/dIm7rHDiBu/Gpqfwolw4T8t+pcyrgJXrtFdnPRjxZ
nyZudFcQAulyn13P+z4jFb+EpV1HKP8+qUS+B8cs2dncSe+aqbgoLfPnE7vgsYAqIUqyETP4/zO/
SvyrpNJ9Go5Y5OGNuvq74Q4hlmivK+oWYIHhp72QnkGnHtSPLCq1F0pEOgWk7ugb0rYp8nwIXLJB
XlKujIXhcaNGA78BuQncNaM65qMRJnt4vZKkptawrGfnKIDbziwsydscPahMyL3CMZg0lIy4A9Co
fU6rkOYGQNb5sntk68FE5GiwLDhwbQFV7NjWve5oCwIR4m+E9UuZ0zGelOSffHW/FUOYWTsYXPg+
46S8DzqqcO7IgkrayJ2O63RUE2AQbapVH5WrUoQjYZEy426GJugE3PZbv+aH1pY6yUQONFSsX8SW
McLE87Uj6WL/5I3eGb/XADk+dgRVYpdYRPF8EKzNYHa5RngVUBD3SMt/2YbzF2ARFXiMZUxeg6Y+
jKfADr7JoZNRwIQzeRU24iXWR00W0NppmAD9hJ6Uuu3fsCen4miHdTBJuegMkH7xtPJpTuOvsXha
LNxrR4MfJlkapzJ7B6V1Dp+neOgqJm+LDuddtaesEeK9z+wPGllfoYsakh7zmwJeeg7zfAok2ab5
hoYyZA93ePPF2OnwKJbsR+D1RWpZ9NJOsfpWcphNzGqnmb16xMcZmNtXziwymj7yZKOQ16p70VVS
sXxjlyFC4IdouyXA5JQYt8MRVj8rJAb8OzftagqUlDZ9P5JaTWvlGj6mBEMlgA9XpQCRTqfn1wto
IMgjyyyWEto0zHxoiYQtm5IVf1zZy6zyioR2LleAwLTpAyMzQcAReFMp+PsdtY6P3RzAoJ8++Hk9
tr/vLzFKkpy4AlporWXzc401rYPXg84c99lAw0TE0a/0BVTtLC3GJSmZwmaXvf/NLc58Yvzm0gpD
/IfDX7uPscEQHVzeb919nZXRCniTFcKwrLr9R/icC4pEcPNPM+7BIG72cXUoZWhP4WZsIXWzfQtD
fRU5ijpgkAzbHPyDNPJ2gs5qL4M6+uW2bedr6QHInpWENAeKaPnRflDxhWyNP16G4Qb72eRdao/U
pV04FShzsz45pBp8GPbl0HlB5wLn7EUdulviQMhlqSAsbfw5CsTNPrFPlymEy317LIKQqzBQZiHW
xuBf4xiMBVvU/RXXwdD+jIXdrUpheJuOASVs5FprGzpVFPqvEhr+TT1TXkW0Jo+SPf5wBkPrKfox
A6zRT497ljtkAMcIbiE5nKyrsCm5EQmKjxGoW0lsXRuxhNjjR1Ycr4fzOk/4kSOA49yw2y4NW5T5
K5dDldrYGEcZvyg3w9o8OLe/L+qumoe19D6mdEePUOObjjQ5yn0D2HHkJvdWJk8nvc3gh+j/Lx+y
9Wl2z2ibjBQZxa22m/GbGecmKLufF+ruSc65pc0svGBcA+njCH8b5xGIoNfSOXe1BNNncpZTWbyo
II5266h3DE2ZiBRhcIt+qFo5s05jPf3YeB81xzAX/2QSC13qebqCjtNkrCfqoG3NqHjYIus+husx
PRegHpl8FyQarf6RqPoyYtf9LOvH3VCCnG9aCxLtAW2IYRGkveZSixCm5HnG7rgx8OrKqawf6vGG
MkXTgukS4gwGpRmlfN4Are2e2AjmMLqJKDDb6GASIgHsoqJlHjvNkNxVfqlYfXRhat88bhIy5Hra
vTovUNbvOypAltAukv47TP61yj+Xmuk76FP26VikflNpWY7GLk6VKs6dTnZGncdWeeMY28h5tH+J
w5GMOk3R5HHXVxGQYxP5gKe0SLAhNa17Ey4KfNRCXNg7FpmO6eHVNtjLPEsMVXn2CisX3o2Xdx0o
QVeAdBaaMKgFX80MP/F3HSsAh74puyVQ90oAfutReBLqJs7pblpIs7APz7NeXBYOs2g9jkRt0uiI
ygjbhLvEV8bZx7dDW+LRUG7iYX1x4Jo68qp27hTU/fV9wY/5r21ZwppTazdWR390UB08JpikHdMs
4xMLzR95gniYMKzX7YOye0o3/icuWU+nWQR1H/f3oj5AVLs0P6Po2kJDA0q+QG+cztlXuVURA/+Y
Fsidn8XwjcQo9RH4oZOJ0ZzXLx5lvH0k6wUdRtKCrpruhCQymRUrKmzXk80GE/o0qIGLiTBNCXPF
OlD92i+aPbiOSUVhzhPjiyl9Q7LPuXU71DmBWVE3J8geEt3PI6hNNsH7IMpKVMyCKw1DugADtKx/
fD2HDiNMIXGGi0tqTfjYBzXFZOyqQEDLqYvrNlLE9Upa0iPmubAWPD/M1W7S5CmxIi/7hkzp3XkL
clwn11XtatF7gk4SlAPGaSKE543jmr9vtWuV9STXtyix4MagCd1ZoKoY6u2v6j750i43884VX4+g
k9TVOoMWUGAxBBfzZWaotMSAK5ZKZK0RspsuvWFywQBqdnHeDmtVSjX6TtnJ59b5Ao5X6gBj3KLD
/6kXjpaGuALpczFkSn0LMuSJVzkPBoR+vgdzyxKPPt5RnU+qw3ewJ7Ji07HFM3lCOndOAl03whyV
NpOA8UinDsqeglzUA1nYVkmGEb3wXdZCcP3iR/z+HBf1/2n+e1ycsXK/SULO2qzfrPzT8unKFXys
22RnfV1qWT0tDx+YqKXlC+zzL3MSvZba8QDXA60mraeOHZdorkyzoIBZLzw2th0W4JT0gfxebV1y
0XKuZysQgGFqH7Oql3XrM3aGEvy1z6ZGb3XpoVrfmj7hEhDU++Jjg0dVUeA4JeFNEgRVpgLyh+ZA
fNG7/WsOlx1lVWirmHSxsDDn4fy+sUQHZWd5YtC/RZvwpSeJGB+YMzZSMFtNcVBAS3UnZblmOu8L
c4Yj7NvAU6F5Z2MgXotb9AT9374ez0zWJVNgtRtcscaxHvxMCVD1PtJWkIDqaFt6Jh8qGY+EhNjq
LBUkziI0cIk3Y1fjsU8XLza9tktDqtVWL/Laglp8ieKLt065tufHXqOwPQ9vToNyXkEGXB3Bj9fK
rAEPz1h+jO6nttVaNWByVbu4c1+DRfvd9fq/L829c1q4/aIdRT+bs1nxiAGe599DUMrV2xCISd4U
LMXUueLEn00IwxMAzDPXEW2F++/DEDIpPjMf6bAY7AxEjXBvZ2rE4u64rw7jms1HVmsf8AQChjQ7
7VQo6f9moKffyxVtgsXgMnfPVilgRikpmGRwm5t+wxeKM1PbekPtgkakJhdO30/FZxw6a7Iszzwe
KlzTY2IAiSGONDLjbruOzO5EHBzoHGmTFUz+pcayVQtkEOZVlFMRhDrKuT24j+ug9Ad812tjkmjF
CIoe34JrUTOOAjOxO7iz3L5ZZFzlntBagG/Jqyf5Qt5YpNTfMeyGnBU1vswrMNwX/qpQ8auTR8kv
upfhbV0tZPtIWmJicthcbc5Lkg33FIlTPeWIBMw/qaemEx6sqDWcdBA9c+EmmzrqyHWH1rlFw0gK
aUE0BOuKfsLi4U2W49wawyImii6ly5RQCjFX5ZX8SklraS+tHoMyShre9cz/saqeVK/8/dKxjwlw
pT/q2sCpa4MTSKOW2+/MfixYCqT1hZT3XHt/f3QmVptFCWjKsdtebL2DaPYHKhsAcqhjkWGXP9jF
k61KzwOmXA1JjZNCZmBBJcHPcHyH7odytM5Htsu5eksc1S1p7eraCDymjeTNS0HUkxnYGUsKr4+k
umcv3agYwZzcx0loNyFCraR2UiAvId0Y/IGaPW6sOYAoC2EBU9mD+pryTG/71zB3vhYM59ENY4E/
6Xa+WoyhQ+Q9vaMObEYuScd3Om6L9WUK8rWPNew3CJWsoX/8LSQJjmnB77d2g2pCz9b54XO1GPga
8bgl0tsiibv274043ira8yw4yj7EPIXlSeobUQkiKXvRr5rN0b50HKpE9Qb1dISrAejpsXURyEd6
ev86PVtt9CsFTPkmQ1V526ZmeLUTXXvwr0njTrv6UfgIa3097wDeYnmKPZA5OSfk6M8z95NoTuJC
WsoxSHx9HpNj15V4KpYki93KNpiWW1iDjq78HaZ+/NFH6mov1xd8vtZRCs/z3BDI7t/NRcanchc6
9Mlu4CeVAyyflAuufDJjjDqZNEBAQTQXxVr/yzg1LlwZtohdJKxXGiAneUYS74T0UjFv4h6lOfP7
pTF8ZlKE42fKgFjgk8+rzHVJjtTSqrW0zT5cdQ2wZwqpkaJUv/PD1IA7znEEoXjH7N+1RLQwsHLb
NpiNdSrSOFlAeF6EhJwDto01cGovluem2jPvkBhkkmtpuA5DgpODdXgi3zdcgF+IuNFx44qr0F7J
FOn6wRN50fgwytFHO0FMITc9BhT14kavfJQHaDoEdFhrR7CzeolTuthdpa9jAhKN54OY/BBplKIU
gDFz3zUYQ+Y7ZQ933hX8L/WMiPxWscYN4lwps8I6fboZl7T7NEI6ZzFjIPky190C3VpX0VmRLmMU
1nUSYNBFhSg0LlXlMK5pzFjBH9puXhPRbIlSbHqPNC5XGx408Nf3ks/iwNkOXMkcMja7uSP7CW34
PLRgmVOnyhuD3afps6N3uboofwgZz9WJpL1z7Y0Dsgmp25l0QG9//Qhr8iUnKrkkFS/9KI5n8i90
VIYDXyCexCTutvc0SEkFmW+dEjY17gs8j7wRNS1Jzk7fTZJhWzY/5hoeTPgfeTin41hmHrdgX7GT
LnPHaeEU2Zv88wUHTXQewlubN431kk0CDxifGVRjg0dUajj0jt01VKqvMYquQFCxjtWD438IB8Il
S4+ZuNr8xPrK+nYSyDBDEz8KhJ2VXAp4SbOhoiJDbr3NphmQxW331LqycM4xOuNVX+rcfO0ipRRu
lEQSOIqOQ2MiuU2EB5OEAj2zOh9owJWtWSxL03lvQDratnB3WmtrnpSM836I936q/YVbrRI/1dfq
X65eVQ5dWpARd1ccAEZPObJ3KGIlewmguTsybDZXCiPhvWn2lzLZmhvsix+sa3eISItm+rxvdplc
peSFLXe74Q5/++FA90BvqRn1UT9FOIoqyEGf0T/m7G/y1GrD9/IMrypnQt2STfnNLTLvwwGyFUfo
cm0DKy0lcSNm0H4/WW2rYDQ3ayvlvaZ9ypkqzBEf2SnKHIUbsNRDdrtnlctB2mlip0cRdY5Doox1
10nLAcCYihts2PwuXytK4Cpe39ZtHLbxwwzybN+8qhZC5Dw8+twYTrXaTPhSncCTzm7grMPS7n6G
i6lCAtnNL1X3CqTgamt3YQV3meWwlA/7lF7VTLZlgiq2xNfh+sBMgZUx3XDx4hxTYT++Gvk88YBI
8cpNLInXwW9XGolnSj8RhhVbKAEf5udp1MUE5OLhyHH0eeWHHEZ85GBe6rWxA4BgU43ri04Co+jb
gm5gpIqvqM3yA25Oy4NBp2q7oRbm5A7VY5aDyCfF+6g5jd6lFu3EC66TfUpUbrIjfgYU3LJy25e5
Uu5AkfMPMyV8qDT2nm+cuEH+ExOAPDtWBYfogXzuU2XgyTln11fMo3h/fncnrf0A5Zda1z+fZ/PR
BKNhKeNjOV0U0jkzEq7TWnOdRQiGn6UJpUTTs/bIPNiCP5FYQ/R+Ab2y7R3PBiYYTtGkiTTVZl2k
kqPi0y/5/hdWX/WYqMUU3PSPVtIoQzZdrtsAEkb37gtiAeTqgp7Sli1hl47H46VooJ5NNKMsI9vZ
cPIZcWT/lPqnciLc/DDhvuJEKQ1MxGQf3/sAJYP0uHR1Okl/29vsBf3ecPJoC6vutD3S4MQuWfkf
7e20LWXn+2oFcOcT6Hg75ZLzC3yorFOAM+5I5UAfwY0TnWV8uRzKfLnIkxs2AYyHZUYDbvfgByKj
2b9TCJtzR8k3Qf86/x4iNG5L41HuP6ZzsZy9JLbEDIQPKH9uFRX6cI/tz0cz+dJPEq9813wV3ftN
t4ht9WOZWZ37bUz7QztbedMQHO630RzLFb2ba/eu6yhXgfXeXVx0XmlacOvQeKOMTkfi2NS6RQZs
BYk3b9wYwDU55DcJ7HBF+HEF78YnH1ilpYE7Wfo3FdjlEaa73aTnAJWh/fSADcedztLjMMk08L+c
0Zi5HvK84D6FJYSXeAzNgz6TTmySRRVQPlpM/hxOkkDqegy1dernUwbc2lJTcL8FYfkdYQfsdI3j
5bZx8yNMTpPQnel3bL4rtHPAwRU081vJuRQCgqErvuR9LnLCUUUjzd2XwqC1eTpe8pRcAirzCski
k9MnegwWUILYzEApuGNr7QhhMOLQKph2LtuJmU2O5s+flrkEbcU78Qwz/yjJqkKjs6Ml2qCGKyvJ
e4pABaIuZ6EHzhmmlr7Q7/2eff4RdcbUA3w24L9l+UjryofnAfrIR3lxf6zkuRYfkzIXJV67tpse
DOhb0SSUKCt4i0BNcmbKMZJlZIzVYofXhC/p2Z4tBPlHIlvJkQBQS29eu+dg7uLjOnxn7Iduu9IG
UyVxyaHKj+KAmdjThQTp1gdzX/muXJC3crKHfZQdWjASZhSXsXtLl5AYFLAwGdFr+oOfAHqLK930
nHRGpUVJXeH51Qe3/ptHvmM5saZ3bS7ozNLH/16ZV3OZg+GwdGVTWRAgaRi9OoQi082lW7MDH9Yw
EVvnlJljhmt+PCO/ASN3xJKozcNrWvDp6ey09/3luXdw3yIS/OHV/DgK+yUP9EjRJ+9g8z2Tsvnl
2oFM1GHlOW44nxpTZYXHQ1B7mZ+Op8oaelfH6Q9sJbPSU8fKZOuPsip6XgEZwesPm9E3qTuopLRx
cztzk9bAN9KiP5ex8NbV+1u3K4vSYvUkik+wZwO1gZWJvMDtduEPT3wKUb23gGAeNFcoe2L2fffN
XQH0Cws28bsFYNsbmVwlbZY/wnXWkTI0/hkhxyXod+wsTj5ce7/dJcrKNcEUBuCv4e9uYYV2wsBq
DxG0tIE6iLCzJgIU0zahtwuqtO61f4yaBky03mKY5YvrCnu80+XZE6vGIa/sIpkuOCH4TjpZrCpk
K72muPMLJbXNhofdnG7ZfMWqM2buQRXNLK/KSN1EdYe+OMMcvEfd4o9gsRGzYSQPcboOohS1GniK
DAqzUT/rmzvUW0mETNvarUlc4ifCEuS8g1Tz+n3/Ivd3xaKD1+m8zejWBZYG+I1Q7xx1l/czScER
BfsktXKKd0yUKQUfIDC9WTRxa4fhhq/KLBtg6HUvAttlfNM28wCmJvBF6pG2W374ONqJlm+Bl0RC
SAXpfP6AkyOjR7eOpAS58Rl0Wd54ct+LdIgYvxPL+fRJLlxSJmcMSSvyAFJ/obGteC4d0pzohkw7
D18JTm/kYIpK7J1v4Lou/QnvUhOOB26DXDM13vwFKEAtn3F15QRMqtIrSzxkogz5wohIff7vI/ip
qJzGLm55gNICvj5xw7WniR8RNVP3t0w/2PQvKi0yiXwnBRCV9kBvfHKNhJP4DONS7xEU3lumq7oT
apRoTktbLxUQK9eTc+poKNkdDs1rstpH2YcnlLWYz+zzNnzfSo45mvJqJbV/7TfcuYLI/IMuoz//
pew30tlZ5M1n15vY95BkjUC9oSro6uw4VJ/6AZI2eh+xOjb07e1TWUGmcQwhi7J0lRBCmNrOOSVG
aWs06Q6/33moKUewxBlf3EjEUNaECXplXktD0HKb11o5tALQKUXn2ZzKnUFeiJxLbWiB0I7SihIz
0dsDywSgIRwXueJ4y//6O03ZAZe9sx7JDSV3u8BQnVx0rPez/B8Uvk6k0YAPmMzwrL8utnzB2huQ
Zg7nuu1b+6m08v1BfuX0VbOljQQCcNaKNLOrZ4TWceFxdbh1gZxo514GiultrIJArJDIBhgLD4J3
B/PpdViABraiNOBGNLrJ8wsIGQb1t1XvNwnv8kUKf33DkSDc0JCJpi8Ewpkw85M20SX8Xw/R1b7D
pv3G5obxmVt5Jge5a24bye5Fx4NtM3S3voVD7rqk1kiaXfp+TglF9x50sGWQVIFmltXAZzS5ib4Q
HxIXXi6WZmt3/y51+XmU28INHxa8PFG8PYYRAn/+/pw4Pr2Z1EFLlvpBB/CJXubdXLz4Jwf/UkHV
XvlAVfEJqt/ZCYhVK07h+ycNDv0LHsRdu0cf292FmQSP/GV9mhbxRXUTMfS4SGS8c7Z8Xv8ppd2j
7Sw+JIJK4Dq8rx4dtclgRf2uGaTdLg2jcWpLn79pGwV1DYLyZbaUaGJRZTVcn9k/lO25XnxiwU0b
34jvluT8+wrezIggd70WvAWybhu0LGPhOiizhF9FPLXPqKuyvagELTXUDkQta9ULCKePJdNa9Xil
9BIUiofayV45CEJfeWRSsbfUXizgpItTfdb8/JQuXzTURsAAbdCaYjpp49hJXSNkLUxTXbhXK3li
BVGy1LjmX7FnRZp200wjAmn5Jm++pjruwlp+m2hGMLHeewWweOnSaBIydbCqnfkdp/P+CFVvcwV7
ggoD/kCvMkfdsIGJVgWyL7/YTlshr9YEjYE7Iq9nof/EtphBYNdXoHcEPfmINgCscramWpbyXz73
PZgvktY3gm5QDUatTLtY96z92Czs8+MmZJOXxCk0ICt76zQdTF3NhOZdKF40kmyx9aoArT6L1OBO
vlUEq1vEk4tKWtilfCEXznxyF4MvABJlDTWMD+uzSBywOv+JF78VVt3xDpuZFRGGAhXDdYTQ8j6u
ok8MvYyfKqH/wQvnyfddE70PNJInEKIKqZkBfIoUuUfqbcAl/+dkCCzqYxVck1oXIoQanGRfrGqX
Jf83k1lzR+k4seyqyq0ClHRVhl73834vzG5gAYURXB1lI/SLNhSUpmnkuucL9qZDoRcuPMsGKgfU
85fSuXek6gjx9QhaTU23SjYx7UGiUNSyLQyLoB97zm8tw43NDBQ0pHoPaOwr9hj2PgzBPirDqSl6
Lq1iN/ebVP2nnjR3Rhtw0uabTEOxr6FBfM6vJDAiZd3GVZkAHOF5AGW+Jg1IKhbZtEn7JqZv3o3n
PLmp2aEBP4JdP7lX3CKE/E/I3OsOpoRAEmR2/aOjyPeq98fg3yyUx+JWW7xGeJqo9fd3s1a8ROht
tWLD3kfuHFb9G6upN/pGLW7PkyecS0c2KjO1PFqF1VkFvoj8UaFtkImjprFFO5ft+L8nLf9uvQSH
0/pEyHeGz1fdKPsYopWy3EsipcGL0B33BPB8jqESci7xkqRf2khr0EYJO0U6eSA6Hu1DG0sNT1yL
P23RctWimVAa0oPJ8tlM0DzpvWREqrayxUtBE6YqbsYI9R/j7SVNH6e7dEcYu+MQUIsMGM89QTmu
V1kMC2cc34k8rhy52EkLHXtEKddXi3zOs4f/IHQPh79ODx7hE25A7gva/AyGaR9wpzlrMFSSkK3X
ZmDeT065oc1ZeDGG8oqISJTuWu+iSsi2X3I4IXuJsgtW5yRrC++zOzpbYIEc0FcnBIumSBL57uW+
dTuhRLA1VSaR+DHht/TrLRpr7Eqi0qubgID/6ukX6qKmR84Ek6YzBr2EbeKm/NKyEtYBF+toN+lI
iWeL4xnln5yxxyGbrayEmvsdMnlND43MowlzKNVdp6a3ePwL9HMbrILAU7vT8zq0Jzo/eMgZYlPH
R/6/yZHbUr/15pS1pbZXVXekifLS9qy1FXgrVGo19HVGFMHgl/BmLtlDT3YTKDPczq7MKYhInWQ0
3/sGUf0yZ691Uc4/3Ciz3w8KKGSoENEUBiri56XZD7Y/BgFCcmbDYBXrEgK8+n+h7GADAGZivM9L
61glnk2fW9wQFqccMSi/w6e1dDGe5igfF+2j7w4L/Q4u40YB6Q3wDGrDYUHv/4cydVeDNocVHKVF
DZNwMUpc8KCVHVqOiRgPTrGsMXk30UjcNyhf+8hqUwV6pjvZ9zdZxwGu2LTsJbpbTo9KKyHoMdWl
NCaV1L+r3IVyrlZ0MYnBhtoXMeSvHHguot0zGoMdMXMvuqb35XCM/REpQ4TBCPaIOySKfdLZdUYZ
lyYfh1GWZSoMB0lnqMEVAwmXlZiW58ww4Pn5kykPTqKfmgdOFiK1YXn3TIBx8ZVnvapEZAOvstr4
ZRYPN1+L2BjWVWXSuFfsnm5N5pnjWOIB2lDcHmEfX9A+CjvMwV+iPKVZTS8P9JNA6thhCZ9eQOm1
tGFC/dEdRcZeTtWXPBsuQcYzXOi7I443l4g4sCC4uHfbdPN/YrbjjPuB5xvxA5TehKpYXK34V7n5
ATeacaAuNYi+ht1YRQQH1rDyXAwcoWPqCS94meGKg2u2I833uIetEsMvShu5DRmOgKESsElaZILF
royNwtO0mxFzG0t3tDLgXWRx5VgHLbySlZYbOkCG5Vvb/2Jsi2+/UPYDJyykcWmdgnIVrEvcLD/F
Fr0n4/aA5dzEbam48xoKpEcqeVooFKaHDdKL3lGm6oJxs9/Z3OGsaKV9ufxoGP8Gx6Svm59NJf55
NJKDB3juAVzVCd+jWTjpRrlftbzC6KIBtKApfwOJlzSa9eHZDjGbP7hHqOJ2rJtgYsPgrCPCKKG/
Al8Sgv21kThdmeVYnDOnWMxB/wSrr1s6WXb1pIQLEXMZdrHksAXq4ha/WNnaGfT4D0mnx8K0O7sS
MGvH5ZLqNvDcTII38/QsPNNHePoPLkBGaWuoxi1FQCKeIo7Sjv8nhCZeFRKO2e12E3pOxJj9p56W
IdhKdq8tOIKUuDCd7eoLFbQMLDedB8mf09Z6n1+akEemXt9yDmuTdat1lBmcK4M4NA736ckI9ykS
XhmadwxhkUQNKC1HiYoec/nz7WdG32CyWWbBa25MLF+pWizeIT6zMAzWOAEyMXGC8UEdHJIShfUQ
WzI644h4T3XG3fosiU/BKFQ7by79Yw4i6UBMPM7Dd8Egwq0aOPM+w44jqBkCXsnl5UR6BWkZB53X
vwgB0HAZy8TzHjKQNN0/jgM4T4xSrgIdxEi7TPmenFw6AUS+QP9+JduaO8fW2AQsV4O5AHk1onfi
3kiXBim6UGorl2LH7nt383Lt0MjcyMPgmLZBZ7dWlqjbvxsRLCmjHhopfioLmxwwWXIYiGfz9exA
uwBadNYLx5SOBfQjfI0l0/Nz55IHGkr3Uu5rogVKlWdQOY1NLaqSxxwI3vPe/JA4Hu4+oQ0a9SFU
+24vFOrMpyrRR0WZEsvrBzCyeSbBVPOUCYzCAROOyQHxk6eUEhwpyAALmkKONI4ohAmcz7Bnz6OF
EcfUqGY3fQOE0i5ImVAevZhcf+PsCmKybkPYC3obT0ln8vkNTFZ+YbQdF+nHMCtsKBb626RVbSfq
aDBu419FOfiSVIWawpQeFjNmMzVLkE3fdQWzqw0pda7bWB3ISMEndCo5vmQKeimUESx8jJYo9+BY
jgRVcdFFWVoQTNYg4zu4xe2namF1XRUfOm+2MJMgkW23jGRKoy4pmwdN6pOMkOWljzZ2uIdEYSGC
SP3lyb5npRFa6iA8hGETOIy1+FWA7UyfeZcKviqWyCS0RhiyHHD1OJwpi5F2a80WcU21c+wHtsrV
cTOjTPUdwEeRoTovyo44NRHhNs9DcDtlmzpktftKE2W6yiCYqbOOonB14hRtTA6T9aOi7+oBrvbt
cYr3ngi7mJgN1iM8KEBI334NM+epB3rFQCrecWiRI7TnBrFM5nn4Jditms5ZuupdASPsGizLPEm9
aJqhHUJSX4gRtVaw5roblj4V6YBF+hXGI5l8s/VyhaPB75Kwsoqj+OyMvapdE8o2pU2zynlL/5mn
G+pzeM5WvWTl1kelUQQt+PMJS3upxXbSUDPFsFzPNc5mwWhX2AqhHMoI+LjIznKx7k9PxRFwOlGR
NvvPttUTZplglw4i2ybFpu086CPCPck01cZeOgyESeG3R2j68r/1nSebTRApOc0gfWohbhSwKfje
e+/fyzW7mbpfVrGxk/JDNfW928kMxLjI0pf3ofHLp0u8+r9Wu+l80kFcHKXXSxn4d6rFwYRCegy3
J3HtyHTzjqcMAp6NLsagnySg+ffhIFvoHXgGygoiRRFf4St0DV7XkOMGdQL9dAhdIj7qb3HymYzQ
icQ86faCrywEuKl55y6iC/iiWNYEdgpIuQDR4eVUGf+PW5N4i0RAxwHqNTMDi3NlsPgtOv7iqaD5
LCUt/K1Tx8geY6ZjmI0/+8XS02FeB+FM69TPmFdi2Uif2cUDqulk8CO1aVOLKoaFc04Krp63wNr+
Bl9BDVPbVWqbDnICjDlRp68ExA/TbSRm+vR09tKVUgChml9ntPaesHlpo62KHiBZm/z+aSlIfrRV
VNFIdtRlMTY0BrfyaCWjCPJfv1VzgE9izqEqwDA9mnRdS7zL+JR0M24auRwdx8tsGdOoFhk6ye1l
/X9DLh+Eo6wlsmnL5bmX+G44gFHlwaQXCCnJFhCsQ8rzKR+nh4JHGufLXrAP6QaDXXYi7cvJZ+7q
t7DDNtNqVx9yn8dJbKfCqktQgJDTUuL6e3sgxNlcVvxfibVGlMi7GWfkXz/HdaMipEMBizImDneU
DYIzYW5ApPuMwHFw0cxefIQIA6/9TPVP/4zTzZIMHn18GT58CwcN5q9k7TmCNUWfrui5Qqvx24OJ
BmoXeIPq5/CX0c9EhoVV/dAZsgXOaVvC9xq7rOuYDErUcfDMB6myC1glWLo1I7luzp3hf5QxiTFj
RR7BlQjuUsHde8Fp8hz5/gy7iTo3p320eEiYDV+sNxBCQBqrIy/Fo0WQn1ukPPtQjbyWYd8g+P+x
/OFw4/BEkh2ALbVN07wlTMMPUIltK9eoIXsSqrCy4mgYVLvWYDsekxwPZ8sCLlPbXASlDRkR5pNs
/V6aAsOW0MMMp0PmwE5XEwq6davM8O2slYd8Xa1xo5k+ErkhflrngqMtw/BqBW+ddlZE6OYPrTpe
h4YHvQt4PW//DQ/V8P1jokA5JqkTK3K9os9FMaeKyk8wlultRy7+TF/928NnqhYiVErOn2Ewt2kc
Yrbs7ZMnanp6sfI0ycTujIouA9QmzrKgoQfKk83V7XaQgVHgFZZChR7GBOrQ+/Rn8yjFZsctGDfP
oQjI5SvTMtvqvDUTYd9eKKZTRc0vpke7zQCn3Ju3t/okrN0qRA0d0fDNRZ8sIqBW8SCafqPcF94L
X+cLHclCJOYKE1Mr0fZsB5Zeh8N4V6l6xjSbS+9xLi5Lo0vd+RHYIp7R5yU52Ya2IiX6m9AlNLcs
f+fD+6i9C+uD8t39d+yibGYzKnMGAz3/t5iG5/UmyLAZEXiLlqRx9cPRxQowclRC3kzxnnQRTz1x
lALoz+dVWFJDlZJEoxsGVzPXhrMfSPeH+qHnvUydDN/cXabA5t3cpT4YRIkfylF2rRwvUPtfAXcu
Zb25IdQiWAx0FS3PU05+YWVRv6XfboYyHDrMQbu7TmRG8Vi0PZj90IiO6I09fg/SY0voh5JT0GYt
/7+DMAtW6OvEXmWjluQvU9v9fEBreDev+XeaKQAFru5RA4r5Y7pC8UCZCpqFmkCJE0rpjglzl/KS
zI8iQZsEeIezL4/EB11TXbFJbNWKDoAkH4ixWCqlki8aAKn2fjzEIlFZsshHgtRvjGlwR5Fx9hEA
b1oz7b6L02RCxWpS0jE5GSqXXVA4NugG0FZeVm1aKHSch4f6wmUXoImdkGgmDCz62Lnsf4CE+Lnl
Hp/br6SXsECKdmj6DXecXO/6VtqvXRMYsP/oJ14UARU+oCk9r1AE/9Fuj1qDcWGh1CXrUfwEBSFd
tmsc8S4MjvZSF0gaYnAnELn1a/UdTjoqmSSZ9K2uZR7q7ZN+lFs0DPhqbqGFu9zh2pjuc9WTv6ul
3UkIg6JDKtOLcgF+nK7LVsKiHoS2frQlxlSax7QxlkcDX5/wB6FFJZBvBT+5+w/NbjLuc4ObmJIp
EzwQXl4SZdoXR5eOqhRcF3acMYqRVoG0ZvVMB2ycM+iwFCYgkP5wCWJmvgJchOyN0+xdw7tej9h1
T/Kg8J1W/eKUbJ3oCAm3BxsOlfsozKTqNtW85gi4SUWac2PtbveHDq7CQPgVb3WUbUfyB5bV+VG3
WPdMfC1Rz62pcfQQH+CBPn+gPmkpLXzLoy9NZ+zWsOyjW7AdaBJ+EOT6eMd3R2Lp36x8sOaiBc5Q
suse/5Ms1qMXk2XOrfauYkCUPNfF1z6J1SSTR46y/FB3Z0r3kmUIiILD06Uu0uOIYGVaCh7YikdB
2j1WfOxt4SXgHWxmYwhHJGfPZ0PTRvtpI6u/8G5Tm5Pqc1qYp+W5v0F0V83qbk6f5rFN53SHSscZ
LsC5XIGhXKjUqZbPv+L1bee0lpM89cFQIhB9+78oIqG2OlSQiVuLL20m8MgoFgK8euOTY+FAWZ4r
bli88GUj9FQ8ivYCPDijsamfPPHmWMW9sh9kuHanlD/NESD9aF4H9a+4QRTXEwdkpGcEsGwHI/8E
RN+kvjD2gXM1UH4zzHba4fbMa1BaQgQZrjYm4mligLoCViSRGa6R82azl1BL807IiYLuLbsEbAyO
UtcZFMMknD1AIJK/FbHAFpUQUx0uh8iReZR5sf0FHmL2kODEMEFo4RjqL5hPx04E82hGss99buta
5bUyFG7clcalSjaCV16ZM6vPkbGVxeXo9kHU1oSSTN1LER98w00A24SIj7/sCGKJXMcalG9jfjKk
JZG7GNQGR542U8kRP1uOUNhbzeJhYm7eDvrsL2jq/xUGF1xhlEXOvfzz7deKs7o30pVsnRx8Cwh4
h2nZ3gzBTHJV958oolFUCxlH3QpejhF1h5/Yw282zbEydUsvwdujoAa2RtFWQtnf361chUB93+33
N6dRRzW3luQ6KJut6/9B4DgJa2f7/y643citQaRW9E6ZeUResR0RYE0RrO875IhFDqdGMAAUfb5S
85r3siq7ZRB/nB9tz1eQ6HCLkGZblaFySPnEsZRAvgS5C9tJukeHnt62aHXZz86VCN9t/i1J7IK9
tK0ytjcp7U+fGlClC314lFUVIzCjidJNhS3GL0LeC7xp4FEFFDeg0eHCyuBIYfvgUm5aMJf9fF13
wtEpdNX9HGwsINi7FtqH+aCrHOLbnMnj0QBHlVOya7aUbZY3bIhV+jx/tH3TeUMpUgtHPmYbJPpv
u2YRaCl9XxGeZGrge23chHXWvMeVQnvZNwx2aojFalnYoULPQbMkVjNNCCeQ+R2ZngImGc4kpnuM
MYv4ND4bphyvKGIg/vmGp9em27+upZqkLAuwPQDiDHhVe/sMqSpqEksVBw8xuwF/zHdq+5R25/Rp
otVQrrmwfCJ2k16zl6uO6OkQt4IYMQI9gYcXKBiNgM64D+GAKuECg+8uFn89SEu/499MCx4NUX/u
7k/cecul0bTEadqSCwdk8eCJaQbL7Wzp/s2oaG5jzn8+Ugsk4vz0bPZL25uBTp1OXMrp37v2dxfv
NlcjfUd4w5i1o5oXu8IPtWCMlcwBXmOKxTp9EZCQNZuUwgr/b+8FERD4QVbtS3DB/DOovoBA5Hr+
FHCfN2ywyixwTJ5ZPHBqytlvwjBjKMd8Jxhf8C8PkKbpedIOJR2wOOdS5mfmmbFqD8FgkHexVbvg
cUZe21XI46FViK3TgmQVonXYgA3nvRMlVPbeFVb7KIGLttS9cbWKVhYCKZco3k0cRBGQTL9itx08
8mJP65SZ1FD1ID6uMLrsJl9Piq2kgHDtMdwlWlHll5GylIEY6WiXY6oCDNRIqnTKoQz0oS2bz4QX
IFF0HomWfT/kYEulJl6apsn1kUDhp3L5zk6WemgYnWhJRQDbpyJhatLwsjXdEzT2RzHtpzxczA3j
VAE5pI/Mwjrnzz4vlYCDmglcCmvdNv6Mt9MxQXxwnP4HfKo7AoHo0VdvJPUm1os7hZ/jN2n5ShH7
XPWY5+7unNLgUNW+HwSuDA9v/G616DxIffugpkj5N6sNDGsqm57h2jTxrnK3pxRCuclGZ1LjouBY
Hfel7gvHRlvT+2mPgTNX/eYZw22y0ewhyUrGV9kBbCg6qOrylLNlsGv6eQsNh2aHGUH5gR6RlfmT
t5thHxlaEDIZ45MwsqSMEFjd3WnBlDIBSGJBabG4KflUh2H3/0gGYt1HwWmvBiwfh/TWjbyohONx
lUVMYrU/pjj2hmCKvMUeMvQvx3qQNnIk8J7/JG7wQ57/KgybEskAlJsRGfezvHs8uXHW8SZbGSgj
K/rY+1DHAY1Mppt2SXwxffYXnAJqlT8TOzQ/43ZEuU8UfjceiyuGyvWmhcvXGUdNeByi2E3565pV
XO26+SxWtyflldXLw1mcfkqVlwkGrL2q+DgyekiBMQa33uxnrykcFGn9i/RABstK3DTu50lKkN+L
RncwPqDW5RzkgkPDx1uc+kMHKvUePudI+USW4ol2ykrC3f5rrzQ5+dWFkXN3W7DekeWrjce0F+yk
C8N1XOEtVa6zpCyxx+Gi9tOThmU/X4ueH/rGacBpmYKd15oAXj6TOMtlyYUFVOVk3KuDoz4IE2W5
e1WPlLyM6zYlSRsW4PAqjI3av7zPxtLFE/HFVVYItcmAqvupyjI5WRjsCab1yw1/v1L4JZMGAZBj
Q9hQysjmoCoDChVKgAmkOgTAym0Xy8UOWa+6cKIxJY5tKvUit4zE906aT3E5IR3n5Z/dvfxxfGjX
vyBRSvTu1sRCi2VXKkM3T4g8PfcndaRYsx0Ic1tgXA7x/BuWorz2Ni7dLtdQYUBfvMi7kcB13HOA
NDT3DxMzzTBQEMuH1N/YBSrNN70JzQc4sZQLFbkHgy42Z0Nvi5rE4sMigtmSli2nTfIPqWTNvVjE
AWSOftbrywKuoTpXrdLKiEaYbxEz6awDENVuOF9p6QUc4HZX7dvjHnUNSoxVoO7RRjvIPAQojl7s
/Ax47+qjkusCU3bYz84fiyXF/3zWPOPz2NTAx9bHR3dSwkKC2Twlg55a6C9cAQJ/bM+xxlX+bt4p
FRy6pX858by4PR1tLwwyQJn7z7ITxaldcB+Wn6p8XDkxikiVKfuQhP8QaKN6KWiLxcyzvCaeLds0
7VasxsPj9AJ21Hjs/lZa25U+dV9+STRmD8UDpKhDnmD7PcfP7bWowGguq3L9H7UMgCrwdfs+RBnV
1QEXJn0ZQoCz2JzRY+D7V0vkCCHbc1RZSOBF/a2LnQMgsv0SqXqUgSXBsUg2xax2fIr2uFakjcIa
+/qaj8kuDyqDojHfazSKLWfDHC/7zMXwd0L44OSeenYxVW/k3pm78qjVE4vRbBPFRFXrM5hG75g/
AkEcPuQg/CAIVZeb4CsX3cpCq4sV0oazxrE+MvMvdF0MqQWnHXT/SnRA8A/PMp9BevgGMVp2+szG
9AycmrVQ3Y+k0ujMAIonjQHkWEemlERxrYitqHjI0L2JxQMbCXGAKekGdU8+Ffkt6SNMZXncuZLt
xQoLSwPdgT1SBLF+aX/wF97Qo8OxpIeUJUQzuSWpkE+HMMMUx8ALbR1G8N77o5qhyYyOgH2QX8Dk
H46pLZD/rotJL1pK6E90pUKIMr8SZJAPjRqHJYEl3SvXg91EWpmzGT5LrJ4oKsqgsmQ7f+540967
4p+W3KxsOTHFwB26HrtSEQ0FewXQ3DDzgR02MuUT3lO/zZW8n6dEHbJk10Gxo68QunQuKTKOBOb1
zwFg5aTjtdaEqe6UBGzLKXYUrFsShVWWa6ttsRJ5R0Mqb1FDpp6cUKC09ug400+9G1LxV4tm8VGZ
Kv33mj+0u6AlkxThWQ8hZsLpOUivf8OsFcYvnS4c636ce07JyDD8rKpkZ4vudsLBUSy6nw1Xj6eU
9H7nlA1JHNzPQzORYI+F6O5LKc+h5yoFgrQmED8/ORQXddTZ4/FfeYk43EXdVqozRISI70ixjZvD
4/8yIPfnsvTz3Lj+1rb3YgIG13iRbRwM6zLSzSquL2nyML7eGzn2YApxQryXhhMJ1sHIlsl6voyQ
wamcXtChJynXZYhaidLc1bsh6izdy+tTrUJwNwWPfR+WoX06HHMKX/T4tEt8QGRlnqdKf6FpSI0H
Wz0mUGVRFog6EP7vJFTtAkRAdE0S5MfU9zYAQbrT5++Ax/AZv6D8dGhjniaCTxauXYj5rYFpjFl/
ezYfNOBAKP7pwWMtY3czdVJkPNymF1TkPIK2bOchOuOB2+soYaYHzzTK2FZwD6ZiH1pNiIzX7BBN
aSBX6qjQMlolG8VHI8wacHMuNNpyxZ+orWQ9WfOtvq0ddJJaAXA5tkvESRQhryw83tu4Mw2jz4Cr
o6xTziWTzbMEMd7nxpig/gxWL/hKNEr6CCGMvu30YvgPeo2uO0W/IisiUzlmy1AJ8xF1vfh+cJzd
Sn3JnV41nijUAQ7Q8csBczODxE5tSWbYl/tuib4V5ddlYUMoGdhxw6kgnRYm+le+Hh6SShHBTPax
+vz7qgyV8fnpKadksIYhx09xgZFtRvfEp47c1Vm/fUz2B79kP6s9xD24gwitXuweoFBn2kcKIV9o
xwXKGBkw0/AO7yVN02etc0/KF5npdCQ2H76DZpvsDKdeGq5Jdt70JYAyJ6qBTtaTS/4HDJquJSbJ
RsWhY6XIh94bftuQ+9Tz6jCXJgQbcfDj3oBTWruwcmPPcwGfe4ZKZy6o/4TI3Yg5f/0OVFoVg/+d
YgDg+i1jXj/djUnibZ82FSg+N3nS7VIzILNkExDGcCmculjd162D3hQ2JVL59PG8afA6J5+gpsN5
9z2AHpsaNI37sDhZm9bzsbqO1eCO0mcyqH9igqIHlTDhgaS2/1J49uBRBSsTTw+dZ1Q0W5Fkgs1p
WIzZfji4WGR4EsMLKwJ/UGpvQxclVURISaoo0v/317U9rYfF1QEN5WAUiQXRcy1dfZpjSF/K8GEw
NO2vAfjexOEV1KQWqEwxpHAQwzdMAJYuzkarmlSGbSS44I/V50nmM7Y/YSFqAlVyCX9x+48W6nnH
5AfOVQC8AC2yksxGJJF0dtqxdafMjVLqqFUQJTxlUqbc5tl+EMcB4xi71jBdhIOkvsYffRYjr8vH
5ieEWq423d7VzuFmC7El1Rwhxt3+BwHyYPRi6xUpbUUHta3LvTdxA35DP9OY/HnbD7zRaiMye78N
7948X8eBPzSx3x8FPYBKX4shS7f5fx+ERlAvICBcdf8RUIJadRphgQJ9qD40osLeQUH4gBbpTSBr
ZdwZV1UD2OhXU0EfjAuAFw0m0o9ltXo/QqB14KdUVvbN7rBjVZFktB65Bl38Zwy7/f9x0jYFAo48
ijfrvsRBD9jF4+gp/8nl8ucJXVxDBM3ufCuqtz+7icdBXaL6lHISqoKULxCilJoDfDXBXqWKmMJi
ZfkLUyxZ9SHpRoT/bRe+x4+FPHKXjD5aAOQJII6HTJz2KvVDlzYCWhwSsThkdmxMOhlzUEL1mfz/
1N+ROamWVmbFt/JizFLykkjjRglIAItmkNxjObeNrOiw02j36YW3TC1PT9DaXu32r88WIW7/w3UM
W3XvF1ZaFk1vEqckIMUcpUjZGEbD4iLYfr182EL60qGOHgg/XyyTSWqoOYCoFZ/JuwiNJI0iCrxC
tVNM44ZAILIlecCSp0BwjwEQaLZ8XDW3ZLzkqH0hV2W54kBJTrqpq5mHOwjPcjV2p+idCQkr9/NN
VzuHMntdngDuPOSw+4VYlggeieuyW3RvjJuTkQJON8WqjGtdXN+9FTzT0tTqW4phoaFyl6cQfXae
BgAzYlMvCNxyIJP9CNsYNciGw28iFNZ7jY9hptkBvvWt7m/T4cSTJdZhKuKjuLgevrDgZEci+Vev
SDqXBqdqqHdV/B7kZpUNT/wveNQwnWU1ZMltDy0aKdZMmCD8gg1wh5cNgzWRIqZ4hEqPPnRlIQWI
A4J2aRcWrRETF+FrySDHwqzN5EBUlgasMWKXeaK8x+nh9zXqq8s5W1jI5yy56tU0Rgq0c4IrwWmJ
oUJA5ye8RedcZbGmmh2b5JCXQ28EFjghITNS6VmJnufmult3TmmX2FYJRbXazVNQ/U9Ex4VS4hzD
DjZPRvBPFUvje1plx7D3kRZNExswLMDBkCKc1NGJ7T1l+Dwgszxwh26pA1vEHNHqGwfJPAM9jRAz
QRNPQPZX2e/G6drt5CWS2VykDmZtXjGcb1NhtxB6bseeVZZtctx/2PbRJlQ23c53kO3Yya6QViqt
kWwo0hJalmvuBM2w7SAYA16i0qKc52aa5VuSf7d8udaej39cr4uZK7MmJPQ83+BVdWvraSN0VYsl
xpjmY0hcF4p3SyRgFMxlZhMwGqlqRVmi+u+K9v6GJypgLQYqAWuENFCRHccAWHGe5avPnQFhEu1I
vIVCYDY6o8zvjGUdP6/XY6qXQX03NhkaHWIK0LvOREuOLAYBlZyVOgPLJZcnoGdbV22lWqIiA+mj
QP676MaJxCsEDMlNJM71LjGoLqg6C/sbeWdSu38C4JHmiH3m/BP96hRVl6Jpd8rvujn5agO/pown
TRl6CKN2bY9VfHlwcD6grkwKOWzFfUbHO98mC6QM7LiJF+NOcTlkeC0vuvhLKxSjfCU0dbGmdRgX
MLXIL05La57YTNzG0FZdBJcr92zjyExJFJy5aWJL+D5X1ckJZmQQrKntjNNJonJehlEmwO4WIcYc
UzaJCTBUcIlw6crEGHRoTanT48ZwBD+zFypskGU4D0QcAixzOWtApeLLAXCSnqB9WLTqbJsDfe53
Sz4P8QDQX/Nc2d+kt3scn7gTQg5EUXF1AFxudgMzlZvFE0QIHMvSUm6yaC6exl9GmGAmxGeiJXjF
vk8dZd58vsFWp93fodSpg3mISz1Biq6h4BrOVAKKTMvRu8L3YTdWfaBj+xwP/rUqD1r3Qp3NPQCS
fh/Bhbskv17hxHYkCVJmznSIOp97bnWRdpVBlx+xIg34jvz1ZIxrO4uxloqzVOBAly9wT3ab4/sb
SWj0njOl0kknK0OLgn2V0vV/hmaHha61744CoDEeEL54l9LNgvCfF3N3sTG3w/NsnsFAeOXhBcvh
Gd5yYiBrOtuMRytv8mqicJYr7iBzB+ztFLrBIQSxFLTdixOcdDZbOSWP5sPcfZmfHMBgsMxBpcV2
w/CFCMPMLG2ltuno0sLu6P7n7XvI8Mvveh8jwv5Q0FSP4Je7jh4exK1U7pRbRCIxrEEjzj2jW1hv
lL6WluN7Hohf4pMqwMtsnPlnhdurZpQObNy0gCMDKQ4h4kKZCX6u8jtEZ8u+qucjIHA/wqP9WO/c
ICgP/iHUfp4ntc0KgP3KvAkdlQpfkVqZb6rXm1Ttw/WK41wIlZ2hht/v+FHFJ754DtntxViJJMCb
qcpJc1puEpMQB3+BSbprbYe/LUfrYZjqX0rKKf0yCTVOGsNBUpso0s04i8zCSDYzpT6QsPV11X5P
34AGHVI5hlxL3wpL99jte9D+1rfpXRsZNqfG+IXL4lbLPu5nPKw4O1Two3wmKjLVS0e9SLLI0QOw
+cdvLgvwothkWRhMz49FjoMcR6hf8TkotAACzFPd2WTzApsMtgqtWeDC+dVB4Blp4zrblN6reyK5
3LncgSIPCg8RfF3Sb/SQ5MtGe1qS6mtDRJc59yq1afhhptxQuQnPPihsVwNT76StIIBhXxXt58HJ
RPZE1dscWxoFOVv7+Dl60AbmYQPV8a5RarGzeqELgngTALMapKNuGg+lA3uCbaj57JhDvLd9tzF8
hE+DM71X2KEro33oHHfhQRaG2ryOBkpoEHd++syfdAEGqkOcrDzCni7IkSmdy2PoKBlybd7Q3AXA
V7dKXOkCbcyzETi4XPP2onHiSVUaZmuTRCXVNFjQgDBJnbxNeeU2Z15FrUHbPpYX8RiS8xrKxXoh
aH7RMdrNN4IEzlFX/bzac7NWbKkzXcc7H4gVW463XMLLtLwy3WQ4QtN/PqqNoQJLrgmbPyUA4FOs
fwiwPgl1nMHKfpDgN2j/aFhDctdWkoE3LESIq0k0FuA5s3mACtFmlkU+m8jfMxpt6VX5heeDy4yj
X5xAYCnRfu4Zcv6nHq34ivCuDAG4R88u0LXuiYGOwl18hsmBHm/ZQP0brfGsNlxmqfDpaPk8/BPs
W5MV8rZCD/+hpXPZDnddhaHKAFSDWpVlOO9kNBbGPLlEvgN6LcEru98cZ2GmJpKNKGBeImxU+1Fx
YCM0T+QMlsf4zjDJR3wbXpVCNZcGjU73f3+g2kVDHnv4iUdyz92Y3VNIO7ALmSChQntt1tdetQ7Z
RFggf8URfFoSr58Gr8oN13vGGa6l1xLo7YCh+H8f/7Ju/RdLgRMvKGAyg0kKcFC8nMYXHPvvBqZw
JyS/PoE7N415ZCU19I1ibLsc/2PeElirtZDsRMICRqc2GbCFH6qIwj7NpKFRNcJA4y+0oKklP7dh
bEAQjH2hEsuMK0pIt/nuW2+pNy9dwIKgNfRiEvqgLAjcwD2mrc8p3pdptsQBGASpdBfhC0NMQ+vP
KcHksNv330VgNPzwBczwBQBRldgDx631aVd+9f6e6nySPEi86QPv+3da+7atYSIsyBOS6bQPiILQ
xlqj4AaWm3v7fYu/fO1Yfx7rnceWLvR1PKmeCuCVJSOXJbhJDPWl/oMUpTbbCGXLklGFRz6AIpeC
RWAiFzgS1rEaFwHdfCKwXL7nLLf7fjJotj0iQl+C8ihs4s3cBfmCQAK39gpkAx5ns3e5bGLm6Pnw
eogkzTsEeV0WIYcr7hBIwvey3GnETQ4C7jmgc0ILv8Qj9rTHqwV3LEx+PGHk1l/KlQd52ckDd1DD
e/Wqt1K6H3ZblwK2hSEC2nKfOiG00eRogBlGMHW8ZD7bek27oaSBAtzK7V9oIvTRqRc1NwbbAmFT
AQ0eOWV/vcM7UL3DNrNfVeRMClPaZtvVTjg1RP/KtLTJa88dcjpQAjhiSYbBZqKraC4o6vBa+Pml
61AwjpwESz8Tm9o9DKA9RBOWxV5fnVFAitkt8jz2zBPifKBASR49WeEk7+V3iX1nOctn/LGGr1Pg
CRNDZaks3MkAj4MIyKsRoznXWHNmlZ5YkxHJlGapVnxd3FCQzo26atEVDlW2EPwcshsTAteFju80
5k9O2Ee1d92OxkBl3sSmr/DSHQyxKHtwuiFz3Yf7IHDKD7ZbwMQcRoHEkrE2VQSUXdvxO6Lv5zFO
fQF+xVYJQIWPwvwNphlD8H6NLEjIma5zF86luvTD2DROIKC7MYqwxGjXB5GU8uMIZdfIdysGK/TK
R/VTb4ZbmkeDiMJ5QbSzQmoiMvbQf1LD4cOol/C8jKZuLocNAV5Zy4QV9AU225fCu0w9grawf5jT
ioD/yeh6IGih+66glYVAZAVeAxn0ZBTXD6WN8AbBqW39fZ5KiI6y1MmaBBzQSTMN0A1UD1f4mvbw
g0YB/O5aTebwww7SjX7+Dbiy78flljQ6sClUfW+Jbad0lOQ/5rpEz9XwXFppnkjLtJSK3+OaDcaJ
sNGRQ6MnAqMz1y95j9o5FkGof1SWHEVSV5tNo9/ZDCskvYT3uJ6/vEFlrDaV2CjbuHTkDdxuqVFD
9fENOjlrHEsn+x9lalWYsRoIXng2bNNhvnlDiK1o+chDj16bVON79ejVJ0FZ2INnMB0X3lYsXM9G
0Vsy2FnJqb7fEE2xgx8KKz7cpp7PjVOsKa/523f0Lo0YMitEX/lB1gKpTZp0EdLnLRk3s36Aw5Af
6tUWWKxm+nT4TSBobjcYLsS6o3giAUbNRC52RyeJPr0yfRIk1mH+2QR3ttBALB697j2IvyTk5PUA
De0eWA3n0MckTCfF7vDRaobv97kONQKrfnmYluNSLL/SkjxrL4PEcEYsD5sSXlQQWVVtDErrbBfN
7GaqpRkeClgcUNwrwpsZRymt5Lc3vffbx9axBWFhm/dMrqNBObvjGcK+Y1o4WewA9TUwBv58SYzo
zfehuZl2ruZf5Eq+23LEiPLLeWqRdDyWPylE/vSYcSgmX5qrZbtm2SwwpoLrg+i2G3e0fqZreXCa
/JXiF6OvYSkPaGkd9HlJ4MkA4R7UGCnCsm6DWKXh6dUGVoFyCyyQvEe4K3xFNr98O09qaVbq+Cm7
ax/tjPpZYSyfwG12hSmMJN7rKfNiyCGXG2LJ8AdaBHMeYGkknDN/h3MU0fuGQopyhcvkBsVKv2Hd
ghFxEzGI9ROOqxqcM2cnufeGrv9RZ9Qrzv6+PB8AosKNxabpJpCUe4qoPGoHEV5oHiWViIxBbxVl
JjKVjg1+RWwmvFHfqIFyeWgAcoOSlaSKN/2jgVn/eKeqFC0vzjN7Uj1HlLTByHJqElJYJvgNVoq+
W7Nc85bIonGF0dnBNUOpvFm3TI0J9bK8hysNQvtI25U4met3Xc0DsQ14cPCGWIjAPTRdCZMUW/mh
alk08NtW4+h3jJ2GSJjV8fGBkLRZnpCpy29msqgrJEOwkrMLiUr+LTLs7oabVKi8PVfEQiBy6rUZ
6iVOYNt7Hx09sLG59u+g+rNwzwte0p0KaMOvH0d5meHH7lAxkA4vfbKb7lvkMz58Q91GOa2j7JV1
Chn8EFIr+A7RsIz5E+lgGRI43aHxwU7vU+yumM8tOrPyB+Q6qWjIQdV4n/4cC6FcTFDklGiYzeyQ
6qDENdCa6u9u1g4j0sGis3aXkqKO9rNr/GV+yOtOkOZbXutsf3frTS8e30fBZF0nx5irZpiTf5/5
BAaZmKDl+N48o82TKvhJjiDLPATcLYGnbiveMIiPtzI6wnuIrUJxtZmFf8mjcl17uIxVC6IYozb9
9kJQsjd7jnG+90vQzHNCoDYrhxpg+wUm0rTCoBvAAwk8tAHB9O3pmlgE++DmYJzGYDfNH/pb0Kvy
XnYUn2mPn+EMwjkm2uvbuUAxV4Oz+XL4nmaJV0iR6GdZzbb2QZgEQZiAjPGHcdHiGevN46f5KEtA
JfNr6VTQ4KULMk4Mko0Xi5kAXrc3wG9+9QmRqDPwaI0ipFDjYxHAqH1NxPHeQwf19nto+8YMM12g
V5ktmtBUM3RtdZz3LynLbIC3x8IZzpTnEo7XMhnaS3f+5HfStLs2K/CJpRGNrwj6e3evzod3AibW
BdEduuuTjp4YmICa/udntlXZIiZD7yM/Gpr/NqI81Tgj+qghfF24KlXxJqQ5Z6fYp3pD/JwB27E9
CgqxTfWhXiUJ5pDp496nSpECELgXpFRTxsgWqaJP4YmA2HMT7VbYLZz4XP8J6iACyJeuPaAqNjeG
FXLIV5VS78CIlyV1bShDWWI6fzpS5YuCQiHXk5AkARXMJigYuDNu41EDGt3Q5ldoL7Z5ktcADDTV
iXBCJPAxZldxjIdraSLnnVN+wHk+uDl700XO7C1xbzdUcoK78Nh5gsbOXRO7t7QuUeLPIFa+Wrxq
mJTXn5gyHD4o5aPyIYVXpIj3+j2Z59CpAD0dKgpl0kNFAGdKpjSka3ZWKvLv2jP0R5Pa7iRHJg4V
O5TZD/AwqsIR+wDd8T6CAn2KuA+GLOqrB5QZcHIlP2pj66JKj/ql+dtKXcrtYjS9XiwDZ+xs4Yd6
vEajkJEKtwuwg4ATtAgjXjWX1fk782AiZgVmiCnhqQkn8YmIx91qx7PRi0tddjG7d7Rq3RQwDCUy
1jVNTjEpOTaLv1eIeS9XPmMW/AMZxcF2PSqK8hlnH13JpqbHwjZOFF22Bkbb9Q2X3eO9UPW9xyxF
r1PlhwUXt7xb1H3rRwPZbCZy4JRNgvAeFe6ReVwLYundk5E+agbNUq6n966cSa+dEYv5uwQKTRG5
b3FJx1u6zqlp68HdMcwlfFespfhunL01nq3Yaa7oSkn8UoocrGINw4QhJGmCURM+gqcIRYmWCS5t
hUbaqNMWC2XeMr5ZVrSQ7Vdl6A2llkx/bKX84Ribdt0zYi6nGR2ytAJ95UwTeYPyyDgct2NqZc1j
X36YDfRdcn3JqKKxSOVeueiSHLIfpk9Bb1kvZRCWfEV6Ki/p00h92CxxJ89yJpRCCTBNFQcuCy2O
dtM/vJX1dJyC3OySIpOcSymYMICmsbw/SzzQXg7OVuAr0/dAXexbIg8aPYRfNUHlGK8rIeq+fE5/
6J0no8A3NHINhaabL0fqamEtck6rqgWfjEX35tzCmN7dBj44Vv0JAiiHo6OK+azdf+ufjAXpbLSo
N0rpsLlQo639mbaGtNe6SetOgvd/PasI8oZi/ja7tfOgXgCXr+FI/811Dn6F2y1DgwZcWd+fVkpO
8vEN55sxWTL3ERDKuirGxt0A8gzYj2sc89fRwXdVqi1NW6bdqb1iFTkPw9onOyYnQH95JW/t9oFj
in1RNxmeM4YUsQ9CMQL9evtz/z/Qh07IjLXGVoJwb2JFbV2gKtuHlUwoSH7qvg/FlujdHgjaPrgW
/jI2NxRoYPqS8iKHyaMGtvKFDIiaLaq9Ip5cfANaaGN5s+P0NA/oPpWYAR5vyC4LctOvJZTup4hY
2jGsCHXw8SUgsWp+3vE1PUWmImIbGT5pnpp1H5iy5H58BXK/5WZe1v8AU5oOMEQvf285F8emM+zQ
P/s+bnYwDbD9/sLQcd81rAy7busE7FEBV3xf8O2jjuCX7tIQbNX8hDsXGNJyBvgVPrxiJRB8kE1M
rIoI+JSj2xRRIggbzrSP03ybjuukvAv17uRLy/M/RyMh09ZsEbfSmr/JyAGb0UKyKwptJuolLoeK
uFcVqQuJm73n5Ld0qurXdSr1fhrvT/ljZBts9/obveaS6FdRNB8Or7v5e7JPvcISw5LXxQORgV2M
j/odrIbMnMYWrpoP0p3he7tQ9SgQBBH1gyORy/eEEieB5f1YwM0IMs6wV6B7SpWP/D6MsFWjkdrt
ajhnyDepiOeH38ZxJTVW7Y3ARdz3ApLvJhTYRCOHjPUpBqYSrdX0bLwJi09k4btPmPZy5InOaemz
1wUqcaH4ihmV1sqNyRIEgcX560qzKYguJ4A5Ce35P/qiZx1QdB1sPouZOO3eHt6UjY1s/d9JLbsP
WnPuUW0o/TE/IgW2Sas6seYZKtemvKn977INrogI96RqRlmiPjsyudcnqXwjxfCDUVDAMeCQnnGa
4Zszotp3jkRFmxbkkdSHlf62MSxyI7FQUWXhRiYoCsz8vkObUS31ED3CPii0MtledeqcRTx9gxhH
8C5ldmxkKmIDfIo+ovthLtN2HpZ4jsuRPk40p6Bb4wxTWo4PHPn/X8BrYjEDgG5f4+h9otVzsVxB
0W53T9NhqiuhOrruo/pKBEOkaLCWYD47cHcZ1He3nqz1xlYz7F0SoKaiL5po3yJzbUfdwCjqPzRY
wx6DZQ48wuLahZ9iZNV2DOYI/SCPjQP61WbV7qG/1rW0cVBA/vmALdjcGWFOjv7ZhhDvDvwbZ6mt
1eL1RfjU7rwG6nkShegc1pDvj0hj1RWS6JNdZuA86NCAIH6iQnN+jjUX/CEW3THqc4Ar2J9xUtZQ
D+3kneyl+5aA3biThVkjf3J2Wa98zO8S/pmCbbYXVqVLo1EjNdf+VyfuPFPMVE8fgxF8Z5IztiqT
Svppj9lYPVEAgdMgyNXuLuyrcmKuwBOvYWdcI1lJ7XycqQqxkvfoO6Vjg2oqhbcjAt62eyMuFOpw
VI8NCHONmHDK+URz6HKalcxedhMjMW7hPmidVdrc1fwHKzDaKOQFCvmFV6VcqUCxQI4ZARWkfDQC
uwQK0xP7GZGG13sY/63ENc712ABushgxIWdnC0CHj97DscZRMyMAuEnHAG3T3zHjvPLf8PfpV05i
bMExFGpDcZkysGx4fbx54VV6GxplwXzqdvcXJkIxJeELryHN8b/d9LW86eezHIrMLWqpd3Gwk6EV
2qBD0W55NmcXJqgWahPllKK5hro3BwhQ0nt6yf3lAoJOA4okQzzWIwTeywi4BHOqicUnTmEXLYbG
b48+H8UxGyAs2RMWxK+ccaaQ/6tPvayjAEkVbmYki+nAtjbz5Eeq+Iev6G8G5QEAjEZgjBtp6tpN
aygc5dH2eI6y8KFEuMaWSyJ3HDL4FSYqpA5MRJbjfz6VxkzfbIyfrvqN2SlM2+k7pMF7f8M1QCWu
vFYVe+r/U0ecxAdZRq7zCIXSkFr5oy82qAaLT+AWkjfD2RH5tU7IFOYHjwegXwJrONjFyeS80ygP
JyJskEhCQl25iaf6QGdjb9m4L0HsnzlPJKReoHHrUQHflYlpSee0NyDv6Vst2S9n6g0S1544XPFa
Cd9w+jkJErjGjW7kxQV6bd+/CB5ZmcezTivqVVTyCx9b3bQXX55FONsAEoCF8h5+PcrkpIOK9/bA
t+7YOw8mp77AT1IewoPfyQi949Lvp3qSWaKz/eyRyVdWH8DxTY3fIGjmzBUtJGsR8tQL+DMY/9N2
KJITyQdY0QoeVGnXDms03QVf/xOsgDyyJmGscoFG1/vU9oK1e8d5DxWxcsCIiDQGJrxEhBiCSX8+
i8Zp/mVy62MZLMbK7TbGnD3CmkvnzuCeFd+6b8la0sN6zgM5E395CPtK6X6/uqxngwYanSgFcXc3
B2ykVLOl4dnlF8GLEBcGFjX035qJumvZgtUoRlGiXg+5cwkhLaZ6u4BMcxUqnd9/GgwGbVUCX+1d
Ix2MvmA9MzVc3Ssij28iNTBSUqv8Ic7n4UAAnW3Ayt/ddG5gneQun5d8INMwJqNxUtpX1KtDAESO
F7fVsDlBYHjoEZQLJV4Det7kHyYs307aenSCQywBRjNHcnOlGIeK5w68GprIBJ74OvpBLwJO5EPV
iD40NZACsZ1bwHIzDnCzbBALdDXS4EKpusdHYKU4s3tTyv7yKsYPARk5O+L5RMOvJYmKCE4VN4mG
88FRL+bWes+2xIEwe39FHbvFVeS+JDjiF6v868dCHIgSR0STmh7DPul0QHqwDFO99hmdQ7RUOTZX
3lWJXPFv2BiOfhpAuW3KbYmP+999huvOw9IKnk8TJdqLtO30Fzrir4nK0S1psGegXcxZHu3dh+p9
WFJYENwV9bu+GBFUG/zXCtzOMmjICjGSBlad+rW4YKKmTFo9vj5eZRSWxzLranysHniY21ssJjES
xFEDq1gVQOmmAp1h4gjlTz0qQZ1YzYNWXTM6Poxsi9M+BXFlEvajZ3utCwC2+Iv8SOuDZ2H+yF+r
TA0ofywTowM3i/XFHBb/Xw7YSbgHhKK+8pOCxmZeOAXHSk1jJOJzZi5fTbhmgPcqZkwnRsoTm1bh
8DafMrAdLTyHkKYwLSIZ09WXST/osl6Ld4vRYwVrZVLa848tuQuxRX7w4KZG03Hh4gkTFX/I6nPp
hP0WUV+ITxwl1LzLTF9ZMMhYYo0WOZCKUzs3lYrCqMx8UFWBAvq8oWVl5LeU9u9WkZEXIrIjDyE9
g0c5z158dxWERQiU2cb1vngVEMiWUrdzgLhnimtbMwqlQQ7sFkxS9lnesMNHRYcIWGiZ7Qy0KXWz
N+OOYupbeMDAcYZfDLGk0ic1p2Mz3WYxDzRUpf3dJJUG1nDHYH3/SC3Q/vuK4dyuYNu3KN+SclSy
FSKOVvvSvOoLpA9uvQdgG2y6jtrVf/fBJ43mRhXfeoCxbRWaFyruP1x/ZcafXH8ne+Iiuo0yJs8d
GdGKq5svABOFcNq8AAVMXmqNGppQhKY9RV4ds8GkF+gEkenjcuO/R7LVDMCfS60QVR1FrdmPix0C
oDvg4Pq4IebzDiL1Y4hr0IeGt3/Z5pMg1ukE/+oLa8U07uuZowCTYpGUsBaZT4XYCGGEX8W0Oj6B
8BF21/ie9kLDD0krxeoyJWgK1EObNTVjPlFw9G6A5z3CDcPtprlVto+bR5Bv6BIpcLAg8qSnf0K3
IxitKuBph+7MA7ZaRjAK9wo1j+7rKwRrRJ9ukawNrzM3KxdP0jnXbnJJ9E+PgYPfOvd8i9QofmBu
XV1vSXSuxM9lDzd76dv/D21XtUMSeqYfXaLe/j1F/BQ6gnerT6Yi3GBx+1DigQSveKX2fprJJyWO
stZSAdDQlheGLMuHfJASWMEPIpMx32/d8i6aF/rfYD3XBUflmSeEe5xzSJCmA3G65A5Y8bRUJLcU
raOFM4Zky2kY7iG4xuZrbxjKmwtXyN6gMei/P6xNvU/rpmjmF+ndFBDvSHGuOgUj+krA89rFvAV/
kUeDep9OQ+HEezTUY9iDXCWaycx3+H/0W7M64LTJEDxt9j2elRZVFI1AvRJCKzgaEV3nKuMbLTBe
TJn6AQ7mq+kosSe/dLxi9wDm0P5hgXMevdgvz9pdlHUbhM9golIBDzClWm3V/yQ3OzurE1y7Pd+d
0+SSJEn+zZIHWZsBRfh1U3f3hkALX8Sx/YqB0jzoK5sjVoE+LHAeES3/jBIpjtHokJi2POTxB7vw
MTWI/4CuTJ4VrPOCFxWk9glYjYGSIbOyDYfjobS2Px0yaC5EYg4xzGqim2eiaPSZe8pPr2BL9223
kGOBOjGcJ8Vj0b/Tt17Qt3foox7lopMtdS3cldfA4eMt9L9nJzoE7khnVT0WLMi4HurcRDuN5zvf
7Z62JhtR/iRkYBsFWZB1iDm5df6c0FrfLJbI0kz2wxyl3YW6HEWpdAnyMbLtlq9tGuAcuHiBa2gQ
WGVfxAKKX4g9TjQjXr3ypEZz+3Ps7PMH/gsLGuvseKl4+xQ6bxGmqlH1hcGGDapirsHRuW3b+O/d
mPadL3zzQBoxDx7erQIzbT+h21vMDZXBY71nNMn84Jhxk+QVAboM/n9HxjYPaSdhFMFcx7/8nEzx
kQr/Gr6JgbgH6HSh+Irc4K8Ys7GQasiZGLfKMnHTm8vHDCIkesdcY3Fx8XjIpWc4uxnUunbQnPRh
lRCWEtxRTTjvNr4urlKN1BBNZpQ4bm5WviA5QULl33IaYeOVLKxKrn2DeZk6Bgv9vlvo0kydt1hG
w9a2UgLR1+vAmxbRtt/r9uzBu0xWgLKxUTRwHIn2EjSm052PtbuPgX9/11TSVAVRJDjh7kA0MdFv
WHrR7NwBy0a1htDeFJBTy6/WkCToJR+zgF1qiFYahqi8sE2Ske20w2YP1tZDo/DrqA/Y0e/NuhMt
XXFFV34XASUX4wzyyoV6/F2QG9Xx/VKlKnwKq174K9Ajm962yxwBXvsup2eL3CDNnDJrBgdpZvAd
EPhwIXG4egNKTn9/FOzciDeFY/79y0c44HM78BDuX8DDGzW5h1HXKi0sUhYL6jeYyuaCDFL62uNv
YQjt93Kdne66HIXQ0VFyvFK4hmvGXwUyCoCdG+NJQnBcIOsG1cZ43IaDoMy6aaEQVPqb8qXEvdXE
ME90tOEopo1CyX5RxsguAgne6RjsUSXOQM1Qgl1zHMk14Fhf8cESRxR/52sVKCgyunHE3P9nk2fL
9zn5vk3CRhGub1l7EhZDEZV7/rsxn6ttpaAEbW1fBarOKe4+xcIwrlxtb1N9fhzCV/CJIikLR2/u
Xs8OwuhKWTMVH5xa0Gg+ecuuuaQSgCQ/iMYMc7TEc3K6ehJ8CmGf9O8NxA1iA2A+v+P1EO9zsSAs
Z8hD/uD5GDsWUsHBEBNCNFsOItPLDEejvVptthkbw2uq1UsnfmDHVrpW7H/X2K1Rg2So/SBPiqEC
onk3jIR1X+YyR7w1Z3pMezJ1S+qHv7B8ml0DlTl0omOeMrdKTNxaGV0fokDlOoFijcIf9kj6ins1
D0Df2E48+48TEawnRm19QdDl01LojI9NmD4ipmGpK1hpuQGIES3mADftY7jpD45XKHe/Nk0rs8PU
v1qs0AIGG4wO1nCH2UfNPTyejrPdN0FLbEI2HiSTzLJsTNRXoOuaEH1v6rAgMA1gt5ZiRM4eMcje
Lmzx3sae9d0hHwPMA75P5SV8V0Ekaq6ulqcRIyz2tfEnX1Cp+ONCSc2fDkCv/aoH45+sgmTHCs4g
cHmYGoOXcV6d9/jy5jZ8JsCgyVFyaJ76mxXyLxgXnm3f5WVYjP1K+DLPfxumv/tuO6PT5IcWgSsH
5BQqnkhd7dKNHwM0kn6hgFtIrnOXA6+2DmOqwENyQgr22OwGRxkfLYQF6CNLVOhDVKbbQdEAWcgZ
kMEODB43L1sCBmf1/Mc2o+G908s/NQ0iDRa19I8wzjUMYTSyPgYl3YSqfdDQlS0bS2lyCtkrh98F
+txT7h1bFQwV2FN4QmisYiVPeBLNYoCwO85RWED8iio0lsB1GWbTbdYQSSRxlBz26uVOnNsiD7Di
KC9PfA68n5pS0rkqtc7bVThdCS/G+fVF1P2W4LBHRlRQNuDH7d3Ki2wsEVXPmCgsgYYpvpMRjlxN
jxfIkqhigj0S9N/hzGa8LiiKircmhPlmby/bPAPg3dpliACfr5fN1BI/m2XYN9ad1w7kjRecn/mj
dfG59bvkqkl0zGuJxTNSum58mfdO9tUqRAU0ZOxcn9QzNAu9B6qCKdhn//KaGFtXemv8B7HNNS2U
QLz0ZptW3mdt+bfJwU/dbqT7Pqsnt98czA0Qqt3gAzNVrG1h/7PG6cGH7DbSD9Lyu+RAUd0HAFBD
9aiRgK4xOtCRM6oy6H5cD7gHRjtxdb1qDk/DGOqdIEb8UoEi5nH7zDDP80l6GMFml4//z6gJ96Ww
qG+pTDlkc01H2GR79/PGuOjOXS35D0no7hWEf2CDhwPpT3DAk++GjS4MYY9/rX47AtT4zXwXxOFw
r9GQV7NIggA8W8br7qYo4IlH2gAPNJx0N5YLPCJJ0buPJkijnld6NNBK3Dedz7rWL9DIEob8j/gT
I81sm8LyFMTzrh/UcKSaO4thW4x757cO3jZEujzzBRaPmVAmrr91FZ5VnBYIas8ACMb3r4BI+/o2
G+NWWOIR4eGONAlPm6ywSZ1NJwU0MZLnl/R0nodaHFjoNW65SgjZ/fwwPip6JLZe3pA30DpmRb5P
YElzuyPr6oS1LNbMNSGuaaNqUd0WDwZ1CfFNblvLuUBrynjS8py9m8OPvjnIeOZ5WrrfotfckOvb
IvjvT8mrM2pLk7YmAXTjph7ApsUBRKMzHPZ3flhutA7WyOuGgptUX6MF7E97muD5qVgiA28Xg/40
XUd3tf40UQljezGDCV6PXl9/hvc+Cw1hHH2GZnKASrL1BI7sEUuMPTIALAmjCp99hAFkpOuXRhuy
lSGDC0hms0anWoN/3pivYlinxlhNkFiwt2LUyF8FL0FQzn3e5ooBHaESMTA7ezQZDs5Cb1t/NZCk
EfxRV6L0lW/VxS4dBpwD7ShEDgO/4wOeUWAD+nVf990jSJH2L0bIbgffUFSKxYjYkIqennlC6IFi
NL0pZXghjxoaU8QJdnaKk1TSBJHqmkOffs4hU/cQ1f6JOzZahT95ISkiyha3LwOQEo8LMc5G/Z+O
qA5k0C7a5hNXd7erNBt+exjY6jOwVPbu9RxBl1Z/hod6vSUezUiyWW3JEwPQ5I7wUTkJM+cwtTqJ
QUAQodpbAtrlMZPlG261Lw5l/3lfiQfTCh/THtKYUrvRSzsQOi4qdck0iXptDo1Q1sR2PF8K8Uly
hDse65aTmPkGu8XjGkoAKZUQSEHKnLRVtV8YXfG7AA0H1Xebe1OCWzM1f8jptOHuXgxtoZZ3b9JK
yslIjIGGxz3TbrWg3D3fiP+cNVy51Y5w5psLmNYKi8xHUb9sgrYR6ZxHG3IDugw5AHaUmZM/tHi7
2B5WNBcnmNzb8t1y+M3SnFLfe3ZxnhcKjz2wJ+y6UkzTDAyGg7+j2J8BDscZAxHe5YWx7w2Mholx
UBDeOv1fq1b9j6ZrGkhHXJs8II0rwa6GlbPLfsYV8ItMH8oWiiXNI/crlsW9qwYLtvqY0Db9VUUt
FfdmILgBdSLnKCa7YOSFpCW15dPfcMYX0h2VrLPsCc+9q0DpY8M6u5DwHFGzLCJsVKA3MH9ydFgE
kVCGgBtWKuuQdNtUCmBSV8f3/HaNRTNsvh8d70QjxTQEykWycq0wOoT520t5c/XvYC8Ccu2QgBrw
rk527W2rOenFJXCM17bzecUKSzAYUAM6nwRYhsFtUGaOaCnf84Uo4ATP/EIYDSA8biPTFyIw1Qcs
40DDichEAj/he9ZTdG6Z2/A7eWONp2H9zf2yjzoCyHZ5uqGDMgKT3vgkwcf+MnoftFB8PD9Dil+6
7yEyVAJQIuf7NQ8Rkq8NsKwECcKDuMdjz8T8f8kPU7m3pG54+70F6la2uMn6QeQpFK+t6rDidpjp
lqWnI4X+yFNskUfWmHgZw3qKk2nEaIQLKeUJWIx2XzuPeMiOoS/molFc2/K+uuF2ixgL8WH3JvV9
9v+2V2LiEv/ryOgKhoUIetOn8riNDqXWiEWQIVX3bRvo0HYTPQg8fPOdyVMP/nAjrV2uL4yQvw2+
MuEIPeHBCB/W/boBsUjEBweGqQcHPrCtBUdxZ0hNqg0z3ehc46fKld4+9/lz8FM/YqfTlQPjwOv+
mVbi6AFejKusEsZ+/Ls1OLlKD48b81o3Obz3fxNTVeytGRoxS/1ib2ssb+WKFQ+VND6xxrefB0oL
n7XangXb7Ttte0IHkxPNOg9xl1LpQEAQPuuMnDM1asVazBKsKqObGpgW3X5D1URemME/5KC01w1k
iR1Lgc0CcJG6tsmJ9IxzM3T5ZomE427RpgypH2es0JBZ9XT6LdJVevP5mEZ0sGVSRY/CYz5wEWmX
h/YVxSQ/Xsf0PAcCR9oeXkY4EaL9TMYVY2PanOyPBwZWHCZvExvmE14PcBUmxzXu1yZNsDAB8H2w
xuiWwyG53PhO/2gBmxap0aaj3Wu+OKo74NnEeH21FybQdovkpRijag5I1XR04TITi+tmoQlFCXVt
NKsn9SdLKc6fg0C15ICbJo8LVKphP4J3n1Zr2z0A1SLOc8X/iXOCbkXQw+xCMUkSrnNjg8/vQPyN
dL48SPtssJED2zImX3xYTsSg3YNY0gkkOIq6Py3B1iTDYebIAGdqeHpr7jDKfTveJWWBpdicFBmS
VttozrvqOpHk8YkWeQ6l6dAyVl5ia3QKx7Zdh5pqXLk0kNm/Z9hPvU6MWv3XoI/sPzkZm45dh4wY
bYYybx3T8pgV8RZYQAhkX79qVCZPVY+7PeHgWO/6kBWcsBPDPglUwXHMiTRHIdHr5eLyLnB0Du9G
ch1yuCI1bSXVmjE3bD/QgFM1c3IyeD/ymGkYtD/2ZumE0b/J8VtbQIndUXJPqJO8lTVRcCws9Y74
bnSM8md+X+nZB+bsbWzEzUETTm6rwDmfMVgfvxVpfRoHF5z5aTdYQQ95RRY7pyrZgHAaAonWnMog
5n0EKn9X19+PTV4kC+GwCdUG+d61NqsLmg+p/GcSZG106o4oUET3JKE3nxtBP4wZIY92b0VbH9q+
L4cqoMGOITF79+4A0XNkjgeufXovEMsraFyBJXqUmiYjK98/F3QMPDnvXTVKaFrO1WuuRHKN+3r0
nAIAIDCmKnIZt98WVWVbNTPXTA+k4iBgKJoBJcVMdn6BLdT9vrNimYkx3J7QWYOKtw0mCx4pGFEY
IoV18LwtnSSLFSyWAOZk6gMK2BPXxtQHpoq5gUos8xYFR+L9vuhy0AezSW/qlk7K/tf0NP++aNDx
zA/U143BRXhkww1TDO1e9x6YTZIElh9nKNvuwrL7vCqRDBZCn5fHGyqwD2Xq7ZuKvWQOT2asubPX
pcyHTyetL27mIf4b2a0Wk1JNd1oeKb5ckKETc1iY82Xn1tRY9RjRt258PPYIBnVxbq6HHgv+apTV
6vvWzcdqtUUo72GGh4HluTZ2LR4Vx7kYrzyagfsZRDHhCjukQ/V9/v0BYLHn7NG3OA1qvyDsBLz/
VhRwn6olXgnpuejz5TcL5c/NwzIQDXPVdnVFVw9VlKPF1HVQ6oHKQ0u8c+uj+tUJINioqnV2M4vB
MkJNsPBbXPDqygPCCe2U3x2PmFgrL6PCEPcP+2urmRR1/jNOdJ6RtP4TxR95ylAv3ep4OuFzcD3q
1dXT9O1uEUaUbCpnsEtU2AEZZe8EuNfPTvWeKXDlf/XVX5bqdwqyRfq7k2feEtQnAsPqQtNJQ+Z3
EKx6XAl9JeQ4XN8W5UxrHCsJQiVJpBNu/nzgx5P1cfWNdJDYkywtcU+gVe/JhYHuVDZD8SVafSSX
kAG3DkpIitLu3FJYjN0V1v+eqgeIt4N9OrnLOhVb+a1jIx8sFwAQacpw/Pr/O06622ob9eNantLo
ELFHzLshBTdyzh01G9r8KqPdOWtALhPVwvsEOR8mkkdw62nFja6syfUo6NGW5yhlnjRcGwyELYZs
u3FktYkjK32gZX2KhmMHnqhp0KuOLf/J34vGBha0yJ0WwN/1C9YA9TlBhFxuefqezcjjtz5JZzmz
vHkUT+JCmC4BJqSTHW7XpsNSjrgAqkNpGqpsvleXzezSAw0PbMdmchLJ5zHwfW9JsQsQVYXQcqwj
w0yLPV2y/ZDxl96vRtJcX253TA5HzeZQ6DYZXF3+c20WlTetGEMV/k/KqqTOVvGZ+A2fDItfif8S
WYHPn3HW8aFE/RzqPjJfO/aDXrc9ntlSS+SgdgS7feH5j06F5UtGHtwzDyoV9XyfjLV1fYyvrIWt
zB6WSoaU/MFtnxoxDsu3liuW1AVzNnRXkt90dObSDQQR9YKNNZu5s5OIyF3bUZTfrlCEMm0ylQho
qSnPZCFFxTiHGhuBWe2Uh+7l5JYveM0LfoF4oT0Wg+ELYBORQHvdRialLDv/n6ON8UIk6R80CoLg
X+uQR3f56aTT41jrjNpyonSLZqvStS4TVbXyn1ybd+YdMfy6yPRBinKeoZzOG/S9ywYJIY1RRmzz
L5dgF91zfg70MGAnJ2rl7vinOLSn/MmtGM5pYWmkbQnKL8a+Y4/7A7CaFyOlBc679x22V5le59Ve
BiK+ua4C5Gmo89MSA/Z5QPhV6NWIyg2CX4yisXEheIVFz5Q2jJOYPNL3Fq/AuBDO6fDxY2qwjHeA
KJzRRRCm1rbwzGSNx4vU8q5lGmZfIHtK99z7ed8ATuoNvhFb5YEbJn7H5f30G+AmGCMs9MqpcIMR
N/WjcjMyLhpbq4pFIGV4YU0+4JyZjxJnCOpz2Iu8BCOTfbcj9I6qtv1eowZjZbeoUv+XFOh5ebPs
6H7Ia0A0c/4u9y854RBLWpoRv5ScXxabyoGCH0rSxz2/w4QpMc/rF/Ew6T3GJP7xbWwXOoNkQ2x0
yHiVHEuzG8DP165gqKThvYcb1bvwub2SRWeCIoHdLtdKEdyoPMa9/21m6sF4M1dtTba81e1mEpkr
heNoGLRDEzCaGQv7iDMPt/jMXeKHvH3xkgiBJVh83B+sKD/kNcpHubQXdEJ+VuTjydZ48DEXcvGK
j2i198PqDSFLMA4C9XlQJABqqGUe3/SJM2F54yEC6tk0CLuvOD9/0IaXwBDZMGhtdQUkOSNEmEFj
u2EZ6yCWE5m1LKwd0SJigsmnyHuG1PpjfOCQHhAT96Arm/euPsS7adJAS95SY7pav+TfqeMLjo/e
9GfY3IYjp0K2icUl6k2d1bMeQkuSVMsC1rU86xAWZjwtKTnUSmucAx0GI+VjHrIcfEHfcK1dbmE1
fVOgVzJS4s+YuQjBsVru6QZVCazf1N9mR7WPi+pbiV5DRuqXG+eZkz7ouYY+MTEqjf2ixa56DTWH
u+mI3vNJAICm2AULqOGgJHvrT+vxACZjezkxZYwBRgOXc957+/brMb8O27PQ5B1eBfnuagOih78S
+bS8n+gYE/vTYSKFlF8CkrxqyrVfy3n23S9sPgWSFKidGTYxwBKq0OiEsKGwzIEnR9RbznrqECjP
XsuWinSuBFywY//H2u6rlI9/EOLgsia5g09GHHjFABwaq1zmQWtvAadFA6UukDEzS/n33sbmJd1n
8QHdcOsbxfIZ/5rF4b3cA8CBGpep2uREDCtGD6qI4qIxVfKLvRSf1e4SlSD3ecXBybCdl7jwth8Z
LYbSSDBjoOwehakI+yk3D3QkKN0Tz/VfttQF5gHt+M5EzNUPRmsbKWAgSdw0G9gBgBmDJ82cotKJ
vQbvR+/8P8Sj2xtKAA5e6054lfURgUlBacA0zTp5tvKBbanA5XZGqTFIsbOxH3Kqs21gH8X0ruwL
kBbB8/jm+jqvwg/GUcSApwuOGcW2dMd/Mi8UYKl1kh0yCfxMDseu9ZC1KornyX4hs7wyo9rkeyjU
kSpKHsqQsulaSNVBikIJqMQ90vNcafAUpBD+P/o8rKiXgbQpIEjKM9Kc9Dlc6bHWZaRkmyUlieXG
PNGOhteVeHYqb2urPYh15EPFqKGE4QddxtuaqThBwrAOSOrSrLqMTrzYSrc9jw7q7x74lqRlEsRY
oRlB0y+xd8JxzD9wHt7hiTdBQquqbRFRBD+jLH17k0rlfWfpI47DDfq/xCI0qLfYOQzsmblv/cBt
GbOKdFml9I+rdMd6/MJ9Y6KuWGXASvrtHca4MZ5RpT5cSHioCbMFK0CA9MmQv/Xu/gYUijZ5Qdpy
dY5cSZPhXIs8wQeCSCmcsrK+SsiEjfRtdNwDMI9pQcFkzfKMjxP8Ma99tXqoh9Oj7upH2jdnhJxH
igFAhMQm7IVXUHRZLq0k6vwSNvmSGlb1KQLvAU2aNcUOIitRLbK2QA3tsNrFj9DLDXsC991BQ1N7
3iSOuM2YCgtAyob1YoMk9RmAgpKw/IY4MSnj1cfg7Zw0dPbrtjLGv8QoJvrUpJ8uF9HtZSvidkxu
yoIC2RtyrPPSZYpeOpR9BkodgFaHJnf7lKUFFoEB1ouIaA4OM5/KxpQIydJlIB4/UQKjN2pPBpqV
PvgM6IkyV3wEDjeFyHC0kqOwT+SEy1A6aH27AehyczewZuzjU04D9QbsF5t3RFQI+ia3d5gi6JkM
HVehTFsegq18dPSqqSaOfsEepCmCJ4CRVIqxIAzJ9YF4jK+8+joKICPOelp/dqJhFjswsDuKWgz5
ZdiXD3alHWhd8PL59dlCfo4Lf/4+YK7vg08Ryxfje5gkMcIvHp7YqM9+0uJ56+yrQuxIP6j2eskf
vdDt3ycXzh/QNCJZHL8/2KBPQ0XvtwmOHxqcPqwmT5y5qbC0IAqDBuXdU/b6/jPbCtubW1H800aq
qwBybPQO3aAWi8SiHedDj/psB55FxCOVC9W+HFwA60yrmuV0Ctg9mvsPs9oYRmlocVF/XCTpSsbZ
yxJ7E+Zh8I01jlBhHrMCStsAA5cL76cr8/H4N6Rfb5fV/lW+fmjZg9mJRoIynlwlfksRa53awn25
WLJpgVZOaKEijE5zwbaRVPYE/9dsnFYM62tnt3oPC3IxdNu6/crN+UZwNXRhPeR+EJcSBSnH6htE
Ry4Qf5rL7WOwPkDa7qbad1O5UCZkx6ckUlylAcoYn27bCu05nMROYceoWcsO6sb1ye5biAPhbDZp
+0Se3h4kCWhwj6rzldg/vI9rlh5E8EITFdKE5gpv7WEFoPare16BK4rz7uCs97Ykn2yiyOwNdWiu
iAcZGH/YMUYE1WhBxVgKiCwSYB/Ho/gj7ZF3m0WQqkeWk1NO9zO/MnOf44ShuQqP9VpNK7XJWxHx
iZEeWzsa1qH6amBAEnSToTc3TMRg/8y+tYzvPIiuW/xMNbuYcZ3Jlg8rtfAOJWhc58zx9xvU+uwX
3WeN5zxAxxPHXXUAms4cP+KHs0bS8/K9+2zmIOls1lfKdkT8eu9DRim7Uxl44cxEklBk7kzVPu9Z
zVggzpRRnnXi7hdcFgQe4+2uD5stfhFiY08hez/h/oiGf5ep6aJzLeMDFeOpKR+Ii/DytGUlakwf
nC58/RYyLR53P0ZDU5yf34KRCYNO8pNT6fPfIQXItjqELWF8XdXJv2EyUiAw/KSfjoL6PYDSNvMS
71fQ/wzFHKqFSczPGzYOAXVHfWfttEiyab9M5+fK8JJ0Krhc2xw4JtBCCkJFLLKZEpMvVmopxnXJ
FpVG4eQTt/Wop+5pRhmsHAMbGmcpUUAdSn1ORQGKF+SVbxsUZDJtB2o2gw8QYml72Mun1Ie+aRNb
QXXkoa8jicgNq83Y4rGeVdNpfFFB6PXdnwQ4zIiJZolW1ZB/E9lSN5pBj4SaX5Iq7Q4w6ka2Oltx
GbC7SQawpi2Eik52fjuWRDWtCpzmWDLQR3Q+hgUoO0o0BkcsiOP8xp09F9FGPHTObeboQZQl+gnC
71N8X64CKmIcP/sNvvzXBoKH7nijdFOmXKECH61vEiuTxWLoWqMInwUJjjTVY7aNjQv6mcM4eoBu
J+Ifi4xGjxw9ngvpPtMp0wiOil4EwgcIunwlyLQh2pJwjjYn6mNlJS4OhfB8nKjU9AMANIyyNOyL
8xLrpd9fLM33Psm2gS0a/AskSG5/fimVOUlXlD/DM+TMZyy2rZHJSFMCd7D+mwT3ow6MWNk2zgnR
27d6xe2rMl4TP6Y0xRrR1qr6kucegQRi7s62UIMhRbY4bkDL3djYf8ok8cbJT2BwdEwcJA413G7R
/97g3yTxv8qVADkpLYoj/fGYcbSVyAEPwFFvXw1uL8+PQ2Zy4mn1zfMPUcrdA8kdSCIscebyEFZE
cBJMw+9hbShhedKI+iMzB15clJthGUzvAfOwm8u8a33OXeJWfTz2TpAxDmZJJJdeQ/cCS3rEi1Dg
tn+dm93pxmNpJV0gRmS56A3dEwt6Dr96cAiaUrFkaZYd+KpWlvdhkihSs0cXg/piM6qqKAzdqMnn
NAm6UXsyO7RBgT3tM7g+qMWTTiAufb3909cRtTFFnxuhBv8FPu/rTJGkd3YdUcfbCZPOPySb7iIc
2Klhpjnd1O5p1IC+dxv72Nf0+o2m8udNv9xDsm3F1C3/k0nZ9s3SnThzBr+eI0NWbHOxb4qvYoKx
XnU7hCXMj6ri5jhzPuRCNPlKUGQwbtsplYVM51uk7VqiWy5eC3wQzyuYuY5v2samLE0+6TVsq+GM
JIXjGk+9DS5ycF9FnYm0aZoMoXky6zYf6FML5iRjPr1o8wuqybVSJAS4Lmu5izRhRmqGewPC8AGs
aAEU23b3pkqcf2xMAM+6HOgk17HAeOFyU+tYKpzrRdrdXbFVIwWrIoWBV9U7wJKeV2qq4Sq9B1vK
x+FQyZEUJ8qVVi6IlXZr0emp/Y3630EHMuYISm992AGVf2zyvPawyR81DQ11BYatK/gf3Sb+Idzf
SGXU0KyDakzmDct3Wa7ivB0m/DaWxT6UcsXFhxLADNO9Q4G8E8Wqaho5Lq+xusMc2F7gFcJ0pvos
qtRK7LoULE1GHogVL/s3FcDPHQwqJXc6syHgBsPrvK0uoWgZzp+YnoC+Qb2arwWGHi2Jo+KTdqA4
7on2XcNunN7MxazZMKLMrtwwNfeVLoYP8oP5JGJxWSV0N/G2mhx1X5ZJ1fDcugY/GVnh1HN+nOE5
04xL6BDb0gFWKVaM2QDqAuLdaQIwSd15bmy7gxXDyRT0QWZbd1sjoU6jg2JNqI1YbFrc4HKrwgJ6
qmQbsG+QIAhcc2eOHnIASgF3r6jCFZmwDAGYzl8kHN6BG74iHJEEXtLAySYLyfZpPvYqeRjjZtnC
iRNqT8l+hp5CxPFT/PAD4FW+MliB+TfwN7cX2DmjmZ+k1pML78pjnhRK9FxmwskMS6fWsZqngXgF
K50B32IqxJuzbEEZh0B/cW6iScb9T81b9tsviGkwxf7LtJrTqi/T8DMRXqecWvDkGOrIUK7YkbDt
AavkvslGkqTrJco3oYfjA87S51H2qCALf3EThMOgYOAoSFyJOtypcnHIDXpepy+FYk3NDSZnOWr0
5UDzMHw2Zq1vRZhKAXf6WQN0yBuZx6DtQNMMGOxOiqn4/S9Edm+Hp1vFLuAdNhuqK6uD/O3nc0ID
patm1yef+ZtIoJTW9n+GaxBDXeMdQUMIAqNUZtrErJJCWSxAbwJvCfgnEH/lP5xR6PosAdjO5r9z
SzAe1GmcTlMLDZuEjxAKh+8qHkKvue0K/T48afzJTvs8+kluRdorsUry9tJKUe9PhiFKCDwOX46S
cAl1XE5x71WkZpKiME4CBB5PBlsvwVdCRkqsLIkqEMQwABakusRlSZoNNjPqUT9Ij4GEBo055cF/
3Ks9hZz74jU6SL2zAhYLhRhOpPF7XhRYmg9g7QvvriMgbXXSwm/ZX+vtaQeDQF5OKYgSFSNgtmOw
8OaAXHNgCN8LCzo5M4lglWDz2M66A/pCKaF2ez//z5b++gTHR/hbq0jfosgnS2XZV2DIhDScLuN2
Ku22iyO21xeQNdjLvtXje6WjRrfoSB17ETIRM+gDKVgxWibJ64p0wPx7N1ELArvhthc2opHN/Jbi
c6X/mYms3H1LhsJcfDNprYUNKWtLjQsKzi2T2TZEM2fbiAPqviER04oStXm0S6tHVhp65OR9ua6i
JyHS5dz9JD3mof+lkPKmKaH2p0pb/NN46KDwCCr4UBu4jJLG/W5xD05MkGGIPB7NhQQPhYtqnpA8
TgF/qdIO2Tqd18KCDfFcoy/6GtgkYuiO7BE07XNdHiigcKnBDyF9/otcgzYEAIJqV6TknbXbajwt
biAz8OuJt8GE4AuLcViR7M/vn1YNjqjn/azKQruxCf5gKmXEFldXhIBHATw/e5dLZvY8aog37QyL
9WugLW5hLraTRq0pgQROEPgEKMCEQodgcZ2PS6foX1TQ6ciIf6QohIyFrHXl9qsNpeodYON9hJWS
+xH9kXxwprzVFBUXOlmPt0IyP/EoQ5s2W5dCOjLns3l/4VxJBlDn/IuZpLqlCXC3BtDvHCwDc8nK
jUbRT2ApwSBGq1up76Jc8E7beV0l+1GrgSOwx/Qyws4ZfZCC8ALabfq6PqBWhbumloSNROf7Zw7T
vLHiqZ/fOSLWy52jMbvNAERJoaUzxz3bMXARU7K18vA28ZGzc5VXJsikpMx0nqLrSkN4bf3iOafC
GAbDoe38+O06ZOJ5kXmfS9Ef5mWqpL4JW7ZwjqMHNd5TO9PNSf39ndhx6FXaWsdhoJpcBucALvpw
g00dkhjUF7tWADLHW0PYJv1ue8kOumlwKY9YiAhj9gsDzReOBJD+xt8BWr8SKCvPRptAKAMxLz6w
RO008DAPBwR3sD+MrfAj7rcXSpmj0xNdXHL8U1wqb4nu01rEwhfbxKQCxrUs64YW6sfSPxbJUS3F
bIDqt15vPTbBzUG6AfpyBYjNoh5atF8goJP9xnQqL4wBS1RIuAGLagvLUa/U+FtKXXRm+w0dU22L
EmBeyUC4ZCeiaKYJVt3tgCbBB8icNAzkIRbljjoE6f5s1m3Q0s5xxC8o2rdtV7j/ie729Qv4n+rm
U9d/6Xo1v1Rj321x0pjwDxx+ypiHX1ACLvaarhEx0pP0mYXoe2BINUvA4tbGDVET2lhK50DAzhCy
PhsSaSg+uBiTugzQqAcLadrGE0K0H9ByRKxS7J3nLz9qMUiB89dR1UFZqgqAZGLenT4SxCgO7Vsr
pmyr7mMyPgvFe0/lEI5b2/oByTEzKYE2p9+V1vdbC6xKTyllJ15FcWT+S20xG/5ufUIJd4syqvp0
78p2nxDWnKud5kO8CcQAck4SlwdTa7WtGkPpGrD+kNyxn4iDhXGg7QGtr9+tCLzjzov2bE587dBs
p1oMbPQVTI4OvMG5u7aN42ZJQQDCCW6UlYDhpEh2WpOHQ07aQnqs+O0OWnEDOF4J31aiILVzKgVq
Bt1Kceqt9+nw//XJAtBqgMwcyzDzlPupm9sBO+oZA87LXDn90DumdJ0OaNsGR3xKr6EeTICZyxAw
un69xs8Yqwcd2cv/IyemoJK3Xt67HCQWZMz5WQSJTM9R1DQ+JL4p2qwZyqwQD5aMHuyZuC04zjFY
ZjNMhatCYxvo+pbhzjr5J+hxDMNL4GnuZ2Klr35IMaCnz4gnw7rCk+fpFUiW35NlTPibSdpQke8E
MmaItCdBZkDo2q+7RdcUg7ksRgksARI4kidUWtb3pg2xyVSERFUFI7t5njEb0IVdNciPWUmRi32e
svjGAQHvhZ9xhhgeYRwdQhEbljzeSFyyYIxyC/1LqXNK4+HHGcSR1rwegpYybC5sPNdHLIUGCD3i
/shIihR/b3L8i1g9H92Slyxa9l5cAdnbz3ldeadMKvkOL69z/eigTeyA5KfFSPA/Ab98ZMi7jM/m
pLSly5ihz9xzrbVnEIHG1KQpiWmeT4OfqzWTXTp68S1Tuu4X+liAijzfNP2MEkMxycXh58iB3xAR
50Gb7OJAQ+ZGOaoCEgRMN4KNiE0cF+l6NHetTfoQMF9+qsFYqC6N2TvLZARvSIje5up4HPgsBWe1
V7GcDsHO15kpKD8kEB/m9FPUdbIR/ezneiz+YkOAn1HHhkTOjK46hblw4/sCgryuKN5S1RrWyn4n
ED9Y59UjHJhNoK7bEyxKolHM5P6Qf+LpAJE04/OmxR9tcMZoIg0GpSHwPBGVIFSlJMl68Zr1ZFrl
bTypoaKMusc0e6ZPa2hJj1GdbQOHjWPmqF32rwZrCyLa5em0LLJFe15NvhW0S1yGB7zKf1jWzc7v
TcjBq+KRtopMNqzt7XaqqaKHyiyHqG+VuwaMZ870t4zJki9LTc9moj2VJ8+XZL59gKk6TJC+LiAJ
g8KJHZwvgWOPB3MSdlGKnXDyUYopBE0sZw1b+w9H1rSxtgXCYingeWSeH5hc+IZ+k6VxM4EvTRP6
7r64kxZRMwNvW1Hg5ZLikQPttt03/1fk7CwO6YBvnTeWeXD/DbNj8oo1FQTULC73TOTAvlcyc+DI
zmYHApcz592XT+eH07guS3JGgpyYAiRhuRYnh0NgTZRE+v99k8dmhJTFccx0xHCPmem+0G4rsJWI
pEo0IoIBqAvm4BYQR+pqKC7vtzm+QVMRkUs+v/jZF89UMX3fTR7JcJ0JZireMJLBTsbrEPJqE/Mk
vGwnJR+CGS/pyFtEDTYwPq8EIcJDitv90SJMS0w9y42IAzQ/obdF+2tQh1eJthF0oyI+fd/iQUpE
aa7I7CdnGmbU9kpekSN235A6erRMEn0KDtCg5PBUMd+wdEW+0/9xqNiWb1QCvYtob+VPkSEwfg5X
JR8RD95IGCjbrhfhpL70R7rMmHxfObKC8FwzwKN2IJ5POuC2MhvT5ZR0EbNJi19fpPxM4d6aXaHM
pcRUCObEXz/9ze1yC0zV/KGT0DO2qtaYUUmkmra5zp/zZCLKVhF+J+laSSyZ1yona+oPnpFf2rfH
T7DgDLikbVSVnV9Bxb9dj6QUmg8gQ+a166eoB4T6ccEoI+W72565VPw2uvc3Z5l0Lj1s8iqs9Il3
xmvPV/t4EO3Mhwz0mTb2Fn/dbha3psVdWxdzSvK8Vp0f5uNVhR9j1Cqwk5j/onWrviyHYHu5qsNg
+rhF505k29wU8rialSKVDVvJsD0i6GBJxLnIvXDpmB4Iw91+7XgQAlhX4yHLt8HK+pr6DYZTr9uy
qvEhM9t3wL4BDLkafF+Ypywq/cOVg+YoZJDI3wSHHy+gIrE3wbZb6rsrpaoifbHpORt/A7zGsYSK
QP12kCjneG51f5r3sxKXSgQqKMhs4oTtQEspd/+iBiJqI31KWd/uw71X+2zKFCnlSM/bqm5geyIz
9pmOdDGDx0xbVubYWMgdK/26ax3IE0Yc/ibCt+VYu7w3Q5O9/Vpu7kojIBypn1CLBjPC1PeAfI6N
PfuPfmgYoqVczYPBwqjMnyl5FQt/kH8qOW5Us5vbZ5ZPwsVAnA7mQzFLc3e7ojfA2PLU4VEhFSCH
QFCOJOCiM9oUn4e3i3bNRQLLuoabNsiY/5muP1VLCh5QH5ju4AGb2O0GWSILFd5z2Igcs8PRknd2
r4bFVJ0C6NZviLretYoxgaWLe2WUg+srWYaPB44k3i6g0tDQiBzPXLBIZkzxxQvp7aSMj0t0gnxh
qpUrQ+tEWaACezaZsZ82NOcKdYiCgQu5SiUqnOvOWXX25wYZYfrXRozyqSqvkDxBtBFJ7Hi8EoT1
iMflZZC5hRSKIryzGnwkEwYX6PdLQpDOGWnRpVLyzt86IMGk1HseIs7Gz6XmZwsNxib9pDJ2i0qW
bWYDriUCZ2VdHPVzAwoM5LTyJIFzc8BA5n+6I4w6acP0LqtG2sYZ+ZMJlZ7X5SvnpDGsHKD9R7qk
LwvGqY/BzSEn6pLixTYtoXiMEllOWsMUqR3GiVUqWMhIAu9Bi7bHE9Q/Kbh7C8E82tvfTy67591O
Q4qlD7nhl7kagvMYzhFGAhTqIMiBHHd0PBOdXZhRlkb3md5q6CCdOlfjqsefdG6DvDT42dJaZfjz
j8lIPNXQXnRP4Cf6KAys6s4vTWop4TdIBIbj50xPMpfO83Vz8hKnvCsYvqfvqMRNptkseufzFFoQ
KyON549nzBrSP3lbKPwrkdyevpBFdygYFp1P7q5iGcAWo54Zd1hEax3QXV1GFKgIWuDtHSSWszF9
TBdrv6ofXnWza9/qeoma0IjiRa2u+9pltK5PC52Dku7sXQwZmN527Ckkube7IbgiNzB/0KloFdxI
uqdbMkJNT419tn3HhVgYxU7+tMUlv8jMYv44l35h0z3LiOdPZGuLodFTQxR5D0O0qiE6axF2x9hf
E8UbzzZvRiND3BI97Qi93aPle6xJNm3cvxndcoeQAnQMAp4Si5ll+c4o0M69d8L9xzqiC6F9i4rp
raIjbJU8vxtg0lr0toQ8Fi2IaXuZDvzQypAA0bGoTfYNEMlnLMfyMj3eUBZR2vg26fGr6QiU86y/
PZJ+rNPPdTS2CIEjypFW6ZlPs613zf08MsQ+pCkpZpKD4wY1e5mw5ehfaKy8ZWV4o9d0RttJZamF
YFeIrEcX6NoEzXle4D4x6/IfCzdYgMZdPQHrsA+vkFxdzpJSejBtETeM0w5u+OheGSXGEDeze7fO
VORnO21JsxLdheXuZSGXye6Xm1oRcSdws6t+Amykif7Y3vpqSgefvdXI0qqjRFiZk0rUNpfwS0BW
TY/O17RYbfBQ4V7WuQveQEiyeyW1duIQOQO+OJCsZMAoApt8FhslpvNM9wR4jJcUHbf1xJtMSzLx
BNVVWe137/yKuO4PQKtgXME+VAK+J+cSndxQlqg7GzPXkcv3W/D9FssUE9nTZZTejXtpZvFVMx6V
hw0kRAjV/9EHwDK5LHcrBmP0xJ53KEA4z34GpADo2XUy2hGplmOjPrO1RpVElO8Q7C2T3k5qZvxY
XhZiXlbKZCQudA/Fo7BGrZebuiC3xAUP/qaZzyW9mxw4ZsOIOyb61362GnNw9YUCA0zbtjA9acQV
afQMkEdwcYqpO+FLwe1l9jLj5CQc49SHHZF/Zc5S38w1Qwt53d/YtZVLbOVyy4XNNOScEkdpTTU+
W/3e6T7HI/5S8sClJnh646+aNk+WcE45OTIiCgyaKJtgzBywTO45/np7MkmBtliDBu5uVgJPO/Ij
BIfwmu3HK6f/KRwU09Wm4D/L8h+YlDWdGVy15LNVpY6YUKnjSrwjo3cK7y7yc7kYk+40v8h/j0DC
3DSiZ5acmckkP5pZsl2ZjQPCOtRpnnJzD71rlzkaSl9BZCBl6sb1eZepASUuGymths0m5zwPli1f
Pa3148/ogNRpePtxb0OF3uS0utkl/h0ZY6a8dEkBwgJsX6EibakdTNeykmBOzWMMkHsb7fQ94dOo
ZEraIWejJkGmGKAboLKRjO/4aH+tShtYjGoAIiLv4sVrPhLF6JjosOjEvZv8PYWxTiBJqyWCwBZ7
46nuZEmZQRgDzsNnPX0qWAcNyFJejSTrBOhQYbne43hjCHhkER9Uaqwwz7C0YRoTZpOIo27Nrcsd
S7EdqkxsVlSN1PyQtbC0giF4S5GTTFsF4saDwslU1sEBDnW+T941kR0rWzOIhIrRalLra4xs4G/H
2cbWLanMcd+6mCSq1pKV5qvYjVnCD/o09h56XxqnOnz/NB3GWF+3Q4kLCr0rWAmcJ3k64dzdHS83
FriimQ28MJANEWAgz7OK3aekP52JOAHZ5WfHj9VgmtMGmrQB14hd4RRyx9vGOershORQ/Q19BfBN
6PfedRJSrPIoSs+kSqkYzykdLTiuIYQSVJOc9GRoaDPUo0PeD32v9Ern/JeLkdhpoTrHwn+Dnny+
UQjtlFOP2PEf9Va0bh7b0fKR4BixYDmT6gKXx2SGJjSaglZLSKQKjiSVLOpgQtBr7TBDpdgFG1AL
ED/eeYybS8n4iUZxZtFpSQWkfOZXXFf17IZnrIdb/9L54sz0+glGzlMrZnisgHYOjia0/6ugFL/U
g1fB3uoTSb5Jg8ICcys8eWEsWuEYoM/jDOmwuDCr72r6KR21ZP8Mn/1a0/MnPwTc0dzaOpYb/Ac7
QKnbcqqxNCI50mNVH7u5iXrJ+jMkJr2t4lLzcELu7uPYC9LeC60yvq8V0BK+FGz/aFeEPVht9p0F
+FoDLIObFYDOKbeGJjwfv4UVmUa1Hyfzo8BS0maQdYDTCaPQcykUSSetV2mymTvLaFudvl/+Ymtj
zt4NEghlDmDRLBWt8hYU2ig1FLXMS2BdsrgcdGz6zOQ5WnUxC+QNAktx1LyXB9hjhvKVQfy6niF7
wR0Xh/+vhTF1HL516fkZ5XPM4SAsOqLCiDh5JTJsaE+81+gC9JrBWQghxNa+SfnrqUk6g2u0Lg0Y
Khr4xoEQ+Du7Gduu0D/BqxTNbDpebjbJs/SoEiGgTkMxfEdZ0V2AqYXiOeNtgvDvOM8uxziicLVJ
BukQYXBPSE7ZDlJg13b06KT9fsG98Ix7YPsJcIzobvgVpo2Q41Wz4wNZVcuxp1JOQ19j17FyufAg
WxBadarAfU2Ym5byLD02Y5OII9a/zgGvRbBQBgeRmaqgZbkhtnYqwMezHAUWPs7gPSoWZeHpz33v
gETZTyZlJpE09D+Z09PSvINMSl3aKI2V57sDIeByJcsTO84l8HzZQxh/5TLLhpeH0Rc5++9hY++Q
ovjI3AuFpIPz4MCoewUjcUB6MDfVypJaL+2w8ZoD503m9o5rLoupl7o7nidkBC9hfEwsbadCMOzk
Aym5R5X2h+TcJttr1TwSJZjPyD0ciWapGmic1irpFiGuSWBGVt5s01MNKtxvSS46zmPhOevwc9Q1
yV+A5hIAf2ZNjpy/kEy7YzyhhkTN4+UcTJxp1jZwDsFPDifVviXVLunUg1tSoDjlByGMv18yzXb5
5dUEK62xP8SjtZ/Nku8IinDlzhBOq10apiSp5KkZVb9ysO2S1SjJ//9N8vqli1tnRoyvfMsKsA+a
4WkN7ISBPRw/WxzlGzqqrYzjqS484ioRIQ64yzQMeVuOx0R9VPvdFiEuTfuQiGVSYrFj50ywYujC
kv2FfOaWn4j9QNpdQTrJ0Z5lSUEe3LF1qXiiVCDHdZQp5vQqNH9Own22x7Gj1Tmeup5M5yuu8D13
AeDGaAR4ztFanOtObXXqjUSs9myO7qNMLycB+8LE8JKxsTV/CdBNgKLtuqJc96aXqlid/E2E2Xlk
B7uLG15xIzTGiVSth68gKg7gldyZBZHxNXBjH1K0V1UW01q5BICtlCz3GI58LfJZ4fWv5U4PLSDR
iC0tUu46m4l8bHL/UfojxdEh9AdAs+kTjUkz/sf21p+mP6VuVxrTdy1DqpY9E/xt92imDGUTQoPg
wJ9/l1xGVSH5pkG+lgI8EKBFpSSKnlVTjrRVA4+x7etLMpoz0i4YZ9ArjicK/IYD8lahlAJYw0sE
CGdLyr4DdMMiAp+7XSgHb5i4OmrJbzQOsvfnUMuMTfWJC5c46P6OcijS5ruQ62gGX8p/u6lIpGm3
mBEYZydd9AUGOT6nPv+p0UkKUJj5bx1MpnfCXA3YYQJD91BPEMbaMPCoOIderEv2fqX/dLUl/onO
rbL4EOULzHAOm0eBJHLgfwsWWiwolY6aLshV0D3b3a+I26V78j1QYW9QkcmBYZkbnNDI/Wzm6p8L
Y++wtvHnOqw1HoRIDEvIHXgtM/9qum/tZ4mWwUMdxqMK5/e2KMRHQHms+erk723BYu1u+e5QZDBr
R3GIpfMf4xS5bmtO5oCzXKuONYbiLtHK872xlJ1RthEjDd3tZMaT59MNR5WsXNQ+ztYjHteiL43b
uPzpqQ8Irw4jnGlDf2Yp9kFNKvtpKaR1tKQrKdL1G9C3Mb4FFIWMj4+sdUbbYd0HqYMPr9oq5qna
Pl9UGyzrwR8CoXVouLk8l9j7bUCRYFesTzGJ+4Gr+y8jD/eAC3jqpL74xDIQYmdH/eUzPXryb7wy
nCGQqyEhArdrLvpAo95A+/PeAJLtU1LBMLYvqoxKK8NlA00DjOJYk9JwZY8qX5wB/nhBrMxsEemS
v6xSKZ+ydJNzI+zBj+tZ6DKuLru+IpUxWXVt4gsFN+GcXRKGlr8MUa+5V+DyHbKh1LOF8YnbKuoI
ntIkhlpZSbXHDO+KOjlofngkpdmmYMfrZI5+MOKldNbnGEVwZD3oVwQsvXb+u23mN86d5Mv6WgdP
G0/5NYAVp9jkTzK3KPVWkeOIpv+MurzKiUidXORv6Yq4JDUKqVTHHqoEjgvwGfWVWxac9RNteYp9
PXcbZwh04wFerJcF85xW5MaDbICRkb0OEQCtnl8hbqRZRbeFmE4SdMLiusCqZ4gzFgA8Ult6ibpN
HGglK7bYi/tY6UFPayyNV3gVdBO/MSe4a43iRZJG1KsNKztHO0pNfhnBF7kpZjvzP0bn8NRq1kNv
NLGE78FZQdoJwiVXrTrNgxi8Wg86fIE+W8ecrAIizVGV3E7n98lCCyX1SKVDgx3nF+eI0C8doWxH
wNhjrv3ddqeFNfKQYJXpX95v72Nn7dJDbQ/VvOg7Lu2yizHGNJnFIap+oeCi5Mf1Wv/5Tznkn+OG
PP8arTMMLRq/OzL91/FDBBNTgEu1v+sQ6ElJYRjM97chCXh0QO55cA==
`protect end_protected
