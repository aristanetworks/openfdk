--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
HxBoLn5Jqz+zxa37VurvX/fOKrFdKHVhtCb3O6YitQWBzklllS067YLNNiyGBcz2Lcn/kMglcKzt
x6yWnaxNfJshpPJcnTE1p1OUAdRd1ys+zFMfLp8q2wwzdxOBN6BIDqABpJMg9+/3q3BFT7j3nxtO
voRsuDOb2Hngw1LsOOkOAR1xJSJg/lor6ykTcKzj1tMrMLJm2OER7Dg4N2JbnUPTBWZU88ePQxfd
2LJ4uG7cBYKbfGTHcvhnvWWgZ1CGg5Z3bj0oM4c0xefCo0xy8k6ZpWhdKf58vEjODpJkWFMEK9Tu
LnjWYfPSjyEB2hLMcd125dHh5NOS6ujjYx0mVQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="3+9426tjU9yv5fB5PJr0r17cM5loJKhoVOQKXIOv5TM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
tI2ERYMnENwLwuQyG+J9IKekzji9PJoKT2sXzDLv2rXtNJX3Ec5fD7LJIDd3uEIJ2dLdsHcwsdO1
8vHxEBTxpgnyP+Ud1EtbE7WE1QRI+ehAndheBQwmZBsKku5TUK/obT+xhzh/pRnWcvKs417uiNFh
6j13e5jqhNr5glhClol0d3f1Wb4tk5N4gJT83cGSHUUil7qXpuNjc4vaQGvajHLuD+eRTZNVvZlw
ALAtQmIzDfgbAuVmN9PB9EXgS657mnoYxJhjtWZZW+upkVqWDYgDwg0tfPPDl4H1RG+tVwBE0ArJ
Pg8FXhJQtuHHT/kdNiNWg/QQpJ/W94NWftMk6g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="glQBN7VLFPVzwLKIkXYJkqQZk3GRygfLCFGfvTHq9dY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 36560)
`protect data_block
MmcxjRH1SVcfW7ReIZPDRAhFS7pJhvCMKBSlB8ij6iT+Flvmd7nU6JatS5+WPVNuHPwFWoIO4vsZ
5RcsV+qc4UK3LBDmJu86SqQtxGlWZL5EvU0+DYivNe2WLV8QyouCh1l4H7oKTqKl1SvlgVJlwvGL
b3Te4io8QRCyQAmTucfsRHZUBZ3NCoqFg8H2PzBIL02qYZgLsc5NS+j/eYbJzSfJcnFZLrMH4zlQ
KwPodc3/4fW0CXtBt+kyJcp25uTWZWsFw5ej/4b9zeULOfrNFIJW3/ImTCp7KlTrZ8HUV1tZpqdD
FvYw5VPiTgLfzLmJIVW9bj8vuH5mvtVxfQQy3Qz4TqFVpLfpBH/HXxsKCiawZNK4vtYNvZhalCet
xzMjw6LE25+K6/7WI4dvO3wVmzqhJXX3LeYpecWeYgkybzaiZ5tLYH2ZLO30OyXJY8gBx4UhSzb+
t2vr8D9s/LSWrIlqR3RSQw43NOiHmXkMa0JYgPwAVeg3uLSwiq8ZFlp4TMyw/pW7NOjUE/xCYlJ0
bxOZw7AZAOTD/tTAEonuJ/2LqA0VvlJNyvtw458ilL6OID8hKc6fAVca4Rgv1i6WCP7XD+denxYi
Tarp/vrQooMou1qOPXBndPIAe8Gaglrp1a8L6Jt3BQX2S+tWopZhFitsKRvJppA7FOT32H6KYvrt
tq5sHbTq2mMi+J/yurGqr3s+arTNwdB3ZWijDDlBifbJ7RXFr0tQYqCBjwIPexDvO55xDX6sBfuJ
PACsIlIyOiABparIgXJl255qswgf64qkaqtei76gr2cvYyeF4iNRFU7vsLNS3LvAdLIfLJxzphL3
ziQnz5BccqaJPCHi+sAvQANJy6rgF2FTCsd2m00uH9DeulTP7m5HDRwt5Hu9xhzb5mcpx1u8N10m
l7mhJyw/1KBrybRP1JeLpJ9yXRfhul9FYCO7+JuJ4SfB8t/VQ4XK26F2QXFZlmCqsLvV79uLJBbh
ZmoTagXaHIMr095XK5zl4+8B6XdJXzkK/LINE1OPHouMjX2ORDXUyknOwnpXbKlL6W/SvPWPEDuT
5nt0uQaKL4EU53cyU/156PTpw3d8Wq2fh1H9PIxqTLv+sfckFiycVIEWhOVmtHrofxlo/ElTUIhF
3mA/vu+Dh5MA+bh1p9cfFksio3OFOfVkhoaxAxosgd7VE2sSexiv4kC6roglooYyqcvv6Y1r+DGp
bDinMUyvfDfkpb6ag+MuKnt/XT0b8jWIKfvJ3yGyyEUvQWXKjBSxImLkmAw2xs+LIBxx8EXDQ/m4
ivF7SERE3mrzZvuX5cmxyt95F5y6jf5S/MQg24JM4geHwDHm8ujpx6WUnA5LXIXhCgiRjQrMrDJb
jCS/G78+/+2TYepAwW//8qrOwDHKOVIhU+OZ3nBEHq3p/PGDC9aGTKxBd9cagP+cabAP5dCUIeZ1
dzhJiutQvlFxOanVPDAYhDk6icwXwAEwuP23h4W6ahBvItHPMMb5Qd5IX/9hfFKfpCC4qCHMHnP4
eNJD/gd3UpVWsKbVIN2QHorW7rcmqukGpg2FRTzFxfUKkDr8LTX1PCm8Dmf8ftyI72TJYGC1Rwfh
fKE2WDRpEIbGmYffcW+ny2Mg27I9RYN0ComFeYUYTuCKZ7wo64U54MnDltOjrm3R8Rh6BifVyu9g
349V3Mfyuzce399C/ATjQGgrN5iWVufM6er7jE04qg7jYeFMy4IV5AWEioRSd41QkJhLN2DCRT29
fG3Xw6bZsHhr8XkG/Spp7n+wEY9yvAV+q9xtuwoGInufIw+wcl03EXC0bWsr3+K5F3Z9QMxLl4oO
CjmPpCjkMUs20lUOb6DC1kCZucYY+A3S4U84Yy6r8id6SxmYDEkfAVgZfZQJGex8ejjShPdbJ6WV
6bR2ptGAVrTTax1qIV2bxrTyVi1DfVeXS/F5UsL5cBnZ85imXcazGisPes71VnCHc0AUoX4TYSYX
l40L+B9SbqXLw07i6HLvfDuseFOm3Fd8bEeN70LaB2Ryt3LA0f076WeOnD+o2aLeIkUJ9jnc9Qcm
cw9B/wA7casFwz69GgHCzLQsleQXkQ2rps8Z9fpcIuJtWXuIGMAQ70hu4UGJtSK5U2oUnLSR27Ur
sdQLwHuATWGqJIAO02TJK6bWjH85baqO3n7FY84528EnCBBrBDY12L3pQ8ZMMMl6QCephA/0Q/Bd
szxT69opqzT9h1MF8Zz++maLJ6hJ2EnlYacx/Hk9kZRp2CxifnRBf1bC3ROOyytN3nZqMDaxmYhc
c8Dj1cb5VQibfBesTSJPFvK95m6XWTh9dHTnX7wiF7QaRIH22+T/nMOKYZNapVlFn4CLaeYStBcx
ZyrYnXP68sINLy9Bc22+tRk4OyyZXiy08ssbU/IetiYWsHUrHtDywVX/nOhIPu4ipVjH7JspigUu
kXskMGTCphDZD6VahHCx+WzTTgXuQyjC6XupfRYzWh/mLK2X3YNzGgjlQXHABmor33aqHeDO5WM0
ppz7HIbbbCuA1+P2RthMT2KF2aliUleiRt94RiI1IEgHQX3ATl+US7rjGijZsKiDrERzuHo9kqgy
mE8x/EsoJaXiOPIF6QFd4YdGWYuagX8+V/vfzS78VkX+kfG7ARyT2pP4LtGCVNXB6seYdv86BuyH
WaELyPCRVRNg2nTu4Tfne1EkbI3/ISERD4JETE8o2X2jaLAvO32X+xzBBsQacxjLGZ1BSFETqaJz
BbFzl4ZPLdYTr38lC+qbf/ksEDXVben5TRYJJE5qL7WwxGkU59wwPrPPKWRcdEGXAECNACWFSuG+
KJO18wG68wqBHoHwlRtm1bZFy7oa+EGwOTNiAA2t7DjIIY3CMBdwT1oXwIwbseuEpNyWfHJY8onA
0xsz8sL1ahNgR7EglWMFtbVAqctDdibnWp06dsqZWsabtB83zEYIqCG4UwjaWN845IbnWdUSiwvz
EvyIvu2wnE6pbwvc2DfNQZEItj2xjHKqwy0ksGNChZQdB6UVAyc/X63UJEUPzJWnA7pSVwMsfW5c
ZxrgvX7O83CdBWoleW/XAlz7SX8/iM98S5gdGTXTOsBfErw5wz6FJEwBCmGXO8R96MtV0zppt7Hu
IwDy1IxIkKG1t24RkV10bVLcY+KghxyxPMj9jDDv4DHxuv/LEghnsiYnz9v6LPgk7PJsmUGIt4s4
UZvddfOa5e6MLnjjg13j1KuGoux5Dxvtu3IoCSK+PTynqFj15uko9dYq/zFLZm6FltN4qRm2zsKF
L6xcoIa4kP652fVWkd7lix2Nl/GsuA1IupjCks5/WjryynPLD8fH2xzR6niSBmZZeuEkfbF+2k33
tLv13V9yfH5tKcmsjc2S2ix4+mbjU8Alpw3vfbldVPOif4fo42iVDNG0sfXYS9Sr0goCt60hs4iM
DSDjfLd45odZludep+I8C/nb1u9xbGeXvf6B7do9X9iMYlLbxEbzBpEkWmnx2B7A2mubnMZB0Ega
i8iKYWeYXi5qehGrZOMiRGZibDheaRJxuqkZ5TCizwTKmuCCrXWpG/Jmo3dTspK66CqHfqXQOEMb
VHmLc02ZxyTG5PHyhBMbCu55VZpDj/WO/FnmfHJN82l5dC2JmP3HFRVdBUgnLZuQTtEvB906aHEs
e0bvBB+/VmOYUuMBemOnI9+/KvKVYO7W1/jenuNv3W300cle6Lyq0eCLdRG/JqFxZocnosn4HZNy
5e8PXgt04xK8U+07T/6RJBImKF4fIpM7PrpjvNe4UcCw7GQprBHYfCc8kviyjJ3m7wGXwgnQADU4
1yi397ISDST45Jc2YUO9ArFnCc0NqVVK3QWOcKIoyzW6/rnkZEjM3FNTYXrRrOGOIY5eNGHecK78
mUO5PlSa9rZ7ZZeeY1igGlKjTVFwx5shBMOCeO0s9x981eFPplS0iCyHEqQbHyJEgD0NR7Yb9+l2
WH7pGHkE1LIX7slTtbeCzvHAdglCmR/vmJUdxSRPIznbDWQxAKcNzpCiqgI2LP2NhXZgYUUrslLw
YHzKA/3U/OP4OrrVplN8f45jEUwOn4l34PT/gN9b76dfO2ucaPXAIzIhqUkRPkSi9EiThdM6jGs3
o8QjBNaMG1S/3G6NwWykSkYHcK1OXBNBwCk/oyK+bd5s2eoDIlcGvay6x79v77jE8BieZF7XNGOX
NWwDA3HxP3oQu1cWn2nT2yHcdM/v33JOvPydvZrKwDrZUXF7LkSNDamIUwoGRj2Tqh72UEwafrlb
2X3zjHpWmz5qlWXQFLp5zY3cO47NMETe9u8KjiKhX6H8WyrGmSLUIuIlvYIe3drm12GSZAo7GSj/
dsgMXn9OppppFqxmLO6+Z7z0zibD1VtOPRGmE5alh9b1dme9TOQQ1gzaOK9yK46jNK/Ch6RGy2Qx
9UyV2cSj+lwOD+iVhSG2l1gtABDVQ3sPPvZQSMTVo74O5K2tEvlCiDGXc8DahCcXHR/TvAkPLZwF
FhjDu7A6v8lE5xRdd/3tgjDwqeKGYAtBF1EUPiuQZQg0lgucYWuzEMtDa/KRkawtp1Xntqqr7xCi
OlMpmPlf8rHPxnzQNMDCxcoe1zi7p2fcac9tl4scNQaC1ksjuvsl09KBNVzuydL6klVHsQzoi8PI
N9HLnF0cS5BBhIbEOl8AUrYqItJXtya2MXcuwDP+6TIwlcstQv/mc/uCVla5XbMd+2fF29jIuxKB
YxdeWvsqi6C3krfUU9cnLiH5jkf/YTauGXtHVHi59DLaDatwHoqW/xObSBFO0mS/TWYaGlUmARy2
jsLru5nOiwQ+INgr7QRZSCbLGy/VhCpA77PNbXptbTiszE2kCUdVXKrB9HNimZe8i2cBZ//GLgMC
mjVUWlusRvuVd4i/fohfi3aUWl3hAh+Bf6zg/4bgfbeBWNx1IXhmmtwWnWBb4IjO+nsYZe8vkTmQ
4qLl4ZE//644IyTa7YCGHpdxYVr7KAeg+BEYR8ERulgTEfLRQfUORDMw8/5omk4t0U5MMSi6rvbu
muTC6z082TwJ2OZ/H7DVBVHWkr1+QKh6+l0IHF2eGsLcwwtBl6UOepKT3y9U69H/hh6ogvN+DBO9
XBE5uC7azfdZDVjEKjtqCwUhRwnE3I7qKqjr3q0Xoin+ZNhr+aBs5y37GzFh2v9kI7MpE0/8Oo4J
t6K2t2rndBUh3QuVPHx4VSB+kjTlOhQ0FiFww1bmQKBAyaoI3xHDUGMwBii8HHGLZJ/mErukpdXe
f6/8a2Zq2kk+gGEM4vV+GIerqXwS8kGP2MOgPWiudVPpdEGlK8HLdxlYQQfXKhtqrbK6uu8CM3jH
/x1hpo6k2ZP6Rp01ynLr/A/vdHENEx/M6nqG2xFz6TcJ53w0AmUSgN/OSqiCuLhjUdsUHsh8iHDR
2PISWGKQf6MteB1rcqwW2rCdYg2NXTw8qBU9KO6YRiGgKjnrww3fOL95lpDVAz5jVxGqLi/MrwQt
Id4bC89RCYivKIrjhY93BH3gwILy08kEmsdtitgslLtc3v06wGSra2hUwCQGlq3DcY0s2IBV+vUE
IEqB+aupd8mMIHOgLhzgW7N3fahiMalAm5QJR56CyxcycBkp6dz12i4Hs2Xe8Q9ux6wHKVqQQuHC
UY9MXMTcBIgAvVNAN2xcJcp47P5KlMxtbiAYULXsPLyKf35HxJHJGUohJJYMCxXA7DanPqgHR3Eg
MkEMhR9yLPLxs4ryVsFS9M6u7LV3m5Ft8jvwyCCAfogCPFUPQkscFo5cxba+TrbXdpLnk9bE6Jk7
wIgpX6WBcIN5qvxBMkslFOy9NFBykGIm6GDjkzf3L4gYiV1F5/SkeuKeZ1Ppn69GGx9wOB9G8N3s
LhyoqausxA0eACJQgr9v9uD5rcAzurulw00xbZOl/o4Le/cgEiwvdYWsK+ezf0MIvFwaIyja5YUb
7cyTHlY2nN3EzLzIv02VCfy95Bw+y7kNSPpOc22QDbU8v9cKHOjHpzsTWDOsVl9J7SevJoAqT3Ys
zb8fyGyL4P9VV4Wg8AqQVQlKQ4nVNrPAZqpmD32LfC3/JbLYnG+OnV9FCg6wJVPEh6WOQJ2hhzbZ
e/+5Bay89m1gDGrZglPV4om5hn5Xed7D0aeamLBgmdG9Jv97/zE5Fc7/vjafUUWhDn6XHHLYfzJr
G+XbOnn6VR2luDd04hsz7H1Wzk1rzEWy4mcHrHCJrwsVY9P8jd0VJpJ4o0umF68l0ONu2P2zzgqb
uPeLj2X+9jBXKwNpY6clcyzZtjbzLWNfw6KTnz7IZ7itnmDsEewfaBNJlog4ENuu9i3thDYKpJwd
TgdbeYFjA9Cgxipcxl0Ay764yY4fWsVHgydxwD/ndErmnlysAY27XWpl1nSyBNG4y1L50qkNhElz
TE9GZ6I8PEK1TnVlWR+R6in5Q5iwFJdAk50qT12yqtwsZG3zocBnNy0WI1An44Wc9AIvhPDEdYmj
qfhlQfjLwY0ni2ZMNqE5WHTwpou4+p6KSN1REylFwTenczbrqA+F26GVsjqJICxmz19Dft4fx0p8
WHEKXEulAA6gj/a/mAC8WxPCvi180NNyBk1Ip6LZNJsCMChnFUHKaee7PagR9hoAwGbalSwzfSHI
ql6GDibPmc+fLvzxcu9Rjzpp+fMBnR/vDJOjo3uX4qyi+O7A9RFgL/VrXwO4FnEltiQX7UUUSUBN
d3tATS+HPt0weezRCxg6QGkMRzKL0FdvaMCWg80XdPlhp2gU/FYY9ReQUtgzJmLV34kjZN9tGr9/
phXG/29ouFfYFNZsJh4IcP5Gzw5fsVEDImbuQQQQanelTHeivr9fgrimVulNLcSohglN9Yb6x++0
AYpbAf5rsJew/DtqSfp2b5fvlO41HwS1Nn9yg8xjgzBhEyr+JZarNVOHRm+pABKlfa1IcZhDjleb
Tg5FCjpeCiMupy3vEwVVg0law9YGZZRnYW73NI6PEWt6HhPF2qnNxhIwcXNkqjEcv0XMlUcIpyaa
FgEWCv37zYlVL8stThVDm7dCxq6S8QfOFvGnE7DGP6xEFnWpz/G51U+ABjla1G9+xJRCD2V0ie27
3E05xyNTowbNZepgPPgcXAA0Q4cMx/+YVCGuCORNKxVaQS3NvpLKWRkZtTD5B/mD9cAfKT29Exvb
xiacZgq3NwJ0TkwmD3SxRSykMn+PO3Q2De+CNgV7ORivwDPmA+EWmhfE+3OFqwPPCnSIkdQwNgPV
/Jf1VM2RvGDXTbQw2BeiB4Vxikt5eWEy/5Q8gX6SbiuZQU0yGIjD4+M4XawUyx92DXUZVekYIpn6
abPLoHyhxMpXg2MF4BbPM0lqGq6Q6xRSF1fdG792PxOKxj2P3Woynwy5R8mRgzeuj5wZWbDNtato
XlwzqjiCnY1H7sK35GuEbYYr+vk+5teWJK/dZ9WOvXf1rCPPGYKK/AKjTHfj3ehErdMn+DYKo171
xqmRsUmzR2iqEx5cKIVU7IY7dvW54OCXuAZljvWquksAEVloh9M7RWXo47YNDXwtHxPdZvmOWrv5
Iu8suqCeUTQBdHXVIn3YLTiqGJPltF2Mfqwpwo77rIhM/SF89D2Rjf7MfJu2wji8WHs9HWZetKqo
BCQUYJOkwej0cKwwOUZTpiXrD5kwTZwxBPytMe78Zu8vYUQLyhu+z6MhzF6ZfEzwr42Sss5Z0gk6
BA83Gx4Tnu84jKwrLBe+0C55/PAsM7KcCZcQwZL8+XHNvhnNEXlase83H4spSYo8Bgqzr9XPjj87
wCyZHebu0ycqN2HEcQHVGnou3FOFq/5okDAlkXL5ipyvPo0ZSKrUUmS+IidHbE0GlnMxDtRjlfnO
TAwFAW9dhkT/OBB0E36zpPqyx+IP8ZjYzMzEkbmKzyoftHgmgrp2JrtqvFaUaH99VUjrx6e55qKm
ZgJcMEFFCK6eJ85bqQPbpQFtBGwCF+6Z25g/5e159dfJjbe2x2hdpZ8sfkH5DqSrQUNMa7T34JeD
CmpPdATwKW7NsnUHZBuykR1gIm4rEktyuCBUmfovaW3XcP4Gc0N3ekuB4tNkW1iPypRk4NlEb/uR
c1gdBbx8Rz7PQWt3iIWbu8FHh8cjGHhfHDGwRVKGtaHltcp/4pMd0fmnoudQPGg0MVOIhW6B9LP8
rhCIiJQA46r8zFQ8DfGTlHbc4zWKFU+vFKx+94QJSEnU/xcizBJDL4BIsL5fFDRgs19MvnoXfJJA
+s/GgbSNP2tGz9Sy43w99jCqQrnnFuTBdt+M38eZpBmzssOYUM7hn4GJi8IOF/LL9dzzmWa03ZVM
fctUnqQMRKCnJQWVzDBhEinVkz2sXnX+RpMy2sZaghtgTFbOqLHSq2OxMSC8IPMhzqPMa29BtxcK
t8JdcTeKpaiYzp88QRd/Sfabw/L2SdjYUgoHqvrTddZoLfFTeJKYgVsltV5tCR7rZNUnBaEGwF9B
uukQ+AjlzbKeGlclDmPLSiwjrqT8mas/1zLqkrtKicmCLRy850QljIYm3qHHqrHWy3hpGE3NjHFY
CLbNBgm1IFn/TTBRumg91/oXP6Ie8q+FMKZj4fXG6sivN0l8Bb9ZTLtcnnjozLnsFgQ4exSiXX4K
rpXlofAWJu3wBz0sO0yl+bZ8r9ggDhCACXysu7YW9k/3/2XNzT6Ht0+wtE06W1PkCbm/sL4wQpTg
bTRKxdWVAQW+rSDFa3vAQuP2IXiwInoYV9OIMUL1HViB2UihESqRkxwIAL79YSjRVEGqzpWI+xx+
9sfsRrUuDfmuKRzoP+9vcHLJILAyjEHHJv2pT9bOrjKIcqRkgZ9FzIe+lUxr2qK2DY56OhoM7/UA
yDf6P2NRtiP1C2BvRDO3HrCuuazh1LG9LspNPfSWrYr7RYqzJ7h9TaRdDAe8QlLKlBpCWIO1eUhc
sRX+gWIaTx3u2PKzXoJiX/96ACAwhxYJsefd1VOW4vPuz5gcijrx/T5B8h03BFjbip2btlk9GF7a
sQQqwB4r58VYkcQ+0Ar1sgAbHd8tDJInzKyZcxgPi+2mjqVCeRkcEuAU8l4011nIa7J+FBrGb+q8
SNoGAWUlgx/c7xbfOqvLmX/Rk77bV2F7hBcBEH1J5U2KB2al3yfvxqFijFBXCDLNC0815HTPBEYM
x6wlch2f3DA1swcA5hS34iCCa0TeaFj0mjEqK0g4EwIZmuOOzQDxu1XPgXm4+M9TrliIyWEvtbnj
UGbCn0vmfDE/WpGCjsW6bslmrLatDvn5rWtlHT0rZnQeo9UDkgY/jqwrVsD82pM0AY5tLQkfMkun
577awIgzwHcIFgG9obpPV14W8/7k7xDZy3qMZyFao6Nts37OiLTlX6Yefiu+BbyJ/7WMPiN2hD3P
RDp10TrOseywWhJvVQFbOo26MVR69BflicVyRcEEE0L9TcWd2EpwkAIC41wkCGbNKfI8jOOz1Mx4
T46OGmrJNDGwB0PZ7WNttZH9T2/2xY07MDnvZdmxoraeNMEuY97d/1gA85tIv9AaIBC6Kmc9MCyY
AOI8DOJhrxyzYsDOHpn9BLGhoraj7R3/+NBs3naAysXj2ps545agxvynmHr6RpCAM4tNOTS8pPCE
MpdZF78x6Z4INgIrP9ffI7479DZ39m3YP+JKBYBAhucUWqcxADXQXqOJ+aAt4uoG9CHfcj6ycg8j
49fyRKpk6RhZ0/2TXyzdVl/VDvfHPfLPV+jw+cc0yzg+ZY3f5g/NeqYkNl85TnzGHrxnfFoChs4C
kPjt+1eHP7apCKM+Dl4ZXXeoP95g6tGQ9u5I5sY3hIKyUks2aLaYSMGcd4Vtv/AMNSQTXDpAcJsV
jPOU/64ZNPhnYbpNuB71N7USaaXpysjccC+NYovCI4Vdrx8qVRZyXuBxPyLsYK7X/SYWLR9zXC27
tKtVcSU8apbHQiLhHQ++GPS8JCPDqQyrXZJTMTOZb5vmo0cpWxp6VwdYYDAvn2cnGS6r5yqI4NAy
cnq15C51wkvAyqCMTuie95CqwE7VyAapis/Z+K+OMgeH2kFtTeQJPHvLUHMtEgnYLmGrXt5CTGms
ng+gh+34QWeIEUzLw1p9f1WJNhs+vfh8J4fkaVPvo6XQSAcSWkuHK83xSUwckrKF8mnGYQskSxAY
I7r8OfT8iSeq/KRCbqSSXW50qsFGWLTewzWr+Vlq5N2IgwlUt3TbXtL/46K2J3nVdSzN1JUCdLgp
d8djxdxZ/iTeQx5E2YIQyttvn2fC0flRPJnHsyompdNLWte4ApnLkTIYjbwWShVctwncdHy1S6ii
xqnSU7feb8VIV6R4TR0H56wslNjyAqtqgZyTjvOT9DDy0QNiGUy5oAc+yZ/P6q02AUHk5wko0DW8
Hk5sOFRCp34uWKTgzQOo1rJMLDUdzYNR1kjQPpsE1GroXQuKPZDLcE9P3W3z5ULCjjxtSggyu5yi
Q5/rWvbo7ijTbjbMkayl00NnAUGx6q9H7rGQLJEOPuwu8MmyjAOazKB4dovH1Ln0Lz9kpmix/SEK
4rvei8ldm8mp7hoSdO4L17BqF3aImj3kItxGhDpPtLvNb9+PWZhpOT2MEGNg9L3yaP8B2XEADQYy
4iTwAtIsoBTPfFUS2jvSXpDCFNKzkXoI8GhlVdjZKHHjpLXIbLQrN9HBew6vi8qtIJo9BiCPunIl
lPPqDf8brUGpXLG5V/UVMWCtFuMV6fRVozdLygbNiTxvVueYEiitxBPibTgtHhfEbP8wht3At1Ai
mR2K/9l8aj1SkF331PRqjvXpyRkSicVoTsR/871HlDhoaA5EQ6xMe/60embs2QwJ9gjg8g3Vucfp
uc7TTvbgPTy7Io2/ZyN4UiWmPTJ1xemogghdUck/XOpQAQppDbJIcHS1ZB9B2qSYlX/PCGp0YGpr
tS86H/Qi65PoWH+6YsRZ8+huaBkTrNLhQlo1//KxTc/oc3+Pgaj1yHHGUA0NsBqvrVgI8e6kBiYr
vzqt+i9IYiEVOuLmtL+HyW1zuwbHEWKqG1PLjyQaBMqotmq6lJMdourS5PqW1kmp5P1Qqw4/QR6x
lwXprLjM6jsw7DmrUru8vrasK0cZM75naWe3AAO6iGHNIDjurCbx8BRcBkRtxBmKhFy8ypAwKON5
ZNS3mEYn6apWpcNQS+Vns9Mux5NRIoSo0HMbjJnaSUXyU9HNbW0w5M4EmwEWS1ppo8UlhpnNe/BW
FjVTHQhZ/mIj7R3OF22jQ2d5dLQ9vW1NMpmT0OhnRZj9uP8oRtpmZisl0HOFReVh1PiKpWi5twxR
poYfO4wf+hKfsYC5JagruOw05lgihXIyArMPZXzA4WPr3UTj9OieMzLZI+jyOZqy6/139Dm0WvxT
pliob888yyx6U+zF2nzBEnYKKObHLCQo9JdWNox7kYnIBia634Im48L+CzlqXe/qDf22uBEYin+x
XYyK8ahCll4ImXJ6V48Sd2HfZEYfyj+5DPM/MNL7iaTVO39054FCYKlsrx6THsrdCw0i6d0TQtot
9Ekpy5VQEFpf+xqmG9/jG9zMUUEWvcrE7vIt1XrXAprG+7SKKszOjXspJsbgDC4XPJP7alEHEZDB
sNq6jdmTcHbJ3/yuMkTG1Y4lxAvmzO5TFCPazrkCwQyUby+364m0crzbTxtk9v651QMb9+KxHFYl
29AlRr5y3A/o/90PVe/g8v8WBe9yMHAvT6zl1Oj1SwauYhKOl5hnpgnEnByhygZDWV4oSaGSNYtq
bKUKBUqx7ZplRcMdZROXB9iRiKxZpyINlH1u/esc/IoRG+96Cd5YqYuMUMwCF+B2ZILfq360Ye2c
qKMyU6drJQWgf5iDr4UsW7aGpWzhkhrtWIdngW5wKQEjshlfEXt+NxHA3944uttxCQ+as9Fu0Yj6
VRIdS7jWwvSlcJj0UP6yvqwv15lI1f2mBMh9+TGHXJgJ/WfawGgFsNipzn7evQ0k5tAD6TICGubR
SwZgBBDU8XoMpWDfjwCJTfE+SFD9UyjB7lluEm5qew5WVm0v2TLSeQ0TpZb75rOnVA7dXSoQqqIq
H3Y2XAibtKD1Z9Tq+3Q0HdLuVVSq1loBKEUJtWsQX6Q6z2SIsV9iFdr807wtUZlbyXMOJ/toNFkU
/irdcjeYWHXVbXEYout6xjCT0HxrIzGIKKc0ce/u2T2NFoD6+Hd35oMukYvBfSVfhEJ07Gj62KLJ
FtWtaoSYeelu6TWBvSMo2DbkYZGd5Wx/a172ObgYLn7K0fIuHrTWRlWDRefvzNGdBivuVvXGCd0C
z4DdmaeDhXJgynp9VghxMTqPs+3huvJxytyBVFJHG0pPBRrcOfy2RycO2f9xE0wKE1HptJ4B1pzB
b0i2ATmQS4vK4DnuG170q9g/7cmQlHz7DuBnQjEiactDiZ2qxh1jka5nY5kbFyKcJQO/rrPLaHdI
XR9vfK/5OlAn3oB7vKqUHUum0QkDHBrXSNXUxCTnVs5qK467qmwutbOak5Cq5KHdajCaEbwwIQ7H
dHV7gtRcNY9j1sYAQKmbNcNfR7jhyZlmGLvnJ3CCU6carC1Sxz+2aMFcC3IvJHytUhmgD5YZluBa
lmjNZqMC2fw/zOKQWZvH8cv0vXTwghttG9Ry+DpiGnb9SgF52Oatk+V5qRwSNRkNnT8ze/P1kIVE
ENk2ZnX0Q5cwrFTB9PIYs8NiMp+I+VtF2FxVyLQadtPpFhC81kQQVWwzFn1K2RnaRaH+CstqaLUR
yNaWnW1/nB+c+C5uvSK619iafMZD8/OxuaG8Dvp5WB0UzKb3ILwVvCvj+kD1XEjImdZp6kpXqxC4
x5JLlY57XaWJa0W2HMwdAjfmCIf+X5IUNHrUJwz+DGxwpBvHb8c77OECwGAUcXQU1hRGX6Rxp4YM
SGGifaEFzjke/dw8eGHhFGEshySwqefCVrh3FuzBPJIhvgCQnFtm5Rz0apf9QVg92M7WJCBb6nvs
YV0WRD+cPhwL5nFn5g6ivybQgI82LwX7GpsNRXeNYCf3ALPUohdCHMoFsf2XEiRNHKWvc+47KDmG
AYZgDRju6E9EbuX40XLCs30tGDDOze1TrS/vLn5YX01j1PFQNYHq9+2GHeZ9e3gUCjImPk1XtDDl
/9hPjOlv8O3rjQdQqQRZ0AmDwEgJmnnlHAx0owXN+4kH50eGYghc/B65ufii0JdIWCJm2/Uhb42/
pLtwLmzDCUmwx5bhCl/cwzpyVVD9w0FS1In1ZqocWV4UbcK5UghCvzjdQn9OUYWd91zK6//+QWH7
2sHIP2ddLFPfB41mKWYQf9PxdjxA6tY4iIZdos9yf9T1c+i+Lxjlp+WxWchEeiFJfU/lbHYW0rCr
bKu/MeuLsQYy7LyAvotV48Qjx88Mkka9pgnmHxUjc4rKW2gsrHNfuBE99Wcq0pE7rGWB717+8hpU
W7D5VZ+ojjODtEkzH7Lgongf2CiuRuRu0szSTla5Ma70jcSAQRQNOdAAFL27M3GGgBw7GQb6m8D/
PtzGNJ6XTNsRXCLZ9Gp6jwMoaykxoljUiYvMtbxQt5Ow+JUQmKFvXKtaV/H9e4rKLp3Q45Xy7yo6
cM9LOU31B3umQLOJVmbvCNqRCmDriOtaf1ph9+cR39z9kpO5wRZv8avf1V1I/BRmUCZY01hJ7RK6
WatuLLQJnqtQMK52KooE9zrH7ixbmrJrcVTrATb+agp3j3qOeTwFGVOGbriG4kIVXN9G/v5JchE8
miuJUUalX0t9oSn0zKwMKnSe1NxlBwaeywMCGbIsN1FeeCo62A4Od70d0Vw1Nt8zoFcMUjKtLXtB
HoNSZ06b23LPNExxdIHBQu4nL9SPWPm3QVNGcUer36KaaPi+dx37YxxVA0qO56zouRLySTRa2ZQh
DTNkuVVBezxccu6rB2XQnGr2gtcK9yWHGWSdMNk9BcOawROTD61x5gxnwnW90r7thg1Rb0rIHE7b
Mi2pxO3MABsYwN+AftaxVSGpCzypAJJ5Ck0XSiyJgcF6XTXUx69p5nvnJjm9AMfnACBvBtpU7FWU
ibZx1V6oqn2Q3ikHFzEmOz574ZtryjnnjGfYaRpn2i/ZF28RMqUvp1lfhcCwK+ABV7igPORzyHiK
CRzEYxEdaPir3j4d9HEqS3tErBpnNUEoD3mCTgyf95Z3jvbb+kS9Zp/93vh/TaUgGoGBK4187tG7
8QaeAIXA+xrNINeAJ5+8oQ50UjwlQL4IE7KBGTmj3rTlMO/CCRuElWe8BZBiwVP3R4qbrwINETYe
Nj2kQNHWFh/eH3GceveaArx1coK2+wZdwCt20354P6Pqc1edXAXsHWwqkAw6Bxj6m4mEv/+hdzlB
vHCnJV8jZfzbpl5v3Grf4sb8bxCmFtTPm4I5o0+F7T2tuJ87Cglo/DSQ/6i/AA3BHljL1ZqH+Ip4
a8ehGgompM/v/Adm+hJl8424wwhEQ4RxgD/dutDzE/nZL6sWV3e1Yw3Bm68vvGoSO/hem6fUY/xG
Z2ehQ5mouHGXH8j1h3TBcu79Uy5J2U0RwSFLURRglrLp/h7GDusLxniD6fuJda+ro/KElqq3FVQ2
epcREnQRrMTse3dpM2shodb3JgrJRD48R+rXbN0nQZid8ftgz8uKg9ZArWIfy6+EDpvLj73IaW/J
BCJeb6mPEqsygMDahlGBHVpNbIlsrb8GQVu64eIkJK+M+ADbWh3kRmUJDhTGljx6eNJ5X/HSvHis
avWiivAp9PcrEdcsJViryQUJaBlV1lEIp9Y0kQ4XGoyt0s2AOZiD1Ln/wT671GjcYHpomGn433hz
AXU966leWcrsVglkF9S/962dUeEJWKj8shuJ2qTv/b8iUHEOxJSba8F4ls7bM4uSliYFfX3Ji2ce
m8p+AoyJ+unIliO+mVzYSEy++kIfoCVduP+aIwhZe7Puj51/q1LhhLHCvGGg6+hl6cbDzL2hDUZa
mef6ntqISgzAaAbvO9QE8xjXfQOJl2KFLN1GISi0lpP1UuIHE/0MMVtwW+xbJ1fXP+EdiPUPfFWF
TcBfG4kbkFX6QRO94YJKHOZMzJqxRv6ct14Hq5JPOtR+kG+6SBDlbBkAJChsm9yI+IFexh+wZHIq
sRzc6FFqtT1WHGwA3I13RZg8XSExMdTb1kZsrZsSiWwBWFKwWS4tLTT01vj+72M8iuFdE49HOFYa
ExMMux0M8YnorlWYX+MYq7iKMaefj5NfVA0bX3DQkKSahTqvKL4B8O6rw0ToMo2UruCyHs4iK3i0
ExYd7CRCvoS4k6+jUZ92lHyvVZXqegW9r5VX5gm+H29JFso2qnzfBZEyqQ2mlb1KM4h3IIgby3no
70kOj5u9L+nbSRuqgL834Au+tNmCNQyvCT5DBOW1YcpVzs6W/t7OKRTvYdjMMvwvcR8cd5A3b3kU
0UU6QWocldEAD7WfQvfF0EeeTLnBct/doHltGpKGHlwU6P44ifFw7nVNANlGIneGF6B7MzG3ZoyE
7NIrJHkCvNXjGDL47dq1brBt0iBzgKEbJznZsHjMYhZj25i4fre6INhMBWIQpU8GUYCX2amKqIFx
B37cZl1QRMNKn5Pk2SJeJnnXZ7n45MAGNLyhjkeoATSIJLNrGMP4x4oT7cSSMAkuC+QdzaHJUT7D
eEsUXyZBihYlc9QRXPAdsw/+INbHa4RL7w4fPX17YfV47jHlZ0PYuMknuznjZ1G+m9+SMPTeJIh6
6luvHpZhXyILJzaIu5KflxJ/I/Do3ROqFpVBZtDirLJRZm9Ib1rCIaOtX6pNtkaiBj4q4L5kx685
pX14jH8Py1mMqeTHK42+3Hjsv1+wPd6p0iOQS2LownHH4VGsieP6uTXdV5NWFjwUoDvxcymInv6v
Q1FUPYDH/iIHKVNgJQPtxrCARh9waiEkBq/BJGZ65dn/ImkBa/s4yFWwdXyEt/pR5X5wrIf53mO3
iEoaivNcD9WFSgFPF6Yj2S98tzyzp0AdlEokGjhrfK7IzYkXuqgYHoUZqWbMnwEG88Zn+zA4ZLv9
ApCj9Ek46BbXcvLX4Ju+AtgijkjzYXD86aVS3aSXkLeCCtoBBzpEn5BtCpBczshyj/y8TUOjTzUv
XuHPX16tkEtswZyIc9Jq+GQdh+/QiOUFh7pOMsj8X7kiXW9QlZTeo2W1x7hVRo0je//QaF1Mnb2n
9pE/7JKTVJjh5ga0v2kZ6o/R4DRExMj4zHSIhTwId4H3URsEMFwtBjbnm7F3aSUovlx47qCcgb6K
km4KhWnf+l/d6o8CTGBkSwiYPaE3zfrKtqu865gCkxYhid51+9AjEKn+FVPDm4u5eqe9LBnUV2R3
zW+xtZwkFxohMh2qjNddWngdvIqoesGo1SgCs/pZUBU8E+RkER4Vc9S/be1zSh7LYg4uMPZaoW+Q
2alZiyBSG/t096yePXLzfCyJeMQAe0/GVS+KnR8reVdNUfEzCpnCvzO6b5os56KPnaIuqVicZcaA
/dMSGGr2d66hegC3W9pIXJK9ko6Dm0wUbwSMXzh/BOJaVutpWIOEIf7/rM636N7TWF0DZ5LYyEJ/
arGrFfVycTZ/7unUQmPAGbO8yXZ+afMyacrRupcQAjiW0hl+LiRR4NLH1GigCgaYFLLPVPB4avrj
V86oBOv6dW51/72QkOX0ZpxrIsdE2VHIEuTZt+g7/quMECg0ZncuIpnO24hI6VF51Mh5WcuxfS4h
hrHi8QDLj+AxeBwn8alrWvCec/qStLCt6Hiz9bG0JRXOA/gGmeE4NKxH+jxzqw34xXST6XEcb2Y1
+itDjzWPsScZy1m9wPa42mIqb0i92H7UiVAo2/Et6Inw+h1prBouUWkIUBCdLphFe0cNIivxqLU/
oHyI0zz7xUYNLry79vmcHFCq2ed/AqzLY1C3OH6lisZOzvdE4aY99Jeszg1SrQKQ6c8uTNKwUzRp
AKTSqrgWN6hGQnvwlBn4WsGygzPmTwUDlgvdc7KHSKR7nB9DRRkijfOT9ihQtW77OynwKhcuapkB
mk4H9litb3TY8hyGCaLJOO2bylO94iL9Etp6lFACn0bbpSFUt5PFM00j+i9fyXzT/ILzhqPVDNUB
sEgEtEzPR2JliwQ7+RDO+Z/eF3rVOz11p95kunFTYxY/XgMWVTzHEU5PwuLQd2E4qRbFNsdiLc9l
7MWBsfW7Na/XLN6Fa8GPcGzdi5HHM2ktqmuYtjxXN77dgGhFBa6tot2F+eO7R8DkzKbBZSZaNw47
IGbiygSBZEMYs7vVIJpol2tEsgevXluS9MBPlknVXZRdaqOanHVmOrLy3A/f7tNYoCOjDQXf8Wsc
FWEsgypC3mXaNNxcdQ6CyCVh5F+ef2brqNdYTGAeZsUvYOekZdrKi2SDO3UwF3O+G9nUZ5KUr9s3
RncY29d5RP2ASw+FHy6d27mIsyDfZFhzAC8mKO+bwDhXXvlqeOS/ZL5AzDQXOMg+ZtBcOeWpo3dS
ANgeTnbu4uoxqiNDjFKjPSOcgJiRhr+JdEAhnUIeFuxJSSxJV9pZ4pNEFK9J+l6ZQ/jy0oBzXGC/
jJlLEPgclmi8lIQArtyqEo5DPHyXXQe3xbH5T2rHNdmAHCeAsn2KgWybO8C4oewAN3eZ0tYHPTcq
SYJpk3uK18Pdtv4cnnh9SqxuGsaX2o4ZpikyvbODj/LFNVIxP5xac4uieus4uOdiQZGW5+6hPQ1t
Ip0k96rpNtPM+NFI4y9VGJWTqsImwoxZKUnrwTRn8TeXa3iBap8WcxlmaJl+xsstDaS/OL/k61fE
z3spSmvzHljw0zJBfwYt121wf8Rxjg0qXEb8eBnYwX4OYgQILU57g8b0ovuA3Y+YMJijH9/oxrLO
XrU1Qj1AEbX8DjelDAm+p36hIodWgde6/LA2scJWVzD4r+BjYJ3NEXgBfF2bNTgmnbV214SdJDvt
BHtQLE4lza/N0tAxF6ZlbuxCmd+xSFyx3DzO5EpiGrGlZieUNahddtWZkoIqXeU1JxGG73+Oj5GG
+LW1n/wOg9ESEHIqX8lHbFz/RwPldbrGBKBT0QrKlKUHBaEosAFgzgGzMso3/ToyFHmbSqg6aBDC
o2l0DObAmlMXgvqPh+0FtQ4uiEXdgNdLVi/AK+n8hxdvbnfZhuXwjkz8Op6frOmT99lcxuoXuVh9
KIjw29YD5rL17JMr1frerAlNYl7+tJbWiCQMLv1gDdpTPDOg4mYa6M49WRs1CX8eowF2EUVPUBq2
GgHxM8krpr3U3KCjD11kYWbXiJykKdWWUbfJrmV7Pr5iVrZTvsJhJJ/uxp6pXfpnl5yEyeIS/zar
49Nd8pWSDAUkPNHxlq6HTDenPmoSuGYW8Mb1MDPNcdghbOs6lxwr6ONbTV2SxULzzX9Zdj7zkf2/
o74IPu8oQo48yRnisgtK+meC/Pws+zXdrS3Zk2yGYFGYl/17voGoXtKNocf6SHpuKwnnasDmyIZ7
cww5Fgb81nwf2BEXtKA4sNTaIT16uW3xps6qCzqwgAaiAPVjmwPJ/sMWsgM2gP5EAM69HET7UFG6
nAY9RnYAScDTVbqB2rsVnvV1uI4WMWuYL95UHoUT25TqRJ0g226AxLLTrErU2a4zQfK7ZDo8rwGX
x629b3pYSjaXWntEXMc7rY/fEhCc/IWpFgwQDaQ5t6WmtwznyWeYVEqSiDJfPKcQLISv6VoLikCN
NqWPvoP/+VcqAfR2lDDWAaf14pFmNgWOsLxGYabs7Kl7KEDoxihREEly9QhvQA659KtMgQFyO+rB
U9Az9gbOV7h9Swm2/BDkEmJ3oe8TxTd/0STxJt6dSTh6+yirkF0HGwhFT9cJKf4QyddPfHW7F/8L
HtLtZ11JAAIQYSnqX9ckbcvcaCCAd7BgGkhtaM29yY7OgzaRhMnfuTc8ZOfG4g5kWIJZ5Wa37ian
bYDSfdc89wmINtA2outvxwRVEggVgm2uBJzs3t63yeygrDIqs/UikzU0gHOHbddYKVqVsjmgsF+S
2prCPnDkPhBJ7RJTIzF02XmtaoLEkQeGMFecpBhSmPNUH6HDtB/3vgZmaPfrVtPEGDACS8SigoSC
9b3DfwfnszbSYxRGJPNqhvSzPskAF7m0q1inQD78OvJfojIDgOc/7/MJovN5kbF43vqLe4nKPP5p
/HvBMjeJ8dtJNn7b1ipPMYmG7al6IjCBs3MfotW2nvmpWWiPYhliHurJ9pnJnWed7DF2p3cJzDlw
kOfBD0ExFlo3RWLj4rrENNVXegRboIWU2wx756lxaSWoFydZ1W/97BmVrVm5S3NxLMA7grXgrMeh
VUwb7UvJd2/59zaZeNApbqGjs830wCzveAI3m7IdPzA6PZd0wZ6OzHb7rrIgoZwiGDUrX0GNvbej
ukJyehpzxGb6weqfeuv4L+qVG1IvH5wKmhLwbRSlMaX3j0zqhUbem/QFoUIwI2dXgS1UfsOHDkBp
XAyWAplDnm/N9+PtqAv3FTHry9GWmRraxQEwcyz77o/0uR7u8fM05UFF1o4IJsaH+ZyRadjYuy/O
IoQ/ZvByYb9dJlU9wtTrFh79wM/VbD3EAWAyCJhseq5XjXirOJ9QnlSkxGDHyU2Y1b5HWdVKygwT
+0/MMrdXrkKQRAKDJmloMlC3cjp3N6ciNYe4/JcT1sWr2pVB60m3XIBdi0oqVFZpEeOxwzo9OV4L
91XYSKvcAG83fz424smTDi5xpPVZzL0U3LadSIBZN8HtOa7UgBJv1oM4HIhGzVZFDAMxcx1D3xtt
oX/YFkGCko54DiPRiGlGQnh5lJ6wRY2EJ7c0Dng3Ryv1hL6Wk1wNqS2jiPWaGuzBNlMpNO11mbfd
dYyLwytJ1u4yeG+8MV5dQUlmyKBRI8I0SZouSR8+/28iKUTSn5ZO7LJUX4FsXVuMyCy1NhWPKwtW
WF6DrVH2+e/veIG3DVXQuHJVVsV9U2ODnM86XLdVmDb6XYTQgtpDzkPiGRqYH+VLA3RZsiu8DRAy
NXv4RZZwPwaAb1p9I15xpHhuqRBdfleR4O+DGn3N4j/I9mlzp7/IGov/nyIS1USC4Lf1jBcrHzJC
rqpM/giaGmBKjCXjTxq9dc0ODipuuhK5LKBnqeHfkwl6BFQeAVDPWplPQX/MSfk0eH4gRj8f7ZGC
1LuJXNBFTA7LfVI2qk2IcxzmxqaU2NdhbeQ03urlzbX5Ltfw0w3c/9yAcJSQZefODxnzH8gAbU2n
rBc3NxPH+rU4RtKiNMItyQb4dFmiC4HzH+i6ZywyYQliqJiQsGubbXYvlD9K3Q/A7lYv7y2In2pV
o3LjNuuax3u/4VXOlCFdT/CdaV8QJYIISy7z6lOOVufEkLgthKp0mpIpJJaZVOnYWv9a7yQZc/PA
nSnebL0xR+6vM6QMRwpMbDiPF0a3Q1j75SJNoJGh3XkyOXbKgDhZNVkp3ZtxVa6VcG5SiP6wTE1i
8iB376WCiPIQB8/uhtKHigcCOLmThkIHEwmafJIArziP0Yyq4win2UWSKgz4DqLHNMruok643toQ
LkFSsruRyyzm7RDVIh6nD8ixpDgMNFMiBFeD3YrTM5jzPRR+HD+x8ILf/Rs6xCkH8z7Qw8uLbCdL
gDnOvo9GpwzM/00fW7kAtTIuJ+8tg7XJiQvP6MCbYd3osalBwMkBbA1eeZXh/PiDC5fMn6WCXo9+
LTwewZq/Q+KhP9VMLwztlHnsCNCXeAijQa/+QDVOZytVvRC2FUpc6CsRu5FQ7ZAp3Xar6okumYqA
B3f/yW23Ahsktif+JWx2C+vnauddY+PUXisV3Mbktgj2YhcSm6EgARWK/HjBzTkHj5fk3gkXbf4S
HiTNOxhkFTUPQ1YEoSEuUwyqfwOFWBR3z4UBsppIkBco4l5GnodmPcVpHUAEZFrUohfrYBToXgkL
BjZoATbgKeVofGDmvAkqwUVL5/ohjigmDI5j+v21Cw7OK2IRXsCNNZ/RJfx3YQz7QCLpdT0nb7ng
HsIxZa6Z6WRCWCDX8Oq++8e/jPZRq/kSeGCNpZln/sBf3vAb//cEA80ZKpGHMeZnG/DJl7rC81MM
B7F/qXJMuHM86WK/bg8lxy9GF3DARWROKsFT3m+PgCFbI/jxHjb+cFkANtTdeIwSJYL/M73F3GK1
NKDq7qIRG/N2qL6XwyiXsV2yohfE0KHTbT18ysd/y1zJCVDvnDSdgNUgzA5ygoLIUCL2TvqIBdn8
XEqQgZI8rcEpQvaTCCanFhUAW6Mn4Bdo9qYQ28VDspIbcqXuowvaohdNCXdozm55GhJZ763BGrG3
UnQqyOco5fKiF4iUxIwXQYy0ybKNGWif4E2O5/e45z5czhE+XVcdj2WItJODrZbkMErQCpa+w8Mh
Qt0od0fFWUfF57HX85Ua1RqnWl0m/1XOFu1fVx43T6YifdMHmVZKgX62tqK+8FYO0cJZZ6YtxAI0
9JnUA1iwcOahg44P4UhfQMdmF2D7m8QQHE3YUsnrNG6m2OrJixE9+fNxhTOCkIvwCTnXkkmiL/y5
RtrG0h2rabHl0fcLyOZBF52QArGyheDv1DFEZThtP2M2WXCky92Ynrv6rpxTk99lKfkHGDL6ztq+
0w37nG6cyjyUYcet6lP0jFgVdF1m0O2ca19c/6Xc0XmpJ+SEvDq3jqSdaYAjSYFJyuwbHehuxg/D
KlGcjJ8B92sdAr/CYM8Ppbb5qticyXm4LC23y1TanONJ+kKjdHrN/TFr9oBGD77Lg7P0MUbwJn/d
CMs7eMjQjS8uPnDKmyuejnM0vVzw7jjIUOUZ1n6yZ6OY1kmi2Ojma+68hIMnHlJ7h2sj7hV4xC53
8c1LFBISUWnbDqa8v4UDAxa57wdg9CpqtrSEr6nzfg6rAW4S71E0KfyHMCYhbKgNBHw6ewvFGBTS
nLWVgUM+CtGDHTgDoDFcTYMcDjo6iKfwEIW+QNLZs3nVcTdcj9edH+HxUe7a86UV3GnBJUi7VOwy
NxA7Fatl4t1ifnT2PZJuKTEcwbSMbzpaq+1kU/beObDVggtQ6i4M8Jl27Br4FPhbdyq/wbuFzX+d
hE9j0l0mbi5cqCDmuRJ81v5Udd5ITlP0w3TYc8J/OHWF0o9+rMd8N2aShxSVUxs4QIK5DQ9P/XP1
B55YyLl26r9W+0bhrjEs1ZZNULTHNpWVj1ZteZaO3VMpWHeMC3gQgpMTVniSPzZdlVUzJhXlVfI3
r0rPk3OknbFi0RUrQDyK9sbB9/O/qKhlvgGmExpZmHS3lHy76W4PQJY9VPwQfjIaVkM4KKKQ9Ftk
mLf6r4YFFz21po6NoHbeLP0sBClo0TbNDMbqsHTx2AkSsRz2N0+g1EQ4zzs2Gfy2FR5HtrlsWbYN
w9l6lG+mqaQhVkhtYnTZnwPgivgNL3LQYDZAZfpJx2WeoZgCgZWJYSrqoOC2yW4dSIH4pHQXox5G
IDEAomRKH8nGBxeoU/w58Jrp4SCYKXDOhW3wHGVXvSdhsFEFQRyvBQgNaNgA8/HckjJOZqF5nLwU
BjoqhinZuuxtTnGvm6dLVx/MhfqI4RAM+fs/plciptURZsBU57mX+nBxbov8paJnZBgn3J6vMIWp
l6g9p1UYX2Z+yn4sdybOt4KoZsmuBuApzxt/KiZIa60i/ycrHQINgHf0uaUxzN3k64RIUxtXrBjK
yFDVRnEqRFlDPoNDYDEiXguC13sfKglxkaLcNX5OY3s9ZbFgfN0PhA6wJglUBNjQd6CZn4b+afGU
riQfXydTw/Bzli5wB5UvbDoH1Njc8TkU4t3gUoeBjzMmatreV4YN1i8sxT6EKBeR1/J/M0j9y6BE
Js7XWcjjwY3WFBlqKACG1P7wsA4bcErl8vG6bJjbmmohtINu25E+z1fJQRun5fOs/5OYi7In8LZA
Q8F1atBUCEWV+FmFa2GX2i0NrGYDgmhibH/dxMwxu52ke1SIMBPKZobPdhYHfLl5lDK8sMyE3D5F
oVgu/gQHxVobhn/JdhZ225YbX7MAAWdgLHPIp1O+ghzSOt4IHs33C8qMl3OHSXN+IEJJ4wbthIku
Mvm5nG4UpgF4k/FL6h62XuVRrQacWcYpTHVmrlaO3g2wDOu/L3IYARfnEQiRPGFQshJ2Ts9Mcxrx
yDyvZBFC6tGKz4EDxZQAW+O3pXXqVuCmJhooClCBVX5um25XTzQFedQ5LRq1zjKJtj61uSTuTGbV
ML/gSph1XEwS+H22ukNjk5JhuACoTjCxu8T/y/LSc+Lxq3vgOzBgdG6C/2/QJmgFkuiA6eHWaUNV
lYywoxQCV3KgykLDqrBqKIUHTAw93xSqquRhLnXHuSyB3noLbuwhbK+odl+M1uKdcDNNATvihy+E
9GVpOuJBPtaOFnNrN9bGeqvvrIsAgCV/3sojDSCqwx5fEDdYzZuP+++xdfhj9vn7JKTlir0Qw2al
i7WnFkQu4G7912oinEMxPJJp6ps1J+Hr4w2AE24P+rAJWjp81Lqe1t+8VWbM11A6Ii5HPPEU0x6b
cQSfCYqHbakW+NCHkGsquJsWjcGxaq+unVYnf7MEpHWYAG1lX14ownIV+s0p5O1xH5oGmRoX4d2V
eB6E2PcU9hC++7D7a0ZwEUnlcCH10U6cK3ZfFhs+Cx9JmLqutFyokO22jNvNfEuUE5UU57xKZZqs
CLMTxfVmOUCuq1LXF4U6KFZhcpjwJEievGEapE4b3MK85NTqeD+1o8dl3fjYyhyf4PgPMpKRvOta
iFs/D9yQikTv7kWI6daehY9HwwFzmjLv6owoflQ5ECONo7PRAgA/lywuE8F+Ioz/xh4c8GyMx2Ba
91rcYM1Dvz0/nEocc2H9GHQXtdia7ul+w6mWQsvlMG+iQKpRtkOngr32rZvRcPhop6M1FR3EWpVv
7RIXLmq9ttea7rOf6U1Pv5Uy0wg+XCHvuuqfPjQmR8/KBIqMRwk6ijJc7/N1rgAR4NoQmrN6Qo6n
oaWHwqTnBmw+lRvQo2j0th7Nr/cy7EzzsjUuSJswSg74FGFPHVYUGfcu50QuokOYI+2hI2xxNx3s
dDddlLqR6TCWpptQLGmuYdJL9DPJuBn2JR+sgpOWePEMjHZYHGfPmUOvHpNpHBl11l2EofVm1JKw
77eRpZIYI8uI9q4PNs/xFVi2dcRvvHt5ybL4Pd/1WULXTuTaLOarWNkZOTJ7xIEuD4CbfXbXanwD
INPTQ9Djaeuw8ih2VSvq1C5rpsH8zH8+XrOr6O8Wl/OxYNN0uR8kNsCsGZfL67xRlgOInIvu5CIG
0Xu5d3ZqvkptYzr/VGWvNKf+tDXyS8JZT+JVGB7NTWb74texbG2LbrzDXN7482K2npPLZ/311WRU
rYyW8AgT09EqM7KbdZV5zbpOt1fcKpNZlmHK0drB27Kh+cwWHoQtvRwonPplKvp4crf+dLBmsLNL
p9BsD9h2JhtZLI6cfAFsQksbsYHsKb879LjyTX0gGrES0ev5u/6s7LJJtUSWXo5D4SE+NpgBTpum
1xRHg3qCPhjfNljgU7sbuKGws6ItwBZI9KnQX85RTxm3MfM31ZnfM30wZP6CkBDCgNL0hCJ+0/LX
vQER4ykjNVB9+L7Q/15sQys9PqL/yHG99mCAIvx5Mq7frByGtj4fyth3+5guAhN4hrdTM8T1ywOP
Bs2+dts2jvIrjP0HVgwxEbrNSAvRsxeOpg/Wv9M4hPakAVYdQD0841fLwR+thYYAZQKeoPT1jfp9
v8mwDrfTXevdAFAfcsk4Pk/RJ+ele9W0sQplBoOlfnNV7hsLsPJEIs1xlLBfiNuffyCwhucI6yPj
LeAnXEp6/7gVP3ydB0U6Z4fUq1y8D3WOhRYo9ynCBJu9tOpjUSQBdqWLoTyWzTOTe5oo+hkPtdes
/AZsfwNxR3vqDamoanoNc0Mbhp0xNypIbS/FaGCiHzmaVTnu8SSRWcsYRe5LiMNrgxDbUp5VF8WN
8liZQxmi8F+RpLDcVLc4KCuk06o6JQGyubMS6OVF24+6LEJqQFssDzO8cDy6NsOO4WpLEcsGzqlJ
IWmSBTjnToYxXYUKybH1vJgI3kH4s4oZFVMD/rKULI/5yQ8PsoZSTs3N7gIJdSgh+NbxvFimD48l
gVNd3vD8pRK3tYY4dTZenwdGh76IFWhlZ4wCpUGd0q27F0QAdwWgRGyuRuLUYtDvGk72kyY4T+WK
CoKBiOnh9356bFKillUIOVUcXVXqXJTtjJIeqOe1XffGaOqzctW9Pf+k5H7TTfqNEN4s45+th+LY
hr9yIHbL1d3YztGxOj5XfRd3aG/+95wBgH5Yt5KUtHMqESlpc7/f62Z5FvTNwD7ljuLWxD+uZtMR
w1L+kL/tpM0H6454Vs0I8yMKEiCQIgz00s3MC0LXW9jS42qxeaFc6Gkew2ceHgLUwkmDRDOA8hN6
JoLI0Ydj5fOtep6j2fwLJmn4cNwKoqvy/uLxO7olUMJT6xJSx1exp8CMUBPIkpMoklstcXYVv3QB
yZnQlwfhOPo/SCf3F5euPi8Sp5Fged6NyQWLwvjefd1hwB/1TJROPeZWPcErHxM2fvqJjLwYlnMh
6SFZtXFKM6NEDVuCPPIST3eLBvPWogLxVawvKEGYS6WLeEJn31xMblpmtwvhxiSy4p08jDqif46e
LjO1Kkyze+JO9A9A05rf7L6QzWfJB0/g222Q/d/rtodWHxaKUy6sQLSnbg47Vv5+jSNW4MqfCDdB
sIojALliAYz17KJMTdcvW4Vn/O+Jkf23JIJyiSqml5RsJd+VRhWZq2xy+54h/tcUTpEGuj7tbbyZ
L6e2gNI2uqQsGBX5ST0OLbGjkAMBiH8mHWDsvvT4w1UUw2dRMzRz0vvotU3lCpzExMa7MNNzz29B
vcFzPj6sMCeq7dNOrJX9OXhNn/kleWp/5Q0Dx5Dx8BiWAuHlaDvFvvwMXjRzbEYOkMVJeDQI0Row
5sQgbf3JlADiyii6qwMYfajby0pmwZZA2lypQ875/sdR+7HC4D05qLiFgUDxvwna2013dRKj/WMv
F4bbjiZuDZpdmmNHb0HrDcL97TSSt1QnhsesBAeng6bASYunowa8s5i4QvtmWbnl94AveOyYbNZV
Vy0oRq7eLplsyrv4biSwWiCQtEb9zKfNZq5Wb/Gib4fR3UOjUM+Ua6+nJMMw4ljU/Cd0uiTmCRng
qb9QeDMAZZSBSfmImZrVAcjbmcHIy53czlGaFoXyBORkJqSuM7M7X3ED3aXOutm00T+dJBvb3Bz2
CFa8VASULvT76JyBKy8RnmVNtVxvqV36gZSPqme2BeO/vE7PMhmPPGs3ofhlrfvwce798anQvR0j
Fh4PBXkHa5hmneKunZjWE1Yi3Lwhwva9ITICvCgdzjgcgvEUSPwqzCLXYYqAIFS1Wl8qxvL/nTzT
79tVJmm8uQFgsykM3QANSJDcLpqbUA19KvxRs9sNBfs86s38p5dDWqnp8dxPeIgsRhgEmZyOXWFi
XilJoV+t/sN7OpYigNS+lYocMpT5dD+ZMXPmiWpJW8DSN9IgMPRPKEAI+MxAJZ1C4s5lkjXjo8BT
3lNLCbP5/oLSKo8JY5sQBAO5DRLUThCgoUnMzgporaJ5opUGqDKcScwLvOZp0X0ZMabxkDjDm8X7
NL8WCbEdxvNOa1/AZlZX5iZNqP2YjlClZ/1N6goy4+u7kxm+Hy6MACVicb+edPD/VCfCpyQ2V1xT
Fzogjygw40eU7xWSuJoVycSR3hZvn62NdJMQJdspvdW2PreFHBP4xHX6DwBCRCfpiM4sE8EvGCc3
cIhZysMK1KhPROKo/XWxZzSLYzboInQNfRU8BW8WvZciT2mpnG9BXi8qEOH52lU2ZBTfiQoChg7w
9LHK7hRHhvOhJHzKe8LCy9c2+9n7rXHhSTdMK2lOfpTdW8KMvEEdBRfxGFff/IhS7Ac9qK/38loN
vdIQgUVQpvRkXaicDy5gJVp7MsIBXCX6y3vtJwAM0lI+o5kSlvAsliIyzuIEDA0y1kFX8oq4SJxn
IB6F9jl6YxmzkdqPM8pkJIQotLi+O1WrUUGgOGYBbG4Be8DkMzTfhw0bs425mUlY3P2qRZNm9wMG
WROXxoqG1QOG3XcgGUXyLZvndPhW6DI8fYxytmpuQuiqZdlyirjRd8wmI2Xhgx47oTOMOk0KNk5i
X/Eac1ySkOyBxptkMMMryuvgjpwXW7uGsPJwEXjsLEmMEbC97/H0HfAmbc+zaylOSWkPpT2Txtfl
HAOwxF2hlG1ClvOYveM6t3xGRGrKiq4zLyypXmKnipVujyqVBprSrFdi/NHcrZJ7CIxQ1I4ltk1+
YnYkFPQQRyMElZ+/7bZAFA9oNaUfgyViI4yVdiEkLAZ3vHczNTEB7dq1z4Cz36HPkLEDaMLOBwhQ
Cxynx09qOpNyCvEeWGwA+/gGQId7EM0438hS+sESs7fPnXhg+mskrfETU+qN0TQTm5K7tvHFOHsy
iu9kviy6DqLdcJPEwz3UaGoYKn6Qz2WDhqPmBHgwK2E+ZDG1NxrrF+sfaOA+DzV8AnOE5eSs09lg
Xu4LoDmDM4GcZHtzkuLVaN+WeJuqScAisy+g2Aw3LTbYJm+2HN+XZ8/SiDdJFYjxAYepxx5SPZhE
WCyLFDTV5PcouwCiqrjNff4Qezk7nl6dcqgt8TtvRsxfOgm4i4vYOMKNdoNd7KDlZQ9kUAsRqDHZ
NTTXlnddLFK3BBHL/LWeqXbhmAFCg9VxosiRb5NNqXSEj//lgsYzrGHZ7o/CZ1Z95+mXks7G0sXY
cDO9EXnYvwcZsg74zCn8IWCP/o38i4F00k2nregdaaRDftJmTGzj1wUTXmsVqDmeWrv24NXmlKc5
Kv2Jdcy9jKPjlmhmBAMzo5akRA1In8/bSCntd6oXaUQkdFGcmyzsyOhgzV67mdJR5aOKAYkxdBAQ
YmEiZuSlLJ9iy6j5l51zzhE8K53gdplYXOB0xmBYiL+q0qvuXx+sg91Jdm0HS5rEs0KPNQHFazpQ
tkWtCnWUEUndLS9v4nV0cl+TTlBXRraxvyteBeErazwvM1iKgCq0GjettTLq9wziOUa9THPzEzNq
M4XeVUXuF4l6IsOHDW+/lrfCFJCH6u4lMC8Q2/NcE2ITvJiiuEMSAVdksFO8vBmEC9qp2I8Holu3
aamL/6VjH8jwOgHRki5QmGw6aXmFBuGu31jAV1BRhJfOaxqF6vmbn3noL+ljj8CCYoqApATHUaa8
5as5ayGGNMOIh5EmAYFumkLEpeK+mrkrC7RpTBcA/2a80pGo/lfRKtuNLPkT/aMgGZFf6omEAKQO
HvikapyimQqOnMGGYdX1saFjGA2bp2S+6GfY7SYN+ks+7TWFmA5NLw7cmW4TfEJAzfIpYCJtsgxC
6Pwzp9uEouFa7reyoYC+EjKpbcq60KXXhI1Fpd9uWFO6APZxJx9SaM2dKnfk55zktu9dLBVj/lkB
4zq/GFVMG2sY2NXc7St3sB2gSeGd96Wli9jAt3XkTgP0K2rZES6rET0MbPSnehk1EfN4GusYPLVT
2KQmGhXng+J+L2oiRdhyyU3Li+ts74wV1uIxqZWi42alRpfGaXbr8XRvEesbBuRrw5cBKnsxSF50
ndpGWtY2MDz0z+TRkJ0EqYUXQjbe927rj+wXuaDs19VcN+Z7lifpWn0PZK6Ma5ujA0P9VD494eTx
rwdz6rvmVI1VJXjqXDj4dchhtIfdciy8PBZqT+IliKUFU+r1Ozn4HLHN4+fLfpePLVvFcNn/xn7M
7s7qtFTAp8aQvU9TYa3mVxTJ5yYMhiIPdHoqaEhb0MDww8QmJRHeY9mk1BkDuibdhGge9fMqVQ5n
GAHGKE4iOhIF8+A+n7Nf9oT8SjtoqqTZIuqwaJ0lRBQnEfk70a5jI5+X268rDRux4fghIyCz+rKU
372+qFQAjPn8MjBHuY2XyGKU0yk8ElneaGEyXyswCwdEWw4rhqCSep/H63H6SQhPW95XZnwzbEAR
9HGFr5C15/U5kEgzCw3I3O+cW9plArbMdbtS0GybxO8ReOm00RXXV3Lfh48/75+Il7bJmzA1nMdC
E4bzG4J7QH1C9zoWqCsOEiLVuxt5HLdroAbsFJWgDs7GDlC1gBHZpImz05QizYDFv/+pqdKtG+o3
sf+g7NOiahxO643AewTM9Dt10eZtjq7d/uhqCWD/9FN1tGi0NZiY1hyxw/l5TGPFkdYWLO1zV8V9
QTBCEawlNxUEp1ybgsKpugb+4jtcCxgnN2HSHVztkAWeizQENBIWBOzxqDIbOErpG/lhbhlZwMdH
RRYAaEs05bfE7Pqf27sTkHKTMD+2BYxK0pHZ6sPZIq2KiOFqVDcdDO59uM0qvihcpwOtqW4PMs8V
tsY4+LpJLpDjeyOFnOoWE1doOOpLAhROhP4nQfbgn5Zgj/5beOaWZfxEByMYdkHmnKo4bBlmS96u
3+J8IQxClgxzok8Znyjwi6DNqXFAsfwjYSywx96WzBOExtQkZpkKPmE1IG4H/VkSK/mkbd04vm/p
PTRbEe3SR1gxzeYJ3z2ZOmy96P/zvFF7KGj2yYbQsGYNDFep7axOBpCdbyrjD8oWNj4S/a2UOZKu
x1kFMaFEAso87NWcn7JW/eVtLMiH9jhDiKI46UkiVtHcCA1xHIAeEHMxJDXSd1T+JMvKKE0r2uO1
L113ez3WCXpv/qDho12GiPAorLNQ/7aglSELtNPjUOZ+9F0eCo11awHVi6i6JDQdCaeMe2qE9thO
aAeGX31+Xl6yMcguBOlXWeh6Upb+dFPJaMgHZ6w8eMQROX6AUrmWFA87HMmtbj5zzCu3U/oXBwr3
eO0xNMFhp8tH+0tnSSjDuvOzsI/CWmIWICRExnlqw7urZrJmnFtLjuM6N3kfGsfXq1QNR6oBXJw7
OrAFSbNrmvmWB4wkdHeWspdlpihrAiXoYuWpoUSCfNISJBEAZcAkE5XCs+ZXODip4fiRM54SStCG
t6gWMkjZJYE1FSpQAB9PK+Lmpc677Cf8webC7WnNQtApyplXkVkOuoUXu1+A3k6it4rME1eZViG6
dQFuAy8YRsawXKMrZxiYcGzh4hB+8e87sUFBn9Hmyh3aGjefhim45mW17JFLJh0/RsGs66WlSnSm
xQtMNuw/Oiwt9RI8y/ZUv5yVVnnFoc1kfiEaU53/qY64d2U4NxcfF4KjllZQ3bbf8JCxCVa9AtEb
xvxQZkpUojrGkqnCTO5KKKIfgDNWwoS8KELt9rtjm1aPtk5dhHU/jMyJ+ynhcn6h2dniys6CUgOu
VGU/Byw7xz84iMImDJbI/ZQ1RzOytHvQVNHagdd4DM7rjmPLIYm/q+97l6oxf/T4HC0nCAnJjZ+g
wreZ1beZ5aW1rtanpnC0f5mbKYKHzayDxlgqq4jTmF0R+qOztqqxdgeEpijG/DDrC/1ytDazcvyI
1utmMZ5oWiM5h7kbIphtjthvgcFOYyyZVaOrflYq+XMDuXj1gk4i/e7c0JN1sH1L057dHeqtU7Pq
nwUhVtZ/N0SWDRrCrnmnU2JZl2UNFpOX88KG3HrROE+DjpdmFcikK+TDSJA8dY82dSPFBrG0EjoF
SPcbOhGonL7WKJR4xuD+ttCzk4JxFTmegMaKc/DLd6Xei682VCnr36vdNhYvZzftOVqOdsc1SUf9
/mzdgnswi/L8BYxFrqVQJpoltaDVO3XA0UjQf/c7CGaIQjoRrOSQsi7MJ3coq0VxEiH1nzEB7MVb
KTc8xpALv9z4OVFT5EKBOBfsyK9uZ5acMQo5X3+75U2wP2WU6Sn/Dfc8ju8VCb6W7nGnMrzmyO64
PhpKHvDYa9JGp00DkxRFyjenFZOu9+6G3JMgruPNu7xq5zOwrsLgKgim8+SK+ZhgxgK6j854hocE
V8IRZSld64nulTLuPF7eFjByYX2jd2eAeuq0FvCwByp7kkOoAaPPfs98GHIL/esgORMp+z71oN7u
MGQQNuJU69yRZ4/EToCNxKmelTemlCld/5uS26MpK1IKpqyYrISeKBtRGfTzVJ5zeytx41QI6ST/
/7T7ciGk8oeBi4E5T2o2fK0r0DMmMh/XDIiP2mcVByjLiQHz7FRpmjzHlXuVGvYDJPXsseiyUO0d
yY8MQcf2XzM1vVQVkvEu44Cfk+KQ+OanJGsi5xHQtNM2F9H3w5K347mdkAUm7kHOyJa+Rz93bBDc
epy2e7ZX/f6QBdakN9+cHB9oW3FVHm1AoG3FKBF/TWjkWdkp+76uZhgQw8eYa9rOIGCIGO7RKdBR
Tmdw2eQJkelCtwlRbyVuuc8QNYL4Z4Dds+BCQWSbkHRvh2xIZlDoqHNGD7PznjjRNVQG4LyzFH5+
JdVBDJWVGeLwWlAxEhJtkUeqnDHOc4/eRkVWHwwOsnyl9Re0CWSWxmS6HyRIi5sSOeJfwf4z58sp
fyC8hvusRvwwb/1DvN30srAFnaxsIpyJu+boxGTLz9l9SMnwfo1cZ2B3R6AiDRig1F22P57yybqB
zsJ2g0kkCaXLKpDqdnESQDRlfuWJjHJE80hRYPpqqB6HKJGNBHX1OXKdvLIxGooQvddRyuLQWhOJ
hP0PudVe/ndhbHzsJ0Dfq/oaczyqRl+DgdEkf8TaONy69Pds1K2FvJLNLg1SoBCar35vAcRAr8hq
tf+ggGWA3Z3lWtYYUZIp2i3YErcAv8Q54P5h7lsMtmfPimio26eywLNzyEgXLSZ2GiaBRwIa/pJw
2xiBgIrae/qHXXPkpFIijOAPoYoCnwce3BA/5AvDELcQRpdfSfU4hX/Iw3AmH47zsBJp/O8TffGU
JW+nWS7Ak6OUPH90YBcJo78XJpQsRQtRvO2kKkC0c64yc82wm2escAWGkXq0G9CX3p5U1GpNMJdc
UVoyV/jyzl/kg2zuuMKb1ar1WCIts9LpPINBQVk7XA1runOmLbWq0tmK2d7WpCPrEMl9XOwSkgqz
qr7UO/ERvdUkl3iIIId6RSOy6A3ih9FAa95Z3BDoseJa/qNDhW7WCEp+jLyxALDhFEGXp1DNqL99
WWcyl3IE5tQjLva42S0sYYCKauFhxXTyuGTZaGz+ZTqCybcs3WxT+UHx+UXxUy56p93Q8wqk2PvJ
Bpgg5XtHIyEuWve4cc6Jr9vX1bU5fVtNZRvDHXWhBm7uUOabkrPO5bF3W9QJ/izFZ4kNf6Yv62Tv
Z7ARNJz/AiTy25lKnk3B/Iv2dGJV4uQYmNrL/28IlHOnitxg/uDpvrR9ATzsUVjsJhSql0/6NNqK
6N5Yo9G4j4ZcgEZWczl0qgdpDXXXObA7Yu4h/u5Z9Ommu3ajAY6Id4o53V+tXfLdxhQ5Tyk88ZXc
vwB3FojOCyyw42dDLtThkwHkgx0dHrgkNMAyz6VsplqMRkY9bXdchIxmddnu8L88s36IEi2xRKH0
QTF5dhbOJJr11OO8PDahI7o8K7gQEUTrN/tmlfidEkpT2zSUtyzpmrVK/8kamwOBwhVLIIa1PlRN
dIblVfIpUrAbu0/szCYtgSb/y32nhNeEn36nCcD8IvN+y2m8o8C8V1UlYzkBbS140A4L6Q2QY5yX
HFZjm6/Ra+O+gvL36+9X+NOynYd9IVTbVJ6VV4boiZ5ldNPGa0IuVYrSne9D1ruBHFi9a56J6UA3
pG5lUl5VJE27Bvxf1tWh1IsdJ4xDxPLAi9XBwqUED6MtwJeGMXbG0PUlTSFg43le8pJp+7oOCqAf
KA6el6j2slhzZ0sss8gTST0xmw720eJBF0Cv0gWMtPSTu7GgE84HqLV0RQXX89zoAdhznJTJBplk
QBcXzE26JobeY1BfYjIDnoHNFmH7h9sn9VV+RusU8JBA+3fBYQ2xSECI9LzXISEtRnVvnvjZatG2
VnSlzDGSitqEik6dQm0p53ecCUNPfpNcK58gDlU0KtHBCDVrcDHpmrNaWka210wfwnWfuv1KMM8O
BlinL2vbji3FrPVcz0do1JsrYPfSndnNvGoYxjsfKbuAQG/8P0evT/OjH91tIHtmNJPy2PBYTCrF
ldAcWY46r435RO+gzCy6Qr9Gknx4z6GemUYwwo3S2XnNSD74aWJ5hJKYDbtwVKczlQ6/Yd1p1p2S
0ZygHIjkvFNThyPIJ32KLiAzMSONr0cs7EyFLqbFCTQ+FfhIG7Yr9clk5zez8GERLNLEmM6q9hcT
IxZx/YYp//RJea1Ou6dlg6Fm+wNzVlf3tbG47tdkPy+HI8wl/bnuvGvO7dasvZB4ItvsTjEkZFGl
UMilk4GtctDdpSMBdODOfxeQAhvT+FHWokBnyuThl+wX4/koMQWgTCQ7xq8afkJIwTJpM3H00Y8+
s9TGw75EklaxkyF8R7ObAEsoxuiq0u3xMlTPU+jQD9hm5XtEvZdU4ha8fOPCI6kkop1/GxOiB1d9
RE3xiFLduUCCHEOvslvAN+mh/JbJWLG6V0JxNVzrVEHvYKOriWBLu8Em2vtu9JvTB1rqPiNKPBN+
iX5hiFS0RkaooILw3PrnxnMrtamhtunD4LKLayXYwJS1GFKMNyt4a7c2v5nYEK4EtFrnJ8kp5pF2
EN9XmDp5Wj5feJhQnjR8pS/xGTXMnROQOLO9KiPuVoWL70WRB+atyf3Q1YEVJrH3lkgzs8jdDpk2
ZlLdE762FyuRd2AdrwD9uoI8pEtzyt+E0qrzL92XbbuIO4h97q0KsjI9K5FOWTlZP/NFS/0OeTFQ
CUGdZEQenKtB/4b3w8Ak4nQ/zuOFyQd57T62oA3hiDIcTeE3aGk9sk+MkskCUHUsSYUXDh/patFe
u323U7z7i098H2JgQpQqGvjC+60YJTqeu/tEzZobX2WhuRalZjLLjxyEc9vIQsnKLz7bH6AyN74k
Pwl3awqWuxrQMcIHzadLbp4niioXA5qu3/0tfpsKPjcgFK67VM5S2xcOt/Mn9ybGgotdqUkFvUvj
MbaaZKNkqM2Q9qFrAshySuy55HMYfG7PVpYsc0oNMH1xGS+FUOrZfHzaBHcryfcil3wLVrvnysYN
7SyT1cAFnnaag4UPb0NJ7UVowjgAn52pOSXhGSaso8/Sr75L/4R4gSC9j7zCO4L+yKl84FRNXRKo
qdhLWD1HPN6WmfLs4/832UEUv3iqziVrYcRMqdClD18DcaloqkHCk1zbtiKFLzCIxx9jj29Ra+eB
00kaFl1OQVEloroOhSWtAZVtQblhCgdbJMCeV3xqsYolu5mrnCLFDNnNj31Kqhj49x+Tpkheheq5
/gLVpF8Eb3XjA155kZ6SaBb8yuJa0fIXyiM75kmQCgc/KNyKsCUj1E9tlL36x84quSAThuodfxFD
zVbtJRXAUgLsXfo7HTJ18B2Q415oTNCSTVxx2bB8DvQp+TJkRZcZwtAzhlCXvcKV8OK1GlUjsawQ
8II6KeVdA7RoMpDsDBrL8zauZcGdNAxHh97vqiecKEYOj3d8v7OFvG7U0zNV2SuXeKhDqGGQsX3R
ESEyqDUhwI0eluSCvLUIbMsGv99Gk+cosIKorJ51r/YGPZfe3/Sw1bhMu1BFzLwdCX8deL/XflTE
rgcIhhIWm7zc/fqHUo2mNfzsbpHRTnhLHWnmHegMvCrNQNzEd+26Drys9HVDZRNsiMg1VBTdpSWz
4q5OcXE5S2w7w+yl9RZ3N1gopco8SEmpk7sL2+tGpI4kkXFUyQE+Q7IgdUAhSc7pT21lb4aUgjqh
nPeeYyiopEMWW5auJmn/QVbaNTOChAQJOlVHVBBHCZQTOnaykrk85y3So7os1GiLgxUtrDugKRo/
4wKWHx6XUk/U3l8H8HTVJo+rxaUZ8DopmnSy6+qafEs7ZXJ3lDBYl81Ath25etxKieHY+er8HGe0
OTNkCgcDv9xOkQPgZDjvPr0uFYyRV0DMUyuorTdIy2jquhBnSVyONgmrJT8I0XpvYuId+wdXKb8s
3LuzGF/PChYR6odjEduo0nTqLm7GR9uVE+1FGlzeWAk81umAev9Kbzya24AiVqizXoJK9nzlYeK1
UBZK15K1Qh65z39FYdxCW4HP4VA8TdoAdrVqqgfi03+hD+VE71xfoMjcqDFFuZEXbACnry9LUj3T
WiDNQE3QTNRZLjj07atBopHd5vnvV4s7L+RjA5eKJl0DukHpBinR0ka7FiDAFBu6/QZOssZD/KRL
UACagM+FF4tkggtcltdbXr+djHV70wUm9hBe4/2kqF+K3UDo2Xjuk+iWADO160SgvUHEhzqkhauE
2o1wKF4gQKWuGCg08DJkYSxr7L7VUE+Qi+GtJkAkI2cpoc/GU/4wVsIk+lV0ENd0+u3QA882ixmf
ehiuMQK7bYswjn4l92pdLJdxwzmV3awqGD9maQm0y2hqEnMN4a7CJgLYvJtVJAt2yB/mInAC2x4a
0ddIR0vxtK9C5CNnTf88R9V2vpB9J9qsB0KeQ+nrskxshNq7M30ZbicNPgicGZA/nEWR0nGBIbyr
96LB0U8Qjvs7yhGb2s+pri+faMaDJICMf6afIegzNdgs3S/sEozLaNCUKOfUxs/JbMMUzg4apPG0
a3zW0SdPeaxIgjzEhtVayLfUYZ642xOi6wfI17ctcbpE02LtxbaN/6x1mDTebalC4qomtQVg+eDg
EbOVqK9JWh2YDUEof1oF6/koPTocB024R9rLQU7NejmxuBhHOYyfnPfykeXKM0jVhNd0R8T3Ska4
Wbr/7wnAqbpP0eic8+5QBl6O8gblkDl/EcGcW5WhjbSSw31Res/W8bGJiG33uZtNuFv0pBYiyKhK
ZDeGgMrdcWzc/eMDGRhs6SNgaHH10SZ0n1/T5bsnQ7yJ7+VXtrOH4ya2Xo1IHuj3z35AIq1ncULo
cm9WVglGDOssszXg/V0Vl9ks9CNcrJkIccheW/wv/jG3sd8iqTRpFwCO0k9xrhpDqK+0rz8HoS2t
6ry4uKfcnvoViAFVt6/b1NApUX8+rj2KVBsuNWtyaNq76AxNFFY/BsYsG8/nzGaMyLf5J+1f2uSe
ns2RsL9l4VjK94So6qJQUxvFpRLKPV3/wuEjuPWjqLxxdYf5bXMSWmRFc2iDH0+52iMzLpsadY4l
3lwk+J1kbGRCM3/PlNjukjJEUBeZ5E7Yef/ccImBZxVUV/0Cz8VvGs5KxmwnIdazs0FGmwzVX67K
R+P7UyWSvRkzSlETPGsi3OQPmPAg7wwBwHDRKC2KER1zhfwyKPpq9brLedeaKw7AVL2FEYeIBqpp
b8bSku0fsMirwV8ED+VpryKqBvbRqS/iUjvNgo2K4s9RZpxHi8vdJUixFIru3HoxMSEnloM7C3TJ
xqriyjElHNC+drG210rJJhsGUp/anl4tcus/DXqwbZxfhOR01t/9Q5SAseHBxrthW7GMrWeW+P3L
LJzzfTSvA4g1X2NZp0oxuJ2P7y8f57M9nWC4jevHiDb7g3Ade89blZtVFUmwSIrMutfJoUS/cWqq
7tb8eGmjOlF0UZkPJ56evEZd1mOEmZwBdnUF2PhvK19ocGi0jjR28QauZM/R7XzELFDotBG78KbA
dTQr38EJRbNvHuUv0m+UWzoNjZ0SfoL0Ei5S2NPzuphAQF7yXa8axivd6DJrIXpeOnoRW+hO25sV
rubC+zMuftCzhTcwTdO7JF8pIgCzHBwwE5tcUeEeyePlM/HfhjpyxOBVzVIpsa/2LLbp+CatYud9
LQmHnZfVGB80Xxe7Y1dSL4JvbW3XliYNpaF7YuAu8Fzd5w4lFFI7uL/iZt8UX16wiJRFTEni+a3T
32uhPWXBQMj6soMb94fhj2Lff2FVrJa1N5Nxgfl3Iknhf+lzliBUsJJlqtEjBGtAIY2laiNEeJDX
R3Nb1+RLyivu1avTsWbX7d9ydCmg98Y9gileNiSSihn1RU3n0xfs0b0jT1sggjTXAEQ/U9N/JTa6
jc+79f5Lqit+JNicXAbjlbrjU/auqRFfq7GXmzsDggG2EKjZ1SDsGIS2uNGGPmAPq0iOtzC38j63
KcQnnafyiNNdPJu237Zg/OcumbO0gMss+/L/NB5DwYD19Ni6pn4LEJ91754U3vziA/yj5T4zttXh
3shNFVpqb1+RqzRAQICpmjsIe3VnVT9KsQ5Yg7FaISIaY9oV6DTmYzNAXjqltyOBchTk8SWvJhMm
Yuxqo9ou0y5dIj30zGae2adSyT/Eo9Qi8ivhW0pPjr+JY5TifS9nbpcYXCPnnqNRG7hGBZJzkWHF
So/bupkXmFav1xk3vhM+PcHsVn0NESHNiKrRWgt2ZSY6uz5xEv7OMkVvcQhH/XRjRdwrX6C5BGx6
ldrq63ixv+IZxRqZN1ZpLlUdf0s2dun7sw95o7DivZJVZeOeLUa8ZmquXKTdZGZzaalvkveZeBQg
9O38NuMoTCPm1Vffb2zrfJkODd7iV0haa4wsryxRyy4eW9+HkJZnHxLTcFiKnmvkstJoEPXkQkXn
1pdUr/ZNF8txLVqM8r+4Cv6V2snU9YnzmnSrCQHNWyOQsSxvz1Ir1nnGkLfhEvCV3IkuzhpnSWJi
+dukNqjiM2D2J6IzwmAR5AG36FfR3GHYHnGLq/bMBBMXz9fQ+Pva9e3pMVBvXt7pNu+FUh7iQTvT
ABQWxHIyDZOEpt9P60JZY9/bShGrLnzft//ih832YGj1Yb/g7JoxzckaQTK4TeCZJIlYolWoGXD8
wcM4AnniagyXMOlYEktMqCm+8XA1W7S6cMRV92+C2Kawjqi3UvaV7iAklIf91Ojd/uis+ZKiLI9f
As4fvAr1bn7HJAwy//accOqAy2RQGJYoxdQOxWChqRIQGrVHIRxjOFgGGDkwZfGx/3SiDeBLh+1f
o3uNlIdsFXsPwxVEdgX7GjnxMspjBSOPBTPDnYpwwtaKu0e6+bIlek4mNDFV5B44ru8ZMhDri8TQ
Q76POWWL1dZumM0AngcsZ0y3gnkuuPNY+Iwru8JAqKviRf7+PSEMXICb1TXaEWVqBzxShci3VrZt
Lbm41driag20MpWJ9beVCzIk7EVYg9Jd4mEKU2hsUsHdnoUUtk4c8h+63Q2cWc/ZnFEgmB05O7K3
Pw08lcd2AoekuCjJo+bxSscSNv++9NNHCfjd0ELfietW7NhkNWCzyx8KI02bJH/aS/L7khAT1HgD
aSFWIRvmMr82XXho+qnRGOlmyllOphgBqWKRqU94bpSOjiH8cBG7dh2aIxxXP+AzPxZpYgfhYe0d
cOORnSijJ6fIl0PFoHlLosn6daPhzxupSoN4CfG5q1D+K733GKuQF7m5CEznoiXzZtEjuR3cGSA4
K0Bv9F5YRO0fMObKcvdrgz7i4QldHawlSOEZ/ACubSHrDgQA4ZeTDFkXz7r+1j0ud6KxOsSiJUpt
so5wlX7EoU+Aa6M05j9TJ6wcB0QW9Sp1Z2tt0zEh7yNCNjbiChwWf8vUyi2EMpBZrnn5SgCXIYHu
uxRRTDf/BQFMwYbyrS8QXZj9AcQlYDgFevzjtqBNjfFVm5RygLspmiGfPKqDKJChIB4+d7Tdm2BD
CwWd/7kRNwnTq00Igk7fUvAIKZNFkgJzsv3Z8Q/9iIM9AXhqkmJ0n1Ysb7+p1lhc86RqPVOH+d+D
2qkQrk5q5YxMEmsGPaDcEl/BjqoeWZjdaOxeegqRp22+SE9AEwMGHL6i1WZEhAP8FCCtMq/e2Eyd
vSrMxUXrIKLy55Nq2ew6mh4miJ5E85EzhD7NfCsJOvVNamEceF4lgx+9dPx7ouSI377axNvCNRZi
BCWhnyq2Pl2+tNovM6PRNrrtvuxNz8svFGO/M+ibzhLTTwAiBbriUHblmTZyzVd6hAVeomaUm0do
O+utDJe5QOcOQb2En+akTBO6972laMIpdhG9Wg7iPIL27gZIjc4QfRzreZyhGqeHUmJfFBXewX6s
KC4rYORbSKyhB+eyx0TKsZzICn4T2NyvqRseY4f/LPFeyL+2tdCSqnP1ceQJOQY4zMxyaxhP7ILD
Dh2ZFB24GyKLRnV1/kIHc0UxgMoyJSRc+Ot4tqvaa2uxBrRxhz8LuZCG+Gd2oaFEYY15NnOUNJe8
4pyVmZBSNk4jaQs/5voG0rpPQ9ssLTpcbG0mjPWo+2dkl74hD3i/7VbrUktynrtd6avjXwjb9cJe
kR6IJpfuN5VP0ckVla+Goz3lr7LoN674USbeADUhq6wD/IB4QhunQO7xV6cGX2LIMrr0rPn1LCBU
UQjwnVu9NkK/tG3pHwHSu74ltYb2Rt1YIuk35XfRm4U2IG0CmZjk+4fGKrkiybs+0Adje2Q3wWCi
1fkWeqR2OFxvqPhahNryjycTAA9CLZ7jSiRo9Lo2fGFQO39mZYys+4xOHg7zTHq1ss3bbgGbtlYf
A90TTMAJ/tPIByo+ZGufudvan+t8N/txSKlUlGHEy+5uvY2HawrqsOaoUCgbQxrD0oEENYKEZZW/
UTBs5SjjGFU+v20AI10ZiJ9H8BotGuIRyTRIArBROkcwGjL3u1P0adCU1ZDeZ/TNmr4mV9ls7KkW
wAAJ5ciOlqkdCsi+taZfpVR/5C+B2IGznHa62+wVTk9KOHDjY8QB0paYXK6KjddXRfvBvFGNeem3
bnTcYPsyu4fQcoYUCZ1B9D2XgIaFpaHVfuirELpQaF32k9Ibe7g3BFGCgtNSNkiFZYSyPJXI8gdy
baCFFl6+WjN+T/W+SI6JG+H9ySaIUieAmEAQ92G036DJad9q+RRxnHj0FaTO5umIiTjyJuO6VEqH
XZxTlQuTMdJ6an9zdgwmT/Rxltqay8mvLauVWy/6aAb7HoIcswT9xHqxQHkJ24UIC6lTQpz2fqlp
ataO0Kb9ayV9crixQ59IffQQcIHricg0nb/GZaDTYwhBGlAhxywWs4ES9vI2nwtB7yQtWyHEdJ9e
jUEF8JOdtdv9MuRxohuIIpcnbzw479egMxeAa4kBbroAeu/ShrOOCv0guhXKJ1poW96u5VEqPESQ
Wg9PPqgsmva+Yg9McArMkJVxsJhwFY+mSV6ARUpQLZnQjJIBTELP81nlI+boPeLMXrthp1iG+LIT
1lB0MnAlK9dUMHfstoqoHOGdM+jGxguqV1pJXYB+qmwEJmX0aQvrYVTYdjK64pn7QI9+fyqsSgo0
QSf4vR509v4OVlB8IsrLLR/dGHeT4C7G5T98ytkzWLMiGFjwRoOUjs7MBonuL1wnjyacf17lbvCg
s+rNBnhP/lPz5GStmsHrD5zFUQcwyfrbYCUgRJrXLeOfvePl+xcbbBuwqge4N0ZD5vIhvSeCuhpW
FicBIN8Q7gpPYlaVptcHYRlpkmlDY4dstNZZ4vCGcObSuqq6VDO8e6ICkMzIcSWeA0LyYl69NCsG
PxxJ1OfR0sUd9ZyxmnMyNdSVhvBULk8550VtLohv8z+sB1P5kvFWXw4t2Y/ZRvnAS1uB8hzvAAbw
z/pACj6sehvRTphdA4rMTTzwMtXHNSnp44/TXogTzWlZB/KHqh3s3Oiyhs4/g/qrxZsUY4ep4i2o
5MjXIwEUAcUA09aihlV2RgLSO+/Jig6LCKffO835vd8igyw11xMwvMFkuCgioGhjRR1zOeTCEQGI
C3JF0fWY7T0k4+iFiLPEVYayPM0DRWrfoEAQDy7SKnZ94D81lPosiV2xm2XDtYiAgThh+xvESb0E
g05tB9TWXM4LaPWOt/x8TretFpzpO5Lma9u9vfCZ7ylrLTAcT+KRuHhWYwwfiHdZRLGH74oPRPbC
5YZpTfvEs3pyp247tqx4LL2d0j131e3/LDcHFjJ6GEfDbbc/DKvOD9Ii6K37tZ05UmYyaT2JKgL0
dviBsNqxDSXJxLP2DGvpXyLbi9LFfiBIilA4negPh0ZbtlJwZjF2Dc9UvA+Mucc8rPhzUsJ5Bgf9
H9bQ2BrHcn4slJXvJUuc0/DuoWUIJQ9uZ0Yxy3FurKDBUr9w+ElFU1Hh2s4UJwa803JRuTdw5gCw
vcHlor8VdG/7LNh84TlK1er5hw83mY/oHEZFP+WSzZBDAXvuKkx4pjdLijZxi0S30HeJskd2aOyz
KRGl8C+H6JZeErYWepH4/2qKid2tKNxKMHmcQWlSmI+yW0qCHp79U6ci7tsyVM9Daf+4MLk6FXz8
AGKsuwo8xcladrlEvrKz4gsShLdndXZzlgIAs+mwmZUccNqK2X+O1Aw1t4c+YvbygmjMlm4nqEE2
NC0Es4YLeXfRSADvdNY5Emz1JYCvSaAOR6m4XCxnhWra0wP0o7dabIqcPV7NYScpfYoxUih+Oc5B
NShFOwFO4Rp04++Aaf9IDDculdGhhwy8DTI24JEE+U+11JAyW+lwoGyeN1gc83BFfe7/EnF9QD84
ES7d51o1oV5MAwBFMkZCpNX/oKJgmTPkZMhyWtU7uc9vLYuqq5kWFhRhk3cbTVqgbdZrTAlK1/g1
WjtXuV9nvnfH2cb+nYTFIeVmR0GupB9QX676nACXNdoyjpMCnTT8OhrYMxmU+O5g5439s6wYqwT6
AaNBmgNaVdsX4ZH2sjAPvJrOxBTMMJYyGkPvFFgfRSbfuOPZ22LpXOZ8nuyfjbt84H/nAM4W5gs+
8CKm5aKSUdGm0riXpX8NoJr6JxETRtHGTUsavl2tbVB6407OeuXfNt3tc/rYOGjn5D0jEpM+0XuM
lEj4mbaJqKIp+Xiu6AzHSXaACQCOBFPoqCdIK/BPJ1wNOV0pNtQ5VmtudALjSqV+GboHhfgdnZ3U
3iFnMm25h0qrY/STO7bGr7qIe1GLtFJAOGqaLgMKW0Wycuk/Ti8rX36oB8PNS4BsQaI0NZPhD8X7
6xM5QX0XgyiS+fj1PtWByrA4kG3FNhROqA1S3myFeT3VSpXLbBnnTcsfLIHlvXsogZmJ22pEDQDi
L0dR0szxM+Ep/T02XdJiqAo9CO2eWAOBZGfHlelb/Q22IbYHxg90W/IsEjAotBbt2gnmMNiVwWma
7cM3vXSHuN/NC7AHdcFv922u8ruMwH9Hu3+RBR0J1HrkFcfYvRUjXN936B+Tnty76ZZtbR1nGIoS
EuMyaqszboF+IuQUq1MeQyVjuBIOcwybEJjp/L8cVmbbBPjxu3hF7ol6+/VnYwR9TPlqZOx5EGOC
tdzMOo04JOOfuDHdLIAH0fhH3GkjyP2v/vuao9GozmMzTYUqZYdbDJ2Kpt4/b66LyzE4rHDDfTrW
1xSl0zitorMZI+puyAdI1jLA4IcdanehVrYhp9e4BoLz0Zwa1IHVtCf+C2IOtDIOoB1dK/NkW3mD
eTzFGbFPEyC5ZvP/O1mHbE5erTor9mUTzpWOolfLkYksks1FhC/Q+esrYKOEO7Z/i8e5E2mfqfu6
GssklCjqfIw27ojJH8H8Y+mahsMMZb33PUTdB9Lo/t/08o6YwG4VXqWBZbgnkUQ9lhu6aXHC0bRj
s05cjHF1wv//9MfBN5USn2DE25XNtUwcHvS08QB3gpp9EETUNXkjguinUysWmMuDwI4qX/HOUmMF
C0Ju14BUHRiNhYkq3Q97saLZLtMFgEN5kYllxsiSuVpYHkuf0xTo/RKCQP7LDkKRX5GKMqxVpYvS
XFwLpjd5sqi0YXq7+lPRpbsET24xL3ALH3jSzy8q+9USjtLpDYb0fu/SPWSOFn9ufpVMD4yQfxzG
66gKk43BTeuvuQiPDJ5/4Ga5+zwtazJQhl/9vxt4fu5/wSJNalVudWry39hvmsqTKCkXoOC1JwMJ
ergxN0jgjywieqKHFa8Llr0SE9l+p5ybDlDfzzXQOpfzZ8wqJzvjNVtNpN3O+ISrQHSjXof4UfqI
wo8qq5K9B4rq0X1wxhQ4L9ClGxqy5qjFsYtQN2UBIM5QeLu9NYk3qyDOx+6Yf4gz7Z0rXrcIQ6Tt
4WKwXJLm1dvd0D6lMDo/ADcM8qY1jeWLe4ju55I9jgxGX9goJJkamYg0tsm6cHWxU1iHEhD7VU2l
bsoJkYW9mMK+JD1eaJIzRKObwwW9Jqu2U/13vWLvJCSKsKYxnsea4YRN6jNFK1DtxQh7z2ROmu0N
PqLbKIPGwCYXhDFz1TV18/8Tk6JuBUZzEYkwsWEXg4xd+lqnuDCfzOVOmnd6J0HSKfkuoIgjwkJ9
ZtoCGztRrnJgVSPfv+vOCnO1RYguXrCBHtugddmskn0vocYB0tBxJ3fwlZG+LEjdo5WY3VwnIvlV
yQUmhQ4Nu3aaapRCvA02o0ma2iZsjAvGVPtxk9rUsXKz0K67P+udgUbNIoHNEYqF/5aVRrtQZGWV
y5yWRdncUGIyWp91NEhDIxWQy1k+n3F0RZHRppdyeUYfVd/0avJcm3Qcr3fD+zZDw+kPQrogPEzP
0x5MTBk3ztjBT1B1mC8uU8QWamtnpGkK3v8MIigZOZDOpJDz3Q+fm5LGmD4Fnnw/Rhf3PB1AjH6Z
FOTYHHRwZHcKvqOpw8LR3Qnp8yzzfcALTgC4VhUqUmDsTHX/lfmB8E9M3aJqYJ1vMmxRfxY0YY0U
9R7IwLf55uFaCZ5k6lqIoLAxeXV5rZ4i+91VvHnrSBj49fa1Grsa3VH8qJJezJhvTi53lrzo4Xki
tf0O+MI2nE6ShdDlY0UdZEfEqJvlVTbTtEVyR/Fk/5AZbi11IaWZpms5z2ZzbvfsHlmC62z5aiOO
vOhGAx6ByZ+3K04evXZ+t71m/d5bIn1+4qw1VQPDKmmeJvFySYFw8S5Uj+o9c7AreOXwfLfYpErY
uI9xRbGFr1qAL7rZjpL0zeOeA+Ei+Zx2cVMfEznPdGVq6gvFdlym0Hv+88Is66LenfQW4xla/lg5
gDJcFA1TZJQD40nJdWSnt4c8Tu9nzwZAH7U/nodBsCjn0DhC+Of8lkryUF6NkZ+jFrwHqpeyqnsv
0sPUnwSB0ko6SCbIMEQ28hm2fWJEkL6NfXhyp7sO10pEfzAcxN8DenwslLh9vKocr6glQJWqwM0J
W4gVPeYMFe7t4ihrlnt+hAfbn6qzVNJ/w4qAjSWtykK7EZn+9sg7Y2bKLkZYBuWBXOztpeXGkr99
oe+9PQc5Q97K2WLxRv7gPkqBlBk6trtd1pvz5FQ2xr1+SXcXw7JV3mQays95CraVPwLR6uV2H3Rp
HJd9JoQele1Pp3TXRwhiruFQL9Kmw++guLPKg6WMb758LoXXZslPnEShQoF06JquIlfjiqDExXwj
Cj0F3dE9uUtgGRz9xBQ+1198rowJvugUW4J7mkO6ql0oo43pi6czj4dsQEZfHpYFkc7QWMpcgEl+
rQasnDP6kcaRZ+sTw75zM4jfxf6Uu57XM3r53z96zk4/zkTyJRrZ23lH8opNw9gZtYQQ1fRoTXL6
Q3aDKx7b8taFNR0u7MSS8BDBgPvXQbDFWunfLXbCVHQg+ga5rkbldB2MrWKVOtl4NDlmaNh+Z2EQ
hMRLzIQ3Ttep6+O8dbozZ6OrnmUItFFhhgiwgzPkc+33DdBv96aZHgSYP6rdJ4ivc0DOni5THT56
++2/5v1oMfimlzgoS1c+jh2HCeY4hBg9DSwvS1i6ZW+6vM+RcoaUmDyT4awEodCS0Ys1sn8GwzZN
80xTJqwpn/Tbdw8ZI0i6KMeHtEhG6NwFc2l9fazFi7sbN3IwcGvdzAfdD2aAq6uvQvXB+sSA/KHm
0eOZwzN07SNTuqgYR5l8J3LB0hJaiZUpJB2q06Lfh75m7PaN0n6iZgq1mpem464s+v6TTKGpUj+B
Q6L8aJ1y7HWm9JONMZ2VSl0fuNM6K4/70tS6SRahHbVTBT/jh37oDgSNySiI2OMc0ou/chQU3SAC
p+E1jlU26f1tJNOcsfVQTPAn7F2eQZd5bhX8TsnXNKol3nW/XhGALKTNNgPdkgDLSfBEsiY64L/p
m7T+P/KIgtCGOxr+aIKGYUOLsHOxkK9qIysF8KytltxBufhL0szCdyNurZ8q3ORCCQ/4//N2sG1h
6XdzvxrJM+XInhp0pybJMTLTIylZTH6x3qi0vZ4LJ2FMdPZI6624UO3j8XmlCLtH55iHjtuYITgK
brhaPTBDstIYIoxaXaGiyFGJGdAJU67YvpQuOVcf9Pj2tbGF8tCNaKvOmY60wAlsahQX70bLx4uP
FUFrrjpRBN4U2dBeWqsnwBoVfKhxrL2va5AspcZQOh2kuW0tp4Gtznk6awlHX91FTsRgloFkZO3N
pCQ4O5+y+psR7/7C60qz8ogdAqbqyDLX9m4Xq8CoLkN0Rh5AsM/b5E9YhezpVudrtJEsmE7UDtDt
xUWCZ7SAsw8+L8Y9hv0G+oRA+wOKHun9R2eQCjnQr6rcMV9Q0kD8zPiPHR4t/siGIwiY6qCFX3gV
kiJBgKP/OQgug+ISVE7SEWq4kQ6MHs6dUbPbSvWzHIaoO72x/75/uhKhCO+R/POOx7Tsa97BsOcq
fsKDlb2ybbFQBCunAphykAcLyYX6guB8V8rEKyingvG6pFGSxCciVJvjwlxlFufUbzLm6bkbuSP2
QT9tzcTwF7tswGrwCNq7pqKXV4eHCBupUHzKqrs4CbHl1ZJAU2sKjX5A8goDubZStVv6/N/U+V5X
MBValsSd5yxeiwa/BoG+bj5b9XOaRg594dp+pt6g3oND6LP+qc33P6jo3/9xwr4kS7mTR5mWwo/+
rpY7EjFkt3E0sYpOmzXjQeVL0bZ/SYVR0LobDCETmKJx1Bx1RswR/kONA9BFfO/XxdKh40nCfQai
DWTMIq9rSBQsoXk6pi1U2BJZeXK/DMEdwwY2pjBw95kVQuZ2G50TS92plXSVdrfF4qsY75SOVtP9
VrHUmR4aXtk4MsnHtwS+p++VvNm5HdddkF8kz+TbqD3R7wIfyQlpqa7/vxSIcQlZYJxdhPwmP3+N
ZQfZI2kgCk1j6VRP25snjqpVaTHT40edKz9fViGvBJejOwBCoL1lDmpp8Hwpv/Bj4eLi21jc8+Yk
lChEaqmUP0sXfSdX3lwuFfu31kxAMwTuvfMiV0vIJ3ewgu8N/Z2S2V/QmdO4ZsejKBlHtMcDIK2K
2pHy1qPMLkW0kPfxktrug0KwstHYMm422Ord/WrgXpkB1svSSrqoFJpBNnjbUS4PzHJ73AVVB8zA
X5k7Gh20oOgyE411jBhznyV3Ac55n0OGrGSrM+N/G1jCPdwNqTmCZ/mDeFlth6pq7UagTfa/gFxV
QlwfyzFnJ9dFIAEvGk0WA8xHmDDNXqNSE9F5jF0Id7HGHGY5dyZp5WsM3ugt24otgiQXOp8iFXvs
RKT6gGEuPVXRlAHBzLOqfth/WZXl0kUojYAvHUciBHR0URg5BQ5hujMDBWgMDdLiQWnFyGWhrne1
euftfoDAbneWFmoA38yHDMnbIMszL9B6oKPGS11V1gpUlqKF7kadqh1CJQqaKgxW/dxwcPeAROQF
otKP25Bnml/GajQ5jfUTt1Cf06epyO5eoZbkmINZrKDE29IekfCcM65we2LP5B3sbUoX5tXeDvuc
lRzpuxOv8E9R9QIX7QGaF0w/UFNPKTKczc/Jv7vvl1FniFFXtvu5YpOpVjT4wGp3T65eJ/oDFxY4
dHR5H5ZU6LRpBL/9dAeLmT3FUiyM+BWqdfuArsHVtxreikOH07rjWBYWG6lRfvP6grshpwYJ9uwE
NP2NoqCu2hgzi3JYKkh2QfRt5b/Sgb+KEf46gRe2oAFPozJPhp05CGL4DbqQ9K58munOVgqKbY7o
oyB4rosry5IsJcSeYYyfsFqZvy9s993zH8frxihb9it1VfUVRYm1R2EsbMLXX0tn5UU745p44AXd
QEwutbo4J7RXJ5s7+vNu2HKiRXlg1f+CfrcRjzcSI1hBSBhgbtfBc4ShAiWRP2kTBpK67Ft3QEcC
N+XQ/B1RFqJqd8A4Bts2qo7s3lR9Nz4qIv7El9WqbDf41qC3rHkhvT9dGsaW71vL+Rip/+A09jZJ
A9tQkHCU9oA1ISQ0UxDVhcVBeZYcQU6B5pGf1EXOCVSgsBLxvBZYZ0XpYeqW5CN0uNm2Xra2qi/a
U5Fq1PmZGG9Ii/wDldJkaGGXquqbduIflp1eFKZYMRCZUvR8YaJICzt7LJEfDpX1HNr2d4pAbRTL
sUAsA4y4KWCXz8M+tHv0lAS5frD1OibiGNM6yvtKcRvLiJTq3vQ/FuXx+IOdDlJZLfZZFgbHSl3+
gJe6g4LUrAi+R8WMRdiD73xtR/mVpYuBzJ70FuUi4yqI6604c4wRxmfkz8GaThd3NA1UC7sPu0bH
ykfKsgn4BXSdh9mLcKQkGUd+LEmcz2J0mCFLWpaiDF+ic3spA4+Dr7YkczLSxgINXEIymrRK9Hrh
9AoGsjNQNCGU5Muu3zgaBy1C+Ky2dvYsybJEtoFfOk/ZZvF0CwUU7dTftFY235yog2XgvUoCCxK/
Tt3oGA7OH7qZ3e4THIhbvqBl5YTDob+V1MDesd99LedBCq4O6VGEt8Sr67B/NBSz3vraHrCrrGDB
2D4LBzz8r/ETxL55iyfPbiKgIcWBl/oPMwYCJSaRWGw0frAqbF5nOWVBr9KKL+STWd0OI6ukDu1r
9IU9mm0LYMX2EbqHkAdVdZb1ziD3ZCO1GkzWael184KTpAx7w3exEL83302e3riV5Ey/7HKVEwQc
V51M4Ow8jcriYCpuOnWDbCgsTw8gok76W8xSgroeTyAPKyeawtrwpY6JGgrLisvUTtjHY2aV+L0t
OOMJT1nsvtifQfsp+UkNiReywv2Zbdjdj/YKq2tpViTZ9pHoelXNPA2juDpVD42y/SCCCy3VMnyk
DsAk2WyAm3O1DUf9CLF7pLoZLMh9Ex5haHGAI4p0JLSrysWleFl40gTqHH6MVORTrAA2DTuZsdFY
cqBt9+Dpi96WkVb/yZ3pI0SPuwKL+OUa+bnJB2RVPBJhKLxKdF7z9XOSXqKsd8wPCrkxIBZzha71
ep5UDppZSlAr32F/gTnNFTp0U2FJb0veLJ3+4hcIF/MwcvuveUDIuS2kaLkqHj3iLSm/q3hZzOEm
hW4qeWXKrmP9S1qRLFtARarhWL4Xn7oPzZCXyq0v6BQ4SfrXIj5vhW+5LQBHwoRqEfbpaH0knWvk
btxbs/se2eCGGjLj/CSL1LosRVKG4GVPgKorMY0DKHLrVJAWZ4x+rrwwlJX+5de2U5sRqDIB8ba3
lz34Mrnt+7N85Jr/aJ6qS4MGickrd3bdXui7C3w5bqk/uGDz4ETpLIZ3tvuQbwX+rN5jQ1uLA7Q8
lP7YQ+obs0imo/hqy0XhtpAc49UuCMIZrZVKGI6HJDF9ttNCjWgZKsVKrvsPNf4tMK9RqWlUvWPh
3f0Cza0PBCSnr4I3ysPbavnaD8GLiLCesV8yQOYbqsrX+/WxasdzhsXoBlXrD8jLVenRC8Nzdhjh
l5Omsm34sjzTonulDToLI5MUlN2/cVy9l9X3xObE8BmesqUtoUQbpITJtR4lD5+j3wNaxqF/zjqa
hph8ASmaY18krjIRmJ9Ptf4J9nioVF2m1zseoo8RuU/iAV8JKC8OBRk6TjJpLNs6lmK5bc+GTM6P
d2n9V7ULjO+XTzDp60FGMLzuzrLeejjR0rIfRI/nNWifcMQm0cA8wRO+FBaUs1E2/whkKSUMl8BR
usy6XHm/iz6COKwyfPitGI24srJ0mvXKmN1lm01Kxpl7ksi7PHeSi3/jHDmFJugEx7UAJn4xNFDC
GDwCU7I1ULLNDFE8b72g6kTZIt25jZwog0j3JR5gQLigdI+ZCPisRxbL+r1+DzooOUUW83vfiW4K
qReYjxtQRF6q75boQwIc0edrlg8sZb6LScNsBRYJIHhN5cVG+fyx3EZnaArUmR6MCeFQYrFp4Pz5
I967+y797jTYdO+uLH39ZXopvT1eSbeoQ61L1/o2ez4FfLKYqLp1jj08LGcC3uziDfJ7dcD9FKP1
2UE0JrSab61IMa9BFsBmJaHnzaNTYWs=
`protect end_protected
