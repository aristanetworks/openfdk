--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
gBai8vC8HrtIXuYyQxMmLMxe48ZEekBcYltIzDVlm4rAPuBs+mBfV5CI7A2Bn7I5awJvGJUNYR3l
/HcGm4YebouDPPfMlQj9IEHYHkj+lNisBbKt+Ozx9DOOFB0/rVmj/pOollQWBH8iEfzZWemd0CuY
UahFcrkoCpuBbYgzIt1SP09vP2qZB+3h6pxSfgJswJh3Yu49PX5PGbtX21IoKdgusyJ7QfQBuZcD
Mx9noOsvKsYXL7HjfvbGLgel14Ogm8CpB9ueJkoSd5/PFx4nVU3vaVlLeLZLBksrh+boVWA0JpB4
07R50EXhkYnbdxVShfapVf9EJeQQsJWe91OIiw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="W3aAYtjvMpZ/ZbEwHLdpCi1pNQngyrsg0UgvG+bn4gM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
pPtBuh5eqZQbIkCGz++eKXKG0sHaCFZBVOYpMxTfFTxRwRztWRn+fBiIPExgvQeTOKLK/OMBn4VR
Al7QDcEVB431MW91lDJCSzxioOkts7q9PqxeeLs5VZ4es3QRqZte0bLrqxyfcTYT4d8hPYPuEkBk
8wjzTdEtOhcpcvAr1ryrWjeMVwyRgIAuNOUo4q355p2ow2RucgGv3LpD/J3EEko0i09dfHnXtiUW
4947CaHwFpuJqT5PhcwclnB85JVjEMdcgk1M5rZk8KQcF74SwQhS9Y8VKKh+T0evHP4063h15bmi
RSS0MkTHM5YZgjvK+PHH55SxMPTexRGM2sjO+Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="j41APodU4y2a43myqsDefATofZGsJqjmRo3k5lTZtjQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2576)
`protect data_block
cZMjR2BNUNTXHKtdosSvs+s3muCtkcUI0/GXwo+EsowqWGUT9n5qj110lRUThc1AQVOVvt7Htz7G
GvyoaGuHPVHczC2Nl5iG/8pKHB5zFVDojHvVy+2ha3leLxqEPJicXAW6OvwEDVQQG8yXmtGo4raf
SGM+tLxix1sXM5f9Gko0XAJX5XpId5wN+uJxbxTQsaPxz4d4QF+VOlwTKbMk5cXk/eLqjC8xdltB
5JNIkGJhs/1amqeaLGSFKQWpynDVt5KFO9DIW0sWaEV9TNfQVIproLV3g3MPddg124p2U8dLLq1j
kxW67Jg6nSoRUeJuexXlppnImnX/1B0aDytgqkV6Zb1ka3s2NNbrRr0goCY/87+RdAj5EW6UZpGK
Un/TtObOQPjgdKFvYq2Y135TQklaoG/4wTe9OkQO2LNEV6EkY3ppeCDl/4RCKy94jlHH9RF5hAD5
fbTWZ4NglodpSMg5fEVjJW0N+IntOB8B3bPO5Dh1RiHnFGAAxjT5Jn61wD2HkjEDi1AogjISqb4T
v5oeG45dWqbxoDd1UGVBFRaG0fK0XAM4N/RV2gILjqqkP6C79RXeYoun1h1VM07OTGIMhb5vuVQk
URma18xtAPysiKgaR5yUe6fIXjeZ4D5M4zsJAbvCzfC0SEyBEjusJNn9O57McJ+wtk7gd1sYHCuh
XK1Ahd9jsASyqELeOsp4qm1vqz0BtT4/h2Qs/rB5YfmJ389qsYd7uvoZmV9r/jMqskJqGZdJ9KW0
FdNffnHq4iG4DY2kS6I0RyzNJRyV5BkADQsqi6IM5xldPEPod0bP6JSou5yhiRQVq7xLv3ulHl/u
b0G6U53BUCg+4j9rAFg4/pmcVxyqnfBRYihCRjKH3MwaxrFbVNqxqizeRuHAwogFubbnEEiLHL81
pnk8LzjBJ5PbjJciz/og0a79n8ncf+i9cXKwD0jnaatUG2uLlmAl9cGU2L8ohBrOfNIbe7oUmBWQ
FxCzqdH4w7yYwWTvE3ohtS8UxVj/1SYU9UKLPAFrs4TYzlfo+mqD8z80xrrxFLc9ArteIO5OWWvO
eHE3awy+0VmQUgaUaw9utkZBVUgycdT/F98cGMAE5J6KEjNL8Gjr1oAc1uI0QtZcpAW3/XIt3AuT
JkP97N5x6ftbdsoy77BsoDJxGaW82/Kr+rkUXbXYho4vy7KSvdU1SuNclNzR4VvLBm20+Lr1ANt3
iEUSPG6lFXgg2xDx/cm/cdHeo9CZaLgoXEWErdKdqN4zQ9w+RfHEo1MYB6mVav96e/zWE56HDQBM
Syqa9HG0CtIGcMQvQMnjWi3/Db7u5xoMKwLIBFN8jnHU+c7jy3LH7TZIP2gg1F3KlTXukO1ErI/7
9kEOWiW9agN+ruOvEfOx1VZPl0IPCqlVTBb5KTNR8cJAdI8ZtJvLMXedKRLGfReO3lvEaUNZvgfR
dJ559Zzf++oJTWiVGSPmbCRO9XA1FM5tfsW5xFXsClJig0vkMIkTvdjmwPD9bV+V7k1JwcW73p24
sD25sQ0EW4so5DxQQHJINOylCCFzJ8mdmRd9dqq6kusox1p6X9z/+0QjjK94E+gOGd8Ejz3Wdwxl
Cm7KD0wqB4VDSKbOLbiVEOCm1YIp9vhA5PX8YpDDmNyY7HzYACwbHZ2AwNh77jqchGofCcLKhlTP
gwTvBKdxhtUQCWy26U+v1VAkv3BplBn1ECsJ3klhFIfkVbn0LcPeqckn/dKmG5Cr9Ah8Isza6XYE
2+VV9m8vcjoaOdkMeiF9RjygapCZUa+DUUcUgV7D3kUHpviul/gSmvP5QIrjdmWZNGDJsjPtj7lX
AshmPUK18jCuxEbWmUGo8IaQrIwOFPHXsJBo7U8sEqd7GfC/h4/XCBGJqTDfbFM0HTLVUbRgdxss
Si56ZzF+bowa5SQypFa7QMFFjhvYxms8YCnflzH8m5nDWRkTWTePChoS7qWsYL8Px/4x2jMicwzq
BTTxbqMu9I+TM0WOoXiKWrDyvJUWdziTjpb9dRsckfPwcUgQb22TgEFkvwgnz04uRFJwQMG80O2k
qIOw+bZD3+kpi2VmVu0OYSHND/f9pDg0dh5DitolX3qIoy1jJ4MUWTDkMw7cl/TIGY9ovg1zz7Ci
oxnEIzCbjXHseNHaIn3pZSq0pgM5OjS/zkE3QXfi2TyKxicJ6pSZZ5dUWnC2TCyve4/NO+7wE+nB
ZeLvppsej8zqbBBsSUOBdOxTsim7SEhM10WeOasmoxKhl5VcFTjvDH/KTk21zOvhjfHXVJoS6w2r
LoovWI+D9d/bzo4uI0G3Pc0C+jf/3gigj2Q/1ci3GVuzrTbOhIhg3YSTm9wMSy4TStKhXYARQOYk
EpUX1bCnSdhm7qHJXZjK00U1y6FLBjhGMEvx4kEtfGTWDMRGDpO48edIZqvrIwuuekuLsFz+jOAV
uPXL8xzfuwmucNLrTahp/M7za5yjaX5/irO0lHTsyw92oDIjqpI0eAySCISmPd4oHqvfrhb0rxGm
0e7xrHjpnHwGeDj9qe9DFwac6iOREc4/+UWPBXsbND1OUVlVC9hSwjUO1TWJZuFtL0KFNwCIuFvW
O6XcFiDbVtwSXJQs/ImDT/iQpXEGx5CDiAbrCANIhx6tw/MgrA6gX7PTIqn3W1/XKfbTzXJxAVfy
zpwUVZMxiIoFboBBhOmANL3W8WeGXTXvnu8ONbtSNtAKOu8hM8Dfmgi4z4ZgZ42ap8g7Ax7yZiqf
AxEZFYfpg88laeDjzKm0sZux41J6+5nxVQBSEwDTfY8Z0kZLVpGdDUBkkQwj2x0oOURcl83fwEur
Mqh8zvjLr/Pjka9KoYki8YM2YYyG+CB74MV4UnpXOB67BPji67i9hbgbLg7cxIzOi/0/r4z3Qh9+
XD6ZY/x4Q9pvYjT32uy8QdfZXyvZcjvg4eXLbBw/jOHvHfFylLa0Jhm5u8d9TJ3bUYz32oLGYThA
6gVeGh+pzF7XA8OSHUgfwL0pxgYGO4/YdSxjaSkFgsrGYl3D0RJiG3ZMsjgPv3wIRVQ7Nhq8uM0w
yT2SJ35z2VmoURklNMlLkfjqJdy+hpGSKtXhWf8E8McarSKkSiEaBVK924rHgM8Xt97ujeV31xXk
qwTNomKD9UDLBe3fFrU6iNAGGkqI5oy6B91MGLlj/wohQvZTK3+/w0AxHVIke1sQbbRFvQr1yMhL
FDNewZD2SsI5BGhoKI/Wz2/j/Ljr0YJcgUm4v9326VXwxvJQTGDMPlNS7Nk+PHU4P6HIQJOvpjXg
cyGrMn1/7trhcd6jzck3fGW288TptUTMUNR7ETkSs4cCBLVslUnZB+xbw6gvQ6kNkdXM5bl6gyya
/w1cRqbDHGzFHaCd/vbNrra2oCtRi5Vdcf8GwBvV5l+NwwYvQ6/tVstU+KpSTgZkIbPPvhZwIzLA
uWidpnidhKKGJvI=
`protect end_protected
