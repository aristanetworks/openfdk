--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
NXP1ttHo/zb3r55CEkbNKHLlxy2Raqqhu7nhnJfPSt70KuVOx1b0SV/PRoGddvcp0Z6VWRkiCTyF
dxeIhB78cNAPH+IFfVLoitBs5eITTkYyqjmmciMXLnZ+mvyc2grOR6U/KA4Om4qyzZ7ePVeWvPf8
PPiXJMhdVqx4jWL+SVTZTATPD4oAXKEs1AJ/86WTQGNvCGqugaqGYhA63j+tlnOGgljifp9urZtm
ZULLRnJCFcoEwLiSASNtNeYXNPLp8ON44rb5oSKOCIm41kKtOh9GjwYaquGDfReDzEBmxrbkSI3k
sRfrZ4ZjRu67sgkYQuCJ5gSTYy0CZWJvY7CIgQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="NA4pkvkFpYePaBjxrPq8EaD7iN4cN6GCxePossoVKbo="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
GhIfaJjgiHzwgQyhHTDY9tznSWWQPdwuoPV0yVgTNN6Z8MX97oa5HVCsGlalShV4Z7QCcQK32I1D
LcQhaY35zhiwHYyQFkG2FlPxHsF/iEX18PPc3YmA+S5+cNMHXAj/nXg5lPIS3RcGz+KS4ztW8Rv1
GhYjGLEDNYil8O+qb8ot71qf62Hobx8guVtM3L9FEWtPlt442P9Y/MlCUjjdAKLgkP5nIl5mBOne
Ol+ogxo7392LON04wry6m8cpKGU3kVNATeevRiF+wVTK1n7m2qrH7cf9rO76ks+RGrXKfnQNmHJE
O2r41IWkaPs4cC9xIO/1IehlAxHNAnqQy0rFqA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="h58cm5Ta9snVDj+fqeN9CNvKwd441GGyVU/o21FVVDo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4672)
`protect data_block
SbH5a9HBjgT2ZuCdbO4Rm/XjqRYxwRRnmaTEctqV3FSLpog+NwntzkGHSzMg0y2WEjRgXF2CorIE
vKmeKyezD/e/8yn/lzIDtVBUn7NM2j19brVfTzIzG6OvTzl+mOKUEC5CqlcChsK8cmJ2+pJ3Be25
xgY3+6W9zK+VDq3iWpaI1jvQmNRHkli69AqR9C7qw2cXWp/5FmABTcSDqa/u+cY/2cb7mXpKKSxE
7c7cX3WTZgEo/faWW09Ev0o1PMNwEmC3YlsZwRv60Nl4GyuFNz19RZdo6SIKzd27XLFZgtdzZF0n
cnnilAJreOwNtxdcHMj7a7a6tQtmjqkSQL2NHJ0IWknqjtaQOIM9Ul39fp16HruoQbfBOAcnHzk4
puAIXUB7K4dzRHDDFOQKqWlZzgk0jB83yo/dN1ikqT4+NOYKe8MBLlhF7USw6z8nfww2Rn2nDKOt
aN+jNpcaJ2+r75dIDhScVe8hKhilLFOyUyA6ZSCaWy5YjfMpUibrfAW138OOb9VNMUbyVfCYq12w
3xBzub8mC2HT7MNhVeEID80LNqImf2Rll9Uel1I+KtFL3CQaLmucTgmpKgqof3Wbh+RqCi6qTHEl
hbusXYa7jUWQv7os0PR7ko+zphbsWFwlAudJd37zSS2t4ytRhG4RYPzLhgAA4i3nsCfYbgngHdSv
+9o2fTVLsmtmogo3bEC+ZzAKG6hPZgirlXZOOU9GajtZtK5Ul3+vAqcXqyJgtQj6M78IZXZOKHlH
jSpkdJU5BIN0NdZmrnLrj2qULYpxIB6h36fGJAo2WdqudFbTdGU0qIzMkEVrjYt8cioiCYzf1MXv
QHGj8nNZYtm/vVDGtppQunJ0Q/HWUa/HC+AOyAqOdjhSu3jxmBrF9nxP70WP+k3ZAUnEQ2JLLexy
4vhKFvWS0c1T1Gkdj8kzaclXg05Fo3ss9bUcpbhR4YrBxxqJQAv15YcCzxY25fnra2GaOrIKrnmM
hw88ZISLgzc0Ll5jGLO+Y7H+n+fo19Td9vqGpLurUdymMmHsH9lYN8rKADg1GAd4bmf5NvErNqLs
nSfhwQFi2B2BZsNWSxsIj7tOV7xYK4kO01ieA8tVb6xaWluytJBgFu4nSHtZkLvBK1+wREA3QZLQ
U60ER65PJ84xqWrNRbAvrNYQRa23jIbMpeFLcd4nQXlm0TM1iTGvpWa607u6GfgzQW+bBWnP/oUG
4LIVtw1cqQnVZrP1tJ+BwREtNjPSgXrAu9qTWbJcaMIDOjSXHCAmSfmjU+6AFueYec5HjR6f2w1e
dYFZ1mk9bcGnzHIjJf6V6G7X9+kfFZZRCDMzrPqajCB8b00WqdfbxIPUBEf3ctRdRB3US1Ya4CVh
VFptaMoZjUxV3sL9hdYo2ZoqkfWaxQEoWCJ4fH2dqU6zIKdoJjOff5xFga4yd7Lh8oISUJ9338bH
zdfo96VKVc2KJ2lc6O32ygn/YCzlHsOmOZ09fT/q4+ibimpwhNoSDx1nUMltVgw79q+umxe7MGRR
Qs4xqmGe+Zrzpb07OEt5lqZA/ghSUUduGTlXLqd6Yun4dofqz7XpyqWuskKQcTbVCahDxKnqtwxM
bH01FjjhC5ARRhRxU1fot80ugotfu+ndjPiz0p3i0BmaH+Cv02DRbBrnuAkngQ/yb9CKgXI+v8CA
aU3QeUU8o9EC4SwI3hIOBp2C/BXu3zQq+f8bH92zmnVKiZ0tintGL1mqvdGQ6WiVel3bL052TRGI
OSZJdIlhdcsluR9VnwYGL5ly8Sl/9Mz59lfOGxwtEbeRnAC+3A/2cDHwKwPnPg8Q5buoKsgZJBDe
EAkwM+cfnww3yMtpj78ECuoER/a2RZ74aHJfQh3MaORKSSJXPlpvPFXFeLtztGE80U7NQclFKt/q
irNB9vXdMcw+K5RnzCpBDeqgBAF7gEDfkMrJot14YbQS7wj7AQNcI6fMLn3vcIVYuxnEfVNLZbJL
O8nwJUDpcdUJBqiWXsNl1o1CQ7W8IEPQ1kfto0oL90ESutGiScG2JdRBg+f0CwSUSd3QPyxi2tVV
E53WSRiG4kZtGSGIgL1t5JEI3fgOOqegMZ6gFGIeT4rfsMo2PkPZ1ZWIwZyTrlrZPiUqI4xp/7QJ
g+EQ4itLig2rvbTDYSTCt5qKFgl0mqqkQlQRBsOEP9QgzyOsoytbg24Kge97R5N6JY11A6Uy8/Oo
R1txxJ+0Sj9E+Vk8Jwo98THvT+wSvl5aSOcPubbi++L7aPaObBWcLnjdRKdbvGylx6AlCSnpOPMp
6O5iMAOQlMoNfZWkkGINgDrtaB6je7/6+OMJ8J1jCKW3IuUD2Z6ERJ22Gn1NhKUJY+hMgeDn7SM7
LUAZyoJ2ZkOsLA112GnjJsWuQd4dFaqKpSEsVQnFSYKnopxk2/Q17ieR8LU12lxu1UGUtSEpd+TT
r9QtmDJdVNnZEU+pAmp+fBZKFdFBPBTxdNtPsuzFa6OkJCMUEYav1FeP58I3KV+oynOFaFPmgBI8
Zd0yvefczlH0drhGPjCidgtvgFCuqL8WZP7ABZ0RWwQNVY4imHTmY8xqA/U4xbGi46rm6MwtPiqi
lvBHFDvl2QHw7xLYzoXFCadl4cHyAdNuJ2X5JVHtTwG61PvL5p9iIxSb5Pr8ZLPPrFuX1sn5QWIe
oExGSZi0gSbOiQtfrG42LPTkK9WJ2B4yUqWVq9eBgzTt49WvV7wf3B49/k95dqU7uhM3EUwOv/0M
zUis80zqn2+3gUiVSjNHftWrQSsTwCvFNzA2OpApeWvr9ksSr3ii/sre9AEu7qcHf9jnWujNsNGy
3fgyh3J5P00ajVjGFkKEudWErqCefktZMLCTI1UE0WKpJmeOq63HvoQ6RO5BMT2hXhkH+rmqCBC/
l9oQn7Qnj/Z9yUGsTBkG4dRo7Xbo+P6eUnCidcv7dGRpz1Pq7eRV5eKp/z5UMznhkl0mzF5cQzQq
zS0wnzoZpigMBMzToIMrmI+Vg8syRNYbY28ZHxM5iY9gFEKQjUQG9actPr4lqUJlNwvTC7ut80Bh
2tlwUtPm9s1kX8Z1Fys9miayeFYaY2GzpSTEoD0+f+AO6ZGTRuejgxDUxq2RoAfzKnvLTrhFTNmj
9GLuEC+9UHumqXzKlX0Ij5F0GLU2CvJolLMYqAobNMmSEjKDDW4pYc7WkQarKI4Tf8aEJ5k1sqdu
+xUTDiujrQt00QIoT/IZARIlPRJzQ7SdeqXhqht3cQj1itjwGKdFTxX3OXICCIA6Q1lpz2oWAZqk
I/jStb6ucCWaZHaj3EFaJFMc0VhU9hYSiLyMZn4ybMi/8iCrYY5JnHx2UM6XdazjBmIeSbV3wZBg
OM4ypKppAaGx6YMYygNVHEHPTxsLfmANY2CCK7PxU4W4AB4rnC9wOxcgyWVQmijHkTb4MBRK/Aru
ZafFmiRSkwd0UNkdGtfdrYILVnONRoIyG4WdKOFoFqGH7MH9mzsVO+M9QltiY1sVEtp5fLtMO2FB
b3BeLbE8tsSt5gIxIoG3fTszS70yMQgimnn9xVNDNke0JDkCv8iQz+4wvAIuYlcAmBbZsAuF8Ax8
Wk1GuU8+88UpbOcqbMq3WGD55TKj7fV3zwzvDB4kx89GTeJG02nvz2OPxzIZTk9DWY7wXssFkn+f
Fj5zHjbIPGvPPKj1fTHOMkuVGqUnQSI/eRnN3XT8r0fXeiof1fzVLohC1vy1LyPdYY5oYT5QqTbr
+B2Cs414pLIBH4VLGeGt7I7Iv0hJsVEi6XbqS40/hiN0QjXgelgF4jGMNoWWxvt51D2tDLR9mYz9
vIdfXip3paScwFgq3Mm6z+b24YEzMDmgx2iE61gZtFzfBHJD7pF3ErtCK0ov6neEqGNqv5g4cC2r
asP/hdKV7myF3PW4fZIc//519X0CyxyhmV47NNCYi9E4L3yJNie1+q5oZ/ivtGHitLdQRW1G6ERu
+NCs26QnAF3j5DEWBarESAY8JboXndN31IY9h0ulKdMRjR2zvpebXWTEZJ3wzCe9C4JORVbQ7S9f
B8+x9bkXRbmNO98kbQbebVEnaTS42cEQz7t4wULPFcR7Z5v8QD7LiyTl5E3RXyiXXeFykZnkvJfP
Ttxsbry/huhYjGtbNWSvTSwPlaeTz+lwaZwjA0jxyxrw7Sgb9FwRtxAN9tZXD5abpb5x4n2qzsvq
Vb4AxKbhNeKouTtt4sQbQM/W+hx2tDeJ+z+RpSWqM8bZTsNeNtC7gOKbx//UHV0LOFMVTxYrJjYe
/I7KlUW/BW5E4n0qivp2FfGSWyZDSgp3PbFCM+v1aYLbgOYjtWoNqH8Aoq+TwSGF7QsXjRMkxVd4
nWlLNmWLtQZYVN0/rZmi/T0jswS/UCVXAISp6Vr791iCrP43nwH2yQyoNTzWVHJFmj2uLphI1uCU
ZgR1Xx+k14G6SAprTgCkelHbiWR4T3GSK7Gxr5dyq8jVuJvE4InbGLhoHaEJaHeXT/KjRq2LZ+uu
+UD79DfYZuzgTPFclCVq5stOndY5b5a6LvDSpMWD9qW5zmqZxXDEiByt0v3yh4Hgv8J5AcYd+luv
qcpBXQzF3HBxQJ7Wo4Davx7/jEjiVv/81GA8Y4CMFJ1Z7AKk3C8Zoxzm9GC/6Xo/ynGaTDIeN2qQ
2kF5Mtu/SDEOkD9fX86n7QWWggsWgBN4bS9fosd5X3Pg+4I5O8iIxNqmsdHjrExXexwjwhu0bXC2
v3xIGDtP0KPBFJ3NRSwFR4Y8hXCghXC0hwxdrGtIxLCklmagptC+8ThOIdAta8D7f7+mG3K7BIE8
0xKgrQJNYrHSx2K6m+15Qa5Z96z9MLoMYxbe8qR4WHesZQ2G01pru6+yPug8k3Nyu73Ht/vffRTT
WGdzQTUagpEOmk35pF7Yih6pLxmv+qzLiT4f0SSzcht+/r7YuDB/WXRCJsfO4+l9glkS/2nifb2G
Og6FAOD6hxYFHofmdB9NvZ3wZ+aD7WzVJ/MYKvXeFU3gMJOcXah0ZzazuFFZpqZ907in2sQtGdNt
6bxGHoC5+cXcvYv/+2b/dMMm0ynAtrx2aXFcmVNMNrmUfv2lFeEovjZdY30AOktLxakYWYx6cqQ4
/TCGPJDHKI7OM7DLc5D1jqqUBx38TVg2eF6dYSHKSPy7E2yMxz8Q6FejW3R8zWAo5IINaJCkCAGP
kAgNOMVxUVHz3tICsPRCCTm8eLXIofMJM4MG8N9VNoqKZ58LDs03d+urAB8zcNYQYWnTbxYrM7T+
/+S9r/do34S4Yz7TB6i3anskvCQniaGCkAJXKBj87Up3bSPSXsN6+7U0rQYq9+41Wora8a4qyKel
KZCdoiL/dFEzZ44ULSPL/dkjWw5LAn28K/dOl8EEJFpwai4orNLNPbmuh/QKSZTLb8sr0+wmJWN6
B/mhNg6PZrPGMMYx8/u84+kTakReT7TZ5+avobO+1g3+zgQbWWiiMlCz/UOvr0QV3eWNi3zxTGWo
3UgrQRrxPVUl/tBrKg198worw+i0X/wgKJfEbmZK3tJgQHoUc0j/xSCs9omcFmOhn5Pnug+9GYez
LuhdEY0Ldcr+fZbnI7lMN8lNNG75HTKo68EKhpLSGo2nBS/mii2zLg0RBGwbRIxA4o2AvY2qhNV9
FpC2fT+SL6E3TsAB0MweG4l7QK6JJfmlg2SW1MnGPF/jmIheC7QF8nAADAT0sn2xs3kzv6k+rHRy
s5vsEXQHAiJbZq6OL2vi6Ci3J96Aq9ILj+4miG81yNGWSNeRdpBBeV1k+HgZGIWtPdyGiRM2n2sS
8miVzgHqRGfGvylLC1VLPYrkg5nQpkfjwiPlKKkPsVupJ9yjxZdBE3vin15L/MbsW6w5Nctd20sJ
Rbm1dpSY4695dq15UJjeGX+AwPjpk5uI2Udc6XOl1VG1hQ085KkepRDkeI1twuUKJxwTuTfdrYyP
h6qTD1H4IU5cfRYyQQ1NyCEc7JTm4VE12AE1ki8FiM6btqkRNYt74ey5e0T9CYGCQ8pQ21F8OQOa
jmO2A8ridN2Jvck4PGUMFzUlDNQLVCI/3tvVIILwM9P0NG16JNUmMukeoakYlcHxYjCoy+9nhf79
BR/mdPMjh5KmIiMWqla2ooi6cJSx8p/ACTVoEAJ+nvw2RyCaNUXxfBQC8x/kB8mWVLPYTjLcZKBB
/31NCh8R1AsqUqAQ12lwOQO6a4ljFHOIRY2UlWjl8wJw8XiddCD6fFFwOtdj/IApeTXjXVtD4g==
`protect end_protected
