--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
WZANZks2fph5b+aro4tRDYY7o51ZiZAr3Z5p1uyeyAzIjJ/AN2/ynMldHpgIaTGtFZT+UjC+9kDn
1IhSisujPkdJPjMVkgVU1UdLaIbyrrBvMz+cIuoAtf2yYoJ26Elg702zZ8GCE4G0BYMeNp2ZjmGm
iGqJsB7GD2z8AsXV3ZGAxo+mntgN6cJG9tpUWJ7NrSqGHaIYgEv9yFe6zL/LvNKW4lyIFvGWt05h
yUHNLlu76nc+uwoZJPUmI5OvtKNQEpYRgaDtRYwAZ1lJg1duTO7zptn+kiYlMr7aXX9/twMoDsc9
RvNsco0xTeNIg9Q5DMZhp66SrmGJ8f9zm9OcJg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="LNLnZqeM0juLITZlYeO7B58TYxqBq4lPaDKSflWA4bA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
FUGX/dEMBLY7GEhzdpPAA9SU4CJ9LNftQjWanRn0cNf/9deCxBlv7KhcG4zXHR8NTQxj84ksNAL1
WvfR78tTx7ls5iFZlNrBjkZLKxmp5CT7LcOTqR/H0dEKBhB4CF48joiIe+B/YR/q9Bvyl+nf73cF
8dS/7oqGCA70JhR7EnpqaTawW9pK02YDlhZwYpuvZIMjGK2VDZ/n83lv3fVe7NBapkDeEe2/jy0T
8naQLkV00oVpcwqvZMk43+1VkW8Bb0h6xpvpvrpCA1tL4n8ZQ7hQEwYbg77b8zlvprcl99MmuYau
ytzBeZ1J+jERmW301YctVpnH38Clig51PnMBMw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="noWe/wG9SIrK/mLtX18Tt0L8eKYWepc1q4I8Wx8OgkA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5616)
`protect data_block
RpXBv0a1806P/suiJLsQ/jfM02/qzHe4tfA7snMBfP/wLSRkIu+Z4x/H41hxKCv5p52EZlQg7BSa
pl1/3046M0sDBmzRO/9x5jqSuZY/PH6w9J/2RMJi0axTCJKttu/0Q/+S5TYWw+72wCxnx0tMYoUJ
Spk0VzjUhDctGZag0uH6ckKla8LBumoFs6AJOax2NDlRyjmUZvQUO5U3DV7sHAm1Gzc8wsYE2821
tIOopdDV3BG4lGEidov3MWBDcYqLJx65fmg0aFpPbTXz7vKbH/YqgT5fCRrZtopMsvLPhhXpXKjG
p6Z5fdjHynn9LLYG2JipR7DEaws5yj44nJtJeGFfWgnsTUW0OySUBiVl/cLghXpeZBVlohmyA3yC
9uaGWZG2qMSvlcIyvJUKpuZYcbIarvEFbObqsyXU4EZTOzgaFv5ZhYk3YBN6NE8EZAS6Sdhuh8p9
DtP/iDqYb0EeSmqGz5blQm0J7s8nzvBypkdL0Vai+UdU6mCvXfp9bghT8RgKzz3sELhE8DcH1Yjv
uKyRODV+0gpNL2zNVK1SgAzhZn9Uyow1Ny0dc+rcAC6ZEHN7YIsWypQub+xb0/84nGTR3t+d24pR
WfNxfJDXukx4iTgxrj3TcbJrOrDQBq4mSPASBhkEetrZqsdWB6B2wwkouglb1cU4G1UJgKUZmgYo
lTzNCShC8n1de0vEo7nzryQv3uTK5vSzVvp7UqUTZN5KVz3H4rwGhsrO25gm9Tb9QM86NDu4hIeV
Ing3kwxQNrkFWXJrXiD1H6B+4qifNi30tEoRjGYbr0TIJbTOlOuI8fttgUouH83yr9+s9I/fIDFk
d78amhOZ/EQ78r0UO+GcGSlB0frm3JgHgfHQuqASEuJoI6VwjqmRVpbtI1K2eDAyZL3QHK3kSQcT
+zdoS0guXN3wA8CtDWc6hdZdiV0eu0El25XhWsTuaN1llcb5Jec2vyjmYL3be3oIIdlojtqIPzD+
qrzwzP940fRu4XImoCHlOJTK8w2Jng0Gz/vEWz8ZnCNc7iIj6jPKaQ+x+dme5PRCdfZFYhzrcaWP
JHAev8/19Js8SZ9qC0gHt1Pn3cn8a00DC3/qCh8u81GZR7nK5THh/LGDemcP41FqA26MbrZWZ5TW
ZJ2Ulr849VUaNC3xWNhc8vixHotn49tu6Sb0jV1Yz1VOkKEqdAYn9H1DasqnoyzJIrAw2qTco1Sr
NxmnJ7eU4DOuARWPt+9VNXmlUCJDtWiacnhhmCE9fseDl9ucm+KkQA/H7+fcbnX7zERuPWKV7t3G
F9pCI76apf04w+c9msdmi0tzKWewu3GtsTwVQCta8U+oDx6K2f5R/WCsvpD3Y3frabbmW6QMNTaJ
vXNwefqmONFV8e9cYCIDC9kV8YgIARz+iJcc0hg2W5V1FWZj9NzAuWOcYoE8ySLRQoAOCCYGsB7s
v8pbPcx0lC+UGpWFZ9kO0Iv3FNKOz60+uIF3tvLm8JmN2LTgLHHma/fuDSVRNoaxCifzfb9kRY/u
4kTWPNB14Qs4oB1W8tM3lDYG6qInp/Yk9SL3O6mLEWTkhp5v98XxIg8avT9SYzybd/TLsaIPGM25
j/jonTy8zbSMY8okUGJ2YRBj5NDD0eziSFKplB/otHDe93CQ8rp67QP2dc6Cm+0oEsgIqYSEPWL6
Up6lKjYFj2eaS6NKD4k6lSuzqixh2GZiSap9p3BIjanvKN49lwKB9hZM8P3q8dUEiMRaY39ZgTOA
8p4STFZJ4otT9CBtaMT59o1gV3SBnBZj51RcVOgj4Vbuwl/hQS1qHDPsOfNoHDkB2ebyGbwzWRNl
lDMsMgcHjgmEVXgyU0gIq9a4kNsHQxj9oht/pWqYTmdUbvor6107R7f55OY4jC6/a15Yh//z/a6S
iuavp3poRMLTye5zLszA8MAS45EBdJ/t8E9k6JBPFPZAN8rK+dOgzgRflEihk5NVGM0QuTYY4TyT
UiisOgsM4Dcyjn345vmThoU8bN1QGq8hAl2huPFiUrDFxApH47IpPiADb4LevbLNCoGtYgZsBfkT
InWE6+8ZpVnwSDKt/2bwKr5c9R4rtDeTZ16bTevcEefAmDNFeLSsk0bjND3z2IeXADRywflsYZPf
aLEKOjM2a8g1sThlcEH4B3A7S2SMjfWhpn3Q4SuKLHLr0J5CBAGBP8v9R9axXvvEgiVv4+k3blN/
KZu2lI/O4K7Ob56E53v4nNZsEW5ZTOtbQOwtjVueMJ6kbz1kFNvx8PQSdffuKhJkEcejOG/jN4ul
JL5bBMM6Cl4jG25FP0VwoK+QsbTaIkOy+AWViowG/W4pqlYCD7ikIMhQf/CJcXrd5aeZBHxNeF52
MhJEfazPbATOnjem/F3RfvYRzSPrHKS1C8NPEaIMZtHmXK56cMbdBAYbbjhv8s0EGvp+Ipu5SZ3V
mqaOFtaHWb7tPTbYi+hOV90VcPb8frzf5mCi+QwB3RAQXS3xJxq0WGHu+iNxJUfLHHPX/y+sVYyZ
5FLHRwgPpDS8+b4cPTBQay5d69YBxw5BC/8xVR6lh/+f1XpmaH1wodi0DeH8KrQZaa1daflX07Mm
0W/Oc8Dtwp+U0935x7C6sB+zfu+81mVRyU9Wa+OcTffaLt+fHVF/QBJJ+ObECbzNM0xFtMGht0M1
IYt+V6dfKcYOCfCJaWdfjdFue9zzWxMFNb7xTp4cQxpq6An+fkzaFNjhxzBkG2nipYouaOh6zWta
ldoy0+tuhrBBlMs6J4lZgggwciZYb2/u5YjDzbT0j02swre9VzUFcYAZ80qInjVDvOIuenaAZwzb
uE7IzPF5Hw3iqRDrCzriMcr50B3PgcMo75WvucYvisaiDbiwZCoUkXbdxsvPfhsCVibmoTveaD46
ju0yrLqyrtIjqjKU6bqfAn/zHCMwK2zciRbnZ3T7ViOjl6m0A5Wm6lSlZIvFl40rtDohEH3VFUIt
z5ztUcrPoAcLooD0p+ZQWNHaSM1AS/WamzWH57At4xsVBW3ZToSNLuURe62FYurfyVebgyVwM5ly
AaOBnizMpwkfGna4pOmkH09zYPd8AvZKjR8UkhTDOrf9VbOCa3X3Ql+G+v1+QQldmYC0nnNBcwFU
1+eI77waVZIvLz4sZVMvZsPC2N2bPZ1hCWAUsk1B7ZFSNhfptNnogfUnltt1GmADsZxMSWFobRPH
XpwknbPBxMoz0IkhYlyjxmYLfJGIVaoCzazh8/Mm5MQPVeiEkieKwStYbwZieV7mmyQwasoE5eB+
iwkL+02S35c1zLVx7YrMsKYKhcGuxgscGy+leBV8bDgJIuO09UmE0BN9sTM2SvpSm9WlVa6rE1zA
Hsa+pst56XYoW7NTPneKsZFE84jRnwfgw2pwExCFw1SaLqGGaliHuqJOc32YmedJTpssjmpxuzcS
RlyHLrOUOflW20R6VCy/Mc/I/+jyWcNJ7MmRji5gj+B+h/8xlKuqEkmNCn0SYWqZ6LNKjnod8XMO
Bse45CiEoZLgJQDVZSCFSGyysfglwy79hAF+rOxFAld0VbQHo+C+lATN3JUA8ie3JZo5/aL/sCdE
8f52r4XRf3R5eFJiPhVvSOtdWbkszCQtLs+JaUXLte8uDToDYisKBLR6L8pwnHzJyPPEzQrYTNph
gxwuHnzKMCEBXXUG141YADVtq0t1YIEM9onnbZ+t/KleFiLQUWlHsRhM6/uDvebDlrADsRvNXcFs
QI7TB1vRhiYjKTdLSySFQAecNhAsFvjKXE+PL0xkZYILguIP2xfeoVx4F3/NRBe2e93HhF08Az+l
tEcODMNrk1hASCRk+c9uwOHqZoIyY4NnXZZMPYJ4pa3SmDBRAicFKu5tKA1FhV3B8Cn7czwT3Zse
oqX3rmFy4DG/i5L9XN0KbwShlG/c0p+0RZkmOrFp5INxkzFKxFiHaqNj4J3zPaQoAsbHhk3o9xSb
2Rcj0K/Qk2j7tIYfv8x4n4+Pdw7L3uYzs+SJXl+2w3aCbI8vDt6Cnh68dEERIdi2DkKVYubldvYR
aO7CW9aiiBEV14uXVDIc7RGB/atSORrypY1mYTzu4H7drv+7bx+vCCcATDHPEw8l4kruf+fByIAf
JebpQNnM2lmaDDaB5sUx9jJsXbUVrwwtatLROMXpyr9+ijthyVmqpCgBq9FHbytYMsd+0c6WDMTt
kfjZa/lvAvcZzkHmF349ffk7+NO6BwjLcpkkkYOr/cXmWny7Eir2pkZJkFS90uM75n10w5y5QaJd
nvNfYR+gJ6NOKaTW+JCjnI7mJ51Yq5oD0D0nLC8pp22JqPoE5WsMPc2Ka7JwN8fpzhFn1YC/H7Bo
5Cf5LDOmD2+4BmOa0iADEuDQc2ONKfNThjmfuyyfG3RGNQ/jC9+3E7R8DQbTT5+Am7kD4MznxEYM
hLZxstyNfEGbGRhDTUdQqrHqNmze6xlEbpezg3szhXY2/Bil4No1/8jLy0nF/P5/sEMea9in9xI7
dHvRDADt4YWaAgbWiMviRmrn4kuFqttLtpeYNeOp99e2+Y4h1ODBbD13bOp8Xo6K69YBc0baLEZT
EEFLGjh2YbyMmS8a+186ok2ZfwJVJ88UObpD8BYDWF8Pjx8a4Z4NYV6T0d/Bl/d/Lbnj3CDpbgpc
77zDWjlVh3xTRr3ATf+VqVQrnqmwta6wbu5X74tDCQeT/OHD5tnIVSusc3qSW7nMo82bJWgSRFAs
9BCvNzaO6SdDJh7XB4mscjAxJVoj7qhofd9O9Ut4aegKpi5bs6Dw7NDKg3Id/+l5WbUL12fQHB0S
XFP7Nx8SgdS1ftkpoT5ul78nWRSFW8JKtuMVkrlabzfp1F4jpgb6J8UV6A0JLnF1w0S8QLdPjtZm
+TWkyJNIb5piwaCwWlGvJnHAuu42/tLewasE90oDIjJjHxmgUaxy6kAXJmDX4xibvJoZZrVE9FSQ
oVZMls3AklAzUTrlkmktR3eTD2D+m9Saj9ygcnjUH0no6fppjYOPKjCYSzI9HG+D1syOlunaO99A
TsuU+1c75Ut2zmewLXaA7Ml3BRYqW95rXlEsbKNg6/nOrkppUFSeAx1OiIUY/5+Rs5gcZ74efagt
n/BRnNF/JCIRjrROHwRdRrZBqHcCpMJSuZ/rAZiYzQ4S392kZzFMzmGDYoYj+IeOiaCgahLxRnf7
2J8Cl7sNYZroq0D89s/1bY6S8wtdACyxURpu7t2GFAaZU2bzehBvEf6U/qLYjz4sneZY/nnDOvCv
s8DgVle7QfvtEvcoTe1Cxt3ZbOSu/IuO4Q77jR0ayyuFfOiXihV4fZ97NiP93kSp/8wOFTt7lYpn
N7YZTqQX7JBTY//C5unGpkO+4TcoJ6QSx2AWNX1eVqcxkh+4NF6KsUyhyZRSoHSvF0lUn4a2XO/k
8ZmY5R3XNz44Sso81rsOjZgaTWUJgzmE/GA0EELykc9elvJo1MUVE/Bbv0xrX6ZMhgBtcY4H9K5B
/Ftmw7jC4+jA9jNRXUl1lVwea323XkeQ8ca+2pIvydWUhd2YpJR8IDDG4Yeqpiau2CGlnNdzKGve
Ja5RKABDkiVarzrY+IkZno55p03MqW25a2yldZiVY5pz5EkyXd1ctlelBCAWJ9ZxpeEtR6MqG5XN
kPhumo4J9i9fZS5zl4cfwATwc7xU5SapUzIun5C18WntKj5uaebvDtMSlehEhk+qQQjhTWuvzore
fD4kfCvG6/BUoGt28m0lSAvS1V5pYHXDsyeT3jsxFaK9zlQRhfvJcyAdS2F3bCYK5PSQLALvQu4H
H+GOMmqM5W/uLz1nCnqCrqX3BwLUBdncf8xigah5LwtObDd7PNnXRDsgprhuaMTThNVqkOTqux4g
7F5z89fTdDUDloNi42dl8z2Uj4vWalTJTbHbAN53Rt6hteJJbbzirSpwM1myRRubVlsKZrdVgTyO
vGaRX7MhkKUSAZ92xufO9wBJM5FjtrQfW9m42YdFpd91g7BXk43YcQshjw4PCCSYJKbxH/P9OH+D
FzayafOF7LpqB/P0SilFMFxWmWoMiqShF1FPOQ0AZRz7SdItnXkvMiQuG1K9zpWHfNK4K5ZMOlOO
7atY7tHHcYAugsB9H61AVm/60w3pS67ACkuaVmwEK2tyAtCgsKXikrR5786VwVn6mD4wm+MvQQ9B
pIUvis9UcJvFPZ94MTjSJO34ENOt2fqa4PwjpulPTcX9olC9wpzrxf/h9VxMA2W2+wAvqw+ntaBa
HCcgjs6oh4wVY0oWJQyhCURe7l/zXM5kUnc9H+CYtx4fvIgwDhO7OYKoRHOLXWDYi/gsA7xql4dh
kF+Ufmu5kR1TyfxLx8wuUp/pkIBGPWkw2iSlTfUjmpyNRFrh6tK4frYnWDXPp7G7wvrpXdIGeZbM
FwRkPwSdxxLkUT9tHY7hU/edP6HSeO1FOe9lFmieUIZwh98DYC4OFGDbMQ7UEgksyGezYt1G71fX
4mN+5IGHnQKed3l75kFjBwkaDmxaKdUq6v2sMmEscyFTfOWiZqnoWq9YQy2frdOzEeqeVt7Z/TTi
Jl4VNeEz0kX53jt3Ug2oXz+FgjJvglOP66ruRTRHyvu/lF63xdhbkT6HNO9t7nY1QhKCSTALMhyF
muMZr1Zc558mLJ/ZprcbCSBPzpPMQwI9iQuXyR7GX32CstoWbollQVDUjBni7NAC7r/ESr4irJx9
EKK27lLyNyXjxPns2xIrbinvC85LQE31H7lYRGu27I1/EuSEDihPRL+DWCiGLPpizk9od5rOYX4a
g50DKvIee0FYS27u1JxeTBHTTlgQgADpsqPt019nYbL7Q+jCs5UtBTCKDcZfYMmGoMWptLtwIKCz
2h1/07CiV2bznZzYu0q/OGH/m5CEoVRAMTR/CTJvbaL2gPhDs/rkh98QPo+ksh41n/Tjkk0Wyplr
2YfrAOJ2z+s9GvDOkaUNyAiOqao6E8kkySo0x8uDTOVSifvpsqouBXGi9E6F6rbjbMAhw+BgxlCE
6ycKTnuTjPTeolq0iqkjQUSm6LHRx4b2JTHPAWuztvgw8T53D/NcJOreGWXslAhbTrkKZRWcR+2i
aqtE99rCe7ZlgJuZWgLLs87KlldlFk/6kA6fMm1U5REQoe21N4X+0m+qjBpV2ExINI4ARjycsrb5
y9tctshrT/d/ktlDxZ5j51GW4E9jRA2kPEFgtAMqeZttt/VtJX/8UTW00H85YZa9zJuBGou3+xX9
JTZ4IFWgzcUVgwCIPKWInYozHIfCSWbUFA5lUG1zzSRT/UTJllBblurA5IlkwmqfSXtBH/u4EYlV
5m3m0Vhk5gJDLkzt8jbRvaTXC1Bwlxl+MwEHgILEM1jq8Axw+1Gdxb+zhKmYJtdKJsBma2KoW163
vOIigL1Iy06QAhLoVNmouGdDppwzFoL+A/UgmYU0d6ofPxNl3i+c0wziK2kO1iP+NmxA6CkoGpLC
kSaO8Yvhg0AlcijWB4KrKq/2ZyRXDbKn1FD2wtmQ
`protect end_protected
