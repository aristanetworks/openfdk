--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
iV3kuwHyavRP0UCwfUuuALTvuA/UUJiYxU5JrNppoousXNudgJ2LJe9sYDscEokwVexwwxTRoBs+
1UfvvdTHZs8JNCzH36f2Jwi2+GqosV2oRPOJQA/5CeqTrZC7ZvqqZgofK6Axd0bIxBZwqe59Qqa6
UGlgoz9Ih0eFnDux20Y5se9JSnboyOQr50bqdobnpGQ1Vq85m+gTKXubzPIa5MeuJ2mJ5elUzjzN
t00WCCLR04D99aTesEL4njOMNFDmHgf2gO+TG16hl4ZhSP4/VIjOGHcwoJqGWIPUaffuWCR1wadn
BDuQRWC1CNPiX7nujcoz4ag+1IWDsFGjg/GXtg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="n7BqSg/QcGbA9YSl/q5E+Z30DO64H7pdvRWmBj037bk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
TIjwDEsV5DaYlxB2fzZ2c2IncPdfYmzD6vP4NUg0d/kBfSNr8XAzw3e4NNrE1EJ7wIOTQd87QYbD
NhUr3a2+5cEEpObL0FLWOskZUzmeK0p/R4w5K5I1JhG1oDHkyUHDDDbUKZwkEuSmAaLQ+hiBjAwS
0xPuStEfYjG+12dm0ts879itEU0Jwq4LW6c+Ddhd2oPmD1d7saKQhNyIbfiEgy6o4Jy1fiNGab0J
nX9J/IUSplpkoyqzhD3w3MWJ9elv8Z7FD9JL5QQtFhOTKtD6Snnw3JrLfaKCbfSMN3c/GBYT3Hx8
CGuVTstIIyuMAxaNXOtc0c7cQ+z7uGos4U2llA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="gslZIoFJI6wei60R8HeIgwu7zejuGskeXDdsbEm05Ko="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5184)
`protect data_block
VztcaVp8XR1rO1NkLxI+IQoPUkoFZhWZE9r+daBDD43CI8DAJEdUA2q+fd7kW/unx4P2l7Sx0WBc
I4+qyH53DWs42xQOWUPQrpVSvEYaYlb8djY5yK1fC44oj8mYgxn2Pdg375XUUlrXAtRt4uJUiKKT
MqzMjh9NmEm5KHi2NcgqiU3UMj9HC6ju6XkcGTAdG/0Zz8eC63jMrEdvf+oMIbkr9dGNvU+Akrtx
5Owjd0/qOyIX/IRxDPD39Y0tLptjMe5slyL9yxvhUw5ErSA6GPl6eH27GB/v9PbZUguFiU0rfwKQ
ffWFLwkyhqpoUstWCSa5Q+e2SenafDtsF1Za74L81kL3199L9QKdeLy4qCejj2MvXh5g/rkWdzpU
lLJ+hgNOVlBaF281pmAN8A/OrkBK1En6eB3DnNuBMq8krStRhSLDNfpKGLvF2r3lra8+vXGaB2E8
4d7rAtKMhgEUJKB1HPYuq79wZsFhznLr9wAUs3tckl9071Im1emL4cNvgtm/U4DtcqY8IOP3eSU4
kBIMEe22K0F4GwlFsqGopi0ktUMgCkzNgNP94sBzHsqpLYNFF/IAd4evw/OhoOMmKkbZD3YU5L0v
z33j23iyCf4VI6LUUjRWUE1mlcsN23jECy29QiRbb/XRbNEM0y1o06n7quCqUEsDvF9Kam+wzlnC
nAtm8kyUFOT6YXUovW20rGjWl7pVJhkTUApxd1FK5B2kKah8XI0BWnw56wcYkN0f/TaK2gf8piye
NfBaNcpxwe5qMCN8XaBNXSPR8/I6FoJJMLBkoOEGlEFYDrxvEXvr3g96VVFu1hVsJhWukT4ibjMe
Ki0VVOfS9chZXYk4s/q8y51vaBPUgA/M+CJmKy0VZPjCV+SPuygSkVevF6PlfSzhRnH7FSSPx9To
oGFkUI92/kNTTfYQhdIdorz3Mt5bD1cSVlDqV6zQkIoXWUVn/juoHEZxZCh38cKvc1d1T6ZMDdYL
538dIMj/gJJwIqaBU+YdKeb9WCvCTTEXPzbtjgIIGKA32HXcNRGUc4mLjfvabq7UhQVcx8WLULo6
+UM2c7i9i624uGLzpN8/BtU+CTOWbafzhgGhfpcjtr0bMiYpJjVv95giso9iRAwiAWO5L4Wj2D0F
cYSfSj7oJATR3lV5Ofp7nsQeh4TaJW5NgMZTtwIFLzdWtLCgXOz9DKDeaGnLeD/vzBcLLfi/0jJ/
rgD+2EuuTmHAoLFNeplA2WyhTri5xU0SsMJZWbVJA24/+rYKwrVcZlfSDWjajoveN5acRKrpvRTT
nITDoCLSsUdrxgwHSGsVR+4uNJOYHg0NtyiR8FZwizvnTEnhpuSyom01YJX1dLRzNh7zHNGv3v48
Ex2Pf07WkvukxNYyHVO0dOReyHX7PPXYX0r9FJgs7vPsbt8l2bP2AgGcDxrn0TO0w1WyV3SgF9pl
AdW4AOghZk43hjyGjFOROq8qbv1nGyU3RG9qqro4qpySFauT5C03zo/IrwCATmpVTSUvh88sg2dB
+AEvjIZAFxRG1xO3BQE1/5HNA9+ReboP9nzHzoCq9uTTGGDpimcj3I/jfx5SFiLn4CUAEirZCkkB
vC/AtnJj70TDXLx92xP+uJs911uVpGNKfzohNzGRyTbOTOb4BxN9i2fLM2oQ/2VHmXTllPAfpaW1
Dwom9HUj7nHmQDBWeZLjlXoEiLaIS0L2VERiT+VHDC2g+kUBDCWpYyjvvfjRjMzXL0zpqLYyVKpE
wevRhaOxo4joti7BW9fH5IBYdYnEcWxnZ/cjYzVRlmqg3EP1T0K3Vg+SCx0id3sHLgOpduknwMx8
ZlPUWKTmBADT+R4rmjizIY674z2S4DogQ8r7RP6ImXiw5tscvfyrCQTlWl9EXC5PAnWLljNXok2A
jP7T4btMycG57H5C9C6xFcPVn0kPV8QZu43c3QzzirfHb8AEvZJQ3mM/l+uVFmgMn/NnUyoITkE6
tjxpUZ+KI3jNJPyfE8/yIymylcn66dHezuUOCQvsCXRz1U/3wMarb2TiYyzva2Y3St/A7bmlJSrE
oVv0uJCdSjhpZVALCdIh5kWl+TGHJxBlPcALhTmb33Y3PjncCoI4gcdtI7Xhp1j4yqGKxKMFworA
76fp+YE0omX4dDOmg8tIRHn1dcdWzpgWA+esCumaYzLZYWPYue89W59geSiNmXaSGBJlAcBxpbO7
9U32+5qinOGilPgRwiQSKSaYaGAo4qZGW+Bhb9klR0DYe+GKu9PoYORLURTKw/Ock9Uu00epceLx
WY60uJeAWTcrCFUWG3GRC82ayAoNf8fHaCEheZ4a/06ez1gYyECOAfT6PYwG1VQao1mLqR6w2Ctz
rJ0mDjKqEBsh35pl8bPatkcRDQA+d0OEsLHChvQKTj23Mo30sQvCVuqvgBloiVDV9lg3UJ62Vwyb
xmRlzyt5YyLuqoaz6HGeW9WDb0IV9uYWs8vSysXzoupN3J7/6l3UrekDkA+U8S0piFxR6WonBH9m
msYMUmqLW4NEkBDdrIucy0q3NvwLUD/VYJ/f8w08P17RwLukfSSCyNj1n+t5gUb8+9a8PiiZ/XWt
CQR2RzSacXZpGRO6z+eeCi8r3xalbXn+IC/ESqT/gigdOo9fpv9mDeGxwyWm/BhDDVMY+dHCuELJ
Qz8hH+kQS+JUNRyNgclQAv+L/i/Z6l7eiDBIo5xGdW2Ytv7rMVirWeBiNK+50PTIzFMCI685BiJ1
soUfal1P+ZcjX28jzoTR138iqUA+CQgWt3kxZmuRpJx9h5K7OtdTkIyPd8Mimjc++UeXYXGuCYJg
f5ethIiwMYzQv2DnxqPhg6dsJrkTS9jkP3KW+ZqbobnoTkDv+JApSdnQekANHoh/K2xCfLy+DGs6
Sq0eZZuFfq/rLEFd+tNNu4K53n0UCiggOr9em7+zPz5yvhTj6iCRwh8y58GFHfyXBlj9noxr0e8f
ZU12JqAFSp8kVIuWYSuUCc1BYZKdcRbZmC9x/HZn3ImUfdK/uQH02UF1Iybm20+1J+UubyU3KPYw
Ik+FJxh/NENLGsCRziICGqFIvOlX4z+JuzhYfrI/NoXpeGpgOJZnABoJkVi3RT/5+/AU0FvfBbn0
Uc/KhfrsqvuEWO3ees7qBDQPcuKuqCE/5njuvMlSJ4EojM3tpEn5IEldxzOZixdOHS2Xj2eg+ubi
/d4bfy+Vq4dRR5DDTrDJHf4NeGPR4psle+WzCl0+oQdQF6CHq9izIgfwAeOu9a+k5yjSFKM4aMQt
QcW4tPUIOlUNNu/+IUEAbkRtxv40eMjYSbBrjnsvkkIAqaGjuucmSUoo/KayBmXwd+pS/DfUfW8l
nbUBW8pmqVwIXri2pTXz0whmpzK3PbvyOWAUPnG/uqHmv1RM4mKUXQWwS355JiaL9uxoUmxfGVWP
dZjrI/3DDfHzVrhA/w+fip+2U7NeJirF7sYLtTJco5z6V76+NUcZ1QPovoDoWlwZo1GPXRk84Eko
p5u+VN7lEjjE47r6RMs9H06jlZdv5n795KLtWKDjB7mHkTL0vj6/J01CkMOX/fnryxGAUl0zj5SO
cUcmH09nog5g2WHCRM09odDwfbyjwmjqTlQYegKZWKahcCjZ5mD2rAe/WooDkdgKc1aVnr/Y5uV4
2eKJbsCFV/qxiRZ9DbEaAkj7Cpj4jt2EfpzkaukcJBvb5IPZp4GA0QwXD8GG8P7fe3M7NaTdiAj4
9EmSw8RRO8TB3k5Xpp9dmxK4WpqZHSqTOhqUTjORu+DRvRgz1jzq7kDloZhh1uhZoA7gDoyKa/U4
5ZpZzr3n402FS8FtSyKbEws6O3CHFagSAuxGo8qhxJB2DmtQ9MPvXDd4lH4+jKaSUkhpm0cE1Pe/
+U8N4WBx4E2eXcuslwFCvGz2ThvQ/UpC50GQF04woBLftRNgrZlM7JCYfsftaEXBlN4MBv+Tl6QA
aYQUfE82SqYrQEbgOuHSPOi159Bi6fRWqo8gg/2yFq65bICYNh+G6ZO2la558redO6PZXqCs2PIa
VJXEddUaKK91v9XqB2SXDv2SrSuOevawwAhBZP2IQQ+opA1tKKalKeRjQj5UE6vI5zrw1OZCJcmd
J5w+bR22eZq8ckA/N5GQlAwNJp/HRD+gT2EHi1+l9bzeWF8XCpV76JP+s9/qKc33+CzQ5HKa+t9S
+ohoENwJw4Qj1uIaEgiIuaUmzNStW9BchRQQh1utOlBJF61CYIW6Z+qo+Sjwd5RwEGswe3FKiywy
KfzBvVW1a1dOI+/k/kkYgXSUJ84LkxbxKMGZmQ2PHJsWpsoc2l7aTJ7fY845j+iPSA2UxC87K5u+
UxZ2cOsR3fAiuLtLZlg7xeFglhYBRrer24y5hzcjKZNJBomx0jhnj/2d51itqc2nbhNtBF6LJAhm
yUBMdJaABjGE1/Cuir64ZbCNy4gCdpxDq5XbS0qGx2OWxro4DKz63jmrdseF0hNWUoUMRYzvEI7H
gxFK8myPRZFg9bSDibt6hsNUmw1Y2dTJsiFINQPAaMY/sPLEnDQfv1SjBOl9DHekA5k11aEM1I4l
tOaEfQkKAIhwZYcZ1cxqNCJ2bYMJe9VmraOJVeHXlex+xlSfep0uz6AHAhClE7aPK5bOK3I89zLd
pi2XEkY8teqSUXknSU/0bnAmOn93YTZMlooXFBPUeUwuVYJqcG24kXJzrykQexy62CZ0bkD59h8k
Xquj7VQC8pD63qQuXa8Fh1cXfk4vtiwI6YIYy1n09to9v9mRYZgS1NZDGMixcuIqWF+AIKIxPU//
Xk1+slRWVGb5eMSPbgGUIJSEoXVqAN+iWyMGRgbwZeZAIV+uy+lO9svoF8c9tYCqiBGLYKZC0A2S
1XTCUwW+MeBKtz7oA6+i0V1ppqRmmm9dBLpKHR2VKzC2Sdnp03/x4/MnzwP6x72olfSXbEUSzKFG
UW/8Q8UGA+hDXqaYRFbT7StU4/MAmhuvxJVJk47HrLDFOilkSlKhlPqIxDznF+10gVbg8imuwG2r
eMv8OxQvHwV9XesbWPlfevKNqVG+M7H5mGmuIMhlEQJywLFocZm8OrQlw6OtWwYI6Zi9zQ5q8thL
HrCISCuOI7XkbZ6qNhj1tzgzMKFFxyXamyOkgRoV4wruqVR0CK4tVBc2eXcWGIkkw/XbswZ1ezX2
RUqINi02IOiITqLtagYgpsWmA9QAAYEVx8zw1nxpdwJJSTiycHLWc82FUdqOG3od2KJEhIEs1hgb
Kuhc5XQA0LR9mR4zxwUjqF8M4K9d1KVwBNF1x/PeWfLoqwTDTAXx7xxil2oDAEN/CQ7t5imqiyAh
RHAwSBY1Bb7yw8ljzOlRP9LHXY6+FGg24Uh/JohKsRK7dIZHxxR1sDH5xGQ6ixbLYFSnA8fYvgjx
x+F0LpuhAPKQyXvberpU0CO8sSX59OaTZMI04StaGq03naeKSvX1naUvmn5BOnCjuzUBerB9t8jk
wpqQi23XIo9Z0jaYyImJJNAd6abf0hDrpcbSgdlMX/gWbDZNoQ0zhITwq4MIAVhDBuyHl5wRUuPL
kra/CNWuGlelyroVixrDvBOL4oahhlC/fKaZ3vZkdla28tfaxn5FWrmMTqFRCK+C7jHapalIODvK
5q7rZsU+5LI/6Ibs0LwAhKSColhVRUH3auXb7ZobPAIxN3yDlr++j9QZEgY1ravwbvioU2zwJJNd
b3wa1c2QzqIRUqRftBaH3FxM5duwITmyoOj8TFsf/hpe56mleY+9L+zQe9bifSU46pk7ZAZTxAnp
KFgBoDWr1JUhZh/8Y5msV6XwUzOOxC5q7q6499rhpj1URREm7vJQj9y7mGIMD+hNLomgMMujLaVl
fR1LAFChQluLR1ZVEqCSs628xJXE3zqrjeR0IQ81LmItRmI7ZJwN81gTEUHa2OzxrYpTNDzPTya3
u7MfB8XpHVRLLkAaq2txCmS/aalysc1H/T61YXi/8ONTN9vJ+/E1oElseyuu7V2/cOgBFIpBne4a
UZmlfxxv/PTcez0inV6dtW6WfZsuQy3eAhY4Pko80auRYOlmb/nU+oHRRgrmU4ZNjF+JGZD6vLqt
N5ir2JNS9DTDNtTg7Zp9Ku+t0HQK9ombvV6zQa9vXNbjcIeg2B6+0FH/8vJhJn2radzT7wr2xQmD
QxxE2y7qwodp1IE8rygsHwseRmYTM4KXw7C5LjzOHJyFpeQA6qIaELE8ZB+UBM3812nAsoLk16HQ
KR2FrQBE9ThOU0Tejjtg+wgVGk1LPCpsOu6VP1KzgP5jyM66g/UrJmWEJOwSuMEQ/+sFw4XXb0XM
qaGnJG9z5yiBrn349MLcrHNsojMn5IAc7+hO8bObcXOvMCvAhfmCrDIMwnmpzQmU+NWicKlg5pJs
T0RcDWDA8IZwpLMEakCXEX3WYZlOmrlmVr5kg8rdivNMzAY06jq4UjZd6ShWqZ4PmV4ykI48cOfL
VlZ9MUyhjZ7Ule0uRlrjViC5XSEyub8QkUoMiI8rlEXyCVkuIvrjHVIqzlEPWt8DFw4/8p84U2BL
Fdgy5fzZjDMzMCLf8irc6J9+mFEcep5PYMj1gRrDuYyTodZcOhDXaWcLXOrchIamV0s+CdkCAJQT
r22iDYZrmY9O/DvHXK0ITkQuWO8ZLfBqePc+MO8yI2LErm06PRsv53hg7KERvGYrdKGZBSDRd2Jm
iwOFTY92zE9Q4n1cfqIjqVkj6xNHvFrVrrGxVJIMy3oa6cUOEpZZ4vvCoWtZIyhhDuFOIvuXycmo
9n7bYu04UAMzm6RK0Bg0haq71chLmhMlfT5YC82Fd8jsL33xaCU7q8Rkkd9yo8z7P2kEfeczN7Uu
HBMWQ7gf/Sx+I1cDwLP6VcIimXZmAK7LUyn3WmKD8U2RSMbkjv5/BXmKyCKGxuKZqqr3mEaL
`protect end_protected
