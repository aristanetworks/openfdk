--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
KDFgaEhGbR/Iy/r9aTgz12iNnbXH25itgQAZmqey5A7Ld82+yvaaRk9y1rqJdMY9ioBcOZfrE8Sn
8RnjM4BA9/oF/79+z49wXO28ty+SPmr4cqW8Ybt6Cgx+OI4lSrFNah237aIVW/9cRHTeBwoxvHZH
cSM/cSQ1chHETjbuy9WyGUV5GvoxAH8AHZ9vpRm5F759kRh8K+E8zcdEn0BYMdoXOXdqK/6/y1zx
r3Pp1AR4Hmq3ARoF0lx3fdmDw0Gpl3UVfFtsYKXIAyoaUkHzeQoiAA9DRCu3Zp0YY5Qu8XJSqefo
6x+9hucXkB95EporRYZy4lNzYTk+9V0rDIX6fg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="IXMASn/pjSKH4T6kdMrdZLiXCxiCLG9L1+ovs/yYABg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
j/8M9dMR6q+6YgcNG13E9lyc4aF4u3R8l24uhSqwd+7STBWAQtV/9glFpHAsgaVgJmWDeMs8ytuP
i0xmy7WyanW4QOYilbgOeJNF1TXoDjNCbt+f+Ev33xwjPQZsGN7WpMCAefP6T4VSb8VULzZpZsA+
bU03e5VN5BEZtUUm7yCQ+BX33MXMOFjwn81AF1XSXqUgzVm6A+T4DFdV1OjRoIkubRTO5tOie2o9
EGft3kGfuY5IytDnwkiGGtUSyVuID3vTORFGzXT6G+K++9mn8lQLGzUo3GEHymX7KmcYfRv5l5zF
mzn5P7GC3B78dAYQvTjMm/Wyy2LQ+nuXhb0cJw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="3KMbXPxPnKiNVRiistnCW3y34tmG2s9EdfLkBCtkV0Y="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20192)
`protect data_block
He8+Urtu4z5fwFeu8yI3oiTpMdKc6NXnsOaD5z8pjkcptIVYrm2EcOsj52kF4G8ZATrXOAY2FmWV
oZrWFurH1Z9C/4u+Ef6LmE9AhB5C6jb6BnOLoj998a6Ug9pNa8C9bDllf4sbGoVeScASyD1WOtho
bixos0ookndLDaUbv43DPvfybUOMbta1TPqVwi+s0fOFQTyAMAI4azC9oW+l0yQOzlDHeFBBVqFm
ioXTUvUgaC12egB10Mj2TYHnhR+worj27PdjWT11ZnxJQoxy7kPWWZNTMRxna4VI+/ooc7BFQdAQ
DxsbIhucTj84QR/HbiYnBeH1p3n0dR5A2abWZh3SoaL987xlnixqyeIIX3eYrcGqtupONUHpgI/A
FUImvxjWgvbZMHQUARCqyPTwyLHNRM2Si4g1UYC7h1g4nVhKjZtSa/gZhLvtTnzsfGj/jN4cKTOr
ABvZktrGeKWxdnNBWpZ2MYp99DOrfHohLECb/D5nW33NdLHZUG5ZWkKmJeh9PkY7Jo288CwewA4r
nGnKalhJHXWx+tS/o+u23Z2nuH58hEuFu4rMmiiJGcRypbd3ZSiBflK74j8Q2jJe6Ziv4Jg/bI0m
FSD88SUleeRO7DR7vjk7VHEE5mPvQ19fgzgyLjaX0Xc/Z5Lld8F472wUln4dAhZrQo2NsNJdAPzC
v6PVxoaACFYZFkCVf3Fy3PTEy/mpwbAAettQfekbcpPd7l9Ls604lMyvu3aH/L4HZ37wvTOj1nz8
DXSQSSanzPDPd+8SyVty4dUcNNY94fuQzBMWorZtcZfgSjuAQfIjRmyVTCUvaZJwwRRyi1eSlRXS
hMztXCQI1dlcsERN4TizFJtAdtwwtiuT1D3YCko/PDyLzW8UfXu/bjn21KlxBrkO6E//EXDghqDj
Exhkv75Blff39v5Ja/9RRwvuPxBZkQo0NBUEdGHMsiWLvJgxjDsoIdOrzou43cvO4y7/Zs87NxMy
Seu3nyNx1HbR3s1aQnO0jnlUgb2TqDxCVUKwEH8RzBCZnbySjvXAWmk5NpNGQ2sIr2iaUchSI/tJ
xewe2IDOU/mClrQ2O7NZB81tAG3OX9JuasoTqRPc/ePgEvkaEIO2DmmFlo7ckbw1hynYlOznI7ia
8MtOGlOgoee5rLJryjgDWCVrlJCEVfZK85UsP9D/LQGnS/jteCVC/ZyRlGOVNJ9x/r7u8G+qTgTM
bzLvZqPZkPPIfMs6ictILjGnL3ESUQaF0DQ24OIS8qtGy97bMnykI3fIQNpvnOh6dRP1fLwRYg4d
UhM2L/JSl4pUT6Uzg9NVFuLkUUY1sK1OJ2z+5aSkAUGw0XYlrJcYawrP/djJdeMUS7LDt2FC4g02
xuRiGfrf9oxQHeKdyTNft/wddLVBUd8P/42zGbqAuP/LN/c4NCqH/cTkwtR4oKaJmeRBbd7JpW7b
9s4x8be5iHfF+6Q72LTHaYzZ/P58XMV4X2k7ygbX6GuelU75AnrwK4NDba5OJcbSsXVn3cObjlkS
8ZhX8h6Q6bn3HHcczNJfsFJvd8+XS1TyLObWNWUllSdgNoeoS+j5wFYJb7QI97B00TMjtC10NzGs
VRF8yxjfGUy9nnKE83aqkrd7+Rutm5fPsBDJJb6Jh2wXGkaOri1cUNa91PdGd6ZRkhUuVqLcL5VP
/w3eA305/sUkr6C9P/shxbe2hRWDtyyu+kKTQzUXY9W21DKULoFtd/eW7jIe3QMLR+OXagsSmmhl
o9T9LV895sMYso2x12ixpVuuZNYtfR0ycSqDlG43tlmU8BEEszgDBq5v7AWX0CH9B48vCMLo6D15
jcs+7yPsEDuVenWWYRdX+Fk9LGMAz1A+bT1Yj13sASiy3Two1dWMZJ4xeL/A0N4+panLPc2fJ+AI
MzS5fqMnfn2PPQSk6bQE8um//snchFiy//wKsduRRA50cYEHpMxd+nJ0qemlZ9A9Q2yiiDPQ9aLl
HMDvjzHYTeHI4t84EnAugxlfOYpffzVXJbHiLySQQV3eb2jmfd+NgLwnFiNReWEXIyKUUUJwTAxc
d3hJ0hpOBCEpdHtdMsa1NM6S/z+VR5egD1rYDUxgJEjrryKUxdqniDIBoDz07fMRIFXagnr7HeHv
29rYxYClXuV9QBjQS69zYYZIIjkRr21h8htNjfLHVDSBuyxRVJLSwlvT8tscWBvMIg2tou4QWDz+
A8rEwPn1Jntu9QgHzOSF5TmcbCKhwO9ubT3wddWrvyjvCqSSF6yy7FA1KO6TUTrURUE2en+g8SvZ
29sYX5CTeJ9aPU18QLQkUZp3o37rM0Sdk8mKw6QnPCGcqoV1T63w5/9c8vszruXGuzoMUGml4/ee
PU3X0Na3VaDv2X80WGCns5XP0nDH20rPSAEEZEVwuufmNOgYUlMMrAxBjfoxV41T3RhKXoIgrw1j
OBDEsisaQuHFCbWRDzcp8xO5gwEyunZSCITSFCw6/VrA2v+A5AenOVnpZknPMQaW6l1TuLMY5ioB
Y/kw+/sYvtFs7xiMMDNG00nvNwF+onV1d2XKCAZILVF9GuI44HC8vN1crX1jKwlGhPdEwD73p6UI
/sz1UX6KtPKZ8tfTOr+u9FzD/MbxIwNdM7Pxzw/eNr3mq0ZKyvFF936nSlPRKQR8G2e33ZO8E/o+
hH+drAHS/ocBDP5SpmBKbtlEGg19BKNEejHvSOKPqt3mMZ5z8Nq252dW8tXxwisFZgn29UkO95Ie
5G8xEjmDNxirfl6oqD4yNEN1k2YK+YfzwFg+mOXaBzROZ3eKCyT9OH9BuycFWMIIlQp7yGkvy72R
j7eiR8Kq4rTscJnEkYamrMFUe/HOVib2cwwIzoiVUlDdzNNwseXRTvKjgv7xJSuKbJFxUeNQkVls
pGfXREGVAbCsEjXvw0ij2mtDwUOnZVnxdYsTf+cUBjRtM70Ve0Nef5vDnFqGq4kPQtQ8LRXzvF8u
T8xPJZzbXNEuEAwVWAiYSlqrYRlIrCk2as1Rhg+sFjSK2kB+zF1md5FbmQEE/37UDWWkBbpEk1tN
hAEF8fV3gxmQwnITaTMdrwy6joudwsakqQR+6zlHAliwadl+C5CoYFtfcWKjpclYitu5922Y4QWh
ELjQTdyfdJz7l60aBtJLb6m1acNqGK6AE2YKX4s3qSOcRq7fg4ZVn9jZJ9ta4uy4jBFXfOVvw3wg
NNlTu94thbYv2//tpOrK1CmzVL8FjjTxP2wvLMOodWzdwajaB7yx1U8Ud0zu0E66O2Tln//5PKOT
b0BnruD9aZHcdHd6FelOceOAItN3Lk5/72ZZiFLl6wlzjPY7DE9pPwFcl53qzxz8bGkqXY1kHvf3
BCFDXiowv+VRMpFvbZ6BHfpf3R28JnY+KzIR72T+VNiHpuslyC11+zrpttsdstN+e5NldZpiqf+S
TCG+h0VeJqWZJbHVlgsFRZC16PFK23RFDcBPT1YPZ59Osc4Mas9xEEqPbjwxlSsx27D/nUyXyPkx
ZHyp06XTufPbcbksrj+N68b5ezNnGKzNLbHLBbvfztFt7sovsgS/opWr8/uVkuHX53VTtn0keunG
2uCI16bxF0WfmnHSYjsANIVtbqAPMtmVHvT1aZBEfitIibdfTj0XFIoZONxz896+X1CO1pHYCwxi
2J0DTinuVQ5LluL0fILsuDRpVk/D2pFL3oU8BfAtLwTaWgRoQqyd489BoUnOHd/8h69w5xn5lW6N
DujETPp2NRPKekxVfNI+GeGGi8C1TuSa3McokweAkHXniEBKZqMSeizY79FXwZIQVZULtwPAVZFZ
dTAGLea87+W5zmxOk6xyQhubmrqQA9RBIdP23dFSslmjLx7f6wbK0zfmtrorf1D9W1zdsPgdC+9c
2B0CqDuPE3pcriGQOO1w1rbozV0mfAxaZUwseRBwjEuCSXj9tRhwkJjjmr5kwdEbaocgUP+V1vjX
IpIWTBmi9n2skQ2jcxrStdQ9mnx4CXJSBNN/d7q0b4oyYKv/FwiKzkSSyKInLWPT6rMQkPX08N2z
6ScwGSMOM8QJQNWABBMZ90Py5kSc/sxjoMKJw57IMLKPjR8jVTfnvzs+r3R4nz4Ssh5A0AGH/Lr4
FSOHilWWGt+R69+OJxDcLxCx66HBCEYkGDGPmHAzWKXHdIzVWbDr/kE+JXy87IF4pADVu6N6mkx/
L+z9Zer1A5oiDRT6rUexHRT8Ha7ZT/w0W0XHRw9Yui3l/nJWFgGuku9x/XsTtswFIRE2/BTAfMXB
Q2anSJEGMrUwr5GhdvQY0EKD241J6SV+aGMBnBS1gyX0AlBfhiU0s98mpxkWIuek5JwuUd8iBmH6
ULrp8tJL7i5iRMIGULtjnj74B/O/lPYf6OShOxgWBuCnJpOPb6ry5bZaX/dyEtzlYJYqz++972mj
FJARk/2KhcyJN9AZqBUMgwdrKv9AE7U1ogrjIOVWM/uDaAd2onh0c+rT23jpo1ww+VnyhpJV9K43
FZtbhuQOSPHtGoxGjJWZOp/Sa9UCS6LjxqnKLHYWe1n1Vkdun0RDMV6298xcV+yuWoZ9rU1lhLfO
sXm5QYkegdMFjyOVKpi+/rtbEstZ237clA+rMqSYQyj2/uLwLe21ZiLYd573iBZCqbaSa7mBGk5B
C9r8aVte21hy+7L8T9Osb37cC0mLljnp7af5qyLnkU/hzEKEG+IYsAMUZ2E84Yi2BN9d8Gmav5L6
9HUIKW1ZBzgVdKqjoJ3GhENgI4znjhGwR4pS17Q1saV3sEfhibd0OTFJKI6Z3hVJZ7frhYoH4axH
tAT30pLhdp7Sg6QZLI7VKMasXaYXO9NcLyn+GmGyk2enohg5KdnHBnttmEF3DYjV4IOmA6kN66Qj
PUb7zSZQxHuZ+PKpe8ooH5mMfxNCSm1OvKQr+B6o9cMuhVeShneXTZt0YJzxfcDQ/Y3xmib+vFn9
51fLEN5DQ6PiwgfrqCBq0ioQFN1d/bfdI/kjmUGKDspWEi519jxGErJpQrbFWd6s0fnUFWd03IeF
/tU3wDZidMgNPwPq9C7oNblt3TJiXg4Fk5jYx3efYKf2zuYUkezN2Gjvr+X4LwPirHGArxhauPsW
6yIgSYjABBQKIOHuEZ2k7Lb6Wb4wxcJLDfEpkjAudXWrSutf7f+0CGeBdUeKAIyMDKnkjaXN8A9D
abTTBV+UHwzdRrq7Lh9+ohmw1fljAW1EsCd8nEp7WIuC96/zlyJZGpyWa4BZ2eOZzcNmpJ5Rt1gH
d2Q+PT8dXTsiUUYg7hgKV4v5lTx9RtDD/s0l1VQWRbHcq7qbXZYmeTuw03jOXzerKyWvGWkFV1Ze
EX6SwYXJ0/duIPTDO/tiEpgXdDhJoueIJHZWpNZKlzFtxbl90I8FadLKKdutyjLkHwrNQ7o7H4ro
uxQ3JTphhYBbQ+YNsRARDoOa5xSuzqq3umEmBCHwdLG4uAvmCkmtKtKEE2v2lng4H0HYwgvGDXs8
OJ0ddoyhdXvMKVYpb5LDMYSOCQN2Xxz7x3ZCTrIJxZQY3xPdp9FguXdKvJUBMcvRSKxp4bcvedhN
vZ3wnj8sc62yqpNOIcSMRbhsDQwiPuDydxI8x1xvyq6e5A7ETQWATAC6gSWEe/sfhLzsYMg4zYqD
4XAwx/h6GMfyhCtKrpoiFIIrqkfeqOE5hT5IMHiKa9lDt1ajKsbrBIrMDwelAZOIsULUvM/tUD6W
9+2zphsTdER8KmOGSW928sw8HJFCeyXDwEg5M+XWluxtO59jquBvxwu6uhHEN8W+iVdSUSBk/1yj
YG4s2Nr+mO/xzFi6+u6V/Ivv0uijL9RsD51+hEcxvu+PnKib5tJeniYicpIp7xJBagjsQefr9rfI
IaX72WIvD0axLLD+uzh7i1DRm5zoeLUSDdZxeXuwX484QqSTy4iEQYXOE+HUBBykg6s39wE3dsa4
rsibka/j7OE5iAiTYQo1HoJsyE/j6KgGUNDOz2G/31dOAwNAVNoWYBWmX1TLbL4/T/IT7UCOwph/
PBCvelxnpdDr4WO2kB8Qt+xUkJ7pkW2NWQAam6KCTXZ75KU16uC6N5R6lgnhctr/xRYcfZ4ZBcKy
menOHl8AazyEdw2zeGenyZRVAJmeLZbktEGUQHoYANRol04Dc4jlU2dGBhz2wAkBuPHTrwxec1EQ
AI2p20LOlEDa8mBRQy6X6LVboQeMaHC5+/R4IT0DPQSaFbbpGPQJpcRTS1KRRgodLb2dNgH45Dod
XqOV+Gm75GknsAIWeQxYBaIDoAJWo4+iytduB+/X8vIiekODPPcCt9Uy4wF/z2wnUIWkGgHFFwZ5
KySl5LDK45XzrC7y6bXE0uJUQFBgfQz6P4oEdh748h613XdYOBFxuSu1Z5arFsLZrjFDHbQ7Lr4K
5pckWf4oTs+ZiQxzMutIRymQPbAXP2op5F9CNwex/ZfAnWG5uHmg4MPGrQx3eIsfJIjqD9BnqAMp
mopRL7McBkAzqY2LnFr21hZE+pCh+5QeHcxkEwJyB8OXZJuaP7CjinDYTOqV2ejUUC+gSCakT1IP
DzwUqFjjgkxYDcgj7VPoA3IZkfIj7s2AyToGh7f0DjTRjbq2yE4n5eHpvCzG+goVfDT59s04WTOi
9E0DmyhgTgxZ9A7UMNtUiaqQvvYcbcpHgO+5v1DbwvxcMEfEhNaVHWzWQIQAxKe8tbp1TEYTxMJM
cgQBVaT0Nidg3JGbP/gMNp+nJz0UkcmkqnsS8cFSVC+r9WLc9KMzjVsW7JHKDP7cd1Fx1Iv2vMvQ
8Siht/4N/6hY+g2POu/KzlGx5p32dLyFsdSvS03glmXdS/MLmqX71d+z8Zja8xha2+wW7sN/OJ8K
3C+lm598SkMDUIWymdmlJHOgRvFRD78vFS6gQrMTiDrGvDNHqCSJTRpAn+zxrLNxTXpHWj0h5aRA
8w8INXsSyta/4KeIxsdT3tyOOw8qFv8gpAdNEKh4EHs1OYjlPEaMBOK6XZxlcGIT0XCCuDQzkVnE
YeNDbajGO/u1BPYq3K71PTIS4maVSJGmqowDD4FOoBziBrf6KMIVoruB8FLwvxT5utTMzfZFz6uP
EBTilf4c/TBVD+seSICUHUqsOOmVNzbkpjLG3tLqgghu5D+V9n2fByCWviEQ/w5G3z0MSPu9gS9O
PMM1JutUOdsFkeyzVYEXEWdWbiWRtTCZNzZLNBLI5bhiK4a9zSQTZt+woh/WYaibl8ugJETyyCDT
xA/4Z+cBmhr/N1FthxUzdiOGHDS1R2UgzZZ/jLePdeU26w+2+FMowRzsYdn95FFT6/3I+R2UP4QH
dzdDEGYXxnkWcJ2js80bqSBWHW7KENc2EykWWnuqMfY6CJRcLLkNSrS/hFzXAqgfYeYHtgwLRxcA
KoRmdgT3oJ1K0KthvoqibwOpTutkqx90YyhytuTDJQCwVTV9YdIZUHPcSyAtaJEuDefiYACOPYuu
RXsqYQOfpGvjyGNK4KRsDmpX8LyBekUmu/44rTm0SylphRq2SGQLVikRzijTEBig1up34IInC6fh
Kwm/BqwYNbITuwJ9+a7Z5M60hA+IgJQ3ogvjlhldjm5yqog/r1tcypux/M0qyxiiarAmnaMWAo/I
HaRdrwISKixKjc+0bWnExGAwIw4YCda16ckajb+21xH00nze2QsYrDwk6diwfcguJ2zlq7Dl52mH
4VCL9ToY69InzV64xyV+L9zF/BBrfQ7dk+h86J3J0RoI5T9XNWhfPOXXHYJmJ3xd/g4Bn+BcRS8P
n7KcEV4iuDqkSx7D8WDCVkB21cfoHJHXzYslFjeY+bdBRpaXqjmExhLYuUv3FT0bgPNea04Qewso
OUUxuL6bOc/t/eU0hdo066OmdsfI19Zmov+AszSiH0y4rw4K/a3jSyEROdXTqfAhxbYXbICOS+NO
OjKiOzAWz/hYYK26BGKuhAbUOdllknlgwzXGxZM9FLOgkc81wJIA/0CcbLaYskXoSzhFM8C2iMAi
7gNwQ2kIysknp1aNGZDjKBw/rAqYibr1Ob4GYhQ/aNf4/A4LlXkfCLl/w+3m8nufci8pRgoHMFzW
LIjeaXFUL7MApjo1OKbtD/8/1IJLAnfX6vI7qvdejuKg6TRCj3vmGXsKQy0ej0MmZ6Eh9B3OoHX6
brsU40/22w2gYmhepSpDOT9/+KxYRwi1yBSq+PPh++GUAw3yYdc+T8lhXfXvT0H41fQwkBXPqyG9
YB2JZmt097/wXNGyw1T0wMVcnUfvitLPewPWXxzkhtU+E8YqSqPiKLy1pPilbzikU46zWSttakg3
l2V/kksqqqYf+svSvztifi6KKTAroZSIYwYp3q2gfGzcqtpByWCw4fJFyzeRuxNmXCxfB+jJ27WC
YLCatLLo3JXQeJpEwv3/5cAEcXLR8RngDJ/mImq0TBEi/rrs01m3SuqlnAbt5x1N0tNgTketXz4j
ZP7p0vSr0DknBKFvzEMtSTw/a3L2fq7NqvFBOatv61KEJNG2G9ZLPBd5W4BVxKHae/Jii0YD6KkO
eJij80Ig+gwf6GO5qVbIMyo7jYgJYL+bxjKDpMHUEv8ZaE12is2AM6oypPb22g/5L18sqtegr2g+
JKJO+fJAn0/fuwrKiA2DEHIOWmiWFsUsOrnYAEoh3o9zVeRkuJZ676UEtcs8ntMCFUDcnqRDqOoH
GoirR/fkFLzFpoff5ea4gGwOBqEYy9u+z1XuwWviOKBEHR77mgf/tEerqolbiMV5QezUzyyZ/mfo
PVC+IttQIKM4O2HAZ49bvlTkrmwlF0qbMhcfWWtbY2N/xS2njIP1/OR3hSK2cQLz42JhpMpI4V0G
PRu3VjxaF/WIdOTgN1FELpBYQ1Y9W9Lhdej40CBKA2zuIL5WjvpRhgjYG0nl+MM5u6p1v8KSSvH4
BSmbOWQi1JuwFDRyZt0EQvYCy/igUzfBfLOFItrDVdqh68+uCRufz9pqyPv41YLwIHNmJYjVjiJm
ub+ck2bqps0B65+QjpilF0ZWDnWvXNSRECKU2bpKXk9nOZOnrPDHR/2h5CLVBTwo6+DjW1IRuKKm
OiFik0g16pXAQacU76e9tgHdb44NYAQvWKgqcEScBWUeGxGLQoVDl0LHa05PpYQeA0pN2040Gtqk
rXBr/jpvDTRWuhZsFKzMSTAqylefEmFwuKB6I5Fdty6g/Q02O+4BAF3t2gUlTn0XXhRR0wGqWcUX
FbISyiiSjrIsJQozzqd25L3t+bEdPReAtZXrX6Ffl1K8CbUvY5+m1/cTxHbbCwCotnUVjEvr6iji
6hMmMUxTXemplkpNQkqAoAdKZEerOCAM+hx/G0RFPPvhou4HZIjOIQR6R5iSVoL4mSNAapqchTrg
yFOtlnZNev25Sx6FkAP2MSsckNMv9B3gUOj3VtEqpE3BxIDieBUxtn2+mecoRgOh/fCD4ltPyJEM
MhFc4NIrJry8S1WsI8s+3m/qwic5e8wawhsb63H1khJePLfjmXTIhRVoq6tQOdvQjGNksh2q/6Lx
lPETPaHimO4G84UnAx9YcCyTjR/2wb9q7YSEpxsVGJcNyUQR/l6ZGaLCbkPuI+2Y36Y9BlDp0XNB
+djLkV+pV+zY09p9tmkYq8q7pOKamk37hm8jadl6Bx9kIeL6GCrNDb0FZoNc712cO19kGqM8XsH6
8W2L7DewWvn8x1oRK3H3RHASKeRD5yultqHNEQ7AQiCLC+PN9tWX8N8ahOchi4QoPtDflpz2XYBG
MHFP/AlXItx6bQmK5cEzO/+ZLc2B67WIoEWjIGvac0JEOPrIixrmos6YFY2BFnxLO7u+tvXNY9Pw
tFwsR3pTP3Rgls9hL/+lbFomYWs8EbedacEU/eh0LJArEzWgNjKstMcigafw3Xiu/nLQV2Z7QmJW
TVWJArMaDCOkIi3fxK29ZwDm4rm+liAt2hdPB8Xn5RZJQj5wOtU8NukW2TsKni46vWZOH1r6CPDC
P5Ay8hYykpNtaqjhv7GjqxAksnFmw6ZO5L4APtHPH8yo1I01yM0sPQXOq06/bfabD8DVSys1FdkT
zoGuDYQXRb1V67VFvza84VOntjHn4CvWLgFWCW9xZ7O7nzm1RbrITFGmDHZ6FAxzWfG0lubVWxT3
STFFPS+6rJW+7cZVIQAbtH6P84Um/Jbb/0vsa5AwiCZgUJpBHFddozw4ADKFoL6fj1xezSydBFhA
abEDC5JvcWiqExyIqUpUi9hNfFAbXtLd899DPf/WiWpvsXTfFWUJ0se6h4thhsL7T4Dei2mDG4yA
BlQJJ6KhpKIzEoCheQnaN39uvqFPcaZLO8NtaK4LzWkAYLar0lQCwfrPSCVt4PO7afr3twX4XM2L
/UpB91u6ONzR+9voblNHyQOIVfenW8QbnOj9YgRFsr/Hp/2IwqrpFWJFHVXFDn9aew+58svdu7mT
0Omq/RthUuauMu220Khk3gs7OvkXF8gtsyEaRhMUAGLbXPaFqE9fY98TN1hJzyz0eZCWyP2naFgE
qWYGQaYvv42GZLDj9Vhh2Jdaoaq04m3Lkn0TxnTDIsCX3ggRhePf7mOLcmWXKAhEjht/6Vz3uxVk
AOZuWEsmg0g0fdutwvyntvhSI8jgazKadwJiZhTLEqJwyimlTkeXqDUcLarBgi/Z+bJRsYqmKcNb
lX07KZwfsGJq5rWSdgy0QlBsy1FJSPaX3D9/fY6XKNmH5MQNifxNO7tiGf7Z7MXfM3Oe3Und3TTX
P2VFH2fkjUJcL/FFrhgL7KzSUIEJ7YuFBkPrHkL+iJzTXBsTVQgRlDTaoaXvXy5kOeapZg6KBVKg
crVfShGKepGHswymq9IQF+fxYadMn3EVOIYb/6/Rb34VWhzKBSqM5O4yLrgM2YlwQrpHHgO5b0wo
UJ69iEiRjzvLX+yOSId5dKA8CxLLLGde6VyQRtRu1ZiCIjlQOexymF43xZ0wC0iXcW9oygaZWtNC
iQXWFgZNUIZmokC1onKIYilrXc9F+b7EwggmC++FRSljRpwEn5OuJ7dV0+WbNImGfM7zyBkn7s4M
nwZ2NZ/SJzHgmJMeg4GUtNx13diHMZRvtjx32DnjE/hNG0WphBPhujGaWr6PGL0NPHYprhq1QmI4
Hxr8MNZ8o2Qqpb06dy1QOOdDncsdLKC1DxnYz04Ci0H2ej6nUjtFqWVCMorZWYqKPQr+wNhpjIwX
qmNSBBT6u0PYwqJhzK7mo7V5WSFC4UuW/ZgPLm8bTmB7SFVJK+ti7jVtjxExpR7yAHhZvNdaA3bv
TicGM8CcThsiQADPBub1+FLRuznJvDpJrG6H1bkfxNEbcEsNiavhcZ9/k66tQEv8ZkwegXFXlhLr
1TSKXTRF9gRl7CwhCqnjqaelBByANPxaa+X6xcGsEk3Aq0BHhR/JXXD5i4DQG32IEd+DbJ8GUMQZ
RQJ+MVGWqkYh3xF6RP6i3EaZspZkxff46tcKZNjF7aFvzcFujTwr+jxUzV9BhwqWgz4g19zTKUfx
nybv/WggKveMyV/TScmaBj+aAjUmVjdD5avPryjXDMMjUgCD8UNDlunikQlsBhzd/aL2jAhqgOcB
DqASFH9iQUybRt/9/J/ei9gcO9UmGyhqMPc0f0MiDb+/0aNrQMfLOpO3nlIBuYDpI2OkyZnesuiz
HbkvEXvGZzsRO9182v+fnjAR03jItC0ZKV8aVt+2QU8fQcFks6ZgQ8yU2m7kKd0vWMIprcJFI7gb
eQV8q1VD0cOy0Qe1a5siSd7dljpCAmBo6X0BTx/E7Mdww/ZldYfdLM2kMAlketQKnAuUWopuJMTk
cr0FEu1/gM6Q0xgIEZVINAlJD9tORCwwic7NJYIlGhjWUBgQnoIIBUKPIJFFgbZIJBGXevXaYdTw
0lN9e4uKUUjGM3JQeQSBLWGWfQwFsVzdN3H+eRr1g8kRvIoEmn2c9pu5kH3SzUBKHadGsvjpXySf
T9AFASabZKzOVv2oyu1vqkc+vtzQkrpe5egY7Fwu5CZyyKWpg4L9M2ozkGYMp4Gc9/DlwOLITrwM
OKU3PUwj6UPWuQ6XovtVuTdiD+1FlDfoW/qHQJOCgDhwAe1CXCG1foKP+gDImWWkSMtbW+ogBaGQ
WHUiDlTZ5HQkpBSFc7r4MRmxhAv+ktkVi+DEAjnxcul5ghvyXSarvpssjoIU2mqgik8lmX72oD4H
1p/nh6PkQkab69ZETCK7PmpSCmZUITfHqDNV/64QgJlSXSWYjL93SuHd3vItpRZXGfLdN+1e+lp6
kZD3hSBijotbfg7e5fJT/ynRipqWqYZ2YX8frrRsEr3NKWNNF55LZTMc7P+cGPqWbDh5Y4wKUWYR
OA6XoiLcC2rOKDWfmbPOGtHVQ43f8kVAAMvx3r4PL5uNUCshmZeU0eZqSc6+pQ0mUVDqmywfwWs1
1en62HzgR26qaI06CSAs56KDB8j/G9ZaUrRTUHlVQjEWosnUlMbqsNTPxPCKyxmJJ9yzrGvT24sL
GUMdW8iplLVfS0yY+otWu1HATHGfmcM+6mrHjAJR2p3yanHyNuULddzFTsnBvyNYcqs8kQnRDk4m
i1t/K3M4rPQzy1Hlk+yIc9ZggEsH7TbszIZNyxMttrNyfR+napYLT7f63LtmWtyJ80Y5YlDwD+32
bUMdfdvayaV1hdtHI1O7NG1ivF3UbYFdk5FfIIDxZEcZKIxtYM1r1zSaBfia27AiBzhw9klDoV+n
pdI8IjbHisAtPEcb0qKUN2rAivgc4xiJ0rRX0s8up+xxMtfDJY132guZP1ZuGd6UAiO20xzN55QQ
tFqLwBUjwahK5hib3TlX20ACF/C8pmqGzA0afSHfxWPdXyzM7zwtusZ1LQla0aeJQTeFnBbgCGPI
YgKsDUiSm6zoJkdrcbrrBw7XniE9dERlbyyd7BEeUa2zncn4vwndjTbmgVm3WmOOtqCs+7gI3PPL
XlTlBmK59CKm95UPCXS6/RQ1rmd3f3Zk3mtHE1MVTCjuuIZ8EybD6gL/JTNb7G0txLPqR+nr2WZU
Csa9jmyOCXlnfu4vQ7QmHWj/2F0S8Zm06/ULCPUvzEdIEWMAZTehVkcxXZkBs5Nd1bYzLnc/SZRQ
ll5qNzLI0GxnwG4Zl7tIlFD/YomjxbJMo+Ba7Qzf+2YZJKioOxRFkfYoXXtOFRjiulC8bFb7Tqeq
KfKjTbvsnUIYW+C3of+8n3ht8DdlmMQem5ucIfW5fKbDz/pLneU3kLzq7fWcArgXs/M+lC2mZ4qT
nZSzo2ZBrvsb0z847LkKterNm6VTLvA07AxTNPXnXWysVus2HmId6EixrYZCuyhwGSs2YDHAjUSf
X3LSWGkgM3ViuotGYfDofjjSqoxnslsjn0oSr1gJ46MdNSLm4RbE/IUs0CMoYLI+bSNEqTxsIcjZ
NxOmMuRtWWBExPsXSCgloU2GCo4QAfOAqE5LjLaBRwB6CMMZwoqmCB4GQM9Uf9vcyl+ivSecRhV4
o5gR88TTM3nU65ojvg4K2x2wSUPRCHEfoWhClpFxezh/iWoDLVoZbVUSP8SCS1kRn08eF63HObsP
BMf0+G94AZfmbNEOlXuxDLYeCyLaF/+ypcMn8QlG/7kjODESbQlirTDMZ1jjtFJHnDsEI8iRXRZz
Iodn8+qf9yHqcuwYiVIo0I6+aGabRoy2ZD7KYIoGbZ0Eb2rXoZKfL5gQXD0ehj9uSCO48nHq88Uk
bnYyZXNyYLPmzl2fowidCFumxVOPMnfU+qrhXbUanU/yYV8rB5eYimMJAAXNAHxdvo0JCSOGtjs1
JVaL0wECYEkuAYfaM4MC62sYnNVHZfPuSWwz/BvUW4kBEIzBpfvKOJrJlSdwgQzsu3QQ3SZiP92h
YDAcVybOfXUZGp2IyEcYoqWXsjMNhuG/98L7aqjztxKb4sjyel5SlvDSCHR9YQ+7Ijs3e8xl53mt
FP2mkz2r6zZeWwkazTbAW22SGrwZzsccAxrA7G8v3o5BtLbLCnY+SN3XqzkN4UULqaBWcKiZT0LE
xTdTpIAQMGxofuvs9rBfLvNfUZUjOKh/M3HJxp+w2Xo6ARGIkuk1DHUXCpv54NWplbWdO4VmSoTt
b15GAZRT3wNDddOBu7vbsWKaXMJfJmo4z3VeCPVaErzu9HgsqOfhp9mLm/qnQ3gqcSlRjIxFIIfR
cf+S1JZS1Zn80y+cFyxHrnQZunBzVcGxy/l1Y6on1Us83RKOf2HaeLUX/4Ye1p5/H4xphCSGNIC+
ZEFj+iQAggaAK3yeUsTJtyXw9jVyuv862UjCcCsL00b3PvlOUkeGw6zgmdGFqLUO4Pi6YkawxtjD
/s4/b2xZZ5i6yyQYqZmXQwv6H+t0kvusEc15Owax8AFzc1g0QbYDDwWlTbw5/q8yPTDasZqG7TW9
WsyTeuWht/pueS4UPZ2bDK1PkkQvCeNJPXGcnLJqL5ZBX+3e7IT9nLRd/5XjRltF5Lth3uy/NWq5
HuE0mlpR4WcyIAJJuFlY6judRCpF9VlVCxfYKBULl9iTfg8jKEPr+utAoENJ1hCs/jJ+02FHdNeQ
kGXfg49ukoNB8wXX6GhrisdyVtokTh047Trs8RCiQ5uqeWIU4Atc1LhcjzjdAeA6NOI+xjzLR/R2
oGf8TgOtfrosmzTv7ZKsoYH0p3kdcl5OSlzxrsqWlwkVy6zLfHkVu+fMQEla28TFz0lJ0+cOHRAr
9CnnwhvbhVThG0BEjdgYHcrJ8F0W7BoY9hxbsvIGuzKvDnyraAeRDANnmD4bSoDrnMHaKosxUVF9
GDvVLzg0AOabShKcI0CXXBIIBHztnpaYXSIEREJy1pMJuosLIXfkRys78Ii8ZiD7LmH37l/PUNn2
V5gFANm+tr08J6qhK2ZOv/Sluj9uN6P49tDxs9uylmd0TVH855QiXCyTSohyrwLMm+K9mvLvVIRH
iBEVgK58JKUIlKidsLUAF6A/Ne4YQFsIiDRKeSLiksCS7uToJwy2//dz2F/oesLwubXy6dHR4NLP
9T9Z7Of5I3asLvg1CSExlT6VmRvqo2AuzbNdjMx9uJTzdcLWxNOl78QWx6cx9ZHhtk0x8JCRJgCA
qqY8l3Cw7n9lSuAGiFIdnMVCLL1VML73b2bZ3vpmEe60v1/I6lxxBf39Cq7P2W2x6iPiI9LHBFNh
McUl4CfAy70PpJ5u5dmpEPo4AG7VYk5boQdkG/cyx8qVv6GulWNOk9bvIDDkDY30Jfqz0z4vW64A
JrTxuX5rwyj62Yy+N4cwmcfWbvTHSejoacw6a8Ckg2tuG6kmB84ubkt/ktehHvRCuqyNTJz9hMxF
S2ht0kJ8kyMSlmAKNqeClJ+4MjJFKBgHM4lbRNt3a/KfkB1RFKHVGcycggKN41nwNNGjq8mAMPR0
w5PABzuYUg6hJIXXvHdUdYhVFSMfs5stt8DLVy4CQm6rsp8R8ZAM7obGnBxAEoCdkwRwjye3ZJZz
hvopAAkXjvOqBE4F3AjtDXNq/V8sVKuE/kcdZ3gODrbWu5WYidoPtB8VDEvC7Fh2gGnabgr76bRh
PS/Xp1Cq3s1JAEyCBu8WC+33O+fKmjlQNCYME5T9t+2mGjycD8U5K0ByM60wRs1AgxtvuVQn1DxJ
sbSpG3YmKZ0nXoYWdwT0zmvtG6x8PcTceALQeZzQqH4/6l/GtBVrej9We36piiuoSDH5yoZaTgvO
EC6jHsAF78NmY4x8lab3LbNIdZCTiER38VajpBjwfd1xNbxBbOTBl8P1GbFWbV1lJ59AdAGz/csN
yRli6hIrUA7Ch70zm4MJfkhWaVzWFt+ji3/1is2pZ9XLgHDTLpn8SXYn3ItGDdbIqnFIe1Nd5OQ1
etTB7CMDD2AEhg0sdhMQcg+SLTZgrYH69l8pUnOiPFp8yzvDUVSQ6wO74eozmEHCG1Bjw61tqrPF
w9m7TXgm/QmlQ7/sJmDR5Vkk19cAFG2zLHkCh0x8gbDAhmjRCwz2rQaIpvEhzYvNPZHUTNkCQcHE
9I1GGb1fHtresOtNfMndD29uv431d16BwfMxQkfc2CJsZLrq28uBn4iKkTY7cpHYOptjRTXyYniK
zomnOx4GWpqdAQgMHYT5LkGcPgfY+58rKH9Mf4kAEV92QGhmIueSgLdl/CM91WBrdcXybHAacSbW
LJ8X3t7tWDAnsL+RPHc0iwe8cGCIka0Bw3XGp/Cl/ITKM90ImMfrZ0di5yclPBwtda0A4al689G2
ce1PjzAGPmdWiJoqswetV/D3v/1OGSgR/mC58Vn5ZPSBKBZQqgHjRUv9tJ8NtdF8ymu+IiOrwVBS
WEfLlh9h0fHnwPxzC21H8aPso+UBoikMmbS/ZSkramkEjOz33gKYOw922TjzZ8dA6GbVAeVafK6J
rcJxhDCwNKdy5HUUAkE4Th9pn3teZsiAlXD/rj+BmExx64hONmK51q5UrhG1eAhfLzdiPfRTattz
frdTGiQObvyej+/iQiSnaAvC2LgG/di2d9x94CAVWf52s3D0auqd5j6a/Xp6zE8rGoOQhmgXDf1M
dik5QdW6iOkphdbEt3r/8P2IOvpKGF78BFcPJ4dGW85S/DuK9GoayPqASRdShN2FKFZ581dPQocl
oHqrd0vVLg7vl8pIiJSL5cJ2ystIQqVj/C+l5RzUtN6nmMTpuRJvWzb6OQD/OUH0Ca+WbhftOpho
MVZI73Pk+Ncr54sl0B5g9g2JoeMwIl08R64nG+Cnag4xdPATzzvXMQ2fyKaLrBsVNaR+Au5fMcA3
HqjHSfQ0qmEgWbCtHKTBuK7VnRPPfXg+6PBaeYP3LbQcYUADjo4utdo3DhoMLWw93AFBYpFM8zqW
vIVvq4IH+n0XTYx3Y6E3KS5Lx3M3mSR0GWHXSXpYXMNBckurn3uOb2Ka5xsqzmkEvziyYHdI09xS
HupKz/XJEZT5+UoA6DroqRkqTPcyjn+pZRXWCwKLBqGWrAvY1pecsjq7BI52W96rND7uhdysqt2A
GfeqJ/RjCVyO48+2TRyq9Fwwgh45wNSHHotiLuoCjwETULQRCN68K7f0ReHvz62GXP9dZFPLKc2C
hpQdf5Fi0K64NwXmcN3SkeeiFzT7O6CwJjD9fzhjH79d5qdnvFNcMmPpapNawVu0g9XwilVu1GVP
CbF9lf5j7WIbu0l2dV8FsOumWMKmAD8Wqs+NWa4zofmQpvS9zNEPuDsmJki78fbr7J8f89F1pust
lnzd6SrVs+V4U4vICMIwUau9uK6cIvxehVbWiCDzluvZfEHGZq8t1MeufB+CU6G0uOnJzfkuLe1K
jbxZqD8f+GtI6t882X/H8wOdN1dY8M5M7fm7zG27HD2Rp9qmTqI+ANpiWx2Kvz/qTdUwctMLuOJy
ITbQ3lgMum1/hJsSjPzCexJJzkK5/3uPXRTvEOp1LmSEa3Z9gUu/F/zMKsNSgBvprLmiIvHhklcg
jaCaVmREUjrMJ1RMNfnw/3hQx+/6PENO8+pS/hFVwkZSiVvHzs8NG+CIQIOYVK4U196jfKdn1tyK
+TBb5ko3vdXcOjKsZIWWZjoR509MtLAyc4xdsrHLRmJRBeWjilhnZ7Dnxbec7QsC5i5ybrbaUgMl
FRt0REMRad5j4UnfyVudF1sMslF88BFVEP3x+nvUkPQuyH6ZAHPJHKI18Nzu1IJyRYShli2n0zZH
VMWc/jUPSUsgse1UtKodHiXK4q7KF2Uy7764qBczpuJA9c0XztneJQcn39FJHJwOXihLXyU51C6N
3OG78+SbhEmBZqDD1mdLKbKtzFRKcFgdbRcNRVBfzpqAKPgzIQWuIVg4Pnu5QqPtOVyEUQ0rpq0M
TtuQSEbDii5Ydbvr5w4GAuPcz7YOCO2UFOxiXGkimiDk/NC/yjpGXO/KQl0AisOvY2uO0bRK26jo
iaorPmnZKZA7KCGnPaeIHtjhbdS6nd+JGnJB1wEO41woXIKY/KWzWrmSmUI3EClWsSJCIS9YEKsk
pV4fOFsONDeWnEBY9Lk/S4G5Y5DNECvZ2Dq0KV4n4FkpUhMJhIC5rsm+fI5yxsudayDXn1dhOpWT
NXfoAU/l7bk1DyIXzWjnBbmdMVne370MdemqEuPJWNt+/X1X6SFii5c1DdZf0LcPKbFfudLlCDuZ
/Fkx33WsRdcsPylXjHcXJo66lWXKaKxnqDT+fjxr/kuwhOY3Cp6u4bFEDUEBUQ5b88hWdz6pNMjj
iFWSxlo27mIURXtNZWYwkVnnPcw8QhrLgz0EMtU+nRtTReyZUQ+RMzOawJ9wAl9bukf1/aUwQDb5
aS8KthjSDNnjlwFeh7ZEyXwX6hFbENJ15ym8ydAWJGt6/LS0bTCAR6vby3INTNGrYWhEtw4d8RCT
FHbP4DhiU/dVLdoycuEN45aHSU3C6kNRfqRHImanMvvc2vn304Mwg8q3SsAZroCq3JLUaeEjAHIh
mJMkTCwARIajzCes9KoEOtN0g/oqDg90VlV4LypmXOW6jYvNzoSsf7HEwqIEFMIjBrfP6Gg5LBq7
LdB69BMzE3VCXWenxbJSwKOy21qfBoBpU8tMI6fij6G13XdPC2+SSHNRDCRKE4EK+xJmv7fQoD9F
LExU84hF5Gpc02TOq+KKMYGZu3rZu2tErtIE3mfRmIelzi6VzcE0HtIT8F9fNhbuXMAJNakJY/Up
luo6lv9fq7PeO17P6zS2FOFnAiPtAUwJp1c73oXtDFWmRw1MNEY7V6IyePEns/peKJpWZ/R6ZFOA
yqiZl95PV7E2IiSA18k65tFqVCTnHjhyqeQUzaMp+8gIXE22DER6Qw7VgiYyJJtMXwinQD90K3OE
GKt5F+u7dbh8TlCCX7plVFnYQoBp6o21hOqqY49kSnejdSy/VqnU0Vroya6nw6VAPwUyUuqKW9HE
C513OPeUEeLOethi3AEY2d4vD689CSao4PcDbYhae71FooFRfaz28wfrPf0zsyy/mykJBg7YPdCN
cPyq2/mEuwNYohLkR2GhBVxELFLMpxJlHS5HoO3alphPCsOxVYMUlvNE7MMlKFiS3NwVvUuQccWo
MkLrW8M63OKOKnu1agW4LQxfvnagQDgmJjiHYRGgzBEILNZ8MdL8cGDDgJk6nBaAKMd7KJr6vwcq
0ZEJIo5ne9eujxSi+pUnX17FMEYghpXjBh45Ox7jAQMUTeui2loXYhUdeqA8jx04I7ViuOWNK4SM
YtySFMp+GqdyQVa7yFPq6enRA3BrDw2ZoBcdW4VyhjIAKSIYHic38ykVXUXT6pDjrY7hY5lwKO9I
6FT9Fa05grIImXHbpY8H9Dyg5iaYbxHNvgL+SrSQ6+d/b32qOj+mMT4ZGoopbABWKIC/BAfZNXz/
5EMICG3yjpttmkzmt8R+inFntQSYg9qGE+ROC+oWrl+DtT2kigmJmyc5RCjDROmloz8TeKT2MwAp
C2y7DXx7c+mwOV/182heDMZytdAIOos5S4zTXJnkS8WKBbG0E3AXfY3rGe3YcHkcUOpDHOPWchto
Zud5fDd2XAI0HWdTv5UAXbCZvGCg0blaVKgJRZfdToZ5+9Plx/inmm3alxUsCypUENe1yCoPK2KZ
FX4qLHyB0Bp+q0QXZ+2ctJ4ek11HoG2heb2WcERmvKnMIxXVYr0m0mCHNxrWS2oNv7nRJheyRyVl
QWs7vpVPLbts87XFcA/eQSJZyHnZqwTxMWGJ1fknFw2lkOcQ4xYG8yvb8Efwx5roc7q6z4I6/p6k
mC+ETjkSpYSIQimPFuzZOlMOvp9nWfjW0w/gQRCyjPkv9LAQTbt+91d9LDlJwAu4Lv/I3bn3PHHR
VLGyVNyKKj4LsnTGnP6ug/5dr380VWQ8ed6FQgK7Mv7WTSD7KA//zceBtbvzOIxI1sL9WDXXU5Uz
by4bEN+6hn7r94e+YgjiBZHb6RKpJgwLM6orDlzoN9J3KT31ejqcmbmpQYrwE1lPl8E4Qu0/0EdU
Eo7C0N3paoePNwDPKDyc3ApiHaxjZOxC4HVlhssCNEyp3vsav2dZ4dvKuTo1qQjTqA0sjn/prx/P
pqqBfFOWLzIH6v+i0UO+5Gx26UovV5VrddRga8Fq2Q0/c/977BU49KX/+HVssH4G38mAfdOBDUyj
jFeZVI0IsIoI5WAlQOx5C8YgXttIVtb5fEF9ikI7RAQuGYfpKhOZxIYBIE81rnrtZiOH1SNX/BnS
/SIQ80HkFT87TIO2qL5TqB2iQzf95qBCdXqroo6oJWwsjdvocOlJW94M+JiVobrhCkTYPoh0ItIG
Xkhbs4OdCW7vNzo0HqnAovJWxoVT7HK72R3rY6ziCTaE9/3y6u6ODjoSKoccizwbK9d3Zu8l1qBh
8Vr9FaNJ/637VQQ1qc/Y5Eh9zgAnuzAU4rl+M8wTMEp4j7pYdeVYIuGdYQ7X+/zEQwb7A/ARucf3
02IogeCrYQI6OTgRwqMxNdQePh4QZpLx0X3Dlql1fhitrnFRwltbZQJ37vqnKsxoN/x/bAuTRF46
LkQpVma8S3Hp7XSEPIWRwQG4YrTDKfUpU7KIZd1dRCRZqWjaX/c/GXXyRxacrut2iZIM7ha+9fKJ
l24xX2aXW1PvH1gNh/mwsAzKUyFAqBw0+h2gW/GknOOI1rlDC3VKlCbOuOj6/xOjwIs5569ElDyT
Jn9jG3m113H1tWBTHMJ6KlTRIkjxqZv6O2AkIQ9AI0t8ZQ9l99hzTOAmkOpV7FH53NZAhiwCVROJ
A899UOJINIIUzhriqhHvr7rbFSDfcxO8bHEgwBwRoGNqDMiqwgDl/Vb0nep0sF7mt6RjiZsSpBBm
t2FwsgIHyz8Q3Cu4prS0kaIMm6GbGov0fBTG73I4ZrR1SzTgzvS9y7hdCd+arlcHGqbiBUGC7jMa
GAd+dWYPHIUzTPccWDKbFaUfZxiEAZqqQraw+IR7dUwZNEuHrw3GO73C14VI3+mlpj0qm6R+UwjP
Aql3QeoS1oFc5WcprEjaYdQDvERvAhKE2YxivtAq3ZORRzyILLIot8fVkTb9XF/q4K27MjCGhc6N
A3aqLWOHVYetcRmg8/JBbUrFm+q2PMEHaYp+gr4zW4CRqEORiR/n4/Zf2sBEY/fkrAXuuLe+5UCT
nMNtWb7+SQrGjeDuDeaQsU09RxYLIHNhZvtwxtlyS0/bxrSwC04XV0qVHPWVjx3QS/TQdWVlHrJZ
0+Sx3jUHzoarJxi4C8GaisQG3B6ioGYm8BMSFK/Jzesdu3XSo6FeZBkrzKPIPfdMPb9II8dWiy3P
baNmCed2eFEBDSecfgaq8I6RgBX2tcR7hHBmfLjpHxWv4KmsSPJDAxsXSH6vHJ5PQe6AD5IWeAaf
hjca/pXxwjHw2eVIgkwsE1rv1dd4JZ0RNr70evSHJYsc8vfitbgJbnzgXxWKKzwxljOJPKzhksDi
vnw1jAOVQD9sAA6I6coQatqMEIhkehLSLkSIQ0J5I1GoR822ZnWQv2rMyNYdUwxrMvrRFJRV16wF
bnS11YzJIiRa7u0zfPONUCEORNSNSkQoSOL/txCuf4Z3TvBYKLS8hOAGejizynecDLbxxv/399wT
v7oaYc5EJds92PRFLXtUluzeWHMKLI+D0PPkASpY/x91IjmyJJ5e6fMT717uXMl6f4QLs5q9YpnV
Oy0tlbDZVo3xH69g+fjEYGZEN5xE/9hRe458dzjzo5NjQUMtyTOob2/eX5kKc7sS2o8hpptzBoxl
4wFRe4PXifXZAb/rPeAaD3Xyx4mpfHV4S8zWf7qBbyuK5a0OLDq0B1w+JFnaWGBn2VyNxZJd6PXn
gtI5gierBn7U0fOtKVsFbZizWEOmwZ8j52cGKz56bhziolX+GmMPo7lGHsVfJQoSKzgC86Ina2rE
DWZN5j1PVjo9frd6gU6sCCfCSDwX4gAjgkt2djvcq/9uujbMS8eDDIu0kFUDgZrqbHrp8Xqt32Ik
clQPrUEsHuDSHPYBkBd+GIcY2dBfhjcGSJ979hiZ528IR3QivNW0rRwNDNAGnhYzf2yKC1eeHwte
qccCqf6LQwYRq+2UFUGQ/qNYEB0d3zXgMRvv4EcLdb08XwEYQH5oof1IbZloZI70gLn/qYYW0oEm
/iJEnGGIwa6D7x3+tICzKGPSYNvzjREdB3ocy0Q+ehaiAZKKdsxKFBvuwuEIBU/s2XYh63sW1O4g
OlDwE0Va6lgvYrE9/Kv1BHKSNnnxRBYEu/szM4I7H/6YBM2c84di3L+c0xy3senc6u8e20FpMerS
jBtd17VL8WTVLOnhzOP2kEcMOz6XpBDmNFYQnE2uS6/jJSGnCVkFN5s279oySo6CdI9cBZHQnkjH
ef4zE07b+cA8MQnaYpFRUEDEAu5xG2JBQW7JgAUDXw2X9yhXv6n/HLLf9gQqYj+XWGqVzQvBwYzk
Dby2XZeklp5hUKAAyGuMhP40fKklq1+mJbOwzB85jm4oNmAO10iVp5YGzhsoW4/2hpzQlvvuYmm7
rI8B6uB/d8Q/6YihdtMkksXRx9oScXG3MtoCg6EQ4S2C+hc+qamd70AMntYBww5W1qMy4LpvkqsB
7If6BKPfp3Bw+MIObOEyR7E9u43mFsW0Ch5gcncTxHWnZaqUQmr+T0/qVEGU8X2hPydidk7ecFRP
xB8lwUuVWrh10UitrVq7uUO1wLJQ+nto581P6yH6P+Sz5zqbarmD6CYJZLRGk4MjDUA6CeqSZAdI
Ow+zw05ZqeS8Zkqpj3bDy8sAeOJz7R7wrdjq9VTAjFxJNMyrX3/VGKQQuwf9KVmVswtXOkafS+VW
VPGfxHsPw8nl4VPatQtlF1S5toLdjW/FNeURBUz6MfwDQRVTaAxwh1QFnsEKobJRuMG+uKRxdW7P
+ZCOsW/moSVxMPwn2d9RH6Ognq1K9vTXgAUkzj39MlXzBPiwtFSBHu+M9t6TXrpzExHtqDPRY+ya
e50CTKi576vJ4/slQa2fm/VPFLDbcgBRoD5B7LGf/kUa91MqtJHtCqJEiH9JYRugEE/XWqdrlTdG
VBZD3DsZu+COIe6Lys4RMjo5zx6USfElO1lqp1nFHJbNIxoM/ODyXzHwgcRDmD/MGdOWqW7VyOVh
mwOMLSDhbZ9WF9EsPQ5AMlbkEkYKjziJC+qTIaV28+N5Sgt4tNeM8Cid3TV8cP3xHgtwWHDIr1tY
BLZ7c+K+oP4VQ8ic4jEt488ZuJaT9dUoDz8KP/qCZdDctXvdFqJVQTjux4hLSs05eJegIAPYnatW
GQO1ahUX5aLrZ+noWYS6WtHsMxXIJWFBSdmCrcpCZ9/imBLV5fe6wzGLWHAzQOjO2WFeEizHQuOh
vJbIhrAEo5Zdu0YurVPevWSBw0prkksC5vWKBxRerdflIE34nzK73c7tr6d3CrPjTW0uExAwzODi
FKF9Ssj+Nu6+zYLF3tlHdZPZrDAN5O+OQtS6rFpeNAgKoOzeRthdc//EYmzsi6gsVvJyXd8E1/4q
25PVbmb5eOgV84TmKyrl/knbW8rbQTUxow6HOzbUqTV+I2W9tBBoE51J/+EJitjBcmcMNI5EhCkb
9hL0cgDqL80SY95VBcrYDSLYy2mp2aM+xG3GOzzGttqCnETjsFQR/DFdf7C7dlmWJBJMJTmusZJb
ZkycMK1g/+bMFfB6478JrBdQyfQeuUCPahz8bBaJKBDuvT1E4/DM7Tej+p1Me0aSppUDDOZuubWp
A/wUwiL5nJnSV71gFSh6UzYrZGJw8HwGw2WLM3pYj8Z4m9/cIV+u8eAbQRPhXENx4vUtwavA5jfZ
1EMg4n3OY1jOkw0ywc3oH/932rdK2nOoe6u/9nwuSU30Ku0glnJ5P4ozrD8ak0i7IRGhbQkxw9E/
8rcIHPC004h91HaqnEIRgaFDdA7Xko99tTPVr2REruIy9PVixFD12k94382yd+Jmt5AteSj567DI
PreA39TPr8rHyn/ljoNsijPXzVDhCCLW8UPGclCTuCnLbYGWMGKwz1UnoqsNP6i0K/5bpkOceQ45
dhyXnNcISMBcda0DDy6Lixpo/lK2+2XzmhIca780VF70RWNSG3GS2QNFnDhC4J1ww3XtupajGesN
I423HIbqUyoAUXekvL5eVFiapp/FbVCUo2Oa2IlzCTIffpXc8TpGAOzs13h7xpDJsSzvSikRIimp
UZ4OjmsPyJDcAwlNrS94sdVkRFAE1Yc7NX7yt6s93gwJLQLJT9PYGL8iYDC376VLBTbatsT7pLqU
ysqmSU5gnE26/2MM/YwhsCP3kiZ7DhKCcQtJai0OjGcM0OOql4nek+J0g2Ya8bF3KO9fB/+YtJxD
ka7704snh67djyIgwc4szpfbv65zGw+lEOgCoTkWutHiZ73kxpqXKCTCIe89BaY34S+svBFuBU+H
ChIARG1vQhPO6sfPXm/zghRbyjiiODx3DDMhwGal6zQcfdslbZRY/MCZ+Z41qTsLTShPGZJbHoGl
4KqLGXAwl5Ch1d6ogaD5RP8LHdaP2lK2e5ZcoL8pHinokcf4pArFjOKmLcox92KPF3f3xhPpgQ6Q
HO7DZxhVkfoOZgnq6H2rxg21pl7A2OhmOVGnYMRSPB+NajTPziychgIFG1cq+OL2+s/06zFU7tGN
U2dklH9mN3qY2w1UDalbieecFC+UajyvGEW610ZGrZX+FiAt3f72P+KRWILzQ9aGv0D5kNOt95q7
blxGTGVs9xHiseFqB91nAWLfCsC06S6cO1N4q+quv8GTDOrBjX7+E8pzqs+bKzMTxeU8bq68zJ5A
WemjfasfylUMPPfjpFjVMCrpaga+H6pmwtvXjnefsjQzHgS0ayJmuya96wb50bdidRK9pJUb9S9p
RrpbBrxc2duhtPDtgnatEBbD0o4aTzhlDJ/6DF8w2YLY/V++WxVjKdb5AeawyEu5dMmo+i+VVzP9
Rx1uTc0rVRu0/rervgguym9VEfJ/8FK8ZLBpY0lTBUovyKa+RcCn6CBXFhkAOn/nA1BEfnWzRXYL
qkvcrYJ1nCVCpXXHLLUNmqLPzFQcqxrdiTJMjYrX6z92DrkaZ9wzv0WkfjojM0hxclo2Ky/m4kYX
PdUhyYNGCTbffbli1vKlcc2TTryoRaTAgfMmZsJXfQSJxA6gjDYj6041pWWriP7AqP/q62i0iXTx
Ya2JhnJCz7Wku0Nrv2Ob3fDOLiSNeEnOB6y1HUrCPuMkf9fcDBPuIFf6LofZDYKWW15U/3X7doyR
AdCmR4yI7nt1ykSavZuiAJYhNrya1pGVLn9AQdIqlLLtR0enA/uXTtYmzSE2W5csL9HmUJoXRWOP
qEdo4+w0m67l6bdcUpFkuBn6k7w0nP4oLqKhF4RPXimPpsJ+Ps3clXlvocDD/olAqPrUCLVaEpnZ
kVofvvAF9/AdK2iGuYw+bXvznU6RM+UkGpcFwPSeGCutSznDT1GA5BbZZh8jZ6yfVODM4Eerjkyr
Xm1ctV0n4P7qcxaw1qjKrmaky3Tfwi1nLzJsiIvB3xqf8pbYY6Pc4z14OUlRkGRyeDTt9z/ZqcxQ
nE5ng0sLq7INRS85fz+tq5keJ7EeIVH6/oUp/T9L622vfyqNCEyhmRGbIRfO5jhe08jXfUqWF2JM
VY35RJmfSpDUDwy52eApn6ULdXFnZZG0gwTJyTM2r21jeQwQK0p0YDiEBIecYfqsBDg+WwLAND9m
9CEzp452QmvKe7kYGZYRYEdrT9wXYZMe1p7UlXk1nrUKZF2xkdA8rkGBk/+wW5J9YBGa+GgTN7kt
HI/yRjajNq/yKAw/nu6sDRWfYIy0ytWs45CHb1G94SSRtwAuCJAOtmdbb9csKECRIWfpWJOxz1E1
EijczcZkQ2m10j45NgAz8jgWfyzvDGAjisOAxXXkBKbiqGpEZNOe6FkMOYe/wBRi5FM6H1iL0kqb
8ZdL5ccJ6aTPVHUhXUOs9mye4iFX2NJixQfTfv6kdvPINcTElDs6fConsROlXXI/p56l4eWuF6Y1
FFepibmmc4+/TcB3ayrhvl87tNmw9Z/Jc70vQ8ZRPOG3eZzwi/U9bXAjqSX8FSaCQ7kxd3nbgDmh
+0knUSjWtd9UM4gWYT9mivxgzV9IWauyLrH5vK9IVv78L/TpPNLAiq4fLiBM/gTq8XETFJksGDoN
WM1RCIT948XV+Ir13vJw2SEKSOLo17wnr/zwbvqMXn5wlSle/tzWINUbTIe6rL5br+mtFkcSIPhs
hzTbzO2kxHhJ4S8W9cJYXbWDSV/PQkbmk9l7Jd2KyYQps/QCemRTElHzAyJD/chtjA9lu6I3PvTA
iIUjXsgPvWPcqc25typm5VEmP8aTLvhSUrvx5q8gbKrzqAtvd/3iF2w4wX+bne/HdXLFG65/+cM7
ePAyWYfmca7zH01J9swsSUqyFDm+BW++4xcEf1pZP1zs1l5zhZJLwM9nVqNoYMmTqXcVmBjrOTOg
DByM031eUPP79L8FVUmjY/6aVYtc+XEQU1soMam/9vXeqU/58coCf0Xa/QxIIND++UbtjvLyihOZ
raLUfazJHoaeNFmz3AFf5ePwf2CENRUVuADh9G3lf5JvIZSBEIpG23GsCqlwOEViGxqjboTZnrRg
YG4pCrMmOG4fsmY/Fmts+zEMIwEaosllnQSBo8p8OCxt92wbfIbybVR+Ejoa5Z08dYcLW1dXZeqi
7VKbZZ+MUeyFIS0CS5kt377Rcr9lE+47wOCCb59XW0joCXM2801YLbbavCZD8a6aUsI0SbY1tcAt
4Xf+3OJLl+eYliEh6slY30z0bxAk98nGK0xO8g6mxve3w1ooHrGw8CZXgBXhGg6praBha6zc2sIu
2UQhyNXuZQIWy4yw4Yb9F8poS71GaNw6snHUIc3gEn4bonUZ9V8LZmL2QoQgjwVWizQiXpvQCeAe
SjQYt507cVWh9gp2GnbBstsrCyv4d84f6/zVO54CyZBkKP7mE3Tlymxr/WZAodc9WOkvKA8z7lyH
1WbgrOx5qFtD38jHDeY=
`protect end_protected
