--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
bG5Jvlfp/9AJKjO3rfWElHBvr96NCAc/gAh6etUOLEseeR2Nft+sSLb7gwRfO60UL5Oz31Bqxlm+
RuHikIvg4TlFuQhnnV+RUpYeswPGdXt3nxnZTkblUVXhf2ePxydcdfhLDu9riDcOuKAL7fc60Abv
6mzFXEUFSv8w/oEwsDvftKGTnRjZp16jKwOlgUiO36juHX48nLQQC0WVtOw7IMJawAmS4H2QG55V
dHXLJTGkd1Xl0Ssiz4FnGyaP6MuVfcJYBoZ948J8PQK3CU3heThLHEkl5OBCJz2F7yucJ1cMPx9c
5Yh/MW7sE/jgejug/GrTB5CD3GVTcYto5PgQSw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="IXaMEDuyQZ1noK0JXDVb1MfFj0uyOOzlNY1mfSNaX/o="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
MdVeDhr+69zna/xM/36mCjeCnKIN07indrT2A6OJ/KH8oSZLRGUw9uMKvRkocPIFsIJ8EBGpZ9pT
k+FvyKmwOfmV8C89Zxcn6xC/CprpEivgn5Xg1VUgxA+PIHUGOjBtmymntTnv/xALVUHwd6ubh/2a
w43zg1lbdfam1u270oJ+uXJ1hRFiPUlO5ukLioLhpOm8gEFMsSL5lUbDwM5/+AC0k7WcRfUnQtxZ
o0ufwt6YfvbVj4QUzcgFm4dHbJpuNYXoBL/g0vS/xybNPp7yezkhzRgIbpUQEmQA70PIuYFd4+qf
MEz3tPcmTXoh5FZjlixODfv7T++Llflyh28QVQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Dj1zYXqm3KNMPX0rckl11ykdYDu2wUAVjoe465JMKt8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10576)
`protect data_block
F9tVVutrAyj7mwSNosn24aex0DG7RIH2hK5yt6CLya8BUclZlydmdR9pX2tXlMFirB5nAkZ6yt6a
OL6gOQZdjANkSUlu4lIGqnCHSHcuzvLtwOsbt3zMfKEBb2jYqJWizX9+3A8JGNpYM6iRygRUEUdP
kqzDxgk1eOipWKpU4+oOXfkShkcscQVps1Mr4LMnZy3J/jJzm42sBvN3C8QA4P4Z7SdH8j7/MbDw
AtaJU7sExHxRYVxLVDGjdwZvEDNzaguhIHudxjiyGuxUw+FIT1PfFpCCnhI/fZSvZZ+EO1YjJb9p
nva9Uyyx9G2Pq3AWpZG9eB+GmRiYcuEeGhdU8h14YxAWazP5TIlwNAJR0VD25+mxsNy8rhQfT8ON
oJfW583WIU0SgQZiF+lFeIg3xh9PeOf5tfSLGvU5hSS0s86lviN/HA+7k3yMmKH/dpO7o05aH7+Y
Z0jF+0TgThUlHeCZUzDYwxOHxl/eb76aFvP32ttRIp59kiBSoY3JJeiEqk1E615FTsmVUUpIMv1X
VQppH/AMKJD+ZK2Jb+842AqKdvhKNRM1sIA9Z2h1LvcZnHofdfwms3gARLjXZgLWK7UIKdZhkLOj
hRIzdy4rKhNY8ZJ0/PQukfAKOthp9Bm4wApYrINCqWT02k4E77MLr/FVj15Ic2LROq2u6fKYq3VV
WKH6bbqdu3jWsYlhwvoKx9fga5cFnMfkJm/rlszYDaQsZUl5ZoLQtq/Mwav3nzzqwt0Dk1H690//
j5yhOF25nwY8E1S102gh1wE8IdByGwcJbY9R1ZfFWh8pnPveR2Ua6zKO3wgjP90Srx2aLpgZ5T6N
fSrKXiRQx39J37if7ACFuxetSj3h5LlPWPcHh4X0EOi2Q3uoe4WEg1GRugu8QVgiyIl6KHPveBEr
mf5q5Fhvq+5FwoZmLX09VpzwF7ymOvXUoqE2KFG9nk23EV2sAxowAzpHi/XKAfpvX6oBMbwRyoww
psDVTaw96o9RaQgf8BYyEj2saRLJXAkSpUs6LEqJQrnlIV2nRj/Jlp7s0GGSB3O2NTqjlPIC2G6b
XGwrxsZBqr3mOe6Ms21DtMVM88UUyPuIgtb5tzJ7kyCRTJaKUAFsZxFBb4I29HugCd9NnpqPkkhT
/BnyBmsPA9Mayz52BxIrO2AhmFOLflJW1M8dgXr0grwqzldDrL/H1gkHecBbL16Nr54G09X1xxQv
LmObeH8NLrio5cSWymBvSMrC4KOlUyYc18QLlhLmjGahyO25euBpCFGV78kci8KmXi9ZCzhSuQGo
C1D5iS+8h8WsrBMa/MIKDs+0HWfAmXlO9BnfUyHxp5aH0VUyy+46Ev4kPAZu0WQwckMQTbMCPS8Y
FjO93Wr6yltv0HO55WmugfDJmCTTQ+ongHMelXyW3lyqKvwik3IiOAQGXrfTUxGMY0+T19we3dMA
X1fYvOMGdUxG4wUdrh+tm2jvxx5NF9WPJyagXFGuBrlXr8G1wdT1/vnDYIY8dbzi2C0iIhGiIrtY
4C7TjKMg9A5qDudL+d8yztNmqFY1xQ2yF7Go9yVWjG+JDcOYSQEyK/Gx3Ky1lFZLEVHuzBEAEfGp
ChfDcen5Owa2V5dW+V/aH4T8IYSjDExKWLpqqH0uRW6ZRfc1cPe0nXmm0OC+QuERC0DmuoxfFe3i
r7hq0NzjL6iCyonQe6txxKC9z6JbC8JXhCZKLz+omRRT1sLvDc/FQ2rEFPiCaLasZxyc+eQUtA+8
AiBg5rnkaVwoYaiWsZKRmo0nh04H2YglVQVtgb2JyU6tSTpmpkDMV2H4+zl+Ka0A3LTTkBpR0Q53
CfqVtaDYkmKo13JCTw/AkxoDprSLR0QNYFp0wXsm3stA7FQsqhvpAlgQ5RkGYCSNPjfpg0MG4o8c
j4BsopxullIEbx5wFfmqp9tJJvqE/mtLkN/hoMXYG93BFvZsOBl1f480oa1/Cu1Yd7rLBj5/L+Nv
FZMY0jzzNdOZWsAIlnjOsSVw861L0emhp4fr51RbC6kezsoBUJI4AHfDdxQjuwhRgt2tHHCfy2BT
ZYgcrLDY795OlmTfWjf1lzkkk4jlKTtzOs8xzmJIt6lwa+t2f+AoIzOulMeoNkvTx7SJnRxCimAg
8FaI4sH83siKc4M6gyQOCQqKeq9SeD+8FfP2pN3CGM/ItGVw504YpE8efyQY2lk4WUsD7XZ7BY4u
U4RoquoG6vP6NfqevOot/IQ98wV4uB8pQb1l/As5emRj5GzYxP9omQfH+/yRGF8vv8Y00o4l7lRW
JXlx/iFEpwm0SGQz/iTFUU1tKkTJwRqrXE7g0+ygYLtK4wIAfYV3xbuRwekaMwdF2Ta96FUcmIzA
nKn0sZW4KqT1sT2dypXznYNm7HYNZIkCZLfD3jPjJH63fZ8anAkMOHyJ9MlYbWcB+LzeEQrxl7Zp
fPkHckFwuCducEyyPRDZTmvJ8zG0cikzOr657YJamajAaleS7CSxz+i8KhDB+9DpzOiBQTmYDf5p
sXAr4rptfRL2++dQk43cUlqPPNpp1NaoeCKV4aLP521Ej4ns5hxRnHDT67imQRtqnkW8JCU7KFkH
K4NxFkJs29ZTq5eelurPK4dVKPQ6wn/MGirJfkiFBT4UwsA8bsMI3BmNEvOsRPhRUaEs3kEgkG/l
KMeY8Am/5iVhXaaRNWdM293pSIwdyOm6ZFcwU3D5M4At0Nc0P/XBjzMsbss9Ri+vKRdf88zukr8d
/ntKQJGNaq5jWIVKzgpnHcqPdNQTsAI6v3ZG2z37PiZP4p9IvoF5Eyrv11hUTbPART7RkrhtkPIh
tdK5xDEl2lrksqN58MlFanrZiww3GKjXmdFcxypmnVA+MM+gFAdu431L59BIx7pEr5+D0Qj9uHAE
BY4ZLFHvG4DhXo0ZE50ulVuQkA42BXDyAyoQHtJRxqZ62PhWnMDcKKaFnUtMoT2AJVqGG4Dj8Crt
7T4nGS9Oj70V9tQw1103B772jUmLES61m1IeGb9AVoOWN8PmGsDou70fmtwavNn8V6yo4yHQEU1d
C/VXSFelHYjHvCOP+WQ2v/v4iaUrdfp94hfbENWA1UwsGQA+bByAOiCzP+yGVFZIIPM+wxupjEIf
Gs/NxoAQYy5MbcVb6+AKct3qsviUInL9aSYc9siSorBvLFNqOI/x2O/UpjHw+QFFLiHHvN2Y8FYk
u9AUkBsag/3RJ7c5atZnYY+ppkg6ipB3ug/rKvc4blPCvxDMYkrS+HiHyVQfiv4+D+IQLbJpKNgd
62tm8XxbsIisrBv+IgKMr9+xreNcO/zmXo5kSILB3nkBsxt0P17H3kbj6zrXHGw7c0VGqHLBVw41
0XggtWQ4PwNJ4rMXT6JJUl+7AMHnZOeBhsFIRbrUsXK/zJZEgluNM+bhQCS1DkZDWvXBWIvzL+p/
1PYg3CbCXOgk1Z/HG2dB4FNtMX8AjY/ToB/WYGk9jLns+qJSDl8m7shWxkGPK8+D2mzGhIoU4PQn
aTsUYWuq0GnkZAKZ0Y7IPIAbb4Ifv202ys2cB+FztCTffYvv6/9MM3JTSdlF3AuNRss+N7DUgyx9
/qAYdVIToqYoezoxglRj3LVhbjT5o5P9lBzA+wXzMTfxvYGgtqQoqz0RvduTpuNi0kOUGdhXVbkf
wD7VEmMW44C5BEr7mYyPz2q3V1So5G8BTUT5RlBI8NUA1Tn2gNMVCqd0pddHOAa1mqOmTuYetNhd
UG66WofNOYl5w8xdgEomDV5pzItEb+RpahMoy4gQa2fvnS7g5tZYmPOx3pfpNgUGCp6hhhKx4jA1
sj1+qWE7lgXv+EwEjVQx4gnGone7oaDgdjVSDiC4JhGIDbvpU7Y1ynqzDNxmWU7jLS9yVYSiD3w1
g1MflKiuWBs0zjCvA7CQpfxdPe0q0BL685/8BU0ZwiitAnxHtzhQNytT9A0G5Tdco1f4qmJiPu+r
zQX4vmr/OtVU7czn4L0Z8YzVTLQC+EspTzDNGJYrt8JHc/diMDLLRq6CMATyowuUMtKLktludJR0
2nSMWfP3a6gSSsBuFmCe8mGDO6TpIZhf1pfRiszUMY7hJp9yv/y8QSoQ8KadoKHWO36uaYk5jcV1
xwZEusJYFVRlcsqrHkiUt0oxytVYDsmHucommEJnyDpup/9Xe1f6NQRWLRXec6okfYLI3JAV6XwP
k1hhemPt/4+vJaeY4XIpDzGAzrgPavOzo0bjviZNNOic/VRTwMqOXe9xfCGt7ZXsNgubdGL5/cNv
IdqjwMuBTQz0XKy5gbD2tRhmFBBjhZ4PvvOYjPx4W7VySDaJi3Zpgst4nrelpAcQrlF94hJqXGs2
6MZQoOBdAM9itv6QBzaFG1O1F+ODBfG0Ifp3gaLY4+QoIIof4cdYidsZpSyOXQG03i1GPH44d7am
1b/4yutCVKKYV7DMSQWgPoIqegu9ffUCujNGCzfzTly3kozCLlEDszqmXVQ8EvJVRFmRH3wYfBxx
MPt5t6BLe0muLJuLTtIhpgDBbmZkVCyGdSpLcce925XMsDRsZhHZ0SzN7fABKmw6OJVr6p4Q673P
lfUjjxO6iAA5hgHMd6nDy/h0oFXGS6YcSDQUqtaxJsDnnE0M7BonX8+REZtXfcpDQzVo5wNM1uA3
IFOysEQTElWxoSMZ4Lqft5scVI7YLMzl52pX+9O3nX7tmktxTWMKABZBFOK1PKAp/VIJZD59MrdE
eN9lZnsFlnVp5pHWEMMY506NtuEb375JsG6/Ysx9DUTQjGdYaD2C9oXC8DH5V1gnUrwao8ExEIMe
PX9UYalgiaruqpZ/VIbVS9m7WgEU9C8JTR7F72Qza0gXTA/y5v2NlDmBcNQPqNes5myg7yMysJTR
juOkzmM3uHS4GG/rXJNoM+qiFYsHX6SpZwRyI9XSxMkSXixmJ8y4rq42B7JnDLEILcl3Pwm+0lcj
6nQpvqSA/RrX6SfIZUY4HhWt5ap0mOlFwDFxcp54Sehp1TUO9fzegdKzG+vAk8oGtpu0/HP82+NS
+dEx3naTzazf2BRcqRqIS6wfmqgLt2UxY3+Z4jTKl7SpJ9Jj5jXvgn88uQaqsOJaqVCba/1iO0QZ
DXaLbWIE2JBDzsFmc4VO5mJvsAHizjcgbN7uT5N4xbXA19mmqV8VCLUqpzvwBMU4Dg/jU1vO2Qen
71XqKyxcO6FnvLoeEzBMm7r3AszhoP8xGKxwZW1j43dR/GR6tyyYd4ejHGoquQF6t0/SnjemWr3T
2n1UAw11ECU6qkFEijrFNiXTcMkysrHArhENHbLRIf6pXOfj/ByJUPfaQQbrRjhwqPl3x03LGs0v
i0IxjvXlG/6gklUK0LJDdq4KZcFLWN+Bze6GvD8HH5bgyA2S4PlKiIdtVcBkOtf13mm8SnKgVh2X
y7JgEmi3z9ejXKU5Yb8WuTSB5Nezp4KTNRFa2cX4Oc/evvsd2+8UkDBiQkef6P2C6TKoSDszRNzC
wIXx5Seg3nSkcGjPLQOmVmfqh90RjD54Y0LYupzpnqaxkX1S2pJGQk54fXpzRCWQ3EyUYnLB3KTF
8PsjBenKTbz35p5RUWkNDm5CKZNPZE7jlstMwIXGVFdn9LBNdR8XfsdofHSsuDcCFB1CCemeRjcQ
lObQwRYxY1l8IEUSQ3W8ieAIv/PolHt8vhArLbSZJpx1XQ1u1tl2DCsYPyW+RI9RNm23xLQ0TS9c
fbTG1nGJMvTmWDjNzRAoKVLSTYcIBiRZi+amQEtXOj00nPl7up9H9pdC+uUvI8cqqW3JtNpO2oRf
z/ier8RoJYzzcp54s4qSxZAn1c04pGm4mP5J/mH1MYYwoWECjE3gfATTSCj+cYnMbnfEOZuPLn2m
NUGzhVP7hgA65QCJ37rEo9HonZ6/3msz1Bt8U2TtXBSr7ReorE2yTuGxz0LanHDxkUnT6PP+UD+H
MTr9/V41tM415SF+atWDLGBnMVJ9zhuQ0sgeQGc4lwHqgJlRISPvoX+SWQcZe94zQSOAk+XDMTHf
hbTveBDvw27DQkyKQJlgLK9fUYTapj3DHzhMVnLqxaCjLSkPn15z5LhmJLzzlkMq1u2HXr7oSpbE
23OYDXol2IOWmOnRONy8LRBGmavRxHY3HCgbk2vBURi2l3bALIhepGcNtA6yeVK24kQ0hD+WNZaB
Ta42KvODf+u5RLcj4OLuTTiPu+wNshiyM3VelPWP7qG18LI68iE1eCnmx8743TEOg/LA9PyWdDIf
WTcsoFV5rbZYTAEdXh3eO57I9ANgMDq9zjvNEhrpXrMU+XaKN+zrkVj+es9UjsA2cw49ft/1SCLN
ncl5yRyEEbC2lf/RPK6Cm2Xboryx6PxEh7Mleh219yM3NADQfNQXy2rC+Ko+dU8TV4ZjmEjYXIYU
kfjxa/BeCf2MmYw1FvlpoAIn+2u/KvFnALoWHvwZEM797fok/GD5cmTe4ItRQ+LXwIfMRDRpImCt
pqSg136FVKFCA6w+EFMbncGIthST5SVS3AoWkT2Mp9bWy2dphYO5yYzgsCQ5U6LRzW0WDwxAMGNc
QwwfJ1ulz6q7lGBFprTp54QpGze7bQdfe4x2IYiGHnynTfiZQhq7LRmC6/WMBzRHowoGlLIrJyWF
VzOcq1NpF04hBLNF8OTaaQtSkfvxswZ7aQbV2CX4R+x8hdImfPo/ehskMkMq+TKTWkwnZ0WYjmbH
iHkF65QL4IamUMkGx35kADU4oihuwm8q5nUdAdbsUVBpWQXcxYPpGQUpClZUqsUPDwvjRBXpXQ9N
na96BtgVMPiMCXKzpsVHmniPHCHv4ZfzSuXxTgHIWWAUa/gAMvX9sPyGE3K1pQBHi8m2Z6SC35vO
UPh+eG2w8G6e1mS3FUFNCZU6VsbfI80uVqQ2MIyHJXykHvkrW1QpURRnXpt0ocDa9lazUPDLW/iM
+Sl565JxliOjnFimFOnWXbcE2t6tqOEFq84D9kaNgW5MCqcQlg6itgtDO4JyHn3pJG43eRYXMrmf
BEAvO+5pTVI+qLiYFV946bMxgUdEV+OQDtS6YIKaIpxBb4zTQ45bq/5cpD1L2ZSc5HGv863iIjDz
N/DCVsPNC0l9ZwpeScUDOrydM+2B6y+kf3ZdFkVM3tZg8vgTmhVuBmQqDYA1UTLsXked+YjuxA4c
6CsoCy3JZwOJicodFpOMCJo2KIyDkrkNDXDoJyI5tRXK8xhXGZvp/CIeI7dMKC5y73nsSBa9XNT1
dKXYOIyVFJykPzQkLccFdrxNJtjCLwOf9xGKqwZKFGJBvWfzXVdspfzuJ3NsRzn8Pc7RjFHjo327
Nuqq2kf28HMSuTsIl7Al2fPnlnMPauP9Ap1IziE5qFIiQPtMqq+v0FIrknRMqTHWiACiVcPYOJSz
FlWaHhK1ZyzI2MFWR1A87dnQ4ZQq/9jX2UARQ0ApVdBFjsmrMjFZ3JjjimMOMw580F9TyFDcSomN
xATRBB/Yh5NmH7DoGzdiFtqH7j7iEdHShQvAvYQdhIIMTogFKvF88O4NmHQIf49XEZzPOjd9W8yr
oJX00SCXDBT08XwE5kZCD6Y4nfxXijaJy9Zq3342oGj6nFU/CP+D0AfPEzsAPR770zVJcOX3wSDo
bdXh7lhdYzR2dClMQX8gmSArLNvmbMUo25zq5AgY+NAok6sdess0CIpffuSwAHDNH5WPciVvZasB
Dymdq9NMJV0oQXaUngnyEBp7a0basiq4UQ23x6yABSUaR2BJDse5ZckDenQ2Gfy/6WLE8yrMjOk2
ksWk5+qDTQLZhfL/eBqb6fAhV6/JBvsn1lFw31WUUer+HzuUqL469VDPqhSmsHX1a/Bf3aNweukJ
ySFN/1kFGwD/bl1DLMbNtOw9to9TlBGiI7C73NuEM7NQBQ2tE+ngOK94mVbuazw+zjy5JhCr42Cm
Ody6SMuhG9ZxDF77iTP7fPBvZmryJCXbLXFSI2uT1hTCe97NqDV7y2/Mm27Ry3BA/YZd1pN5RLqm
0IA/7Gf5DqBcv8CepFtxySQwp54/q7Eohubz/dyfV0L/vgqUdmBwq27RV+UozbsXuEmQqWzpoSlC
V7PK+DL+csJ9jGYPVFo2FSwNat6PZDC7Lb1BgzA844NEf8+QMWLTQTeIWcQbvXwtcfFZi4lnkBOE
X937TZ6W3rfSeNqHSSk+nBe56Z3Ag/LGbUSYjscliBbD5e6vWyWkOcIQpGPoaeq4lNyjKqGzBA1c
mhirRxZ2XOsh8SECkonW0ZDRufiprZFXiFcANKP7zGgb0RNzv2xznXVeGbllDNKpLUI7LQR4GuYL
1X6Xo+MG2jR/QSaOssw8p7z0Hb3S4BK9hA4amEscbmid15vT5RlbDzAef4NDP0lzfSyiGu85h3Mi
pAfsN1+tyKgPHeO2kCqfXuyFDm9pAL4ewule9cApSL7aFb1X2+1ypE6HlCdB/Xzyc3PwbIVSghEX
choyRaXUXi4xG2Wvhh7zKTeuqHGi81Jrml312FXJmCq/41/YxAW2M6fyl6BGdxYJTv7bAPhyvigz
NlBEaQOwnuYCkGiGeTbdCdUr2CO+dKaGG/iqyFJpHeWSJpqrqCXoITFz1Z5R01U/l0nCJtUwq282
JBHY3Zozmu/wOMkQ7xIXXuXT9o1nuSOU17NyAhd+x9+3exhrt6tNBD+4pVA6FYTloQYFz7p5nmuF
JS2uptHwulyOqi65yuHsurNTAy6YqrvvRZeXEjKmfaVX5p/RjFxKqvpbIQ2NoHWl+lS/yzIQhjOe
O5lMJoIV6U2TUrOJ2wYpwK6VJ5k7NjonUSjGEtJPcz3hNJ7xfRrqZPVgI4evTqz3nDunfIfPfgku
NFi28/ABDnVIZKRwa29RulWMNHK8X6bM/ApHkVH9s/T2X64isANr/SrpiuwQeyjc2eSLPfcIX94F
kDuPkEj5YaUItTHLwm9Uw1M7x9IkCIAK531lV6IxorPqInquAoIJBiLKvctqF2e14JYgAu6lsvn1
onn6LG8Ol6/gUUiiOs6O21hw8OSKKbT0btyzmQXuPnHzTLXuZcjB9RMnMxzlKGaBR0bzu6Vonl89
9cX3mDk2uGx0fsRBsIA7U7zK//rmPGQOCCPy27W36NOtguyFUPhfx3Sob7ZKmt/q8RcwRP+0i98c
q5AVFWqnmjP8OgMwbSITH1QPlCB3FjfnIqj7TLHyYVjdV1Sm0iMimi4JNy3X3R2EKNLvXxo4iI9e
A8elAJzAcZ0Y9IZC29LM21a5I9vGHOdXEEvVYe5WN53W3kAnxWbFs3RCyiyicCKtXFD8iGT9VB5C
OuJTJ6apbGAkDPXjH54FESNeOZYD3LoYOFkUnSWOxumeXKH31uOKtkJN/GgsM/Rg/WkiYIyxm7RP
mRSrHpiQYmCNIZSFbnRKLLlSEFMQR2fJDIo9Y3PTDOqbDV77XuEBihqqc69BDEj2JEzMJPDlXepm
qcJJESg+WcutrULH3/FSXCL3ghcG1LVDu/+YGdGrBsIsybcNz/PZ+rrDCpfAGGLhXX9N/KvIQcJq
+t6sz3sVakFk91hFnK2CBV+XgRJspg1pyHsjMR57+1Jdyqppt9y9340e1gPJVDL9PHVcOsQrTa8R
CkgI1I8OD6JjEb0xNqhU9Lz4X3S2XJLu3111QvCft02I5ORzTzSqGs9BbLKVklVpg4RMdF7XTx7y
f2UJaD3bQCO0m3D2C+EH/tjv80wb3nYRY7RJEqHsCJ5BiTy3wQBUaXAtCI8fq3MHfnxCzzPGsV/O
pIHhIdUjPBeUNdMKg1KDQfZBm1ISMECMbQbkDq+stACxv6AkyGAxQdLJQ7QlZqwymbv69XB0yyYU
dgNzXuzkXigaPmLA7C7sjFOzU2C/LKRKZ9Yhng1ViJmHNcuvQ3hGMhXQS/Nnh0NpW89FxSmdjCpw
4eJPumPDlzrNYgTinWZjmOkZZ+uXvyCm8L39NTrlwO731Rf+VSCG8MO6+CmTyJyaNtQpugmby08/
+Yt8Rmot0kyCpd1VEMwHwgDRCxEUaPCSbIvz2wp+9x2L2lojRsBa0F1A2HV9HPrPZtH7QO+elijM
7mb7Wjq4TNkl4Sh46/hAqRHYob9k+wUBUdtJKAtBGgH2f95jx31sRGnjG4xbkbaGcYo0kJh6p9qm
PvyACtOEXZSj8mUTU4TIjW3Ks7mwSEWc+DMoZ1lYXLLHDwt3aMVHK36xlp1SjiIJl80+jkMWxtZg
8b/h+ECuqq8XFxITsda51dk4Az9XfYT3IuYffxqABYHEhNc3E+/NBkhPgikRuzClBnizT1DP01cs
kLlVkvP9oBp+eIPshwp2FOJd1d2NxlwgoJCrAFc0a4gj2OtP+wbRhmJzThn7bs9xTKw5MGGEYoJQ
4Re478AYzHLQVVBsGKiakDcJpY1/CEqPToF+Qo5Jg1zRyt/A4leCzLOJYnAI3iOts1zqwAaETdrV
yWxKqYYXcRITyYzHV1uLPqbg0EhLDARB02/yADdMjSr97WqWt6yO5Z6dQuTKWeuRgqpDptevDTiF
Ed0sTDaqq5ATAYXpKZn9Cdui083q6AOJQ/19fpcbPqdp8U9C7tFRcNAILxQU54JuuLlFd3sV/Eb4
yOTy2IgTbh9rWUYR3tZ9nzDY8+SVsiOv5qOj79nh1XB9ruQheBzpNZuZ1gTjR0TzrgGZp8AR8p9U
/EKUywRYD/BOpYdrjScr7ppvs78x6bPqWeHod0HBGiiAJ5zxoQbKB5JXt6ecIYOskxF3ZeUduJkj
oKs/REyEvWnEnhMU/e4jOrFJrSqrPIV8x4xTfU/DT7DTzBhXEvvxesuKBahXkul3qYbcw5mAI8iO
Qp//qMqNVIZX1tdYQUKiY4/eKCFQC5cJfJ3vYjRWskICEvyBybak78IgZ46W4QT7DlscsGJ/OOfA
w/z1NMIioDknI/hXq3vRUGSXbN3lmWUoUFkp2hJ6vZdJH/9EOZdkoZleUl24NF0a3iVtni/+013S
7nwZ1GkKzy2GcOEmWUKz+D0AROUNplI9xPkJUcM2USs5QU35gTLsV2MVO4BJgV5vgXONUyOvJHkz
2TDCG96ILCSOEkT3scl0NreZaBwicBr6XjYImaPsWoKCfLHAx8ZnnTQeYefBuwTUk9zei4pXZFE0
rj5u3sLux4oC6TS+PpXcgxw4LlTnHbMbIKxxO/QEuPfjLAcSGVpMiCfGMLQrk1qpHnJzHJPHcN9B
phre0DO1T3wa6aef4lCNsj8TSsKnywarOD2qkndxeOBMwUO8ZqoEZ1mymuq3Kn/RXvOjHP/9CYv0
7sxnsX3qnMN7n3SoZ/HcN3XScxcwA/FvJBeDAUzT1nMMxnuuOdWRffECdM/homeWsgxy7U2EwQ/z
zsHyIwBKNqLyohxODBA+B4JPwnDkth+HZ3E2D2GD7ArjV18Awrm+u5qtQ2+w2SlhwK/JG8tbIFsh
it4PmF3kIMzHf+a5mBGj6t5Vpa+5nPkUeZo/zCmpOPzCgSJ8UDSKsVMcN2HWdqVuQBUJ3gK0OR82
fe7K7ARh9AwcgU05OpbcujG4FxmaCHwpphpAVtIQ5ccm8unnkcTq3aREp7DYvdbO+GHdTPf4mHDj
P143QaBhmRqVXRhtivAvUAu0BvwDsctP5thEUwsODqcvbsBa1KpWljqdwuKxDudASMtsgotFRc2i
Yb5XKlvBjrMVfQKVKdQy+vlj4GE+/zQ5UZ8QQwN/mSxlf7SoZHSN3FNDOcQb6QUM3/5pDu86s5eh
Dk/zQQunP63+dV98do0pccblYyJkgZeLr0LZ9OdOls4ekiwn54tmT6SIrxM6CRthUZ390QQgxped
RXFCWzNzd77iQTlRHTEMfLsSMee7VkvI+Jp9X/55Tj/eC4ki1q55/aHNAOYyuQeGB8W7FJeXgJ62
+XM75tku75fZWim4jfh5qKPOBaKg5OlziwjZjI7DBenpRNfbP7689mkej/UOxsrLq1ImZs48r2+T
AXdahL3cwqTi722yGbixpK4pjuSQtp62mVvYZovagTaRDRiIae4G/XN0wRLPaWLFo9ZvGexBCWO0
bC4pVZ6U8zUDScTLB7r63hCtvM58f4jYHjk4NStC6eYdA6Opa31xa2aHQV5KKx9d6Abg6jMVhCFt
Dvp1j8WeSn3UR376JetQTTpwM5Oo5Gq+l7tmUuK7ERvfqOClNqPwfdnZNtYup/a90HBZuhQ5DuoP
A2J/uWQn9uK30BKwXqKtmMAb/AdyOrIVj+KC/lbP9j0aNnpzWXz5NLYozS6HyBph9ys2spiGY2q2
3rJCDarCUzXynGtaTOXnkdBEcmtUqX9CBjBFbxiBwQsbGivzT5ej7n9pyhORa2YwKiDBeNKY/nu7
BF7GqbVY8rEZCva9zYqE9gu9g1LHG/ulT7yN108FAGMKw0n6B61kmE4PW/NvJWsSTG9T6a5TW07f
YDRauOCyJQaUvaHBR5lh5H4HuIXiKGZM70kkxbHJ6buhBvxzeJevfPlTvPt5XLvpZO1GSvqxETiV
0RZ2GdAFnH50GnzdUXLxFsBDuPdPbvoIh91z6FXcZVV4Ph1PNVDfpJGRZ7Gq128pRIHhvjsxsXSI
dzMbdoyW64rhgSB94GUVI0dE5DdQ9nxKsgWZ8t08L6DGJ8cEUK3bxfX15fQHstAEl5FKirOfAz8y
kkInnpZ9JY40VdODCfvITXJb0d4Twrg/bGRbJ9CKqT4iIhPq+6yd4TKya3sbXASGWen9mJhncrlP
HQggTDYyd2k/IMzpyNKwGyebpSVfBd2I/ITB2KvKvibL7ypvomn9vRPJkabTDMCjiGicrbD/f/6v
TUypYHOIS3E7uZOEUjuCHwMHNzJBe+8uzvngbVkfwzTHu9cTYmP7x1eS7go6AVs/7wXy6KsOv6qF
36UIsALOgVS+rPFP/Vsj/AlSPh+zfm1UslxGr+tIBza1avGHVT4wGnd8ErR5vzp2/2q+gVF88idj
aWp0nH3wpIevwd8UAtclOVa3Fwah4OX1LZeBvWjL9H3p/hXSp64y3FuXMSWqwtus6YHE6qOvTisZ
axGh8NLBq6KzuNNT+R7cwnOvNsrczXAJTEHCSY8sUlFEIQaUAeQ9Hi7/feJkI+F3Y8uECcYxFZzG
tOdTsDCXy/rYN2IlOBPIsjrF6Eg+th/v1DYatwqGXpO3H0/x41QJHTtjgyDNQwAxD8a1KxWpZGJK
pY5OB8JtWHYwvNT4Ss/nmYF7AX3BND193hXe9k1CzY3CZshxZsCyZN9b6qLrzRadJy93BO9nTkRw
+3DMiTyeY4KVxbvQIuMUivgRCiA+mZA+1jAnYVlGejWIJvniXc8NT7BcZDPJpXbjjdinRrue+uX9
4phZrd7NOKQnaFq7z+OxzFGarhF/6cr9QN/Svca3xXfENSOZG62M1wBbIdB2jqKL59Wapr8k9ENV
xG9/0gbKSE6tcBNd4n7KYtMXadnmp89/YMd1ZPtM3xwblLQOAVhW03GYgJwxmea+LtzDJXKdTfWG
AF6SD8OdPlg0z1nqTZGjgLUauAKzI5X7kVPjUPi4sF4wz1cW9CS1WI3KnASN3nPe5XSen1ni3TOW
7BWp52HJ2k9Fiauz3IeeYTkfyBZs/oD/IfTTAkgTeX6mltKIltX9zYNhB2qgP/BBvQl7dleBaXMR
tzbhgQZFM2KmP8Qv9s2OTGpcDgh0UW/3iiRGu18rkDDEEZYMzsYCbqtIVsv/1DrriXqYsRGTv70l
pvz/leZ/hOYwdoalaAhHV13Lzobdt8SDwf4P+tiItjfrh9p6PMx3LuIFTMNwm8w11NYysYEKU6l0
sR04gayMd/JKrd8SLBRMBXTC87SM8JBoMGnbBf6gBhuUrhsTEPWfmZIb9bcRWjigt78D+HcZ3QNq
twW7gM74UnZpdsV2nG8S3jb03n6oHxciGKnDTmCkZ6cqZvEttlPRegZ1uPj3neWmrAbcUut0TU/o
obZUsRyCaL3jjnaygvfeDWCSlVeGJmmNvs4E++aXNAAECx0gKy/uDe5svdrU01pzfyEZUEiH5g1w
ooK6YmGPRvwO1JXWcq3zOYl5HKKsm+x/MTICsQFRgHbg+NL7jh1xPWG+HqRwrpVtWtKuE6xSCD6S
u0AXU/ftDp+CPKXLElsuBrwwU8ChRTO+lD7Od5aAbQ==
`protect end_protected
