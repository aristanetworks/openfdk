--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   duplicate
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
UQgiO5qUwYsz3TKk4TWvi9ykX1RHywZKoa2b5yu/F32iV7mAeC5/6Qz+UFjNhnRMcN6RGMUa4HT+
PYdSFtcXCWe5tUZNYuBT7l+PzYswX6gAmBMVyEFzUygNhFPXjek6lBEAbTY75gMDaUOxxP0kcWV2
SakvTHbEWY6FfbMXQ0h91ae6Ow/ZqeUR+OEi3Ub5tkKAxo/CYrS6+WqMOyrnXwgP6gtohQONhAxF
mEHMJquBP17CTjgp5KLNzhZ2zU17+gnX/BegrYxKOMBBrjODwi7vcKAj1wYRbJq46ALLPWZVTT4u
7TJRY9wb3gcs6jKHOyisB1V8vJrm/4dZrjgy8g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="pTFMMhF1twZmyB70sTUvOogqDRfugSdbKSjrFEAnfwg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
Sk4TqwdXC4zj0yygTcye1GvJkLAFPTiFdQJr3rtk5fAaTb/i6I9jrw+a2Dw7kB2ZRT1G9B0FVonh
fTqlpFqP3/RvalcvJccsTILahrxFh3K9mgxEVbzeZd2wPe8gZdz+bXxAdSm0+xEj+svall21LckV
CtGoLTD5LoDkaK2vm0Wj79CTH5VzuaSTDHiKQd0Xm1BuRLElIzSoQ3Jyd6nhYTtUblLNZT6MCzUr
VqbXBDWNq4lU+iC9vOdqU8UUa/8e3NnizpxVMfIyB7ZmD1eNsfh9PfL2xIZKWI97Ng2hu2pbJud7
S2ZGjJIRm9/5RhKNTqDPM+/37f2C3dxEBncU3Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="fj4KIBOwIQ+/UgLUWmPLCRcIQ9mW1Yv6/0yBO+feWHk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22704)
`protect data_block
GSXSShEiGGfgsNY+qNmlVmWkfzm1sO40OYmE8S2HZwuNzB5Falu1HBXT/KSCcW1dUwgFR/s0tx3R
oFNnYNR+sAsY2SbQ4ZW33NyonbHmwofzTctgYA3xs/dpWjM862PX3ORftMJuIw/UlVrPiw3UXdm2
LAXnCLZeQc0Ud6yuupub/kj6GcQ/dxxDNPBMTwSAl5tfxfITOMU2vfEQeaRW3LmSbgILXDvRbO04
MlXPm4Lz9IQwtpacO9/nTW8OMOSECjQcrNLQbgRw4F/JfQw0Mv1wMOrAq9bJ8xEYO+VHUHi0zP6C
l4QINJ1DBiDZSqze8uNxewMTjqW60m7ViX+5ZNvs9c+UrrM2OCHUTbxLgvCOKAFOZYC7jEqWGMRA
sjPQnBY1nQPEPj6+z7Mo3u2HLtern3xBiC6gXhYWqkVL0qZVKjMeaaAoCdWicPYYpALJn5448BzU
iIbjm7gyfcR6M4ApKbLkxcnA0zfZhitjDrBQ1b0gDmXJgF7LRQeGhrjx8LAXAlDtflI1w7Ie61Ui
hjdetexZithNyljAaTkg07q9OFzPDEotffWCQIcApinbecd2TsHE3icSsKD4f/jGPjgWzs4F5KCL
pSNNv1zi1d25tD2MIcJGHFZdTrOqPkxWOTBUL6Xj5kvHQkxK0IU7ugaNxXh8ja0ew7Mk4t4GXhIJ
vfa69i2uzlZ9qbhQfUhU14EGT6XbBefusydruW2Wm0iTgkpJOb1Vkw2nwz3fAyF2uIiz+c3dJHB0
wQX0QqlrJZ8U+MHgLIPgaWKI06VPhoDTN8JtVO/HFiyBhplr4wAqSLSEVkKe0pxpdjwLX8xZQdaA
8e9iGCi3cAOnXz9Bt5kDZL+irA/6dvvpk6f1f9eF5szSay1AGAKMDRKRMfyUlfkCkQA7TKpDyqiR
5EveBDWu2mxx16sisYegDSGFB5pO6jpgG5TQm/Mi3ngXdcktLI6Lkbof7092i2dphnPwPBiJi07e
Rd4nti93T/AkyE00vOL9PPNylywp4mQE+wRCl4n5n/9pgU9QQPXnOS4R6ii5Px5xtjaKlU+rngGP
rOe4XBpoIOOQLy7ibB77uxwEsRrkPv+y8Ma+HOOP4K7aViXCea5Nfbh3ZoMGplwjRRkHtIBlUxAG
rLZZUBjex9tUnA7v3+mwTk5BXWrnurVM5UG+q9zrio3mIMM1tTLpzIV1iwPrDfzJPnOTCMBZb5A5
ASL40/f4Z6+c8XuC3MrbUPTmQIefgQeX3PU1prL9HGfWa3OK4JY1ofyOEAO7ioYV3C2izfsyW232
3B7sKDXFa5rKEQzPA4yNKObTwUIdzB5GEohMAUFlzUjamRlb5krXX1JcAjEmUj+OR3DD/p55EgCL
Sq0i82vsffbNQIEu36Ot66VmXgp8T86PRejPmX6l9gOx78TGT/rxd+CStUdoQz0vv9GJg2WzWJIk
SXpFJIMuATIoe1RE0c1Je8f/d2MS5IOuKh//kCz1R5Yve2HRFoCyeJH4Sk9uvkQ7B5Tpylyp/kUi
Inz5sv+djPhW1z/rJyu+p3fAHA6R3ZctFewO0eA6iL9Why5Dvpne5DZd3Vgql6n2Ki1rFcxRHG/A
0xO2qduLYFhhohTT79FJyoIsbhuN4I44YZ+LRhsJ29kAqCBj9fcIgogG3EOd1mDfnGy3MxZtSigB
JvzQmePffXrEokXOQt4aVIqex8tIiblWdY1p4LIn4KGBTYO4m8O3jnUJUiz6zd+UsHwxPG4VRI8u
LaAWRlHMQzSSUgta7OIYxXxdbQ5sRlx1qIy0d7ZxBxhcltc3lB7a5LyZHikZbIFMj2+ZmggbMr43
EpXtrbDJJFhrOMKLUPMvtMF9HBIka9X6LEoc3zTmhH82Mt+o+ZAy9lpaxPoNvd5CeozO1Tt2wFDS
GbXJyPTHVEucQWl3sYNiJGw8rlbRk3Mi4UAzobgPdBYbY+22lCYxYx7UWZxaYeSwHToTiIiCfp6P
mnohJ9lrYiUh8edte95XjN+Q/YnhBUnjw8G+pqVbOjDLlM24niBJPheBFcMSlXYWlHVJhQgqmHsJ
A58m6x9GHWwoHNS6H7ixiqPnkIG/f8a3Z0m6Tp1e8jbPzziWs7xOAu2E52Xo2f1v28X12x4mvxI2
pmrdUpruTclgFgHr5Hve+gH2BZ1jZAtE0k4Legz24GW1f62ztUv7NdCMF6b9HSttvxQ5BlXYvtMm
J3ke78p0ByYaHqcmj1IkQ1qP4kTqoA/EHfYX+fKyEdAN2IVQvl0VDTK77lYvHYjVoz0qlXd9Ck1V
aZL7HYPXzAk44VZ4YqCPwoPVrM6N4XfRYC2DFNZ0Xa87JvJu7E40NKtmQKW0SufKms497zKke5QS
Cvo04lGDKgtF14hodpwxjTEzefB88qwSlPViB2ir5uVL7qqx3PjNh/78en8tB/O0BqKnZevqgPjZ
RlnFp55VywCnGNMfiRbT4Au4F9cx2Zf+CNW9t9jjMbiqIORkyZBjHbqoDgQhoI5NwEbAyreSKl92
IPhwwex9KrlkB8wov0UOR9PFj+XOfPOLdzUQLFF8COs82IB2L9bZD58DICCDq0dKbtv50zKahw3l
MNPZxm/K0RvQIB+p36BCnaD69T55SvubbxJMuGsHXhPsBvK/UlglbpzB11eMcSYWGwG86U4tYHGL
VhefOX8cVM/ROxmZDSqjZWGKTsAKk0K3x+N9b+KSUfmHC+gFp6DtRHIZeXZV0nDU7HqVSURUjxiq
5KGCTfvVjWd52Aw88GlfQpT6IIof6qxrCkIPcG8HxevdNHwuQihcYTkA2J7cbuwFyGHEttPoc7pR
OC0UVVeBtW3MfqmeZv9DHPNNMKFbu6WXYhwchdOaooNTGxzZAdn15NtCcsNaNKKNCIlIikVDQMeu
kJRAFIgi4eQjPUukPGDACU5WyKc9JaW6cwv6TjT93js5qhXQBL/rPIzqiSV0EsmAf1yLzK0fy5mQ
gFZSgV7agQWBYQPLVbGy3zDIY8FpL4e25fpvQWQQzB/d6MaxSn5yz2zCaF5LrwrZ70nL0Z1xmxEK
YWiPpttbNwl6eE/etT/YWQX4z1hCr4Qj8369355u8fawQ1JZgJZhtADzwa7Qdawh+eNU/Bb+GzSG
cpMzsRRhyj082FJQwDohI+RfEz/DPcB3K+zL1xKzxnluXZ3L9IeJSowTTFjaoYH8cEyOcSA4ESe8
tyEh6qLwD1YMaV5xFYQ0vV8pVz8BTIabahsiHOtr66SrCSM3Cb3rdlyCly+fP7F0nf4+Bwqd4nlJ
awwdkZYsOT59ff/szDm/SbDwoKMPss6c+DX2N9rOffoHB0+EHrmxVDQsRU2p1NqIwdPQ80d+lszO
beAmGRHGOBMalAzlNziUALb+SjHE9XkUgsLv8y+Klctu1P4llv3I0956ZJN1HTnB/7iHWl3fAqi0
pZogbG6jo4FvPaJ9Wl9oFlSHnIyY4JLBEQN3ccTQcZ5yPqkvn1BG/8A5w7UnUOPHkiUiEDywRdld
NItEH+Q4rAqoj2fMuhYxukdvcDCza3Mi6IRE3k2ohkWB3pmw8ecxuhxsUkXUe2LS1spz/HhjYyhC
6T+NU3L+huj/Opx2KKPKms8NOoWwOoou/duRKtuGJH2POUO8J0ig7ZbiW4uFtqH4n1pQJvtgme7E
YC98YM/gtcEv/TYXG382mR5AcszCxF3LhL+k9DPXqNCbTisTnvEMYLm8WoSb/H+K4ev3Xy3NeMYl
+OORp99JAuTz2JtyOrUgD6wA3a8QiSBQm2itEzLo9dniej4+Yvupig2x2dUXzZFW8hjKO9+umIVY
aPbmGrRDqqbZCWi7u3S+bPE6Paf1dqtbsqTwI6ajjwloMIEiWN4AF/lg0bA4kF/m+3X1Dq3Fmjcv
UujAmBkn5FqWtxcG+owL2gjJh5uObKyDA8mfHA81tIo9oOb8F+F7jzE/ZVPCmahl/6Jeo9PQDLsT
CAnHw3r88aFqwpRDGp1kt6FWVPhHsRbFjv/8r0PUzVFDHUadSKKGbRcLWoCn8ro1xMrfVS3OU9ax
Wjm2Y+slNOjk2eHBE8mkwNjwYWKzs/EK7S/zev47C60/nsuikijJwTkAtidY9D7gxfmiJ5oa4q5S
V93eaa7uEgYHioIQQaXA/MElLEYe4ZrdSqyx1Lu3x4VPPnDf3klj09tN3PLhEJZVEya2nOZXDFID
m4x+/Yf/4zaMc0hwH7D6OaBBHb74dlkEAqw5EgV8+64q7o1dhNbZkMjYwHEMO+gLxnF9tP64SNTa
TPMFYwdy0J+D5W1YrEjaKH/xH4HssBwOszpR9qmgaUT8W9EWJ4c4Y9Y8xG++7Yo4td/Pd+FB6D95
ix+2qN0uLxLLhlQuhk4ZZ3NZ8R6oNHr7JjnUNuGrKLnKaZX8xibheBouq3d4QzjcaxWzjT/cIH62
EqwnsIDBwBZCQ98OjX6CpiE/qKz7MwnG9sArqwb46L092j5Vori/wSLimlAHI3kMmdkJWi2xGrhH
MuH1HMvQYtAYTrMlyKdbiQYKsPH2Ztg4I70u5ZkTbuOFqfMgPvnjxGLwa8vuRiH3ZOw+bbK8XV4M
5EYRiEMIe0Kjrh/i6ASEOETNmBDeHzCA7d528Add0PYsPoihiR6EqB0YJOkZfvfp/grewGkx3low
HnbG0unFiw10WaX3/eAUEaKThaZ9cVfMbLwChyPbzheg/C4BE5Q2EjKFonkBmN5K22ye57oaV1Fm
fey2chy0PT3BwCyy32HM/Qz+lh67eLtpicsTbU8wfwiFDFHeciJ2K20H3hTO23K3ao2R2um2iEv5
wo8l39Yw2Ws8d6nbrg48Ejy4ZDNAniNvQFeXA9G/yiOd+q+hJ4M1JdVx2HyBVEXWMhsBJFA+GWs4
5GG5qeQdS0Q7PdNXEQh7q0BYwmI/5Bhb6StJQ5DWFUz7KWMacmMRyI5eSD7DBaA03JSgVWcsk6JG
ZYneR4PON9AvNKAV2JL1rmUdWWf5hhYUhpHcwmUnC2szHNsWyIAc5UWjjg6n+aJUJ9+by6tU/RyJ
XtqtlbhGCIO7rQFUDfDnEMDrUgLzGuvefc7BfXVm1uUhqB+RBRxbm3N+tYKMblZUj17hgo1FrnX6
1T7EPFI1fOPcc2FUqZBBYiyaq60il4SF+11nfZog8U/j8y18KSpzTZPXuUU0D5vyN8hRhZ3XE8F/
P+199hnYdBefPjrREQyE0I2wbIqNJR52BUmXq/lEUwRxquQBJhbxYSDRdtbrXc7l8DIQCQnK8kbc
efDQYZrH4OGQfTBGJBgUURx+Y6dQHIynQI0VeeWaeLNJu4YeiF953hpUcItHkBu1cEs4CMmfvPux
tzUqOH3O2xL+vdmHfd5WbYaDs6eTZs/EYHDi0Mcox/jsnnshc4wUjQupkO1hzgUUVTHofjzYevPu
a2wSpa3txj4pb+ZI7wUtAomWZq5MneIHNCF4DTm2dg+CMXwIRWgyq2ajHwEOXP4XOIxKjBiHqeeY
6VumohE/P96+nW0Xopyx6hp5+h/EfG0MPZlSwbQkKwHj+xL4QuRDKmVvdxWfzIx+2mRNEjvUsT7P
0Oz1oiY5HDV6AK4WZCHviObTMmo3SqLsQBVTsLeqCNTbHlZZ1Z7OQNsCo7jQPt1aLzVPmjpPYm9w
j/KWoZcvuo4eZ/63qrY403elB4YYb2MVBZAoCZDpM9S082Wv12yHi/svKUWy6RJNNYI5w3SsJiyX
d+5AX+yOFccu+gXRG00PGcoeEtXEHHtUirSDJj6KtzD9pbnzcyd9gGGydc18KEMhqkH5h7aT9NoD
ptfdhO6nF4MFD7Mi9yd/C8BxRyOMwfsarS+tQuDC5tBZb66i9iRh1Z4KPpsJp2msrE0mSo3SwG83
rgKlZo+tyzFsWiRhhb1+ul8PK8elADFztIzoK1SGinepIgsq6MXp4hGc4hF//2JiscTJhUy17EyM
T66tycBWJu5gF64t6NqIBULJ+oKntp7YVuywcWZpI01mmKwFpepL3M5hUbhbl0fHXL6SPbklGV09
LPTyq3kC6l2sngdX4KlG/m9uv868n5XuypcKM8qBM0jqvltdXsjx0rh0cliwR8HGmaNNyDTxul90
90uG7RUxjxjhrTD4wLLOKs1Ar2uoRZGXasd9SfuZ/jsJ632srfxKVtQn00XcPxdcKXmHSZ4vVa+s
NEnS4wJ02VeJYe0fYZIIyLTlu49m9dUhHjN42bWU4R+ysvkcmLQamwop+Cyhvo5TlY1h1+Sc+5c8
lvx8wiqmvKL9NSGSHSU2H7WtwIDNpMu9nbu1Eti6QDDBqRF8nFPYoXmKx7XDwFl+/4r+6E6brO/X
lwj3GQZfVGAWVYy+Nv+US7D1loQrnPYethRuU/TqBwDBupMrzMC9P2I7n5hvK9o80djgaAjvazDS
V8aR60GM5NWl8kDwiHh1ZhmczVC7vUWAO+iR3ACMWsLDj6nCC0cv8kEgVQdGdCKuP0BDvCYmMmjI
IzdPmOntuWzuFqCtXafpFhVz2nn6PWm1vg7R3J+2Bx+CZP1CDgCEbKN28KW6bOg4xCV0tyXDzmsX
UdUGZ5XfJfmRxaVyqaFYFrFPZ2FX46sUi/vIQgWOJrhmkExRwQh/CDd5HlJ7BsgKWWh7Tm0zkIRi
cp5oITlHiD1nH8x0xBvGCDrpDUKXfYSVWfHDus1o0ctFMDhk+SWVNcUdco0H9zgRNs6nNwiYaIGj
u+/vsXnAQ7EnuhDlQ0JEuvV0GMdGgTDp6BLKY7DygfiMAD9hfPpBoxEKzjwD1NaD83TK/X3cWC7H
PYxQoCY8l+25zlL9wgUci4e5JMAPafESNsztmDRLldpAxKMqzNBPn/MVcUB7bG2LbB/pynvKZCaW
82GujEyVXaX9I1H+2v5aADM7ys1PPPaFD+RaQfGfDRJckbLkzbOJxk5ipgOawX6pDWf3P/1tftNk
Ke+H9J5vznDkYedrJfOfKNUepbAcjjwqdao9/gbpeGAkRzSxu2l8TPMx+xdXkO5vhZhLshx7feS2
iZ2epzM6j+FHw8wFBhCkQCFVlhk7fU8YGFp2+ZQFhyMtb8TuGYsVATZ3uQuPl4S5pdr6rQ9yCdCf
8kgz7Uk5DbmlD2QTWWLHRF3fztCxabN38bHEL0mUHaOPGvOkVLsHWDyo+HXVGc+QhbNv5jYAiARc
i8I+EisvcLShDmouyHvb8+aEMLISxygXFnKq4MWOzEwAMEAcSpSpoF1s9mo7D5OdmcOXBAmeTFIo
RF4UY4JdFDRnWL9gFE9/D3LkJZjuZn+5pjqlMzynrs5/deqzNi+iOAipHHZgi8lM7Lg/nkkaasTR
/8mzTBwkwxURXKnJvJ1HWS0azC7mtQh6rFAXKkXoVcv1dzLqvmqgLy2jY/z2+cI56koI2LDPCMyn
MCHv6/XZNTByDrhzvtTDkcOQkuBwwd/gz7GppI665eMGYckuzrK/ZjIFuQEHz9sL5beZBBqAb4ky
5ZULeE8m8JcI26ZLumuX9KBwlgDMhm8wAELK2qG3Xj3ZMgT7x8Puc9eHlx1Xk7yFTWjT2OIwzd9L
LaLYB4k3r5apsQMg+HjHLPkkC/5kgikL3/WMlFI3cFZ1LJCsU6hgczgljiMnRzwkYrgn7qZ3u7uI
hlKHJrgAHeH+KjrAmnDOaoptY5BrkDoC2e53XDrhKeoy7M5ubYamT0ObGcvLcmLC6SqaOgDwzMmd
jDvqb6sttN2bTEfkhl+5Sa83L2R3IwVoqVXG00y3NB+Q3NEtZShVI2qcqKvncEVcnAnEbuyn0XCR
UF054w+vhad6HqWkCxhuXBf95kwg988tdkb+xMATzKsZ/S+moFQD3w6qyqYIFcsG7zf7kAn6cid6
/sbdgCyJIeUKZp3evxw+oJJ9MBXOqtjjCTtRxea7DkbCDDerahicUkwvkKN+f87UwxlQx+hF6Ivp
UvHvKClJo8W5Np3MZnMtZWjwcu++CozOKGCP9BEiolLTJhcayfJEf9Yk/ikWESlEnURjUAq70qJZ
b7I0OrRMX+y4n3hT/nKOaem5MBWMTV0TsXrk75R3bfXKhxpy4fCizWklw6wvT9PLN+GeJXFer35s
VkL77Yjijg7nZlG7UXiK+lJAyJ7U0MZjKK/cv4xlljtSVWtaKgBzkdbFFSpbUYQKwNST/TN2Fydp
E48d0RGvfv7F8lIT8fJ9o9fICTZPOaq8w3BFquKXvz+J+f4jcBuUgUIMoGct62HJBpyFI39khMAq
AB2KUM/Tc9ggTRC6+Q//i8SPouGm6u5lgw9mE9/82WV7wZeypikMxNNYnAbnwKZlIpVhm62CEh1P
cluvM2CB5cKfdMV77anoYNdUA5KMIlnluG17xt5D8SHc/PWrRcDO7S2ed02MUI9DMYBnwl8BK9CD
TPUi8v+EluV5FIZXAskeDIKC1OVdsbaCUu2XwXjGAD9eqGHuWxMENNz+cqf0d8YUkj/gLS90scDu
VbKpr8wxLgvjM19Z6kEltSVeCwaeMSweWKVleh7MBAAG3yJbL0zfej7T9/zkEMu30n54Qm16Yg3H
xuo57t9nhh3qPfAuByr1sQuJFJUaebzE73mNPzRXv/zKGcq0aFlHpo6Ygv6DupbInj0tnCzbUKAQ
ePOHJZNMjQgddERpEahQIbVAq5pa7uSLUCsDwmLL/ejzvOoen4kaHKvcUXR1pC/Xh6oLyIT0tijr
QSOqvS2T+lEgCCWE0rZjupMfd1TXqVryb3tdhQ1MOa8UX9/zY6p7dSQ8vUvOxga/Cvgci3WNCg5s
t3ZBuemj4FxEx/q3QHcD0W+if+Wr6wPLT9wxQ3pDnf1N2VCo62vrNQRzFYcvnWj0cWjopnYeGZTM
+cFDPcYOL4iEk/9kSm1EJWfbHebLgDdzPeccEz7uXkmIk+1gf+/P9CK/QZvYVAaIzBMoRwK8UUzB
8HgF0eJrqmspalbtSRVaMw0YIo0qwyU5YgJ71+LkB2zgIbUiMHNOrf+YJJMQY0i023LP3AMRjjvu
HcxGZkHQvkNng6c7/jbKPUo9W/tQTBWzeczPRxa6umQmJjTCEXfVZlh5s6YlNNZDXEXs3VRlWDIr
Qj/LeIIGNtZEm+BWLpRkYWl/KsKavS9lDBQ9DFeUM1qOlWjOYSTYbMIMamS6JGuN/yiLJgKBhYbt
i/vVEZrf2EL2oyOdo/rNLpOnwKAeUCzmykpqwYCWTyPZuwTYBtHpQFmL0b2ulkR1CS2D6s9kaUgm
nXxIzRUMi2euTWvhmN9QHPmYLC/waPmDazpzyOAHRDt7cyWJiuCHYnfx9E+NrUyRrywornmvZur8
AvxTsN8wIMq0IzoGVNpIhBzj9PM3ZHX1WGEU3NwlSAAYBMe8QUmAV6BbsY9j5hi3qEZ/STVVgs37
uVB/zhbdkcBDmV0tkCVutyePdnM1d8VJYd5IkMLTWS3VJKVctMR14MgkY1QkXRdx69MxQ3YtKivv
2pPuu4JL22w9yn5myeCnSGStjzxX0fsr/BNvUwbAHbzJ8WZlkSZPkl2ymcpRHWYZ2c6jaaqPxtBV
AxnLTtfP5NbBDkSHtuuW0swq9K8NPY1sGuFD5LdC/swszkLW4wG0m6KkQjH+X1AeXocojujIOe52
1jPl6EgbFMUHI1HWey45jO27YuSwtZhhhaw7HlWvTWYsBhl2yyJdKhO896g1wY3mF6z5PAZXnkrX
oEoRuE2RVdD08qQFrQlO96RCamQSkgjpkp8p5aAeAkCbLwH6CVKr2gOkzTsFrTfhRZLBTz2yuy2Z
n/WISSsQ+/wgx1ye5xdcpqAuInUWdlPi5OvBofTVevEoQ5SVzKe5nGRlLgCoB/cvLgNiehphe0e1
iEax5jd8OLm6jgULj7uqdDayrNABJrMMJ4NAZBSazJzrSjJIo3Ae9V/CB1KIRwLLz5jgjxkS+Cu9
2i/OCyJrYFRwxHlIabEyD9oY2FtMKBfqAk9Ltt71Zamt2vuI6+aTujvu7S5rkDrriF5ixjo23PgN
ZDIOGd6ZW1+PWRynMLpANHdalsOBI3+WwfW4xG+/exZzEn7Owf583n1xdL37VmNs6G2sc6FZkRFb
I2UM6mSKuH0tvx7YARrIWADgTK0p1yqZEU9tzCK5mflLorM/qAISNWkwm6LWLX0eHxQKfghA1LsN
yJwFaCa+RT+OMh4fFcmZ+OnRQ6FN9o69Pg5X52mAwvhaCtOpULowBc7oEgbybhDKWZIVedBR8COC
zsDcG4uhJBU/PVSEDAdaLfaUspfkDtM7ITFRGOSLdz/XB3SR7On3hT4KrQsP2Y5hDRXaSx7TGVBj
BOny0uhfGnPpdRtBRVpjQqc4qy21uJMPaAoz0CUDPBuZY+V8i/GF4JVwkMYOBd1d0Z2xaP3Szez6
nbh/7Xo0ELkFieohfQBCmqWHlK764QWJ+4sq1Cb6JEc7YZevDJTtH9xwAhiIx3JgrOEf4Go78uv8
+WEJzON1SHn2YeLLQAZTPWok38pOPW0YhDyl44wnf9et85EhCro10WoZbYB5dLg/2PJ2Zzy+nQS7
p7ylhzWwGFywfCCMQk455+o0PPbHH4eWWZCmJiv6NEftmSQO6Na5mo6gu3k9JDsd3SCqZ8vd7uks
U/Ew9lqtn/dGPzLw0klxYznJw/ko78lpv+eh2TsgEYQ2RHm3vOswUaeSWToOtTjj+EnJs8iWNmNO
yBZmTWbEMCFfD9oTnibHctDoLg3t8AzL+04Jkb1SpfaogSIpx+//xKA+02TLTcAM2qGeJUMkh4Gv
qnOjrhz+eym1dChe7iae5d+AV7L41MPjCsBtpDV8Gvhgoz2FHtnC0FOqKsM/LyMSoctlO3lcnzRE
ve+7ViZURiEJQv1ar+Tg+zCcXJ0/ZFx7s/cxuRaOTH/qDw62Lp2waJShFdafSYmAO08FNYZbcRhM
nCx2GGGH0xcE1PP2fifHAs9MiAjmCS/FAlxTKZeTg1VYdRf2CTQmtkCZBQaGSzr0Tp9zG+vob2lV
5vM/DEmklM3AkBPqDwDtpmdbx7NzXhqkM1bJVSV+wRTtGyixpiYDgHplalDpp0NEu48m+kMD7hKd
YQEwUVkffow5JNzSmn1KG1KIWn7dHf0tzEKUCuHpS+zQ4LOguI53VkXniEheQA9enkCsIqDm6Tp9
jGkEJNG+4l8RdvnWuF3JL7HVgycTO9wqwh8DR2IjlqBa67/ViFQZNoZRA1O5TycDjWIYJ54IkBDD
ICJ+L01G001i02cXFa2VUDER96ODIPfRCJxxgQ15fWsXsqjmolfVVuE/NHKO1lZsDXmZcOJx7nmL
nS2WEh9fg1zckZB7dl8v55m3Ma8+C2Hm8s0RXsx2qkQC0ThbyjO/ftWgJ0sbgO98QB1N++HwpJ72
E0npSnylEzwruY4/WUSR5186mACzp351t5SgWdwTP76q5qYZ5wAazd/z4gg7Y5sJk3G6Q4LuobaK
Et1e1UOTmiKr/pO4hSQApXnUoiDbKZSg2X+I+lEcRLNykbm+oZd6FXfqvjCrmK2B2QFfDXz0S67v
h2qSzg1jtWVfjrOublD/F1KuXiHfcP/ooI/WvvZLcbXqQbVYdblR8/mfSj9ECOS0hVHgD9PhgLqK
qtOAEl2/Kx/HBhBrwlPqHltT68phBSfN3XXx3l8gTBlZ5lGYXTZl/zuZ7tvE6EXVw0NxNLsCab71
lmNSHSy8lsdg+fPdtmD8MmkeBBkj2nTMRvEDbMXd1vw9IMwDfOTBg8TujP7RqH/6OvoWv32HlaiK
lIshvW4CpmoHar5EPtzxE8GOgyvZEIx/sB/viXU7aOlQuJWloQUCBsNkOWt/EVqfss5AxKegzJYV
06hTv9nUiDvsLPhICWLLnvXuH59i8cqj4uU70cNDKmcvILmmq0SlaUKkQOyaL48tpTQ4pAzR+nSN
effpcNelgqZFcs8szfKs/M7sQ3b6jg3baVFywNDtgaWqfGZu2GbVTq1xyrcjbiUOhtxQlGRM6jtQ
1fsI5otJfde5OoGq5RvDx1tBVfESFzUv0mRK7u9Kk6fWsOIUxUjwkRjlTwCgcsahZ1V2El9nfdH7
2/V0O3UAmkCkFnMS8TW1VvuQ6Opl6bh99dZQTDFKiCKtOyR3aHZbugEZKYP9m3HzmlWKNGjv6LkT
doZyNQtAGb1m3GvgYQhgrukWvH9iX3dLAIJedW/U0qSIdT8WPeUK+rJQP7VsyLgkMTpTwWVolt3z
4bpeoADOaTPnyBtI08L9b9H/Bb3zYvJ9MFh0CWlnM6SB1KS28s+Tl3KNLFvJ0Z93TPs2+Irk62bP
J0L9f790QWG1kBymBj8wm3ZE/ay5TMnrgrQLY+c75IBsZjOcZabI52jmw1LUFW0uYV5snT+CvPYk
rlNt6mnPSTnRyGGVsSPjZGEPT6F/dO3jSojKRm1dDny8dFFaLyU6Mdgho19vaJ4nCV9laez59/ps
Yb/kquTE8o05ZMTtaHcBXfdj2CU05lHdPLdPGdyDktTABlC+nZpWTuxIQmDcoEQepHurbQLpglKA
b1xjXoIXxP+ll0MDXlWADq6HWttikB8Tx88mwOkKXy6fQQwh443VyObHw82s5WPFoOXlao2WP+WZ
3S0agStdpSve/Lnm9/BGI+f3oVWgfEx/0j5nHmN1WcypnPkl4Rn9S2eyZyiYIo4cyoZ5dtnMGy3g
7d977ORQUGOTO4TUZSV0BBGALbBS37A1Uj/NPtGUWSx7FSdl0WyvQcnYKcINDGN+97kxctiq/ivR
5ub5SxVxdlVzSWwAy619BaX3wnw07gc8/CflmhNX0d7Gn8w07X3DcMdec011wKvVKI/Gg3tFednM
se+wy9UmwT7CfdPgBgXpdHrYFV5VZRDBKRTJtrnfzUxiMPawGEOh6Qw6mPKwg0XpyxeRjx4qKo/H
l/OzD7NUgmdK3oWwoDk1gy3RQknzva1QrZgLkxLh8QN93ZysDHa6Wbe1i5tVqyhOPwsnyfBCNNyq
tXbwqAn21EPyiEYEiC6TQf9tTIk4bz2LKGsNgCD9fUEMLfldU/uSdYNqQy+1Yva2SvxnYa/zwH1a
xcrMfZa9A9a2uFGuzQMJ5l9aIs5ni/XmF1SLxojplsKGp4nMkpy2dJomczzgD9QUjwY3l8X43iCL
jCplpoTktZwdTSRh46YBGI/MKVBZSQbXZrmtSW+dcOkuW+BIqQ6K7R/K1eG/FCVs8Q7iyXoWjrjS
CUnqU3IuoyUvNqlpYRYr0dWY1hrJ2KkCI7m3t9pjc61Am6eR/pCZJP4oyrNrz+Rb3hEHw/a3GvXv
JuVjMtdCaGikiN1mvtwJ3mj+Bdl3coAJE0KIg4Ynx9oTqNGDXlybpIBKKbDDy9Azlkii2v2FCF7S
YUtZXdsgiGPSZ1Yk1av2jRAOD9nQhfunR58YKhEvWbMu5Jd/rxN9TukRAThcSg/YGKk5zZDGAHyv
lLOGtH68nP2LYsS71Tzf3zWMlQeDGM/g4rc4LIyGFQk+rPloL32PBnGp1nF8hGnDBr9SEaO/DIOC
jCGKQy57nf2Z/RYZdp4EQLJzFpH4SfUh5B4RdzNwPlwyAKG5Ik0QakIsCxb1U0DkENp0bUlwn7JU
o02rkIYpASp/Wbm88Zl3IQpqmcaNQKPtTaB/PKsACUiFLoum7u91uvVn3ZE5x7ScPpU45DrBSk2e
MYgJaKeR9NNCn7dsHnhQXMcDpw+/7OnLnv6f/EZS6r3T9tX4DfmoLOF4271cmvZE40rMegFSTSan
SztNofH64P7yMV8Ra9nuIzijd0VXONbC9WsQAwgzxBsxprOegy2KFgzwZLmXyqyC1+bdrd7pUBNO
TA40R1sTSwvM9p/GTXNzHNs1hOAZnM9gtSpIcy0XHZQIzdbg+5bUQ9obpi1CV6QhB1K/v6m8qByD
LD5J2/f9qdFcASXRqpFzIO7aqNXIpSGfeyI+WU7QD5zl4g0QNOpcWXfiVajzuGxxFETzstGtPBfx
8lLZ86ZoHVcpbeBEVI7tan21LAty1/dOfN3ohxv1X+GHc6M8oCSH1IwUaIFdisAnvrq99KZQSSaq
kmC9b+hyEdasmWZXwcCWanyQBGVDRP7YtE1T7iNctlH1/olNUWCBJn+t4yIoIHe7AsS4Ice2laJ7
/tfRToyHlOBaYNh/JjBuTysQCj5s/tkGkHelMdy6cgcan+iP8d718JWMhW+SrZ0mpGpsi2YXiz1R
FC1pqyzzTszCu1Gl0LjEPV1dIforxi9ReXd0aUSc7W4RMEs9vI9O9AkQ6544mrHtYgaobU5Y1QNv
5g02+i5qOafbUg9CBFHZoJP+qZaps6ULUSYCNOWZrUn//NGEkZnVENOpqr9wywACNxrEQ8VTXOWn
hpkLDG+DdenCmFQT1nZOpwCVOkXiRrzjIik18fD+T9/u0ojit4SWZsVf0S7bSmjzdt4Ru4SbYhAW
GSyO8c1NdLTLvrGvEXKvTMALQp92l+qbgc6CW8W95yHNEOQ5MTaxZSNa/6HvmGQzm4A4ewgRMDX8
c8zhhxxUtBhWk7VBO5yc7pJjCqwrdKyC3otelsJPzi+Vnt2Y7CBJ6GUgs8bfXlrtUvrcttVB/i9x
C+w5OdIenZwFr15yEO96d20jAaPU+60v1rt62pbOSsBqgAD7QViKpy9LcOa9DrajXDyntVy9c/lK
zNVMfv16T6/44j/U5nWwMY3bTGzmI43khqKpvMz3ZpWWpojs8lgHuc7Yoa76Gs2RuMMazfIBC6UB
WQyZ/NfnpKFEA2rOBpEcPbhEqIEeB+v0Q5QlO/aXZI3Uh0EtKWN3mPFYoLotpVpYLp6NNhkqTEZQ
92Pk9Dk8++wn53X6oPtjdKX0SoO63Igh/PapV+Ek5udEXZZ7rVmZ6el98o6n0Pufv60H7vlAUTjW
yn2ix4833WWZjpbOi7Uq0hDcXlYjaizcH8AjXxn4AhwTHGyUqdX+jBaoO5LygWlMQYGLiNZhX9TP
jGj+3awG6BM5QBheJXgjgh80Yh9zdtSZ0lpmO01kab+GkhHiZooo836NP0QeBqmMgAbTa6MfRdAb
p5ooj7xOvXaW1z/qIABrJcn7pXXLkBw3vbq7DoahyNlEQeHelgPxIf9CDKthEcWzWo+flX3KOXVd
H7YPXwQwAk+mc7lTimag9cCtrSqgFxz3yZqL43iFbB7RD/xAXjrelTzOs7BdGjr54ZCe1A7PNyaQ
dovExaTXKdO8VH/j43hY7KaDnL2UPK714I2mEg0OLuk7ZoZ37q9boAuhADAjKWFDH74usqC6ifyG
Y8cDdVqPWx8/URDtiYAH0fSqHPuOrD37Szns0a1I0QzuGbW5G0vpCNS9ShrrKTpwyr/pgdbFsxgS
IpVKnMkQbo37umcdbyJiLQcBL1iUS7F9FkAOXyE4u1pKsN8A6vPP7nvEuMsKwWf/pqk2gJFcC0jQ
EIwKQ9tdeYoQ9h5xAVCUkjdJqh4kOqsOShM9xUapeSrvicN12yqUhSAdFdq9ViaSyiqrFRbI3OYD
14PPHfqO+3PNZQNs2n8It/uNlUL2CgMJf6bKXFFY7ajhuIica2Q4tr9GwJT3lw6nlCb+kfzIE8DI
W3YuPJ7tiIB1fiIbBEaMKkFgu71zHMcJ66SY+GJBSglNxwFGROnbri39LwlFaH94IDgq6Qqj+Gwa
YtDMixqBuLCSUlghHVtyLLejKU/PtEHe9rl7pM9sEIJvlP5xNvb/atMkISFqLLZm4g2muXthx89y
QNLugxBGeEoHl3NLu0Om33O15One33R1Y/6ldATj729rZLdg5vj0dBOaj65eDAwq5qdQH1lQKcYp
hmnd7evaCm0Ej77BC6D91cnOaLVCIYbyzFbDWoaIPJanqUvvMsW/NFcvS89HhZuNq6Hu0hfluDv4
mwfRIFKbf7RJq9EtwHwvZ0A8w2KE7Fl+aedJFEaFZ3/Eh//5/IQrTI+v8XmyDYvaKLOUGIDXt/4C
bJtWIxakiXEnKmX+SZeaYQFpGW2oZHTpyQI1oCMJNs041zgWS9Y6Oi4EOCIbuSH2ZKSCn2o7lVgH
Q8qvmzcuzBQ/uwcmFjRk4Rglb5dIAfSQymKunIXfSKUBj/DTxdfdvVAtDrKDY+JTmZRH5oKd357Y
WbrL0QXcwmWiGtmbon6aF3L8GRKkZkJQWXGTKfv2lZWnRLugdjYpQDep39bfoVA9Maon1qtUR5hZ
thn/mI6cVSBLDTXxdRy/ufnSp7Kc2d1K+miIJCAHo2JL0Hy/xMpjKWppl3eLKnkZxDIdwnd9XZ1X
ocsSNkMYO3WLHdeO1YlaRFSMX0TuD+ipPsRovtt+kJ+JtKEqITYK7tfaeop3C4woRVfBRskwLH+O
9zeCBbcuJlCUi+t2Fc4Qz+1v6bCjZqO1Cph6TCqLqIaIc6SlgEg9KjAQfkW6hj0ZobiNEZlR7Unk
cerrz2p4a3MK+zK9hdgg/C/swkY//C7qvUxn/IDr/PgHiR3CP5Rm7stYyG+pW+RrZ4JRohtri6kW
GipenpmuhFjEI6iTX5UU9m7S1AsiKAT3mbzK+ZLY4yIOEFRFsQBEVkzZ+QywHrDSQLoom3IfhAvU
jFGFlDYG4LpeoJlYL6fxt2SIk4TJS85Em0UJFF4qvK1kSM8y/kM0lYfmQ3/8xoj/sV7YkxI6fQTd
dgNH9X2TWBj99kqz2L1KbwSs3ZIU+23UHNR+ID+m34W5k5YJOZglxdRDZiT7YpDAx3GDK8A9FpUk
GUNCgbfBXc37bJZ5Alc8WzFV7JNmjaLWEk4Ykd5E4uFRvtlNLFXDhF3qrBFoocU5HQMEAMzptTla
VT++ekfsMthzfNprNP8QCSNe/pGfgiE6Vbm/FS0RvwlNNXPmQc1N3lRqr0ngncjVAG5roF9xKP//
OBEU94z7md1DuEMJNug36IVHZESOHrXBRv7iyy0wbg3R0WOq/t/f1DuKt1uhB574bY+m0bjrQ0Sd
NTCZZ2FkGzKK0vxvhu+qdv9S4IZKREIWq6KWHZBAjA6oTcOh050k5ml8eMc0aQCtnXuw7Wi8aijh
MLQfL7RbUCu8w9ZxCLhCiW+kLmPgVY4dOc5WGv4ZrqTOUyPbox4HBsApq+EI+VVKg9nDGl6zf5lr
Ve6gyorx+m4aRBVnjvILHqSD32DI7XVw08r5lXEvG6RGnxor6OnoLVIv40xH6HP79ObuFoT3x4LH
l3M467ICT9fM4D4btvHGl66qvUSFiVeP27p6aiEWrsqMBjYI4Vw3rxx++ZjkgSVEIUtvbR7p6bNV
j3vIoGNaJew3tTOJOZSU5hcIarX/gAGwq++CWcYpJiyClNqQmLvIdg5qYvrgq97K0J8j3HpSNTra
PujaP8AJPik4nPwqMxqmrkcwAj4UKfgt4DpVe4gAzhsxwi35Wgvf7QTgBEj4cVCzlVrCmmjNjFpX
WKwq2EWljC2vz/pzxj31UENu8eIVqm9xkg16870+B2bzeB5pZfId7f1/wTXjSYNRu3RVjULR2UkO
ojDlbmbyuekZJ7E45xHk1e6oOCCICtuuIdUS8UkPTQIbGQdf1DowTJxbpR9Bm+apAcclp0C0bfSN
stOVuRzI0kraQqYyBaPhiikdRTtgzjNWElDb+grAem9RZuq1XZdGWXRv/ad9+gza2K/9n/1s0VHC
jQEh+QJK08MWqOC5EoIf1Lqvl1rwYB+qesCzGo2RCLiGKVwHuw5cOgvqe4VIDNQ3zuXJhO0zs3fL
Z1VUmFveXJDzLq0Ul4c3TbmkaXOGasiXzP6S/NPCK3GoNmEbzVoKE3uzV1KxpkvTkjY+qzAG1Pis
ALcxtEtYm31E8hgl6+h3xOb9VfoSkEKnh4VP6YgwcqumiMPTl6HWcFFcKI0AVZWjf4fvi3/FaDyl
fi7eqKANybK2mIYeTFY2MJ68QfCgS7/fSN6SZWCIM/E6ZHhJZ8UbsNpaV+LKqpiL4R6S9Nq6y4Uv
lZkKwbSQZ0BKHdaSZR5L6Syb5W8XanLwAaE533jZvnezAvDk/iBdTBnW5i9VzBmgcFioS+UuivNV
JpQ+UusZJHDfmHswFsLYspZsxs6xXygECzkhzQpWt0wVuovDUZBlmhT657rX9GD6y94jUBbqIC1f
ZN9Yb6NXMKY6NePVf3jz5r118cuXYNaSiImF8KAhSgfFSO3MaPQVSZpjuyZdjJVmh5ezCFz6Leq6
VynkPLZX3PHz4Av8YmpSmqfc+ljWkDRZz5DC3ChdWPayGtwbtaiurIBg/ZKGjT2/JTuQWA90gUlM
xvteWcNPOyPotvgXjr+6hzpmVYj64x/K+Pk9pSJGqF5ZMQy570nGocg2yb/2QFkz//DeGhQoFVY3
OCy3cXjzaYn86W7LTsUb/x4IAr0viWEzT4aqzSYEqVHXkJ1E8TUo47D4/P7rlUyK7K9zBIQGlWPN
UvcB5KarVCEO0ExwhZoPB1KmsDPWG90jX5fot3IjAog68cvVUU3NNKipyxSCwrgUImFMREoaOIyl
p4Bi2bYnqPnkhzS1ck2SV7Ftee+xDiR+j2cTeyz5nL33NxvqHxOQis4muclaLjHxqKvr9lvBe9b7
g1UP6Z99eKvWmtoi86QDXS5+Jdg7N7ep3EFeTfqVVpLaHGZiUX2o6XHi3z5k8sd6yV4Y98DnY+4c
Lt9Xzct2KOA3XIJaa/WLkFrH6xyMkTppR67VZwxqCKDoIaKX3SLPBVRT71zfY/kAbPxSVw2lHlqg
W6ERzREcOHE4683IfwIrFCyr222hXESmV5VlXKve2wGFLYOskdUzAVrRjdXZkIgmcmcYUkvcxIVI
7a9cWUxOn1a6yizBXKAALrL0Gtj0Zx9wNdjByQ+Qnj93bd3nnpagf7E4CC4c4FtIK77t5/zO0hKw
ka2vdqqY7AFIlmhwk5w5M5qAV13FiM7mCXp6zw8gvc3cJvJmjD+ShNzgYoPIIyBNgYuXMtdv771l
lo8OeI7yP/9FOeXtyZp35jvyvL3J1OSYcKAIzFbqcrLQQn2RYzrVDtzL3iA0JhTiQ4+dBwnnyety
hmvLmIUhP6kbbUXSzgTrDzNz6WMBV5iGUW685XUNbRl6vWoPUXjIL0njUu2e9hu8SkBAaSlfns1g
M0Y9BTgeOPR7N6pKg7mrJ4YFDXDk3L4aX9+NziogVzAM9f77QO5WNzFWpHLCDR4H7csFdkUeE+zO
5Bq1tR9BQSCrhap+LV4CBTXqd9TNFENuwoUJQU0dILIs1cpkj3tt0iSfxi5boasotr4AwFkLo6W6
A4HSoV/vTohI0dPxCi8c2M/fQEpPNV36pleUoRyzzHb33phLZ127OIiTLq32bN8Sr2d3yQAIgYPi
wHtGOvY/JWnixldKPbHeeUxawEYh/OMcarPS5DG3S/wDpnmaMr8w2lmZLBHD4jCKCTwbXaHyQB8m
72B+awLitTmgwHAkjz21tozjlN7U2v4SZ+QOLRF7GtqTvGPfp0mZ/B3JYan5KUR3RcT2UYMlth0h
pUy6PTSjS+m4cf3Nm7kPmV284Ryn5Hdg9NV0XR15Eb0mG8otwNPFy6bBQ8SNRlkeHiEwyJDCt6nu
XfamCQ7RgqS6x8tgxPI9DbqJFdC1HZcvYblDGRwfKdjBYJmCJsBccNlE2V9OP1CBKajHtV7bf/Mm
EBBREPxMoHd7XKpMM+MEM8hdKYesC2Z/XendBNE9eC64cHH0yQf3yGnfKecKdCznmu71TgRIaAUw
9RgF7uWqYtmhMRe37z1z2B1tNkpjcBFjtTbvGSVN6PmB1oEIptsN816jMg6oUpcapfofUHy0ZNTb
G8uEazuc3GnYxwDwX/FfOx+bsFI5W9qFEx02XHZApKZtzq/J+xUdfUh5XTIok/udm8oS3TFFpKKi
ZNUrUFMMsvCGWdQAHNcr1n9jmOWqT+w2YCl80JO2bRiYue43p+xLJA9BxOOVJQZ5y0DwYQiwzXsG
fiy+u5SGBIbcxODe45wP2qOQvmNGdVQAwr+BpQPPfmJxR9lJe87Z+dxYpN2X791sS1AYQQcrvUlo
dJ6ICAba3v8iR50VU1AaJveQT9QSpfzSUWQkjvvblHgLg71gqDNmq2If+YYypQJdaEmKoRIDGCsD
NEzcB4BqWuvMHx6tvU5mp1vUARFEBWWcrDyXAxguWuurxmtWKMfDio6wD4ccESLimNMtsXirZxNP
bQDrGfYsdZUSHm9Rxiwk27aa/7LrV4R485zG+UKA6woM63uP6CGBOKNlihz0v2JkEb5p7mnyp0jd
Z7H0aFk7a6uaPy4qHCaq0ZlLyw2lR0uFfyqgEiaW13J8Px2TBk0KhABv+3uoPHJDTifO3Rfvn89U
mEBtg2tW1Dje9sTdmoT+TB3LgLsBZJSt9n9zACWQxnn/OT28/ykaLqNljgvmF5J9X7wpatUXZiX9
ktZE2fBZ2+FPZTPu6gLWl3pWPpaidC4AfSkbH2kVwObtUB32XuSEq892SY9aSt1bBC/wjubmckKF
2eW08QDzzw9/ScWHbtejlxZhhwZ9zFgDKMw0O2Oer15N0Zf180cscqzQzwwSKE7smaGkHMsgQbP4
8Y34UuBXdCb5mMO3wmFZIhzHaD7a7CoKm+KR3PEqz/OsneUOEqGGXymGuP86YjTtcGkCL2rRkSnC
AGEKdlZHSfwlB2uPafAvBoPWk4oSzzQudFbdjFMDhk86yqtHrx7bb+lDotBZ7u0TnPK61eeh7g9x
1/mzd/TxTVnyR/jjqnRHw9tLJUwH9jnjC3ZSNQjsUJ8X+eBkH1QuweLMW2Lo8mflHkpADpBTF1yR
CzcgRo2jLIrIoUwDvQ4I6JdWRVXLxnlXENfVbny4eJeVDltEt1D4w6FOvR7g8x2WcRuGG/MQLJUS
KFlc8khFkeeYUDMpzHjlDgEr8liOS8qzy4nQvfdvigdtsJd8V9Io85QRx0IgEex/mWG7MMkqwbmR
TKocHPlg25E64Rw458iNGxYBb+X8f4/OANMoH2ToqfhZHKK0lRqtaYk+3FE2Yu+8XVC8fk/6GfhM
A6a/w00NdgteHWK0LMb+wOTFGijUhY3LYayOKFO+yO3TBUiOJ7j0XyUgRF9+zmhayKbxubSVY9pD
/3i4ogFh6ip5momWm44Nvq2PWa0t9OZiSfwTu0d8/ro17nNRT0mU5NazMI/iXOqy1FteIPjQBl1m
Y6cqv49d2bHYqrOVXmLu7QBwe0frm1JRvv+CrFGmwSgoG+drzLyE+QOI1IITJGAWlGojUgGAtbwW
mOuxAOWreax+Z8IlgTHzcaIqyX/Rol1rIgngnyspmzKSM8vX98VOlphuqIzPc/YBnKFx12uiXnz9
z/4dnAiEdN1JElJ9CSy7Hqmw2usm2a1Wm1ki2rvZH93/TEDOf2HcVE1XtWgjfJGQmSfVsXBtX2za
nMdxdY2fW9rMisEKC6+TiUkMVN3KAhvwk3KYh2V8dPp9+qU2NRK0mAOVtbv69Eyoz0LLymiuDOEq
5q8/TsNhtSLVevOBrrhdDFpGDwJuRocfU2F2oxTQyXE2+W3wh84ZyAb3/TqpdvluTiXkJ/9U45go
SftCC2Jh/4fwht+ici/75fA1gnXX2C+ekEcnsv0s0iV/XH72bogrE6+ae2rF5BDuy2Y1XrKrlHCg
QTwxDfqmHWEMljFE74PmS6wvWtr0Jb4p//iug5goKGz/ewopBs7FkoTjBopUPIHr1vHRDkfX+DyJ
voZQQJpUnTlvatkECT+3NnGmPqrxvIVkygPCp9pjnWFmacu2PrYFZSEDczYkuhaxu3kyITummuJ/
BuJGOCV54RC+saLuFjsr+O0A8LOFGyP8wgz44wDI05+WxZvHy/BOndpUOA7fvXelpYSQzEBIeN8T
wI1tCMFP4YX3F27hEs2gMgRd8l12bQ3SnYZr1E6pCD1IBZEk5ivhYhDntJgfsn1nCIUSNRQHDFfD
1IXyH40cRV2075kYsoqUjBOKTmYgTSggKkv2Dwl4kpqUsL9L+fzjwGjNUGXoOvbvknN264FU9ygD
PlOqNNAizRqSHbaPei/FtCGiPXfr2tLGaFADcUfMv2bBx+p0RdAlJHGEjeSjPVihcodcFei/6HsM
jnbXyNwMtzVVoZmQx9UsbPhr3l/Ato6NkaAku3UzS5JNqemhG7YYvP91fAWXwgJiLi6yFFJiIL5X
xV9mHQsipn3e/ROiIoZoTsvYA7jnVQCxN0HRu+kvHRhaWF9MQVcC4Dqplnmg0ho/FmO44jyzvcp8
tLGo2N37PKxKo8rpUHbUlylBsPT4rTWVD01wX6Syr1lO6l2egGkG1zVWLwu8SLqgIvQ8leaHfLml
fJcbKe77YrXxlnKtwuLq7XC6pfjbiRIXbtzHInCRT2M7QoG/yUac/m2uuUmsHH/iYy8AGfE+6R5F
Ylnvi7l4KeZqrJDN0XzR7oqafsqQXB3rNgP0A0CBNUcrHrovwMJeIUa9YNhqyqyAUFv079Wm8sqd
7cHBwQHy92GCfvn3FKQRyot9K5VwvnAJtfpOnLKYADK1IY6n15ncREXAY4URK7w/K06093UhkdIa
LMY/7NILJtp6lqV4vhG+bqJ/2udF1eqcgedRzk8bFJf/tAEvo85RNahfROISwZ8Kn0XDwMtM+qNK
6yj8j5riOmA1aqk6KIgm6fLKp2PKH0x8pFp6xA7VQB/E26QLRi6mahg58UaE/2XLBINKrO2WhgeV
OIS7wzFu2VBpo6t1FjDzaU4GyWloAfn7ouVlP8q3GV2a2jkFE55KY41/FJyiMDPWXicleeq0pwoz
1aNWU/JyLqAex08YVcLiMsObRsMFr5rBrfAlhuOcnc9BFyqRukvlzNq/Pp1/7dv4neqwXpF+58bK
VynL6OPQe2NEfZ95Dj/HFWOvNo5JPAKxeWykWHrNiscYF+fJjkttY0KrxhK7os+AJU54mDpcFMjt
YlchhPIWl+3CPY6ECqoIwlknhp8siHKL14+V06pMQHWcI4gTGGSMY2M2lEKYdjlD3goFBYhfLsLB
I10cnndVeuFQqV79VP9iQpjGadROU/ZmifQskaGnTSLnIaWC7KYF8rVYn7S//xogdqbWXV7H9nB3
3eSGvEDnl62p4cxZwMKn/Z47QDiQktPTWMnE3sOG/9b88JuuMrV6Aynthi1XsWGtGt6fDbJ/bt11
NKFGrvaCD1lB9NYcWTisC0/OzCDr1wz1KCikveprR9ORTmiZdfHS+cXLZ8eJY7KPwt8Zdx+MOmvT
bSTi7+ElxMR0I8qEQghwCL9Xnb3ip7Mxiasr74Nnzva9tdFho4oiChPrNDLIRpPsbC4CNb12b60N
y+NPHWEpXrpHOPcTINuvvXQqxqMhrj80XwC7MCTix6bC2ygefNesmCx87lPtElbiNj7BN3Gw+iV2
cAMqarUuYt3GUhHdxabbLIEq3CIy3iiC8X3byzIiQUUe3IXfLu5vzJiXA5tzGu9J3rwwLPOOmjlH
BcbMIla0WKjstjawT8I+ABy3wVoSEyacTjoR04M55ViKNdcr0+JcTATlQHJfbp3+mbx/0Wcc3ULa
h39jUVJPp2uXTgbdprA4QYnTF+FJgDuNingF1107M1EGEazRLVyk9Z9SAwS4JC+xbspFajTl1WXp
TjU6D+vvaMemx+KqcgICXHJmb+Dx+yYux/rnmhQqw0lU9nDqhuORQ3DMAsc0WCNZgi0vC7pjljtr
9LqZ0Xo4HZ0Z0Yoo78uxtwbyVRw/aVhu1JAKKryayadqLOrQQkuJsrmwOX89s96z+PvEOVt/xwIp
7eHVFXb2dvrHvHL9cz13zRU/myG73qFdJvK04nW101mqIHqEATEzl7RtuKJQKt5pZTE75WAHyj8g
EWL257bR3tYBpc7ObHBuciiFbqARH9XbqZTpFOIiJUnufSxeGYcU3BMw3udDaFDRcQDXa9bqpZIM
+TGv0B8pPlTeeUTnNArZ5DWgchfitc00C2KHvRKbl7zyIrgVbpmhmmuI7jGmnQmAI2dO3RkcOYms
PKaiAnxFQOytbpBVpdRfo2NcoSUAr+Hz32mZwbOSZjqKD5eXRnTrlhAzywuUozUNfPPjYoHFfOZv
BobhvKhfmlsRvXHMt26IOzSjKmpVlm3FcGMa1k/UuSmRNeGlE1brM6pho9bjw1Z00naFj5a7eGbv
o6z7tF4GeZyDgk5H4MUKoEb3WSqSWWHPtdQo8jsWeBvEnKpBkOLgKFwkOc3QZcOygH2FLg1gEhzm
CH7KX6GbnR4L36OTfI7rpcuaG2470zrncUSp5rYNB6d+7S5L0B0hZzxwQ7J9kAPJ/FxDPbR57Xs+
MlN/hXUJmeGfMKO/64fRej/OYpIAVTVKsWHdZKeg8D4fqUHneVN/c7bttn4bW0nbpFQlYFRYQALo
dYgGeYMeUV7IR8glgzcvlFLb2U48LHsbljja0IxX7KVkt/XiKo/WD1SgdFmNnGzJNjpB62EQQ3z4
Odyhe3poV91g6dfHSyB40vTkhDTZL5Gu2S9H5qAEDzp7/HpbJo7fLbh5TDbIUJFRX9RR2UJrEGHb
WAbUjPkkDQaHIUoVRvAuXzm0TB+nmS5w+yXfgOrCMzuvJIO5kalSe9UJDXmHI+6eZXR1Yl4HfUhi
m/B9vhz62GrbSJ6Cnt2FFlJOqy5TZJG8UAmGmc3vrgdEXFfVEu+popz4YqXWdmNmqDKfgqKyiD7z
hIwFeC+yjvSTRpIgccpRJT0jZrOrsdCHvKDDvMV9iBdsilHazoUJjSvTmkFA1HH3YHTqL8HK50Cc
AcUTTwjfQUmYKHytg00lXK+/LIZD1TueKkAXM2I1gK5DdNpPEzu8wwEFWON2pdvoYx4mQBsjb9yG
yW08SQFJr2A2dyjIU0bzEu5EzWOQ+Qvhf3mr19jZRKNntVtPVaDXsyLc2237o9BdPp+v6dw2rPuo
tLlgqZiFnlBe4sxAm56dfF67Y8qXAiy1humNU6KNAEuXHPKqzbI+KIQO5CNAwEOGaT7Nh+RZzqHv
FmxBSqPFmPu3ZHzzA2RQks7UQWUpmyOErQ1YJoz3XVff9C+E3zFMR0dpKCfanTvnP5iHy2O49MG+
VgyvY3sHGm9TWuioxWV5RvdYNztqjbMFEYu4DYSmnz3h1icvlA3jnAWDpchO48m6PHZzPrrxnu8R
CstkflrmJgaQXGbPIXC+mE2NZbnYypauDArn5PsVxyIeiTbQ28iyvzn0w2mJOzSBFVhpGHvzLxVY
oZ46AxbxtHb5go+qe5hHMEFd6MHa0wsnVDJSdYp1W+rCcWaszdN+YLYkH3g0GTI3WUbBcqmszO6c
pfpiRMRQc3a1T1IGuBylQ+dAS4VmCuSebrMZcV+d3/2ABJgIFEu2KHdsFjahrpLL3Cc6hCwQtgz7
1xUH4ewCuIhFVjbY7zL7VaA4T39pyGCUdta1wiDCwOBjZ4176VfD3uwWze7fn7cknPMeg7RngUcn
6WG+ixpopDBfpivNYNs4iaDiPsLOkKmHAXHhJqR6OUqfFn9vjGRN/Wdu9sPH1khrKq8w8QGtGiSi
ROEM60rQXRlaaszOqv6S/FA2LZU5BD35Ip8UBDXq+J9E8pAOdfi00Fp1YMBXXPRjL/zVCvt8X/KX
dhiq28EVk8RmbPXumnBaByGpSKxkXNkv0DPoHNEl9dzwjJ0KZ8coRnjQ3pgP4+PN1gl6iQCO5YjP
Wif2eXl4VEF2aHWwDQrwA385TuzGRp2JvqRvuueTzcGU+KiwVPt6ereAVpS3nM2ChTHQOccLaDHx
86uRW7TRh0wv8kiOjTc/L+aVCZCTTkU77YUL5SZKe2fv4oa6uMTw0fMGeLqCybTBr9Ibz1jqJB6F
lkZB5ZaEczGUIejWCJDfGKJcHGq1yE5KnoojFpdh1wZZmA1eP3nE2U8fi/XR+fK/yYEWf7z+nn8k
ROCnkuqckPocmLoDcqUYEEAtXjbDpck45ls+v41vu0W8uJzmFK+jKsFMUJQEB0Vz8zh8vfv3tzwu
eUvzsCkHFTb67Q8L302gRCNJYSJlQuuoh5OZCv2y0J/Z1XWZ59bHd/O/GjawITe0CRtF860auQSt
LrOmnw3QjniOKTnDVS++VI+OoLLs2XRapdYXX4RJBWtJ2cPT+4aA+kDVKn7KltXR6pagr2IJljtQ
WAKX9l/O18x6TpCvD8+SMojviqByZyvDWrXkxcAUnmjkB5rLPSJfrFBzNOAGpGqbZYeUsBrKQ/Lm
NYioC7d9Pnvlp9PyDTgVNz/Y8vehyUm0vH2UKWt0Spf6NVNK7WAPXQzw/l5vkTRIPFtEaca3WthY
kJpwOYLDmL31zJYSsD3Sqz3PDZZs/N8yoPe49n3dk1z4je37G9cAyHe3Pq1+bUw6KAQRZdUpL5fO
sPTl5ZcBJT+y7t0A1qrCiwSmtMeN8LmxIfL8do1/RQA/bAgM5g1CMyHc+D+Ol5moK92BrT96qe8Z
1ksInpZtcOETjytrVgajWeDh6AtVAzFxI+P3GvGhsic9BJGt5AxuJju73ROf/GbymD0usphOdaSm
5NK/kGU5+5YkGET9MJWd90x5rK9eveT8gy7QhZkOCs7sFtCdBKDcY2NqAe5H3B2FRzYf6hIdpg0o
ihVpvg3M6VwWCnpYKRWCT66oluWQGZiPq4NIaXxWVONXp8SXm1qEaYD8EEmSg8nDp8+noi8BBals
DwcwNUeV9RJC+LRH6FuixjuTVM+JjSZ8OjZC7BuIGIea85hLDJ/KJJ4TpcvPXcEyN+vLoWOQGyN9
Z17cdwjbJOznw1DLJmFbHhmRCbyywdxf1j3MGeGH3X5NG9cSwC5wJG8CZ1PHgjUKl9TDNElVy9xI
CNm0CEbX+lYL5eyzWJ+6MAHN6UZLXpZppYPmw9x3b23E70XKuMpc7//8VSHtwxPWn2CHuSiU31zW
u45jZgVrQlmxMb3SeaP+6yj0x0FuwRgRwS6GLtxU+ajKBPYRORqgXd5HR9xqgd5BSlfH5d1p5Nh6
deWFT8l0DOic4NWAZtLVLeHmYOJG554Un+28DtKa5nenVlMBCxG7wcNnrl6R6MywcltzBvOgPwCv
mDkHOmz19j8EDZtM8ahaEwkt/uHtaHjNeTfvuRdHRxqc7Tvk3qsKs/diBgZWABEWVR1/nrDHHOaD
ZOVp2y6i2k/u5RXk9+J5fpdiuI1CitVsO02oGoSsjVJrYdg1ddEX0T7XoaDsEbarWWbzPioKVwR7
A8j+4ii11g13cEI2LvS7ZDU3LmbYG2n5BNuLI4+wEf4GmkzNQ+1GOciv3OCW2/q+7uMZHjBmXjqD
Ol3wTFLY6niq0AkNZffljbtwbyUB2T5zQo2y8fxpst/gKNT2UeexejKzWp3G5Hf7nGYT4lHQzsFm
TAoOq2qtnjIcBaltkL1TXLp5IttQkgKVFnRwJRTFqT7gZ+M/FKtc4vUdG9Le1ia4CGyAQhg3yXI9
4CMHLhlf7qgTRyqaOKc6AOvBRCgj8SENaUWsXIF+ms4mDO8dG7Z758JdiYRcd4qS6UCSzC0kGBPP
41jmOL86LnXf4GoIwqwrWXd+WzwyIdBFfoV5LA6UctZ4Wmo7BLRJeEW50CBwC9kXjopTgogkB7Gd
FUmG9xzTuDeR1f5KTduwa8F+BtVWreWrGto5rNGj0XHKXLukBRb+pV1Uy6MnIDvteVzOaPk7Gsr8
Z9G7x8Z/ap2BfaTHagvprGsWn3LrxxBZQqf7oRaLBOiJRH1e1OOHEuoRMBEV+9/0WywN2UcJSnBN
byDRHRiWRdIl4Mi3Sg1KoX6GibrJwHXRO54BNQJk1do/JFvENKTHY/FU8fEISUCUEhxMac0ZYuMR
13WnPDkPs7IIUo0tfjMrx0drkXZbr/eqRu/Qm88ofEJgjouBitVsUk6Kmh4B6OSfCDqTbSBgkE8U
F5wf+/OywVVx6lWI4foVoIcrOs92TezlfBAgQ+9DDUQSsuQHQukNnvhxdnD/AlHWN83lo/YWFyAx
+kCrjlbEsMtdrvoVNBv+BTbl2k7379cJD6RjRG0kGSS9gi2s1S1BW+56f0tZuSPhfHY3P+B3Rsk2
wNCKiQV/werWoIJ+faYqXTVPtmUCh8bthlGwGbstP2iP/4lgTAiNV/Taf1JHg+hZTmpZvWLdrc0v
vYpUppLI53cV2TmAzZmj7y4qqn2MwQ4HabNyJqMwZiCitUOgUXaPZT+wVSVjKNGag+UA2QfiC0xq
fZ54z4Z3As10rI31N9OwAYWcWjt4PjmdBgwRtGAkE3T2Ag5p2qlTVLyVnQiNzgOSyQJkGA1q48xj
WIZOhos6Kb4o3rNGxs62ReTOSWdkibnv8v9IZO/LBXBz8LxYEPQUP/gzcxi+dHEJ2EqOH7zt19vC
tu24RQJoHFz8bq33qkjCmTiHEQ8GELT8esZZlNVkhJcy2zhtNSB0eCL58lI2LXOJo004CXoREtR6
OLcyr8a2jRNng0efA57QZfumSujLDyx1cwoAz+1WS5PqpnUTzq7dpnzE0ABY/C8iy0Kg+0m40WNm
j/gmmJ1T17leRrmleSyP/oGj+Ttu6kUEZhRifRyl2Wpellsq+IqqXzdIB48s8C+eqv5hRKmUDXPB
icMOOE9UEZKxss0ToSCMs34d6b/UxnG1CAC38z7eAWrPAdZyyuMsGbB2Y5gUTs/Dbjjtj2B78BiB
9bouQ6QL00gJ18q0LZMLR1efJAnF/lNUi/J0gNUwPouux35ZJhqEhgMj4AjiUXr5hbATu0C55hkL
XJdKqtoB60DoULZ6VJ/MN4Ep/mjap3nLZEdPkXj6TBfvIbc6sPdPwyi5okwC3QyFynRbFawQkXXQ
uW80ohQoUWtZYAyhEJ/kFZVbTKCRrHdRr8Epn2I6KCSXKMj8CQEOnEZY1yEWj7f0grtapgrE74SH
SiWC5J0R6gJyFHzzrdpqw30n+2WcZG0zJLEWiitGYxG/vn/q/L0plTpAglA4ui0dy1Dj7IkbB1F2
Sb66etOKnzuuwh4L1yknYjJSf69xUXbCkBnrGMco19u1BqKGsE152aMeVU4qQi0J1VZRFX6rl7aI
IMPZhwjf2+Hm7YKRS+H4djzLUtn6+XHQRBaAnfmBzEL0aBMV/ygwVusPUWkjxvrcEp/Sbco6FHk7
TBtSNS0L8h6fCeU0oN3kAiJrYmbXvrwMg/ymIGfqn2T/6XB0p2QDubEeAHD63dq7YoRCuY0BDQh3
aAP8nl+wEs9x07C43LWCCTx1SL4fMFRQ1f/g7fn5Rr+mJcRBWgOj1gqA2ayr/nqiU4411pnFS1uh
O6LhlHQLKZxd7con2/wtsEJYulUqWYudexLAfprAArk4R+/Ro1f5hQhX01w+jCHloQXAb/dzFGnx
06G5yR3AP9hRQsKbfgyvnni9Wq/dRKLBHzVWJ05D4OWVw8CrgA9H8yVyqss6lDyrdY5+nyMLNpzv
CXebfkWHv0oxMXRmogZ/513mAC4fhCZGNH8tBIgk7OzTw+4eeWm+7PSMd53CVcCjTw+BdWpuFz0T
uAbCWDm+P9A2BFfXDihyblgdR2ScPck5cjvAqbv+Ku7/Pf1he50lxcGKAm+aH0TKMnmJB+YauB/v
Qoud7dTOIroLXPpz5/BqwBpDKJynf3HEflWPjs3HWDKvvohtOrNKDyG4wMLmCtcO0v3Rngx4qE06
ZGID5vVcbdFr2bAwkntx4HoW/7wXvPcWzN3tRffY2jL9J3r47sdYNUeqt/mN88bDyRaedJmh0obh
/5KuGotPADMGX5MLPR3kVtn5re1me6aO96xpLnfMfePsm7Ft0vqGGHkjYuQzrm0Setm0/tgZwEjN
VR8i7AP+Ee/UzBT2x9hAuQz9DyfsRQywQyveMkGh3sepXZo90tBMDFaUj400lThXnfXNdFZ2nMFl
L/qhj9uCijQ4/73GdkOQZgPnWsuJqKJ+wZiuoNvPzeGZH68A4DloqyCSt0xpph2dWo+5m98bEfgJ
wge9NqQ2g2UKn8/h/RZPFWE90o+Hk0/tpcx3EtHglK9qZZ2aA23oA1zr5IfPahdc59dE8V2hh7JX
Zjmay9XEYcSEp3hWDyx8qiFRdp40ErF4i9xkb48sxUkiK4NK+NRkAKymsLLkR0JD3r03FLiGgxPl
UtGujlmb8VJIKoNXmLwP38gEzQ6ru6zVRuZ8+jtl59uCzxA3ZCifWzHSR5gElGSGPJEgZ7aezKYA
qh0cxcafJKvxANcRrBQ6o5VqHk7cFkdzifmo+aalPezYCHQz0B6aGmhaPGfrjIZef8ee0hgJl3aL
0E6x4zeXJBP75JUtMmj9TFbC3bytesl0gWqGH7y2HobX14dHuoG4axBjDQ4TBvhmR/EPxgWzPvtX
EXMRgCIucBY4tzZ3Y/21iCTO1/ltlAbeKRHb85T8PJ/8EN3Ea69Ltb2wvkzfIPHTyXWTIy2XFAEY
AdpEtCD8It7mLj15OdHyj2Yy
`protect end_protected
