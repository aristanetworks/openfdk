--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
kWRyMwc95EZLFTG/YKVEjCwH11+azQLbxcDVPeXjzAdW/vWwPyg4o9OVBcua3KcnwkZsS5wMkhY6
y1a924eUSmrBltV8jIL8BWjFa3TPa8VtTwnLLMVObjNesF6JcSh+WdEsWsIBQwU7ZNwHYwtFnhJP
joOE6y92dSJBVAwnj+ctCyEr9CWb9OU/MV+/SNy0QZiD/SosGliaiMcElirXzLZ8G/pQYUhkSQhD
Beo6UPjXYcuOUf3o3m/q7U9FGexpZUjZp83DHTURBq+L55MzSLRrJVZz5hF0HAnsYf1uZg2O4PdB
OWAf61Fi5+ghRsoW58lB3jqe3WabtfX4YDrjAQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="rb2Ne09BK0O/LLSgIqJ8fCSNBt7O3NZvrcAfNQTQ7vE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
MLsE7bhq5ftywlASmkMuEtC2XMtUg9ffyy2GqK1QX2JWKoAb5tpStnKTrn66kB9QoVYY0nv7BVYD
gBcIx7iW5zUJhbFYeFOAp92LeVgMVhfh9gXQFWHz1/HJ5DNZhXv0ARrLeY+OHtYvKby1xVnJQBZK
0VRYs0dXni4N3IigJEVCgEzJr7C6e2qgDboLaGiYkjUtnupuo1jr1kLIu3zsj3AVjeogksd81YzI
J1UjH7Tc3PIneTLzZy+tOf758ZUQHKEcw7OkE0AkZ8mKQA/t5ZVX+fZ4cBxzlEgoR7RFPo3oGiaB
ZZRWrR8SzClRMxL6EP49A7ZMZKjtiqG6i0Wynw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="foIUQWhB8mo4xcEzQQMdG0ydkUxAv33nZGGVhwJFHaA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3264)
`protect data_block
0CPXhFrJrwCsQI0i7fjAb2OLTildqqCZ5ojqUodRIahEXkSWmU2aggG8gf1JNr0e282JrdcM/4dZ
mhhaxeD2j+vDSE8RhZrW4ZwiyL+EYRJhTJUf2PWZkHvzLPoUpytfu2YpgS/iDWRUtttvKnI3d2qW
NxQxn7qOOvUipUrjzRiJXBOx7VJaxxekE9Rq+5eIRrXz0vbMbnavPYDKW3IGm9evx8Ri8SCrHGrJ
aBOLJXGxF1az64XTO24XNaESPnjaYWS4E8bt3aw9I7ZRO1xzaAgNeE5s4lceY/NBgpjtBwwPudMP
FV+ExrW59J8kx/KdfFV5QT8W+64q4qpWBENIHCUMiqCjZ7dHXygVBZnxbohx46kp0KRHb72xAZl6
ewlrjO07ix1R5hzWCP6cQt1EC43LGB7hL+SaVAQccb8KKLIMr1K/oNHjSbhjZ5te4RhRGu43WX5T
nG6jjaYpyZo2bcvgQ0UwTi7ftJFanFOIF31lVx6diU/fpaPz0pJim/0L4VHO/Pn6CYV2vmNvroLe
ThFs6J9PhtQKetQBqGAbls3/xUIVdL7Pge3tq+dtAgaziPDecPkD0b7LcqoOqmCJlz7CeLX77+qm
goHyNtmwOKW5Vf/jqVg8BvI2Fybj6eGLOpgfVPxKkPYN1kNg+g50n6t8cvELKO8t9l+0Ihh00Wr4
U9RSP5oRtTURhYpzmKxCccc/cSiPBEV70gNKIrYS4MguUjVC9dISv9tiU5mleEJpZ9S7/mmcEEj4
Wee1p+Um42QPpXWOlkUaMewXmIeQXYMDiV9Y6lRy8cX3v0S4JPn2Y+YQJAMZRPoEgxI3zk6444xI
eX02MGOLsH6upBZ9kcIoi346M793XTW9l0SM+WZWDHBo/xuXkovBizYG6Y3mOIWPR+Bj0utbCjUh
P+W9XNE0OllFOwzPkiIVG8IYIUAJizsBEulbQWD3eEWPcnOFuEXLneAYi4JJQPiEgGL1XdLyfE1f
d2428TvnFqB5eyEFw0QHTMayI/jkP2LfwnNV9fDcOWQ7stC2h8Pc1e0hqfx72NZylD0Xvk1GDQd3
L7TFLkrmhon9N7LzbN8Zjorofjj1rsK7IRZBrc+srQPRxfYMOExHZqxKBD8mStnEC3PS1OsIi8Qb
an9GEOT0OIf6IgsNbsuFsbv7LmT4Mwew4D1eMyd6ce8L+hF4dqI4wrpHpP6ofR+7Cfz4TnSsU6l4
01mfNoRfVC85bwWYKT21Hv9aeVKoqXqA8PzoG7ZD5Fo4pjRxVtEKgy/w7kMtFTJspP2bDmFVF1Ra
0oEQH3g6ikYtMBs1A7lcuamxXUVtJSwmavE91CPLdOBwdXTEqAf+LBPoh2+6QqB3YWIrXyQNRPgD
jCj/agOHgwGVCj4OKx48UyxojjqvjY9ciMicUmfZd1zh9URpYsat2oGVd3fpIrWJBE0kGpR6Qm9A
iTJLiZcsKbarrjImp3FQDF1zXukF3J1kR1IC2zt4pid+I0mbiMdGNDvzCNHKgd7GAhN5oOnYusvf
3ucyU0D5rIe6/58IHkW7Z2pZHz5mX8ZHiYrzjA8Yx0ljM41GsmSKnh3iD5qK8mqV/p8AXALCc3Pu
erwd5uR+62wzaaW7iZPbchFxHZdrVVtdLNZ5pqW3peZHADD7VG/h1pX0/8Snpy5DoLa9SBjnaZCy
1FZFENwhlmFz3xDQIMs/K9VMNUpPg1TfWl5UzPwNA6YHRl5YDp+eYgbvAA27sfTTVFUTEP8NOQZT
KgjtID5PWvrplenNPL4TzUD3eWXp2cJKxBGHjNIWllmcuHoqKBeDp5rVTu+2qHscUc6CVQgHQOCd
eybFPz4Vrp3Wm3K5FnKwidVRKREbjLrPFveVMaxZnxG8swgC4kqQjdUrskjkJ2pRMgTEHZWEz9NV
9TyKbM/xDjBmkyw9HJio+jsDQINJfwedkTaAG9tg+w0ZNFdmxpdxIN2C/kI4h5m7TK2H3PHhqJ0w
f/UIUegBztgbELZGaxDUAWYvWfN+K7jp+SlzqP4lcqnU+ksRRrYM3d8vF7ocFL2egDyzVXuLqvwf
kF4LO5kx8bSptG9LTJQWhCpKPM+rxPttb4CCtwf2xchoM2M3//eff3emMYmGw8Za0JALO8az3drL
j3ZQopMErf5hivFvnrdhTPg0rjBlTNPrvPGNqO3geDpnXW4GERgd+ZgR3rXgnwxDhEp+KAD7RuLd
/BqZYgA1CtbvYNgaSZv5s2XxVuNvfjZxb4A5TSdvk5ZKZ9yCe3DvoK5Crohdjr3Y9LLbiL9DspoN
Ft7R3OItfjt+vl9Zx08YRaewrONuSC7t4SwDMrNdFTXZNQ7QcIQNzl1cFWTKUL32d0gXYNTrzNla
vQ/4aEe71BbDEMNltKW7E7/cn7hSUoskf5SXlPZ779eyS6fZtTxmNBltHcKI4T+z0fW9uLlxcUM8
/fu63ZjFfkfg/D2ScG4tllHdFWMR6qpJjblWHAHkQNK82S0MjlDD9cIEDmLrckojtlzZ8H9HlhGj
G+43jsxrV9ZSNnZOhal8rSgDos3Mc16E0aMNO+D1oIi9+D3aT01B5L6Q71aMCpYwbJWihlk3VOVS
4ylHgouGk5chgWgVhR78JW4rhyYWWQs4okvE5AX4b0lco6zQelGlm9RBn264i5NESA3iCW5r7OMw
HmrNsh0Y0ujmKeVOGw/mZZ5iLlbtCdmISKrr1BQLJjYQgbZQzGMPo6dzRyGZduwerjTIgA5xMUB4
ItctcstH6Azh0y3uiuawQZqwCGZuHfMTI6ISoAc/yE3cFFk+x73oSlWVbKmcpxEIvNS4KhLxGLeI
FS2KQAav4nWV+0BsrMKr2qkgB+R4TJ6WsawFAJ8Ma95cQc1GpU2/Ya0PHsdZ1FMvzDZH/bVl/PWL
k8c8Tbmi/Typia7oxUwbIxbqIlD7UoSRd220YYZ7F6NNDpScNtBIsfSknVQ4sbEozRk7JwNhwTyE
kvUxqT7zgEZiYCjIzDpHHD78PTZK5VB6/RJUbsflWGuGTnlAOX6UpmCFv3Z9po+ldtmpSQ1ggaG+
ifBAtqmvXcOcdCsy8Qm2DTWf3GMpLc0UyKU6dQBQKmZ544XexMp0URsZZbNemqgp86qvTNAJGW5+
P5DiWIOWbtvQRBUVqHlQjAKXXw4TxIUAE91+JjraEbjlHfhe/YU+qdEGCUilGozdxT6bcdW5z5JE
Y4kETFOxCMCxacqizrTpEIQ+Ej3aEr0GRnwMRiSoVPS5iRmd8I7nxBM3iWC+DV+7iKAtqIOeywSw
1KLiLL0YloJzpbnTAsOmj70ZkV5yv3dpMNyH1oM6gSPn3Q7n0axNTiwYl7EUW+Y7b25R5j3UgtVq
izIn2mgffCw1QMUSENbD4maTfYfOuKnNck8TBNJ7T1Cp++7WAqcJ5q9INDnFEtffogwG0DvRMMbl
sex1NMUmN7k6j7snOiPQS6URkOoSiTmKn+2sXxT7zIslvbJQE2WNy63RnCiYMbu9fJGwPum0B53T
dK5mMAJ0FSzNFztolbNwyjIQ2Rn+z3+96BYiG49xuaFasHcU8zJpXjcPDJx3c2TTxgdg8XVIN6xG
chSDSS78Wo9P31D7gxbMpwpyZk0QkZlirWN/rTYDSv/iv70+3YnM7x0qCHC47tKpqBjZmFUlOzkz
tMYI6HB0XdAy53FnC7cETXNFue4mKWKazZVcObo65CTniwsXbAiqxSdARRqRHesiUtUbbqKpK1OC
lGcmC9jXDsH6SBeqV9Lqu499xkalJ8fD1g2zF+Xl4iCcuggpb6mLdXTckImpwltp/ksbqcEkoEMW
4eBk+vlAbMAJ96uuvl9+NG2q63qset2gQpFUgkU/U3WThoREhELjzHVwp6r9cIqnWk8oZPxxS693
iSNTuNncfEMULgO/9LSz6ZTCARDcOHlWb78NWz1rkzaAOb8qYFEuZOc21Px7rmiT4gzR683VX7wL
UkwMO+Ey2WEpEDTexiv3b4UZHGREd4eDyfhsmHUsyKSIABupZmIyixkH7bW2IckvibHD+jaaEoFS
K8YZwzKC1Duaj0TkBv+Ja0WiFMMRBfzLXVtLKS4PkMS3Dug3Ah4AIKsi8fozXwOgT+IJ4v7xeqHn
aj7p9zPFMe7ODxMR/AXt6xbdr51wW66OLlpjPLZV9MrUsi0wgX9f7j/QavNr+3suOuo1dPv1SsSQ
LQUsACcmfb/0dgdc5wmhpZe798vmdKu+kyrZuZQ4NUnsyLSI9y4rvyGatGr2dE1sHOEyYd7zLoKB
Tm6cZ3YC/nNzvC69QaEK2hFlCgsJwnhTo6vhrwccHGgtz0pfTJnSD0OlXUH04o9bZTpb/8Vborn2
46utqDHfuAEACvMSWXsi
`protect end_protected
