--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
jCHu4Mxb4NPkP9JQI7WV2MQwWXkfw3pOHoxP/+6QFWMqNqjvsfbPIbeMOKwvAbL0p43yP3Z42QzV
WpiwvZScCyprNGa8E/iFtk4T8dtM+heTs4teG015/wLQun3+QoaEql/c/EN7j1G8V1sSU0w7FMzD
CnvRoBf/mG9mzW4hl2XPSWmbESPyr3q3sSMq63aKDyuK0G+65PWN0hIqiS5xIY9kB5guFy8IAFFc
MYEpnP0C8pW37tw/tockGswYkooN7cJV1w/lnfk/mCT41DVXy9mC3HVtPZwlXUA1ZOJD8mD4F6eu
Y9gS/IBJYBeuGt00bw/taOzNUnl8L1r0VTHM0A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="1EjzlYkxEeGQs8h2MuVgORZX6aNllS5ydqLZFU+fw2o="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
qSyepaEKYp+IPoT3KUx6cqFRuSht0rX3UiwOadMiBzb1ygKoWnpiSOl2J8Iw3Z0ugC1LwdM02EMX
XBBctzGOpSFyUTDbGM7sjFqfP6WIVveIFEq6C8TvwsBLqUOIo0wWXJc/1ApjJ8Vgb/RsAxyn9gAO
Mhvjrwqx2cpjUomVE013ob73cqFHAuv/Hc/oxgrp/MFY8n95pyX3ADqQwLdnYYGVgFkoFApB8Bvv
RuP5Pt5PCqGX8Do5ZZMHxxxnhfnjJKCG6CPNI7iQEMGKAjmezaWbcdiqrtZyl8DszKQ6lvFDL8gi
thfbLyZEuZeANij2vzGq+nYOuUQJyULlxich2g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="z3f7UN5L+4JVOv3lnoBdzihbdIcm99aIE17/xncYc2Q="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17888)
`protect data_block
hxD+qLcZ7ioUaEse/qeuSFhomx3j08BwUUL5dkp69r1EY8qioySRftBy0ckJDYzYTJAbhcalkl2W
cpaDcnzZ2w3MYxZiUd5Eb3EQhjcXP4I+9luYIpI39vRxsO1FQZBahAZAlFJX8JQi/I0zVzo8Iw/g
LGqCKifHKuUGk7avX7gcT0QCT7ixBwrXyLsXhOnLjgmIKjCrGugFLk0CyDSg+RkXZt8PEeqY970c
hash0fsB8L0YkuzDBcBnn9XspQ7kKCkBzQvYk7D7uN5n9QpMPts841ikqGzgKbyhy/xepqzPItD3
Jz++ffvpcLq9UYVIof2qdJlxzzKb2P0nKqU4LDS2djPoCQsNwmDEUT9197w5iN7DoAupF7YX538N
epTtikHli4Ct6j6ZOPWayL5NPOsVVVL1RWbrv24/OCMD3WLL2ESam8mDxSvzYVHr7YwkrOY0cj8l
1cWvnsyK9wa1XikM6wZ4WmBn6Siq3X6wChMNVr48OmFsa/r6+zwqit8EklygxgneDhgiI+7D9SK0
ZCjW+ieQca1al+VbL2FUESjLcsG9mijpz3pBNVwM9cpZPBj5aYPMwdhPrmH2vKkj06Urxxk/+450
aSOBWBAfH+EUvn7ypBg2c1iVOAypQwZatN0AOluoGDwYRBZusyzwmyWdTJseh8xP2liYUz3DRbK4
U+uP+JHLvIvAkkhrTPLxUvZ/+dtl6a8oDeS8P1gGRiAXxrRWQputZZ0oCHzMOawBSBe/0UvMrpz6
hSNy+zTVu/vv4P/h5j0ILAz+IIdgJXpEoUrFGgr7ICe279QGkbs4Y7UaDIH9SgS7v92Assan328s
VpqvjATUuu9UwmoI8ehB5jrgQNJiK8BMMTE4P4o1+eZFnvWqMVJulR9jRVUVFz+F22kul01TtGAC
ChyfVNEADaLn6blwv0OMozfnihhc0Sz6XOsdpWXcUTMb1GCulA+6Y3bKqt4Fyd8a479ExYmpIN+Z
9rI2H//scW8DypQOn29ipOjeKl+rXnQps397BItCq6LmAJtFkmjTDoHg587s96KFWuhhY+YT7VQO
HvjhWhMKkeigO0ZKdda8CJBHthJiEW+n0o8clCpjBjZjBlZSlBhd/JVtwX5hkzTMueGe1xAHNZte
LWSYpM3QTASCwiB/rs2tRM27BE8wC5GZ2Xcsh/2DZbyjUmdGnmryK3lZu9lHQwBKJcvpAy8AyXjb
J2S0k4/mA1PW1v0dW2EMMKswNgve3csquAnIC32ToJSaOvOtF+fJn+PU/jhw2pDwV3SlnhcNQ1eR
/uneQZrYooB2SwsYJRqXB1b9kbHgCbJR1lBcv6sQQBm0BwiLRmLmvurTR5p44C9I2bgMTrAg3oa0
P+AHwHJQJLGCO8rHD4DUIS9C1QV1oNPoPG0An5zZ+SWY3pJrqCZZc5OMx9xJ7rxBbqq67q2RzCj6
LiDOPcH2ZYrgSxdld+Iw4hlu7C8VC400S0bsOElYboddLaJOMCJ62yVVAsRLi4fZqgrxJIBpGAwv
ff88Q4B2WCDJMK0EU7FAaWzJN6hQG9b3kKEFrEF/1DObmE8GT/+0rpey/mKD5EGy3UHbTNx+haIB
HrCIK1UETlF7vgy/jmjmBi6WuaTzJ/9YBvlGw/XOAkEikRonxunteJ03Fbu8bxenRnpeGejfIWw1
jYl6B5WW/gpuUPKFnVBH8QGWD37X9gzODlhGaHs/5+ygY2+JGsO3yI2BKo55NyN+Na7gXIKsSsdT
3EnuRiHElyHp0np4njWr3aTSTSc3EiaXKW+Lxl2FKrXTagYXF+gpQT9Xhr7fHZLtGlTyh9Y++5cz
ZyrBOHWoGmS5zNxIKfVccyxjq0/cSX6TQ6BSYuA2tV/l/riNMLoTxJ7vz/mKGtvWYtjvXKsw9SNv
rDaEeCvK8GUtBGZLP5wyWuZKR6D0sWwDQWLxinCBAylFYYOxyEVIA2EWBFFb7WNgW9SQRL3Yqqfh
azLSOIlIEkfua0gG+3N3MNwEQBUgfy2gvUPXDbUEwNFzqNytfXAkjEcLhqwjLPE2cWd/OAZ1SCND
Q5jm154zcq/9IfwLCOrWccgyyvY9eBxBclV1euiNnPt/YyNVqWtEOTYJt/OVsO7yGVDcJTzzu594
H6Ky7RYFrl9dnDoFQumae/fNmSLxIU6XqKaBK+xfIgZU+6IL/9pOhSHOHRb0zz2CUouxqCe1JDrf
K/n5s9wDCuVCTRaQB8mgl1s7E3JlUTmSk6+HiyYBEvhrx30kKiGP/3oPyc9WfXRbc6ksO2wNhiIj
U/DLEQTWaJYzssYmfhLKWfIyGVlyNETF/40YEkI46IpXGI6pxfm5dPPGwnBpxt9y3O71Pqus6fty
OTALAytbw4bEAAdHKpJ0qEruQimkEn6gux+abvh7fXxbXoEoCityP8XLsuPflXjzKDoHHkrwHINE
l9QwuSeWAUPl1snjucEQapq1vkYgZkKlITkYCtVbFqcYfVfi/gNii6gap6qZOz2EjLyO1pOhceNJ
+D8gvoCagkddlMMgv/dpZ00mrQypHuh6pbyvnwiIX/QAusmEl8tQwmlmenYmrejpqoJGAocm2BQ8
n7FpeHtJjjQeM4Ei6sZfpl7kg4HsMDpaT63RCe56YeV9ErGHixFcJs1mwR2J1FRtLI35sc8wSGyq
nqyix+r4IwunjSRGRGSus1MxuKqXFMaNnm+DLKwQxJvMbO0cprzk5Bigu4Crt2c4rD3xGhEwh84j
Zpdh9aB7yPGoEX/WQlfqLEWkAJG+CYrRcPIjUNQQgWPOpE140V+Ra//AxtoGqnBufY34FKq1ssuJ
sTr43t8NxBa6lgjTYGLBFramJi1YAECIoUaxjEDSu7OF/79SLKxlyNisDDyjH6mvWTMJnMNQA02M
KhPXJhD+EaBh9UXr6ZScJOCnsnrqxUrUDq7lLgDIMAQ7wQKF2xWR9tO8GX9YosTFbpvQiaQc0Pzo
hO/3pCWarWpucr0zLpZQCM4AsdrP+uZanVTHaYAfdTGs8Qc+JHnGq/zVoSJR8PmCtgLrVush01Qq
bTsZ9qbjmLRpaw/yMXRXaHbWwVOsZQ8WmsFLMdYvlWo2QqEqD7gePsg7sm4nbN5nSw50JlKPh8JG
kPuS3l5Gm+ETvgxRKAcz5U0aKptftFTUOJG8hiLOLgJJq4/LVvP6Gi1uaHYTrGrOh1KbE0qv34Nu
ubK342elQIMpxPKsnBDK81ZTWm0CaQeWhfu2HU5TE3s2dMjTOXy09ntUyqBya3Z/MOWrfM3G54lr
0MtAvBVAe/9BDo1n6R3lyK0rUHt4mRJavViPJ48iDrxtPgmH1K/uGnNKnKDen4dyNg7GDFv/1WI2
opXNN4anE9KdgDegF85QIu/WJEB0BXHx0nKvpkAU9cdQyAmbQ0CyGg8Cg4NB+6+51yodtI5mTz6m
2I3sjHC3o+UuAQYl5cAVF+rPlIDBuzTS/QY+x476RzOwXVvZbFn7R3VXggzPXZIDNF3/+6x0Kbco
pBA1dWSTt8VA3kfhWOBt4BH+kWpgXgssC2lyZqftdnN7AXmHHGqj57kti9donupwvjNu3iNOc+kV
gRnKNgNwI3QgrTpake5Wm3URrSCDOehlrd1AAhLxTCRPA8bz04+6bbUyByJ7NVR9phz+DN9B0jfk
vfoqyp7oLX9RaffgpBPLYOCY8XGq5jqKFoglfqEw05pERO1rgD5i3TJysr4eKCuzi+vkxyplgZGZ
/XhYiJ+eu+wq5N6QU/fzrxwprOZYPmEYBBHKmur2YIrbF1F9crN/WkikTVxM4drJNjLlXkrSkjyG
rcmeFOq6TqkipXGno/XXBXNlqbncxuV1vnEy0ZEerF5YaETpXRQFALEE3TctIP4oPy20n6lq4MGL
I0TMyHiryi/mGK6xT+8htniBtgRElE3aLl2dOmHm0Nn3uc6cgTdlUCff+FOu3atXlIt4b2OXdDqx
dygSo6XK/5hUu8D3CM2s+wMgGEcfc/5mUyULMGP5x2IKrWDn9TKLY40AVRlZtqT0lZTUouhYXv/a
RKfm+sCwyXd9HPbqqFmq3/HjONw8MP625uosenoHZcriSPsC0HoGuankvhZoDB7CC54s1dS+bMHs
/eL6nggB3cPS0p2wJFmZSTa/qqEEzaSTEDODXnyQ02pUJYU0PoXDGgVK0Gxe3fciUtcaUUk0NUx/
v2irzI8ye+DJx7ynIDUUcdmhFBepus+WPz9z2zyeBS3K/hDyTuEJgMDteolElVTs/zUMi6BEiXLG
Y81XZDdaPQERD+6CxPSqf0rqZp3sDxsGh8bdNG/xUJJAUh0VEen4Dnh0/Kw454aihNNmD4uaA59H
oOrW+DHtTGTLP9Igf0rinvW2wYZ8yMfB7RlkOFT5Farapgmbjl90v2gZJTMNHXWhibvBNoGbJmG5
MlTutuiQzSNomo5WCfNIFxXPbeGRYVQnNJY7XjUK9OMtG2Ip2vFIz/wAACfefihO43TofoaypSCi
WD9QdzWGaJzg1598xdUv8wvZa/RSffNz5btVWHPEeLMO/r0wQhPylapfUcaIR++Yi3hNOvFIo6ad
y8PVZ6aU/ABSBHtTOB1y08Z/OVJbUpmCOKvphLXddFjxZdFaprDQL0cgTcKqIMcOvJJsRLK60rIG
DWR2fmmsn8KgC1D5glg8mTsxIK3tjzT84yrwLKpmONtQPd3CVM+8pxNlhZQG3EoYoQtiMnSlf83C
Lmin/aU/5pr5Og4sexIghsk38lQNPRJqIGieihtlU1sbaYFH8zUFC8jTgr6KJ5x1Hhmk9smhrhsM
UH3QtN/lW88xZAeDzSoeeC03NjgKtztDzZcX667rqPrs6UjJn5yHyFKODclnhe5n3XxFS/42iQp1
4jNFenAMlroP4oAp8zg/Z9LGOSdSPq7dHPuC96bHdTy/lC6BvBXQmwSJ0nY57tP2AOKFAJT02vV0
ku2sasVMbBIzRh+fUe66bFks09o1fQN27RT1SolYuiIW+NsZXdAKa+EIGo1yhHzO6w+VGp1z3dBt
My+kfvXQ49SOE5C34TK01dTlkWNERHoH/pjNCZQeL5uJOkuBKLf5TxmopM9QH5BDrWXvmVllBvXP
raMHeNwI5X2qw0sGt99an73HTj5iVowDUQBUg7xz1bhoYU0a3h58ApaNyNEtG3r4wlOJ8ms/31+E
ai1XnsEqCT02N2BqA0ZxAsozqf8RwpgHPBtU8bQ2SLysx6Cxo8LgoAAlADqnBWT4YlAY3Romygtp
+vEu4zf9y/6BMVFU+X3O8cleplipYtDFFOLaGcIE0KHtD3KnhCyfHQ/Kr+7bRzw9BHw75UFhnrEx
bBW2uIPDvO6qXRWa86aStRcYEj+vLVs3yQBeVoGixUkMLK56S0lLaSLBZqIOC2TJ37g1mB3b82Pp
Id2CkCXgKx4VhDJemQZ3f2oilppLW3ed8VorjbCAkQ07RWQ14biyvaIpPjwvDE7CBpP9PoFVkpBM
zZltkVM25WDEmtizVt0pBkfofNxQcsiVQEvSnat9qghmrfOCWxR12SgHjrI3rRLMMwZlOMtpcKp8
9ys7PizfrnI+Hy14wStuZHiVzC/x+Z9EclDcmVuaSAUgiYMvj0z7g1/uWmhbEBeND8o621rytNIx
9KvmCZmeIDtMp3XsekcGdXhCunUoartmmA3WV9hToRYO6CiiMspywgeRFiyqAFZbui/3XUMhptcC
qYebTyk+aSCoyQhjb4GJ9xZjkZoNKQQO9AZXC3tbpiJkDb4ijVdOfF4KsT7kOwzUulJjGbAfxVe7
QYLkO/Qe11hMSbgOptBhTq3jm2P1NzlMwv9UQdFFriJCsbO3KESRQ6zZ/ToHRqC1jTHY8poyLWDK
JC4VD6MSTGyvAGdbHQT3T5N6unSgNFSRLfucnOv1ENauzeY2B86EELKM747SHsypvbR1KWmL4tWB
pLLjsJYP76nC3QJpcYbcRkfGAIzIBVYZyIvum37E6WgKxM4yMWj346KRnS+TNJGotaqX9bgvPHSy
nfP+yBwcpicwa59rlJj/yLyBHOscfES+xsh5f9mOJmB74RKXjRD1u/YM9i5KbChK6Zho4815U8Ru
5KD/loRu8IOsF6U2tgSwGnFe4VBgAayU33nUQOVTH3alkxS4g5WVsbCi2QqPq8R2Xl1tSIwXKLaW
EYqH6ozCZVVa/jxXlLo9nDYETWrAqXuskja+BV9xF46BC4GQ/4SeDLfQZ2Mz4iMuedl4RcCfNbV1
n9dMtLf96moEhBNLBFjFVQsSS08xhTA8MhEEoLZwoPahFy7US9KEwrEpCPLcYoEeLp0f5v5kYWcx
DU34679BOAcOPnubB9iT1MXS1ArPpcMyWzz4OJfj1LhudUUEEVwfqpHUWOQr/fZxubbc87d4PRur
mMb53Cr7YF80YaLwSed8cfOEv9+mn1h3apNgPNDlXz0ldqOdV9iyJPm9jBKxNkaIvNmbUIYuxmyF
E0l7RqdFuEJ3CtIwZDucLygnGZbifN+GmJC8OfXSHq+9bgImdx3ZkcY0TiNVA33uq2MbRqdSAuLL
JRst6jUtr7J2BWQxJJ5MN88MaPWBcdszf1NW8X88z1ex+xo10GPECMj22wdaKTb70G5i/QCRuw3N
+1gFqvtUCV4qg4+TXY66yr/fbYSqknqTN3JDwKJdcKFNwqw0n/7vWXMbN/1soauzWb8ZPuGKoRxb
35LqAVG7dlbfolzg99wc1DhjxfRp56RgaNn+XfRnuOzeKDxSyfQBPhREFkMZWkww2M4LOLdIm+y9
qRYcnWnYOSolcmWfzbzrhEYwI5KBquMduUs+T4CaBklQ4K262yvbL8ZV4JKNaik5iboS6e865mts
af8Qu4sLtKaxgyTqH/GVnulEZ6XIJ4/3GZnlO3EkeDPIs6ce7hTfBGaOKijN5BFDiMKihIZDR6wb
CDNXX2bwsClcmA6KW6UW6K0SZMTq7fPjdZcF2M1JjtDX2ZkuucPEKZq0GGLegTuhYfNolxL2Cl01
9CJqarxUwvxLmRgjbGdLlKLwb9d4AwHrAVqzeMjjkJzAOlPZz4DzLQILJKRCOu/FmE1EvUvo/AkI
KzuLh66+uT54KNSMzqRrJEIT3p/nQVUGIFLQHptYj0CqvVfT834msQpo/RXgxhcnQiHtVDUOeoYj
SYNA+L5IxndUadLyRoM4Rj5d7R17mi+Q5K8+ov+R2D8GT1G3n2IM0OyfrAKbYwtsET+PrXpELJM1
KY1shZvnZm8zz1f9rCxJxTqSNGfYgR5p3XfqncNbH3mPM58Y9j0C6kqST3nNRsGIWI6eb1C+QNSc
SYnIUvJuHBkWueZXS6enyZSW3UVR/WOg/drey9XVUbcdTLFr7NHMVaL/QDa0mQmTRzK5c+kh7G+v
Ks+tFujqfWY3J8dvHymAwu6VHZE8fRxDBPlyCdHf2PRHlP3eMuTKR+hfOkcHV+ObheqdtTDzFPGg
M72+IIaJvl1mHS7xHBRNQu9hLkX6bgLGKqAY/7XJzzxbRk/F5eBIYEZReT7XGZ0eo5n7i52OWMVf
jszQqkPrpxDa5GWQMatzKaE1YNKFfvziu3xs4D7CqVTi3b5V5zGgrit4mCH2DYDVNLDWyePM5A2u
h2zIosm9rhV44snkXXBszf6//LVypz9uEa2MaRjloTu1ZHMKm172SNKOem8EkD+pLC4/lsq15DzY
DAhcAvKboa/bBncnFLAdmIUrhzLT+2wH2Nk4deTdTVkUBwvQU77KTBniD75+lpV0va7YPqwW34r+
Q3+9jTia2E+em35ponu7R3q+w6ZSTC/wMEwk2CfUghLuYQ344PH8D+jVFddJnlKVHgAGET1+Pg/b
IBIB/xB1u4BwxGV5Q+eaXGEIQbfb3FRvORvTZyg10nLIBl/CK+tc0sICNp69WSLIF4v811e9qF3Z
v0k2gtwN2HkuFKlqGj+78dU+fj1F/bSi6Rx/ydFgqvzEcYTHfjaPYz7S+/I3OJL8HG+z11o5aPgn
0ct8KmA056yZciyoWepHLPFGA+FBXDcZu+bKMZS6pq4H9EqdQD9L3Xty3FYEqyMPk4NnLPAbEpTi
2yOT5dbhaHkojedAinJO+b0AeolqKxTuWt/0jPfoBu7ERwJMpMpDLOdRFbSECoJcWkYEFihJc2D3
T9Easfy0hmydsqV59i2BiLMQTKks7czb5KbPZTAcbZ9/egfTI/i60oNWjjhr167j8l2DeaEfPKha
Vgk9WNq2blBCO4yz04xIisRh6ruGTuIh3W+mplfVVdWGGmT+vidMjIjlDe6vXIRJ/J/FSwmAHIqw
vs3sTazbbtFBq4yBnl3PiC3017bxNFGXkzSpUqGYq0T0E8rLX550yuc2D0o2/s7PoCtyf0wXPthb
MV+VmUzb4CM681iJ+xPMBTs0ssmY1VFJzGoW+n0+wPCSx0J/GYoBg56K87TIIlEVi9my+AHAoo0C
5tpioFmMxYxdhUK4z749F0VmSe6wOWvB9GNTJ/DbwlM8ZzxvNg1CwPG7lHRyOkvJFr4eIT+WR3Wl
xNFi5eSdz+FI/CCMS9JZJ6QtFOx3DC4MiOBtHgMso08JOQnl7/wmf9Q33YOkJBDS/pLKgcCvwbwe
aYUisxF/SMPjTnDiRiqYQgArg+a2PIgYkcwmz8eQ6Yrd50hgj7XaQ5xPwNCfszKQjCjvJ47Wb0J2
SupJUBw26rx3+G9WzhezF2K00rJhT1JBKxM1zcXhldOuYbqVrsnrwIRDnP41Hi11aqMQlo9FBmSf
D633YDhiib7CGskllirxs6p/m24H+DFNSZHAF1XkyB/Z6PLzk9Oj3IsX6tcscvvWaSu5+p2L6waJ
kN/yOmjnbWFk4ajGEUoZ4+nIzAxEDUW+R27MP4fQh8x4+zOFi6XuEOjmcYdB7LMR15HrVFvyiuon
fQZS9eniYTA/RxXomjgMSZBbombZCHkobCgiV/6MbGx/2rmlm0J/ALe2MllHCOIRMUyTMvTLhKhE
ULZ+hxripiyKhXmFDTlqEEZlbtn/oX3IGueb6EvwFy2NaSbsyIs2weOgomrDusHv8Xyd1nKdQ31Z
t941cgfsFarPu9Qu18OHShT0DDaSxWpYEBeSwBtoWOPQJ6n+Nnf3Hh47lFVrFoDWdchevrDkLhIY
OJHxkseVxuTi9lAfB3OlywdAHpntXczIQ8trBTHZBSuz4gfb1vgQ1N65c16yMYGHY5CajfwIW4hO
MMXTODHqlYTQ6t8x9KtS9BjbIDcorwdvuFdKTL7Mh1UQR+EbxxQFLVcDM3EDvPh6r7Hu/4qYA816
NPm3JwoahWno8CGWeHN5btpqQrvu4aYtB2Pep2zAsANrI3+MIDS41RtIohPm+DrAxRPU4/zfLc4d
G/MnH0t1zoyXSL9/a0I8ySl3tJoQ0/4zAwQ1Ae7G7EMBEOAmpt20k1SAijxzyf+HCSpO01RpCUBv
Bxb5yHRagtKExggytXFJ3fj4otlUZM9Htq1YQFFOzO7Ml8VD7avjqOGLqwjVr5CiM24Kl64UyQU3
ItIjUpnAAu7KK6Vx7OAEMa36DfaKpvqzaf6np1AWDSG5+/5bJhBoswNyXOm5CMD3wjM8Gb2vBZJH
8ctFnu/eZaHrsYBz1dv1qi0cWbWRrHMnnfQqjVVrtyAbkR3wWCn2P4ocqJ1+ZNbPkNR5/7ct0yA+
KrvoOz8B/ov4LY3Dg4Qu0apJb56Xk8+U4sUzDriZQVvawyRdxNtWiaHSJiAorg296sid5/CBOpqN
3g/LuMlNOXE1pgAW17HW2bFfl6e8si9oalZfC2sxCV/Mcv2ESJpLhgcMmsXaJPjbQ4Ei0+Hm/iKt
r5CrfOnrtIwH6FWhk3m1l0Eo0qmGvbl6PVsYXPjURRTn4NmWXESNe1OipFhsijXSDhtb3wpbWjRM
UIakAlYXG5eUZKnJ/w96CGks0ZbP2JqtLqKny8dMEY/NnU3hhLSjskp/mR+dMB+Zqo2KTWCQud8T
VeY8J2QcrECpHqyIYM9/ILGBVsFIIkfZ2LxBD1OKfNoqn4RmVTH00So/D4I2KKmJsMM8S/pDyx1V
j0IDT594/+RTQr4DfpAp2/EnrMcfzdSYjdXihNPsG7rjwuRZZBQIeh+z8RQzzSywav6cTq11g60V
HArvnox1oj6pA4jX2Va0S2Z06DcKgx/qQU6t+1RIR+f14j1AQb06QopOeRVsE/D7jsJ/0AC+mKQu
3mIxGY09q/ixx/JK60Tym6xo/uEOCCYBNvJMpjAY/PoTJ07/VtjkFPrRrF5zFRggvSeeIIS87WLj
mW209LfM3OuKhB5CYX5/g41sPTIt8GgewzwburBxlS+Jz3uxu/EkbwwedauPc6+XyUQXag7skbJm
bdGPrcpKtYZfqfKGM0pv4oLWvOrj/qDZMNAgxPljb9y3oPTBTfAwaEVzU7/EqjVyN33CAGKXQOD+
BLYCpR8f9476EsVJlNpw6a2UJw+hlSpvaJss+nfqfWA6ZH72OTCBtE3p45Z5hPxs6Ht710Z6P+UM
SkdQykI9CJ1uNnxFbz86pbaTBOqQ+yEe10QqgautPJamxnzEeS60UUf+BFeYNbSpr+rB5PziWf1z
8COPIFREvHZN19ScpSJfMpzivcYEPlUnqAIZE5IzYyf4hnqW3QU0hJNvj3s+3US1K2JxeVxF3vvd
oZkLabyux1JAptILDllZXLYLxXYB2Poc2ETCzDK50nfhUiC3FdT6U9awovAHLEMkhp4mUg0GWdLl
7nNeGCWqVzR/SIiHhYG32rkCIIBN88JSrg96Rgia6AOvRow+d8cC7o4lQsCrZWGW3po897h/Bgbs
f6+8bq8cDMFDB7c+ua/ECsqbggA+IJIbSDnSyvjFr2ueFdHSAua6ClALHjoiMO/krxKbtY26qmgB
cCwV9SuQYjm3MavBC7SzI4bae8+gcg+liTOhW0bZ2Ah+4YMXWytD/JycQHlxPThrQiwIDSb1V4dx
faKjvpCG24NhR5PU6M1AnqPWvQda8R8nsg5cvEekeG74EGMUXORpCzrOSDpY1OJdHfsehTxrukR+
VGCLbdvmgEv1FPMzOgi5wzxtEsmNNQGCSl+UW72jgk/qtP0zRvGH4cXp4FfLqGbXMMX5Nyg2tEBk
TOle2ID3sZMfbkSltVIafLRJDjJcuH6GklBTfpENPig9F3Te3kkZL5STHaSHUXCXcH8U6srIYs/j
hRMpQ1yBb67Qh3lT4UX4SzbvAscDT33w6bwqQ5mp0QmrkN72Pqw7UyjsO4CB2yrjg/7qvrqWXe1K
MXGeCp/S8hdR4g4qOkXPfk5TwrjxGtQR39WG0DfR+AjYw+rAbL+8PuryLoNedAuiP2MakPa9bUAb
GR0hFwNMgk3Dez8ME9ywBlsyDoeLPQcFG7dxLZyUEJeNhi+nLlVpINeXS4elmKshPuQmECQsMvI6
6YwAQTbXRt/nhKABRyayclW/9ZhemX6GFNMj2pIeFcx1Tc3jvmQEMPHEiuIrMGjZYn+YdV3AdwRL
IS2wfWDY7Ih4iL3KJMNCY6KI8vLb+Uz7b8pB86Ujrhj4CDoMF/mr3LaeFN3t1CPlhEYBI0GombV9
gLs0xCNyuzB3Pt1yB+CXWTod9xoaQkBtJM2ejjjFTHfTMPOMrKWq4Akalwk4pyL2klEi/eRWaWM5
G0iWW+2ZWBcXEQu0GWQLjMvKKW29Xr/sOoPNB9pDWq1jgmREUsoL2IME+Nqc0lxiToWBDDeluulR
JY2t5jewgv2raTlh25oirqceI3RbcaJWa5NwoeADW5HUwyqeQKL0CF7IZAtoA77mNz/BnKvhG/Ad
GdvgRTU6tscE0dvLJv7sFfI68r3nfq8aW0NROPrGxshcwNldVlL6Qsz1rHFmei8H2Pf9XFPT4mUw
Ep12JgXBllFFb6KdjdtSsW7Bvhzs2NgTwJBUEfCC6WY7wrXZeX7ueZpeu7miFpJVSRbjOXkn4+s0
8EYRpXvsMHYcZ4+6RBMmworPm6aXDv+Z8NyHdrKYqEgIYwGYLq/9bDqF2GjJPCpVXV/rY+vODIfg
2B6iiwUWIXBWkoEFG06KUzTun2Q8FFgi2I/RzVSAOs/b5QQu5msB+1NFRr0PY4yFTgzxuyX94Owd
eaz21nA1suU8hvaHpQgxC1wuL/TuvEX37vDtz9tq99+lEBKlDPgkRXoM2XC/P/MWs1CJVoLdyAkW
MYij77MO9Br+DeTaJvrroSlSx0rVLX9Y7hPE0sIoiHG1aAl2hvyTE8EdtO/3sGUPpq1HdT39n+yp
eTEkCcmTmH4eW0Io/pFhMySAR/O+sQBk+OH6y1/NO1xbpyLd0e85rLNX5tqUDgECzIh25uxHa8ae
rdEiZ3BuQm/bzQt14w0Dsb0sBsuv7qqjkzV92FYioq6xvxAtCfExzNJVsbpwsJIYRV636lKMLC5A
ciDzWxKak7yR9QTo3MLKxys9M4IgcCra2pI+z0hF/bZuItwUqpiK8FhsMl+PTfXflq6ucJdKpRQs
vMrPVfcq6fIN6plJHaa/F+9WJ2I4umIXks8YEthubPKwlTdPaLDhZC55VTnF6b6SpSxEhQjDgsgR
lV24YH6uSH83sFB50pMidBm0GkLE37xo2xuneYCTf9BHBazSAbtkRqQbNxGBb5drksqyX9P1Whlj
ZBLRTz+Mz0RL9acoNTkbI2xo83hEKboyqYWJXMOFk6aoni1FRA1ohzJLtgXT0uTdom7ctl4Te49w
SuvzvYhStFDWOUfDty1+SemG7Ag4Q/djTYBTF5h8SOQZJGVplJRUDglEAtT+vI9URW9CWaWUTpjU
feu62h5qspQrgdacjhCB/d7CwtoFsV6fX5s6BsRLfmNaMvT1EEiWGTM2ReAkDCZFhUm4U41RZHD3
9/h65Uymi346qjTtP7wJuIFCUnNoWXNKZ6boshhUXLVNZzRSyJTyy0gANMOLevPwUBxch0rV26vJ
lxwansQATgvUKNh3Wwe2RfHscQi7Z6G9ZS9nZJfxM4QeLqAMoOMEoEhb9dcNANdwjF9HGe5XmSE1
NsRj1H6afnhgTQ3aM0+ZVfl8YQi4mfnwBZwLrrxmekSEjHGi/56T8+HxpZOj7JLuXDFByV6Ym8sm
4fYSUs4diPSJxTY1XrfGCp4iuJj5r/GTiz1TTmGQI1WnngYEjL6QrVANnwGglcLlY8sNNRrkpc/W
/rj56l9gE8eH8dYIM5ztlLle50taDXLJZpTenGZ73Xa5hCis7KCHxio6RrSzdpUOll12L2vte4hy
8g1sDsJgaNxixfNMrI7Po9i6RFc5oT/+Urw55L7+ogGhVmbImCJChh9yhVkJhZhTSNG95wqBO/ZP
QVF2foKX++fY2vkFNj3YCjrMbZb09iMS+rNiqTaZ9CAvoGy0q20IcOZ5bKqGU245dPPt44jwiwRG
kJSuhdOX9T4YLG7l7mHo6C3pgqbRLaI7hsKUMYWcoAh6uHuVRmIZAZknXn6CmpbtnoCBh+2diLXc
aGSBmfaOJs3L6BWlHlSyWG8oF2Ox4IKA1b8pw8wtRdOiUwGor8A3MqhpzuhCTosT48ThVzAozvmz
Bs/VnR13UlfJDijgVOva6ktBlPMMZd076EBYCxYI84oi0lNYkJ3y3qW0WjsQQwqsoqFZuBG8C39x
wrGdV/r+wxtQGXeqXzxBaf5zXRMd/v3Of+MU6Amykcikl9mPFVMVxIuwRzyQ0m6kv0SGuDRpbESU
iuyJPsQTEzw5RtmLEWyp1eWdBQeEa+YquLiexTve+mu0mK36SeT7c7igHm8NibHOGQUVaWxhgRyw
7f8UvrDoCdk0xVioiHsaPkZNIPOwoF1XwkFYIgADQ2Ss7becazrr57oe16iPIUg18Df5j2vxhjKM
DogmNRLOu8BolUvFbYcSwz/4fOdu67S6Bnzvmk4Eoj4jGZDjeo00K+3gTlT1wESu2IJgRaxolArx
vFVo4S/utYO0qi87RVI2lMkuDciSVr5XqmqebdulDOWBgks5nY4cNNj6gOZ8t2jLLn1EA07uP2Yl
laog/9DMHbzH8IK4y3hAPsD5L7YXwEvgTAoAHgxuS/8V3U4gZA+mXmbRgrHeuCmryoNMMTV1asPq
vKiXgzGizmD7mpKIjVdLqMSINFJeYMppp878Eodho7BNSof6IeM/K5LMrGuKdn+DIebXyCniaOel
KwzURu5Wd3R+8mJ0I3iQeYUeFI/zJTTTpX92D1tfwM6KEYbLKQpaL6a9xy4p8k9b6GyzND3c/VTQ
VFxGGTRi9rG1qiA6VfRqpWOmscRBawvc4DuMCTO3cJPhZIqKs2YfMNc3UvkW5uPGIPWTRMRtGwny
KHaNB7JEUzQF0CILUAZqV3FRGIHsCbBsWLjI2+LTzLP0I9BFwNbiX8ELRszrj9/Sm2zucF1rou5G
ZaHAg26fS1pYBgSQwW3skX3zCz6KDQGe29VrdvZJ3CIQ2rB8/BmHGir9a1pfnfNaU+YA1q4RWi4i
5hR6Itlg19ViBS3nXJMsXoPAbRdZ/Ng448mZM8nbwm1Lqm6vdsZBaGfNbzGa4Z47V3OFOKH0uADY
NCI0jWfgBqDJOd8o+RIblmbLbbFBcEAEQGxTP1HHow+1Zn8SY9ACW6dwgyT0WVzTosp8iHtDfNn4
GjyHASoXVIXUhBk4SZKgQYxSbKl4ZunOYQ3CV8fTlvns4SM6hBZaiah6FlgGijSgGVfzVHS5c+5Q
biXQjWttj66tD8Fn5X9lCiKeEQo8is45YiuLvwA8BbkzZrriyWRlLVWRtQJfnQvnvk98i2WX79lk
6bItIvrkdGbzUWP4xlnfgdq8fEsaQC9NW1wOrsWQrJZCIwyw+157o8NdHeH3y3NPA5/2CmWJpXyw
2bt6scSyi03AAbGVSPwnpo1mP9cAmD1/5y/f2fppv6nlfhmXGieH7EyV7z2WBDqQrPAN8rF806TQ
1eNCf4FRdIwgdWd5sXS9Pj2Y9h6Kd3HInR9RwDNwRRm57gCcA2g20dOjrH6RSmFlvTJ8Ad3NSRAo
FlRbfA4p/tm+P5wOYOYGd2AJ4DOFmA3urM0T9qePVX0QE1UobBR6NHpSTuJ77h8ACL+rfXIU6CB7
lwa4LEVMoFCFio9VvQMFUuRZAEzjp+VfVWj3CCZJo0DlvN8xLgf5sCq9zsxn4oeZu1BWme0pnhDo
1nFKsb+QY5bJuRm4QfZWGcq0FK5yxTynWavIBy38qL3i2LFensqMObBsXZzk6s5mpTFTaMJfPnpL
kzgeVfOeTqdOtAYVxliQKee0cyQa8vhNxg/VQTSHSpk6oKd5582iCXx8/MOCRpTe2wYi/rZSS9YG
iJlMN95sXMI2R5ExQPjURleIKiE08O5HfJrOQz0dA4GIN8Q5qeiUEzAGKAW5rdp5uTEw6NhzF9zf
r0oWJRpzzM0JTRR4VgZxuuGWEiigB3kqY9kP6VN+H8fPiSYAbb0lnnN8McPiF1Eh7pS0mExasgL2
g59ddQzaB8chTEETacFuC34SJ8cgL5M0Pz14CSu7KOV42w+OOiplVXh+4wBu8i7G6tC9ggdKK6en
R9dIE9vmCjk7WfC4pyBZf7cUUa7LjsnLbJaEYTr2JKaunTqo5+ZZeAwr1dhF+eBMN7at3dhLFAdB
atk/m1+lyAvJ1bXqU0vpA7xuLuC6HpxTirntFwMDjDsZyRTb2EsSpxU+ILr9DvpU+Y/Vr8SKFTZo
wPmuBkYqOzrTv0Q5wMJgEB+5FqroksJHuJi8/Uh49/ixwoXDoBKJdRCE3XQM498JjG7qIwwhaLBA
1hyx9WcRSv0JxAHIaYYufq4pz3PulllXdZCLXU34w21cY+3Re3kcUPkJ2tOWsuX06RC48xLKz5CM
Rjqlg9xPVrJPcOhRgnPYSQrfoVZxopURQpjuE0T9fS8tNlOhp3yXJG89aA+LBz+VQ2XGcL7stohh
wWi9TQNC070VjoI/vN5EhPpFJpddnpBt9jd7FZumOIXJuFXsuzVoXW2u0EmY/LfOXOxHs1+vtdGO
ChVbsHfdokRI5E+cpVJRrPYg/67jnFGefnvtZ4rwcwFGkQVN5FZGe0fi0MbnXAIaYWnHijcr6SI3
w4nhLgv4ZLECsRyBZJKcfMw2vyK3yZ9B61ptKlTN0o4kcPOs04Vh9r+IlQJwLB7yW/ucoZL5Npho
od1/oB4d58kn4FVH0lClsaS+2erlWkC5Xs9s+vd/sFjo09SG5Q7TBXSqJkJC/WBChxlZsln7g10J
dOuFIhROypyOlYUNR3YmnjIuXHpG6HhJg9m82PlgZa9by4rs4rhT32ukb3eSDFxzAabNh77sCWk/
fHjj39A+BlphfdDrhGdOt0KWfvU4vT3TZuzXFCafUByrZYzbPYQ5Tk5XWmTsK4LItBDblf4GGK1G
iAl1yH3EdErlEekQXGHwiYNBg7pSh0EPCO5vTkcpTKy3+Pbqtj95UJnI/dmqOUXVUxu8t90C9M5a
EnmNvKB6GPAqhPENdL68knHbavMioe6r3HGsTacEA/+6+oToQcgna535tql5UlvaLnLlyjjXwVYu
GpGlI/o8JRr+JJDf9y02GrwqJTyO5E0JvRBfNMAQJkEVWbxld3UtZ9uHRilooC9w5gh/1nhPOuNY
aUT8s/7PWEbzI+0mfvbn4FdhY6dGa6LSZ8ByQPHlUNPkqLk6finorHFWU1EhrONlmXVN1pLHwq5V
P83kkscphD8wB/nnyuCdXeir51VLcut684jMVp/SKqDPuEb4kmfAV+3evkFDlAs0SrpZGi2cnIH/
dH9XGetJuOFiYXTV43MDCpznjkgEYMc0aFYLbD180/8iLw+tjujZdfMDkST21tPmVKOhUIVLrLpq
SSbbEb17ui2dQdcJsO3ZJcKu+NU3Q462G/Jk3+1yslsE8SRQkv5w+mng4WlXHPAN7cZOzGvXMDgd
+/lxqeDhRtpf8MQNYMQ8F+SIFuAdJIYzhmbtWUyC7rwmNxVVLFqoOB/gfaNidTLpWzaJ9Z61DF7Y
wEL/8vT+BY5Pl4qg5HPJ40K4rGqztIkX5eNnbLuXhv+ikAQ5fV3dYWRa+CNZHaLapc9zCrV0Adms
Huveb77Ue0Lu7xi2a5Aym3dmK05DXVH0C8XLa+AKzAX2Z5piZCAAbFHAY1CPONPHzVYCfnevWWDM
i4eL3ado6AoPJtPL85IZVACvPLtECjF2qX5IIabbMt7xOxVvcNjuVM7ed3MnFTBQsk/II5sui4SD
yfVMKlMah3wTEqhU1H2KUKYjmRxKtEF4YBCKxlrKr1kaT0ivBjE5KcOeedi5TnJQwGwHDMhwHQ6i
RpM4E50/LlGKFpLhdhbUOjwxfNC6tNn2O+nEN0R75C1kNF5w3X/IMBR1oXDO/g7XxlWzX8E7eFNn
bzkTIxl1lS4fBD7mlxOdlcTQLumOvgHkrjFtjQwXsR9dLXrTnWPULtWEge6Gmh6y9U9tB7EELc8k
noT6X5C9xxnrVr8BEqZQHbPnBzqboBNW5vmdIOjq071t1F+Xym8X9f+DKZgCsfCjGEAC1qJLKWT3
HO5jvBpEjG0MLfl73TH+Z+VjH3azrjo6l1J7KBIGJY5VhmXYxXbi/kOYGxrCzMsuDmCRs0lsdMtY
8uqKQ2k8OfBNPIOTeuMDGxsg7M3mzP2QkFxROSTkeJpiirByWLFhylgGsC8EIwx6T/2hMB3LOA8a
ARfz/VB9pFeImDtC4KtsoPp4sFutWgFORDGP6LCUKD5iwdU4tmn7/9k60ccybsgqkvdgKX6kBT29
X7RBcArVEmSsPKRVBBE33HfZ7q31WNHhYCKZFEuV23ADXy9E9qX08U3wji2ULPA1yy4YEf9bdvEL
WuQwQ080819W89HAnf0RQ1xAVvj1INMJC4D/9xgBqjv/oc3p8U4eDJyTlVfQ7og1zqO/o1740NGp
m4cuI1Cn+t7C4NaJmEnEKQjsWARqaak+eMzVUdtViJNlqwrMTo/KQAfne2cv/v+z2kjcv2FtgKDy
op1ZTpAUvKe5zc+CYiicepTLbSNmEIDFc/cZzfUE7CI2wseQr8qYPSH33AMZtyRb1zjYMkSTWMkn
9EP5o+qBv4n6DOVbKOx8j27XU2Z86f1+vksrJFNPX+AQsf40ox3nRNZBqz6tvtjXGavo0InP+FPo
8T2jnSQVhYF0E0Mm5BrgMkMEkBtTXsR8w0KepNmJpbwdMV12gk4vwGIKlS7AOYCD31HEM8skL12T
ebIuqyySEAlUd9ryIe+uG2VZILNBgnDTouyaUamIj8f+GsdsMcr+j9ZVqldeZr2H4louy5EmoCys
ofNFW7k+nTU8GlgmdXJne7kyKMeDzUG26gWu4AUSffD1yMDdgUNhOux6zE39SIgacNUhvBqABFxS
GAAzNZaJajUzqOvTHaiK9MCwxWZpgKQgi4x/V6e+oALdP25rXud1rJEzTw3ubJzvhUCeIfpwB80n
4cqVyAknirlPhjWjnWVntFyHvacuwFkYHMTf1WrHu8MSoAzOvqGcVSkBsaYj8JS+80iIcfA/a5CR
2UzZOQwBaTscdjtp/le3gAvgcKvc22T3HKwCI1neGbccJn3ax8gw2YLZrg6blFmQ0HzOJ4hVe5lv
H2Wwt739P95tyxN5CVX3mgsoowSV3WTZwwf2GNISD9JKrSj0LRjGsoeidhz/v3DnSdZeWz/kQRDC
W9IwBECj73JYy64IZDXB7L+pGh5PEk7Ilku87UMqCUBl3SQ/4QK3Zo82bFQgVaPgLF0VF1AYq3KN
MzWUCTmw7DqI/qJ95iWxieDSiMYR/VnBwJsiWMN8Z17eh+zx1hQ5FnKO1VGjv1Wrt/IHvgR/tvtd
mgKf/cqYvEoWReWxqBuql5LE5ewY3NJtUb6KMbTdbUkermozV3VCNcHrteG8PiOqJSGK+zE38NTw
eECMLHAkrL5lv3MCc104q9Gy9KbOVtsGj1FxE6A2cqg0xLDn+vQ7fx2aBkQMORFa5bDKhDES+lhl
LL1vK2td2++MhD3I7iXKZE88gv0RvHmaJaepzcil5nJ8PxAgLTG6aEryscJzBVb0XwRF2GAteSV9
Ioaq45Su94MllDHI40nn4a4RSPd5cDUEV9uItcrWracVWQYhM7hz9yhxMw1HMbksJ32u6T81P75L
EOP981eO1vFVpb6kfjSdm7VNONeTtQZgtM37FRPYkkGQ+3VAprIsTm6sCUso6QrFpCn8tSgiv+KS
KFxumJ57dNJkSYzqzf464i6GBuW8qzKrVEhn+z52rCLTYdtA1J6UqnIydzCbaJeLLLhOmWo6P5o/
EIvj2E8pJB2zTHHYZAIresMwyaF1NAbFymmJk79SOSVGuSLALx/j8Tn0gb3XLPsQ8zK/57a0o4fx
IjWOUIZ1lKoYGmgXb4iNRy/QTT+x2yr231psp/gpODD3OI0hRvmcm4JRqYMWa4UhAQMYpqzWWv4h
nkzGUhRFvlpq9cwJIJl1IUzEYOtsGQTwQGUDEnsxUvr6QHO07YAZgI4gx4RTM4N5amM5O9Syuljp
ct8mM1asgLIW9R0cIGYmf9HX2yIORe/+aEyN2jnjfVPXOPSuAaGuPx7v8Urw9cYREYUogPXg6Y/0
qBRObDifJ7GfURsdF3DKKYkmcGTCY5JjX8OiCDR3xLdybs6Dy2zd53s1tsBYvxQS9B1VW4V9Be0q
kwrv54GA8ybOTOVK3IYBJ/4nKaWHRE2hYvr+7g9pigTsU2VTO45QjJ4dcYqQxaz3Ag/cLHnlseL8
MO/rfWo8wQ2TO4ejlFeFxpdXAPea3y6cRJQybniMu/NExjGZuVklfaQFlPSdTKhE9p+gwliT/D0V
j+PauplMWV0Ns11AqyFIXwuacXjFzGFAYhy413kLXvvDdRdfcpv2iQBK1dqMprCTPBQERxjX6wZD
CnEuLXKpNTZzEGf2WZ3o67aEaH3OQmLOF3IeMhvbIKlIKVpC33nYYHCKtzIdWchRSsMy+PDh5Atk
LvxLpGcr2CMwLW4OVe5j3ssZZl/APdmsarKe4oHpy4U8xRE5mPYuWLn6a37genyK7lu7U+PC3e37
EM/hyqpP5WfdDNAik+GxxvWX+YzLFcfHAbRsgesjoZiUwRKuLK70K+ondrzhTqCJjb8jK1gSWDp+
IC28ee3AaCpmbwWcaN8SKesxOVEHCEWYPMG2fnAUliA0y58S6ZgKVC+BTmsodBQ3ea5kLfuBNHxN
4hchZVGbEwahQV5p3mJ7W8e3QlICIfSHkMHbrw0AwjNe0kVJDfd7irMO/EQo2a+dvXnqcHb8rPm4
c2nih8aGQf9T8T6qke9aiW21I1KJYey2PGh1+hgltSZYkKiPG4wO5jkmdTsi3MGvJCQzMgOy77vi
AatnFc/H27mmmsd1inwlH5tBYSwFp82Vrvj5c121qQ2fWAtGOM0/rDeQwM/WTRfk7EkjK4O9k3vA
HFAVQBIUSakZ/pRrV9ayy+yGvtlXzQP+fe02srf5yZJcEipa3+wOGUI/rU5Gm/jG9pCUBfv6esk0
m92ZATxp6f4VUPwdG+H00EbxxY+hJhy559HDH3R3FxtHjuiD3utORJJoP4KB+StxdFWbRFM2Ebkk
4V/msPCkoI+1eJqcbK0ciEEP9QouryTB30s07JwGP0CsFhotIHye/amFlH3YYryUCoP6tRWlzjTu
O6ZV44WmYCXEg4Q258Rej92lfIQhQPT8HiTRvtzVLk9sawBV0hKjqnTJd0AWirYZLIhcNLBzhjBk
WR2XgRfPVLh83tOpmBohAHlr1j3j5TXwlrAP1uVzUg/orWBhajC4XrYXYHWZwCGNUCzDAjWNN15M
a4pS+CRBtiDuyUd4c1FmMugMkiDEmpIVQgxeFjTcBdHmByLvRsg4Wfcl5a1pf3cEGWPGuRqlP1DP
E8Nk5TsJHN3eKKjUchWaXrlwF+bJPVXEbPCAhhvfrUbi3rcBPxy93ogBUKRyZxdnYPt3NHsk1CV6
GOCTUQ/tbZ5blheU4Q1KDyMbObA+mYDD3EiwKQIqDk332PMzjXc1ubvgtn/T084WKVTIP7MBDyPx
AlmvkTHS0DCKY2NhurMdyE3/Z2Zah9coa0hvA4yPECSrJVU39qSJuy6rIjI598jvR6EVj4ywA5lV
nSC6FAoqkl6xnMvk3Gul4zR9ofxTmvZRuPnxjf6k9dTz3ULzisC7ABjf1vhuagFSiq33rCWKPXWB
xkxjFkz0m3P7Jqh6N/17HfhwsNsFw97cRlGK1IGbJILvAtr7UiDC46vt5dcAp+Hs3YxHQfPJd4eK
UuyLPtZypCG6PXaVGkRhVyuykSvf1mZdTqwia8wrrfDV5Cr5Zq/JeIm1earg6rUqQVrrIRD2gazR
jvROUQf1pOgByGRdW5D+DMtS8bzj4m9XrPbRl/z+Gin8+ycDSuUFLKOkmWsRQmQxem4Jm/jXlLWH
o2mW65BNQzeZnH9dFAFQtBup2SAT8ctQBXy9dwt+a7F14UAYKlYF1ZkiUFt8v/uin989OEED4G3z
aSclbqagxFZ3jb1LQD8PMSIQ7A5ITCb+12WK6oJj9dT6vsFiga6pDXkWhFIoqN1S18/+rNRz6ntO
xPtTh3Z4be3sZLjW7r5BMEzl8dx/c7ct0fGlLPlUaqqVX8OsgpWf5VxxAcrmcw9XKaSu7QNHeHsD
jZL1/R527BZFWtEdVqKPx4W1ebIR78LP6tEWX5NO9WEBTXBfCIKrQAW2z0lcDOdXXOBl+SHSx8/e
/05tGuHM6/7NBS4hhUvdE8/dVN5sqUWy4d46ittBAOw9A3N2KASC/OwL6n3CdbQYJSHNgS4q2vCf
OmopXTq4hBTWo4Vre5q5siRg0TDmICqCxNbx35Hbv1G9WPWwNgROnDgZWxhpvOocOe0IbLqVx22o
+M+4aQXWyWgi1dM1RBqvSIYRhgtL4p6SqUlBIS6tdltO7MW9nEgPh2X8cwX1Yhz12KvFDHYxEcx6
NOzN3Pkq3NjS2IIxskl5ZxSGOv/DQNW908wsD0XeyoI3FrEoW5fRng+/F6dwz1MZpIC3kA8gpLx0
WBmjOLV0XxujAsDtylWIdA8yz9CLX+jOTZ5+zu1tWGX6pmMVMiV4IOlfJUs2YPniJMLvZzdKfbs0
O/cvXeKgWEFkS90lSpDzsVFNQ/MaSgSMyb3pV/98Et8/A7v6MqPg7xoAlWag9DMVZkK3uZjnkzd1
ZUTk3BrEH5FF4itgGOFJgRLnkMk/D5jYzjRE107mH5ZWHVJPq0tjZbeXGFRtNhZqhjOq6YXAxUpf
92DzFPJBis3coTfaNj7qorsuM4N+iOGxtz+cVcRViAgxB0W+nT9I3/9Tal6WphQ7B64b/ElYgrWb
6iVCR5VYePyAWpNcmBAVkoWf79yjG+W2StK65eFrqZRdMWdgjK4We+dUKz2TtXo/5/sdkoKq21lK
zYHxyQzYomrCrjd7x4hg4mO7zBYSM0ZGRwVjem/9biJSJTvEakZqvZH03Ns2w3qktHB12MdEajef
rhcfHbEkv+8poAojsJRCF0Dhb+5ZkQAhB/unH4DXo3Nptguq1xdsF6/60b+FAMdVSSc2F9mg+62d
xQs58nfk4gntgyObuBzquNR963gtCgRS95DhQ+W3RoCbjN6tllsdtfjQoSE5YbbYdRuUgqnvP/GS
A7qcZoKHZav1tMl8XEuQ44//v56rsVA/0LWgFmYfSxZjaYs4T52y0MTY+Jeuw9oJz4+iRNKgHCfh
EFXyHWNpFvJVmA5iliYvcjQMlE4cvABdkJg5Wss7x8We14db7my3c4OYEXbUv8mOL7NIIx9lZU0D
BNptHP4Q/wxRr1h5j6qu6mHg4sp+nHC95091ZQe9I1mIf2YGCqYKUogp2WM4+PsHXV7oJz6gp/tp
VA74gw7sk8SFQf2R2ejpN40oqhYzVSw2MFIV9rz/vmge/cjJsW0bAqlOqJ8tmaMX1tdDzQaVXanE
a4Ritg/RRzMrU8LkCqCkj7zdl/Z07L403GH/U4t/ROtSAmhGsQ0AMLf5hAc2odEcLmlQdoDWApOV
X+7WOQmB6gfTQN5ch/lMjHC0pxOeRdmmN4RMvB/GhWEKgxFLKC3nZVKwcuqD2DVGbFLWaaFYNkCJ
xcKU6kgNeqBQ+32pwlhl0Eu6lZZGRN0ylO36sDr6jWP8vIF+EAQmrNxFh5JCmj0HTZwtrSRvhLx8
WkFARn5evqLASf5VNa2WBuoEj8irlkWEiqhwpu30so1Fo48kyga9ukJctFh43+jJRQpHcffgthar
usG63BUrZk3MA2AH06zyG2/nsXLSKf6EpSFput91U+bxA8sc9CJRZ1Jyb8mtTNIll7AHthVK1wLj
xQHoakGkoDxqh/lOa8Qxi5eCHRNoQZCHb1G7DX+lHDSghWgsJtVJBm3TcKuf545WNGkrYkEaIhaf
ZiN47zdL2tMHKrOVkzoxyjEop7MOqPzogzbKrii2V/8gqPKK28sUSMg11P8PvIP5Wc4rI3GfAoFU
Qukd2JkvAHkPuVWUJvdv0p1tjn4psl//jiz22nXLFpu2uLsXp87n1HayAYQJLlHwkh2zHBDVed32
8BcY6InWkV+8xJuvXFA1mTD+/cQWuyaDkVH4fzvyNQVq1EnxyCBfkcczYWVTT+bJ6NOL5TUov2hY
GjGN9xzonyjfi/Js7IDJkmvsGrgAS6eTfbPai6AOuEEAz9H3Rt218zirkOdek8hC6tdxfQtIOW6T
x73PFCqEZErI2PxkYGtSYaMXuqgISbpfKalWhvwjAtKUFmce5To4pswtwn+wI7BNlBsQmP49vH2Y
I3YsF7hiHVYB6vGqimnLxt6xgW5u2U6Bgy4SQQr8vdMduJ/aHBcHEF1BdeAmNoWHqxS7QX7Ruh/G
HaXZXZGCFC1Wx/stDykFiGGcFCMBAjEs5AqxmbVgBm4/rA0EN3QuBB3DzdYGrr0=
`protect end_protected
