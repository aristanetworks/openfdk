--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
WZUHoZWCx/ELUThz1CmfBPMYUakhdpdQZnl/E1hhfwi4imBz3JJeYXtWZwXcTTf5uKQgcGmZsHbU
3UM8ppCEag98DHd3S72Dd2POuqoHSUL9nCMhu1dkiLKURuVGQ6qHzhgQ+WTEBedZLnR3ySOTsuof
wHGIlUdAQhu3vUC3/B67KtpvH5PGJBJnEjKXFmafZx7M8NLJVk7POgfN4jPPYltUSzGsbnAhjBSL
TFwXx6WqRZvO/d//6orB34vg84CCTBx7wPXu+nf5ZWSMb40fMn4Q3LvP1bxchtg81FrY/yUEQGjJ
uR9uVjcYu4HLKYcvWoiUjPGoMD2iqQbk5xMqHA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="RsBLr/3ZFkPd+2NkZdzNyTk50Y1qO9CmUJEceFuEfcg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
PYjd57N5KrJjlIPZ79FaC4Ez0sPsGHbYjvT1LQdWUqJUncng5tPu4GTTIqmSmBkj8WYbPuwZSXb4
+ZHSA674TbqMCGSqWTdv7eL5v4E0JSAYj/e7XVB/TeFTTyBPPwPS8dnEnjyaBPNyqASkZXV/aj9s
SWVA5VvlTexWLiBufObNl+TO7QSLwZXRobia+g2NkrGErqNA0hwwSfsi7hqKCFUwKAyBvoV4sxCf
3Kml6hiY5d7aOlS3IzYw2fntGQeW9PjEg9zQJw0wXll/PVGXeB4OZCMAiSQSkn400G/i3sR1ToJo
SuIZADbHNZdJqyVRF+FWryPpDBKTgcOlFaNx3g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="bCsZ8ifn8XQ+Ln0fv2mVU9M+8vDFzb8zMsTQfCA9GnI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5184)
`protect data_block
ljmXlQEa+Xs93HJsMj/NhWhQwJQJzx+eiOH7QqftOPPLSpmvg6VDOCtRJtZ/dJdZah3za9q+2xX3
I78ukK0tHE2RCzfrjSo1NoinzdKKZgq8wP/v5TPIAL9wueBl2mXWrzVJoo/uwtRhsVLznOEeY3M9
QBeIJbr369kvMuyvvg28tu4g/dalxD1g9jxyqzPSzhzx69OzfoqiAUTYCGTKccrpDAHF4/FblI+0
Y+oLHh51U9r73s4eW0fKUrqDu6inXET7f5XbCj+yKNNnv+zDsf0lrrio6LP0c9xakf7d5rQGq/lH
J/EAgUXf7Wht2QlCAY0yCmfQETmbJ96n+sqLi3NZMQm22fYAp/XE/la4Qgleu+BlSZtHvICwlPKY
jhqQiCqktVRYGfvVLDC5+O5sVs1QiysI81AnZunSE/OvaeA6noyiA1yO8SVW/v2O+1ifQd0h9CLP
CSFPX+hEOd9Pt8aspyM1uCP40tJ04iTCY2//+8Xi2ksVgLj8bDPQjAPAeCyTG8yu5DG02AeIuVgY
n5ye39YFLAEORYeihrG8u8H8MuLey+9L5n6v4drHyv0eh3tc3rQiI4TvaSrCjXGOmrwYeW7jIsLW
+VhoxsFnwl1UzmUkdZR3uNoueUjQLH26KjxWJAtzwxJFPEomOHklUDYa4FRegkrBz0G8DGB6JvbF
ECbxpCLKAS3reO3tkx9/Rvpxy0iPo2xRxjHIhHBJF5XXa4s/1gW/REO1ShyWzOCMc4yRZ7BYxonJ
GKpJ2+GHddvx7WtSHg9qqFQ/HlkleRpH1m6/SL/qMJ1QulidcA/meW66TKvhqRQEefteDPtTw7wt
VJE4Bby82FO7u1XZOLqnInGimwEH1sOuNwRwT0IeZLu2+Y/vI71yqGg+1qNNXg41xOkCqiQnCNJx
aiDANnd9nsB9bL+zF55iIvkDVlrGM1zDvnuEVR844/kdbVba9M42Cb+PtHu0YPJ36AxLID3SnBS/
4z3qk7a/WhKqf2GpPj8v742zv1DQjNQ7QfE5xYjTMD9iLRMyMeaQSgk1JQxzBhLG8RZNbh9Fycr4
tRCiF9xZB+4LUUE/M34E9Z2jLejDU5RWx4baB0sRugNnxvPPQNIoLbQaFzph09N51y5cZCKCJM4C
Q6aKA7NdkQLCOxdGBvj5rGsp/gWp45OBEiGrN/Mm0E4lyhT3dKr0bSqZY4IbJkDuXvXavYqjfMiw
TG6iCuUmD0vZwctfmYqe7cTtOOuV/RdRycHnPajb+Xmy2XgF3MNkjV1Rc637EIj9XjRgpZXHQq1O
Sols57T4zH53xLP+vlXfDDtG5JszR8cI9SVCM793cbq4nEFlrGbQyFZLjtvnL+hoSY8GBkR8UFhb
LQEIhdDycjlONdQT/9yES5fXqpo3v14Ot6VnCS8jkxaalfh/qQ7+vNwYLhLRQpBTh8C+ue+NterK
8MWkivh/LbbGOpXd3oNGuft+pDe7xJfb8/m6TffTNcewjKG/QjlJTNAZIBWBm9H7POwpvAUoD+Te
w2LvRLdlROw693SZKODlSiS1PKViBu4Z7lC+CEA0Dmzow2LExFS3xhqKbWFkXtqHZ41g5TeUjZLM
+AgL638yGKXB5gen1ojOR+Xk7a1rFDTLnNINU63ps6JYUzftJ6nFkixB9C4q7ptMZAvA8d8fybnv
CVj0HCnFGYOiXtv6sX2+EU4Fs2cxZXAtRFdr9PohbwxWVo/WSy38XYpdrvFnc5SlBK8LDDFrdwb1
x8b0kT3nRfU/38Ku17EmqhNkhqZFHDEr/tDkXpz/d/g6PG39+FlKA41Xhe943r0XS9zx4/vuz44i
A+KsAn+a+tEExh+5NWgrs/aQ8kElZNocKj/HcJLZcDf6nXiPj83hXqLg6Gyl/V14aAtJme/LQYlX
8O22k2nhHTi4uadFHfEhgBMrwpQSLVd3hDDRN8kJG6z0qvCRN6L66GnE2tW+DLu+fwMvIPVYw7Xy
g6FrewM3CllOAitZn4InpT5kyR6mT0NUxa3lUjqTCa8KDljtFPgXF9LtFoGKOitlDfGlLxcu7KSk
fZ5Vfeedf+iwgcrM4TKsevW1fPGGLTKbOHWuTunBb3JwAm/knps6X26TBhFmbV+SNWDRx64LMBL7
x/H1XHayYGzgk37YCXO+U4uzctPcRrjyY1+6a9rhCE+VLReXr5v0vo+nOb32prYvs71kihQa2mwy
cCfHzyGyE1AYd0QiR/cyANmJ1XMFOCYX2FgBTNHiD4+HnNv6lg4A6Jgqc2T5B50kwlg7J0qQ13xg
8KvzACdOGuR3+mHYSLIpAsg8/dWOxEWU5kZzPTEWwzGjW6pXlcOpF0tN+zre7tBomZAQxMiCAxR+
iHIndkoFjp0522IThw+8mpShurc7VKKq6JtEbuq88KdXOn36uxGMpfjXqqGtILl5iGfJgJPGgwvW
Fae1imHoBSUAmYIdw/jOROTTpmFVL65bfFrJhEOFCol8nLqpJacsHfIZc4lYu2/B3dw8V/gna3h7
Tk1HoxKQmpPpWf69DMUCQpkupq013rhCenreBMQcaxIHXsjp0iINXhj4wBVo8YthA2hUMFZIrGeV
/KY2aAdJQ8NsDo4EP0ixq+bUh4JJKAo16J+aGi7uNr3R9YxPcCPdBY4AdRfUX1Vo39LTEZWkDDvi
3VAc5aian3PVs/DA52SRPqnfB7NY3sZQZWkfieQmwOreQ20tQvtMzyaop19E1kDjx/DNsAEZzt1s
Zn6KpXE9PGOpAPd+QQnOw7lqaX7fmfgxQ3yn7mjrKvymvvIy3+EZMOaU+eVcZxooziDDuqJ7Q33Q
5FkEQBMmCgvlY0l/dZiuiXI62RGr6g2jq59N3R0owgeo4Y5OpEnlobZgGmuhoZh1+olzDl6ZXT3N
j4orEct4vNp7BvO2rwjZOxJzHQE/V0SS0Vt5qIzURk9Sf6Z6rYEQNeZNWZoWwIbB8EVbdCtILSf1
R2r36hVPRhOgD5VpLMO0hKkGHMuEqW7766wLgGiOlB1XDZK7GU/LNlXjT9iiDZzecBJ3QaFDizne
HMF9I8jvgvc13GOMCVjWbQ551OmVGvFRUuaCxANLhjs+rXrdI+4HNK8AB8a1LtQhVMMxQzFi0r2L
3TtHKOo/o1gQvOCPfVwILHJsjJ4NiFmo6t3dkr1iotYg0kS5jOgQKvMzYkV75M8G9qmPqlq1cxxQ
Zww0kbvqTGMwjoUgU7qgzMh1sB89QpbJRHL6VGiu5nOaLKipXVhyEeuxMUtOZ1spTCbNk0qFpW4e
8DkjOJPn3DVzUzdQVMegRtEDsq2I/AYMetehY0s3X5RMQkQt5V808J/bI1yH6urgUvGxyA8WzwOs
Ek9cHT1i4FFGFtFFy7Uoo5uHkZIU7RgUiyOOqgybT41F2DDFx1/3Txy/FpE/WttC7HHoIXs3xB8P
Cn2Vzr6+q7x2kW7ygIlHyaKd7Pj7wI/AczqXMOxsruPRdpJcWfP9qhujQjeGX4WRk3zEMLT+gpbF
YFsfoVAS2K8zzvZwv/fe132d25nDf45hMjhb5bevygc6GUDJou3F9BP58NEqGC52rgAHc3TnwF7r
euB0gP2d0g6Aj+TpZKkQe3MqYG57929FynmRJ4x7MZ9IV6WHnNpZJKW+ME5FaDBhPORGSpybGVNP
THVdvGCwFu/vpV/2O77N5drdTyJJkigpOAM7cLRhIl+m2vuOcYpzBYCivs8m8cWlQVnoXdnmpRYd
z8zVBYnbNQceFUQyZB16zFs/Yc/pyUZrF9lCeocFa9XhmkaQuq1c93G1Gxl4ucOopzcC2QYIGvO4
gznmsj/8WRhqWejd2JkpENhJssqg5P3A6ny0NUdSJFzN9BX/bT0NtN6H8RIfLF/VPK1g4OKHWbCT
3li7SGehOZb9YIyV/tXHczvf+KES54/ruVDJtD7oK30x2Ya4uUQyeyffnLWbrZdp4/R1Iqa+KXtm
PMG7n/Ak/zWbvVmjNCHGX7eM2hUv/HUNTUm+yNJan3m8C394QzZcaaFyuWKkaFhyZY7TrdND+Yj8
D0vN28OWoyhr2VNn5oP93fKcPD1wvklLyUR3yH64M/N4hVH9ant09ivcJSOhSt0d/QEnKm8Di/0b
4IjycsNbva1PqByHM7zzHvMqaXuHlFHkk8/U2HyYzSEwkRAVlxlRXyEv0mP6yYe8eP7SJXK88DTa
miy325GJU7VXXYYp2WB/BilE0bZq3meACTe4OUZikS0WoixM/yo5XJfJeL4ZBrLEh/fa31z7eups
3OB9mCJq9vjqQlUQCIl8FQJU3UPxqtBm+JkxhnUtXFdKEGDJMncjrX3UPHLAlDakjTpCjzS4UfgH
NGJQ8zlrRVIpcRL+ogxWVwZpmzRNzemMBfEFiNIC0/SmDdKv8EH4hnUPQ44xkcDveL9jmp0wibdV
CRaUC2c49Og4OYSWrRWzX94r+xXx1tVxugYGB06Skw0aAts7vUCwWxRM2lJvgpfZ/t10zt5ywBp3
r1edoRWIqHGt+WC72RTX0qLgpjmiPTFWYZqfVGh9PqpoZlsklYJwZiawCX/quRrUcdFFOPiYAXw8
SNyf0L5cO/emQUBXB1MugIYe52Whm8+PHORasxE7+jKK6xBOq16vB6b/JWETXE+V+BfF/N+9DYb6
bY6Qm35Z08GMLSLONE3k7XnVBpSoPdb8HKxvfElmvpM1V74tGZx6jSZ25tmFiI9tO4yFQJ7Dbs3d
3fM/e3maUNQi4bWDt6itaLiJHxQNAVlMeqa2307zRA5cPER2hceLpAmw1az5+6FwfpN2Turcane0
GkYpTZH1wNSK3oX24K00dcI67C08LQ9wG7IfKrCSfL8xQzzO7x7ghbvsgt9PqSLShBS2D98h0Abh
YUBJrcAcxzGSas4nfBP9a4BbOhxFBxIh6P4cwoox3DzG0xch/SPUSelVwDhVrF4u8t/Hm1Fz+QXr
nGyhtrb4Pbt0BVwsETw00bCvj3f0duD/Jtdyf8Fm3vczr/BxDlqW6k1Trvp63zQqw2s+OQWsFyy1
0QkRR2PerlnZq1ulhoqpWWk5o5oTf6K7E2ooxuMpOnt3L1VbgxFKg9qSQJtHilcEr+uE6ha9oftq
F9UkU3vdRCROcKsQUJAx1/VmG09zEpcBocFWeBZIcZJF3gbs1CoN1OQoRbu4aYqssVTOFb3Us4AG
Zx8900CPMmQ2dh5cYZQ0F7wIrm4Wek0gqN4p/Rk226n02l/8IN/028oHqKoSTQhrtZmqm0+4Ifpz
8mE8iim5BeW5G/4nPpj4FLcxxmydXaI6y7qc6eSg12FZSdkkkoDDv2LHpKytzwq+8zhHuYidTt4s
GodwEsfPovmDLDmIpfgt9WR5gv3DU33GsyLjOs6giFuCU+1eb+uqtCvFG1x85ivEQN53kL3SSW1Y
rxjzmD08B8PGqeBOsjaltq/eExBL1ZuZgpc4N94ikebJIohk7fib9hN/x8sQB/qrpUAPXZQr2/M3
4VcsbywuiHjxsXGKZ/FcBs+MEES+KZ0Ei6AhKSzRUVsUDLATibcKO5+Dnio3pnxOlg5g3I6UXtqs
9phpEprqicJGXz1U1LIhpWkqX7lePUg8KoHEIWsCJcIAps2bv/MknIimtNP+R7IMT1oMru4BeFwU
nNZXB1jr6pIIwR9Sluh6d7lwmIwihytVRkZz7pE0SGPO+0MW91ujLm4e3rv/skypPf7DUhc+TzG4
d1At4dQ9WOJLeLNpvANOPGfYSnIafjDO2a5IwHBEbT41zYYZJ/O9pil6yLnbdSOwZKXqjKfmFtnk
kNTnNpUVTuXDwTAyDqV44fxMWbkvYzu6hBerg6hUQ1bOu8+8ho5WRVADrZTeZ2MN4j0Zm4n6Hbk+
rihX+3BoaUGYcpnk0LawpWHcU6TZVaODmPyGUznzRcg5EQ3hOV0GoZWROLKSDJfQP54cctI9jMoQ
u2uhJRW8KTTIpdaZ1XB3eO/WPxHiEkOOHh9J1RZ27TJvODSU2YKaSScHbxSyRukSlyH65pT50vuZ
IHoprf9YPrG3a3O99s3TMLXKJXXLm2nroZZQvRDe0zFaWoZMJD075JywBwHgzIbw4L+O9ZLxdu4i
5mqT5MfViult9TabwRCmcJJc/SC39bXR9ThefMaNaBNJE9qxRb76W5C33qPOAdEamwJagUZATntq
FGfZFD7j46BqCKWD5hQf5SNJFNynvV7Q8CkV9VTosoJ/sAu/4zcUJgOLp8Mls5igKpCuqp4hYMrt
aNqZOpGK+QyX9+Hcz/zHQl2LCUMI2vWpTqweRouVaL7kpAY7a2PEIxYYVeBKYGxa8ZnqWlnrDKBB
8OBUmxWXzoqFoH942InOhGWWAQcs6uZ67HUCqGt0xgQ3Me+WDDUOJUNcS7h+aiOb3p0SdKbF8Vo/
WDl8rmAOznRHqwSSGwIxD4UOy/GA4ZX3f2DU4aEhBStHDmM/JtuFuWWd/Yofh7ZVBTq138n+kYUm
mGdqJlWVvecxceM4WGQx5HpLkYoe+PC2BTHeV1PspwaX9zbEeS/ay/tzgsqVwV1p7kvEieEy7xPm
vnSRa/BYruetlDOze3GPm7A3LYrgAwq8cveNRO46q6TD9XfK3tNJHoCO6q5a8pLfLkw9t7zjd65W
ZU6NagvQnzi8U7b3B3YttklloCpZ2ni/XtIrBwCSM8omFPKY8aWvntQyE0L+L+C67ZWGdMpqO7cG
l1kfBDX658n5iFj7bx/Ei+RUGHRSBRWDKVw2kOjwNX+LPRUZHkeGPIAa82HOpe45TDdLQAc1Qnz7
R18mPfFWF1x5E0VB2uYa/Bq+FvnLH3TmvGdw5pQlluEFqQidodL+n5yMSdxw6KCW+RO9cLBK0ZBF
U+chuMTbq4mJi9JGPUwbmbQqLrSX/a4vsp0WH8XOq/D3/Ux3Msdbx1YsGeSdyTFfvCvuhCye
`protect end_protected
