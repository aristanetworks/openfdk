--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   duplicate
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
bQ6JWLR3pzfaKPkmy/5lggeLjWr5+MJN2Vu5UMzC9eU2pTmzcttKK371Eq6lo65D+1OklQEY4Oof
EzHx6kVoCK8UwwD83ftoEiPK2BWpYV196OCaEGl36bmEVXIsmgrw0Jog+m+qvvtYe+fc6cbHysjh
XN6oqUuhxEaGpJ+d1mVGRbwdfYakxmrSUcbhSRmVWMrKb0Qkdsjwwm4gYo636c1S2k9z1oe/p5/L
kczhGNSrLKJs3bkSscUxhrwcbcaNC6GetkRpVyzWTpu6PtVzTLeqMSi4nKpCnp7LyjfLhBTA/enj
uK5GubReKNC4hDLRH3Go8HZG4L6hAWOcXoIG4A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="EaLQSpw31rKIavzDTQ1cHAShYBnJvyweFD6395Dv6OA="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
Y9b5+UGVaGfqoP7b61sbRCmxb5Xoqxkf9XGH3HP7bI74LNQ+NZKC2X+tBIwu6sCovByOHsbmkYp8
BmLCNV7TiDYQXlGEhAw8Qc0luA0AL3q2g1NNlrzrN6H7EafTw/9dZG9expg3PRseZtcbgfnPqL3+
oMy5RXtkgNcH+e74Fg4gz3WUYpQNd86nRgjgQL6AFleaeR62WKGo5n854cj0BZqDmjLrebEHq5Q6
VeYFpxLtLVynOHRVnOCypF5bgsiExWJ/Woxd3bI93ff2qMToaYUWlx8p3Cb3xHcDZPqhUlkGnpnZ
TJH+XU27rAVq5zUe0PWgX4QpAMz6itGesc3yfA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="89wyHKzmu9DvGTqK8uHVRVRvw1OokC3NURcqX1eFG70="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22544)
`protect data_block
GbJQrOuNm7ZiLfqLCDoVyA4+3gpvEJ/oPRh/z1Wi2436Tl0aFBXvR7XU/2sDA4r4WeUqnDVMrPca
pSx4RK+SCNZL3SSvR27sThR00/QdBaHsk93O43nqKJtlWivWt1NzKMMcOBsNm1TGIjGd5PvoAbHj
VErQcvbOzwATQTv2xOjeqf0Z0xl6PA19K93gU4Ybd10IeI1M9FrhBLJfp0Z0ux0nAq3UQiOar4bo
iBRzcUMNfuBIqD+1VOYaRkNL9C/OmmszoGFihO6bVqtw+yuZw0hPW54fV7ubpUk1txfwZkEZpgoc
Ee6hkyxtU99ug+9XvVpaZ+rW/WXi4BSBARa5ByDSMljHK8rn4Uxb0CdR6KJdiPS9rkv0GUBw1qo5
jgOraK+s7M9jq17yboKDhLdCofXUA2KB/iChbqBQ7oKBidwxrBLVaKIsj6XYRBsYoWBKHvFhwcuO
7wBuWmXkjXeWBWX51a0MfIXE2k2XaF2CSCg92e01T9vcwcjM22mm+VcoOq7GgpARBUZ42log/BaM
qPHsWvhr9KLQ17akCiwW5/rA1bwOJwVwkVVX0CiVA7dyIn2zgJXaytD0twDq7cIfLYpFkAbRAIpD
ZITdUo/9Fw5rcqHHvqEHC14N87B1kKxMwOcVQqr78fq/6nghvFBRaZUeFlOGp9XVpb4V0r2QGofG
7WkflJPPrjMRyNYmxAB51FCqANGkbj/K+ZGH1PMoP0tfmvCkWnhg04V8Ap+bB7oyhbn+YHprklHq
52fICGM8JiNLrIygwZRrSXb2Mv+uHzR6n46wgGURrjcEk20GxNex4Hp4U+9uiksDxlTAoospFPwA
/V0TXzUkfOWtwAwGZCxtEI21aeX8etmUbQE5XeSHCTzBnRIBpjoPkOu9PjiztAawdenvtdTXsZG0
hAffQTXm/AuS40VeWC2qto/F/EPzapSs6CBkxI+RajXwWdckQNiCTa9EH/nMOpC00mZhvMiwuCEM
+SBck3k4/y/yJApig4i8IsrEDpKbn6ORKwuoG5vjYMV/JVfhXOqPA1Rp5BMuIIbpwjWNFS8SLL8G
gNmghkyHfp+QWDJTG3VDQPlJGbnk/T2KAfQDCNmPXg+7stOIfNuw/cqEjLhx/pJlZlQRwGBCwqPt
/zV6jb8P5XJ/e74p8sIcc/LL2DC7mIZEXcnta+aAgqE7c0svkIIuisIDjBrjPOHI3k5cp5L5Kv87
1dzSNFpFTH1hIqJIUlyRUj3Ok4HMl3f+vbSd1AVHahZllpW2p+GVkuN7Wyh35ZtFej5XSyTun6v9
LzdoJbfECWjqXEokjwtaJYN72TBVh+6hA+wrnR4c4O8jNiEt2Z9IvVRUyg9u/mjvxGBvHEVH+Hag
0Xo6xr2D09HBLePHXo+xwalhzGaItq4eBX7g/s79Kb/TzeodrF6ewgnElWjIdnh2ApogpD0W4yry
YHz6Ng9J79rVMJOPJWdObXKiA62x6vGLyMJ6Jff3RMTBGX1wTxAl6eM2YQjOIslEo5u+oUlayQfc
HqWB8RhragDchUeoJdzv5BW0RUC+U0LY8n9rUbPq3F0YHNEIULRJ7fp5kg1EddS6SKLSxxFmP3MG
71VixB39eVs9kVbQyekcOr4d1LAcf9LqDUcZZVG1Gwa1FVm3SvFJI9iqGmZ48MVG/sR0UbVoECkc
d8L7DwaJL36gyBQiY0rWlZs7RxMi0DgCrtgSzYv0ztCjQpTCMN5XeJx7ot7Cg87bF1FvbE24MW3n
CvzEpqtNn92SEslcDbxBhDhQNaQgPhztUg8vsi+uNT3rU9UMW+4c5eLn5vIia/nQPBqwZ/wSiG92
mg4JbCR0nF3Q+Oqf5ymNuq+YkSOMIsMh/UxGxA8ckSXvFRh+cyd4Nh4i0g5TZ5GfRB2YcUsao1s8
n1VJpbRdvTkzTMOu5NSAD8feK2YJjvgpz217Kcg6jCuBLtLBQzVZRrJMN1ubUsFHxe3c4RS1bCsC
XF51A3rr7zzqq7lP2wnUj+7/BE3v3q1sSb5o6IvCOdTUcS4LPeOWnncjE8NGUZLy6yUvOU1khxy/
d017z0InYpE11VmAfP7am8lmEyaF82+oRTqB4v8mjAYa1EvvdIXfd7gzSfn3tYXBod67iODgJCtG
TBoYiQbT1grSXv5RpiYdqIGgYULAQUexsyOhe9MZrRZi3clyaHEH8wglsZpo6/71CjCfCycCIinn
sirUVNkWmRKRzj87SIhm6vbPSum2YslWc0Dbwc1JdFALbpIVnrMNU0M+ezIiCo5kilzDWTzGgt8r
TNBfadvlsO3R7Nwd9riIY5/AyNIHM6r9nL3BvsRYhosfBeB9JadQ00lfAXUBdwGIoTYpRdyZVT7I
2tn22+VDHeiNHpTFX3RN9djFDvHCO4zs0aWiO/m4qpCEtRYOp7ukETB4xcDXchKmFGMZ9KLWao3g
ainrKsrIS7Mp3cQtrOn4Dk8mA0N7nn0jnHsfTWZpxq8jCMw5sU00FJ3r2kAOp0lKg0/eMnJfy9SS
kY1lvmRWAWqJGA0sCoeL0Ytk4bPnWtqnIVeAIVO162CZJO3PQpMXiin8VMTcqaFvbSdZdKxvBynu
bjY7lb8u8cOPEmnFBiPeKyUx72O6es8j3GAqt5l/ZZEr3tArGRtIH/4EnX4zCh1kw/3KXxwyXGvb
krN+RQFln9j+kdPxNUarVI54TKwlRnbD8mm8zuRcANEsDwLK+ZWQNsG/lYDbxM0euKkzlkX8aZrW
+T8d4rNPTnQL6LwdK3RXG6MkTVVfYgPoaPs0xY03YQFCDsHakd1zR/8RBcUAKlfbwhKynCLVhDl5
lOGPcWyX4Slx/9ImXhuUUhqEfoIXCZXybjOvuH1Z9TYAJCqKJBOS3DDuNvPxQoVNihYkY2VQGla3
uLyhwE77QJJ+UbaBX8uEIoLygy9cgXSWn8DAGO4PKWxsFSeugm4ATmhZVVqYtB6yyYh4J3n28PS8
KpkWG4MxZBHnv9pMXpKF0BhlyqHIPW1YKKGYkNfFYzl0I6A1H1qFHZGYDErbq4VSZk1BjRKCxpel
TypvSVUkAPa2w332YxDEKY3/rYVnHc0wT3iw20UnyPuCPe+g25LNxXQ8pqlenPuHwS3eGJOxXKpO
v5GQU6zW0OjybvDUYhKz5cqBqyXC+1fEWmvgtsce//oG3rGJdfv9XPqvCG+x4BHuVV3/4eO00rya
sVKYEdD/dY5ohq0m2Mv7R4rqBG3gtnOJZKGpcOirmJs71ZDaKLLEobKha1S4qDoFRHT8UjB6tTvB
Uo9m5xn4jtwptBUJI6vd7CG9Bx/B3Vr903mU9CMjxMPQmPTILT5cS0YnL+5crVqFuEFweXocDm7Z
zcmPo8X6ds/kZ5+R9Zn66miorT0Hn3NrWHtBuTV42/n/MEvUmBO35JGN6a8d+IuoLrOXfnjrMQgx
eMtdgFDetDAsGys+RXzb2Hws9GgaEABQBgOJ4SPn8zoKkkQrJfUqCrpOc/Kk/zHlwdMgBrZbzFxQ
pKTLHS8RMiB9IcRFdnNSEvHLIqjegqsW5G75KkfkyDlGDh30dY42b99P15v/zAKZdoSXipt4byEw
rdy1HBVV8pGRFmVKIC34YMVz/wBToKxU6HAZqKDPada1QbSxY/IvpCwbwrsFkAEsE/wo0kQRReS9
ae7lncT4lW+uJJHjWYd0Ygq861ZJiM2rfjTnViYpUHhGfzi8O0AdUk4E1s6/OVpZd07mjD7c5h3N
Jov1XxbTmTkWR3xlNf3QQusD8w/sqULLo90bVwPpKHWPu3CM7LDAZdfGG0A3pg6iod+2DvM0Hsr/
YJG3MDu/xrauV4RXch0lmFvQX3HWdKv9nbpmi9nF31akEoZzSl6n3iE0QjJyu8yLIDY4TZOEz+5e
H4NqwKMUzvsP4NoVs9+B5HfghBITVi6Fofx2C6zOuzqxJg6RzKCQR6JEdrPCK3+BbFxfla4LHMei
FCCLqXeV7b2B3h8hcC4mlz6vg9GLJJ6n/5Yy6LfqOELpAeMzqe2ex3DD8E39QDJeexXmSz1RIqVa
TQSOouJ/O8r11muW7UeD8z8ogQkDCtrFyo1tCbgGRpO9zJuSpMcLgvQpngO4gGsVo39TI0NblzzM
dayEx+1+qWEKs/yItAqo0QM6kqbp9RDx7F3NhgEPbxWmJ39sh+Za1JAA5rYR2HRGAx31nU/69JD0
uXNV1iAwWC66ZMb4spSuP/fcOTjsTD2Mer/Oxu36YzGtYf0zW4wQRRxAsFgaLCNecbG6Ew35R0mH
HKFeqes3AnIfL2XU9LnqstGfSVP4hoX+g3+s/wY7Jd4pJHcUUleBZOSfzM0hBDdZcVtPgvLF/6Vw
GGdcFWoRjArY/EITGsU7AUXBOL4RROBPR0fuKPTgdDtR/3XCAEgLSpF1yoFHzpJ97L3eLO9CFFhI
RswZMn+Rjv8UCNFEnMRZETvH9JKdtsk59FSyDAb0/QXj7fvwk7quRbNp61tUU/uAddOb9f7iw1pW
eYVHSEkodgiwX3KuE509DhK9KsgcbLlGdWHsqEf6TfnsSDFf6ZysBw3WGzbYp7gBKuN79/zqMF48
y/nv+iJ3rDpt0SBQ22pPy4oKG9ghGB4GytVwqLU56AYWy49q0HHfudD4t1yaJLqJLhEAOaxj54Vf
XQNPYXLhPxnFN7A0yjQHiw+LHTI9eszMpWYpFUyS1Gr6tOU+IPeY5fdPnrGgwOHxsVOLrtLFYLmO
Nu+ybWUJ9sHVBKcH9h62jnywGO5N2xSHxf2US/hwVEC9WB/xj0cPy5e+N/daf57S+ttmFSDbpHpl
b9KilTYT97Z+3zThP5qiA5B5VgtW9KoNVODvwr2GZVM/LzoDeU+wKuYQidAOzJw81Ilpk1/n5lPy
g1+Jd8FzuhZGFGzhaKLMsNgu687uB3sA82tVWasmnAXq1wFfmrLzjGmOrxqiU1R4k4YAiAmxnDLt
78f7KrciSRPOKB1q1upka35WGBX8uiy3SF3WGALojg8k5XhCsS8MBPN5/efEpmyOmIngRhHaiSHr
ASrcvkUlCWpWOsb97P+icRQZ6aAvt+s5Y0XTALuSmhWi3yNAGkEXIK2p5NVJ66z5seBhsV+ULqLG
BBzzR4r1dsO5YNh4bqkuzN3+Uv1FS0nq53ao0lEoOOgD1YTSY0X1er7Z5u45jCA62AthTfJKahbz
jSBT/kz9PByIloY+Z/8HjEACjdqAJpBa4W81cqYX0VfBocLwKQftOHC+QKQQ9S3XOv2urjn8ZNQt
gIZdGyYfQATeAxg8mzmNO/O000y9rWh3HZlajzPOCP8gKm+0LmoSoLpd0pzpu5maE9QjgZOlZa7X
7bZWTogREJK9E5P+g2AxWZoizJgU3llD3srUd5ivd/U5H/14bQjOza2n6ukneXBBD0yjF72ZLzUk
M7y3WWqHZxMCm7FTWR4qVHcJRHR8W03M/937OzM2hJdiGaR2lq23FckgXLKFxgQfATcuBfiB+6Q/
6pr2I1paUHvnE1cy78BVutOGyK0yksqy8YHl7IaUnE9XDLyzrDSz6ChA4Db2quO/RP8tF8/Nm34B
BQVkfOFD2FvyzNuQxefeUHlNnBR0b1mHOcSkevbfWEGfSS+SZVZkeaxF7gmGElP36rmcb5r/8oUN
1bCaoZg/atyAdajbM7B7WWVNBBI1W3rS7IvBxrkZeCdm9IwGH8YTkpkNPwwSyVnxAvhf/mcu3h8g
6GPONh3DQRKdr4fF5AXhgNJhajedt7rEjHWLOcIyRdyx4EBGHraEAFgjk8BWmlIBBgkAwLKVkVm6
rCTGdMPDNs41Jtc59ZCLlJOJQrT3uKXGl9hpVyYT2+gzqkjJhghLgxiyL7oEE3qZh4S+MH+ThKyh
z72PNppjxxL18H2bu/i5n/lfERWzad/1pSWnOuHQJXMIbLJ1VuJ7GGV++OyE1HNUEyaDPEyqA/3t
C8G4yagGvEZc/ZnTCdR25O6C9ey6BJVyxV5Zq8/JqRZHggdDk2XxMnAR2FXBJkRpXn157UBQDVBj
x13wKm4xo9MV2pFqKW1ORU5kLbcvuy67Wxxd1Ce0qqLJVVJJcyIT3IzEl8TEkAKAi38Qyd0AMgFV
1ZGWQYM5ymK3/tm4SxWBn0fCKI8eVe1Ui3RrjhHTqttQg+CvNpkhmoRiD4QhAwB+TwVNEu/ZA8Jb
SgOPL9+5fqORfD3Fdmz94JO3wVN1Se/+T2cRZv4U1+2V/2w0j7Q+7d2LSRt4EcFcRSdhHei6yKZZ
jHziLCG2E/FAdbAmms4vQDhyMNgtWOjfxoYa7w3VpdNqFA1bpdM6cTyPqHBKJCkfEKauP05C2los
D4o0axYnViZhB7K3cyhcwS6m96mD+FxDACTK15n0gOkicCaFL/K0+7Ap40z2709xOyjMzsPMNKnX
LYqLZZpTkSoyzsl8416O4tKyIPHRtIOjO7Uc4FDHe9a8mVh6OQarWwTjd1SJKNSNNYn8QTceia5B
owfEM2clmdohkdJjs9UoolVjyyUpwgpfbdqF7/ckFoTltLwpLmTXLEEYk+/19XG//S6Kmpt5Z0GW
3889peI+A5w3o7Y/kaAG2tl6qOGu5qW8+xvngtDZO6So6TpXj5dfGUNdCukYRaBylmBR99lonB8j
SDX38vG++LAS7VKrG/9uSgY0WMhNA8Ubo6kUqOYe1y4Q6H9QK5MQqdJkhWWStA+cO3b5OYmgiPP0
+nZ3DyIr+L2t6TC5TwxvqIzcCqOYyERMxsFKRDMFgzOKracN4yaS5hvG1+olAgeNEy1k0tePZiVw
8xK8DaBlsk3STKMsEfdHl6GFEI4DEpTv1Kl1lelJREsqblAJRaU83Uovp9pdyAzy9ATEgZy3q3aT
RLlaWudFgt0Zg1u2BpObJZw9UkqvGJBaGPJq6oXt/f1GzvmEnFuvKKvzZXoUYX9kyK3xcUf1Bseh
t5MNp41zqCrEWZRrCbrtgXGC2u3hyBMRldQ7pJZDPYBWS8M9/h/zt3bpx2ZBobtr70/6d1XohO0u
ZFUkdMP5i34l/8Z7UlFV6idB+uXjyxWgM+nZC4GUhnk43BMx/TEz8ZYToipnCIThKZO8qFkp+njI
QkCV4jp9EfZ9gibGgh3eQ/MtwvZqvhACwnQa2rlx8jeZp065C6V0+NOQSD8Gp6CFoQHjSE0IM/8m
MrvRoH4ohVM/3LWRJU6L+thWS4hsqZUiZhFPcsm4jTY1wjhJKR/RQSz7FYlZ4ZCFVZcMq1fx8XMN
dNfliyZ+Ht97bcJf0NLgDO1KjVQK356Os+r1VgMpflZW43Rtgmxuh1Mg2ws4nCTTOHg25XuNJOWz
PLPzsOudnqrBtIYedI8yA+Oo6J2yJOWXAZ1fWAld6YpS44Cy2A7OmOxXxPgTnLIqUOn6iAXu//ho
ZfnMjHJjatuh6AOpRFNAe8fKeI+xI0Ke5+0u+CAeAcpkhOJDnqZlKiWBAFcUIL/3milnLJojT+/4
4ckSS0ToiFbtevleVg2pdPXxuw8vZLDz3jroKxxVzVl1I2Odxp4X3pEmW3RzTzp6aCpHIoK0uiRn
zU9Gdkj25hkGHFX98z5Gbk5ocRRo+M0qOeU5VaX9/G/zDGX5OT3QNfM2NyCTthQzotLzSdSvJI/5
DibbYkWCuBYkdnFDGnPHAvAdgWna5+6kd9ZsBIJcUrE4lbdtcT3IoeeTxBSk7DYB9L2KnR1VOKxz
uWuJjZ3dG/vdPwzWjALZBVjJ9nxjHmM50uLM2bVCJrCvfjqcI4Qj3U4nOaqrVB1xENXy4MK6EDru
yeW7C1emHXCCl9kNB+Pa+oCfmcwgbH+mDGb8iVsH10O+WiiqUJ8ubV4FEsXpn+fixEci2xPZ3tTR
DlVLdaal/KFNMD9KMIOdZaXbeZvrC13TzfhwGLRnr9290q5N32LMsmmOd8+PO9UUuFXWuSr7wMK5
kJc0av33W6k6gq3yR4ScyhuFGs8iikNRZW1sMB5BvRZDnEWTZEIViljGpng62q/L3zWKsSKiwlg3
b4NvFxwb8FnxlNmLhXwIPQUmd1CsYMnPwEvM6ZCTM1Ghg8Weet7aXKO9UzUlUskSMuOirLu/8UNU
O1OqvNoqs/o7AbveZs5P8DviqvwDtJ0cxPe8Ub1F+Lqz6rMyqdD4/Pza9tEc5r3hjPMFNWj2ktXr
RbCHLU3PrcQwnJghnIiBlHjoXefe4oMtqYC4qhJvCDA0DfoGOmiIdFs4FwUaH640kULHoowIBwso
ezSxjm7z25DHAu5ptMxOAncl9s5lD0o5fRkA8yM2CK1XXlzzcUZpNBZJgzkjBY7wI9YwtEPlDBbm
4qn6WzUbMk+RAw1+eJMDQV3FnTNowETjyBVv5a5NljOgZTnddAovjMiaFcDtyIaP1Ow+d6JynKLL
evEiolv/3F0hbmdXiHYvXX3k+MDMEwgUo1WsktaLOmA1mb3GBVFkLbdX5+i0j+2HE5cnEqPs97Lc
Mqeq1hYJY2T6jheDxUySKiuI86JappAtAEg6jDKJXpgPdSBJvm/PoSCGXmWKU0jOZj58l+J8ij+/
luFMHxSxJbXsb3nwy9eQp7rnYH8IOSJIP1aGcFgpaUpopbJtkUrowYBRCameQx80z2vVc91a/9fQ
D50XINeApwCuNpuD5BuyUxxM/U5wevQ4gWJdltxNed2pi9+eGHZ5Yrz4VZKDhW4/of+az2owQUc2
ei1RA6YqU+GC0g8kvVJWK+C1ZTHNQgPr+Miqd8URx9ywrdRvuZ2l+zFXvF46tlPrpNjuhCjTvmw4
g8+ZXvsNNdtP2nvHX7LD6ZbDKvFWshA0QAHzP+Ow/mcfwqzXpTcZKxEEtp1phjkpyLQokWS1mOdf
kgRcDd4jxWFxhsIUKYMacIc18rL6DVBg57gaujyTY32+gwlkO76rqJc1anzYBRzoMOgqYEI/fIqN
yDF5ACL/SwNuiivqT+OYScq+lm6nKRR6Z7uo6u7apDvjx80tQLO2umtJprAyLwkY3WAo0hvpiwmQ
IlRu3qmE0NNKcq1Hz3Cipdqz5PZPSu0bilvfbSQN7TxR8Wpn/2IgMOHGH8UsOZP0rVEuAysF1kOd
YHrJdz9K3cYBVJwPzkd1lfe5MEewr6CDJ7mEf5kQ+GJ+X1YYmCMxpTOycrOJzmcYqkZnOc4A3o80
JMjtIs1npQa0662okWwQ6OzuVOVMepy/vMyYFbeRK3IpTXbDXdqQ8ZiEJS1PqbRdM31dDZf+ndtL
BZ0c/Li9nr6YqvzXVVoiyHyqVJvT080u+8ney0lTeN4HjOw/7r+Tou6BVZWwEPCUk5KxZXu5PqO+
kWdPUn10u3zi+i96peSekz/WBhk0eJ38tnQQhrf10JzUxgfOwMz1iG9igAIDx9iHejF2j+p7fClG
qz05XIX+D4PE2747Z+t3neCLNF7/2h8zs0miM43ktxUQGCqVyyZEpwnTS3vFwpPopSWO1XuSHaJB
vRAYTavnihCT5JVTmiV1VPZidMGMb8MflknNc5yziCGRDN3MNCNcDGr1UL5ydh1VUhl8Tc2n8uMT
WcIMGGlCin+4qb76KKWQSv6Qn83fMjiII5iSgEvdlvl74aKWyOyWqo7wNfGzTNh1tY0xSq9qC6e5
mcUbPWdu9RaseSktxhdehmptm/NARU0QMb+pNVkd+Xh+GRvWOeQrLdsZfpm1t87GTiBpMKqNFztF
ec5TAFE4C0pTkZl7Ta44K/rTjnB/87ILijdqIN0Y5ig8UBwqbIyU8LnelF4J30/FAihAwihzDht9
2qiDyH3X/zbOcFv3JH6X2MuHlSJR0yOvb4FJuv/Ep3wR4S2kpnggaGLkTpI6n3ULWkLuuesQAEcr
GR712PHgCzJNvILJe+G9SeIR8iAhPIEj+8qyBPiyIKI9IyBGsXnB9pJLJRL4t/G+9f39mH1+ZOVw
DluKKILB6sP4PD4vrvdBh6VGINtW8fzI+/0VpA5uvnNY5RNNBz9L4IJ5N+7+B7QMZbHsQoNSN7dF
Y3MTLZV8QruBqjn2tslRN/+viPfz9sw3JDRr5V1X8FeuYHYhPQ5bOG9Bpat6RF8q0wbFfu4krE5q
saec3ZtfPOaCx6PXLojiasbcvDqAA6tZmCTonBHpdDAK2UQwWoCef/w20C7a/JAWcAW2kYtxpxsO
NoFPGZLBUiT/QtSuqv00bhi52Z2z2/u1Nr2TZaQfddSS9sbSaREWtbO0IBsABbNgtXWiwj1UEH7K
7pMevDg6hHupBvgeJ37lhkSwKHq4ChJVsIvTaXwVXjytLEwy7pzmoqRbAHhGWVLi6zsHx0P9cZix
AHc71m6xYUOLdBnBGyIKcdvD1aRJ6JL4j9k8p7zoKAAnyTtWUdTpDIIqRk9lvR+qvWIp6zbKo6vr
pw6k0RRGWW5rocpYACUOT40zT19zo4oQ/kMV85TQfe4D/s+MnYdfq0VeSj5pCAlwLTWZWy3aMIoi
btBms/bxP+Rj5qHgGtY1/N4EGp19raL81VRxntLZGHlqGlxPQFxq+NvPJnIHzJYV6Ek3rGZPTGYC
J4OkGovhy2aaaqYG+7S2Rx1Hjts4bawetTcvqeiT8hIbYmo6GuGEUc9w8TdHiX6fvwk8kdfBumk4
cx0iZ2A0hm/i0PzMm3DTnLPxehDknhAQqdKqv9BiaDL6IyMmlkc4yiux6CTsKajcWOvfpxd956MV
BuQpKwuFpW1cdvgyi/P8999gTu908nOSO+ydjkqvJ7ediCDmcU2COQ1xEh/Jpmo/36oOI6uibq01
+IpOjgfZ+tykuWJLRW25zTUFQe0otni8Z8/xWiFe3opDw0KRen6eZXLo8dNmmPKJqnIGJgnWBNuU
q4eP+BpJWvGTyAXjWnZPcH9C/ZEfruEzRLpiE8lVuSIe9Hl6EU2p40r6JCqW1S/WUv4wanmrlGfF
rXDbJK8PC0cjJP+9yFKYsRx/h3LU/19lrKeVJ8LpyaNvGmUMJ+Bu7GTz6NxUJjNfcdddetSIJ3c3
tlRE8im0aOscBJ1WCnO4eiN5sU44TPzd4Wq1C+NetJOv5DVsLzU4iHpukLkRfLcf378CeW/HXUSL
9HzWvsysoox8jQvqzV0aEz9ha28o9Gsbqb2cQxf+/zW/BpS9XfjkAdX4ZU/I/xS26D2MUG9BmF10
0ORx1Wc4LyWeFXgxPk7TQZpRuvIMBub4HGwJcHqyzaMGbyKC/btkm/Mx2RuDBNU5MnnTizwiL671
7PvWuDDl+toxsGvGVN7N8+YOTpo69Ur9ujxUCBNGQ2ervcKVIxqKmcxhRtMs1eTkzXabkbJvozQe
ompW98KqS9uXJSB3nbXllFQeNZ1pljsfvbXw0mAXLLAMavPXD4CFXkYKdW5POQJB3mKv2tEidjsB
NoidEMUfAgjkXjJqtFv1KJlpgQ0X9PuJ2HU3pHopPbbIyFiTAbCb3GGri8nveHNxQ7GzpZF4qfmW
KKA6C054dUvWdsI7E8ZZPSNcDoioh1EtEhAPcnekzl/qL5zD3L8rO3RZ+lkAHLfu7tnKZotVYTKS
AnkLsMRWJY7fJr3dhOoIJh8ditZklaUONdoeWzaKcW2Hm3OsLsqcw1A68aPKc+Wc3n0tXTSUdhk+
vex9O8/gFdhmAWbJnVGLbEUBu4r3zZupYjXaogaOaA+8yoFCB8dfi98tV6AkE8f/9E4kMXrarsHI
LBUSFnfSsdkKN/a8Doo1fyK6lKW5YoxryI6B57IEb7xn0LTzsbhtAQahD+wyxVLQdePWP22v6BNw
rX7/zUblLD4lv8Hh5b3v1bbmXFrVTyIwZBtsxFtVzbHdjy6DRhzA6FWwjsAm4UMBaQWV/RXiXsaJ
J3TUwdqfUyN8sXNJOgYUCcHnB+rj9HdNAXpjHnlYQ4H8n1QnXf6FpeMhl9lIwWlcMsfMSQHybDDk
TqjM0K87EaFJOmV8H4IzWZWDjHEXF2/XNJyot/tL7nGm6P4hPiPCMpwyMl6MK3Ep62alkbw/4AgE
bofs8m4d19JBcOdsCwJ/ThcLEZSaNiMa6vLnb+4tTcdh/Rw6kRfDZwk/JvGjfqrxuS6DEjKTzgkR
vFVGkJfVN3iogs5RuWSiy1QMnvCDUWr4N68CpT1i5zj858uq+gjPF05240UZQwwtXJ3ocQbBuqz2
hLT/VE1tyITb1QFmfjmqKhp3/WdMfhqdH3MQXr7hxZcRTfh9MI0jJKrLqQ8BX/Q/RLXg/1BUeDRi
EzCt2TPBlIlZXlpq7ZRlh7QXi0IDXCtYUaApl2s5UmNHQHoLCPjyCpoWUCeG0UIp0Wa5AZKPY+Re
sYGZZ0Cqo/mBqvg/nLEm776CIelRzUYcMPi0nXWC43usGxu/NkZIGrVsvh7ob0Br+9uE+MWVjeve
nzXtXtig18SzJEcUgASvh12SVDQ5haFimPHYE9Rjf+d8kqOkesSF/xUpqRLLZc38yncQE6+poYI1
7HaffQnbZ/GMEPjHLScqV9i9uoTvLP8RGbaUv97S6FYW/qCsgggnYAcwzqEWJ5t2tgIDgImjba3o
i4X+p4fP6bN4QazE6e+Qf8Dh5wsLf77A+KEyufgrkZZ6e9VIwUW3YE5QlQsinFs91thDH157m5Cz
KM2hl0duHm1Hk1Y482PniODtodUeMa2qWT3rm0EGH9UwESj+ftY18PgL69LF+06nC5nNylDEwCbj
ZjTuTiFolaIaf/2VvmM14CQDMsBOuuN0t8vwAfeylyivRhcTyWRo6t4mdVb9K6Qru6iRy6OQ6QCA
IH1BooQykgf9Ws+JxEqcGjKanr7BqFC2gQKN5vkldZ4PAMa9h4hxdL7QoGyAJXmZueYdh91yodKZ
mo52UEUO1+9eL2Qj8lgU6R3OO+BIvN50XEfl4QkrVhNtXEtw31ykxBB1VxuE0Z4KLqkSHifzDImz
TGTi/X0QmcGPMTfQdDJXR08PcHurF8vIm204iRNvuTi7jTaTfUO/o43xBbGlhixWjtqIH+JI+BsO
ijsF79FDUs1bmZrPtV+PpYnDUsgb4Ck/JVZ+dU3g890FSRa12Zkh+w1HXBMXG0B6PrprdhS67mZa
jO/1fXauP8sZBbRJB4xsLxXbfAJenvQqLBvu7xWpzPtlSKetnR/BvfTsLB4L/UrrbObWN4n9kdG0
t8CGzIdeWMxLzE9IgLwEhpP4485FtEnMzkyNqskPgJC90LyPt8Y9uPKoEmyhXxXnUOq7FwWQ4h4E
IyWEAtDSdPz/I/dm7yfo0KfKDseVX3vfO41KglNMAkHbYodQpU9Ihzw5PTP07tc3cho7AItemF6S
2Sfks9OFlPJCWMzhrfzj2mInDO+UvDPI2CAMC87Evz/AwZupb9j4I6nUS2t4+oV3Bb+jwBHwTKK/
3UHlkdxmqKVFt+gmeAqc7LsqEKkk9LN4/NJuty7m9MY/DGsY36b2s99UgdUY0bgK7Mh6hzwV3MsX
C+x/wQkyjpmRpva5Kp9kC4eyu98+tGbmMUlgU/Ba3A1n8vuHVlRYy4YpFJ6ElsCujbihvAYf9Wsx
unZXD7Lue7dC4MzcXjhQEvRLKfhYvgsYHN2dyD/nNAHXjext0ZxIkJMleMQf3wKB2n9EBgTo1EhW
lFwzwcdtqpDjyuo88z7/I4mhovPYU5zubNDVvkJFLScbxTXVHG4dxM5m8uk4MJ7oOF0jbRuvkEiL
Zv/pH3K6WVcsNRNTKJfP46UUuQDVzQIPe8aSh6yMlfShYJj6YojWec0LS6UdPXeqLbCJwrl1456w
8caqda3ufuHF2lRWlugcgKqMV1hCpKX0o0zklrtZIHASkuzxmU53QzJUu+LJINAWFlqc/o6P53yv
H1a6AMIjtkp9D78yRlWaReelpHMEIl1mCE0A0LY8Er/5DWTFH2J16m3pcWSZTJ6+hjiwABym6NcU
qanhO5he5XebVMHTWr8ss2pnFsAwTZrxuxY+EPoH9m5iniaToQM6RkHRBf8ymrm4f/+3YFR0U8A7
v/XlMgC8xmcHzqBRiWEGmVNjdDoP4QyYloEnKPOjW2K2w2sjLbrSHaDmNNthr9/98wD3wQIuJzj7
OIX3dOi1dmB8/niLlBP3Dbm3y8Qic4tifp9nUrOGzv8OqyK3g3BQEorUPDRQhncfuZjCX9Uztpvz
MQWQozpUHrrH6LT5sSwXU5dKuPwHvHnqmCJ+aFRvoygqI+LCdk5WIwztICf3vpjEMawZVLJUnOv3
BvcYFNrAafPoaEHNYVWMmzggMNHmHYRUMupyGQeJ2bLvW7UTopJoSeIWlEdWeX0K9pSjmb+wQ1q8
dJNC3mrg7b/7UbS38aqBR5AXRYIHHHLr2INbVlb6CpjmgnPfKZAsCWkU2b1ojB6xTxVVt1s7bYew
i+Nf47xjsE6vxHqRN6OqZNQwGUEyFRjxdLTPPipqj4KHR7hqpXWs8ozDo9/sQ98HdnYcHKNWWJZF
pGiJ47vnjNDQDIFs5GXAoti38koQLh5eg/jOsYnEaoTSBwmaTdrbxUdb6Ua45ZBY62GXFh0gtpgO
ijkuuL2KllTdQSCWmk4P2ovS1+0D3dsgkuwq7HBNE1+4bs1Orw8NXcnvlhzNmSJeAhGIzYxBBKTX
YXADYHV385yu2JnoVDNhCyn0NIHC3hru0n4VLf2WKiq4ihWPVNypd9XR3TtNXO/KMSXcvFhrlENb
QzVaf2Qk2SinqeIMsUHJNa6PjNdgKWURlq3In38J2hPkRFFgK06NlUkA0+yXUGy3RYQmjnWoy2k3
j0NlvtIpz1KfBAqJ31v91mFVWwXdFtJ26ABv3uYXSZoil+UIh5wkDfsYRvh6JV8qcRIFjNsl8BYS
ggMVJMq+fa4F7WksxOGygUXSNODPSll3Osr6cxnQI3Ls29NvMhciaKNBBPtP9U00E7HeM33m1nO5
h3fSpMxAzBYV36uHE2NnUU+Pf7gxUPeskdpF0z6IKHYphJvtrfxxZKskHOfQ9glmC1+Lxx5kUNTO
fSsoAjG5eLo+KEHJHHLVjInYEH2DPBAylcUaYqCBb1YbXYoozgSXE7O/AZ3hv42QXM15sx7DDr23
EMOpjHjgJjDow7YFx4Z9B8PUJ38PRczwh0YWG09XxY6bYhvGY5NDdUG9rEupK5FXoSP56oCGcakX
mxFKXQ63S1qvg7mGy5Oz/xQq0wpMOiXtN7lu85GvxpL6aQRBg2NeYOBzpNWLhC2Okyc99QcVu5lG
5uS+pVqd/Y368WkLrLBUAtxKsl19rMCYKr43WUcPDj/sysikIhnrXcobF90WAFrUIl+FSdHiPvCu
CW9Moxr9jrjoxZCUrAKJNu/NUamQyUDDQ9TnOQFA6Ut2q4XyaPqcgjqnkjCcJtc+GuTfAo/ipZuF
KhoVRFrhruZQLmxLi23AZGS2G9GXkwFCqPzMVvbHQqQqQduK/mPFpqXBzTgJIqwXYzmrrY2ppa1Z
OK3KaP3VSKCMtV5p4WxBHaUyrl5nVOtBeUJZ+vXX4aDcb+5qxWpOJ+abGzFHxOqvJXOL5WLbbFhr
k/7Ff+hjdS6vwc4Qrkre7f8+nsp6dslRbYmE9BbeoNGO90T6c7a5BmfjnIPlcqesq3j7Zs7HsOOP
Xl7PAiPLyiUUwsiuCoi9hZBnVZwECLc7D8SjyL3RiB0zkkz+c6h3+J/svFYbZgf6pofVtQyDVmao
JvxftZn2XZ1DucVdz1WzASsVF99wSc60KpUpLpS4GJD4KzXQ2+OHe8oAkGFoO3OBqV24sCrXvuIY
x1S2dYgc6elZoJqhu2c4wUTh8mjIgpDBXPkhvEnID+v/MSVIt8mF+6SAnQiNZi0T6QM2fCm2EoaD
bCh1wBiEYMPIu9MPcgcMzeAbHg6+1t/djhVvfyqMoxZqR4T1vWqcu96d78xcdtO6a60EiSRZJbu4
lbooGC8uvEI4bMkf91yD3BWAo6odaGNAuLf9R5Un6Dvtx0/bspRHGiW0QmFttermAz6Ky1P5LLbc
e1qrz7sbzk6R/gtaaz3jIHT959MwJtWXS1IBahtMLqGDceMMUi4Ps1Yjp7ptWKyC/+1dz7/XM6xF
7WYKf77WOrDrUIRtAmUifSppZhQvUdeUWGNcSzjP/3KNGMHm7l3p4C/OnX9jAr5OCxcrOEu8+jkv
YCPXnNzCAlp+fEJYxCuQVfC6VFBDTHLdbCCMcIGu0zjtpYLrSuphFCwA6TOtRdv6mr4AM9heQEs1
QASocCAKZiSKPr+YkoTdHESsUF1MA0GhTrXj7hZYKZZzfpY6kAJRZFARNRtC9B67rkit0mnKy2ZG
OfBC9Kbi12Z4k9DCam59IeNqcKjyGodQhCp7Q3Uda4O0pJofTL0QnJ8+7fTAxP6hYOqWLypJDBlZ
NQi6rxtdyjEBYZX+28p2tgqRvQ3uzCJEdPDkUaUEjJblDoXYxiOdfSvpMGxMBiunPENRuoU5/44A
9MWV+iJuUtzX5GEt4vLrAOQfQvT3jJSf+YxuRNktfowx/rxda1yv7FzF5q75xDGQ6ZekxCVxHPKd
sLkrFl++QJwNhCBp8VKplHHgFFHag5qyfBSa4JIX+Xj8YHcbcyfxs2Kyiudql/ood8aSfo3xK1y6
NT6TQsGkIjnFKvVKzDnjnCeLaY9M+8tWEZmXs5PpfPkPH0HdT+qKVlm1Hzaxny1akLlMah1+UYLs
uRfVR9Ied9qREl+Lxc7hrX6iViNwLogyPasXaEpW9Nvp0X7Cg+by75hbAnaVtj5oMCC/BZSXpJps
7Ax1gcUcRGGNhL5qdOckw7x2EwbE5zHlvST1mw5QOId3PeBWbbnaboW+0VSIwdNbvRHYOhYMlgXU
lq/rNhRr+wqLNqbT+acmUZ6dQPgSxeISxUVCeapaq8IlXDDYqEkDfAVvBmJiu4GQxrFSxkCqeM7p
i3/t5xl3J/b/hNytmgOZg9bldAN+dK+A3v5tfMz162wVU7rmQ3Z/wN0jppIvh0pJtcjS8eyG+guN
Oc8Hbi3TYKERf2rqvuGOvKuVP1mVDbXNummjjuzJdG4cruF3gyN5MLo1cRmjbd1qldoOcH9zRHEh
Ouk0RLm56v6xxfYVQz9CJcdt2FxLHyZcehpn47iU/QbHWQxbREzyXheVRw3RYcd1cG9InJQOn7V6
Dh+ReuFAeelMyb7+sEYDdvppGDZfCx1JQWRDUgr/kn3SZ57IsQYq8kpZpgFACCrwRIHvjKo+FrYc
+npq12+L7PvWRm+pa+6wZs4wZbBjDHI0Pcwjc4ZjazuTEPoNAZ6wnL7eDpV2gHaP9CYXLFenJFHf
nXjf5DXjtNjB4X+Qbpvy3MgljgbCBhPGaomOhCqf7GPNQWpa+Hi3o6vk+URFEcJ6Ua+EdcAGiWnW
J3DNWd9rx7NTqVyJYVyrzY2GE2XsMlO3eQzhUkuV27753Mx3RXYfEDa52AnG6KaK5bQeVT7ZBtoI
eRdO9fY4+q+UHVTlbO3Qk7qPRRU7Sq2udZtrM2br8A6tnmXh/3EeAeaHohKAi1JK1ZjRzQd7xX7U
u8WVhnckpgO0MZ9DeaAYXB7M1tAFpugeHdEa7MEtJlVT3EUWlRyEPOYPF5qL1iMX0sqtFdJ/gxE4
HCTUGM2fBvbS43RdqJ00mNBWRqG0Q2m223mznuIaexFswMAaUJk7Sgq5/El8VjdH4eK4vhirDEID
nVpW5MN+PJhy8wX6jrO1ibE5xEHj1Wb6G+zFFjvq1J12N2rJ5JzrZgfItDw79L2yAMvPRJwANzyz
fsNvfxtKB6OzOvuleq9QMzQcFQwCmAjR/c0i1GaU92ktcLKAAxPNwyLNTLZ9lAZKLNuWrrGodj2x
Ou7BDZDtyzy1cK3f/683QwieyIe0qLWwUuT4RchTF6mZJRt9ObSN/+EAxwfKqRvHFbBR889XxOv5
PJnib9jip2618xMQB3kFk0vNwOe6C1ESpOPmwJ40pjYywJmAJqT7pup2uCc69JPhYnZABkw7daCJ
ZK81Emp8nudG3MKoqnqYqqv/ART++MO/KMDNJonCXm4hPMZKKjZsoQjP8cEJlEThoXwKogJ9V+q5
zEnCqZqm3I5BCXi8/a1maZc9mCOukKr26c1W3MpfxH5YDEP/fIOALZ+emIF7zyH+E5t8x6GdYSMf
dv35b0OO5ymcoqxh8OtSSMJr6OJX38RGLQwFIwLLwsv0GvrrPtRoQqtR6JJ3qYsvp8tKlmf8Kan+
P8DS3vCB0kik4dyuGB4WYL9YzaKgb2WsgNRkgjGgtx8RQLP9oKRrK+vroc0QMxxO/zEZDhP2Qtjf
KhDm4zfbIr38TUQUYOOR3G9dKzluJWug5lVF9oQjn8GhnCz5u6Kk6fu3J69IDXxa+2aiHnsee2TS
nlsFeGx2M49DMPfjF/wkHkQUWVlXF3IOnx6XnUv+olIfGb5LV9pz0mFn0QsgbJwrsocnyzi+I9Sk
xI8l/OCbhV/fVC0aPvppuoXXCoU4ntrw6bO2jEuD77eeuFQhiHwEWraeJTREgL/k92y/YSLcxznx
iS+av8I6jXs/QfYhHohPTNo7UV2TdjX5jk66MFTUZUaJ8npntTwl8A3oIqTXS2naeX28AK9HciV2
xLId49gG5RtymyarezM91MkpEPl4Wk1HARAbj8UCGC8QcTvDLvhbdOv4PduNDcuagZuxCMUkZl8Q
U+lJfj1+XXRHotvdFat0ONi4XT9lPLsvZFIBECVHznx+0nSuvrBgNTm6xWpvd2z/TJr2KFMGCzAX
nkkNYd8hR3+M2ES1aEVD3e6uGP3hqwZlkfkQavf7gCjmO+PHzOYDNgeeUe6zJEYcAHzWWzz9v798
mKqzE09J2zBXCv3QXSQqF/ze+IBDapNwZ6fcvx+Ni8goBV3C+dM9iW6Kp/FEO2Bia+eTXdDOYuAt
rUnvkOhQ5qNg4OR3bx5rwqFYPRM3NDJD5vxyvh7k9+KSLWHRu3r3SzQxwRNN8gGV/pll1RZJMkvg
6dskYgNKighc2FFRnMciMpWXs2rFnujJhPHjL4KJv/+GrkEgoBRedENVkBftF8tMVKD2ySFqnvfN
I7Wn0HiYnX33m+U3VByzJWHPB2dtLxAWGxTzxWdyslxT81G91uGTpkrUYPbXkQPq5fZMrq+y8oLR
A6MsS+PGGggwcm2+yN/4aoEhhB4r8/FZ0U7BjNG28FR0yLYXJPVbZGF0Ri8lskY1BML4v8hDDVTi
tw7iJ55N1wff9SOQwVh4eH2AXZ8Y+K3Eo2cSWPz72yP69tOd7+9cXwGgU/hsO3LVZzCV9mjgqQT1
O6c5cqpFc0tXn6g+I1vUtfgFwF21KF3hlhNogHhDDpMWpx5385ldaxv25yTZYDKJtQpR683XnH6U
o+4re9xP3KiD0OZbNT5Jwc+Wxae1zGhXcdQlcdUbfUAqLLdXFmX3e7zmHyi9oE0gEVufyjjtuSD9
5YYmweZlY2S3afbygrY1W7QM1Pr8rUldjWPlHczWpH7PqjBUa3X3lEFM3h58EYx059HdttudBAWc
X4c7vaUgiFwSNe/dLgfppWnJt2TU61NS03eg3yCkWC/qJL3Sf60iBHzkyRsB08rXqpLD9RLuWr2X
4RQ9hj5guHb6cKYhjvArV1DFvy6TVcmzNnhb0uVo5ArhgOFtRpWaz3Y+Etrumr/dBO4AVCmjEt+Z
S6nsYM/Uo5krYPtFNZ/NKZey3bNA6FRjX3GgIwYrVERvhaj85csZ0rxQG1J2L98Zzeekj/nFdrdh
RBWF4SS5O7rU5Qpz5REgafNIrmRNDFaCi/aKg+WIsAWiUXOovli32BNgn1VVNKogrCypqoKVNB8a
Pi+nUKpcWKh7G9rtdQsGzbaSOa0mK++eNQZDJAr/qpItyaUSScZnjKOebqZVNtGXnwTyAQ3IQ3/+
IPOYHNA+RRRHIjd74XkUXjR1JxDsF6t9lMloxyXVzwMEfl7Zc/LsXcqjwLkT2m+570oD1In9Z55i
7M3unrw2iFXnwzdTQo3cqaQLt0MoGAqw7tJbueXUDmenNpi+1cSouDrze7nSAvxwJ447w+V8O575
BM9PAlXq5EvwA+OyMYwB68kXCTIxuKOWt2Tfndt65LtSgOZnnNopB6Y8OD135jZmBwx1WFC7TMkZ
TOAVIeORO7uNmY/SnMWhZgeLFTQ9R0ujRp6os9um7scD8b0wpebA97HBH9Gpjk4++H497qFzehEL
aoIppQO5vz/nV1BP0iPlDkQkkXaKuMWk2h1Gsc5PnSYVBjW90X6bRI7U8stdvDsq6NOZ3TCHsdD4
6biYa0e7pXZ7pxYCAwRfj0lWi6BpJzRtjNICyfKDpTB6d3fts2WddWo69bZ3zXmsLqPDOh+Rgw+C
h86k3HC6lHUwUVWk0KKibLBQkvWb+eMJjjCZaG6WEtDzEb4uPPoaU+NOrrn8ZnpJl4l5XhjV6WK8
6zO7mVclzlb71zjU3B9foF5amtlJ6b/BflOCB4NhaYFkl13BD0TjYM8YTILrL/fteOYOfnYwKEkk
Jnq1VjjFMOksIrShDJe6fR1wtPHHixN8XMZyyi5ovrOqclvn4esLF3GPyHmIb4j3YAtsus6uqkd3
0F6VNUrEAa1QzscT9wDBwFOrMfYYLlPyVI46NYU4FcCmMjkRgYQQ60E69/0drCZuRsMgqNZWyio6
hqDDukOYWCpKiRzpbQqwQI82asFg26dIqbFM/DaDwYdeml9c2OzhKZlQcseUqT9YfasCZY1bnWID
7JBcszGISU1OrgzlCC+0Sz3J5LrDwDVNo0tom7qMXwgeOtCx9FGTRZ4zbyZ2/l1KWaP48pnozxkb
+VE5h7I0fB0bkqmHwcuw2Tzq8qdlJun3tnKXFVWID3zDVykJEhkomtU2TR47X5sNc0fvoZEMDyhR
uE4hbJ394+Wulm37yvbwPdMUbcSS3bbxdlWKK797E464seQLJmTRU8ziFzaZ9yc2I13BZqskHvZM
aTyi5aeIzcWGD9Dmv/0RPIxiEBqtbgA4Qqbmh8GbcJmzJ8TH6oKXy/4GjKJImCoCcQm8gGfbl+bM
cXN15UO+fiMQWxLf4e1EJTEx5O6JLghpUNCehOGjz1Al5LymMaCLcTaMxbmIRhaOjvxkpfftbJUK
3j6uiZe9vcHsQ0FD6wH9XQM95+kjAkRA/b/zOK54KfTpYZfDpZ1wjXQvaGZ7tfVq1ZQCJckWX8Jk
IZuxi5T9CcmnnfgqUq8Y3bXCe38f4O9JsqHJ3cOMn3Zi4wJQWGFBFZI7/8RcFLw+hkx0bopjbYO7
hHIo4Cf4DO1NYRTIv9bUO0DR0UInn0R3WbrExEyDHEIOqFw37Pgv8hAU7+SOXXY0KNHVJVKIG50f
/Qm4nWyNZrQtrBr7+fgWJVk6XNxsIai2uZii1bJEz/lNztjN9hyTdQFkC6p6EtVF+n+cyJAoPtve
EvNAu9TdzK3kHh80FnjIgcV0qiFqJPYfYTUVAcEmI2t9RILPRKkuxjDCfCfknyzE06wcIfEIJyR6
0L29M4kMaO4crOL41Hp7GytbeAbrORSKEKWfJv6KtMvmBh4RiY3okzjKYm7u10jtiQEfC/eRek4K
BozzUYhRoadDlQt6AFOqyEKazF6hAMiLSh9j1a8ghZs1O9O4oTUsGjsOL/npU4xTnMuo129Cx9Cr
fnz2YgN2NYWKhbA/Z5Z+8rq7eGKINrD24uvDyS72EF9b7a7GCgg3Hg60AAH7XhMkDeJOO/xIYNTj
O+g0Q56WPyIJ9gMRdbsELdgZZ1AP4HZImnEnBunUq5DGnqwPRrVK6VE2focX8AFDay4BY87RcWcW
JRk8sh13pPYBlwUmFnQAVMjzNiZb1Yr8WuYTFe+2A1YG3jTMEliIK+ylQT/RLDehrRuFp8QRxJLa
b1mK031TS9vJleWOzS18bjgAm0qmd3cEeVE1VUt6YI9ZqgRItPXwE3YJNWbcYZ/p7BL7nwLlHRuy
MyKiGT6Dzj7YCnCgE0Zer2nZcmA8DrATD1QzwM0WAifrMwxpMy31IF138RMl7+Ia+iPxoe1QxhjV
Hj+4qLgpvBO3xa7foUA5f1L4QlRzrKZJIwJypkB5LokfnbrFzgZApClwt0fyw48rVmv4H3lPeTNA
+W7d70nP5XL6bO5jGqh/tIvI7zxLX7V6u8G55s6qRabLCi3EOnCMAmtACBbeQCydlUTU2L3LPIFo
atpng9OQ9l2uwzFkPzI7B/kwQOLHLjCmwiCtJAEfll7z21SfPk8+B0Hp68yRdGswtjwqufCz0mzn
JsUI6SUAJe+vWBKMd7P0XuPfsGBsFLlEwsWSJQDcVpXFUiS5Z/YVIFPXTCz4k8zlZXGc+y84qvwO
Lh13CwVBzxFB899+vtnC9aqpSwQdj0f04NeBhs2ukCsPVq7JiBpJqidWMyV4EufLiybyaxivXIpC
X1QzT6uCoKZSLx6bpvhaSL7aZkCjaO7QUZ9AXK8ad1Jx2LVcBjafV8g/Ne3N7Oie4gqcB5aiRqMs
Pzs3ZiVo+BLeCdauxJuDVsHE5xbcHkCN0EIQRUG/bmZreac7CLUSZBsTsDGlVPEIl9cAjktFiDHN
uF5FfPq+7SU93sWhhLEDVkLwWGbqAg6Yd5aEr0ITZRy/ao1QUQQNvmIGo/LVna9NL/22mwq3lj6o
SETrXkmXiq4Bg+QvfxWGMfqiSrCQbaS4btxGbwuwx+trsBpLU4vNinxcRu2QXF6oDmzNoZclk2Cy
7uHsp9mYdluZK+A3m8Cp21HbCalu57+NK8ccGpr0LnLHx/5M+/pMdB4qsLrkcWVve4s3WanPrZd9
+iii3jNPsl8uKXlMtxJ1czZvaxasBPd+UEeX5Fqp0ZxyefZPsDf/3LmN8cWw0TDuzw/oexOqLptJ
jOJAnZC6RRLY5YjNimc77u4Rqezc9D/9AgUoGlBMwULXQmLMiT3ys8s/Hj78HzXP+YM5ld1CnG0Q
4upm4kKozd7PLbFwt3FEBjcadeQBeHcRT/luwKRpz9LbJidaF1KQAlL9FPqjNFYP8OJqNlIWsk3Q
B4X9QjdtvKSX7X7UJC4/5Bu/+KUfPhMEB9rlohPKKeVKcnPcBuClj1lwJdyH3nszPlby+MpZuX/g
S1K6/rNMm3M12n+kB87N2Q9F7mWjOtOYXklqDY+BPWB3IFPcljfqg1Px1FDb+e6bl7NyYRve4LtU
o0ggKRDA2xc+KQiXMv3SnoHTWIGwFhDTCDpO7jqxSB8te6fPhZCS+g+O2r/YGmNTZgvLRYXwWF+h
VJpX3X9FpWDmmWDmQ2FSKYSL11ceudkzes8kGlcaU+MkWpGSmR4iExvCnsfcQL8KnvytNWtKnKAp
V6i3KNwW+006QScqXcS661L2+8/T0bWUmUzsws4Gk6Zl56rOMV+xcVcFmRu5a/8FyP3uu7xZU4gL
vpIQ2R8ZVhKM/9rfmf5y2z70BhFX1fDxu8id96eepONp2vc/SpEcUbeIPSVIPZRF8Y+VKTFUAqiS
6DunU17OaHbY+dp3YoBCoi00NwI9aM5wM1lA6egHglgkKflTw18Y0/jd5xN3yIvBIa1D5Uj1P22w
+m6NqybQpQMRXdHmH+YBlqcz6jAwQs5Hmt9rdLsluLP6FW7pxRzXAe92rFsmoHRFGpSR2ELb0oYe
w32NzY6CabpPFuxfT9R6LXCbyvyBUVDDAq2QhzgNu1voQWEQX99XLfruUQNBTH44fx9Oa/WIA+4G
BdHNCxjRtzYWlTP+yepN2jlFWIbxjEiuhqeAfO2AgwtpBSWuMhcG0HIRDtNDvLymk5aNkbOuwW1p
8O7VbkDfWK2W/oXGQt+0IC+hv/2H2xT/Jvvr8JYHY1ixBE/g/bEGWZIfSarvbdrGDJFr31iM5E8J
0M8XJ0gUmyhAs7+UaiZPKGmayinihNFFJJXpZpIJUyZogrhpAy5TbeT140OneJ1HB8uP7tmQ23xf
+i4k9U8DRzYYPNYTguqmzbG/xIeLg1WMGS3ykeYwIrtm59EyJEiiJpjT4K0NdxT55ArnTDKMwRaC
82IdhYZo6adbFsq62sI5gZhY+GPebGhXQsuWtdpYv+vYUzwaFCD3bd4LftjUXNKxzI5g58Sa9s0N
LWjc4KbVWQgbK2gf2fipzIw6OXQIjutzsqLcgbq8v/CANKBtiN2+M7qv4ZRa1SszHA/rt/0h8S5Q
A4B4gQhujSkjlkQNLY2EAeGkXSGaOIb2Pc24ljVEEJJg0ynbx17h051jvVY1t+qlgzszCw6qY9K2
8BmEgVNln+eTZqb6ZbNXMMZifxIAAEVuEYoG1hj8ZwY29e07MXF4/SOn1fFBAJXK+la50Ahnx8HD
rDW7LNBN5WpDEd37l/Dl2eUQfFQcJgXhO2Kn/sUtZiEIyfhrCDL9EPMtwEhsFTT3freSyslTqNAS
82FK4LrEplhla1srdT4p+w0w6YWDo2y6gQd69S/MUrEK49n6cq9T32H2y/TKPjQopVient0y95Ar
vBLYlC5CYfezbi2Pbk4q1qczxLzHISvuUXN/wEwX6pnmA5iweCsmM/CH/QwdWgBan87l7B9V9yD7
MHC5WsvA5NmmfBC6JNgPu6UF+luKjtbVwNl6PAPLeqV5rsRf0BrXcJmUopcNBkd05Wf38MLc5J2e
HOiwnUU/+qaHu3JSqkmA80rG0BeHlwdDKsEXznCl7+kSRvqOpB/3BAHyNVhd6XLsVpBk6IyBupHf
CVmIpFyniNoWD0TG/kzRQ2po2ZtHkggWM0Oj8085KvK1+RTrqeLpK1MZf595zGzwtnjd6HGp9YY7
nEFFgT4dMhT/o9xDsw2miaBjWDTfMrVBbus4mag5UP59EfZbqlorjVLIEp82LEkTaljQIw+a6yhY
4gdniIiq84/++md1J/FXWXMsn05nVv14WLEa/K8G0SWwfdj0LH85cismZhBMp0l2tZfV3ptgXoF9
wl97dIvDQqdOZrDdOoaxrYPvrqf4l8dfpsbXTPy0pSLpQJFMDt+jrLsBj21e38kWje1hwUeA+wNj
NW66+RHAUP/FzA6qydVi7gBxcg0AFPRrKOJu4n1sAwmo0EyO+GKFyrn6K7gg6Q4qeMaCM6q37j0g
R2YSi2rwuQS4PCM8cG+mF/d8H+csMn55/67ffYiVd1QcqBut06ZRFUMV382ATY43F3v0wciGSlYo
C9wONYZZGzB+frJHXfN45reTkXGmGsfAjI4/TfsW4Mb/M7ArskUFLm1RY1IttzS5VsUCmdPAdCdY
YKGC+F1tpWUVSedPnTFxYCQxMmXwA/v/T/GHpFf3UjcK2fWPC3Eb+9mVkiR2KJ67Y0CfSb+Yya0o
nnCEtjzTB77pdA00DW4voN5usms9vQZFk/jNHIZN7Uv5A/SHUqA7PsrLQnsQUCfxOYuJ7IEYDWxa
APKMQguQCioALeRJgRG1cXDWhDYne6E3k3L1BBglX7bBEXWizpX9VokehJag+D5O/TdudZFGlEgA
r09/s/547JlP1E73f3FRcC4G1Pbbqlt2bWzKbC97ZrjEh0F54D9DYQhZK1Xer2yRadDTOF9oIcDl
X6EBLqo9B2dItHPF74q4FJngFsxLy8Pa/JmC6Ejq4/axGrDiATYnlsTA/MG48IurPsg+m3hjHLdy
bv/6pPEzZ3OANFzYld8WZKlPSb6ne3QaWCLLnzjUFk3216FyzV84FG+EGOMAaxLL6m+B7hcO1f0D
MLvwQWSWIjGFvYMxoU6tWcdW87oVstETKawFSnU2ga3I+bZeIl9xxe9b6za0qSvVkqvVsGF6gR1w
FaYGVpPkJxPXeUPr7DpY8YLX+HnABgMxM5kEXrv/GrKFm2KOPypz/us1WwIqMOOAmyf6eIM4C/u4
jPG6Qzhqnpau1zlKJXC2AR4M0UVR+mxQnZXko0kvUjH5p3nEbz45etVdMpxzn3nNkszsrxXZ/XIh
Vh+xrSd3ym9g/b1JR9+UWLRrJCrjuLBtSCG5sZAqcarVGvmw6vyqkwx44IrJXkyPBwnEVfEqS/Rd
j2AL8uxxpbNhNLzgMfWJPkDxc5qPQIGzsLLo1GPmPlbUbMlv84gtVciIWZ+us92dwWpq2ARws0sy
YtYMNjM8I/v2sfOyDTjnrLVUddTOoD4yE7u7eeo8g4FW8jyS8V6qGmZU6mwk6lp7FWUbfl25VWrT
FVG6Q4xU5TKyvwMsm0mk1lwytYhpN2yogdyyrCylYARwqwDkRF9faxRyhty4M2p1SFzUNZyRMTle
Iqgm+nyJOvM5mQ8yHhCJaUE89ZZbmmyV+ySFRgb4ezXsAoPO1MGIaG2mbfYRae/7eXl8f+nJupnZ
zTMw/jXJg5faiSV0q2ppoDO13y4nEFFIivUApVr9dJO+OvlA4ppOpbwPZpIr55H6w/obqvHUcY01
72mO8P5cvEv0111DtdfIp7FqyI4ozaX5g9UkajOFo/q3sqa8tGpnlULcuVc8dvW43cgqwyLipwbQ
NOFh4aesUziTnTf7Nl7mjcGG7SD8wEGltOQJYp92Nqok5fBekr6eYyRyf/XM0w3f/ZA+/mzzm3D9
tDwZhz8fIL0M4KQIdDGH5RWtghYi81xXZCwb0+gqRm7blz/qcekQq0yk7lsuyl5Exeq95j7CevPr
jIbFayFYv7/yUZF8R5qnzQjQPygLhfuKmcjJaIpG/jU4ovkdVrBiwzXjE/fAbuE18JYAegn5Ly4Y
tkJE/d0VGvDF81KPwXms3qftEcSJQHFg/q/miP3/d1/6DfC/hOyP6MbbWvc19foJBuzQyR784fZi
0uLy5iCKCmuZ4se8DbSlKpfS6MgLaWHt3qdsa/ZRXvSbE15qApjqNUKpS6+vdNS7w37YfBNxyYEZ
jDtmwwqbXdas2sKJnQuqumRl2uT43Cb9cV1qa488YVQDX/frRLIJ4Dpx56a0nXCNVXCt2LyWvX+E
axNqoq6JvBke3SLExRH45wujpX0WwlbC0SlBGOl3Mz7UgF/RJVpmVudnSsT18nNv/T/i6Z2pMn9p
yzyi2vFxU+urDIbCCBEVRqk8aLAbuwE+x+g180/pQ8eux4r2yTwqWtRfhQ4geMV/yEMWoPepRpd5
mcwXwS443oNhO/Bd/KtjNZb25Tfemc35kj0+I4ry2Y94EJ0ojgEVxqnds/YIYV7gMHDjN2Mxf4eH
WRt5/4X8op0v1E6Ea1+9lW1IBWrLc1sGwIoaJmXaLZ1kUxRY/6ifXdwnJNyUIMbZy84SJuT313we
CRouqWrpEe1ShRbkDKNyC8LbLipd2IJqEgxcTpWZnPVgqEu/bOSCt++S+rf2ezCo3wC/Kk1ZfnwT
jtBqLz6WxC52DM9z6Bwr5XAq428fSkx31TgWkZenapOd0Yxtj1RyzQwlGmDGpQtf5HjavnZR5vAk
noiXh4fN0Whm4j7WeDe8gb3vQma8wPWAj4QfVPUGKm71DG6oNPXpkHgAPue6TeL4fDL7UoCIxR++
n73llfGwO7hhYGVpd5NkUH+t9PZ/qguzezn0zgT8Eky+FtoVdlhqD/R6bDPIBejwpuw2hQO54sRt
y1JkMKRNoV81gloqRc8sf5WhXrpDQn+hrnoDwELluOuzEhrc9p0gxpYBanQ8UxLQnNuYtOSqOlfj
04MsnMi5EuJ+s26Z5ricn76kCE5fmnZgosxTAhdU+IkeB6tkQAupFP9XHtF1bgW5cA3ksDtfvN6H
R8a67e84EHZZ2KEhwTiV9mrgWjobOIyuEKiYSCMv+fwrrdzJxh88SkMqqr7nHl84koZoBvtWXgNF
iLF03F9Pby1tRT2ye71rjtZ4RipLnB9qFYI9u0yoa7rrF/onZ5bf74UFZApnsBdXQEvL9PjQnoDr
OR+QuRYYH7h8ZOQwZq/3a52VAdcs7FEHOG4NIsdhH0JFKyF+fVhgmNyTa6Z2Y2KVok0zAtE0o/Q4
crFcjBmmQTkj5KZjiSOBxBViBzDYFm+Ys8j1qKlCgc1kI956bSRTKFOmccI8bx6YWQoSItrBeMH+
U1P68Ireva6BWCmlcOavsuOQS9lYYWG7U/wTJppWXqMJHZzQIH+KvXxGxZjRa5VkXDO+RI5+u+fo
46jBI4GW/1VqmpQy5C0pXvW6Dy/EpY6spL+pAImEa0qW1tq9+lkqtx86lUwTrEmzu0RaTrLVQzfm
gLOcMxEsliq8e85uE4eGLDUdxLCl+f2NFYmCpU7PjXDdP379jJ4oXmw+gfVp1CpTYFpVAc6euZui
Vzh1oGGF/XH0yruwSLTEfp5ROLzajHp6SJHRnW9xCQae09AlIxqXdO2JpTeoZbZsK24bmqmcV7JZ
Pirn2XWgz3v4VnPqgpEIaB9wSF/6PoyArjR+eEtHMlza3H9tskIn5Zsdw5kyh8VbOfZyJou9vW3g
bTrNhBPWAKSibYG2kgD/NQap6Xx+c6AHkg6iOYIftT+1fDnrR5DmVUfk2e7ubT+CawPkG6bpwJb3
CE/cSb8GDt83FGdKuGC3otnztLYESkdAdEX6lzSWnUQAVhfxljxeIO1f+iONk5PCq1Wi4DHIy4ws
xXdjMf0RszQ+UC8Jeprpo/AcUpLWDx92tPuI/VNgOvkSGxQY7iOff9Tv98boyghLbo1qlM79IuQS
l26cnKQLW1k4AR7RiRPbfz2m+rruSqlYr0EUr85LTYa5P5/c7Iy9aQtEAkTm06eRxza8E63z/sRN
5JheXLp41H1gHFexqj1H3nZZ92YULGtPpBOA0u1ATiL4bwg770SY1T4InemwWCk2lJqHHZAmb54v
0fJMktRqn0s/QozQ0csak2/qAdWNFXdXZHGIOXPevkm1O3DjQZxYmOR3ORfE7Fq9gTlpoXIIaH82
0q8/iDcvwk72qbAAEZ0BgXsBIzfHV6MBXyerIEK0NZFyHb6b7cU+0qpdpDEx1JrYsAJz7Y3Wr2ZQ
1PXxrqtWwrMAX+lVQ1bDu4JWXIbo3VJaKGO1sR+0ijZRnsqDx4XtCgs1gVIuRohpGsPdJ3MdAYdR
eRIKuTZH4VuDyoKDbWxJw6RFQxfzx0EsckjiJaVmwsWcC6NbMQJ3fgeuNt1hIVql5xSgqK7cuepl
Eks/jvE5YRlq5HUWAk/SUqGE3t0nsqtcN6suBlB0td7IgX8Futxua9QknoB5EyqA5Jy6kN8+WZHv
DAhZg+AizBXUSSNWrP2MhCkt5/IVcqtr4Uwn6hQzyAieNJf7zvdEcN52fpGuL6mzvVcRyV41K9hv
C8AbGthY3wjCxHPdq7eTpnDbUj0TtOFAbNTHqcBebi7R33bQeX/3LFduWLgioACCq35zBHAUG3Qp
PyxkVw/oNszigb+5b2zMYnXpYi1gUo11dv2XOWmYAG27VLxO3Zm0QXzXJocdXEh8fqUEQ2eWGrfh
0biOake4HmWE/j1asNnRP0s2xhZ/IFmP2gI+1QCE388D6VJd/+b6APYh1GKOTgAhp6TyljMkLmh3
qtb9Mm3tjLi8RYFuTiyCZro4HXntBbeYSsWARSv1/ujnE2pfOQngEktgvZo2rQi862gIhqZFb1j4
BMra7sr1+XYZDLn8KJphlrEdKBrVEw9O5r8vi6XOLsFI3VhOv+bTtJqK7koNKC4OcLxdWJD1rSjE
755Es+KgTJcRPArf7c1FP6Koydx5MwpSpzeIvSoJlGFG7qOK2l7ZFFgu4jxIRebtkqRu7iuu3hFL
yvK/QYaftwRCyF4VEnXD5RPQCRatyAvadJajtufUPlviidKbWr731TIHfq9gCsnodYBWBj16Buz2
ituSJ2Zf5KoC+VGw7VJWNWEzeoaEN2PccU/+wFXrUdQW9J2hrCUdF7B53tA9og96TWzTE2Y0n2VK
WmZ4yQ2P4g8I2MAtoWFsG8MksjlqNboNK5+zaEHONFVrlIfpYKsycW1CuAwh9+jtYy2iz4mGt0Qz
C7odiXxthDCjxCR132f5N48lXj1Hvg9YAUpWizLP1j/XHFw8kIzSmP5qwE5mEkWlxv1OmM9LEVpj
3o8QCPybmpEn6P7KwQOB9A/y6uprZhp3BFuxVjswZ5IF/VB18nbiX20KOCyzOK/7ArFKnJhdGy0Y
/3U1SLFHyisPNj0v5EcdC6xv7OtJ9KpsAu6+y7K94zYChx0MKoJyIcMwLmuh6xObfdTzPA2vce1z
C3qZrC5NjbbhRoGkFO1+U4N5n7cvwL302b2x/3H2gcxP0Hc91+V4FBrxmKlPAcHecZCQTA2p1E8u
GN/fgtW8A0KQc455n/WrNDDcwbx2nsdJKJZ3ros=
`protect end_protected
