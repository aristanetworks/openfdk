--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
JPn8weYlL/yeVEuHEx9zlBLEkn/hkRz0tmp+GhaVKCcxtlGG6taKzOJg5pwlfkl9Q91s8PgNho+R
LYjCmm5Ud0vOWv9wivX77+Br/EtUHqMbKbJSqSHjWG/B8+wil2nN2DcmL2gU8I/O1tCtiBrdNL2U
5Qa0RKS7EbI8S99SNUZ1gylsQwtCrhYuu5WBmhaeMqFmQCO22MWWXs6hg8kcoV3ELq1VW+p0EqFA
G4dFvDVKlvd8QEU2QwV7if7lnBxNHdR8IcJa4/68J9clsKFzSzzcjaj4BJx1/hT7+nSo1xLqiNEg
05iUZigEuMH16XUDJRlQ5WSI3wvvhTWQlD4u2w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="4sh4riDpb2nDfBSGfXvWLKzu1NZc7ADNk88nYZX0V0k="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
NsRmVk087B2drRPzEP2XBBfanGkjUCQAG10P5r3YA4nILYB/PGgZm7vo/lEM5o4rvBWAIXlOGPwZ
BQZ/lkhxJBJuqjkQe24lzNKq384GQ38pbubRu5eNum2PjKaNJmzz0FJXtkD5V+jrwK+652qvArs7
dfpWPP4zrvJEPknfBEMO1a62CB2rNqqJEeaqNOg7Fb3suvSvjM7lN251LIgWv60oi8tBqiZ0Kfg0
dLv/NvzD3rIIF2WP8LfJmp+jiUPyatKxjtaxk4hgahIqY9pm6sXiMxFI+0MxRmTCsZGEZAL0bpX5
C1hPZidyjV514HmiVUn61xidGyNGGUeb+i5pog==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="7VBlWacuL8ZbXMdtz3GlMsLa/mGp6bYxruni9w+78Sg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12336)
`protect data_block
PxwRSVLeOpGmxuYhpoKPo+50ipM7oF4pIxMyiZcRQhlCtR73QPyNgsIi5K+CvhRvLRzOFxymr4cb
GpQpm8ycve/nU01azBWfvB2P45sogNRmijq4qQjWq94MgwUJuQvcNl9Bn0YOdt4MB6gfMWbKVXPi
mWHp47hGhGafoLrtvh9CfUVSbV5D+CyPNK/pwSLNHoO6ZlteTcl0u3YaH+BSJciL81AgiF13jy6Z
lAwiDF6vAx9YF0rWDjiTwQypYHGOQLrL45WFf6Nd2oJ44qbUwBqAR7ve4W128UOCAIe6x/UToN7Z
XnhfzZvwyoCCszXZAxi/6a+xgrIbE600A7xg8+Trsi/hW2Rlk+zdCYOXavLE5wPpngM0YrGM0pHY
MgAHBrRPrTDeqdBWWMJyJRfG2PFH95Y4Ue3vuOmifLSCAQALGTa11yw9RrZ4aHP1ml9A9agYT375
Xsr3B/uvFJPbSPf3RcABRLZhOnIX2pDHy5TqzdtUSvFJt5WhiYewiF2YYCxXCOysxZFB9CTIXzuy
mJmXpHoFyBJTLgPI74cDyrbu4QXHOxK9HCgaDrz+Jk3r9DFP5TIZdPmWH83AQEtHe3mSn+1W6LhT
z5Pd+5ANdFtXwi6fenyigircRJUy10utDrvrawGLq7voJXommJLHjumN+ph7gZjPaJHm43rnvaOk
JEeenRk7Ps4qNltSJSjdoQQHQcReUDmrB+iZedfNigL1LBAr+eVZjM6xhfj9qKFWzaQqez/M1iS9
dNykSVCYQmPNz0FmpA7W47Nchka8aEPw1T8kBoUtZZSrvPRMnz4VINYxJThygvT3a16H5z1kn1W3
w9BLm5jYuTmPsZOYkQU0Z8cwTxz9iP0XlcGpbuiGyNqtTgOh36rMNjQXdQlk3DeZAsJVg0WupJV8
Z7g6zMkNPzCO81K3/xoa8DdO8g9xgIK/5fudApoN6RWJ4gYORxnTGoSrzqDLcG1XDRXizlCdbrSL
h8LMjPRFPTB8UQzUpsQQaGxdRECxQM/JoQQfGb9VJkMRTLVr4O6yBiMhwL5N4RPNavX4/8qHFAlV
VA54se87yqj0eBFOMtWiXxnhls0Z8c/hnGjPrh5jYJfVUJnYdyHWq6wDkCzzRMJ5710i/LVYU2YG
deGfRNdVJJUouR7x5rVI5WlcThUr5JMFDY8nplsK+oHJkVTE/NZmsP/XQeZ8xX14DvvWprEYs3H0
eQHLVrxiCMSheyoLuEMkiMYxcL79OS4+YvFiY1Gx6nhWTi5Fuyv9BTlc/f4795UV7MWjtVyB9ovU
ee/ac0ksTMDF0+N4Y+EKNeqEv0yq00vL3kBt6BE/ohdUrOWtiuqZfOJZp6oIJBswz6eZ8DV/25Nb
FyVwMAxUaN8ilpGrdhkYt/ZV28fwDMalpn1D1M3hlJ/NT9yZoeduVSsvVOkpPH5OZMNKgDXrgfjK
2VZH6OePrEwLK714pQeBLGBnvNy0uTLDdOI2hWeqK2H+kdRFPPi69c2d4n4B1tWYRIIm7L21CJi5
gDCNYtpJMmtLre8M3Vz8GMfLjC8g6t0IPfja1TjiotSllmdI8O8oDe5K6e+lwLT3Zyl6s10dyHZg
JFOk6AMqhAhbpmvVaNJy4YpY3ByLNoUVAImNEYUru/oK0H+lXTLz+OBeoX/43n4JfO9lqJw+wLKB
vSWIjND8X7PGOpST11xs01LBqqm00QDKAoRfau0ZmyjxSgqoTn5LNFx3ebTyFEWd0oFt+TrVXUw+
JhYm3Z2iGZKtjZHymdeLz5aBA1JXQNZTZmQhs3OxTpJOkXBmaqa8PtkVOHXPLtonqXy/rT7w2roa
fRZibGhPuFTCgMDqs+s8wFK7WFBqMOOT10O1eqBTQVmIYqM2y975TyGYhuQ4S2gFSe7WWe6hCygQ
ljKZdn5bnufTaDgjS+YYQ9mKMA3cV2C0hLXMvJWZ+5ANOFgcMH2iokywi/WQQxRFs+YdS6HGFNsn
Q/DRrXmU+GbDPppVzwYH7NLm945xoba1IN4MEhI7mnMLm8bnmu17OV65VAMBmEqOxTtZ47VXhASr
aRm17SLkQEGb8DIzjekpFUIQyHvKo3dn9CpAsstxF7BRZfMWRdf9hr+qGifG0wMBRBsbaZKhKheR
g/qMMtjU+10/HEB5jLW0LTEr28+TL9OJNTCKmfdXGdvnEm4cZJE4dYH2zdpIDO6VyBPKm+A56pjw
605dzMLMEaeTA232Yup84LUfI99rgv1FR4RF8blXV11wE+p6Ak0YMG5Q+NN8/gu6YcFwV+TVv1OE
KaGHybVJwz7wa8OZ58El3v/K9KX/wzeB0/v7PJ5CEIePX/+qnDF+Gu32GUH6imKl3oCjuZ6w+gBR
pbMoiXWZKUI3ggUbuJEI7wW5ZqFAfuwxRcrXcQP4EeKH3+FF7C3M2e96Xsc5AJP+trV8UVGf8YGG
zdmba/+xPyMUF9ZrTw6aV8jbkH9lpnEzkvslQJJN317SbWHbdcY3bMW4i/PmtHxsKuk1BL9J/+v+
p5kL4wMctV5qluvYBrOJCGICcy4S8Zy+y09eGQLzUkzaxFKfo1zwy2+g3I6GhA/3kj4my2zjW86c
Zhqkx9ger0FIdQXTZbOVxnIOKbmZ2EGb2PIi1UtCps0cn6ZZmb5B4nyAuOiblowl+BLLzD2Arhl+
2/GVemK3FTy6fLTOb9driWVqMdPxJ8a8dQF1tLpzaVclEP4TR2nFCM+PCyF0bA7jCIe5SgHXYEmi
2Y1SeIAmmHLZyDDYIfRbjddYm/c4vcG5V8BO43du/D+Qf6QFJ6jgnx67FtIjhmntUmY7J9tNQ77v
BCb9OObZWwQdYXDizGDV135MXED8f9jEEIUnS4YP3HCQJ6NSqI07zgHF0y4w48OmfO7lmQA/aJFs
tpmscx1tWsXeqBKCpLVsUSQBUTse8LEGLkKXQ9vwudeyvLvc+80vWDWmUvoSqe/BIFw0XM1ISdWb
u4Mur5UnGUAZqOOFTSekOf/MowBcIyBvSNiC0qrZ0LiEK3lv2W8wRe6kwaVc90MrgY9MztpHxGFD
0HteFVyGX7+MMYfxS4K/YNohKZDu9nr14IrXiFQpVB+9EJhFaIrsEA4Y45mIZEFl81IdHW9nJ2SY
7ZU7r8hZJqR7igujCNQNMdIFwcjLbj6JVwPWZUG/24Q80op1wHMJDohh95IfjJDvScBApqKsh1eN
C2kWaeZILTm9W/U/vrDy0jPjaWpgIH6yf94aniUmNTg1Zq0MB/htbF0+pHOm2XroSlhjkTm7LTPb
o/qrz7o6Xr/C2FXbingMuIq/bwTARGeqM0ttEbHOUc3U7tK2hwshp5mrlr6tQOXqYZalCQG3iJK8
s2h31GHy2LZO2CES+BazWUs9Omo+BcW5csi2C+cwaUfw84CSGwaufxLieF7QNsyMRqkEN3FgC6Zm
0MDQOB8kFA6SBdZ15mtuCh/jY1dh0YYU6C68n+ssn6rUnoahV54FbJ0o4isEDpwtl7xV1McfuzOp
qSFxCIg1PbBRJFqbFRSB3jmcJcXvvo8vRzvcv9NKOq1Gd30OC259qT/z0clP1Us8HyHVywcI84MK
ggm1KCucKZDFU2ztvAxh72AYqgYDPJFcDYUeWgpK5mMtnKT2aTxqDesDVkuwaIycUrz4EPVoHKjo
yvsT8WtT6psU09jfOQ/G+eBiHlL/ABkeHDWIe1SNjgXG3WV4/tluNOTNNW9me+F/AAF+1PyGeiDO
l2IMS39T6Cn5WSEfCUJyP57ZcGIbA1dWMoPxR6K51hoSfbvTuI3NQIlktbVhpsHRIHDc/i0VMF0E
IYqFI7wqvQB0N6Vz5HUJHyEpipVUuyNQAPZMSh7yuXY0Gx7AbAkWAQYIAx5N6iRPgmhqFFijBXEj
uHZjQRcE2G0T0lyaIgr69/XmPHy8hYPrvgFdy4QJUVCu33wkHaNkUWgDawDM9ZVAO8lQWFuo7fdT
94ycJ0F4NRjqfKLa5QBAGBWauM1XB+lqH+XxAau21PkwcWXWGmzPIAvQIJlX7McJ3Zf6JH8issSN
wCMagGm5fgkhY1MsPIJW9DOpN4r5c13JRqtZHVvyOmQ+Z9LDnesBiJ434q0qz5RytCNzJZlR4Rxn
rxE0xli97a6guwqqKwLpevjRRRwrquxJHaPyfEeBhtnWQ/ya/QPn0wYRs8/i6MjC84hBuk/btz9B
H3Tetjs6Ov9YyeZSPViYhIImjkJEMtN+EZVAxdVVSeimUQrPm2N0QLX78A4zkCOLkVdjyF+/y+U5
H/scC+JJ9qS9WkZv0i03IEtSLn+LYFRUMJQ6XsgtvUMjYmfmpKsNM4f7LA8gs+26Er6DF5TV7t0V
U2DXjmXUYl3FPBjntLWKH+4GlE6959WNYKulgVKA6Wv8VgWZVAZcFv9pOhVg1Qwz5gNwpARRyuze
CbffKaP+At/L9MzomwdtMZdpNTU77yBhEJixVoqm0uIr4qnZmP3LpWUyZ/Bex5wrJWkhrqzedFxM
zNU5jb+tzqx9yZHA9EvlXsZgqVK8k+0KF4fAlYBZxrH6kQBBkODBYUmOymbz7OX/6f2xTj6YgpNR
Wl7W8KCA7SGmkh+QLuMWyg2xp693ANB2TR+zhtes95DnWfl5Jd+kGiPDEvUW2k399Ym3UTSOuxJ2
2kNGxv5hjlh0Vh6/y3v4f9L36BGA0Pf+sROHDxg9GfPxprZysED5e5ij7Zz5OpBcBfqA7nqwicNP
Fx+rNbCi0+3hsoIruMeLHIJx7Kh4gyNpmLWi1eoVgyzUdCw7XFRXw4D2NgqKC9YjSEgF6vMShKz2
2b1eBAVNnT4+nFob6FPCuKL7XyULZfHLeAzH82UKnhh+qeH8K4HTcO1iNz7PghWSzMcs1ysoVnxw
HXYjnlSNf/SvQjIOpyRWJLvDC8URlsialFbFH+4O31sI7pqerVntfcvjajnPiQneCpegQvcOef9e
hl8Wlqf57nAY8UWrkEXxXzNSa38AX4B+Sci9ovKrsK+M8ozv02I0Ztp3jIn6c4bcmC2QLT4dyzyU
7tbgSnlheEKnPXYhoRS6+CGhdDmEnhxjE4wD6fClWaLww94QrZxT5Yq9pllf+L3lzIhCUSC21y0W
URB0kcXkNWFUS3cC5YRhiAcWPNFDpJmLKs4muhYEJbZ0/995+jmZtCjZhs8hl7IwpRrz1T9H+FRr
8h+oDCY8u50px8Weo22kXJJfGkuCNI8sRGAc0P2Smh81A1B/Kgi2khvYNMzAw9alaZipaZFF3l3B
IwaoUJ4mXy1VTGygNyq+VcgGpwwj9BaHPiMWPigyryjsToHQ+w/v+U0E0QSCRkDNSLYLckqrdtH7
Fgnr8UrravGBc14Jbbv17p39ArGOaGnl98go22a7W61ljM2XlcEk0Vawgt0ApYzE5Z1l5QEIBjLN
VTs5VkXwHk7UDXRvZ51PpsHUbf+VX/fisIdM+s40UU14b7s8T2+9TlgpmRp8dvTS8aD6z4BIyt/0
lcKA+w75o7Mldu1u1pUbive+2Sf5l6WX+DmRcUF+r8FZurpbqJSaMr47fItpb3c7c9V9qY2wLkon
sNo/yD62IQ+7QA2TH24bkwYkcdoqArmYFaYjyATcYw+L4Ope/H1E4n8/1Ez8jqRjs77rTHyuAn9+
1Nhn/r4lr4BDkDMWPAyKH5Brtrkpm+j00JXwsMP4esTKZRChalN8vJCRf2RTuGAsLwVr36BBiDt0
LNdg0V9FFqJrahkzfEzRKDeR3U3QxuEgOQ8LGGjpgDD6bqk5FYvV5dbUM5wSTLc10Zut3vHvKvkR
IIByWPeNYZs8cfdM+eFZ8nMe9Gx5bCtpJfiVTgWmwOnI0ky6Tg9RvjO2OTbhm1frhnWRXY8X6jvU
2PC68feBKzpJy8Ozad0iQQqVEp9YwSuCwCl4HTO0XrRGMyHmKDTkkda++YR2B3BiFBkO1P9So3b1
bTbluPk1p7kpe2Xp7NlnNfP9fUystrPdQOnJSWyc2399ac7UbUlcF5kJClgW+uy86Y9fr61AfFwE
mDRWUBGgwWZ7gRok0ycvScQLUqkp5JYyrbraZNT2T8mZhBJTDM1n1ujyVxcfQc8pl+w2gD+dLahx
YHW8W7Hrz2PrthEhCUmtnOf0u8O5BynBQ6k9GBTbVvSb2kVDXOEmmDJiJfKlGjxq9FSvcpCwNEzB
TY9lOB0quHeGxFEHa3lsYDbmZmLHLX/1YF3r4ZICBBOgE+DD9fkSqLW9r4pOYdeYm48pNiwm/bxM
SmPD8oFnPZxYeAxwM/YnCn0tkBsATDWLfc3ypUqtZRlJ5675BQhkonG0CjRllM9yVmJ4t6qzIbp+
j81ON56Wo5BBKZR2Ke+G8oPOqFTdBnPgeUiDz46UMcvXZVj+NTyCXj0F8wEBHrfPRADPmk29FG8Y
41Ze48d8TwBYHB5DpwSFnFffog4IABQZNqBvqucag6ZMmiJPe0mup0XOnbTwG1s7COYxMpPJcZat
G2/jOmTqn4Q14jAOQn++ybGI1lP+uwUEsdKWnutZekR1xvw3h4+knWDvmLEWZ3IkUnWD7V5XJSFV
tqJ1Z0wnGp2UlAA7VMb4ncgE2N2RcgveGqasQx7ku0Lio78keLP9k6X5/onjUxLhm/e8QdnLjGlS
ApilvNul9uc/OlUBmMbEmf+cwW6oE4U/l2ImL2ej6hnqRWesRip2hnPqo+9IaMFBF212CCR0jATX
pUH8btc52cSlAwXEE3PpaFRNiUUYh2Ek0zGf6H08wZ8ZI77vmv2DKenln1IrpdRGzGOV5uvRLqOQ
XCfzsmtIoiSxlJAiFgjnAQQyu5rj9qoa+nOd0RJ+H6L6j/36ChgegV+haWWn86yynF8/JfVbTySo
Gk+EFs+uVH1NYjSrabY8Gv+SMmegHQ75ZxhxhOZjQKaNEy6/YucrlWMjqnjcxV43ZhRTZu27+476
mO+q5+mBVyG87Fpsv9GpwQPH1nKA+eu4+QRnl+5fJni7Rk8Z12IcwHy/6HJ7tWoMxKRfHGU7BHhB
mMl6yxC8L7h0rWm71h1jPXdJO5wVvC3q+JnvbPhl1T8Qnitz1w+/P/tlyvgbyHtVSoNYXpKPrby0
1pP8nev9hiL7XeTfhN3/s89n4r+l/kNTumT1Jc5uVX95AteJhMISGsrprAH5u+1fupQGUd5rxYTy
fITje9BVlWup3cFqX+ACubgYSzcSYHNIy57fw6/lt+ldXymq6F3CqBeGCYpZ11pRXLUeKaga03YL
Z0duMyj4d3N6EkF+QaqS9hjNaSCnQ2m4duQArRumIDCG6wmA1t5F9KKJJ2pxBED6iAZZcsf3tU2z
Rui4OXuRTT6AJym8D+Y/eUXw3jQ9fK7XgZNM6JWOhlyfBkz0oioe1o/7pWbZ3gck5oR66JNPKWgZ
G2Qx/I/KvjmvphAULdawWN5f3SH/bti9vWWJ3gXXsg7H17GxJLtrVcBKqhpMShGgyZx/52KR/0QK
UQhjpRSvFlCNsYivEhI0LJsJ0A6NCK6td04P06p8f7EGmW9pNf4Jied5j6YSwUBoTSxrB5ozSyJR
w+/cWGsV2cEwG3+2Yj8PlkgY7pkGCXJ5/CPyd+icR645Tj550YfkVVi8O0+61snyxbghVJpaSmXN
CKZvy2KN+16MtrdNiUar45f2cnVuZq+x02nCXWFxWlVxvKUQFVW24YpfQz7hJgskbS4jfZn0sHG9
/nhtf1ivsxHQWypUaiQ2oB9wrpeqPtx2VLVTtLofZDr6/6jaXGbYZxf+5Vmp6nqEHh9EGmSIQvnZ
ua4o0O3yvdMKYbctaep8UnPo73dnutGovzROHvUhGGIX7tD4prsWZNlGMgc5g+seI3IQ2WXrj4yw
fBTa3/gyafBqq09HZwGWihWCz9KX6vEuf8uKe/wIINjIpMjZd4hkx9+b7KQPLaAUFS2lg1m20ena
vHD7wGvra9GWbFlIMnJZlNsLrfnQnVdAIcBmjKzGzDFkUdZfYV7mkoB2KcXDZl/UsAaeyO5VUFBd
eidq183AQS0mGsvxjKXBwqbROktmXjcA3KrdeFHlAkEHrNa4i0UN1CofWkcHGqzMJzsKbVC35JK3
kGvtiEI80dDOsf+a0fDiOxdwicNH/PY3c5ANuLal6UtXdBVli4LukxvM45Ov0qlEofnlM3JFLfMv
yG32cnreh8nqK+XO+yJ6KQZrT7e1v2DvxbNGkgQHxaxFg0YHjBy9T+sMXXGmnbqNNPLHb/b2wpYp
fVQyI990al7oCsbPN/syXfFdY3+yfNW+nLX2yVMNVJ333KI0oCdxQhvBHKr7I9O9y2xm8srMP9zU
Lt9UQtLmW2SdvNziv3ujEYBchdLnGWLGtlS4YEIzcBaT3IMCKbVoDjI7H8yQYk7rbzEZsfFslC2q
0vXTTTFECO+iX/KH5HyU67pEoU+qV9eH8ztMQcl2dnqB5IpO0OHJ44a7EW0z1SkiUgcF5hMntS8v
RcdQjVzV20d9ldvLzAmpv76h0mvuOD2TpfQBEYVBjvti/zFfEzeT6Aj5pyDyImWe4CXnjYMhyhZ+
WEvWG+dIaplURs2YDpMAgjEMLJklhrUQ4kfivDTXlXVGeM6MAGODKXp2OvlPGN95MY8E7bhc/Ab5
kuDT4Qj+Rj11BPa32xfgE2T5YRPq6fz2mnzXrexMQahT/vLn3/VluUcZVzzoulWzogcQQJvqE/au
lj1PucBqAWr7eg2XyhDgVfGBQVTN5IytkVil68oLNbhvDJbKFa4lXxaRwEgzd62vovn8pEYZ0tus
u+Cc5e1tQS0a39rzzIYW+mKapkbQ1+ba0ZYw/uexSOXipg51gQ6Ppo/FOg+ZQTUgwOaC+RdL1/TM
0wzyjQoa3o78iAH3jc15BJe2UAXFNpPhVN2qtgSoxBKHGdUDEg3j+Mai42R5h6PuvunPMigGe0Lj
KyABkOYqIcmGgwZYqIvB1fSp6jJVxhrGsL9gLIejjw1rmVdZIeg+/hYMqN5mR0f0T3m1KSZVkYnP
b+lVYxxfE+e4kaVSoeuvwciQhaGwPUtmDVyY9GEl8S2gS4z4wslcks/YAdJpjUj+olZzx4E7p4fC
vovmflfWc6SpVav27Si0cpbLq8oclttWEaAvzD2maSVIemosGFp445TFPm7FLyd1Nfmuy39IEKIq
o3lfKDoAx1avn1x4KMWtN6zOZ3mZ2YrHXKzKkhjXZ1MuzvpGP5UNpsFsuVD0pr4DMdZR+mJpDvI2
CpFi/UjdTL14RpUX0nsUl3Qu1t9B4oWict6iMODO2j4R7TbBIgQuzCTt963Yg2MfziW2e82kMuOg
e+Dqfk08hGlKbJCqbO+y0oxRm/EMsbQBVkcnKyuf/4cyTLdZrkE8Q0aN7LaI7YyWHHSUWzczHMkX
hMCf0MylAY2hwwKbnR/H/+aEdcM0gTZChAWFHRotu+j+IIqawFtSNUXHHpHmPrmfMlt525iitMpW
58ammDOnUO2DG3BMnW379RWBS10ry0+KeYq60FAofN473fyw3eRMgIf9aLoEjIwUFCKcKdoQ2AIc
u5Z1z1a3AgR+SvJXG0f162c62EGn24hlY4XTu9EeebZ1kPRQxFHGWSB9buw4DvKGS9+JGhAoAGQX
84hI4Jgq4r4JQwVJdwbj6qezQfKrAp6Tr1iRVgqPCAOQ1/q/uVxucWQ1oXdRhiN4NP8cnpt5PfdQ
l4ZGvh+PwaeAUl6RIk1ItFgtHM2O+kFKzUCKRKaMquNZk2sRwcQU619N4lF5vhJxEJ1tzShTnQzg
BrCujKGVDY0pqxLkpntyvLaWrd8kcx3I+io9cGYeDNqHsoNGf+7PPAcqdLOpOrnw/BX1VXcuHfyt
gfWLwJYemHXCHnCpA4kP3Gxc+2jH0QjSinalt02MnJoOo87vz6pcklstimH8BQnYfxaKBgtwkQyp
gLmZ7fKqCRWNynwPfcBKwkuZuMH4R2suuc2Qpw+hMvYEsRzoTV73voh2V99JXQ67UCse5f0N+8s3
Oy6VXFoYQUJCSPai6WlIywaAPfk0sfV7yJVjP3+h9tl287QS80hrJOn0StLUoaZ+pp1cShOGlnD5
lm7MBrAte5Ug+tvkokBGtd7K0ZuqeMjxZwVBPvGro+2S41if/yyvrVOXk3tKnxMaU63zF0HiN/kI
7vgge9t70MH0S4StpWdWPgaN2vhuRWdhBmqMY5534ESmMEmx28kJiLUxnxlGjJwPxyY53xqe0lQr
ImbGSRZ+OQQaDWKT5YEf7atNEn1nrSjA7ScWQsf8rex5dS5jfifQCrWqSqEya8noml2w/5plTUhH
zbY/ZWibblMTqTGA7XgcAM1jMLXcG0epSHb4bfWBQbwqTflb5KJKi57tyGLXRQXIs0N5Gjvl3Nkb
pidxWCB5UwzF2NI33/8a1DqHJCbdiPifL79FUQWLIkFBF5o916cfNtCgr1YegeEp/ktBwM0+JyC0
EmmegdHIyz3R6u0bs1SA2v2uv37nBT2nA9wRVC5lxjwUe4fQ0qagw+SyWfBpzL6uQMwdtNR07WPg
qvgqvDj1QA8fIpPrKjYl19VnLgwasJ7sklCqQOytX8KhGP88U8huz3zoterJ0ssCVq/VMKMAZDU/
1bh0/+DsXVBiXiDbgmNVeSG38D/ufdMeQNQSonRoMd6gLD7h1LqITWF+Y/dD6An21DfanPlYMdqz
VP+WUG4U2KUt71bQOwR12Q8hIfvgT8yR/rkXQNlIP1B8jTThT4OXZjsue/xwt0WhdQdkiEZJcyNL
SSAz13SFLt9TMiJTlIX3EbpKhggc7PL3GkTZc9lWidIP00PdJuKWECw8fkTZyfib6fTaDJNH9/zq
zMNkOqoYOeSq43gW+sibSThS5i/u+IutGUIRx80CLv2BmeNasfdt6GSHj8TZ5vmA7sclTtx9BhKa
HGk/0A6rVOSNiS0Ngh7E5go2A0WxEcghqD9U4JxJVaWJ7cdrURTFpoKXtnLhx+3pcCb/i/olcGmS
ioAYS4WMjB6w+7Zfi43y9eYZWEhDeatwk9djv9HGr6hYATpYkyYODSdPhqcycU3ReXvIjTmEZJ1n
atap21koyaBsml881qHcSay6ECJIzE9ljAHIcps5PZ7hF8kgWMH0327VVJ8ewTkIkCy0Qr/7D8bZ
bXvAc7lGoDS4s+wL8+fZOIhHJ0fMYmOF9GNXKBjrP7GKla2TyjVl5Z8Z/ivoPv/uZVaziRjWSSer
NLmkNn3UhI+O6HGel7E+xq+F+Bx4L1b79Fu2WX+/MaImQwN6iLRvQgGs9DehJsq97MI2FqL1JEe+
qXCjp5Dqdkrtvh3SGZNYTgw/s5Ii2M+naDFK0SF0kDdwqn0Kisyl4UnTyAjf/buYPUBlSddauqb9
gRBu9irqaBPGHQPoBz48cdHP69DF9pJMFYkIU1+wbT9gHvth0I1KJwWz5vatxWmCcVgl3ePjxXtu
7Gai6AQu6vh08cpLukMQrOcQX0oYqI2Yn05yQFMnIyOAA+iLyKVhH9IJPaM9F3XmPIIPfjwFx2ZS
rfyf6aZ5huvR/YdNG/eISBweXh0KzsgEykljOb+Ke41/zBTKuloSuFCYHEROozwNe3mMDEwYtUWh
WlId/El4lghssF8W1FgmuFrzl3NJmYuIQJqfLpnzDjSwKjfTfIXDYaEDaiOoDPKdNVma4m6IoKQs
bU9zVtMG660IotsLKfYr2tAW3/KQKZfrpaZxJYC/7Fxi+K5/kSBtgAXmeL+02YcTfSSU3pAqBXIt
gPKp4y5dP4pywjDdJbguoCLq9TU7yxl2SBiCastjC3KZaRz51cN0wJsULAVPBCiowOmXYfFjmGfU
gaIXvRj0duVVkcaMqDw6yNh2f5O6h5+R1/zK2lfsf8XFv0SLSr7CzQh9W1StThfRJjeHAmaETkVy
B+7SKP7jgZH4zSyvWpCNUKQhfSiTU1/6Hm1AZanJf6YVg/4XZaprt1khq4vQH9evernQV6t1e1LE
bDwVq2eVCL7nqkn4BN+y2zZqwhvCnF2SKfsztj5s4GOQkoTN8z/NtOBSqmIoGy85d4xnlTDncE8z
GiycwDVx4JlFqh1ER8pu9L/YIFkY5chbEBX6FMRlKQ71+DqBZ6LKEsUnoYFaPWV6HS28WLCdV8f2
N1AzNfrclIUkeMPfysCey5neBrgjwz4bz+fghpzgujlqDc+umGmUl1iKQXqMDPSBMZu+j5of3K3e
BNsBYQGkaScbnVtixo6bqfy62Ol5lHCRKiZxlJk1PYPnE0r9qXbMsi17bIj+8EaUaAkBD3bkfQKz
71JEtBtofX5hahf7VNgxhIz5BY0uOo12+1ZmAOsvyq1VutuwoTsNtgHazQH2rByVphkwNniCla4B
1qVz8LINvm7tp+3sflcTq9Vu1ZkgKoN1U82DSoOf/YkRztKmc667SHD5l/dPqdKQFbYpG5z8BZ3g
ZgXwQAP+HhDaUThiciy8+onbz+KYQ6jS/m47TDlSS//fo9ixX8fIKRk+RoExRS9g3pfdKC/5UlVY
/h66nSTw+7yanwXZb4rWt+I4PgFR7H+ToGuFHe6TriExX+CRI7zzXOROdQA9v0U3goileYa2r6/4
iPaQjgzZ9MDNRdahYMvUMjDCJ+yuDLu2HEuOP63DE2D1kCmTuZyO4DFppDxWAsTvzihOD6Ppva8i
RsQ8BhRMWCMuOdrr5XJqwr5CPmlCElzHtsMcb5E/DXB6PGox9P40o7Ut+ewLMDfnXLZfKEmZTbtV
GmGVfsDlCA4wsU9xD33E6B4nYdyChA7TrG2tJjLbxwEs9HRv50SHxO/F2mfBfFdh0rvJ00MOoSJ2
sJOIwJ2GWviPcgMDEN/MFEWfgxcbApHoWlcIBPOK7KD73sEkAT8QQucxP/3RYcso95yizT/mLs2g
udVhazLqmHEdu6W4+2A2k8RoLYRKcnjsz9kIzk5xi9rg1sWsZI6b8Xlu9w7bw1uwGvjFbDSU/EuY
Zrpu3f5mmY/nKb0Re4Ky3dwgrcBskzw5QlVkyjXXx9hXVM1U49xpOWzdbAWndHigZnTuhn6qzc8e
UCDKI8z4hSWw1iprhsCScWF5vU8O9ON4zz80AUsfSz7cA2tw7iG4LklpBEzZk/rC5AIZGP18cgfc
436pItYiWtR7CrPzBgZthPMSu8DjN1WIUeBAQ9WrttDuc+N+D1ChMecNKtsnKpfvmoshWpjn2KCl
GkvJaCu1o3/4O6R88F+eR8M1r/L4IaerSl3UlimkfNtH8vIM0tM+HdLOCZgYoLvQ2HRiPRkRss95
je/KwrfqHW7JOWhcni932Tur2HBsGmSN4V32DXfW28daD1V7w7l0Pqcxgou8MVwtSC3IjoE35Fr1
hfC29wm4zTttCT1P1MLTucn+efi2paHMup4h2BjKvB3hocwOFAue6WBxH1GERv+KjGTGyXvsZFQd
CYyph/HzZySG3tOrMvbqmKQpEMtWJ2YRKmsTqlsCXF0yIoEQZt5Oa0XVIO1B9UojAUhHU9PTA2ZM
0HjNtaY4S6BKFaMMsKkgFS87VhST4Goz7Dvz+wrcrAndkNYDDQnYvt822xNlmhmCPi70Bcq6b15M
Q7XUYmj9U4g3usSi+JMVPMEbvEdIrnCUDRzGzpbxTqTEhP4BnImK9G/JsxGaTyBQlUCzGesGBwIb
QOlzedjIt0nC9L5SJFsGpRUQj6vvvl+U1OZbxxmPsr+9GSjaFwkipvKiM18g9wLmSa6KPvlpR2x3
/GRhLN6QxncsT6zdUxxmD4TV36Q2BFiHkV6FFx5alYh4iRBiwyr2ZgnnCQY2TlVhzl8Dt4OE8iyT
MevYaQ0jnF4KpKB6jWRQF8wPUpX86YdUqvx4VN4Bky49r6RYcbQCDYzwtFdl7x3rg2Pn2PKvMTgi
94lrfFCGCcJMrnFjbRoxPtGNCxOcaiN++BVbFXVIw9uxfsygdsq0lu00UIO+z77Igjvkev8rjTcM
ucC3c1BsVK5ABkkdoGCmxqd1V1e27tUwc2mMk1I6R2UsBchgHhFX8tX9WCwdqNV0mh/XoCnk9YZ1
Odp+6euc2Wz31Z/9ogJSXW5emq5PU0VD0qNBJFXpsRqPUaPgXAMXvq0FICe/vGqQxDGACIvRUHui
nHEvsUMqIZ0DjLbi5OcglR2KWJ8ev88zi+iDcQkiezSuz9hy3BTM/7khCWQdwihoWH2i1Dp/59tq
Ei6c6Hgr4Tu98eReW5VgrMS7cvlVwTV+bFvxLm2gebS/rh0Q4mWEEADjrVag7XDBbrZfFsImoPGa
6KaIoJ5OXQF2+hsGYYG69NGcRwhRCPh+npSrXTPkOSwd/0mcDBXKgJuEuVtAcFRjNxrdiHbAAIlu
Gp6HKP8IF5K0pu6p+CWk6JmWqgM7CfiF2GUVqKCcoeds27WGAXQreb5eoUP4seuLsto1XWuUDkcy
kQIybh0Wqr3kTzm/lOq3Dn8eVGd2IwkV8o4rEg6hV6hbu0jSJNP/IPHNNZ3Hqo6yO31rEBOlknAr
6urgx8BYmOsG3KLttyFGFWFDGXcNOh/L1wAQtA6mL56CZ/VnSqaCu8dJmefliWdT1CILad4WUjFT
BMdQu4wHeI4Z9cmhLSmj+R1fevkAre3VxsSbGgyj4Dp9UQgrZzgVloDLt2ckf9S3tf7VQDkxxQkd
w2YjQWj/ZKuZBd3Pba5+en497ow4b5ZLJG8EzI0I6ORbqG/AbtTWiIyONUCwHwhA0BUe+1r+GlGG
vmqo5cm72ecLHtKFzlNwOmWgePjSngr3R/nqarMTya6inBljV8wSHR1AkuVTeE5H7x7iG6ShCiN6
8SPHOsM9n8aw/nJO/ggtFgcJTVswDVW5R728Hkmo9hkzzcPFgEwrFN7YhIsu3U24i53tZyPwOdC2
0O/DDH+p8Pu1yB9f61OpPpXJWtAQdLNmkSpOjkCHR3RgGUBtnIFC31EauEBFYWhUYkDvn0XSwaLL
PN/st2VDjARNcHAnNxkH34f+kKqhL57lliFlLzBcDQEwOSk71scejA5pSDpO27oYMCwONZ/cfxEh
rf81nQFGjntgqeMFBjUTCMEG95Aj+TsAl/3og3It0pWRGsoIikLhXLdDuwIOfSmmnznBEJbZGkzh
0yElENw+q5gQgj1K/JCQS7xanOQnH0KEnVjT/pOzLtgeTpLvdo862HH+OpUdXzdteWyOCmg0CfDs
FY5NR/BkizDWEcOQjTRXTJv5+u6zyQNs9D/4tlmwCsnPP0chB854CRh1JvqzoPAqFVn5qSbbc9OY
VxPfBSLjdhG9XotgEtKRWL3WW4ax1L578ZeCsMF5o/xptASWqW2X5Hr/7yLnI8+qXyF/JGw6UNng
oI/iM2mKGSZWAkf/oCYhyjk+qkcNETQje7alLUjmz3TSiM1Jc/3Ust02osN9ddoy2dA7H/cRkUcQ
OO009pBmaRhGMyl3NP5JXTO94Gofs2xMxJfjgf8wuV9WfLhcnMpmw33nJpMbC1hcVksSoZVLaY5r
r6+JqMnWgr4lZFBDlX8SZATDbMVph8VyuefPQ+MCU2S5CRXU8ROB/iG+Ycow80e1leD4qzKJv6nX
6BCsroHiq0tpHrZ4JOSDwoq9StjG2dFl5zVtlKYKu8hm9BHHPl5Ix10xyK8ZKpu3kP1P9tf33e6D
VfBD6SPl4lcr75humD9KwMb4KuIQveArqdX7sCtzWV2adp5Onk8bhz8YYGoXNxkNLrFWy9RNg7r/
c24ky27aR7afKnIhhmAyUWWGRE4vJs2xIp45CtrfN6DJ+dMbpzrZJRZZl92/FVVzIAgeqaswM4k8
m2oPtT+ktxIv4I/8PQtYOEvnRai3pb0ms6iX7l15NNPaITLg7BogwBK9euOAjXz9TjOc7OaDG+Dq
HWN3X4Qn6DM3hLHsQu83vtOew7ZgleQoTwxSvDNoVhw7eFdiiIg9yji9WNrsPZNpQI1TP+XVa1Di
UbYeef3CLzZlMLxuBeOzM7JFck31iv9LNUJpt9OxLGJkEEADJ40T23eK1JiMAsVWSHc0jPH+su6k
EsDbEAvZ72J45Lx2LdidFjOd8sHRVUxVLNCeWOiVd9cbe9mkqo8g0fXSIEaVm1l0YyiCJ95+e4Uu
t4ftYvaEgBCpH+7MfGNpOXZov3PsiRKRkuPybRofEknmJluE2SqGrSSZUUBxXAvNHpRedezwCKys
ryFT4uQsCgohasnyooKIwr5qMZ9+lmjn/oXQluSVbNBY35rMy5hUozd4PY9O15ycHXRt2L4+56YM
Upvj3z0+oObkXR3lj49Sl4GfNBwlCoXLg3r/ZFWDZaH3KmGYFcw+VZmAc3zaGFGBsKQkh7gHjwcT
1QuKIrRBjLDOg/yr5t/w4R7aseLigsArlTEAeB6pKdVSMT2avV3J0UYq5LI+X+G3SDDSc8TplYZ1
P2gLLhGUhwpptoSXrj54Q0YaVUncr+rWHaiFRpDvJbmU+B5F/s7GD0S/e9NQTE4nHEi7Lqrd1CJR
ejB/4bn2vbsAlylgB8FqPYApDz7pP2KD
`protect end_protected
