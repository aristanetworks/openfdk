--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
eLzjRim3ntwhr0Rk8VkDzEKDUgFrMcHrqBMstb/WDBSuaj87n4EXExS0eJnWr3Yweah2jMkbUTo/
S1pCzJd2BL+qJUP/gHRiAopRNQhiwwDP1IZveXezVzvA/+PONa0GnK7qZHX/zpc397SCwdmjkxJO
V+IQSRvq4FaCGq9EJ4T/yuiRz3P824swr1oJ1GQmTX2olYsADPKTONgR/8Hkff3rES9n6RT3EBL9
GFNsVcBL93JqQOhLRLjxTwD6aNvgH2SeOiCFafcJtMuWZSEwnIKc44WlJNjtMvgp6q17ajJiXBnF
yuGgKiogr2yooLhGR9CGpgDvq3cdljjTu4V0yQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="aQSBm2lMvQxm3z6gOnBgH9NVDP/N+JFzQ7SJkgOJEAI="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
pTXIq4Xx4eEkZ78XQvrdw2ESA4zAClWb7NAmbqt0NP/1+a4oFklog4rptvVz21bHMzTz86R2c+Gr
Yp1forB7zCDiGqfU4kY7+bJ8YGqF2dC6GpOCZ+8USk3MpXwBqXEbxPWhHezRKGrHrF5u1T/Au7e9
hZIjusPLEEtG7ZgQFI8Rq3qqHvNxLmN3tz397UUvmYCe4JETo+5Xr/uWqwTkT1dBzxFmwgn1orxV
hlzxVe3qq9bt5XFNIQYVEewfWL+Eom2wlxkdZVb4HK0bFSRpqafWzEiGHvW8qhyg1yzezcvuuPSz
rAy7b9Sxl6BmQuh1OeYrde0dAPlBGnZkjqeB9g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="H6anotp+/QigxkpdogkhRtFnfyzKfi468CmHlOnoiH4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 29280)
`protect data_block
3t5oGj/Vpgcj69zRUBJ5Ubw5Fe3jZuvPh8zP+6l1TcWtfngzFGFtJBbHsl67AWWpaU2UjEyWUGdl
5k3QojxbPiRnNGYkpZ59HVwQeqREX27FcbACMaFaIMzzH984vwJyxUVxGp17s2N/ABTlgZBX8sTV
7OSP/BM26m13e3lT/zhXmSLHE/Kw9U+L8Joi7ivjpKvhBblKfdGcZQ/di6psSt+Kku+ffVXy7clS
19hgm+2Tt495qVWIyyyN1N4rxHhjIOkv8tpDvVYsGwtcMfFIQsJMF4tFJfV92jm1Su376w7dzTN3
5qUVbzX0+DSNMxurVc2enPQNbH+3M1hYoludQFcjFp1dKI4vBYEl7c9Pl/ngcOvMCIis8rMSaLSg
iz9IhU7jiRyRsH3V/8k4l63wkB45by3fb937ZKeyZ/+3dFxqiFcyrsXA4EyHP/txblZMjeNhqk5g
Mhu1YAE8EJmtI4z0PBjPy0sCOaQB8eK+fh7MoHIriygxw25kAm1ElGVkOSR3USXKQqXSZZ6d0pSc
+J3pmCqzRCaX3aKe4kDcZjTAzT3aTvj78rPWhUn88Jl4jBRLfINt2F1ZEeE6RXA2d5swbgbV491k
olApmDqgqbSh4cEzr8VpfWg8vhuEPu9SoQTXffmjT+34z9YHDUMNX+Dq1NkstyLIiWgZAhKDR1V5
mEHrj70tW6P/bDCYrmiTEH/ogp6j0jHLxwvpXRJywcPGgf4CXdKizDBcFbLOlCtJbLBx2ay4MT7j
lsz4HfxSbZIc+pgWynFCBkYvX02CrZGmnOwlXxepEUofZPWoQ+o/Za1o/EQauV00hyj3QhZnDaon
PEFdRdLkPiH9d2J2FKRyxy4DbfHBcAmkIHp5pDpAQZYoD+URqPjr6D7Wu4g9ZT33Sc5N9tQiX4aA
2rl+8BR5FJOo58nilrLF8BWggNKzd5ZDwJiZ8Gi7jOq7JMbmyhsSrIaBEUl1OOMDIjRHikn2/J/m
EOpt0dTohh1sPbuKoeXWvEHdikH33O2565RpdwqZsgfuWgEFq9G2ptxNMM2P2mvDaVqkHriFQCla
ojr1F9iPgqDimTCN69vQprtPA31l+OrVLojy7ir0jLsFdqxCVSTLrQUpShJ/rjw8ElYmt2yjc0Ng
PIVzNZ2oT9CroignUvWlSGxLfFyyNwVN/juQCh/yXLG/hvLJH2B39CvZI/2Ku75EfHBTYKZhtoBL
TA7UuR+dQzL291y3eK3jWR3e0dzTi+P30L8Ei1apkFIczBAuJRC81kLD5Ik6RWnsL96VZvQontuZ
kEl6sMCNJB2K0NlfaUfe7/htgMZXyJ24u3eREW1gpyySW5L8xIaB3vOrjKRNWPUT66rdD3VEalte
iiX9CdYjioqSv2UrtfQHnAKuYkA12bYXfsaHEldTeuWgv4YeoMVUFfxF436D1It+PfA7I4XQuwXd
ofJpRoBGI4CP/TOHKxeW/C5nDQTaIKVbqYFCdOjj7Pofc6DeME52u0MO8ZVzkHCNTF385SOzGa21
dSsqKFaKaFvGKWaMjskZ5dkcXEXOhX6pYLEzO98W8QfLIhH8/bZ0Tdm1kteNSvEkHqkGk+F7iLXR
Xwm4gEZc4QkdAR490Dp8VxUbHe85ERK11yHHp5dXVq+L/MpUzJlmwNw4HCLaFUXYGs/np/Xf6kt0
5UBLO1RRXv3d1bnSr9u04TUPstu5jmvQzaYmK1pCjDGdROg3sUs3H7ilAW/mo5vCHYOLed/kPTee
xviH1RUIZ6CXDB5Ijr9NS0EocJLRxgXDoV7xwAQyMcmNp5QRsnDcxF2jcb0uSD6XFrQ2PWGkIA87
AjA0GNY1Ypx0esC/Y/p5V8aHHmEcH/u8f+I0ycWNk8Iuo66k+w/PfSC0Fq2xZWFdU+IgTdJBUY32
Zn04U7AePtG29TTa+pVHmv5oeevKmA9Znx8WF/m8WgMrZtAbbubh6C82OCrd7pUGWmTQjqoEVxWT
63bqt2xyFlcchKgufnT/OeJvbfgVf52qJtqqfmYvyxjJBFry39SDzbNtbyn7S7G/MSIYuqV0O280
8b+vr6f0tS7qLQZ07yzrgiatEH+W5nQglUah9xSouSNqauSHUiXpsBu9sIunCCbmm7FEGvSz+doR
wMVD5ty/0Fe70Pe+Ww3Pfo0FjSrKasQElXrsSE/4i8OEsudMZvdN71FBhe0pW0fPARF1+2GEDYri
HX6JNyptTMwhjN8kCt8amckgLqSM+tWmbULvsd2yx0EYDH2Dt/ZR8OTUjZdshXVl8pWdalwX6E74
eS3ewhvHmnGqm2dtOEo1BumWimsL+MCigNYQTctjjfytl4KKuzL6bLfvU2Cj9tA6bUcNSMGFvR1e
Tf2FozDqlFsSy37H/WIRwE7KpvVEaOy8b7tZqscHZWc4Tl3ZyCNZtiEajbf8/OKBojCtOxTF8sQ3
uUPo2aPvaL9Xfp5YaRFTMdoUinF3ZVVfq7myP61YrXP+fBT7rZ9sRRLpPdxe6EC9XScRCdf1e6K2
PqIc4b8fK3mV2sA+MUJ4z9jcHP12qHAE4SdxZ0Pbk2EeNP+NUtuVqrauhpHb6qIb2By10uKAQjaA
ZFzqNT3T6LYCyyrmGB6lEzYepDUSsC+K1CaieL7NWLItzty0fqMo/lmHx9w8MNF++gk2GayU3X67
hEoZTm038ixTRKe/dMqI2A9Ob8EfaXP+SGDlG2j2neyQnurx9P+D5jZ2Mt1PeItKGtnERbDKHj5V
uSj3Zf+3Le05dHwqH9hviBuheURmF+BfBIaXEpWB5toEIhcBS3ELht/jcx9bML+PZ07Ocy4zupGc
hNNqNfrhpQr8nlwD0vw476RLYA7EVS7+L6/bL1ruHz6v7Do+BJ6B4N9UcnCqeTislVUoEIziWwyS
CvddgnDKB0NXPsI/vN/ImfBgSlRpxmae/umw3Wcdd3ovHK3Xb/oBQTl7vmfZIz1AX/UcqsDxqaFz
9UZJW/VZOnEpjfeiQMeTFwlHLFZcCK2VrDXMIUVUIVXfFf7AZDK5hyKaHb5lBzUxDJSO0UjAoVV9
lXjFPEFwPmmOzRhEw5GXtyJBLSWXGEe98fi6JYHIac8H7xHZ1emYWIjTEL8CiXdErCkMAY4Rq1As
L7bGEmXSUXmqC404HVzXM4wupVKVigI4Bx6XpZDtSVPNocZ5Vu6zhxgctuMOI2qDekB9BOVfV5aB
WgQAS+EhOtYhwfzIsexk1UprXNVQgCNd4uBrDRGHfV5dcr9eNE1kIaOXWcq7E2KOpGA9DwPrIgg8
rAQQeVGBkL1RK+wujGlRCtu/fexfAIoUDexVl8a7OegkrUNAeWapC5dOoOFW0FOvmRkAbH0gj8oo
3TjPbEs5P5DHus7ve3F0dBgGUBMYHyI8CCSWpFUbwAy3MTVcAblqqTw+Lvihl1kx8DupJHXXPC12
EXYMrUMxPzMKH7gj3xqnJtLSgNL8nU7HrJveW3OAoD3QUcB8ILDK/2X3QD0yHnXQMbYgDgUvXWme
pRlbewhSr+0+QBlJgTPJ3h8qmrWwnZwsDBtUYyRoDhdI5BppS1KTQNRag4doUu8kQo3Bwr2J/m4D
/cXrx2ix3PHz1PIz46U4mmA+dNOaXsvJE/Kus3Iv7QhTN45bMl5ecYdGv0BtGPffS5AG/isqv1bH
WKuCvBppnvTorz0xIfobuGB35n/6zUIVBTOS8dUgSMhmjPvEtBGhOQ/ctHlmHkPiRSS7k6S8pTIZ
9mX52N2Cxx3e1e9vxoebcvhd57UQ1DdwHwjZcWfMdn2Ky75KJDDuTDUhWpsz58YKpacNG7dfeKTc
bH0gxoywYd/cVQ0PejPo6nR1F3Pl1N9fCZ86JwJVzMUWYP92VFWpbBpBU1MTVdJUQNYeOiIwhUWm
F/I/QTo2TfuDHyV3pTgyIrzokvxTifPNHGiVSs963p3v20QAVYQ6dBZL3ay6a8+RkwAzz1j2Qdv7
NMP/Tdm2+o8d6vwYMDyFwzNH852dRysylcT5Kc2ds/Vk+XcYMvw//pR8XfS8C5XS8Cb8twbwGDV9
0GW9oZvJAhLdwbOSPi4V6tcniiNO+VHcwQLwbQg52rQKLyvqGMJyc4ZTWjsB3I5yeqYhuWuXGv0l
srniy8KJqgbkSc6Mwzneem2JffQgMkWyGIMjcmgpq/+rV/+ZH3GuE/h0WmLYU+pt7SQrZOUsEZYs
LeglsPVAqaoJljC8to1Y+wgXeor+wQBMcpZluDstSTGr+4onHIhTo2DGfpSBRgmkXMo5GKEZcRUl
vJOyRG8JfhCA5HOn+hfpaMU8Ot7Vg3ErEwzC/25nqw5yXqeuerj/EtSsPHWrodoGuihvTnDKxGOP
DZTjWHHDHwYTa53d58RPAMbnqfJLTifYV6nnoFCKLRW+uwrMhWx30HKRRlZJdIgyGnQ4z9/2YwNR
tOySDgPtF+BYtPBjpjOS1+CdCpBrvb4IqEzXd4ZgcuLJkGgIXX2cCb2VbqbW7GuyU4rZVIzZJ2Xu
BOw13/Psvc6QE/r/jXaFTbFD314s+pVZbZApqsoO2Z6Y7tGMgFmMB2gDalLr/LQslKREX++pUvW7
wyC2X3u+F4N+2y8LUzzJCdu7mCuV9G48cV9IvM5RakMLH6JLiMrpJJIQipxS+FF7TNxp5/X0uGP1
DTraSL6q972guCPDKqXA+QfR7Bfn82h95Y3217DWHBZOKc8kEhk4cSo/qj2b4/flxZYGdW7o6Clt
y4r8Gr8pHpgtgh8XlsAPf15RgkZl72sm6tWbWa8ziX7wTLwmezpmsMGWBvOfdQpX8wodx0bRUPNE
rLSQyHIHi7Dujgg09sLJs4fpn+pNC6kE6XY6u5dlg6NDlTq25h25oXw3xZeeMBZTDscgchuUKT3u
3dGNJbewwVl2tRNbybG8Dyj7A/ZdlxdE6W7B5aF15kPUXuUHcG5SksQRIk6+PYlF22E3AYWfjYu4
1nEVxQ9YY43W5RbK0d3n9bH8agrxJhNt58UoJ+jpfoJWHK9mShG6vwStfuPE5JipicUTf8Mge5yJ
vRySiESH5JwvxGibdPBWXp/+3GxLyTlzfkD568pBBANbGfPQ766OqEgUetElhAdkw5glu1LwA3E6
qsQ3/8leylXaD5x8Gunv1sjfaAalwLmP/s3Xf/dBO/KO2uKu4R7uxxBsw+meB74HJCemcDzyt8X2
ds6xC1kyKvLt6c7i7y/9Dd0y1xfQvgNtbz9f6TYE5wqKVYCOwrPUkoRDj2tW6pVauVK7M1eVOtcd
x/xyVRtH/A5eSrhNjgp08R6FCo5S1Ha1FyaoKwkYID3iyX1Fe/KbUCuLS14HgOG5xafejIJzQeFM
z+SzuIRWr+dkiKGnya1B9P3rG9liWUE8EFkJmwRzEzJAQIbVS7qhWBL8TS4/3zfVg0ccPGIOuvpo
2iOjI8CHrvjgTR7UQo7M9KcqkYxtMvLZoypdHc7pwp6ZRvLbSAmwIhCBHtJCU1jG4ZAO0dedV0a9
PFv7IyajqOFWRwRYOS6f81C6t8nbsixEJtuNJZFbt5lVsA7eoAhAMQkNQMy+JfVhtnm/TG5BUOap
r7VEBdvqrXb1jjRLNAWevMNPCATxLTbjGQHEPNXYizA32xCsYKepkXXja+bRydJxKlUw7RZTw6Bn
yqewAUB5Y5poK8n8jaWn0SSRUhtCVNBBo2XlE5LGYnyiKfJeRtvvo9CSp+dcVLiHHOv+Sj5oSKdI
ft0w57brc+DJR3omM1C0R0JU3Pv2tNmWsCtYZ6BaujPE+hd3Yy3eYwSmSIM/FvlQSzbX2mfgqE9w
tsjSN7kEr5+L3dTuEjyW5D/p4mLKseOr/ItlH59JqqNf7UTiK2qCtIp24JGjG6NhEFtexJpkaC2V
7fvh8HLm/RiZbYFYA7prFrXbrhgAndkTbkvSgfnbFziAzNna5sWCfeVoZfdEStno1QgVBvWFwtnt
hYWN0MAZPMMhKmLRHPNlEW1VorvVPDqsVb5bYrT00Q2gJFzjI9AGYTWm9ual22/N0KhtuC7oM/dh
FZEnjbZWPkksH/DVJP7pQmMxeioRlGv6yIRESSoM0o0gw3B12JRang2JSfs6Ld+Y5bzkkimpMAbM
rXM+tBEDbZ5On6xYZjD2FRRQXUBEQt/4iC9K72gG4jYUPEEW0G18yyZnd3b8cVnwGqblcisJAc0K
IiArYmRqvFl786M/Hq6shjxksqnWHieJDmXYYpholIirG2spEXLD9mIpEboCOEO3MaSCjPW4f2QF
Lao1kzW1RZwIZRKT3CsTgDdHbyVPCBG2I2ejSKv+xxBoA5I+2QGsJFbxZOVYbYYpc8j8F9Aftmmz
TwOsz6MouOHi0MHxnU0RiJ4Ysf2w6cEHLAoEFQw3LVj6ulSwSTe7b5RJuTLJCfLOJpCkZdrwwHY+
1AeeLpyABNmhNVFf9CrvzXr03NNi4EA6ItFDcrc1addIN3VXXessJVnob0CMybAuOzTrsvpqtI1W
81mNngTaDkbGfL9VYmgDN/CPrjh9c/aRNT8KsWxqFzA3c6vvKeeDt97s5IMMCVomqazRvVvE76d8
ApOb4W5/b+x0PYAKFinAqshM3kfWqWSXfWhdGcpAwM5eopHoACVftlQ20bmgcZ4apu7RNUFILGWm
B89eICpoQ8zk7FF6T8OjAsTd+hv17lCjL0Hl/8TxxvWV4PMJ3lHNutw8uAXafghRSft4xN/x4VI8
TCoCOLSkRaMVIMgE0e1zkKu9tcLHYBJGVlSfkNFAg04+xZjuzvMomvrk+rehytM1KJcHeOqrY3h8
gOJMnP/yGowL0fj4s/+eGK7noHLJGJXMeTs/TY/Ewf74xknJIyNlCPAZ+tA539zyrc5g02gS/lzo
bHoa4Nv5r0bgChvQGtMA7idKt5hxHR6WilGvi+q34bSArUtUHO+I7BO1B8LjeIyI/azM8C3QYCw3
3kjlw+f3+2tPjJgXrZdmpUdL9n5E8dHzn6b61aFaM8zPs0wMioK/wAb/k15KPT45dkZnbJjq1p80
3lUtM2ewW5/4stlY2KnRJtVvc3ea3wZ3fWZleIZi3/bcj/Ct1HG91+LhoG6C2C2YuUZXIIngI/QT
pdDFrcLJIPgC8nyadH+7QEUf9H7OTmTzFllUn6c418127A1aphOGSm64AYyaJ2MCajb8fOnpSj8g
QIcxtYBQdlzDJmKarJjrtV2yNpxVOVoqgJQytI1QDb2YH+LPljoAx3prYuhQE7+5ntnFN+TY1Qb4
itEJCwufP87W/UWIT/8vOZQrCdnko+PO+Qy+iJnP6pO0FE6v2/0QzL8ELfdwemV8TEmL1XmlaVw+
OB/E1ByMFV6DEoT22/dZjMOJWfc2Fu7n9ha53VpVX4koLz+nTtoDOWQdfOmN6LGNbucrdQhlgQdq
UrmYfzgo0guCs95fxky+o+bVA+V/XvNHgsdL1Hl/h3PSil1mbwe88O/bFvkgXpdoCRZBPKrDTKfz
EFqTlafrJSO1yYJYSonzaI9SnignX25WY25gv/MWjmEFQ0GpVY23EYSFkEP5BB8v7hb8batMYkTx
IqkgoNiZrjSbsNiGzrK6JD8X4DK8AwGyaJ8vKtfUHjgbGH8IDruvnF5wHzjRlNNF42G6/W7hafW1
Xa0H1+rWyMnav/5Sy09tFNTwVRBuGkbwWw3rUeP7qwQXaRZURdSu69+KQ8prkv2a+BP/K+T4tLNv
464ENcJeBVAcQYkgv0MY80/wa2Z0FUlQZMdIPxZskjQk6N7kEFwLEEjNAelDERyiyaXcglj5/f7c
8BwU9+iN+e3sLKur6ybGf6oZraft0XND/9BqakqzABpI2Tk/lPXiYH1IXVdpxnu67697QgdB7Plx
7ArXxDxEE1SmEzvZ5EWl+WSh+j1tIHxlO3P/ZrKWlsOPRQd46drkgQJRTRlY+sil/m/qzpSuCqls
xRlH4GD9HmCW130mesgb1CC/GYbu76fF4KIHIJzda/fr2V7CjLfxuIhYlUZIdr3tbyqWge9v7YTM
SayF0M+tdFhXrjvUA24/Co0CzoQvhiQtcr2GekwJseqp3ECZOZMy1jZZOeJUOcpQ+jPkO5D7oRC5
0WwUFXSzTu/5hnb17nqO6Wxg7+Qt8Dmfxa9AVhO4K9OPOp0nssgqFg+Ig21P4AYMrQyjnqynBheN
6cZFURBmb4aU0cSDiPcz2ty/e5kKGh6CODSle4rHAr1NKqVXC1g3/zhxqWzS/IAHhmNuSfvkTVEP
fW2nJxbSlfnP1y2InzyN25Ydal0uYWi6xiwofE3BCS6M/5Xw4k3A2QexpBEHmnindrZ7568ddmRP
0giB30lDgQ05QRwHZKa/dPBOL5TvLhDkw6YqH/IizqwfwT+SOs866kMk+j3J+P9Iw18sfymiln2m
Fc+L81kuGEoM7LN77uTyZG0sG4Ae+ErKjrTg/RCOCuqdaLfDW6iQ25REQ1d8DqeLLSZketTjkbk0
lQdDxN5KVDNRc2++1wrcZoCmGv8v7vrr5ny3Q4fxdzV9YpIIoFSzH6C1kQLgZm12DDd416/PFO1D
osQH6cxFrZJfCXmoYIEfUc4W4MTFrgAeSqTKO698iq4NTvRy3hzgkS4z8ES4XsHdaxdS3R3apZHq
5V8XAdlXRZtIYTAP8KoonaTSD1ICvxHqFETw860yrPM4/Kw2oDsuVqFd42h87/qvdnHQxSIJ9UGQ
EBmHvXL6rfACPVY/Hovlt5KE5FRl6mCjM4yx1l0TE2qkxjpg84RjdRkIlzXDtiuemyTKr0n1LWSg
WZvFuym/eMMx33pKadEHUjKg0NNhcCdyiY2pHewvFTKs1NfoxjfIKZ57MBqZLO2ynWXNH1Em7iye
InlbrucPnkZf0QRwmzXK8dJCQrbooMD0tcQVDx7IeFnxv13nsfYMaqwkYiFPzxpxIx8SmIfQXKHl
NsW1p3YArMDFy3vtr7h4Ebc2TFOJEZS439dvFtIhA97CASUv34D4Zz1kV60G4+4A37l34Acfa4Jy
vQIQM3EEjN2xhI0vAIRZjiJSk4bXwfRSKvxi8llXim5dUhtMsvx2GWsfqWwmQF9YJ3ZH9UyVDt/A
KD+nHsX8WcCks1UsD8k1cnMulTT76RlySaBaVZdLyKMfebsOSozd7KUMXuL1/ISUPo4rRWrMu+EI
cdTwNVbeGMQXbTOeT8oKA/Ytc1ecHkIIpf4yJAobYNcGTCub7BkSNGjribGtLWePOlE7DiNRlck+
O5+EThRFVFU3R5WescBS3VDXg7R8Kw9jZwvbquJC6WFLqsvlXYK/x7m/brcfQ+/EO9HD7qsrERKV
2Ne2vdnCX+m/JKYofXUZjLau0fQLQ7eny3NA7JrbEPrt06EMeuc5JFeZcHLsmkI6ImK0h3mJwTQo
+2xyPAqP7Ljf1AYrMVm44SIYdtG44il0/nMGHIQ55sdpYIfbeCtQSTVl9SElYMlU/Hmt3wrbuzG6
7JwjCwxQ7d2530q5I9X2YlB4qdBJm4KfauXklEfksrNhYNZO5FQXNA/btYfWtymmwP5pet4TGuZG
ut+FGyGVhRBj2Au7sxutHnLalZD6xhTdZvRi19zLR1h7aRWCAuY9ogIWqI34wlstg48IU5cH7tT7
R4npbwj609DU8dLvD3bXjnulFV69xDKO8tnoFxTOGgU0mC52ZLTzGeShoL2qjMJszI8dlvHMtv+H
QLgSYRzaBtpg9uI3WkLpuSzCwhbA0Fu/edy66bxw68T9PkjuL9bPwOZ8I3P5ZBOd+GRvzb+5DSqF
hAItx3rS32aGdu36FADpqgyOAih41d5T65JS99gXOG8BE3yqgY4/4/xAVvyXDonaiqQ3Fq8EzI0P
hqKgsx7n10C2SI6MuojHTmAmr8JwkXrKLkDHlK3x/RR6EfcIkuiEgcLQGmXYvrhc49Mk9vmSVw9W
04/Njc0E8jlErpnRcaYLUwWIZ4O56eNc6WtMoEfEHZJ4we48GFLY6FIWRj+tMuyJ08vdMjqeHgkm
zP5/Kvajy33cj8aPy9Hiz0/+ys6tenko/ddXKbDvR2f8R3paruIbArrNmqmjk6bbXcW6XrbrciMx
lzCSLi/09kHUbUBXALRmAGY0vRodiYd8GY/imHSUfCB2OVW9ImEtO0abs/gxObhfKQ6caWwSj06C
TcF52uChvHJdC8goBHsoRmLhUClD0S5G7i3W+sIkocX59LBrN2PkmhJKIHuVjlZ0w1bnLKfozD0q
PtxUf0U0y/GsAjmcl3kNFOTnZFYsDJqTzvn5c6GRrRqHz3650IvpM4cCybavRI/UyeBEWHbuBYBY
06ETp76IuEGv5c3hmlVFH4+cOcX0houxL+JcsBYrRVL0YL5cXXyZtVK1+K6B/n5jb6c0SphOtF3B
PzKRnTaSjakmpc0Vny4GFt6OAJTgtKI81oiVtKF8t8EiIKElMGuNhoYWPyYd33hzOrxVqKdkkjkR
gHZjpHLmtJ39yplI62DjhpX0kUTVW84dwh/oM89x1rT6oSPCtdplLmSpr5BLdA+d5SIXh6vIZqFP
JiRQorQCsfKA488bWjWkQ4L3kqYDFvpaEwfQtNU8F2hWXCzUIdOAhtngUOw9IL08Dvs74dVmz9r4
rOnib2GvqllXiZm4qdaJfrRUv6KMVjg33uvBYvO8tF6VxV9BHY/jpUNgGE9Onnp0Kd5nR7xwZGey
G/Uje9KjDOnYYxGS1IKY4G2630IzWn4N23NU90Mn6gXAayu2OaDX+lFW+nAsqkhMUQMJy0dA/ERO
hLflZPpPsdlF2EK3cUqcNlRhgv65mieQIZUbWr162Jh6c2YCDV3i/lfi+zfvj8BkAAl8Zu60liCm
J476BGC3GiA81UJcFExGhmHzmS7JcmGmRGpdD9mTVAKiZ8F68GUO41ykqfSV9IlcNV0fhgZWxAYd
l33P4PMcWlFIebghNwp9oQ65IIlDfPOiz2a7Rmm4DaQo2nmZLJH2LbTnjNxYOjqV7NorY1c1Ede+
OVKxT7g3owXKAthl/oaJuCw8fTx8Nlmgwp03MLWOm/KqbUaTZuScAMw+pNPfudO9Hh8NA57nvmhT
B8SdRpUklGSWD1o+fsHNiSxr9vi+/bg/8E3M7UZL1s7W6FZAlltlvkPBphA5wNLXESEn3HO5ck7Q
VYNuDTnRwLGMx+3jA85nTWbi0/wgfXoJ0Rvb0Zg/+621daUa6Ps4cVqMgdQ2xLzyQcGs+OjXnG5F
nylAbeDhodBgPluyAYFW0fxj7REuchDPFMJEo8//OM9bJWCWfs/ESSTMPnK/jOJRXyKpmmb+bJHQ
RWyPdTsHlzd9HHMXYQfVhAHe5XCRYcrl036ZanEjHY/Im4Dxy34sXvKIW8kXmiG+BUgJmseHt5dC
k2AJlVtYamCkeRPaw7VECLKc1xJXtFyjVZkWfE35n6uLrJCx2JtJ1isjWNL2RHJ9XsZg46Cw0Iue
5UbGifVfeQzKcDN/tc46u2mnqSkqB7J2fRwyWPdFgwG4I6QBsOwJB+kgi2vpjyM9ez50sKvHheaC
Up6bY8wZASCGCX9DxggqRxo3IutS3CbrLkchsNor55boKYK8Mx9qOAJdOq4TZfzjglWruuSEL7Ya
LslNhs5Yf///aOrDH2QdcLzR+hZajMgB5VI+AzNXm3WnoQPuM4N0vR5pYx3t2uDiTaVIpiFBMdr/
p4+BcwSVyI/0RxkvJ4yIjByJNGz/PvkH0Zi8hAnvZqFVDuvL3mkgWTcApTIb/A6rw7TR8FwH6ymc
Fu5XpuyREAp4oEzv5SfUSKTYzubkNH/N6lA61yy/PMijWGeT2882DANVLW0HtGhphfOPzh1oGbGD
OIDiTqHzQdnGArb0X50IWXuEjc0g5dkj0EGh4D5T6ocVCkie2/9kMYO2VKy5/nGXpsYiJsxVYldX
aT9Oi9yIiPGD9+Tmsh44FA9/dozPjLTTOWV5gz04WMjwETF1cAeOPRr4x1dyGPsvENgV+TaAw79X
U05HK9kOMeMP9MYWSdIOi2l0ifWG/WTDtu/tNfwzlK8cPRcnFN+Dr2FkOcOp3oRURh+Kd4jaNKL6
XbajPdJQ5d7FWb4QkHTmJzxGxP13isUt15lzKK4HA19uDqkuCve5v58tA6V+BRu8KYNSTK9a7rQy
tK5LlxhDo14d0u7Wn8Rew4/U71VZgw5vkbmkuUGh4Sm8WXfnAtwmyScjdyZ9znjWE7fABB3md3QX
m9thLxiJmyqfl0QwlOvl7bX0VmBj3lqyH5wsgeOshKFgMBiEjwCklVsZ3kK7ksBgsCV3dx7wgyZR
8KcHaDynt2y3Ihwvh72zOaqc1wAgpf2aMUfCS+8N3UDm+cdZO08ticjLLKGBpeRqdiZsHbLvsAZD
xHV2U6Q/S34ovlJaGJVoUQMLl1aiGHphExiDrcYmqs4MPv1CMnYr+79cGvJuXKpQuyD0oz2Ld7LH
Q4K9O3iRufioYoNdvR9/bs2SckeZekgMyIisO2BsCRGm9bUJrjB5AzD+1xCGhnrsGhHdL3lBaCb6
SbMMYH1tWE8F/bhlsKcMopCyx7/dHemVslqvBA1Oi7m0iLN4JyeVwNq4i0rQk+5Cr6360+iJoxQk
NyibbLzU5j07jgrtCE6Zuirz5B8AiEW05JbvZmMdt3roHASAX79ElYJFIfKF0WN1HjP4EJbuk+nx
B0WanpM+4Ze2n+JryZ7N6WPSbWs/upxzi06CYr+o7KJmZnllp0yh1b5u8JoA4LI5RBtoGl/CTGgo
IpawD/gFZh7xPxU8mftXZQAnpBmvJDB4iSv2bECbRyvqJiMWrp1ir8KQiSqjTEceDpWKVSUwhUt/
at/nRLcpQjeiMuCojFpSP2xc2RpN+npPcL0iXAQEZXnZ69yjumh+6fNpQE65XzgDwDoqe+6BgawW
sZ4CeC73hNqGlsiH4SRgCYKzUwd0tQQND7iKqqE1LWFVHGrer5RN3AB+T48v3X/rZSYv4aISwN0b
yBYn5HR6SZBTCLD1V0zde7nc5p1E4Lryy9rtWkvBV1jWxAJP76sBor6vEYx8gM30UF9TpPq+KPvW
Mzm0LXwFR51qWbzc7j87PY9oo1C/pVZJyyLC/GNNvszI/LOLT0uX7BNy8QM74Ax7/MuUcxNxaGWc
scLuhokF3JXxI3rXvDQFPVhHHDDE8XKrz7Tkv7UqjfP72aF7+JeuMDyt+JquKqO1M0j6LakpmKEi
xKoaWtclVpLyzjRVBnoXSi+ZJqtt3qervUqt7Oa0qlBBgI43hKTezQ9SWXK+yYMBL7Ld/FUWMKgS
HOxlEYmK+euZs8FaQg0R5zCqgw3n/mIItkPcZcIHlW2G0WUrtKzWyDXPLy25kjvLuAYnFOloyAdH
/OV+wKZnnkSiy5uq8D6cA0fXIsp6m6axN+Id2qmLDgcd3BJ4WVBwlk7iKj5MN9/GGRyh4X/gc3zs
BWiTrX0JXCHzwvGVZGd/tOr0J0ALuxeUHFvkiK9y+Z+BqZyTXXuTfCOPXJDTnMkhbmWAYSpmmHdA
51Tj3hfGoZWbePkEGtTX7Mj3pclv3OzermN1IHWCb9QBue8Hk/XXulL8X68nkRgsGHYN2yDfRB8w
qRHFspyNUI4mQIth46Y2U+TwdWxxWZnLHv5EVoZUUwHYZkNNyv6889Ym2wi2oTLs1au2rKet1upn
u3k6SywzoiOeepQtQYO+FxPp9UROwS2Z0W17i1VOzdQQqVqkAU0JqKm0Pil9ZjYRRYsZ5Y/dKBw/
llqbw2YtXdRcCQzcoOltZpvlu3sJBMoBh+wa7936zzO0aXnELk8cHHQCnF1Ucx5rBC4F5GwnfVo+
M/lHplcZpzEfujlfbSqmieuB6jVHtrH73NKKZAuP7mXwltki+0GQkbvq+NxNbQOHZ/MxYs4gN4c0
ohtuiXlewTCzzDm+53+rfobtAaLeB1mWALTHKW8EPvmqVfm+YR+UqKrpy3lIkqGUpXr5jSsbolVn
F0s2fWQpl8hCuqfJSXZ6oAvJYjqfHL2znpgNm9X+NfU1x6Yx6EsY0oJAm7ckG7DcCYPifWyQTeVl
MJhLbZRjmrft5+lh06JqBYenkKkYd3UxhT57aBGywfRF7/3rCvCoZi8iulgaXCXqPBYBaDlf+1Xj
Q5F8nqLHuJ/TbHrcqfwyYeZDldzxfTePbIvvb1WemknYOEhPLtT9alzN1VI4lFAefEYG0EVk+4S1
OBoZyh/PvfYxllcjrhX2rkq/XQMoflVe4myX1aKs2lYW2rQmwzAs7DBzldLoqXDtPu56KLyad7fj
vqRRJVOE5SufVpbLhklkeUWAImbfNJirON95aITSVq1Drhs6i0WJClyNCLWm6RCVA3fnCDQg5jgk
3e/DHxa5KFwzJoUbaUwcsfZiEgYyoIz9AbI3eUUes9z/W/iXfAblwA8+9uL6uyVeeGmCtaGcRqD3
+/7CH47t5apgvOjzAfSCsuUUKIgDEqII010X5bvgWs5P71Uu/IDW1TqAcx1J55CjFuxtUxQo4cni
z/JSe4ALT6d/NUIwFa1ui/W5/bj9kRo//Pn1jC8bGjw1TxX4VlVyZDOPd06Mrk1h1oEvEvAuV5Sw
6x8ymPUL9joyWZ66Gc3rPhqZDNRgux5MK76b2oMv1Dz3EuKsPoWHFMtr7Rk/y/AMXeinkEmqZIxY
VAD0j9ChtyArPSvQvOw+2NUJdEfG7y4fFnYdH59srL6yBvHdoqw5S0WYYpBcZQJPgHzZ0nIHDBVr
KHQ9z0mKtV4LFHf0hafzh99cTk5kV8EK1S3CGHZQJkJzdmccdonj5gzvhp3vZgb2NsrxyFi3QvnA
6OGd6i2toxH86TD0J+Ax0dyjqoQaDk9qBIc+9ECKg5oYSl3UOjKhLUA1qoA/x3A+Y4pWsO1Q9MSC
G7/GrLWyohcRQgaDS0P17RYRE7hRL4wii9wwAwwsjNahd5uaxd0ofkm+Pr/gnnGg/Vfp7uzrUt4k
uueO2ng5DkuPwTJH0usSqEcyrn7eI04fluV9BA8mxIVNJfYfTy2XB3abNO8WiCncdghtn0BmxMea
ljUTGQFhEppcTi6t8dfT8XXI9fw82TSCPuxOatxH2YUECykwJJbJ9V57cK0senKfh5qBFKfnSDcQ
rn/8Y6DzT+vJTgHh4GAA92tzVGpqQ6SIfH5W0Evi1mv8r/bxlXkAnumBGfwF+MrmEnP9NpREAopd
8L4OkKr4y1t5rvAOGG4X8EboEzfB6httSu53ob57eKqrJpOC0CZ4TfW5qGyGO/NibHP4+EX+djao
sT0d6wNCHpYvZx7IeP2wwwYsWuZb2bHLD4N8x9aYeVazNJlZIYi/DhSQbFJ8a6vdcL1uk0C6xruy
T+zG/dYSuEPRQaH+MRAwaqEKH0EaHeYGmZQ3SZNhtlK9KMhjTlrXW08Y6pgdFiOvDMtRTSe++U9i
7EYuHS8AMmfkLGkR8yvFQ4FixAa6brlYyITqYFQRuB6ieBU88fn5alh3F2+14D1KZy7AJ5wrzpCt
oG9WHWUswkdgbtJxzWydLf4jDs42/IaxuAF/zbg40ODAuJvLlBTDsRwujcBTdgczXRLIa6qeRRq5
aroeDwJLVSm78B7MB/lUfbaPN5yLtNFNVTSzqrkFa+6/NTF8s13YXseOKGhLdE3ROOKp9iC1pVqJ
5x31ZH1FoWbAwefXcbTYmg4vonZKyA5w/ppeg6FP72J8DABjprUzGHobCQnSfSGenKecDKCoOPBf
R+h1JMp5q57k9JX+Xtbl40jGXfXx4CBX4J97RLZ337jlCUtbEgc35/Sq4xwWDgFCmU1qioIJh+DX
1MRl0i7CtoI6iyrWpljZpFDN59OQHkgidHEfkWR7BqNE7g+ChLMK9ofEtkk8ndlXlEabh1Gnwin2
lidMxZzRWI1I2cyG4UB9AoK1zd3wfWlwqiuh05OMiXdVSJo56hF3yXe19miP+fDDx9CdjKrjmKau
LZ/B5sr2NckRC62WWmT0RcfaYEqxBi0OiDu33iA+cHEIecageba+rHHzadT/tyvwWYLyglNb3j+a
V3tGuatvbOBAF4ugfxjVwQYsSW0QYy11U7M/pCX2q84xPp+QgF2NKqejtmNhVUkiZ2zeVM2QDLJA
1uF2V+iYBBm/7Ds4OEK/LcMCrp57NY/u9xteeeH5nG81jfbVXvTmFleXQYOljYg6KtzU6ML08wvy
F0EvO8mPb7FBFh565++jDvvhYiC8HbwqIfcvYpjcJZw6v+su6CFTuFGOooLVWmfB+db26BMTX0l2
4Qnsa1Ac8IG3Vs8wEp0LEP4AzFvXJGCt9y+bW+fh9AJkP3FJtM3MMzrcHnsHWq7MJoR6iwW3MiES
VAixd4AOBmBCScmz0X/hekO/1AyIx/0ZyXqBEPpfD4zkVCGxWXkH6+OGY7zG9/DS25gQECsqGEI0
NnpOt3XsqmK3NGD4k3BR31wZEWBon7KOsz60gS+Ic/S8EXmMEenw3lMEkvsm5lBBro1rX5CGABCg
6POBCI52YDy2Ezvcc5C0hYawfoYLuyrJN7qkQ/K+SEdmvwITuLVxxxv2QqkP0yaomC2miOM1Dlf3
mj4sPoiVtXLrgoJlLYBK7QgkHym84CyKnYforhKx5KQv7k8ZmZa2qO0Zztf8go5TGw25jortzu3b
O+2wRmRwz1mOSCX7yMAVqvzEagNNu3ZO/c3dwsj9wn8SymoWa+e6fRGjJiWEAbMl2m3rCBaEjBiA
xQ2JEyfWCoU2whKSFdX52NuyidNFSKtryg1kpqL2ZRVC9ODGAa72ygYTJ4PfWbK4Zy0IOx/URJCO
D6FCNrPGzbyELD9k1Jls7qbe69aECBKILSiKXi0boK/nmh9PXJ/kyafNJ6NbT+7f7ZbpqamEUk2y
ASYnRCXTS7cegW+5rXTA+D7fHX1HeXrV7cvf65aGrXZfL1B4ldzqshpsOswTgtbqjwkzDn8UOmcf
CEa0crZ9yu21/eofMTMQzzqy22YQg4Jhhwnmxp+PqHUzE8M58b7DseBYgrTXCQSuEMiPZmbs3b0b
UxQCqYLmVt/bK0GSBWEn1xxKJvWba30bEZQ8CKD2l5AzdtPZNdN05Rnq/gKe9xOlJY1FaL24LR+H
Zja4DI9HNa8MoUc96E1lFWt9q+02ZGknvAGzBDsu4SQBzhvKDTo3ej9OTP4UVGUJ+aSe92gfoqhL
cHXkBRhdm5xFfHcmJMQkwJM+Ube319TsrHiQ/cu5XTgzN7jWIZoVLL3E2dZKkA8TTuMPzc14SaOY
Ve2OcR+z/DIhE/HCx3VbGATeXbtQwmZgR437rvOrKXGRv5hhZzB9Uwoxd5d1m21qJqWHKJUVs9SX
Q3lFQxNbl3alQTdTKnF6zXu96dR8/gakj12Lw6QX/IVttTehTP0AykNkiVUJbpqImyjSFD0H6AAU
3s4xowvzcvwuro4N8CnqcpguvZBL8+LjXTRzguzkkQhcSLjKXiul1DyZK1csZMMBP3cmu+7rblBa
0doXK01DqF4wN8CyO62Yfet1SBYWTw22ziMgtWruUs0D6BUQvSoWAppoFLRrdyf9w1dD4MFWzGfw
nkekHXWpuP7LeH8VAdlxlmiSKGeVipkmeT+ktfjT5VHuCUZlOmWaGnbBTP4VeTybJ+PM01HvP43t
37qRhooRmYxDJ+oNV1fZJiemM7fxqtK/yJcV+C6tZZkUfNZ5UZqHo1YNkfr2S0w4SwQArB6erMfd
PD4mOopFkV8+L0h/oe5yO9AHtfSby79ZAfbYtPpOFrqKyx53e31RnJy6Hgatxb48a0f3KzRoJZNN
wWzAcwBZ1VVOnM6BGBWg1ULVSCOsS9tSC6i0HKcZMexG9FP58u+fMe4H0OFfm0Yb8Cu6Dmjvusei
hqafHt46PlAYVUYhbCFRrrMPmi7j0yR51I0doWgvY3hbjKjYenlqa9qK7of7ehIg45gjB+oo1WhP
Fvi2W636qYv2N4pZJzn/iRt5PffjYUMI6DqYXrKMd9kUxqYkpJyIXggQxaeGR5dd5j4LYyMdI19y
rFnvyUAgpn4Ixoekqn2Vnq58oBmU6B+6IFthccwUMZwTNR12h2duVtwdrI7JpEOvkx5OJgDWE53j
VUIvX778k8KCl1Al7J5gAgXomFYDo+oTU3sWlg2801d2ygH0dORtaQbV9NDpxMlU/5TuHZkdry+K
cOINi5LG4kfjYzndGr/PfWEua4qC79+YJ6c9oX4DLjuah8U4bE+VcJFZLM/Gh10jgo4hQVu6tI+T
lIVF5iiMI9LCELdJZBfrEjzCPAfLUso0KiK9p1b4687wV168YZNaErdctJZHMTteoNUQ9gveZ9Qy
y2TVzzbLqRwnhqqswSr+TfLyYLnxw1BX7VjY6L0H1IHqOQn0YSNsUzTdZGtWTrmAL/BrsPpya2zs
+a3nXZtTmgdqVycvL2ddHDXwi/mWP5cIZ2SAAScCxwXpnp2UneDXduffTfzgVpGwdlQM/V+gYxHm
lkwLKsfQCVlN3FD8/psAbkRZ1yRR/Ewy9Fg41JM6cCI9f7jofzr6USRY8qtiCIrJ6vbOGF6kY2nw
7Y1BZnHmQ3FTw5srm7I1wMVpeCArUTFqeIrimoTQgEIv0iFpj/zTFrSsdAFDvxHTxXz6nycgBnMK
YK89iWnnTikFJJ3oL3j2tEFtHK9l8zBB7+kNRc0hw5EO5qrf7bxkQo8YFcTp7WITC9kFaL8vMwEp
OgOW+utgbgB4qGfJqhvoSvpE/7wjSeDFucOl4r1ZweeaItP9PCzODkLG1eIYsKG/zWRP32pU3vlg
5nwPULLhXLEkO4fyr+rLKq+XipHDzwT+91T/f3Cycw1I8948o6NfQn2rwuh3aJx0l/e7qTwpcwZR
Hf52GhnOr0VjJ1u8kdsU5E/C9taAawQ8HyqSfz/FLYd6MkMu/pXaQy98/P/BjrJA0HskNQSVpRqF
q18E+7FDZvqqi2YC8a9EvHIylghURwqOH24m9QFV+gYEY3NkoniQV6yi0WaUfwMwEesB3CDOKF+/
CRljHdRki8zNBuWxNlGvIIxPc0RbnzlQlUJ2DEED9QtbGo94T3LcnZ8zn6nkEku81v05povi1eAd
SjvzQw2Nswv6ctfBNovhHR7naNybAse506KT/sqdhNAT7+tjX2JO+1sy/c0fEAu13K1Ih6lQBu9w
SSY+fJM13AN3MJxsI5URrRHF8kYJZ8gCEaRQQ6z4+jA1DfYJnbHWtGP1r7vIpntXtzm3ISniGBoo
Jo1X2PNnz2cGGEhN6zyovtx1gJqCzVC1FrgKQ4/z9UJDv9WtUDS/fUYmuVCZaLuF+kpOEXTSWfh+
wyxuTjleozm1KR9PSnDdj3AzEkSMOSyWDmBhAi9sMTo0ZAl1iGfMlhP5BaAjJ5jY5iqzW8JR2zQy
C7efpsas+BPyEA4Ac5PDDvb54/t/3eTslN9Gvi85JsMwuuW52vCHxtEi5042kQShOuIxeqtc6lvl
hcFknOTA0VAFCFvVS3ZRNu/uMZlfxh9fZswp78IFAq/eSWoSsF48k5cDsMyeJWRGNFYbnbsEsMRz
HPR0RDTby4pl/G33/mvm9DFfqDGMQjvYRblS/4MGuGD2bGwxhlkMR2VBGr+h3j5Gq6+9p14v/Ftj
pJ9DJcPZLi/+43PayexKNFTLSZ0X2okKmLfS9Ut/RRbQUyVLY1lmwNEyTeu7sDXrdemwtoSz4+YT
YSW3H8AaW0vpTomoFIhVrm84itN+wFf/3iDI5L0a0cnX/RscwOweUhifsRafCZOM1wq1pouTCVfS
ymxYYB84Fcix4oCcxSwC2BJVftGG2tXm1y8cWlB+nAhHiSU5ApeEzRVE84hihTmfrXRQjId2dd2R
tvKOUMNvGv+QXN1SAYqpKL7EF1AY+RhrMA8qzhzhK13MBSvBEXqAkxw3xf6Bc8GLvTNuude7/BHM
6W4OAsZVsSKlvaRdFyuZKwqnuGiBxOUvrd1RMqTOGCoKDY1rihv6zLkeqFUl2OneEgSIYTpjQTBH
uyogJ6z3DvAdMewtFWpxHGTmZvPPcvPEjqytUoAmoP2AvSiUc3rOEaJFQEB21Cgpi82SuYf+fE1l
vjUR9Ge9O9rwzUvn23eDr0Wex3J97lwCyYIdvI1xR+YWcBMyMzr13ftuvOkjnbvEnMyv0+b6kU/G
bInxOv3pXS7nPOQbiB9RCkuQ1ekFfOekQ0n0XUAb7VIyIZvafFkUVqcVsiTaHaWDvi8BUdlRsCgz
Bm2UDX58JXkMMfqPpPRehOKAeLi8qjQQKK3fcVX3TWcWzdbR7nj/d5Jq/GLhbZ80HjjwzVekTgk4
qc+/qZ0awgiyREt1kLZrrJUe4VvljFWYzLjMmn38B4VL32XzLkq7mY6DWZJYflkD3Ja2COgGu1DW
UVPepbC11NcQntwLjMUZosv014YrM75MX+8N0dAQBjsfwHU1DUpHvS8f+hTBgM0QNKIjQzllRgEH
HgTMjAfMi4Auqq3HFTM/z2H2PKVK8DIS8MqS4e3e0wmjKdGM8UdS0PEQvoScVYLmjcGZmZXGrjxy
kc4GzEXF1HJi6mQg4HiBkJy6d7FCJn5OgAgoCZSove0SluE3EejYylMf6mZnCRkCR2j5pc015aU1
lAdVO4dzRlL+hZ+y1sCrSybUYSfxW2qNe0Knt77XLl7u7gpxkkgJq1XbUPqjrOcZPhav/5fMSAnF
UnwHmzG0ALuVKT6GxOZ3cCHuzdNvcMbKXkWr3cjJoJ47urliLrji2fJMxh0JCa6UWgN9HMIbGHZa
64rDKjpOp8m+uxi1abm48RV5QrtY1tLV78iPmVA9V3IiYLrTZKccID/iLJXJARDH/jZ0U1Qbx9uB
PTQYKpIysoeHNjMxKqW+yXEgwvUSClynGHFyefE1t/UCXeMvzUX29hsV6AYEsBt5QF9ELisPBVTT
4KOS88kY4C6Gx9/ks/mW6V6mkhW7paZcFIwYdslLkPUHbjNf581tbcuDSNSKceHlqw2pwDaRwQG7
PFA4u9vteIaKIU8sW2fqyY6G3G+ziIZp1tRWZ7z1aiOinXl5aisPBnzuIA0xr87PCnrCW/872Ou4
sDQ326eBdaJqgPtdpTaRr8Np7TWaerL3DyB2rOLgDcSUypVsaMUG1o+GNDNSjfkcvqmbRsJHJmuK
OgGMoWOfobko1xQ5eYUXQYGt3YaRPJ5GGQLrkEvLI8lWeDI6DHWIrVOg40caGHodXClbgFJbA2Ps
BL8oeIJ+D8fm7UosPsWq8MPENC64FxBuPmmPRUDbyIzt0w9rvrLhI7fgPUSfpt8odwFC8Qq1n8Qa
b+k5/uHLo9chYxwPmqtgqpY07DT20VoL9SejDgDSrPnE9SJEOYfIHvs//VI/s/KRGjrO4ZBa/dmS
dUBLCQEhJkKuIoa1AOuRklLL0GMpqyeREkgcFeXMDBzVrgvtjc6WQoIfAQChDU+p0UZ7cl/Cj0wf
Rx6x0vIgV2DbhkvLE5EGAybaWvorAefUv1z1b43R/wnxxD/f0NVEgsKlt3xHaIoBnfS/r9SnlNA5
r6j/nGX18N6vpzVdY9u7TRLjydpZfbPLWtytMNMvnugEUEcyqpM02G9J+fzxDAblgRnhmX/OXMso
fs3UcGN0AYNWU4Pwul2x0OC/dIGY40ZxhQYnKbB7qoDghdHo44o5vw40Ab6C81SLf53fZBZGOG6h
b2REwkh9LGud5ssiuKhqRapKrxjTOgMiKGvymrNeIms7g9olHs6Hkh4rjEwTEzBhqDLpInBjLWdg
4XJ4qv9OEZBA22lBfoW/cqMrkl/5wfESpFBhswfngvQtE2BkFiEVPhTam+0ZaBj3dkY2zPZkiGsK
MzR1KPM/fVfxPFFqEbeSO+bsUKuCJcFwOtqlKvSydoOQGxsKwEfrKs/sv+kUs4gc9J/Xqbf5Hcnd
WnybLKlwovzf1vlpS9XuyEZLRK80HCr7Y8bYu0Ls1Uq64GXZ59nVZFF9VbVVqIf22vG8bAhi/tlr
Px3bQORV1BLKFsEZ9Op+4CnAOAqLP6ZVys8ayeMPUDICRYs4Yz4w5p9MlhHD5jci3UNJTNcoeUlL
9l8xhlSpP3U1QiM7DfLOqewtbOZCT0cbmBv39CjbDwh04NZ9qwy8mEVlyMW/t6szp7eH09DAv0BO
hsfa58GYNZPNotDGWFD4k+xyC7O7FAHsehW8mkbPw9kbHtJHuzkNYR7QNzVGZH1ttI3TKLGZpRK9
/NarMhAJeFs107XR/cTj5wsrKkoCpmYLT8ijmqv6wXGoS8d+u3oXEFgFS1lOYmNg0Fm+STayysgP
FnFQz9SrgpSPvMvR5iTuLKtOc5fPByVsXoglhYjn7qYrAJomvK1QaaUKoc4v5ToHpxEQE/ObVLg+
Q+/WBiFIK4X37osnMwyJ/84ZAuf35+gQyMgDLlAiocGL1eGu0/LBrBL6sFt1fKUZnDZL3CRTkiV/
qrn2vWy5dQlqyjGIC1wicsNrmpJIMevKnhq9zoSJCp8Q+rhRBSp4HCjgtMlWYrlJnQF+whORGL1R
Lio3BmADFcP+sTgxxmrexa0rBIyOthVVEqr01C/bIYbqrFdRfPGGuj3jZ0Sw4f4BwhEUjKGLBtIg
67ZAsb/Xs5Bt52Ucd6q+X9VSlMwM85SoPeen4Gx1TfjRngWupCFS6Odh7GTL+bnGJVZ4/w0W64Lz
l7fqUpgRaNdJEahl3Y4+j6EFy7d5ih8PLoWEJ13vo0lLualDqUa8ayJ2yHeIkTk4dQtuPdTf+Zko
akvsOtt9JTMKWyAU6Y1vIqimTeLvDbu6YtHTQ4vidklAM1FnRj3gop90HKkczn4sHmpAxU58Y6Vo
7KcBhUb49e2TNPUpmVVib2e9KG1AWY3kjwtvbwwjBqe9F0/E8P46GbESYZWxm6+UuWQD3mr2BTNq
n3n1l8gcF+ey7jY+9nzrtEIO+FldU2HM1KOTbRTA8QE12JTCTdrRKR0Jqn9NAy0r+katRYIpNxNB
Xe7LkeKdFW8N1p+UvntledE4WqpaCi7MfrvRTKOdUpWr+cgwfk5VWD3CzmCv43h9I5eJy9NWGtZ1
SIVkxHIUHjee0l8rDxCoxrKX/Re0Xlgz5cYWGOquFdLM8pFxbc5sppOLJaeSTCfV+dlF5aURZGt4
XTgMMBBcT6xqO/WJ+15k0g2tazby/QmGKmBBVGhLVHbqlMWniTQLe6g8C4j7p0CA+LbAI0GxTna9
FRhvUOt2X0odebxmRtH3+Hs/jsmloMigJeBvrtYLfL0+UXyOnUawPTAovJZ0rsVvkNWOj/o7g50U
aKU5l2vOcj08vK5nNEGvx/QXY63FqaVdjP34gjCAHgDWetOjRDUFM+Z15ICdJkhrb0QaQS++9E6v
CcHDlruONvzFrUgZ4VGjP31en6kqD3VY0kHoN6NpqVEFD70xAHhXDKhoBs7O3gb33+wMlM3oSKsC
VLCYvpuWObJNBGm5PQOjqmrb6804oXvrsRN++wvpJHdsYkw0e/v9Wh8GMjPN84sKetF6y+dtbsjP
d3FSFb8pwaSw97u/8HOa4pE+E5EQrH03yImXPzEn42yGyY7eRBUiF2NqS2lLlIzNGv8bG5uXoiTi
0pF9pkNTQr9Cq+X8WtvnSTtDME0W9XGiU1WW1y+lkwWYyV4bYrVnooknIipXQYQNTz99LM+QPTCo
PwZhCJdhJC35NClm6CSWFH60duIF7VAsaas0yfNuxMp3BpdI5qVD1IUVFVZI2Y7YITXnbIrwffow
PTzSn0zLtkltRwBwzh2yUvvgU8eOwtb+qiw27zYCXD2PlnexD3DMUIdA4Crj+QoXPnF8Lkw+Rwuu
bygiIo2SfcxTOEn5r0G5NpMHP7gb9p/hhd62XZJ7nBlyEJADo+c1xvEsGdcBcqumRKcl10vxhJ3d
FVN5yB3juzuo4/yuh5eazMRl71lPflF2cdBZv27cjuYeUHLRreQBvcma0ult5sKn8p2WMbG28KVT
/pbYJ9i6nX5fBO1GspsZG9xMQM5md4worbw8qPhTbpf0EAC6LlW0aZHPEbrjEinZ8B3z6/GT0HXp
bqf+RoNo3tyTgWrW3BgLTcDjG6F0NAae3+Ml/JDr0Rn1Nq/F2yyIbqW6iWgm7yOVHy8U5tE+jrMM
9nQS/ZFG5iAWVhHRxkGF4to/P+mtxe/+X8U6Mu/q+BhdeEU5WyXKNoPPeqwcKeXxWYYD0OTKLaLy
q49Zx1RKJqFjbQY3XV9btlOau5u+oLpL+iw2SymluWztaFHbOTWueDZ3j7nzzjtF7CTlLBHNHYdc
5YUizTCgEXwqgi5oCkkd/aOfhUdJp53nYb40y7G5otmJIFiybqpRlivSIF2Ij3wFeS65/h9Ot0dW
uSyyz+JBYqmFiRe48xUTMUeCJgXv0NFl7+6GKvecFsEAxVERCzj11LUlTg1kH4BHSYk2w33Sa27S
GEa6dTXVdk7xhZDEZMNqs2MvnZYuIwzjhlCpXQ7utX8jke/jy9FrVQWtG7Ts1taO23P4IKrVaRMj
3XMYVlexsn+9RQhbnaz9vCG8fML7u2DlJN37wNvTUU9Oo+hYZBD3e4xhLz9Z4F9sS6XahGx9BVvp
5XNXHNlTlrhvb8MkzZWJcPDWxCcOpNPhjMl3nHou03mmiIKO43x/bAUZHmv9OK4dI5qvl2jfic0k
vKx/QEE26vdK6YIxWy2mFMvW5HJcQSE3JU18zM9tXZg/nFFGRfMBUn/X2EfvIlU+R3n6czuftc6J
WPmHC0M1rERo1YP8L7tcrobSO+6SF1373yvGquAWzlzKOmkyWkPAGYQGchYEtjq+UO0OwxB3uclj
0ReJM06eTWObYFXhuMZ3Gc7l4tTfhf+DlPePcLCtrJKzW/22iS63WuHnW4snQ7BDg0Vnoz6wM0tD
SyFIAeLF+DwACP9Ir4ALG6+c4eZMETUGRJJu7NzUYkxW9c1RhJH1s9Tkd75FTwQ7ZZ9FUYpTmK/N
ABeR5BS3I9NR4Y6WWwN0R4Yniz5rO1VIZ8iDTdiKM0qAwrWlJHbZPoz+ejmAILSfm4araekgqGQj
SJtDaFxNpsP+9EGO7ZLkV/yOvaEvLv4s4/EtY2mG8OyCW3ZyyQLHfbLXY2vPgoSV3Ecs92J5CjlK
tFPdLZzGax9YA2lPX5UxEDojtMug1epgRWEajdahtvsItHXHeUaIqw5xoy7vmBAdtygU5wkwh5L+
+TvFmXif4MLdomZbR1KtVThr9ZBf44xBWE60YxjmMxciq+lxRZqwigdq6Jv0itFngxsXgwkRxXZZ
VWjyoeSek/rXueZI6Rok32yqQ9DL95v6jlo7SC5dE4YzlX+ffyHRLNJlIWmV4RsCMveJByz3M1q1
uY0Cebrt+tWYJvhBsDmo+K2Pw3fBeIxhcbPPUo5v36FncuuThwCiCCyE0FZcltrOiC+AviF/8ZUE
q8L01ENqO9SNMwKJBHXNO2jqP/cRoHx5cdOm2dtwjCaCKqjOOI097PAqDpRTQXFgIrfc16YeqQ9T
vOCcUKqzrPa2nm/olf0t7Ulm8FKWHqouDzEZSIIGBusHIfr1BV8MenYI3g+g10a9MlVKQay/HDG6
taDIwR5yXvbCMJGzyZFCKEGz61EpZJmazeWlYqliRqccboIBkXlbjk3Nzufr4x1mS+Oyf1FatlMz
wOmWQK7kDVxZhIIU4G26ERwxF4Lt1tqhBAiYUDCTH+6lHqbiZEtDSnWxWudy2GeMVQ5l2f++qSG4
SQ9EueBwMUthCAZfMDoGO93hzsEMVi4Bce80EBgYnKIx7+VmqLhy9G/rKNqQoy8mx9JoHPEY7lXf
pN2vP5Tdydkc4JspNtHIL1rEkbnUhW/pC8wHJgcVMVFWthK6Kw/clLkQ6YXH7IqtslndwT0t1N7m
sRVo5cHwXkCFI0cB6Hiqjll+rPrkGN5T8ZlkgA+89GjiUv7lqedijhT4MIwMAxSLaYBBPPFPfDz7
U7LdefYwKQcTg2fFAKLMU+Za/Dt2enlAb4l1NFfw6hBglF4sPv2qK/+aIr8mr43L+gNgX5r/pVhQ
Sbwr3HGNogOD6Il3Zoso0SmT5wtKsPnNXGN8RTqykIQexo90BMBengNTbYkNjGuZMhw1fP7b+rvU
CXyMRPpmfcK9iG131PlFfohFQ5URpndg4FYIc0Fsd959f0AE+nWBZyu+YhPn19vAY63mwJUHKPOQ
a9fFspaNUdiAHCgs78W7+2bQVR18irNf6NtqBVg7Mu42R2OLwurKIHjdI73d3Y6JXc3uNLsHipo9
ILHtJCWEpvtEgiOQOYFYzpfgNv2wA58tTnNMRxOaueRBrRys2UCo1vQVUzPCgWt691UALJFZ72vK
xEdBXYXdb21ua8Nw+WeqqG3q5azqU2qTcmI6hd9fn+6uGi0vPZPGeQRP3UOvyM4+bu4vC4PXEQDk
xbYrFraO9AhgVD0LnOKFzTjJkRTGidTL6sA/98XsuKLNUI1GRaoFUznEjtP48FUL8+8mlNoosjdA
Xlnr3RhfB4euL+0AEYNUJm6g+aS3vxKAEIFJNgXaQA5qfB+Cdvw/xO3qgOQxvIkPTZaZD0kzBJ1P
8lV1LkGyW4vjL3Z2DG8LOvAczsIaGd5H+6uVr6Ns+k9xjVCMt6bDixAumB99o/ySq8DA96CRbovh
/v7s0SXGqI7q8Bu630BjQ3P5Zs4UZnnK95zjRdf98OsjYco8132Cf6gTgelZdTVSJNqRaRvAiwwo
1eUb2CXtHUFn222fYUR9PftDfsFk3Ghq4hHc+jFek+0ylsPE65e5H/A1cmHGI9EZr8wkTye2Cowt
1E/Q3T/5SkpETYQTR1t8CQQOBwlO2Xqx222cQBoCr51Ie0TKslLzpproFWLvjhS0KthgrNoyYJ6/
il4Jp+Mu8y7ZNKKYedByOu/Uq/ErScQKmrjWz+U/ReGpWlJkd7i8iCDt1pe1SGCiti36+Ib3BcFu
H0MlWEKpmqoihp4gmgup6pWn7rZ2+WFMvAGEN4OVYHrLWGAYsN2wmWHZd9eFRvY/vLDputF5TCfH
nlFW+5k2A7n49sAK7wkheDaQZlWsr6vtPXaZO6AM/u8+2/laUJNMqDadtAjE+PfHf+nI33yJCvaw
i+DGOqtOwJGfni0jaXl2i1aGZCRXsCu7WUNqSTf3CiTnEDZZp/ghyNrKPqgSDDeiwFcLYhPXzlvy
jM8heJ7OFkP5M3rZNNPalBnSMU95Uzv21sB2QHDJLDy9aT8sDnB7Dfa6tkps7majhhasCux+CuMn
J4nY+Ak3daRk/JhpAlSfPureA/ZubbuoalMUnmlmmg9k85MnGxnhKgUsCdA5kufbmjWVzJkE5P3p
A3C4+UnBHzyi3Ffe7f8VULUnrWIkMk5VEMez172pIA5DzTd+4UauGjU9VJFKnT52nhGQFYu2M1j2
zGU8YuXNdocVbCaaEDMOKIVfQl529XqN7UAR4E+f7FKCpIvVEmIzDrtHTTgWGfO3RaPQK9ki+Qx5
wWqTiEaqNQ8BuOyMaSGqI+uv++Jl3mpSLbWXcjG/JllzEQPRxYQztBpow26RFaG7P/Crn/rI58kF
OVTwRbTcBVYR5CBOHShmOrMz5YY6FGWpEyfL2+AQJGyak6082SnWB6oJJJ0z35pNWyvsarBt+XdK
1R0fwJqxDB4WFtiYjtEhzS0f35vCfXL69Lu7UdEVE6f839tO+cPxC45E7HM3SVd/T7RgmeyGspJP
HnmuPqc3/2c2FclEY34x2cYUC/rK0lsilxu0uSyOVi23gwqIpSApL1Amr7Qi/mOIHj00xsbFtm5F
Q6kPCBdWTNfTuZ1H88LvEMFAMAorp4HdzCaQxDZ/49Bn5/DJu+KVmxRM+gvXjGXXIC/BBgnTFme+
x6/zzdogmJisr2FocqcjrivruXvp0DiPtSwlr1YIaqPGggxH1hMVgcgkZbNE0ne4RlYQF9qwxQRw
Qp+RUsNnX59VB03aD/OzHvz98wEub8ctQMXklDwKBpiwnWP7HvDgGpBxA6XGkj/O6NhzVUTzZPam
LaPCFhCaI5h2XKP4H58MQCGzH4D8/YjBE7OtIZLLNgoTwKbrTASgeQzSb4To20wP4F/eKr4VatQw
0vpAVcrH/nGhGdFZNdhQbeDEsVaUJtBged0no5N0wgDqE9cjPD0YnjMllo9Qlkmum+TVToPkLS1R
eIqXJ5W2EGC6Vkzb8MOmtAC9WtwNmBOpcGn1slC830KmFbv/QDiuvM5d1WHWYaLsmK1W6aG2mPjH
EeUQKtJOjAiuzABvibox6+LdnPl373iWLijFvMeh3PN6D/7sFi6L9R9D4OAfP1iJdpWeLZxiU8T4
Lnw/Ytie2l6mEMbkPVOyfxKTyg1gTe16nEutnTifZb8jleAW6iIQUgUXFKWXggRfdv5jf/xJM2P8
3fZMV8vMo2O0Ni8EJfHqxuAEi0SnuEkiyPjm39DrhE4NrkgruntAayQdGhwcVEo5tgSwx+iUkTkc
BMCCozA7Tcr343WMbT4tg7W19IplCRqWdBFKGwFnkFsxGv4GGZS83vMs3lRC8jnnjHGK5XzS0blg
vutX67/jVWtagBjtw5rVdB/NxTbxKR4h5fdIWdfHG8VD0j/EgSATpYv4H9Ej8Ux5u2jRyts7HUDT
n3KMgtf48pltdBsubWDMqLWNaE+krcPtZMVwxz051CH1LEoMMxj0Q9kTdMFYHXn1mIrf+SLr+QNB
oIh0P3cRWZWwVR50En6YCEBtZ1p56fpjTwhC+8Fl2Dtw1v3y6kMJijk2hNyAZ/0NOMpby5YwoTdH
gqhpNsnStQR5ibVHjE4rWlils+ayzOtWiaXU9fGYa/Z61W+MNGuqq2OdBV/mNxNmtcK7DQO8tr3t
zgeTKp154l2J7ceK933GJShipJt9F7ZAbHQntVPH4maHGIolQHuzFrnUfsCnU6MU9DTbrg2GTgSV
TYMw8yU07r6QZ/YynTQ9+IpSXn49jXRa91YYMI74FU6u/9DSMnKne/sn0Wo/26TF8wxxV5dgKMwP
2aOCRTHMhqC6who4bTjecBGh4W9OjlvL3fELbnNeuFsjhSqW427ScqVGA3Cdq5DxkNKQ3UR1rIRj
88bpypRK/jZ7aZvcn1DC9oVhyh/Yn1zuT/INsVTB/xqFDSqZU/HL2aOaC7JPg24Nj2xoeiWhPQYW
GO6IJApcvalUJZubGGwlKaY6ovTivOww/WN3aL5le9406DnixUTMLcwqptKje8IpC4IPxA0mE5AA
rVOGinT7/ezm4EsA+SZsxzAG4HxJ2FHP6IMs9309SzKQBm52drZUqOznm0IIfGzY6pW9dm5FPsOR
9jxdhczCTjCIYskfMY5obiON1N8aFHaJLUqL5w2JRLmVhodZy+NruwFZTLSxcP3O49qK9uc/JPdz
ZsJVwwWQrM7/RJoNhMxdxQXHI5YRWdgIYm6bVm11e8qxESul0jDuMc8A0nVblGw//nezs0fyyvap
Xba+8IbvqX502ACc/196Pof1s1yReTy54ISjUXwul3Wskqex2KUPNt7KVmFANVeDfwdMuVjN7H+a
cmaPYEuI0EN2oXZE9PxlBPFhxvzTLK/B+9YSsJqNPRhbwfDcmqCjwtkc/pIxRL2siW1tPmTqWjMg
cea0exUmIbyftfTvmFV2fahXv4CzaJHyY/llSb+bRx/NNsin02OXhbgObi/J69aJkrP/UxDpIWIe
qWJjVbXu4lKyJNNnY7rYK5bBHbMzRGVD1ZH57VVOu/u4Ib9VmhgsUvAhP93PvBS04d7J6QIUi2hj
etNIGbJzPcl1L9Rc6tlFZXqPah4BL9R2Exj0UH5kFzwnJFhdkA0KOs6so600s+yerF+SL1rbGQZd
K4ZMOCoXPkj80wkJYD993nZ9FRd2q77J+yAAMazM1u8YY2nZJKcIbqR23udkJprRt3gKmxdXYoxt
qvGy4jDDY8cPoSiFYPHKkNQOWQsB0xzA0Gmx/jrbGwP3znQjtYk9yYbcz1f03cnoBwVbTAmXk+af
vO0x/TrRixeAQODbWbOH26H75F3flkc7Py/D4dCoc8+EVjcXLcVwJ6W9Ks+2pLSDv7DOeACKneP6
uUp4r1lTvq8CpCnPv7bnrZzEbxHzR+/UxweoGPXxA2zHA0/DOl5+WLmtuIN051vudD1RVxh9n2QB
/74ljQEGWhLbm8Ds5KLmvLpuff9nnpuSK0+w5NROl4ZvGnvJP79clJUiz9Y4MyPRRQw9JYUc7tKY
91w8+CE2+AfNU6Qp/nMYXr+fNl5RK09AOb3pMpB+W+uRx5ndtBIqKMmNfxwj5zYNYR/NIuL7tlr7
XUBb9S7EvogepH9deQPm4Am3Q4LVFLm+b7DeXhPJs0bc8SmiWtxLHfE8dPfGzWAXSj3ScfT0N7m3
RlzR3L5lVufN/deYBcakKvKxNAHjp2sajQiT8MgrNciqSW9F3boip9sXIwrxnUPb1NN5jDKWBc/z
yr2s7XRTtZZs5v5k3txp3TzCRKR9emYQG7mFZIbSnVrrNiV4T8/bQ9rw8G83kZNxDpi0cELIFebf
Z1B3KJPFodm6HXqylSGu+pT/bzWE+vT93NvEi11DJb9Uia1o+Bt0n88BDbZFYMdqs6lI8fvwzyU/
WY9AYvoN0tbu2/+eQVeumgCpFRYpWXy5QVAXcUnhHnm2m2DyHDZ1YQQ2Nlk9LfXeMo1S58kdSQCm
hZuSPhM6/kmF29i9IShRxklZ/uglud6NdCQWHz/VF77WiJwcy5xIEOQ2mqQkEvuUrlAG9l+sxeEb
6kt4qgBCtvng9UIEO5tDm5LtVf0evQf2db2txt6cSrn4L6RBEQM2pSwuBSwQTOsW+fA6AlnTqVDO
O5HM6+kV+NC7GbV+W/JN9fxdyVIF2wqYCw8NfqVLskL+sbfaqYDktstRyAPiwEs4kIpZkXiacNjK
x9Fa27LeB5/tBe+B+G5+qWgF7eQ95gH7Oy5iTN35b/OtWKKXTjBT9fOYEFTO6gezoK4vjDpfhtwN
/T7deaUCT6BO4fnw1IoXgpkjfueTIHMlkCLWKuYOfhzsY9M9hJq3bs5+Ri8JESE/klW/fUWgqGKE
Ok0xIWFTNozOQ/6ZOEipnCNxqblqn60nRnSAh95cYNkNVsO4cTnDEu08KXId064cSnmFPOqDtddS
EHHim+wUFgE44TkZ897A84RaYDR/8QLKzB0OO1h83N7sC1gq6/cK9JZxUjmbGy1zCeLQch2WPl21
pesnrREemN+pxVAFFYhhkYssGA4SYw/DmXKcbD+nlxhJ78072Q7UYJF2jWZLOAKkd+1iUU5ffQEk
keLKtTPFmTe9dbMyOPSwSDL1kWQNWPUnuCtd45omotJpCmyQnflbsBzR3Mb5qF8ayex4iPjM1qaG
JeeXeTTmMYuuLU5gjs2SxH3bWWpN84s3NTo+raRUlG3aI2sQ4SpJK858AE5AMAt7moREd+uFWtAc
Efp731I+35P2+i0VaXqgg4yFqz8UJlLrF+2B3qmNw97I6lUWSotnydL3cjCDTmPPezOscMgukekz
f/7NGbhGuWxv/PhH3VtV0BIlWrUPNjCpBkDhmZX2jEuWlXoCxxauOn9PnbgQN++cKTZ5UX2S+xDe
NJgr7iCqN7JcVKtUAFticOWm/4WJyhFkZ1ebTcxSzMx+x3oewNw/HZq2OIGHMccMV8TZMfEyn60f
Wm3YQ0BUlOfdoxwTlxV28ijKSpoDX6Zb1bb9sRpbtoI7aXCGVbgmBvuq1+4xtZJ3W3s6DC4CHN/G
wHao9gGj0CMRbgmzRGlwenB1hvi0QEXlWP8TexpEMEyB8EOkHAVhhD3ln1Qd+hlMRb1JBa3HQXvc
/OLK0LXrEKc7+B+smRSWkfw37UNZ3zATHmhKQC1aIvPfmyKW5SFX3b/wNX98CHv8vtCSAZG9M2fv
/F5OUYXT6q0eIgzjD/5sv0vhmHaIdIoLb1/2LmhLBPVaYYsFMqQ3tNUanVhKMoe4t18srYy23OyN
yxW/ZN4kb46zL395X3IkAiYE/OLtlpXS2PdgZedIl2wLMJBuHSFv/jTeTZxPWuy0nuwgHD4A4Guo
AWUddKm4nK961uRm5wJ0iZnQ79ewQf71FFZOKTjrxSbPT7JQ7ikww9Za4E2hRsG/Zs16U+TvIsFp
Ko8ic44Zn5fGUYBP+2trJGddhl40aW4YLRt5g7HCw1f6r5TH0f3S7q4MBR3EFAthd3cjz83Rrl76
q/K94PAZjY3V5cnsSvT+n+0H03L3aD8N4QAip92uvNe8aSPi8kT/IutRbIqxI5oFTLJY1+5939kT
rjtc+d53HV0re1pc1+xZrOU62NocGBvngJMDwSP9Qyn72EOnMh0XUGNviSA3ubrsDwaVYTRSpM/r
tJ+PKCiTCygGprIvdzeAI2MfxkU+pJd1UwI2PkLCioEeVZHtSzzp3RSLmBOCmowFqVULNOZ4wTyw
k6xaCk5W29/aLBoGNLsue2m9swO1YZyDb48Y4eqEAvYO4+OI4t+k1b4GrxewfG6gS2vD5vqfAKDj
HDPjapYxFQuhzzblZ2H3dd9gZ507ax2SSZwviNN/f0KUJ/ebvbbs6dexEQ+ecn2Z9qBvM16Uc2kz
XZ0YZVm2KM+cN/NtVCwqEZJMdXZxpOR1YWdSETlAK9nsLip4En5gsspcurB8pAi3UVHJdtnbEGs4
vbV9RmHe5Oqd0a8v0+gJNJgZYYt02cOA77iWjL6ga0yfeZCPkJTf4QjUfb22DjWKjO5nL7Px2KXc
0zAhb1oxI2XWy/bOkMJshF/q4PjuEC4jiX549SM2xQXghJbcZ+0S1V7Aw+/Q7YpyFUxq/G5Af9el
ARhSGcCeZCUngVJYZStvsG+oSka0UtnJu+LhpgilVzxtRs7xKcHR/KaGPiSe6VLbp49m2te5z153
p6ElaHwFvgMrybm5gvu7cOsaD4AiGnCL5d0L7+Mvh6pI6jMJDScGUarIacmCVH8rwNYpf2LN1998
8duPaMWflvp8VN2FMOuK1mX7qYbJj6u8cmho1HL2JgyrPyeQTwq8A55DAGTTOuxZ0R6+Dmp6rwsV
DwRzqDXcB2yWXi3yxfrvHDqto+XfT2Fe7Es+IiW20JeEtZrF3DjfBxuHkukGFtxdTwjR4oaBvLub
7LV4LQ/kA+kUes6PK7afQIlwMSqJh3QcLT6l+Epv2V9JHjSwlGU3D22DWz2yZSPgRJDG6YS4kuoV
VudYGkA7UsfgoThkf+5/GmOHZtNwKIpJnEuxLDO3S+2kEdkWW6WFB0bGpdZsbFOhF+bXoSCpoOn2
eYgzlTMrwJgcKOcey+WMjs1QooCt2ucqCeHUPZOJeTw49a9jXg6KxXgmmNLTn3CEUKWR/yHdCK5X
VHHxhQuO6kJ82NJYEs6lzT3rAaZffRoQXfSigSvR1e6BdkmyVrCQ+xrk7jLIAfE/9lsVd0Sm7zRw
+t9gLjDzlzxorzVUTn25XFzm8XTcav6F7ksPgX20yldOkT8SP0Yl1sWtx9Ncl/GruZi3akopdEVi
RuE4xi788H1KGHxOuV/Ty5irCUiA4NuR0yREil+tXzKzaa3FO2T6WDpgj2Ok/kbZepFu3/RBF2Cp
IUG3YaAgBf9CrA7S354OaI7/ybGzo0BK2sgb9tLJ2Ax+RvybOTmfLn8MefpVZRi97cyvmqTwmyok
fGg2cK1zZan47VC6xUe5977JXDjKNhDd+XVMxogYZ4wQYqGA4QFV6Hva4qz6zr8HF5/wWLDE9VSU
l+42VmIzYxEDyEmGh3zeIqlgUCpRyNCJRc2ncAAJ5fA7O98X0Sna72t1fSFimE5GgiVrAO3qoti3
mERRebQFe2aciNsH+ff7tm2jYH3a2N9wCS/82dIuSPdftGHDlB7eASEgWRXlmpxSh9cNVJ67hnfO
2ZYn9qXZ96xWN6KJ/FaOHcVAP2DnPbgUCf8JclypF3ec9bEdY1usgkCHPZbd+GAne1VD2yICPdJI
UcJ9ECYJq1oiWLW134zJhJobs59AC/p2qzMM/NJo4Jtk2mYkoh2UpupTOoFOxFlxE/FjePZ4/uCp
iuH9N3ca1I482AZvab+nGF1p+GMmCD+EL34rEvFRpd58CbjuQSb5AlFV87VKP7XGWL6nEJplkkNb
S2QebhhO+JYvYq9PSrjqvfIFGl7m71E6cUtyX7W8ywQiP4ZIhqFtDGWOa9R6Fdk0MPeE3T7OIUbD
16vYZ7wed+ZbPx9YRlmf8l4176lr8zEbedd0XuapLp3xC10ovkUsTcMQ40i81cwXh/cjxU4vIwAW
aYp6cXB3lzundYxTS796RM00giaN2vfffZzfoGGeiN60a0w8OOFL71BNAbdk6NN+OwGHBVgoTWuG
IYOR0ORhTWQmJjWhHC2uOqPyhicO+bfdygUTPitjZ2b7cG6XpqlaI7xsDMepa/NQb/ilw6ARXpjd
b3IxCpjS3nVFXar4gcTikM/CSTIbWQhCbLqI8Sg9E35M4ULBEH7zi475ToT0Rnx4Nkp/9K6KicLo
fLcpq9jAdbr5Ro+h0kZsewmDvsn03n603NZj5zZdRw5t/mQBmqRHAAb7UDylxiBN8cpTwvAeO2Fg
cpMjsj8Ex5/t6nUzZg8eNmS5+irtZz+HPj6HqLKU/AlVWYl/7vKEbe+3TMqrcPW6BHPMGweo3mAT
loSyTU7Ik6jEFJR3PxxHGohDzxjAaGfLgsqfWvh6C/+Na7p5WzEXiYItEIPn97oNStLvL+EYSE+t
2Nw42E5D7oBLbQNV9oEfpIhuD2wHBtF2rkeyMqPf2TrR3Hbl+b/cbvLUTkt5Ow69DOYj7OK75xj2
xlPURSFCqSy9c/uzI7WWKfrxUIdtZt2ZRpmo3wF2CROTxUqsaSNF77oF3nEW2YzmZLcVaL+s10b5
CxCiEjYQkiD+yPidbiBsQp0j8fZ75gDSaEjoImcEgGmfna7V6jP1z+u7DzGMktiBtZDpSb8NkUtf
nRHAO7Ya9P33tcuwxtLy1R2KDuM8Kf9tWuk9LfDZl6A2uF1JRVBNLdn4n/gtHz4OMaz54ytdYBT2
RV7OLE8rYuDjeM6u1sDV6KABcjEZ3tGWsmmIk3stEGStqErSE17XrIy4yhc8BfKNzwMHA8m6dE8i
dsOkariQG0RAMMhc4wDjTe4c97uDZXlI6K8V+81VsE5+3Kq7WUPaGbOmRZa5Xgr9GDUijLyB6B+5
QtzXhn1RrNuBfPk4ftKKTFKDzPe+Q8LSIu2+lt+cppjCD5Ap0yebpg8ks13dzO67pbJ2FiIFzCWK
9pJZBoKF58n740uSUhrRcALxRXVK+ZdjhlFTk8/T32uLxDwUlsclVjCAmSq1+ra+hxUUVhLT6KGp
5IHvosLY1U/r+A4LSCsod2/Mdn690pUoOr6g5c2PlEePWH3x7+cAOBFrXbRjhv986CeO32rieijY
vRp8AR54DuX0urKE6LSxxukK+ZjjSZG3PF4vNLZm+JSoQV4kbewkvbCACuOntc7DUQbSbbhdx+uU
K/vaVSZAgO7NFE5upeotFx5u/pHaqy01wG8cnvDLGPf/VO3o7kRX4MzsBExAt6MnIAK5m52AQlE2
zS2qXOW5l/1bY/Tf+h2wIeHoTz1O/1BXkb33SQRE5JUjvOUHTsNFGE8/Zl5UHx6ZW2OAaPrK56DJ
hsQSl0V1O86fpmPFtyvjHNdJkC/Nb/hL7o4n9dMq5RAfnpCp6RIrn2ojOTjJomv5NwgLdRcKD47l
hBg12uW51EYdyRmm4f0HdM1zsoKooZmDr86ZMlqzOMZed3hMrjmOKubpUhI+tu+TbM1l5uN/A7q6
6MJhhI+QzFiTzO+JcAlEHctowA0Nbd/GrsVciSrlXZ0V4GUM49uydZ4xCW851ZOrYMPqlLNacmjU
GWc+EBRdKzhM/Roix5sYNGKICtwR+dxPVx8nWtYFaz8fYA6pMnrUd3iNhwYtgI+h8f3gSl2ZkMxi
3l2C+dOOgdlrd+cSQmQF/jhDuOvIeBiaoCFUYOdsvKqzJQgLRFQRDN7bgApMzBikFOa7YdvPGr5T
nh2ekvX3ngI0i+8L0d7xbvELV/Wb+tbu9dcvTCtdR9dT3/gVQ8XrXkv/UWFWfQwkl3eDehKq4VSF
TagmhJMGCVnOsxb3SkGSJ3WPqtvQGJWWKCSMRResaHDd3TwrNLJz7Ne+ck7e7NF2aED6FWRixaQT
okRuegHZLB88LQHHIVAPlKmVKmLWuBE7xigzf4NCTJaBhQ4/6rWm/lUolI7L4gikXzIztcEBghmb
5vwI17Eog7ForP+uEhR+d3fyBfuF2Tk+pwPiZ5bw1qQ9L7eI8Mv1ALXk6eLSYKquonsdfghHBgt+
P7UDGV8N8yCq7JR+TpdJ0O+MUr/wGT2x4OucX4GkTR3dhnotMxZBmLy/wgk5OLqEJNvMyao7ZsNw
OQEWaM4YknkMhnpleQ681SRs5xVSvyFb3kTxEItgrIId4UKt/S+HoqLnbTLv4VqaMpQ8+wmTcVX3
yG3TdncauDKeYTycbHvZQxml5JA9qRlGEZMUNVfrO9A25ixgBBzPMHnwlMHG8psZIZk2dUKmitLL
pzE1FDDV+Or0rNfiPqwOpG53Dx2okEC0UvtTkwXr3x3IkBEBN8ibVQit8rdyOiu6ROUL+AoH0O8k
TmNjR8grbdsLGFUJq7nR8E8ykgoBKXkwnRew93enOl4RFLM1S+HEfIB1Q49wnUwF4C1YyDo66J2S
7gcOyw4kK7zpQO9HSetEoun3qIojpUcmimCAV5jYD9aNEfN5JpmaI8c2zVLw5ooC783kgJ7gELJL
4aWuuxQO0IhuKdXWNtIKEetMGu2hfndl9mk34X0+gpz475+ZUd+dC97d7iJU1laziwVRRfF3fC1I
R95wA6Mm8YaHqKLJLKylI7Je9NpOgXV1eCr6EE0g3+1/8n9pyVqEtRu/NSgyTfUK4eYhBWr5fsSE
WtebdzqBDCJfRp9bjxK88WSxvtWONbDtynP84bl/41yy1pdt5CD8f4053tpkvgmrwq5Id4lxXWo+
9Vhfhxq5wXlEU+M6/TgBmmX2BmBWS5KPKUmBwPpQw3uUV5/absW6bzzu3r+UxK9UlakeEWyuwAD7
fWc+r1sBqlXlHzvccNLktWrGSAMVJFkkaBzGCanhOPtQA75oADe+adYwzSKJnDL5wtK1AR5uEgyz
pGKeYIE2xYhe1AqcZPC7jY1pDZl+DuzCdiA1RDyHVCyqu8SFkpjz53u6p4VF3WchiGgX7ofuzb/x
zsXJ5t1MLGGWtRInlf3+LqbMKDBDKUezb8SjQ+XrOCDxGv6cXJThbS9sL1QIiFJq+lCxIcQWYw/E
vwgPlWj3v9/2qzERtXIC9oQ4Zel0gHh+Z9BjjIha71ycsK7ufjGM9CsGdLcNWbPZf0JvplI5qOa+
PWCjyUAhbkAd3DstnKw2esaQQamJNN8nUneAc0MD/k7YOkgASHQtXn1o+vtdcZJI6+2FArkqgSS+
JK5gCbALifqtkx+wM0BH8tsgm3diwjzmTxdUaLULADti0eSpBhsniHAZ29fmizLIjCGcJTFfWw3l
6wqezOlrphZy79pyLfYSQ+9wAU8ndSsnOb7atRwXsL1vD9AHzBZ0024cgAvmmQ48o8w228nCAfsP
xMaP2mKX8v1Bkz6LotZ/HizDch8nyWFyX+xkzIQvUnPwCDnwBE55FCT2SRuDu2erciDs3T9L6P+P
u4pFwDlMdZVubLYYQdzCHsnnVPdm0DAtIz+wXEGq220Dbdw9nicS7mLaZiExXA/qQnNVuVF21iIx
OVT50GgTFrsktPVK3PU8LymLbBntfW5/AsbBF7LDlKG+34qFXEhSp1sW/ws+KuG5UGvQ5XomELzy
wV4CSibMPiDqLoLYvbjuNCvtNfRdl+lllUuwNMeS6Bo8gg3VZ1A2AnbRAX9KZ3mVBfB67mcn8Sv5
7m3SyEST9GU2xHK32mFOf6EF9WlCp6k5P6FRsJEmT61miBcmOvGCbLG9qMmZNZMGyn0GUpJJCyH9
txWAt2ucyZu8/wIj9pT52vSwuYhQw3/Gi2G7WOTTco7klFSzpTDODeNd0wUou/AdIPHUL6sToz+O
7U3KcmXG7kSGfkc8PRMPmUS/XJPxpg5EDMVNMSqFcX4R7e1+2XnJO7xfjRhtgC2tmzrqB4CrTvMD
clXmAnxf9S0AILFh2rpMg/AxTeNPYo96IOJykesDH0d1sAXuUdtqVFe3BydwrfYMr/fua1wRjT07
KqvuGgrVT42wkdrSfFhnUvmi2UVqoyS4QFnagXXDpvhEW5V4RpXXGQ3mub+FVEhdpcAAkOe6M8LV
kRYoi13zHj5uRZD/OIcNt6LyxPGvYw5xc9M+MT7p10QuZWDSlOsAbaSrjMP3vU2tMM+UHaLbzVG2
AzknJO9IQYIqY3Eg4NBAVdgsfWQQi8rNNJGQLvq4/R19ORQqUXduvmf+xnrcX77h7yHyPrW15Ymn
QsPmNxlgTb4eaHWgVMwx1V1GUQPxQwYs8eqT9VCcJu2RJq5LUfaBL+3mhO0a9s/6QgbCYas5DMER
yZwlVFsyz6/2T0FRwZzb4gziDK9c0A+MtwEmBQ7av7wkmd8MpwNBxgKOJHSWk5JnTxyNv9B08UxQ
yZ1/8LJQa7vIyZnIWy5sDz7/RxP8uxvhiRrV2HUr8VR8AiY8mlgZ77D2eL6nfjSyWcIkHOlEN9kt
2MigDRRWj6byR5NqEcrlHshhGDUYp8Qgy6Dd0B/b/b6Gj128bUj/XqVGtlDxtkqLuu7CIgEJUd/T
SsY45J7p2Yg6RH2pjvqc4S3T12RyjP82R2KcdK3QHbOEoaV1qRC6sSiEXHjjCgNqVGp+8TPeivQI
8VdtqdoW7grgcvYcWcv0hQS91A4xLOXlXPrWPKE8uonw/jowgmn9Irta9kYFkrnjP0ik6aPG8oNR
Zrng1+8kfYt1cuF8bD1O5o0LypMee3x4IILgnvpag6kXLdNlzl/5J8IrBMTO4s8sYONLrTBVVnKU
9Ba0LaFRmZ2n3PdkbkcVr5c88FAk+ovfYnh+FQfElwL53CDPYszy8/aA8mZXbIlmqbzAkKSLujqD
jfj3/8O5fpt6cl5ZC9bHOoU9ockHd8kUBrSEIofGDCI4Z1ZXxLnmJP3HGJ3vDz6KWk5gKrnhCPNx
AqJhlIIPNHHC22jQAPmgC9tGoEm/3ZvzyTDtXs25LoCRZRCm473r
`protect end_protected
