--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
bGb/YCQyGHb5tZ3ddRj5IejCoot9cZUVK3rx5C9C1ismglYr78VYY76Vs7uuU/gw2EzK3gwETm+C
FNe0zS9/ct5C2Bkd6XV84eQZG2cagzN8dlikE4jCp4IMsf8+iyGblzIhBzfPppsKty0+tuJ4HWZW
d7gqCeWkx0o5h7vxVsM/0RM3mUC6fWA5BS7ZJDvx79gJtmPxEg5C+p/SRmqCPwsvHQTgOEqafQMm
ZGieWCydAkHqMeD2kyIWyzKzjbDKz4JrrMsbtSYDjZV/i9apo2Qxvymvqa5LwEClVHocJmvi4mK2
u5Er65vvw/lJ6xg0iXafH+kHmVbUZ8e+BEAz8Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="asX49h3Dur/A0j5yxnts29pgNIdoX+yGGhkIkQqoHXI="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
qWKLzMTz0ZTZASVRz1aQ6XP0MmiqfFEnpyKNd6LeXOCZqzlyLTH9U5MX8okefIBNkovSrbBsoNQ/
+D+siT8Oq3OTTXv4QGP3sFAgdONSgFPHEBIJjl2/VR5t5dYqFQ3Td1pst2AsHevaO6T1S8fESr2Q
ca2huAbXXJHb+xdfCGIB0h0FKUHk3zcTCVQSHCJKy9iS9BgnbbZFEEWH7iZn+/olRvQqW9CfjlG/
5QSIQm0baEnS334GWhExPJ3UDH5lYJC/DjIT3tj+SUV1BI5zbeMZNEs5bQJRd3onrDnimw90TaIq
4+7rMrbdpSadTDB3H7jT66CILI89HjPJyeyqJA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="R5wW3Bh7Cy00jAS3+9Uz0Q+dKkcFJPc5fqj8473Z65w="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34720)
`protect data_block
B6uYS8X/b2e63RVaRsg9ci8eo+7dSsL+/eQmIVdJCIZM5HWmEZvgP3MJWUP2il7m/AuyaDtJZoLO
82gOdAXTbbsIjnQGb+bhMBLrJ2DiUNtXDKz6N1xMdJPxQZqufPVRHeoHuXJO4uSEAA2DL9VJCxvZ
cNe6UPWF0ye8Bwg6bBXqD7UaMPHTqe63XWCWKv8CKGBYqZJsHvYMBTJlCNef0Xoe8QEKUb9Oj0A/
TfFLaHQDA85umTXyuyeIuYi3TZx/wzo/Wc7n4YwyYPurm8uWENws+tQAU+wc29z4ilYdzpOITNMM
KAGiKdQJBsrmy4ytkLiVDe1uciGHOja+aPHMCqGePjn3HCe4UprwbRCsQhHlD7I3CM4pT6S4qo0y
2tWPba0u7LEBPXtS82+pBWF0cWefWC3fu3fO66TonWgssZ0/vdzWle85qXxr/rW+nckF0+6QPgVA
ZeIoJX0lRi+Zj0f/40lesO/lh+RuCMo45mmmakK5x/qpmMuYecM9JCRF87agc+c7TQTGxC845UxC
YwOdKtlGwAOq8lQtvdhEZ1fku42/b8Lr+heMahe9YYHl9li+6NHKl5wT8oDwNchDT/cpAZfzsi2L
Lc1mkIKsENBSMUrcIV8prIGusXQpCqEnPsVEku+jyvAICysKDdtHkr6KoarudToZmmfSmq1D5Ml9
R6leGf8O5Mbg/PVK7rxGJXXp5Ervw1Krrq10Myac8+Rpkc2shLVfMtrX5zXH7mXM5fSPidD7h/ZM
zHdYBaY11bGtbrtdwUBEZIBvsM5wb308joCww+Ity6yo8UvnqzXxOMfRB6/2QKHx2l1zWrtAiYFE
p2Uz6uaPRhiCQEPBJVTUYw6oRoiVWLE4K8QVM7pmdSOcTiv+IRrxwEYd/8MCQq077ZmTOd62DDkM
N08Jbqppe0RiCrahVD7YTXqR/+Aw7w7/V9Sct8bVzMHcfuvH6Dr695H6MOVCRAwpGhH55ci+NJ7t
a0UoFPSaMBWlgfU4VNOrwkxB+FjU/eFoRclabMuwNyvFPes3o+UwM573LL/j8OHkJk49HL8n6QSW
IPjmuYN6VRG8ma3PcklTwDdq9DKVvKa9oeo6Mn6OVEeWBZLQKPy2viY03pOFOnvdZ9Gr1nOjQcfJ
RX9/+9nRnaKeNq9EZc6L+EiIPo/Jf/PjJxYvciJvf/0i1CtRr8PAYu6OcV2xr8+j6qrZ6YMk3iZz
BMYl3jpDF4AX6ud6w7UMquoORRBeuQmr9N+ZCl46plmZExStJ7U/0hvuXUcKdF1b6ImzDPhety8c
vNQBt2wB9AJ8N9Kvn1IrS9xc/EcY9U04RToauL4Ux81UQd10kwbdyhQuHa/NIvbF/qizijFCcK5P
QkLxGXU1R15AIV5XBp+g/GbhmOJeUBK44mA0Y8qLc1ogXsc4J/o5OJXDLTCJoFfl3IKNFU/48iYW
UMtIS08YJyTejt0UDpmBCtNW/eJcUlGk6Z0Gbl1Jf4oJLA5M23vaRCpWagWItrI4kYfxqAEybpoI
Nano5jlFkFVA+2I+LDN6FS0XfRTICWQuKFaLH0TtkLD3LR/tvtfI5VYHKuC9mVGdmCPMEs9j9KgQ
y2grXKn2zKuPHwCfZ0n6cyGGmjeG+f7zhhLf8+TJDqCZKPJDGoKykrN9vNWlFJmWPdPRyM5TbCYw
4u59aAqPhA6H/UkXc1TXyuOoCrQMgnOwcUVxT9zdhKnFYLN2twgMobZc7WB+jWPDbOg6ChOfuyvK
WFpKruY+6ELDWofyWOQLsA2Qj/2UNqcnhNxnkAHmZ88Q8GoDpFZaQKlzA+ArK4iBPhfIaEnsCje3
CjkUhLH5MXNRKA+70htjVKYbOE8SL6FycrFcicvAdkamrloGv4+FYS2dVb2qr5F/pI1RgmZBKM2k
q8euEjP3P8sCepVZfcXyT8CI4eUB/1KD7gK0mfE2uFFXuMMC1vE7r/hBpoBgilt/IWb42p3ICYNj
gaOEldvuLfYHFZFbiK/c8eqc+GfRrlAGXHwf5m03CyDgdu3g7Sq3+f2CXc7buyfhxNXRpU/xIJBo
ayVUE6Wx5fKkqu3nW3l2/DsHxpzpAgdip/SoO/N4zTU+vEbt2Y3epG1WMOs3pGXnBNWw4DoH9cSr
dw+lEQr/2rQiL0kHyqeD9fz6Jw7+SIwPQChmQs1L73qvwld6DTTOpXMEU5IfBmnxa6fUOaaY5W9u
0sdxPJoGEkf+EhWUxl+A+opENDHmWXmY/RPeYlq1FNp2FI1T/1t0OzbJM7wk04xHSr3Ky9wy2u+b
K8JfpTdGGKBg6hsdELjvXN1EsSVjEsIPkwVIzeP0NSffXFNHwesVmgOhcy/1jgia6pAxuxOMKxGO
DB0jO1IKIsBGGZPA1rV0pTBDGLxivVm70Nh/ksCOsRpAW0HFp1js2lvTtmQcpcqVRDLSIh/SfoKT
vAKi0ao6SWwZEhTT73RtegcP7oy0nT/8TiBERmh+BJv4ZWWOJ8+KPVIcpBHCltetkMIzjbt6GiwO
cbttzeI75ekNxGuk75eJxcEIXe+2QjaKWWE0ImIrNvtH4oBhfTlVjBbuOtAp+oupapOwWfMGcfr4
9Qv7UJ0USgujoSPD3f9VVY14Ikzp/fmaS8jsrh5hzSKkrRHm52EOYBLLGT+1CT8GeTg6OmqBuRGo
QACICZbDDd1iL6oUv7nubbcxGHhcudmA6SPhyPcX9eoKogEZfABzJpJQFaMXRuRDs8nr5N8LKiLO
zek9oGOIMOjtuLNxaDya2TteTEu5MyGwL4NJF2EPu+DLtXT/T8AOFYjj2/0bBn4z4Mmgoi8eYIdo
i5OQ533Y7cMQZY9LkKYg+5LFt9QGEXlF6HRZKS3E/S30n7TGS0DZBR9X84MIU2/0dzYlP9s2c4WU
5BHLHzaiX9bRXMLtfZauO+WLm+hI/7Uf93xLBRi3LNCXDSTn8LMLDykbFu8GMnt+s64tOaGQMo4S
ybSvggtMn0vMc1u2mu+wE5w7ZI5wXF+sPq8adtp8LmRQU0yTN3C6EUhwcRfNtnE9LRvwUMNsEU60
uUqWhnDA3PuGJ2HLIYqCOYzG/vgYHzTFUPS2SuRdVH+8ifh8n0+RXkAkunchnsmpTKf2kUOtyttA
oWFPylY14tsIaKIKkxPwgc9zN9On9sxjEaw3L/WI4az6+16sCCetW0FrBccNr3U8GqAi8nqbuVUj
slXwAY4f7ieszw4ZSNT3Jc9lh6KloDxcBQVzF0NE6l9se4ZMRzUw6NKZko0NihAA4X5AtzOJGp2T
fv/zY0XTx3922tdd6sqZPlpFXFXPkH7aONBfmP1se3z/k+QTfqSQjF1xEnK3gOv0o9IgsDm9GuhM
xaxcBnF4H0Wt0m/3lWaOBrZq+w40ph6V2Yl88KOkVIyp+iUvz6ZFrwPHFX0e/nME1TzqH+Il/Q+5
34k88nDtWWF01UB0BJ8ffiRH98w7lqNPSI7y4Ab7HdwCiz5/WiD7S+48/8G7R4yalsnGFzSk1ptK
eL8H7DoIC9RMwDKcfGQP82/EmZHTZopnfY5SRLdNKm5NZgJGO1e3QixiElB2oj6g7HX92HvkW4nu
OytqBSise9ueR9zkYRc6mBpmaqW+gqUO4PNVC5tIM5e4ieXxNiHCYJc6W/OgY/439zHuMftnU7LN
PFW44TBsyHMofFkia2+ld8eD974IZDBh7TJlFxfZyxBZZe0UXnHL7tL0d4ve56fFZSTf6tuwO7Fm
hfUX2kTEAV8HBTbtZnIJ0wf9AoGP7kXNDLQY234a7oGfxkZI810qiZNiTIrlBk9h5ihm4DHn6UT6
fhip4Ylltk0EKDHtCee213zymMQi/eKzru+ngfmSGI3JRsD35438EKKOQayKJViSwLlF36G+y+oO
vFqnvt9b5ZhB3WEvVtfWWmrXemSKq2u2Mt2yjyL6icr9J4trrr5pPrL6tYM6D/vR8bJqC3k4GoAH
ntkMRawgGfMTXllkemF6X3UapYxIBnj/k0+ewQvmPCwerv9xnt0E+viHt2UlM+xTokQYYxbADQeu
sjTGigAqtCY5Lw9iwQHjqNmwdlB2lS6xVvt3inPaOk6cj6gtJ3fJblyhx5+/6wmUnHCExNPer0Tj
MSvRUxTKCGVa7spkTiHsYHne9XXzO+56vCaIbkMaDJHcVIPFRlWNgMJEXuM8aXMX2oqms/abqizL
CDyuh45Mc9fTzSQu33TWlc72M5kfrYGL5NLELOBHh8C9w8Abea7yWwe05D77XYYobTvcoCZLHwZ/
sEeYvyApJMBOxJDyaB+mAWfhInSstAwsBNylpG/p5FzhcTeyC6+q80MU9bon3FgALjVmYLXPRpgv
zqBSj+WCg1PQi+wnyRzDodBnROFbNVlWgCEn0XzfpDF3vdc13jHxH77RhpUvLzi8K9bGNbjNnW8F
XlUN7kfqg+9IEOnhAL7uL6Rw6D2Sxw4tgV1IwlIpSeCCo0AiD4QKwIk6sgaQVJetBQ6EJojKtL67
W4THESmdSaMRCcWK/5/09GhXHNIWoKwBduv7vr9SKh1BySuKB2Wu8XjgJMdjQ9VOtzfoAOnMDzbc
mCUX8YY8Txeaaq9DA0KvwR/o3mvuDXlD/ql3D2BoNe0LgVzecRuVPkv7gBRl2QigSMH28ZfcaWFK
kXl4ttArHhAYHgb//rn5ibgdnNx4NsU5ymg6inBa495xDbgg4h72siY3tVk26A3VazCXbQo7bcp4
B4DiT7EznAygqNQQq8ATMX8enFoRIxDLyILH3XSLCK/ogRfrRXdWEob2Dpc+IpOM47o0O2b4fVIo
Xavxr3CUm0C2rnxzAVrcxKgqHU7nqsxpz7seAT/e0i4C+J9SdJ6RHRXAG6d7pyKwhlGpeZOoi2FF
W9WfMpBmyBh0b8zUdXSB4HgRJh1OtoP4rZYPt5nm/BPXI0tXp7yTQhK5XUKd1AjovCBypWeip6lX
LU5jbgGRK5Dsx3BCyL2CHUL4GycV9Xd1EkSOr0QxoX21zro0nYOKb0WaHcLeF4zWqa3JNNxzIPDx
gzAYRtb7HW+SxbgxIulJ3UHdjlAcwEzEwxxifAvAai2RlC2QB1RxTHc9zPYSISJaO6k4MpJQwgWw
KXTISLZT1G+XTcdSx+RRX91+A4FEA/uqt13ml20l25XiTmTNVd29rwfSWhOAIWC8g2RRiOT6kaJL
MM1wAwb/l602v7setK5nqtxTubUyn/CHBvL2biurKhwTkKJOb87b32T1ajlwHH0fawFOGN0/XIz5
scOpdKdtAfxtPTbP+2pKNCwIs98kX03bfiFUHiDebY6SUqlcM+NQ+XvQObDMdKB6bMrV0ArIWRwr
MGWJ95oZ7TrMkYW6HxZt8VZ2Pty28vCY/33Wov9sMnfWaC1mBgfdP6cXYEJ2HSP9gojinvxz9wWH
0MwONdMuhQqMSlUMAz2y0n/G8mUlI5ImS821wINWcrA2nFm/Zqh950btO4mRQ+EvwZjAu9RhQ539
/2if+XLd3FUi7oNcJanUb600aYKecRf3qXRiY9sf16+YF5rmaTtOZanv1rgpwhxSd9hY5ysT8JxJ
Md+Nq5cAHA0+9/DL/xVH0f1QdrxcM+hXKlBf1Syp/ojzHcUF/peEXYp/9d+gzpwvG0wizGKS5jyP
bwX38O5sk+OyKRzm/mQKOv2T2gyaAGeLepzpEacjXGbZ2FeiPJ5FJRmWRIFbRSxmvL9Lvs/sccd7
vtOzcRGLo6yQuZPpUFcgmTOfewcZr3qEdptHXOpmUKR8JgaCRhvyWMOdoa19UvWzMkPl6pPRVsGd
4eA1GsL+k9GMam0XcVZscqTnRpvMRfSYOLBOkhEf6RTKsWjMO01Jy9tm8lVDt2WgA2B/+w1NnSSp
8f113LsGmpuGyNK/p/6baeXhR5piPEw8eeS46kfv1GAylrKXQbsZ7a4vkgwjIDXs/hpj9Lb9iAII
XfHRcmLVjAO6bZItNw4BiZF09RPDcTw4861wRXz8IHHx8ECa27uxD3HCC/dCxpoLQQ31MfBoh2e7
uSUc4XyVindaCmFxIpprOxB7Xd5gVsH2YqDbUkqovByrViK0zUnNeCOheKavGmMp38ZcOdCvejIK
sgYAo3ZWMunQ1lvZB6fKPzQqGOEsqKv6mBcTC9Omf/m3JbVBnCxhRchFgSExAm1HS5Yc1STxsIyE
9L4apumf7EQF/gFKgP7K1dGsqHEgR5ydyANN5asxRMr17prKvEtSN42zrr/tdVkKmBrbGb8/pIVS
F1aEhXFAGFUNoGmJ7IrEzOvO3HTEZoJE1R9ac8BJEAJ+UtTI4SHdyG2k9B+ZNlkt3+xJO/lmQT4O
E9lpVNpARg+sE9aJuR03wtX9r9q3tqyjWcx0W3AaVTIWC3p+h5YlSo3erGs+PML1MkCNLDm+QUpa
6mdDpmDAcXVWURnS2rzBfbfg2FrQKvsP0tlvH73Bt19HwnzXqEnksJmdNdvHQwtQuJkzE01SYpCf
5WOMwdCOfa/ZuzpDfvF4CW+n0t+WMJp2/yYQBA05dx00QOn8o4Lxh0u+mYNXRQbqSEUyaTMLVn9v
xLR9kUyRJNsnZcyy97JXAi0wP3WH/9exLai8tVDNi/uqZB4KeHTFxlKfJe2MWoDnjbwLo8aJ87Ri
ZAGRY3xdHZiJZSqIDhYvyI4RiUKeWNuk+aMIOkkXzx/fQvLmuvK7rolO0+chm2SL1l5ncwfbCiEh
0akzPLhJaBINHWQ9BvHKQxCEtDNtxm6Hfbr1QhqPincwcUU7TBR4tlSFhSl5oSVdHMJF7GWT+0yr
v2vC9SEgYInwFJsw3PpEPn8wEQ1rquLjafKEzY4NIOL5othH//+uPnmU2D4evz9FhXXA1ZLDZry6
ilbd4Ls+ERoG6DRoqfbQNWMM4ui2Nshb8AXbfEhyLReS2kQWI/RaM70/SSbDWj16S7jqCnzhjjlt
X2yZujy1Bnd2F7UhrQxVnWe6Si0TTX+AN2PPZyJrRt7RDeIiwk7OjrLOXOwkKaH+zG2BkjJlg9z/
Tr4llW27cPjWt6wEcHe6k6sy9/aZHsv/yHCwDic6t6ReGkcqh+Xo0NpzGSnlMmW5faVorgYRfCbN
O/76WmHbym+if6LPuRSdTP7RKOBKm/g/Z0k5LKADZN7EPzzeIWFwS/z1arH99ALTYH7kbZb9P1cV
H1STrJqbQiB0TrV0NPTBVva7VwRH0n56nsnL3CqzumGJGzhv8TW2M1fvbQSyHXThAZ2cN1eHMNOi
ZyBxYkivJDsbGLw6yAGVHMDLMJt1lhm5EEcpSaYNHTls7vydPZB6zTVgmS1ajWaYU0t54axZSu4P
bH0jOP2XkWwgimOZFpAlx5qIgjb/nEJwcMrt0WrAas/22xrmCDm8+UxlHMH//UWE9z8ZuOPztkeq
3edyGBh98AT/BtmdBJLOoRgGkLejh7+y6gfhfg13w5+VVRxY3CdVw1V18Mvf3Gx51CMrmQDHkBxx
HeOsnZXrFtvw43Q6D0ahEeM/5K6vguqbB1tbze4WFIy2sdzn8N/yOu7oBduzLPgv/Wq0t1wN4sfg
WMiKZxXmZT+TO4PYiAWm/naGbrulOFESAy0cCCaBm2v0X5+rj+FkgJu/0e11vq436oqdzvNJLyTR
UL7URLn10tkniuLFgbxdIcRhbJLpSrECtZmRcOcjTF0t4R3RTwsCZ46zjaUTLWfg/lo41GONmKvM
vIV9Y1DeF3KSPHOcshDdOor9+JGlrblVSCNN85pT8ZmPVa9U08XQrWxPL4GjfD//ZvQkIi4BLhVU
2gn+DuqdjIwDtt1oHDEC/mMbKNJr4ai3jxTQxkrZpHbKzcpTmr8wdm5E1hqtQFhMR0BGWeUsr524
UbgTK6P3zyxJhVSG2PFsU17+GvaWOjuKBVhNJyIur2nUw+lX3QN4KJTsdjw2YGGYnEEo5ykRhT3V
89qiusUUQ8SgMzqR+swPZXU4L+tsFO+b2Ir6XFdUvV1qZnbj6mb1pwNsCMazqdqhLS/lEd49G8/r
/FQSgBoCnveuLKkq83KYICRAqrgQ8KGUkRrC0BxZB9V5TH/O2RtCFY4EXkr+RPo6uc3kWGWbYABQ
OGcqrk+vFkcEmVqsRGtGVBquqqtQqeufMem4g0SMd+jlaO2bW1udWt/6cJUIagGGkkmGlR2vx5oX
ERl8ZfOAD44DrelWQRhhUZUOtBKJg5ZarYy/nxKgzjsWC5E1CYn8Ax6An40BJ1C40y/7yib9qUJH
AwaTHADRAKEx8RLJJCqrA5GDj1WJbtjtw/Cb3Zu+8QyhbxkZNpnPzb/J8OIohNjXY7kmRf2G/S3y
6Bs5j0nSd5n4MBatPLrx8FpjbAR1UTOftoOuwBq284mt+YgS3jDU/gQFRfl3mr6o7wj8dibzkqVo
RQoDrz68+gJwnlpEYcNJk8mQaFVoK1X+mmwduQKXRGiHIusPQbLsaIAmm7/QJnToD4Flgm4pr46u
2CYiu9NsUrxNnimZOliS+fwEbM5W04sQy19QUPlZOniCaWyFx2aS2CuoUKtvvV9+9IIzcgBKxnVA
/PPxqcIdtNiXlmb426MlCWzZLHEtplctDkghojAk9GR7fMG5/2VQvBEmGEIQDf5mIaN358nM93ex
pskhVQ9Qq6KEQI/s6JObjaBPe3p/xVH3l7lMU4p60rDhxCI50iOp9JDGPp6RjdxKDhOQhrCPcIro
+Uo7YLTUMfyfNCyk+emyXJ5gW+Tz8dGQB1YvR6uEQP89emAwOeEVXcCuc7XunRmh9UmjGacNX+bA
F39u3EODMjK0oZcrBzbhES4mL9NDm4PxctIbBFJM6RIdyglhCW5XmkXx6YWgrDs94asqV2LVVgiE
x6E9N8NIksdn0FW04ym20G40DLGTLovAiZeFv6Nn/zXlTp4eKYXGTuMehedAlYWbgV0mSbYVVaBL
RaeVkY+UQ8/7dbwUKfkwETiJIOGHBZvaWRDtvgWEu470MZsT0S4dRGwlXxCW2Pxds8UUPQxPqful
hlKjdVh5T6ebM60RViNP3TLTLqThX74Q+XI5YE0SxJj+NRDTJkj1sCZVP3Xvi8vGW5lM1k2mHQgt
eo9VI1qqmWaGda4OPQycQfBxL/UesEkIJZQYY/TYfD+xGyEc5RcHNkQ2cNZ3OTmcIorO6Fi+DBDL
BRZcO912nqV262dtL8K598g4Dl+W/VYdK9ik86xcKYY9seVICKwTiq31/YcW6cCwxCfvNxeMCzCF
ZDNmYPBpePy+rUmVJdVlcCHCV/yKjPp4uEfaQBcatXcVPfPkqjRfmsY79pnY2r5TImXu2x/uX9NJ
5I/cA46ZjGXxdQKTIX233RPOTnm919rbIvnHJFilbE/6ntZAJ9nuvnXJ1LMSUeD+BLEYJD9QDbDl
hYViHkBVf8DMja5pOHYz3bz16D0CdeoTS/JSElipnpH0+UA3Glr6hWSIf2np1AXjFNwvZzP0j/AJ
clB6/P1YVpL8f7zsMEnVqQDzyBVH7zunk1JcMgooPXszN0w2mCaOYjp2zKo3vMtONBNW0H7rPt/3
TmkJX5z1KRB8lcSZp3ilvbj4x0jVsSkmP1Ksao9qLxFa+2KlUZfLLBJwvkNxwFdwAhKcwKSmnINb
wcoonOlFVTewK7GMbyjQDDNUyZxK7sEq8Xld1NvDWXUNR++2PoyXbNaK/0aC7BojZ3v4Jsaz75jS
sGDKf5Q/zCcUcLU6UiljKTcs+XCl+D2kjRm33iaLQ0KQM34ViVWhREqgBHlWFTKUIeW7zoKVZdz+
YlloUsC1IbA76TJ12Vi7uqzQUSqtAJY47QkqsfI25bH+1se1cVWm50dSmoWwADnfBb5PQn1jIejI
NKu5VjyiyhzpaH4qitdkTZdrKuOG24h9KwcD4Cd7GG9vQ3btTC7Wo1iLvykHx02EgAOTfEHem9ol
AnJB2XBp4IF+OCOMy5YhazKVJorsMrw05tTwO8gBD2fjmMsr54Hv/e/HRvG/WiwTIzUyI6cSd03M
WtII3vOInQ1hHlExLJ5aRtQ0Ez1RW571vQjNXedOru/HWfJzUvPvVXGZYlTYVvRPIjPCXYCuBcFr
eN4ti5BQB4kp9/9mFObY9fgYABJRQAU+bNt3fP2HfHxReTaF5Xbe4al02NxrsynONSh8w8xaH6fX
W5ZrPiM8Dq60NBrlTeMnTrM2/GtTVZ9yqUHb/XPpJNruf5sz3M3LAhJJrUzA03UIGBdnI7TJ8iMX
D6EbpA4b4lufaxYi4hAkBK1sP6u+ZKtX8GPaLfFLJFf1ZPoaI4LkywPFZ7okHkIXUnjn7sjm3krw
Vvd51SzIUNjOFRVhEY1VApp9kq7AHeyvv4pTvq1EBkWC4hCLewwD5JiSQVHzGDhtIMyoykJ6bNGK
/QcC6vv2jMspz9K+OYPGLUoB9HOvDIzytj+VedZ3tI8S/rjD0gRvbhNKPOIszbCPuEy2i/pu6DKx
/3BI33sOs5bf+cUTOhon5yjcKqhDGaaDdNAXt8yvCJG5oXYMtCIaihhVDl/23u1ie2nkg4pnVE//
jAOnky+UggTC78BR0T4qwxqlG7WNhPGq+bfdzb2lOd6aS2oy38sZ976ZVP3WN8vhgLEF5S9edI5S
NFy79S1z6JLW/91ln4IdBQaQqo58Enqe1WigOqvMOHVX5x43H2tZNlSbpsH7OsnDXHDX6W/Sw3G0
UOVqjjz2CAEI5JKTjFd7BGAnMwyfwI0MOEp34I1/syLkn8iyROwoEoB5P02ct/RuCmOJMdyP1q2Y
/AcL7GhVhgJMPnZeqPjdYO4JzkuYCLisrSL3bpo1pKDxZ5Ypqizn0jbTjtGgxFMJDHlIRgmdYwgr
zvKVf81mozNHLew+5VfZRcLnp9iw7nlJbn54mrL3o/BgpIu6Iutvek50R5Ha5ofZbeIFqWaLS8qa
6zdEICum2Rdto1W6XMZoYeyPd5dUHvP1dZQcjrBY5vX5mF0xuyZZawb1eXCE9nTMQN3jfWMbpHgC
4u7PgHP9SoDxNiufhy9lEvNjnJTuSH296DLB8F3T6hrMZhSU7Y4Y2WplRRKV3GcnI/5a7KUsn4MR
A/qZzR+0ZdqfqvSyzxbiIpvuYzYZfU+5OAYcQdvxkZRM46jg4LdrG0Ir7RE9O9aRXn3Ng05PEh4U
EqAUlLVI0Q+XXA5LyG27o8YFUaeHlQFOT7AKXoovM1IAHdNNBR1Gzn1LoghCrosBK+ddKdoFyLlX
4wKGWLpSI2Ief7rmu+sAhj97l/a6fqk02RsR4xeYAL61NBy+CVJ1wfSfaxTrrghFMG1Sg5x4ZnDf
XpZsZH4s041t3zyNAnVS85T/VxQLIu7YtNuBFPtSg1oCW07oTdCHlzRIJREgYo0CitGvhD+rgPEq
RoMkLmWh/etjIV9Vs4LfCtg7JVQNCIb+YDp5Wail0MEIJcdt9dI6I32JDfQEfmrwL9ZmmDNx5zuM
uBMZFHW2sjRNt463jU3PFeVqLpWB6p/4Rep0bfOy4YyofBjrgZXXrm8JmNLGccOaGWt2kqn/ApgU
ilKYNiIrh4dQ8NQhcx6gITTAOBhYRLtSALDOH2lWN3jGGpzdIIXIB/I+We4Emc+RyDEdB7jtVfsi
IdPsAgXzS8dcXV0LYgXWONbnFpn33Tz26sESh5SIbSeyzh7dPx4Ljt9RjxQvHfjlG/iD1uW3mnge
NvjeGCDErLA7C0LT9tWR96e9K0IrJWic+KnIti7mMENfXiKtB+iYSyCa4EWhUa9pe30wqJ9BZnum
FZgIMpZ10KwplnsO5NZtQ3fQmugLKhM3fVvwS1OVB5SQLKMLi4bPCaNSQoOHiRgHEefCBEMKm0p6
q56W8CBLFrMIy/7LWAPyMbfnMCkYVeahYT83FP5OwRoyCTUV7m4yaE03f9LGZ9V+WaL9EOlU3VfT
ywx4WLlTjhrZ5r4epVoLn+f7JPCRDGqhux2A3AFAy8nKD52ZIwOyN/lRPAduDczGDdhO/ah4YD49
EDOwyyswxQ5xhv/g6hb2hDDYxpe/3NXAV8ckU4PfxusTg0EMQcADB7jRub6Dk6DT74XQChXHxTIc
U9hsgZKqPvGm+ZF3Tv+st4EvWfyVSccbtlBJ7P4NQdLoHlR2SH1hGMD1Nu8f+i2TWUCMzznZj3o/
k1zfksK10ejXBQD0wvkQHkbaFSpO05XFy538DXPKlv2OU1QUo1QEJtNuSg2oaG2KVwslZyTtZlD9
zBj2WmInusg8JyyHQXQ29Pt1iBi9b0/YtKMVffsn5RSMmBfv8JkAKH+GhpBQyHfeAajkeFBykF58
B6aFOfYqX7K6Ii+PTgiJJBr2LsnbVGU3fdEnh20lW/Acd0WQ9PeFzte2T+g23i6/VXg9JPwwOQGy
U8Wosi+0mRKE8oggbOIJheNyrBZxYUvT8+0dIESZaFYk92+CjvVTEGmve0eTG2+WLxQ5df6LXAbj
Pq0dAhlBQApBruxPXFSh5CRdJeVFbM1WCK0p5JHwVO0vzaOiRy/UV/VtamXT4ljRKOaYHnYJboZD
nTvIUf8hCUztpPLb6gjdN3T2/1+2f80COxtXxlR/54/yR5e//jwP7NweQsSXrMrNp+fOj7Q3KwNx
G3NIJD38SjnNQivCshcDplkWlAP2CreyDpISGM6FSeXvE54Rp0l94B5JCfAM6co1JKEPCPiyHVX0
kDNty0+D12b5y41k7PxNSBW0HKmjN2CEWmqm11Qg0Bvfpht9fRU9KlqHnU7CdPt0XCyrx91MRU4J
Gdtaolps1VpES+6KkDy/r90Iq2/EbC9mhqnOHlbenza0YX61GbmJkDtkg0t5vKyo4nBvIqCzrzOw
5Y5lywfePc5dcEmc9ONlSUarVXLtAm7noCttNsKGMFgb7XG9DPdTpdjPVZpFKJK/4cKIQfrWtPLB
8VB19Zqi9kqzDFzECsG73PIWGU4obLO4Nn3TsMrB68yu5hl09mNn8Mwz3SoQRrYJy4eFhiCdmDMQ
odNOMhLtq+naAdBSrMVBxSZYB9p+DYVpZkfKOjg75DrsJnSn6vjv7d8ZdoBdibGtfvNXaMyEpJQ1
JC2bHIAcTLl9o9Vjor9bn/XOkhH67O/GXq/98NoBttK7OPXFWNsczx/VCNqn+Ujbi+4iFEG8igV1
SDL+jNGGuAZoUdEkwgFOhc+QUsjyIjAnE424sqAvuNsvB4LKOAi60YX9SJMg0B+DbtE+Ebf6CftI
CRN6EIX85QwuCZSR+VMbkECaAPKCU2h6TpRMSCnnCc8vrWRmzGgopT4PJy4Ti77sMlE/GfqFZ1jL
UWPO/gIRz9CGQroFtAT5A6IEFtuiPpPu04QZavsfehlthaE35b5vBLmz25UDveYLIa4fkMjIhyxt
aZeeNuCdeqLfeWttqWh5tRPzSoQg50efcXq7dLzEqGK2rgza1BANnhaRozWvYEZtboBSBwdQd2BM
2AG/goxl69duOFmo9Mh9igDVcB911YlP4Ut2BdMiWNUDrGB0Zy6+inhNUvZ4Y1PROO63NtTZl6ts
KjjBBoyIeLFM0pOkjmIi6qCIpNCorc3j3E1M5x9hINegT7HBgqVbrCLE1ZzpVWAfNlXKnm2EXt78
R/+Y56SjCJNiSDvgelqC4EwXVqkyxnbzEVmrPfc2sPZpjy0dRbGyHrqAd224GSV5pRcj6kidarjW
DXklQlyeT1J2svys9PUJ6VUvBq+tnV92youJUjsRY4g5kX4X7twtrPcJFh6lBS4V626clsyeFCuY
PN/8fHZ08jWAd5p7kgPrBe4GyjgDQerd7Wkgj0KQpVinfkzAtb//Nd58X3fv/mUcOG1OLfflp0VS
molRpqYzdWnRGQHN0sZiYjPz7J7/BONTLWSlckRg2bS+RIfJv44qAMzLj835lYbszlY7NchwfbZJ
DwX2JTNFRsYslkMY4D/x4r++DyWLBYWTySlj2+v+w3OSIH74+wHlCmBaYcewvd+f4ih2jLEgVy2W
PVC2ZvD3crDtjrh3Cesy7Bg6IvOIJ7H6/UUgc2t9zC6y4kPRGLmY+iIdljFXmbmpyTfJhdk+hS2C
wI0vZC3keWp/h6qKVYPpmPcWhdoCIbgkHQNom4CAGk3irJcIKaAugG+t7qIJ6/NnIPb6mbLBmAL/
qPczbygficrRR6Z0X6l2x574qu0gm3EtXuP760Gg3bfzevuvArxFnZUdEyUb/cdUWsjWV03bIBng
XdC+vfRmfRwMhZyBMo60ZvlusJbLVY0rx3T0EERSoTa0GQ8Pba2dfzE1HKvON6lGoKpZOe4dxV2Z
73k/ERROnpFVxy1zE24nnorb6j9oy8n2MCSPX++MtgPxOBELVM9V1ja2ODWtMhdwKEQNH9CU4Pb2
YeBRkT094JdbmqjfBjMDXLaPoukviU8rCAu72NbZCNbHHXTVhBGzzW3MLgPU7cyNGYMJFYqMjTKy
gAy4RH6sY1ksTLFKieS9f6vfNhAcLQxto5UbxiWyRSAHRjph2ZU26m4IjMsiHk5J1lcZgWy5qtDm
xo+/70EzwiO3+LEpaBb2jKEggr/HR3bdTLkK6VR6OesAeHd/3SLqswlfG+PkyCWRkGlN2wjteYw9
jD0ABKnnH8GllhQDFTY2ls2gUG/Hj0/N3uIdxSWOhVQ4fS9vuvKHI5U4PLcpZ81GamfzfB6hgD7K
gSmXPcyRD2PZBrBGabuNEfoqZHF9t4Ne/YnjpFHNF74pGfGD2fzmH0bJ+eFu+CJZYDXcfItLn94F
5jURviUFgWREka/k7iMY7Ksg3Mpo8wATAzTmV9vNGqHTExLtbYhIy3ssHcgvRlMSADjv826Q0XyW
PJxtLM4qxNJnEedVkuYwqZyqtTx9iOQe79BIB4xN+t4TEzVaeOGt+I6AN5/8+xxlkZnL/5OMB3LW
DKqB5qAgO5pU9b0aox3BART3j7BsWFHyZSwk73QuvK1UxN5sdXv/5rwOrDuU/sMGQ0m+ADHXxxFO
eRz3qeBkLGO1+oTVnAVGB5/zvIOANrnrCvBTzxKPWBhHcw2WE1p96OQYumQKrcWFhHW5Pxq8FABB
pmI3aEx+ajDnup/3JypjcPkCelib84QohqPJjmZDN8kPW/QaC255HdvSzmiT3X/R8tTNlwWHzjtg
Bw8UDoAF4bPtCGy/ZYXLhI+sVSFSDZt5muyuuLdu4qgHRpmx3s87lZY7FHHEp89NNBm3rRsOYDDv
ZadFbihDAtBGZhfZA75jCz2Qe1zBesRDQFWMswuoA3JV0UCPfsUjPqdw2/dH45oCcs4DXa7yWM0E
74ExU/61gQ1WRdme8GKN8ZrdKsgc8uHiB4amEkAtR9w6pTtVL0eLVPTLjmwCCv6VcrEif0NCwk14
ZgHK6Db+npWLrWZ4TnY0kiPjZVWpqmhwjjis8hUhuo3bNk+0/CXb9HEcyAHTJKYkZShkRZ2u+wls
8c9YGwvLhdDsKZpbrzEOnq1IWW5cdtMoxv04+H3vxYQprS0dE2NAtNserK5/8qbfvcupySA1XLPN
flZ7W9C7hLJHzHeSwVD2q1FUqpDzs7cs0wt0cOcn2V0oPJOkNpsTjhH+7RNZwzP0GdkwqLcGbXLR
S4auSldq9Va7epRHW0Um6NE+f42FUpHESKRlTehu5USK3aI2hJnjuDfGEGVx5D3dNY/fn+HB97TP
s4KykpMJqGmRA3f/DegOmmF0BUEEIJzxuU6sS6DPSJ1QrdSK6lCXCy828IsXVWbetBAohNJSTHMY
NNeA0O9cQ7R9r5zWfFeEdUtgUoIaN7udL2pVnoZRWTpjEjtsRpRA5JWQ5uDyF1XhfdIl6vl9gGiH
Ej/siD6coDl/W6PD8hQGpZifUCwevNzG6afNETTmYsQjSIvYR8r5ZPyC99gapop55TEQhTnBsU0l
P8eBtj/RVYqxAGxJWNbd5T+Tse3O3fSOX1XgebN2NERmacBFeQ/3rBkLrtNtsX34nuQTOKd5hen7
lShu/BSMoMUvYBGeFmOtwatwCh7cRN5B47headQJoYiiJfXZgFB9YpSEz/i59gjZ34Ym+6r0i/HV
Qjo1fQFNJaYkN9neLI6zrrDx8DSQBg+66OZ7g78ou4hg1NkB3VbmFsIarzkh+Rxo2jCmLwwj9IEi
kLmLs1ZjMs7KoKK7hJz2fTnRuCOBdagQn9/P/jcxXjBO7CtCi2uGvuLmARbZzhPOZAm68yalgJ0m
kWK6/RJI75sd4q/eqfszhezBOOSbKp+JeB2CJF2H/k80+Or4As/a5ZS0eIWSAvoaYi1t9WLyshIs
E+pvGeW/BLx9wnv7emgut19Ah72EB3vsb7SDkaAbNASIOi+mzRHjc7V8b+58+4QDLJSL37kkZBZo
bLUrStRbD1jQnZsBbNgiUO3w/zoxQidyxIbRxKXl3zKGVAba5tCOBUAQvfwHImgVJsM//750pa1w
9DgUD4fBKOeTXSi8fQ1viTVTPti0wkhqhOG/t0gs/5xcFzMUjq9Ej1Yj5kweLBggI+zznmvfP7V3
s2ApXxl+rlhhquXGFI++GRRSCHjE3vVvXIRkeFbPka4n2yn6Ib46gOPxMoe7p7pEw+mOTbhdDFhk
XSw532BZwVzhAlm6zRytrxus4yr+kTofQe+TUUshA7D8UauHjeGqaSaLzOUsf1OrgsBDSd1a4rt0
9339SZKFXTkHJnfPciwQ44yekh5lpGjsSxnVQlKqq9ScmaCK3LyrNkgCJmPyli9oPpqu7bNJvBXn
I6Q39UKy0q4d9QmFJHpPeUL6IXOzOSlxIKS2p70G3sgqAvwfaE38PmJNdPuDNIFvWbid1ZWQRUjm
YeQsA2xVJ7R1XjZJpezRr+fduExSrjnCWGBcwz9yRzpUrkerO8hcmwN8BRNXHXAlkQ7PGMC+htJr
0DsNGqqhMF9LgxYEdKIvqq2st/Gy5ZRBSbZVqV8e+dZueO3wSp6A8SnLyI7UNSBH16hHYQqMHnZO
evTVN7MjMoifV5ms3ZQ6SAyaU013R3PRmDujqGnbxwEeUAOCRMkUuh4llMxGaItJ0GQfqc3mzHJf
/uBkz0mXOLZ2A2XmIJQx6JdCVD8/A/N8CIdYyVg7NeFXd/eC9VU2kenr+dxosLK/drYRGbcLhz31
lL7sDAtvgV57DRSzsPmv/OXZ1r5rT1rI6U3FKpwBfemAsyh7j4x4sZ8nYPyRH9ZW3TkXoh9rbEZC
qT92m/UfZXADyG/AtUO5iZjetMdzYS+RhaX/E1hUqW/kDbrAFbaDJk9GYZGfJ/9L5K5bFIpw+h9w
VlNnruHBsgm41HuvvDPx7gWKQjQq0A0URhJ4GmqStu2RU/5je5HfLIbmyAFqvDZZiQ6NY9E7vxa+
x8d1nVCieemN2rZHQtFH/p/ww+mMMu7ZJJ0zbZGqwPr9UctOeKwaWnDelriNAqROv/7emLUJY1zI
ZW+iKFwEgA23s3n9ffGY4eUy0p606P8/sruP6Ku7ehaHuMmMbLiOnaUFpkE6up+rki+F1JLsnel+
bs9iM9pC7x1NXW+AdSx34ZF3TB8Gq9m6Mg6UrJY6Gjm0c33CFwC3vLDILtcs9XhYwr9kJRTXbCUO
rbyOI+BiolFANXzXmqVdIghOb+CNZaN5VGBSWI2Q4la9ltEIMazQqNnLTlsJbLxmqQxIcGOZJSMp
XO26WSxopeKHgG+a3HfT8mDcUqItTI9wxFUklMJysiRKWxNoWguG9Yq7xrrHNfGc/kYtX5evTaq+
e4dyeBCXwe5DwmMFrTKX1x4FIvAyUTGq/bZitbNpRwU4mWV+UlJErk5kk4wfV2OJ1K2ifsg5FKpM
bl9/S4JY7Zzn8dBYnWxaRUaYmKcCb6DoTAeMeibPPlWXj7UuBXjBUC8baHqq/ZhgFZ2pBNuxpOWg
CwM51O9Hsxgd/bMMZhjmbFe2AZm3JhZZAOxJy05JbEYHFttkTxvvbEmXOZFzjr5LxjUw/WB4TzRY
NpqiWjN38DbTDBYRogMMou2+5/bB0LKe/sH83yiQI9ZybTa7yXVJyXwiPV2OXvFHCWRPLxtPNfz1
IcQdaNW34r9EZQRmESn6sz2vEPvU6ZUQEfkXRpgFxj1QYLRr8buE5o1w8rmHgRIn9I+5ddvi5MX3
ZKggJ4XqmS95dgJ9zJ2WDquFskLd4DBgtQBle3JaHYSXGmMp52VwnrHB4c2SM7huuoZPX50Q3JvJ
KvsaeLaiQocgN3AYHh+fCTv0tZxEERse12rwssMhZV6hYXkRItrM+87zLO091WmqOP93ejJXYxUs
jY/9PVuVknFhjoruhtYhg9IVKRVFQWnRYfgF41pbMo4CKzK/YqsMIrqUL0fap2OOv8+oZpQVKuPQ
2GK9paq2Ec+yoW2uHDlPtgAdMLCu4gLk1o0WRV2bk70cSD0kdZ1MjhzTMNiKceqGeDZ1LIa+a/CG
kOzvfWfUVVw/vcaGS5ZLipQ3RdmMXLmHmeMOUL7NMOBNxmNco1qchSz3Ue1axU6eGpG4422Wgedf
7pZCK/pA5zjmQnG9kBJz0wmlaVw6v6yb7aJ8xhPCPrt8vxyJ4qK8gcWw5vmfgIp1PST45R5MWNMA
YkuOWBZqopWnyXNKBVos2sEUFIJgDU0fYpJB7g/y+OGhvb3Q8va2kUot57niD6QHqrFFBQwWr4FV
kFag08bRPdB2orTUNRJoJ2Go8vDNKQKQJetf2vtizSbeGQO0QjyX1/+GtxLb58aOOpHiD64D2jqq
yW76Nv7PNn985nftg4UXnSoVqeL0kY6OU5hOYjc75BdaoxYqo6ijBIkYuGi/MrytkIXfjbYe4qmA
ZnZDO0UJlPZnrPoezlADMfl9SB38aA2UXHqXNjka0EQQauhIioLgmmj5tV+CyKVOYkG+vBqXduwH
obgnTWP8QeTb1+jpxMIvkGj71vpDQqe6r36k8FRhAK1SGKkTRWkiQzBOQS4sOlHVSL0t7jLY7BDD
Mp9yNTQC/aYUv3Y4LRqJohIRP5W9FkXl7awP7EPxZVXGz0UJQiJuQ7sUMTMBOtAqmbBJoP4o0UOR
+FdYOLp3Y2uFz+msoKWfOQ/JhBssyf5yL4g9Edxq9i5tt1ItgyEHeRAwDZCSoDTUaKwuxcZRy96U
SFs4cvq22CU1hJoAUQ5BiAURK8YiC2tHIw9uX6d+x0x9LaTIvECnIcjjyL0x1aiFP0yfHLVd3Dq2
qEiZlv7IZ4EFw44DCfs9XNmVtdbd88g6KytT//pMFBLiD4HwZSBfoh9QWaNhyPThvt6tVttITgU9
9D9OeFvmEryJwz8W0YxMDGd3njl6i7xnVQrXFgg/+QYpi3SVm/+xNyvwQE/WL0OQc6mWEK+Uq/C9
BRzrNIhhiKYahM1coRSKLBdsxJQXhKN6DyIyYzH4Eq5ZAyQGX3nYGKgpSRvuvCtQG/NENGglYl07
UdqA+PuyLUGYFWH0ee2UG9/aEH8CSLaO/mvherapSoljOlixPUOYlvDbe/sSNpafFXdvlR7sRzXD
Qb8pE5FhAl0FBypGIYhEfDSmJbCQ3Q35qI5LSThlC69YE4VnmD+en7+RrQOEIfnYVrwfx9RMpN2D
lrE7pB+YYCTVKqVLlUf5ng9utBmk0FGnER8Llv4+HPHYKw5frmWXoKwrXQriq50BHnjOd3jMZhCl
SKnJ55Ul4rm0Qo8PkAL89cYqk7XS7ASxfdr1v4k2BBB9ZfIZPv8SBWEXHak8Ad/RO3kp1G6j63Sn
O/FoSBPOtFiNIzsfVQS04LV6Cov/4zmAUWrC09JzukU0L7X0Fm6ylIlVL1z3rWxw1qht/eS9HT8Z
zhJWVssZsAeND4q7pjsTSjmF7+B+Ml4q79/74r47OaCHMzhC5gpT1AObv0/xE9mnt6bgBCrNspgJ
CDwjMbEcKH97LXTXCRDMZwgea+12GR5gAsmcGWjoG6w4cyUkJ3SBr4sbvQpZuCUFi6D1731lgeR/
4XUUPZjRt+uicHQMnrvBwfQIZ22Jjboh9hsCGkWluMwN9kH/njIDumrrnpIgXKXcWz2hSFKVmIkm
z+EM9iKFxceNAZPaHopF6Jq5UfeXLBv6RFg8ryoORy9RhOB0LaBMkN23WPc1JWw0lDNj1mHUxvkx
x0z35wSZS1lntNAWnNR2MK8lfBxpKdQWlSF2Q9K53N8YwOoWvpWiSF5ccldh6KvgAtR5G+31s98I
3DalLwbG9QIfhFUb+X7UMDRn/INlHS174WZ1dv1u0BI61x9gyZjTQn0blcIwUAxva14JHs58ac0c
S1kG5ktQ3qvHk/WMAyPuhkeS8a1TA/lELUakYxgli7vr/Gom0WDNGH7N2Si0WrpYVyXIwpzCS5Ij
yomVouTVXKqmwnlXnhpISVxSW8+EMaEj9B4cCG+PZGfCk3sHRF+t+dm3xKGaDgyqykpkYuWl9D/I
PpfKWmAmzcebeF1iDMGd9ckVNcxd7c1Uq2V5ffNrUY3O3xxGQ/MiMIMw20rn5Wls3f0vh3AOUHPp
5Nj6voCgqbl/Oq3pFhzob37B83hNjl+lkiXCV9PWGu5ZPWcAXYfAoc5feAafU7/+3cFta5iEweT5
UE97HI9T/cndwplxZbBHwDSvSkYwX+lnNMWngAA8AiNhLS2t86fnKRGI8OTbyrIKbVvLPF22XgoH
fF/cjyeUW1ayhKxW+TBa6phTTKOdMWEPAI7X4RUV8VVwssS8t9JKJUYAnGfEbXcxxUZVgDs+w5Eu
haVpPBmcFT4lhHONVJsW66hjY6EX6VnzwZTEXJrkb1N0pwA1P3NQ002zRj0GUG5BTPDCfi0d2qrv
5BOw/DN86GH0yBrB9jR4rkbj8KU/KWjRIDZiUjXjX7tMT//OwGi7nYeJdtbRjtZW/l0Durl9mK9w
mh2eCIQ/N8hyADyZongBMWXZSSvmseGltpCrG8hHi9i1SLMAjzjPytC+6ZvW+NmafPKjzC6LN6+U
xnDijZ5l3/4eLI/ArClQqZXJQETtIjD5va8urfGZPAwEhDM7ZmHGmcaZvExYMuRVzyIhnQ91f2Vf
89YBBh8gTAXj5lGU1q0pkY6BBHMwI5J0jg7yZAtmCw0jXpS0bDzgWdm4ob/+mOh+2HV3v7Z93CBX
SU3y2dQashROE9hIU+p6YK8AFnmMXWn9drhPZ/Fod6RIycPZBwok+diX4W7E7XQATzigaSzG8sgY
uO22BjLOLSEyNcy7ZzaOedZXeTMYuVbRD7y/Arymfx2QOLMVCKXcipYxwBmSbmqCizOVp6RIKXXv
BWGVRVvDxQLeTEXh430ifWU77cLJsKidDwZaKEXmdFs5Lp5YO9uHfl3K0erwJ7LJc/X/G8cw4R0z
2ioY9hHiboFZynRVppNF21p2gjt43UEYJnto7DISAFr2cRNs2tC19iwFuPjF33axJ6zHR0L0pc0x
eWJ3tlqZhKQwptqKtk+1BIs/rY2s72nTV+hDUjrUJjhL9gfRe1fj2yJRJ2QbbwA1TbxLk95776+t
kFGBdTlN3EE8rjIKGL1sEXLnFW2xc4NiEIwmzNpnFuUIX9wFzJbKahDiWcRctU6ZeKLxKbAC/Yec
67pmiijsY4eTTAAmNUgW5GD9yj9QjOAfL+QFevuyj+qljEVa16ltPbuGD4RhtHY8PBIxPlbzFjeg
zya/jcsn7x2jjs/0N6Yv9bUmaQCe2gCQF6hMM6STH3aYoxSJ+ug0eOOl7SZpWkgQDTWjfpwn1oBZ
e4OSw5YIlOxSiNoMQpy0RivxZgQwSH70RegzhPNHqURww6GjrDMqha9lkIxJTATX80q/fQMUKAaz
2Hk26ptpKscX8K++E/oAYS5qX/MVNKMiP6ppaxksQwA3gHxydySWjhWfYMwAKsEOUOeEOVd2eEHY
36rR0KfobVslKO13vZ4Dw2bbbJHaz2z7hU9Y9bY9eBppA3qAnAObGmkm50hOstP1PJF3qPfQ1FgE
QhRO7Y5j164ANNHWyn+5QZ2vlNxrDg7KDZ1jQljdzyLVXppEdibIipYuconDjuR+9H1za6lVSNzE
9oh2pOrHDPG4beeRtbEmzAs34JY3B31VtfipemMjMsrUuNz9aLggicutt/04xD5CKif7ovkv1Npk
XRApeU1CsLVirNF7IiZennLmEY6q99uoGKMyT4G+AsGMouRstt2Mca1PEyDQMeJaYEJPOP/tY5FD
o7aIDROtw5XxBp60ZEbPmkYhip/3IT9EWsA+Fbx0lr+8P/9f9FJmp8T8NVntS0S1wXcLVFKSXj2j
for+cK61CtqHvNtGfYdM+aCGPd/PBSBXwXncIv1nVWq73ggvwvd+TIiPQXsVVZGfsAlg4icYNiHS
5UR8Fy7p3la4hkHdZYKh+HcDNvJOvyhdtXyS+narsfOv+cvfPaFIEFGfpLvdS/ObpI9vKJLaVHbf
ZbsodH5aKU/wJX8OV3LExuwx2Z0G8WU1iyfBnZ+fgZeQ6Hhoh8TD1pUxTGb/kZzzeV2RtlJDJrWQ
YtwgN37WxDIiMS5XeqI18YPnaqW0yrrqtX5yB3MNio+KMT2UJZ6Jt4eYcVCttO7Fkww54TKjDOFq
CzqwYomPKahaNARRH8o2+SFTHVHHGRO26AFEnxHfacbr5AJ+WXLW6q1nWi+1Ix9gKLorgZNKUaVN
VMvCuF7blMhCpJBnEhtrkRZaBe4ZpHN2vhmyoHQt5jciZaqjh/k9cPKc+vrYv8zGnPeOvOHB1qJb
6ldH4RrykZeBUllaob8fU+BS8d5Q61VlHeM7OI/ACipynPk3ERrOHvC4WjD6+NP9omjVA35Szizd
y7NDS84IVXbxPH79EeY2uQQ1jdmnx85S8lfE0F/HyktKmXtKKeHH6R8W3/2MFudJVZHUuiDVRQlY
Vsaq5gRDKd1XfYeYx1cxDFL+7c3sd1IQqEGmGWK4wRTFMNb5O45aZ3hCpFUahIi4RrqohUOmE4vw
Rr9jCfC1a9SkEk0kpU/mlFSy+K2maybr+6oxFU0AoQPj2uMlKKTwgWtLMASfmIhBm20oDXlYM2DX
tPJa4/a8EuzlFnU/wfrLni3N0V+L7bRkxnDGp4TlUvZGyExIrWY1P4kdx96KZi7OhHDvTmZt1GMh
aLYOs6Vj7rkt8vAh3D/BrHW5k2c05ybYfeV6ohQ1m5oCydtSy7cqrtlL5Cd9jOkQdF4fLIuW/N89
DHUSRhA1Y2JBseRv1iF/qjvGoSn2JfnQ22aFhHiv7p7MRyMTCcdB5LkEqzjZhdfcGHnSTINZxmVr
DY4ty7pDObo2pKQ5DSScs1V79bKETH7hkbDrzNrjktfbfSel6u6zbnig/34uMmdVfWgjnlDFdq4A
nQWvMyPikKUl0p0SqwsHe11l820auxPlENwNpxvoxxFZKDtigu8F+alB/cgzNBTtoYhQn5LGNErC
5EFxQ44UUJ7NDkXbFvdx5mEGoG3FPWUu63XKooZ44UfW+l96pa5ZL2ZnLZw28zej/5r0xN6CZdCc
YL9lZc8kzZFZyCue47CMI1uAGAHYtNqZhWo/2frzFtNgtA8O/N68wjMQc6UidvISj8rWgmCKa7iz
M6B2ip0eFuZWyw5+ePBp3O7ZVmnULawvEiMJYFhCGIseryJ8MhQxW2hCEZntZx+Heesi4I7xBRnd
CxsUqndK1zUo/Y5Z+6sw46ufpAScUtzACmo3YQkf/sFrOuyrsQuzGt4TntLdOEptfJ8imlcjMCxX
n5iUdRcezeZ1J9nAG/bYicdV6s7n5puAhlkbsxdSgCYP2FYm0fBTqUHTx3hbDcYvusj9tfvjyc9K
mDldz5rr0PauPRfPDQuYovxLwLziexKy9r2EyzEZ8yIcd6Sad0KXoduf4CxBljQ7mIJr7J3xizOJ
x26ghiHHvbrWerhd0ObHCjnlcq8EPfHhNBRwSCekrrlNtpf0nqsE4SN3RgK/U2iZpD3XIAirosNR
fEFKPmBGJk/vwRYSqR/EucOy8Efdid3YvGmrPtl+Gixke9Xty1UEcdZrKydbFb7XYMJyTD6GZXg0
ZH2rJTxmcM7o4nNx9LbbN3lJQ2ExtZyJnNS9y1tGeCm+ln0xmpID/KDjE0AZGDe9pbJX+JZzlvcS
IDZqWi1adbGGdsIJt9loLApX5G79PGiRqjGlPe/h6D+anqaawBQfyhOnzutgcx4pxzdjZZYFdpWl
HRPZeGSvKOxUNfQXISG85SS1K9zw+way9qB+yN7SMVcSTFpc3k6MgsrOym1t8at45DrLh8wcuCRi
p3EzOAgr1U8TAvuZsqrEqq64dmUfVgbyCjDfS9bkjwRqP8gqTOAon2hrH/hyk0tmnekIVrCnoGk4
han01HpWGuGjq8yC5TAfkAi+ajqPxoQD1ZNRaOQpvJt2YL9NKPQblwDuWrqPE4qf4aLtfXKuRPpp
/wjbPmXW0W1FZyIeIA8oj33myQnkvRYhpOBqdH2GWZtt7WyPDS/4Lnz999ZrMtF//xBjgva1T68e
qRCUcz+FpqzTBUFEemeeo0/c05RSoSau72Fi66kjr7lw7BsW8Z5IqDrceyj0+7CEdwzOTI7JDBlQ
WuyHdXhIR9Lxxg4B4H5OmU+Y9k6sd1Zx4MFuKd0BG7x5Ujjyi9tY6Py1tqyOr6METSIPYduVkEu7
yL7NeTxmS9ppYV30KjkdBgHdDP6BL7ycexgm8e+6G7jullQRV+B4Q1egNNwwuGwE3TgGh8BhgHJW
hxjn6tmT3y87LU/P7SjC0VsJFJzwqR4lAmBClhn1CmivMqqkaPfBZKVbzb/oRAhNp81vi7ODAux0
UdwrXl3anHhdWwRkkAUgCYZOjGNhHZusuwggAD9Ku4aobtymRr6OhMukqF8JtsrBf0z7vrB4LZyA
XCoKC2jrimngYwITj3YiHx3//HCnToA9bPLYwLad6/bGEseqWhBSag8eILinqDzVONW2Ux9tJQfO
yGDm+SJiyA8Xk1Jqm0cj10m/7EliUTw90PpjwjNejmk5OBgsGYm73Flt2u+Xz3rgucV9fqQZ62tG
mOs1udvcesjduNC9mASdyub6AKJ+Lb0Pj3aann4P6TWCA8eyU6cVghT9Kiymh7jFh6O0qdp5EHrF
B2oyDo2u2Mze4u5r2aL1FoYkaj76P4zfNF+cvbqIuYL/onOMdgeoG0SW/Q3uuvokG3qz7hF+WP8H
BJ0yG0+HaY7/rroWNPjxJLeoouvJDwDBpr/mlAegtoaPbNGofCszT4Qi+tV7MrPUaepnlYgNgVCM
XsgP6Mb8yDpp8gajbKKrbrqi4yCQk8dtImjH+/ojqUal7RPkb4aeQHS8VCopTWy8VaRVFD7ByzNx
SwQEM8lgHxrojTzaaGPDW5U3X9bXw32526gilurg1lM3yN0YYHAsQ9Y7ueDKvGvlfvmY6VHwNsqT
IfXew9iH6s9UQXMYi7EpIJWjZJwOQfbZrTrJvjMGVSXPMOftXuaonkYoD7jf6x7NIqfOKbO1AEW6
/ltie+yV0J6gbUi+TmCpl/zARxnhVCYAFb5kyQeG4uccXiDOUCaqYw2LvmCX96e7IRzHiJne/xKe
OYRzv8u4lZjGsvJ/GDP1AmgVDEPiFPDvkqV5/i8cxFh4IBdDg5MOZTlghA4pmgy7L0/ob7Ks01dF
P9pXOZUA51NkMQ48JvXVcT26h35UyQ2n0m/WuV2qj2p6O2TV8n9nduHkrF+MRzm/qU2EfhS5awO5
b0Y0gqTf80YCL1fVIQHcsZ/pSgxjXDCxSDxVOuYxF4P4q0Izp8ZE1FZl807o0d7ivNfPy7U3dCic
9V0dGzy0+Q8kNVt6D1SsGw3cmsnOTHrRPYwxuZY4XQBsHGAMUeLbZEByWQTs9sA1WslMdLJy+zzJ
iUu1FCgUgrrDbliLH686RWU0VIwhKc1RHp0WBUaHzpkHcw6zayTCYiyRx/SynSTWsUzPRgiZqFmC
Q4rAGnSOW89Z4/auo8XUbqQ53oPN+Nx9DjPevnQ1JXtkTJtP3ctEGKaQAb+5jetIU8nEUQ/eaybX
jxsZ3Q2e89YpkeJCASC2Ljcbkgu3W8YiwvJsqyjPPHBSJqE/RdqKOdw4Zg+CqYGFHoE21K1+bppk
nY34vl9Lc/H+AcntNp2tzdgue6SRK1Po80oKEhWzcJXCHkyBWhXI6xFcF/CMNpOKrvwsSx9FAfXw
4DFD6C8EbbpnX/seT/DeSivN0NGGeSAesQkOj/itHeYrxj88OY4549aau1l1QXHHd3y3OqmtIHTj
X335zOtQWnr/+IJo6S8nCSSLsPQiaSUHYffQkUPX6Nfdb0PP1PxwGsglTGEjRCsjwTmE7c1vhPsD
WrwHNDdEjaTi/np/P1+Cym6zCD0iITAdGCwHnBx1BRfd3MI9lRW6w5K1ml6grdM9X56dsAqeZBXV
jBzDpfJIf3dchJ/ocq8HQDM8I5AXuSmO3MY7Gw6Jlbr+VtqtAsH8FYVRvAqpyoGPOSX7Af4mhcsM
JENuid5m/25q+Yjjqog0ZmZyXlB1oAdUlUuqTHNE04GyVUeMoefA4jRnezYrSJZDZr9jfD9yPFkY
lk+QscLcCxJZ+ijbZmecivWnQWmJ3h+dvHQlQN47ZlANU+5+i2HmO46mf0lUS2j+OQmOurrNP7sD
P/7swxt+mnNXYNk54ROzA8NDKAWkDPECBcm2mHEl7Ix6/Jin48Q/3+61FQLHrBqLnr6rxeAsVdNz
ud11mItJ4XaRtp7GQIgBUdl/SyG8Jw2z+hhOS1cNmryHGymlKnc3bSgOV3EKTKZpFiocucP/s7kY
mmyMHlUCg9XIqEFGekZyayLFP4zEUTWFgMwqPsTz8CLD1TZ9/2nDdRbT4XtJ69nodN2OwUGDpdZ0
1plLHOF3P1ttMbxeo++ubKpYqtRpXl4Z3kCAxsO+Q5SgU/yFQ4wS8JxTziTLSTaf1lgyjZz5lcKE
i6deZZN2MT37Qx0QKTkO8c91AZLQJdUaOcmFd7J7LEALjIdojCK01M9RRCH2SIdDGn53hg4tSDbl
rgI4YUBqMXrm5/1rFLLJNlVu8FKwoy6vl8C89fJJvW9z/0hZnwjzqIZkDcHld75XMRZp6b4ovUZp
PezND6rycaHlu/rXndHs73I+kkGBlPv9FbGMO+yS/Yz0FCQAATic2H0I4KukZnKkX/uwT+/9Kh2J
hgdL89MDx0F9yiSOzUDn5+wAj/fIIqFUYbhwtJqMomEDtoGx7raFKvZdpu2DT3MM0KmZNi7Yl4xN
bDWsAPtrEv+CwVcE/QW1+X5VQ2Mdtmq8B69ijOzf193y0TXXLRulCyijC/iS/MWcK4yLxqTiVD7q
u694TUFzZQ+hYtv7xhrlCFLbe3vlmxAJe40gTxEo6VEjhYyoNUCuSr9CSfvlC+WLSJEsTRhL1oVr
L2pkYZExhD4xMjOCt1lNSMsUjVWm5P7SzRJvlydJNRjjoL9c1mCcX4zMqc6DSDabOPtlnfk+/loa
16jzslJMPxqJNs4GcQeBj1rsfx5hcE3iSIzaKhG7Btug4h4GTHOW25rLQZdgMmZxbTVMslQuNf1v
c3SAjsugKq0BfcjKEoSn13a/jhmTD3o+TvABWovprGRbiUmyx1wRA8hvpEsOLrGG5twPS5IdJa+V
/jEJxAU/oIV8RoYgCGI1Kemf8/2muzC35lpap8DDQHr7oLSZ9bDwXVQEuJkHie77+afMqhjoFVbh
mwM5CWssR+El+llBxWsI0zfUyuko8gBnP9N+Zn0myq31fPiM97blseitayqnaKU2pGETbmAfnwZA
u1TM1/uGFhgSygD29jolQbYRTb/MKgN8P+TQ155kpPnPi9kQFDGkLxdT7FeTmG28cQrnDPaftX2f
r3coGZvr1CUVqeDcYKhB25N4U1bs1kagp4QY4DqbTqvaY98rDf5jRCYfNoxRKelc9ZrxttTVv3gd
w0qlrOsIcKAtbNXnZGEdsCyQqB7oPiUrV6ZVeSAh+COq77Lv8CciF+KObaqA/gHaGG09STsBCAIe
WKZQhHGhqpGbZN16wAyvhtHaWdo0Gv9tjtBvScmfxGj/B8x1ywT8WDXk3J3AEzIPFr6nQF5t4JgN
w89TCwjkJ5MP9kQqDhV8JIHe8jt3l6A+nBL376rAvSUpXN1cVPNc3D4uUS7HLOzymBRFBwn1VknM
Gwy1dCQZGanjXPSSgChROaam2uCHOjKabWcDsU00NyxPot3Ces4VMk0PcvhX9+dZboghlsY6q2x5
QDm7b/KCUkj/x7RuVSPkB3nEnEnMfceP5eukPkUpdX3TvU3AOECkuIcK0ZTNiT8mDes1D9xgWgqo
r1AlbUTgxTuntwQHi9c6k2fDdZOg7DKdwsHybkfUI1dH/VJv9hYogEQCwyEruG0bShdV4gQ9klsx
4AVQ6sulIKg4WYDhvaS+da86M7wpKNS7V+pt4XH+eNTeie6+Y7jr4L79FuZ8TcBDY059Ajbtxek+
SrJfGXWCCh/VjDQ5cdUEkzlmIow6NXGBcgNyeke4sNGR2SzSyI+02msdGRWzh+gAoVByI1tG70BL
RpZJs7E/DBDyEU6ZYXk5uJZFodRu/2SCDCWWPnKPM7oq4mKnF/SJnp66/7AMXLdiN2uZz4Kd1dj7
Gs3Zbvs9TmmM2ZfT6D8iTTGOHv9Gma5Tq4YnbFHrZADPXo6mBqhyaG8D6+m7ZoIXk4EN5yMUBsVI
g/zi/DaYsP/RVT/DuFivct+fEwg4q8YqUt9q6nx3CQG0zWgqNimdWZ6Q2ngh1GAQU38dm0gEQiuu
c6hHp/iDOjb4+GWtDeAiEFmpLNRVnUe2khe6f0rxgPp6pvVgUIrWVfealaArkLOJMDoQOAPoUw+6
wMo3OU31B44LyUmKu0gfHFhxgEdq+/5tpMjYIzAgoCWvRxt7mNAGwINZE0pudQJ8rCYukkaUwH3S
PvosyhFaeEc7jqkik1lRTnVjMPRguchZ2imEKm86L7dXK+o6yVVzia898BIIraoly9R1GprkEV/4
RRNvFoBwXw0oS4OZhDGMM4YYsZQJARITCCE3GvQXBHRvusOBx405GaPmyOFzwIH0oaf1r+hC+WCS
V5vKkk6ybm00j9ltiOaETSDwNX2Xi6NrkpNBccYEIz73BE+LA4nLfdlKLHdYmyMoDjmGDp8abMMU
P+hUmE140cXzgF3mVMKDVv56OujOTG8zkbkdzxt5bYsplwVNd4ltPt0LhJdvwRzUfyMDOEGsQ4oK
/XfoEAaRi2Y1y6UaZZF5+JAbQzlhbsIzL06IZtkbUJVkQ1iTNeP2vTGBum91CM4G5KfZ0xZjgxur
xiV9Id4p16rW+0LDU2EeTr3VdrnvYn8sDKV3i5lYdd+3Z+xOR1DUEsceNOkgW9MUefw73FYY2nVU
esOGc5Dmh8M6BsyBJeuxTgXc0Fd0XvKsnYPhDUz31knWs5rGZFhC+irCelZIPNHPWRral+nwEcfV
nMYYIlmQIP/Mg/jqRRStb1HQUDDMuE0pG6nBCMK2NngLDN0VtNG/A9Pek+UZl+TY/DaCnxZdfa2M
sey6lIx6jfXdmZQi4k/fT69W8poVXBUeRRObqxdCwb9aErhEtPsOr1dA0Lc9kXmrbiKqwfP7YZ7x
+xtqXebxhJ3n74Z2/f+CCn71xpbymnmViJuvGCKTocpBDDC+f8PwjlNeMJL2+0YqOE0kB8l7IdSU
15LwUgho+66Pn8IU69I9Jqd/9OMQpbMK3P6E45KaImzZmOtJpfev92KiVSGmH7Hy+8QVFpYDwXp/
kxGJc3AUuvx0wB9DyxH0JsWWogdVLmLyvNU6eZtl3BKvkhQ7FinE3D04Kqdl2I44oEtiCri099Ey
VrAISO0qQG8M0h66ru8CSOd5Cvh8U6WBSOzg3hkz6Pl17qW/FH7OA7c7Fg7SynRl/iYuRT/0uzZC
Qaurtd1eEfATo3ukWC8Uj/RnyVSicgu7l8hQh9CQL3N+v8wRbyr2FSu6ps1KAiuLshP1+CBjH8IR
JCtnKKKqLt/F1Ymqfrktyh9fo2jJzLXvjpYMaHr5CEAQ7s/Z6lu1JeM987+QheXzY3ZSaJv/HHNY
U8y51lQcB0pxryK9xDVCzpF/cMKYiVOCWms1aj8wBHgGGC0EESy0E5TNaLGjb6OqnzuNVSUnsU+a
YWKRYlAAizB+7Kljvbi9vnLKgPRF5YeKnkEYjdMMcebOskmO4AnbnSt4dE5GZxSeg7oNVftbYsYV
YiiyTNfkJrOUYcH3un4VwftU0queUMy0h6e6AxREhRmN4GxBIIiKlFmXIkPh9gfDvYvudgQiEsIk
7NHyIc/XfGnWQuP/wa5AdzcMvpc8pIOIqqMiiwhe8uns9tEmQFrmUWLh39yBRIb4KNY0gRTHMljd
t/x2QMoIuVVuj3T/us/C/yRTgheG0Xahsm3G81jVgaxQIJKWeHQyZMc8bmWVVBc1FLaZYaEQJxeq
FDs7OOcc7KzlEtgj78PaVpuWANE6+1EkocbJKcpc1cnH8O2ht/pxFgJdZ7K1n85XGoTjPZdFJnWI
137q+QQ74mdmR3mg8AA/aK0gsbHmkrfILgaDreqLw85sre9FsZxzowaWnUtqStd9vbHABT13dqms
CR3E1S32VETY36xqSLPWX2ELASIAJNVFi/WD2HOADzKV388HSTyo9Gs/gU/6pCBjXRtgCQE1u4Fn
l7vSpAzhaNt4N85Fn933IAMb4Ahz+LCMxz4zZn+2ZNu8+NNmXFAcEfFJ3isMkMsgtKLwc+v9229H
eaU0gAQ5zy3tlEQb/ZUNZof7DNh0LhNUmvu+QQ2uuo0jlEUFU3GDpP4oy8h1DUqgDA0YMUethnuz
35h5KPVCZZ8H5oJup2tUf9rNpU4mRZw38pzE47fiLZE7g0FMb9ManKTAVsJa52oIFSSAMQJ+SHz5
Jsnc/xQn8hdaOAXm4NWjDFLHZOtvL+k2frjWiOuFpW99vjK8ZCYue9gTa6A+sxZwCKTKn4obj6HF
6pK5VkL9AKkpSoISXfT4EtqRReq9HXDw7atc6ehIeVFQ7QezmtQHn/J65BNUM6dskYyyL8f7W0zc
uXdg2z0Hdf8y+2UUBQ8E/sVfCxbOWeP2Fq+ZFCAtxk0vyG2LPJX/cgXpDLn6X22lVEJQ1IHcsPiT
6zyvZpszJYE7Jqg+RdcI3vOk2UGfIe9WgMQ03LHA4IxAyqxByPFalIeYLjY2LdxURCm8yeQrwz79
MJNHgTNuyZ5e0JCjqQ5fm0cL/jIQuVYhBazHYQLNrdJBZCAh9m7YUBauoClbL1tlU0tMBSJ8PL9M
CY4pKabReuJrxzXmW11JM40OKAdVie1k8otCVLnI3PkADuTmaQVgzMz8ljR74rK3oMWz8bj7T7xe
IpfEkglMfRbmTmp2JybC//4okgKZWilnG+AmrCZX5NQImxYeqrXq241guXsH1n2X2rn2DEK0AsRG
6WdTdBAF3nPioOSXcBwv+Ys3I7idSXq0E1dIn1z/pwVRJu6wuFyFTUO+hU5lRq7A0+vLtVSs3PRd
MGRX1rgmbDlDn5ZNEAXSG9OjQdExiPe5HAVipkkBkBrG3fifP0l07LQq88ljbsbe/FBTsh7kG+yQ
70zWGSBOfosLOsQINKOJcMs2L1C7v0iT6QkbDOTprPs+Ljn5LSG1QsEbwFxzJlKFy/VUeBR7Gssy
Di86MbZ/xq+jVrZBZ0jJuBwPueedmbCAS565+cCZXzpSluw1mZw81JKXmN/HKwAG0s6YK/QK0zvp
AaXVxjnpuZdt5qjtJkUYd8oReS1nuVmGIUTL1tAwcge3kwR8sgzElqsaWCHz4ApoQChT3wFe7Uhv
dSxT9GuhDXr9pmHpX5V+PrI4yT3ANiQvYT9laRNBl7qeFttzT0OQYWmt4Wu3cqtOkVnYxBsWC/4B
1hoAVN8f53EMtUOCMBtr7ndw8k+Pw9G8LberMdpT8vhpwqAlTMgZb2IjNseujIf1lN5AqoqeyNyk
WiwoU3caDxivj+wQfxLLPA6/SQ8P4SSAp4DkMRdfBbGmVdP4JXKZqZjI5QoZAVuBW/EeIn15LQMf
LMrcEefGCjRFN4VNBhy0Fl7i9PoyXYZcVdjwMEiQS6od+5Z1jgRP38xM6ADPex584RA3R2Diq6VK
3WPjOXcq8vl5UxrG8LOdZtWPQsrPVgFbqhzqX+NabojUVKHmIfERwiTMmOvqKUSk8HH7VpvW/QdH
rg4dV9J6rVvafADcnxRiHGgxkxQLi9Qr+YPW7xsM9BSEgQ9gcJc9+fRK4UpnALoMDKeSHPAzXH01
KaLq0cu/h1d0i7Lq4ga1664XY9U6yA/ubd2859VXMW3T1/PfgLA1VqqiGrzyGR0VMr7nLZQZKvN6
BYcWkNtnT+zVjMc2YEV1I6vT3dsta0urp50Tsg95M2htiQny8IYBEv7XCiqmxyXUVo7ZHH0520qI
Q0MJR4f3+fAV5i773iy/txy+9TlrRnBJVdTICU37UTBR1AEhCOZ9kmz96nlRrHUJvhTPt/yCC8zO
PYxj9CxpDasyVUNUI6d2HlZJmLPwEkLfC5WLxexbaIjKqPFHsnup5f2040Y4aXsr/ECj9wxZH1uq
OYUJoRx6Xa/pJ2gGCk4UZnnvQN6jW1Hy+h0GU01Xi/RTz+0YkzBdK0DFyRqD0p9MHWacu9JZhiH6
oAmYABz12MhHoJkA+MNmuy7DzUZnuTCUpeQK8SU7XbsvfWkM9qgT46dWULmdEBlFdLDFPLtgvAj1
0gzKHQ1mZMR0PN2SfDQbov0gEjLiERfhTqoiTzl36XMWiatziLEGnSsLJ28jBRLzIcLYpsxp9aFA
WaebNRKf+MXaDJiAOhX3D1mE5+nDDchGs/9opAAe/jG9JgVOhPvkI4CqZ7fPE6cAW/LDMRZcaG3S
YZD9swP32oUZDgToK39BIj0T3Z/mU2VyuGC3P5Bs76R7o+HA923OeP8BTXbIx7GroDtZlvM7bJqa
w1OjEvIF0BtbQ1Aqu55Dq3sugT8ZZpsviR8QZ+XG9TKNxqzzVwvCcviMGlLWnHoKXHPOH3LRdHc8
b/BskEKkF9nOo4LTJ30B1ZjXJeKfZsoreWm3Qs1g2EreCKS1tEdhshNdRrQG6aWa8WmH8czBzo7d
FHFkaIH3WEY7wMEMFmt28LOF4m81Gg+gaMTas2aY+UOlC0Pe1j9T9ZwXALhGM0tIwe3/qRvpjnDA
ps69D+lrYORs9RF1SXOcOCmRvw2g+OFXPwV8BWkcePbssr5940XHkBGuUhagA+JULnJ1Y/4dMCTG
pex6K+7kbcmZZFxD829zIFUPSvtMB8+cSYgFSypzKh0Q42C/z68FTm8QNf71LfsSl9cqlaEO+JiO
rjtIUglOGa9wAgvOsMlOPViNLrmHSEyJI7RuADM3JUFUEfgdWZV4oEyH9N10TAE4InXDR55X3/L/
ic3FiwhOJ81DWvY1LgmjTaz4dxnL+SmgCkmUnPvXV+W9Zve+Bgxust0pLxBA1tL0+/CyysyVWGSS
Zh6+c5Jfln++qYOYiKLwZdnrwtExwSTWxDGABO5odprQyJMsDkRjjAHQE3YlpoMyEYuShSBBL670
JJ1eyqaAmdHqDJgzEOFrTc/S0jul+5MoarVndnllNt/bbR/0fD81K7zfyUzILyDJOyCHXGDVMj5z
6Xom5NFGzS98I753SYQAIdbxU0eW4Tsw7bg6MGW4YFjP7EVihhKJvol+wVgFb40KXYMbwK9cdZMa
PozxoOMdB/mmBGP+KgttqNQTH7VctUvCGufJMs++UjU3EDKr2SIeGgPg8lWxWkiQ8/gGwnacvsk2
hPT0NfG8z7j3wg/w8PBJffzJYvPLY+99XbdnT0JUBZlCl5xwByx3Vn1/z++wDvAEgeTl/EpkBT05
J0AiUAe4CVbg4q07pz+OIelJ7Pnvb48N49LLEkENBwLcAZvpJLSZQ48KKBIxza7oGSG3wO1sK4Me
wYGwn/EEzwzf9lRDwKSZWiLdBqr69gWmwu3H6b1Ue4oZ3hQzQ6+6IxTDS2NTvuFl6twNq/hVED4Y
NEjYaVpTfjv7UNCC0NWRfngXdplZLaWb6qRa9qE4cSLcm9psjJojX2lsP/8221q/5lCGLw7wiZFR
oJAaHBAC4IHUK1o2U+Y7xEED7iFvdCuFsNShL0c3Eiw9iZft0FwlV1jM8H07TAwh22c0m9bZjRfE
YsXV1IRGXHe/H5nq47gy41mpktFaX4odTYRyaTAOqVT/7W+7XlU1LVEuLuGzqX7o1Jhbi6bCn1tS
PCwiLXouIaYwb0UdFVuQQKASbLHQQ5AV/wV41tu3w93q4KTiNfK6Fb3qaf9mS8BtL7s0n7IuxkbT
eH1Z6iNbi7Wn51WZ8o6Cv50Os27w/vluKK2/cHBVxP6mB0joEzVnexdOXqwhDqj915FaUDbQR8Fs
IuYaZ7KLHI56Gioh6NoPZrmxPhJe67C/ntHU2/KZWxk9ZvM5Zy3ZOTBpOWXJpBz5pJR+tevwqV8m
n8Ufj/9shErXRWzlvLVRLwglaD+BgPlq1vKgpF+Cv6LyEkB1jIn9nARCZwRhZlnVueY/Ek+znPYa
xvuQxzkFk+HEq8dynE7yv2TRAEaZth28K45zgnHZM576PS2gFP7Db5xhHOwf3Qw3g6yHErLzyGNj
4GDnI4pEyPYdIUVRgisguX9zSB+CIkQmcdd35nQHTh64zDtoSlwG9UWdaayPhs4vwP8WdSKAyRM5
Qiby3vEQ/qe+UZRWtt5LqpugIv+H/RMHhwXiO2DpZ8Woi7SX0ZeUlg6vrosW8bwtOvqI/mbIq8tP
HWG87ALEo5SCdR77G2OG3T8eK5UiqpS9hkpAtYGkeVOn9910pMQaQVlrzb2CRmcMdb7aeaNRlANJ
fG6m5/96NOYgSDmrTKgt717AWPd85rfNPNoXqdSXhehI8Oky5Pjras1068tXuKoTyjco2rWqNzlg
I/ebNpHczrQYlqtA59bDyB03PFIn7O7JdKCTgFC6CrVKUureLFL8YD/6qH8A0ZpYyu4VPpBL1V70
XTjJaOk+6ZChXtyNmtbkqnlnbH0pNnArpq08qBgZdJXf25B+/G80uV1B0P9s26Xs7VJ+8T/tkE/Z
1Uwuc4DlcnEt6AqYVu55ffE62c1CzMGX9y9d8tJSmiRARI5rnAX79/Aylq86zrJFeQbS7j86E4N1
g2oYyVEMtcdtS38xObjrdRG3s3+6y7h5A7EzwQLL5j7S86p/ZaFdnB2nLWAv1vqMtnjetFCi1OEH
P7HIjeZN0pQ0EK31eDoNNbbSF3DAdVfa0+Hj9+myvcz6lERZIeSIVFWMyBrxXq9bg7O31W5Dp4vZ
rutyIa/uOdfcHFCIQnBt28gGyaa0rg9SOEgF8hpdO01t6peR4+e0rsAqKSrBM0KMQt9oCLcCurhP
IPMZvYEBoIEbY9m29bky5WiEtRdQD0W1LJXkpPGUqxlfbQEPdQtQOqP4zRrsr1DGkBjdJHK8hNJM
iXDfxOstNknTj4kkGojH/VtdTvOXTFNFo5b6WmEf0zw5mKbLX1QZKAGvl/VKTBUQ5gSed4fqwoQc
hRVnwutA4hRWQ9cat9ZEhb01t/amPNUmqAkYavVh2xXVibJzEN1TnFxcYksI/QjSp1bVv9az8KdV
GFwk0su+b2GK6dToyaQFwPyrpLb9NQ9rXsLtdRPdtxqsClNMZvoM5tgqRwkBU/gmlvaqeRhLscGE
5VJe5SwbCKFQB+A3d06FjgeSaMVfZi8y7XgPY1Ov7ARDsl5Q7W7WnA+hQRV6wV1gQ3x9nzxfJPoS
1b74R+UViRvWyHfedqtYTwDT1Dd7YabDt/PoyVHjp6GvkFYvAWLWPl48DLBSRCP7tCchDpykDXRy
xIFs7iCYdoodoszcxJ5gkoaoA4UBEg0yrQLQ1fStzvXjTDUPi1ic6O5VhRZ3Wgsn4jODGjJpMLrf
ACR+8FU2I2x1k7IL1lAy1EcTBZpNvcadmGpQwkZuifUYmIJCJ11on1X7Xb/CJMXnwvd6XX5JZMtR
24SqlGYps65MQOBHkxFjtYAPHcQwCl7rev/LcokwBL3Kf4yg+Q0ZKLTfJrsQGq4HbF8jjFUyHxXx
9+FdvY/obUFLJ+M15Da6HuaUobGcxq5yUjZIO+TTeRM1fi20RiKcRZcZzWo2IHIYYxm6G3IhnpD2
VWpdJPxPf1LsxrrGKRt8LEHZLyYbuPFbIM1/l8MLPUqc4cX60yJmCCnbpDz0Hmy76GyH7biy4Qew
oJnDoykyLS4ifCVxf+NGApeXXzhWDicPIebAn+C+tf2DSI+4QQ0HK+m2ztYe3tbE3mSEoVBPHFlR
gUWvFLfRA4X7lnvtH9+iki9LQ7kuQxk5I41puaBlJjmgxWklERkn35ZsJsaITtWAEZ7/RNejhiuJ
zl8ePYGpUQw2kk0nRZWsds274k6GkEJN912U2A5kwEK767NtpByQhmsn7Wr05EVWKY8qP59euJQ5
W+2TMWbHNTaoAHckm5U0CPZqxp4ZNVldZ0FMEiCU+S6DGqivgcCk/UpqNabFCUEtpM02UHCwx44b
ujvSTLmQ10EZWyeBoaqD2ht7yftrBFW/Je4Z2sSWxkVQOyPQtv/R/ijA+VJjp1lZSz3kj3PdwyHa
4R/OA4f22Lu0HLVXngdDOOkH4Uxidz8TjiipxJsgOekfwaIbb80sWoFRsrU6iaFiu04AapwGgqWt
uxsK+mK5K5nmcUCJN1jmB639bv+jTIfrS+Us2oPHaxBc+ZvFQe75EAjQksrjd8uwzTamUIXFbHbD
7OHp9YU1sWDoR/QyQnqJeYZvjzM9fv6mjPTCbH1mudxZYBaPm7kQnwaaUufuiowUtHUKE2KhuL7E
tt9MPz4sBn8OUvyGj2o9FkIhCI6KmZPB2Z/5Pa5qkR81+y5toDDqA0U4V7cYY4jJbQT5XjjxrhA2
dWxBcQQzoMw0o+fNlaI9WxfbhjBZpNONDvJkVKxnhDato0FVKAF5W/akdHqL3ozYVE4m99fNUoqp
OqFkjhM9fQ1ko+hw9Wj0hStDD2cTkxhTqzBydZkWGqui+aY6oAvmffyHdfURbcRLCRG3CwcJXPv9
wk6GNdOOzMMDvzXES/bu0LJ8ZFOkC+B9MsbR+Xr4rTOfXtM55HrVmUbvbQ0MD1mFQ2APWPb1XrtB
M/NasHlJjpApcR5+WodJLRKmwvTdZTxj7ovm2CVvvpNCp/gBKYjUE0M8F8Yrj9ED58ZALPdICt2N
OCQ96tjQXOCQ/vWh8P/6fGFiCYLo0m4Cr7KTL0ARU1Su6WC9oALBi5RckoMelhy7oz+qiNXkoIQP
QTUFBH7hFCaPYL8UoEmwXwJhqHvw6NdaqXcj0e8vU6saILX6b8zEbRXAwyhOvOP4GBu/KLO0tMtw
z/YF26bv6XxCcOd/z3BKSpQRsWtPUDQhG1qn0i1gR/F15RNv1hY0M6BNnyQLc5O4/p/phmnSvuRv
mUE8FSLuidQADnBWZss5ZXDBAEZzYKluMYZyJmFGrNYusuim9PQXzS3MjJva4qiztW8PdtM2stmL
e6ckrlP7MFPLFzVCNbsb6o73zeWEIvEIgcJamwXmgQx7pjE99DRQnd2Gxp+GM64E+mtYD/SvnAJq
Y4xWu8RDBZgXs8MiRi9eK1vU3iNQyfxNbTrgcuTuOUuD98brt2dLG1AsE8f7gYhuLzlFbC+if1lB
BYP7armBJrQmTlX/5ZK9UpSkxA24tk/4/SBKRhOgvsfKzbivedMdJyJFpMPny9uwFNHA5/9WWb+H
ErWR+JB1GeTNdtZvUACOFMQ0ea2YYovNekKCNz36lqyNnGk25JuzkyiD2nlAre7yehPiYaiYEOvK
aOYwXLD8STlZVCkQBspnxJtEwUCCwGQkwRDnFmrhtk+VdqdTBI3ikKWw5ucFl0AGS4MlRozrAdpG
3wH8cXN44r+tKQtO6y1bLVgnAKXcn9KQVO3StHvj6C1cSMqdFyNSQ9y+dBJmFwihWicCNGuqHyiH
sQ+G325Ukwcadh24pOzauxZD4uIdj4wwARNmGDAZAy9JmdjkVYWYCAvfUeDBJGqUpLR5Wu98moYM
1dIh7Go8HCRaKFyA8kya0fA3/Nt9hqQt9RPcxez8UEfJN317SIDUMGkP9KgcRgPZtjN35elRzdBZ
uOCE/90OnrMytx/qSiAacypfMdSZHv1T24cx8EIpSnm5YNQQBPhQZQ4LklgQeAILfjXCPPpi0OTu
O+UyELCOhj+bH6dY7ACHEK5iOQMg+iYD05MAF7SKzAy1fbciFP68/74vZIS5Vq5RHXa+SoqD15mu
lqgCoqekCqOqpcEs68lY78uigW6hrHiT7RgpETDvb98YtA7f7yinFavYcyzJm9Ak3x7GvywuZ/Yn
7XyR+CxTJhcJG5TZngbc+bxTLJFWTzj/iHW63u1jWSsz8wO7XEjaLZok58k4cQPriDaSbWHLrAKw
pJwQvbuFe9fhJ5uP3MiVH3r4Ea0BPr4GJvy0Tfc/nOy2pfJuqj2xjqDpHsPEr2yybjtGcQT0JaIb
xvO6ZsR/wqFAVCKwTriyg4uF1i0kkCgTdqBhBHkVL6aWUy/RWIkuRcGncP+cChinduWRIW6YH+XH
QRttwFdVAPb1ULfo9LZ4op/yS9o4v8v8w3J3t3JBw0lFqsPnNcCVmTPq7HTmD//QvpZj+o2jsJMk
//1Pln328vHKG6716UKLCcTnAHkNdSCTm2K2qLUhYxG+ml9aRsvCUPxTXfWhdwetqF30/3bEOeNC
K5JHfyJ/nAFJeMcOn5MD/J6Ddl8b94fCmTShYSoqs7CbCm505oUk84YbjMgg60Bk0gwG6YoFohFK
yqNWWS4CeiuApqeqkAfoUlaKOcBDhoizs0SpeDxcdGz4uLTmhlvpTn/NloVVh7I0KftZKLc3QWDn
4yZHl3TU/xVOXll65+Nokl1iTej+p7SVXF/eFByedJEGz/2zJyAz1Gn1XMn2UV9CQRsRpq4hBb1j
ntO8/MuRKHl626TGQNK2JwfHNN+qqck6u5XH70w0PaHx2ZxunFEN3qPskXTu7zwyqb9UObNoih7B
XWd5AHSSSpwCEUnXGXqOpTsueDa3z/0MXP9NRTh4Awtc0XQmlhdnlIDb0g6owD32FX5xCUgza9Kz
JXsjdo00yi6m0S5vuA/sXBuwHr/zpYVV/SnrAOByCb0UQs1uzzVJjADecPSgGW/bvQW33/IM4/1Q
fpgdTwFq0GOChWdC8RUtW/mF+ReOI0AzjJ6XZT5RZpW6TAHBTHQfNG9F2alNDWvtIuU3muIOO6Ur
74YVH21MkzbHksvSAGX4Fqauto84Omn6SujrFjIJ7IprAJ/Wy+V5r6p6E0sgf1nLXQ+Nky99hvjR
UlNvzUC/MBf/zxdr/+MHuTLVcuIWrpEa/kqXgm95op6twj86hlZ76COw9V33IJA5H8Dn7ZAQbE3M
h5+STMkuprpkAovaSC7DLtfVs3Qa8wKX8QMHYP6xHVP4zAuVM4//MVKZI+xohFEOvOYZAmH98gS7
EmJGZWSgBj74+T9znq2G4mZovZNdfAIgWQq3j/otNHz3ph+M0ENt9sy7M+/p49oTyk/n7suLEL1M
pUjccFjx4uW/g3hkXbUrwTBJjwhxw+5WvfKZa6aalH5c1K6HnexTEfuegLTn9urGeF2qz//mnQjx
EjCNd03a3uquvIO9earRgVtBH6dKMS8NhSXHDbFcE2WnXgiRoL9OJ/Gha+NJ9V2n4clvSBx9oaiI
A77g6GK03NalChbaDoclsanSKrIBu7/GcDJOEDnVRYyJiXU+KQbwC5KfMYsOQkMxH02bAylLVSt+
LuG7c/Q26M+0c7yDbxIHreyntLdocWpnDKv+Gjj301xZp5GzxStUYs/RlN2AgTqZ8+PaiKXG3a3i
ytbGpC8XVXnV2m4X8v0YFw3QLPvCjqdkO/4rvLfglYcW3AvoNTSsu+nBASCkYAfjsNTzvtxhgmzQ
5/D7IJOL2X6v7VoLaKGe74x8Prpf7zKrfwlQ3EKvojes8A36J8kjLb9Ef0oqOnK48hteY7JAEc6R
dIcKGmOzs+weYx0JtY6//rD+0V3z8cLgc2E2g9mmBJz/roKpJBikt9jmUkOwoNBKXi7MTjQ9Tsoq
rujnWNtRO6MNrqpxgNxdxGWzRkEZJ070RpuCCyqUZ8IqFTs/gAZAHhePlG/IXPsB658BouDvWq7U
qk8RBDzlDydKFKVeXGpfm1awiRtnsRHgV2LWG8aQYH9tI6OYY3ZDEKNgBTH3GCHQ8aCezn9vTcUd
FU2UWFegknBTrGp7GtFSGwTdcFsPt9N8wbtTrfaqbISYn/V2yeBon/DoZaHYJRkcsHAg62KGbQal
8wuHnavVgePQpJIRZD4Itfy1tspEc551NgwX45zP2z29/uH256/bIEh6/H2i52WkbAedly8wVJ8C
A1WJMAvzaXx8Z3Nfc0QmNCfzLw0CNCbcIQsINdFebCSzuM2eNW7mjkcCv39Mktk5MJbC3qtwjsqn
Sv0TqU6ONijFHtHoiB/biZESMIRrZLwzL3UKT0Oe1CI5wC2ik+UuIKUik0bGozgzG/v+rvNcgFA5
QyOnQP2uvy1MK1kGr563QtBW/XAjQhy3HKoujaF4njORdapTB4KDwdJBvUhpp/xZK+/dGAHthFNJ
CjL+nEmXkkeS6K0F1dc3js8+SaXMe+lCPFKIQDewig3OGI1mh4Ng33hTW5Dfr9fGEQZnSNtDXYGc
DQqKrt+JuhV5sYXpM0Z8OUs/4Fwp/xmbKtj9X3QLOnVYlX6WqH9TCabZROyFQZT4cUu1F01cCYLi
LdWNY8nzJoEawFuqlZx3ru4aOTvhCMKwtbXGnjYU/HPdCAApBxDtLs/eS8adidC7twmRx7ZwZny9
Qz7M/Kbp7MDGsxkrGhbQ17EXT7RDYGSM5z4s9nlWpRHrJvxYWTggKGOUEdv/e6FmST7kAhI3XwsU
lZQeA//9xWJsPlmWhuDt1oUmiTawMqq3V0goU8iGkoNicXLuG76wdp5tLgvpyUPhbRVy57nlHXYr
IMKatNKXCTQ1JjLxTTHgub3xwQnDzlNDYH6Dv424fBHYONyDGoz0cvrpnEYvEkcOj7k0TBCcmiLa
++QO/5RHcPUx9OcYaCv6OYiE/pC/4FpNkTps686MbSckLQcFQpS1U/1igYGE/6xVIqjkyB/ZwQy5
FaOYZuHekCaDRhL24GRz+i1AUYmEtpD0QSNxoiuZ0ssnJswJ8w+GQ39+PAH3WHtDAzIPJPGgNIf1
8Jk4Q8U4VKRX2w48HoiWjP/vZS1nMrOEXX+01yxovMuXtarlXVkOVnoDXWrR5CQ/StTcudozL3XN
ekWOuyRvxLVuAjYjk7G8ay9zrb00baOJRFXQ3/6nIGgGLAoIsGh0QTII9Nkhq2bLfoPfk/S5CSwe
E32yana8LvPTNbrDEVKB0euZnDfOiGhHrcL3x3sPD+CdZCQgsDNduciLWBl49DrPDZbyOL1vV1AK
UZgBXGEmndCOmn/RfZ69ybAoMpo5tMclm/5Msc8FjIT6yICJIM4X1dlVy9IbFiXSxEEYeHZh3PK9
VtQRxIgiS5fcelFY78pDu2hNcBdMg9HTDq2cR7mn7dmiPQLJaWWEV8ry9yjk/SIn1AIkYty18Md1
RZmmPv2+bPAeLBYYIllNxUng3aenA9vxS+UVsrrZ1zqDTxBu8SpfxSs3e3xPSm6Ioe43SepYcvKv
jdBYt0iyCWcGWUOIok+kGrioAq+B+qaDxoIfMjhZg1c+RVY9TK5gagBypcLffhNN0YPPsTSSVMaC
q9RSBO2QBthnWx11OQQTlyI7LR3+uqh8S9ZIFuYY2mponP73TWUlmGDgbCV71SuRPmF9YjcEoiWJ
vmcjqihjYaV32Ey31R+pKLaD/2SSWHo0qdKmNa6oCssEpnRkBdp5VLRHHsL6d5DBI4mOHqFtMjI6
swnoLH4Lksi7tMC591h2Piboh6GEZm+uu6t3WLt5Ox4Ck0c2ykqLvwsrvwVnHCsve6gvvQNOBG1E
PDELzAu0rlTnAXJIRHAydhgWN63E6HZrMHR74296LtTSWaKEEr60iKozofFZX6GOhE159BQ2dqNL
dwdsuK0eWvE1e5fFubHLf6AKoP5eslhYCtoiv6yRx1K1CIpslZhhsSUvJrEr3k5/vX83WvkXAFhl
2rPFwepfebDBIXh9w/T9pDOYyLi1RI6IYXwommh51pJYtS7iYdf/ZcRqiw8x8/HNw9c6c5ZykII5
o9/V1uEKKromoCb++C+pDfRgoEE86nRNKvmxKzLQShzZ4P4s/r7zSakAOBmLSSYhJDK+DJ02dkYD
6K3/GiuJpDE0PdWR5muvyz97oBB+WTftrVQMQTEkOm5fX2ygIwcIr05CIfggg9j6TL5EaHs+Czu2
YxLzjlAknnO5S9OPGt4maqvxBBmo9eOjfwF28XmyPMg1IDherA6ph+VDQijneFkvXY0jcytp5qcl
TdbjNMq1UwkWd/a9u5O1vc7GGtWMWzgXrJZXw7+500/PVi+bYNIzwPiRxwGwi9mFd7dRKj3AQAng
20xPbLlTVKecS1ut41H4ZDNG1Cp1i2KWkSKTsPxmny6Ip0hQrLhOyuagaeN9+ytbxtlLAWOyJ5Vw
3zYx+Y7ZS5LYTdipkjqv9yLRXMLM3SWwmZSgv3rEBngstoApGIb4/jHyBxLbcnS+Q3XP2ZHdFpoK
iDSGUgkc56ldAMcxOdeUbFMyNSto4w7TA3QrzXOvTl4GMDCXjx9LLvugnt0HcLJd19FslrtLcl7J
pK+BHn4TULE2BoG/DZU9i4vWezV3beymIqb6p8Rl3twyb25TwCL0CnhNrNkMkqFmOi/sYk3oHAJm
Sh1V4WN2VARPD2pgna1u1hxkFJdVPzlx4LB/pabdkpRCbDFX7sMg9mM6RcnkC1hsatEe/RAlYROY
2gQcA2yCmiiiwK+Z80KE30QTXrxnkoEUcWFB2xFMsZ3R5mqydXY0jfujIIUkQG8nU7m0ZlPoJ9vP
B73zr5cHnyASJevKMb3I25jg6P7Ev8XBd6/D7GiMoizdUyFae8elG0cPgmZO8pM0ncDsH/S7Kc7q
wTz2byRLN4huZq6WLsXD6bOi/G7Go+awC5Q+XeY8lBb72A6Di/yHMEo+VI6X+bJMk8XBq1qG3wB9
oNrqNOXyNJsgJaNP5NbYpC8XjWFjQ/ZiBcArz80gBO1m52aJsrc0Qhk9LdEUsCDIxKW6hYZcae3j
NfhwSZyi9rB29em4omjJxd1qEpzK7MFo596K+Z5M9rs0bRzEHRGMZ4ESiMCD5cKABHiUOYjPl83v
U/6GCQVfFeJjwl/ph3fCxPdNPDHAfU7prhNz7506B6df1zjOwLP0PpDWlIzQ0o5tsn2ugeN6td4Z
+E+auFGNVgPvq8Ltc31VuupCgqEZJX2Lv3MdNGAe86QYV4joIvuOZOCzITJeLulC103z0m67ItZs
6z+czNGN/uvb1KAyFxj207cXIlt9coHUfgvztGOVdkTjwa5rgNzqMGc+2vSoW3Lh1grXIiZBSKFP
Vy9qhik5MMKSYHDNsjw/RDhsbf/PaTfuCMu9fm5piVPddF3IyNDfVnwkrb7x1BLyW4Adf8jJkNlC
sU8T9Xmg/NAjEfFHv7Pu2/AtoXoV2Nbah/MW+Ti25sfvVyctRmLEaHR33Ey6tVmnsvMZCMekpWdd
1sQkvnp/DblbmWJ17Fg6Yitc6SUrx3I1ZYzeLz+ha4GrlOG1+pIK51CSUoICh8CKTXpoyppcb5DU
BCr2tky63FtT+trjHodcu6O1Nzv6RCnYX+U5aBaFuNw9DZZrRZYXFyaUblOfdgqo+T6CL2kiN3Wx
UDcKP3N530h+iyLFit96NjvfSJBtDVVBRo6fDl0PlxX2Rb29QWo1s+Ab5HwwbW2neF9YbIVD4v8S
vyceA+ls/F7+UZma+20olIqWOZe+gZ61OUM77JI4roZMGGDiRkkU15ysGUnLYXxNUfePB1KZjdBm
qQYQrvp9y57aP04M8RifMlNAPA3v5m+7TWatpiaNP4e6Iyhq7cQHSqV5gLuld68jSf4g1GCW5zIW
siMgmZQC0f6Wy1m93uqB/NoISgU0cRrmfuUUnPk4Bwh+Gu7+lyqwNAK9xyzNI2rO+8HnT7EexyG9
s/czQYusHW7xfTd4m6bB8QgJQatUlf/gazfC8MB8NIBy7/2f15ZerjLTRJrJc83rH+9PuuU6LVBe
r0vLYU1bgx7T8j+Tg9gVGrRxCg/1NZOPhc9XIUE7UXpE58KottWL8IJQLDj8sC1xFBeA55U9W3gj
QuYQsK+8xQKXYWOHlBPw6XI4KtWYIcKG3/BwrHdm/PUjOAfJlSLFRuhqIQjMTuWDBA7d2ImjIfhD
e8X8SEjDs/0UGU/gn1snQ0QZLBvRfCqNxX06tNxUrEferqaEK6HmBk1Mq7MaehBzQVrvsoC7r1Oh
/Us6uMyDbyXGDHKcYvVERl0/U2+hQmHwBAzdUFidnm8M0A61MCtlp1KZobLu1CSz1rXxXEkx7KSF
tGS6KGzOCJ5syXVuPm2pq+mMXFX5XTl2rDrr75kGC0D1ePSOLqvEK47s4soyIokkTS4Ch8SvKpDc
iH7Ua5ugPzIW6eQin0qQrQwiJwV+/96/myV/9xdqXY6I88Y/M2QZjeFt9ulSCrBwUlzNi3LYqW6r
fumfhVaYY4IuYhKAMSY4mDmvCmxjSyCvJAMrywwfyxclyUToxK9kBGktFZCgma6raGVNu/xHN3cs
ZAJQhe/nuEXJ9ZcIo2Lirq0BDgXqseHhPTo1X/+T6UEvtNm4TVWCEE/7sjptWZyC/0SGLa8dY9H+
LB1AuOiVVGR+GZLUy3okGQGT/JPzsimaxNbXMHBbkhjOgiMwlBxzq8GDNC08GY0k5pdxFKbFkBUW
i01vEd3hYlWe18IVojuhvbBM3uA8FrUpSJFVSHYbhvru0jZYvK6pwGeXGxeLSiRKMf6Y6GlpEx5K
9pVqHVZX69iF4rdLluqCxFuZxul9qvXtFzkjynScYyUUrmVzk3DI2gcB2S3HfP3QEuGOSCzpDnjj
YNH94dowmnUtG/UBUg5VdvkDBI1Xwu64uXHo6+0il9R+eCc0AHmtstwWkZXdyvLT8Sif69rbX1HU
7/rZE7AekDyjBsQh90Kaqmznj6xakH49MMmVtoPow9ZU32LJMxRqdIAe8xN5cjDv0rUtfudWeNjl
b83tLA2F6n3tHeVash1xX7sWtjLaV7d+2p4iszv+FyUnndc/nRlUaA+zS9mBC1Bsotq3TK5aq7wp
sLi/PaJaOFriWhQSDIRFAb58KgXguUHEZdN5Wf4vqfp7jQU7eLLtflvbK4GvneMlQpFh8Ik85whG
wVf4n9NnswChprkJ3K5cckI95D5jzuE9duKQiqzIqTgt8bQFSHinFFWJ/F1r/Fzhn+PyUUn3Eqx+
PVyJRkmYC6isGS4wyRcmwZtHpCuJRcvabyjS0aWNDzK+a8u5o/Nfrz1AOPwytroXHF4mSeC2BqLa
bAJFOWKf0H80Zcl71VVovkuVVGQQcoJot2/X9ZV+s4u66pXs4j2s5SEkOqr8S0udA+VEjUbdmM7z
GB42Hz4iW/bnD0mnyzvjCKjnSp+kwAZ5pieGlBMbb/pTlEXSq8s388N1OUhnxwImbVsqZXNvPa/w
1d9ONp5jHI01U2sQezilnNasrJay7jwCXzLnnjb46n3x3e7HkpxiZi8Ya9/T1v0nHr2lw8MQIe1E
QGdvh2hq9EoDUlP3RZ40FtQ3Roe0ATM+6Y241UfJXDh5zy2DUSoEmRRiiZBB4hJDDTKya4Np0eI3
2/Y6nU2VMYnkxvUbvefUYbMuLudToTrbNNEo3MfYDmZ/TKZUbMz4A6QL6bPmcMKydBgJ3bG4kAfp
23Laaegrj4/qdPZhjo86H5zl1rWlx301NLb8jHASgOHzpNuMVy2Ctsc4DNQqP3+WhmV+4le2LHxg
YkzxxIfN1lF78YNXULX7fU6f4W+jtdFutbGgA2Xr5tDuJFuUQqmfarS8x7ZJ9rMliUdCOOoqm0bC
C0OvPj2e8DY+Pb3QmZpOZQ3zId0R8LzOYX6lobTdBfvkzpcA2ZvyxEC9W74iNC33327lp0wcJKzl
ipU/x5t1/qEaJF1FOVRw2h9Tp5Te4pAW3FuyhHjYsB7zYgPeoxEJzBtqQT0V8g7MHIJDaIhp+mHr
Dt/DtJE7YkBwsqnor6QL9tHtGgY1h+t5mDt7dZA9Lpc0fjqfSjXw37cYaZc4AGixcBzBOThZlvwp
EKdu84cHgSWZUsxeqz5zGjOBA9nVPEG4uLvf2CXg9UoyYkduaDJt8kVBFK1v35EBN9R33KKf9pS7
0MJYrMPxkNXCZhhOiM59k4WoMusX4ItCcV+AevQDphfSj69WGdu01xGqbsGHukcehRdcmVh9r0UD
WOR6PnslQFWmPqMOurYLCCuCLu2s2aPsHPmpY3YNnUfsGKWT7kCUyeCFfBeJ148ZNAhXsv0oCCPb
TS+sTqI6zQ==
`protect end_protected
