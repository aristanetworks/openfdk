--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
B0pwukpsVjnTyUD6qzMr3C4FRxeLMmwNkT3JEZikN/lZw2aSNgLHmF6Zk8itLMyeIpOAqmuZveIK
mQxMUUH71vbOpT30+qCbBNBVd9KA1ETCsOQ5mURv2Y8IoB37bwR4rHJ8fYjX255VnSls/DGIszwT
1XuLG0e6Nqouh9PB3ZagzwfHxSWs2K74TkhQe2ffdDRWeO1pPgn5FRn8UU6CzuB6JWoMkda0BozK
dHWPi5TXlPk/J2Dm7MQR/8icquNExmFpVraSMIzFPD3HXi7+rGRVX44gcHDxQMmwO9YjczJkB5J9
/brERJxFhsl0xFFZjV6A8nZ6SfVOoDG6KPNFyg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="bcQ1bxYlQRIm9sZJfjPWRPKVLxIKmQq+bEpR12EzRqI="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
FoJFTaeAtk/e5gp4aTp+TlUujjhdGJvsfw6iXCUC9J0V5ZPD27tynaMYIr4YIjrSw2jHtz4ZV/ej
SETr73/5+R9a4x9yfEfBpoj3F3ggeLhxOj77SPrVtLZR2Zru8oaMypv2H0Kg50v4JUF5tm6emcNC
YlJcJ5gu/SPJ75JQvSsoHG+wkysglKM2mi4WCpAc7H7ic6F2jRhjLnPtfKEMuC3zRxWIRyekQhfD
/1lR4TWQ0hVqUawlaQaGPk+9ck0M//2/kfYWm+4YuOaioHiPkL7SsF3gHD0cR80n7RRBfm1792fc
dg2lD0cFnBEffwr37iZqK3HatB4KE2vy/s6rMQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="VuYB5gCraZN97wehTCLB0c5SBDcKkPiLj0U7mQ9bkaU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2512)
`protect data_block
McCZ+b3apIGhIanWNBPbghRWhZXX9ihAJo9M7bf46G9oG79PW/WgPvhjup6PCH52v1V44lYp1nCB
13yuIdbMdj+rmeq5cNafHJly0FaWwyBKJQTVWqRTzwtnYEKWtCEDRFir99J3bqDelseE/wVn8muA
XDwXAWc7ZPpXr0C2gxKN1TBmEqY+eiCgVJebNyUsRLPWw0tkr/oCrLsBFt3PEvmOYfzsiQo7Sl/D
CqIFSwZZIjvras56kTTP26AgRABsLOTOraZsWStTIemV45TOIGgIhj20yrw3XxQ/JK0d9fe0EKvH
DrkfiEaazU5FVwauv5Z9DPK/H0NN/SEZWihUTZPSoR9x04slmzhEdG9PLTAj81WJ5ARkeLhCWAY4
QEKS5j71kz/IAatPUNQ8cqmn82cir4oInCRbTkMAxmsb+6RrHNquZGr4lVL+qT7LqvGwk3q5oHkQ
pQ9vNO3XcGfv+mjzLlOpcV1dUXgfMW6b554qQmAMPYR1Xdg6oDCbKA8CpK2ShgrcK0YQcqA0Et7c
I9ExKMeH8o8mIOmI/euNNIJgv5cKxCco8iG5ihx0TbV59u2xXJMhYYFVr6zWO1y+jdy41dl9W81d
/HuLAfv7CtcQkQIjvyaOF4P94uFidkSIYptgbYotjUrwVFjZYbKxmkqW5s8Nx2V1HDVHfUUdZKUg
YxkuRsB7fCL1JUwTM1dYn8iyV4e9UzTleAeVzh09/hz1cOAdETMthtGoHSFKeUYsfuv6ZO7peRJK
XK+db/oj4eK48H+gf4Mmf5yED9ezUBvF+VJ+BORnQ5hGdyuteBjg0Ezd+9RY47FuwLdNfzmsb8kX
iv83A5TRxVBOg4faY9dqe+QgR5DgKuOX3QWIW0DaVAz3pzRBQG2pAQqLXJ/Lq3zVM327LZMRZo78
fsAZ/dj7gYNdlFDhd0+34nLBaaOTKnt/5nD0i0vvuD303cJSY81Y3DJKVFiegzi+ReDIF6og6HVh
Lq+wnsi4dW8HQ5TzItHD+Sgr0ryx4zTgzsvIAWtM5pN0O/lrm7ns3cLfa9dmbH9660MOswIpOgfH
dc88Q/dM+laWK/hmshGIsVJj7hLaC5YTicF/+eAY4m/jMZP4cHfFYXZGaV8AIKttFcdKG/gp4hzK
utnZIwVtJMCxGxf2NCy5chUd0LWtQsinENIq3++32YmLD2FAhYcMWuxOosaeSm+6EDoYeFbZgjsi
sQSK9X7UhGsIISfkGacF2P/GFvU3rHtSxFZ0/mzbiNB/Mu69hJsn2lJCmif6iUdzxdyFuozqdm+X
l+tfI8XCBINYJ5rTileFZ+/Zw98p9UAeFCbnrWG02xprK0EhAO5/luiRR8f4+SVomZjCbzJD9SuQ
jWVuVHjPQ3SnpAVxz7VAUVb5nCqIVPp6OLnfHA2CJJNsJc3SQgc0ygyR+O53YpR/Ep6GATjtPaKi
E40ybfUO2VeJmCcNtgXeheQO4ZCex2Qs9KRGxiMTWm7B+kDxIpwH/x6fkllSQyzR/FLEovYjdiK/
64uxQwmOHnM0Cse338bA69LmLz70GnSX6eiU8KqdWMj9V9DFwPQUASPo5SqRhdrhCKSbjJFobD0w
vkPI5KoAyUhAN69My5PcSwHQt85ftBgsRUBlqpJOr5ItKuI3CG6ZnQySXae+NdasV1CPNKQX+E0z
pB4tubZgGSVWY0hGQmPf4oaXRL3F+k6QSIAGZPNwvzFiczeUIY2k5DAkN2Ij50Q/0pSg75aZ3s8V
A/TnucFg7c1GD2YeZun3o21vZ5I0ke7jjfvp+sQAhcXRI/y19LKKLm73G1mvE/53wdNx5lVFGjj/
ePym95W5YO8aYErmEe3n5bkQm0GcMwiSteUZNbP0lALS9fRBpeJjycb222DR3Xi8M/8NuLWA5msi
MkafPr+H1lxD0BM2NEgeqZzdb17UcgbKIhRdtonOPbtVgYYV21kGBdetppD3Dfs9/r1r/+4PAVKB
rlkgBfH5/w1oNfampn7c3+tNUh536TPvUA7i9DRXAY3X2NGiHi7w/Pnea5WvZ2d1cBxBhE+E7dLH
H/EXinbnx3eEZX0YBVD8+gGRxF3aMKu2khycMVVqvdm3NYqrw/g1L57b7Un8Ym1JO/ZZ1d+rOFF7
/NJ9jna5OltY44T/JHpBJrJmqp0eTeQ2ijkXz8eH4zfUYlFPNrwdc6x+oQjEsSqfPTDeXscFqMbD
hr/2NYTfw7nqJHQzQ7aoKB/FDNLlXf4YUpySY/p9mohaZKhnQUgTVaadn4/VPlxgdO53DHY4/kc4
sEn9qVTIGGGJElS23CwRIlcNcmHJWJUGhN84Kmt1O+eOlRHgTaAU0pROJcmdCXw0ARrkv7C39PbZ
vRGx3A4gtQ82N1kU4qkM/9rICVKPCR5Gbd6DI3glC0j7nLkaoLVWpH5okQtXJXSPQ50cukO3lt3Q
FE+WPjdH41oTBoT+CJVvl0mAmRG5PDFWLN+N6x92Il1x30IlZLhI2Qc4YmOAaxpQO6vrPz0pDAGN
meju6sCzAxRty+2WZ5B96w1grBKOLKi3Hbo8RLzQa6G0dccGw/VP43PvBxHpNZz4ePAHqHpp397P
BEYcF9+E0Z0wcKLvw9J8rCjIU4rvn2P+osMA92uB4J4tsONCWzLgRUjLE+2qQZA1MH0u2X/E/IQm
sWpb8v0cBQ6/qD+jBhoHT0PYspyPhbeD8iETm28x5/lu2LqfbLpjuIZm6iy8P+ZHzVI2LQXVJINX
FCr9hPtdJPXTtHw0Gx2xZozvpyGrWcehbm95mWudQoNNeRZU0rkqdtvkN8ZIQZfpju7vib61cg3X
MU0IjwbvoQIObvQnklpN3/s16cFTvwP6m7JgzCLAmXDWewLgEg8yigZumB7hwFTNFARW/rWtq2oK
6Q15JsG+bmiJxGPv5ShUMlf/BptE2apFs2Uzg59nn0lVrZ6jFkuZa1rm1CSLjifq5Ve38brmQfzo
dK1WyeuNVvotsSfdMP7v3wCqV05mKXbnf+KkQjfOdxcfkS6oPvj7340Y74J7HKv5PrNJun5KYJcO
Z8hWg7fx+KSQYu0SJgUzPzE7ItxKeV+vD5NXHc0wSOC1kGFoOzGjMEXM9Tpj25K5Gr8Il78EXWbX
o6TQas6zs6DocVdI62kEC6rHruRBlAk+lCB34ZLhDwE0P+wZ/dz6+3yxLkKmJLQrjmZpu+POhLiw
/1uzSU2e9n9ujWSgNTbMf7sImO+iE1f7r8D7b8q2zhU8vEArA4075FqDCPEx5FX9aF0oFyzEr4pl
bWDr4MwIggMdblU9bqqWsr3uz8q5yRxQ7Vs+amCTCMC3szJKm29lA5CRXwA5bxIAsXuJIKbKVQkc
M0V/WQ==
`protect end_protected
