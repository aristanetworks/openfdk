--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
oG+0BY+AYtoYF/n6cW8g3s/KcWdO0rf2/9Q6tOc3kBsTs1Ghof30UhDWJWKv0z7O45tBmbpT2mkm
sMcQU3i9XkWTHMXLlvw4+WKpkUyhPcjFnM+k/+lE5XiozRaql1m8oj6u4wFWWDlglFzKF/BQfFL3
nJDHUxUcFIeoc4CgWpJ7irj8QFLfaiaKp3F/DK4u5UlYzFkiI39+IA3dk8bdfxOxtNHSgijpV3xl
MBvEIPtIjp8Vh8yPwgseNASUOBQlcsM2mF6nqFV1U/JQbL6ZTJEvGJQ6XaXSsKUQzb8GAN0i7v6f
WnXakqEBjr7gc3+o5SzHwhA/K5WSLfrRVDNO8w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="nkhspykfRTDAz3HcaoGsxQ6aley0vvZtrkK414F+SeY="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
k5qJg10tgGFltYb2q7sq4phNvCyfD61DxpmrUrKZjAFIuF2DkIQev66z3PxT5297nC27T93gza67
BT7GzvTSorJSkFZvdDpaKlMQ62HgPNeNFkppf97x5ZcFAC7+pJifgPcfiu2Mnc2MKLOqzA24GHwr
WtMwXa93GdyX8OzXnBagETNnP/STh/CA0SrnLgW3JRlemsYJftVkr6mCVzerUHzly8V3AigrYMQa
hETC/TgbVBWihzuaxMFLU5Li4GoW30Qul05oWwG9rOEUAzy2VzPLZD5HwiEvvLsRd146U3EQiIuN
oshmdL9VEE2ZJ/UO2r5RHVpk1W5J0jdfHGYugw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="zuUAM2h7wNQCE6onhzFkRw9+mJTbAB5rv/bb5E8/sTs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12656)
`protect data_block
mbrHJ/qM8m+J39gWFJN60p7X/bB+p2lZdG1kpezo4nxm9Vv0b+I9kaVAwd6gyOQkkoR6N7kHIF7M
wQDWIGeg0ggzL09gaY2q1BSO49ND3osfeFklDSR7fSRZ3osrM+q7Q8FaHlQlp9yc/szOKLkLEXVQ
RYhTscNwP3i5/PIvaFwlHKvFe4AB56CdgV4tJXhoAisafdkv76G98eXQGgEK3wDCq3hlxzETjJR1
hWw8LnftXymxQKmvO7pXb3mfY6h8iiy8t/vY2Zn0kovq9fGamCMLD7ixDUhZuRY2cjGdhTPkpLSx
E5dw1RhOtizvfvrOp0GdcWPOeTqxtZ3TMyuAbC9HtCPO6loOX3DW8T5d902sOOIDRpRfQD7RHagh
cMVNNx+GiKxo53TevECgM5wfU/05yJ64hfHaiYIpKZdIFmoH/MYK8zlKZH4BFQftw6gFty4kOV7s
qnTIF7lDoW/1slX98WAnAfg6xxz+YAnmwlYn2QcWdxS5MaBOEyN2upUao7/8Ummkc69g1wU6hfcJ
5KNDICZ98umprOJeeVZAssszuKdZ24xd+JeCGESy7X3D8iW/F95MLby0aytvcAjMF6+XEvZcMcr2
McqA75ITorTFYgHgE2kN4wLKId9KJVYw6OVe32/b8kFAoQYUnfVgU/Z8nXcmhLf+RLgnQvlq3l3F
hyM6+0NLY8m2gfJWCjksiMCgYR1BJl8/77S8UPnmdq9kWyGbxWHfexTH6n/iuo+TiKMjMLHJlzHs
THx+Ba28NN81JCR67Vhn6o25khsoMk3+Uob24WLBmNI2Wmo/TuciVyA05Vn7z9zn9+n2fES3sjWi
mqXdTf013FdO07L5waYZB3/EZFeA+eiiJhuvANn51EmoIztGgUcD7A/jC1FV+1nfXQB+MgwIAPsZ
XygSZfZNirSe9BgPnRhT2bjXytZPg/caFoCh3I6k/lDCJvw9d2mUNd4WGcChBmLMgMgvrTAgTfcL
eSFDo2QDyUmYqtAH0+zr0+Tmpdlb0bxRrL3CFi8813IeqRgu99XUPa4oryf0G1EOxgEekYLNE0su
hlSaDlEVA3fPkTS1dn4QTwVkFa8VNXOj4/5GATmMeSFz/KOdUs267eaLeKwrsRe48rnMuEnerOvc
kP67GHa8SZMd/vHx+q1boxMakMt/Jr9r66kX/kQveMdpOOhamRDy3sd1vdAObEoLdMfOPx2VXjPT
CI+B8DPQqZToXlectVbH8A7cbTV5X7MfVFjz0I6FXvAwJsE9k36KIs/egM0tPpbMtTXaIWvHoajp
+k0eDXU6TTl/vJqkGM6n3dawQrQ1mvmgeDMjj0Xt+wS2s7mtOzEf9w6nbSM3hsMUxthc0P7ap6Uo
OCoixJ1Mu0Jdn0oHk2v+JejGh8iFMtJy50VnTo1Vj1dDcsGCY6skLqDYXlERRdfEi154fKtEBoAr
yfPSWBCyMk6w/VUuoPjxdaZ8XLJUPyYpW59k5s9Ycx+tl2LVTC3ghjRDsxDFASp5180aatK2dAId
0YkQWyO9e9TQKSaQkqTaF5LQcN6wGtwgx0zID0d0y6D76ka8N+ZLpeeLjvc4hOnH5V0bDLu6I80o
KRO9pvkz60rXI0iSUBu9Q3OeEGeKMX5uB4sTU8HJbK1XVW86GPfxkHrFpkf9zcZczHzumJ7yhQAq
z4CXtrTzngiYCkIvFqUWCKxPtRhfqSm6TpfVlczS2OCLJlzh06E6HKU0TrY9B24FnLAGI3A7WT7I
SGbLQ9Gx50vcyS8HX8RRztbgcXi12gMUZdxuxlJ8HRZpN6O4Aq8UW9QDCLYkGlbwnmGp4mDCCbr/
MoI2dz00VhD2y36YAEfSBU4eZAqrOtX+stDalGzhSgfFOjD5hG6QmkKOJaWGVkVN03v3rDwn64n+
XdFxjq2PVfepVwg04hjbsSUkwktDsqtoO8k9ITLpFKNBe6VbatOY+9AStctUAZnJXHAQqmeSviSv
cl4TpGHXUpHTvpko0x+pd3+gpjye9j4HYEk34C9xKIIVn4QTztclXdygvFYk9DC7Lw2lmlu/d/iu
KLl57WKCChjbgNogbtC745Gb9oTYGpi0/Z/m1Ed5+Xuy5GgBh9fbahgNUPSfvbDDBT37mP+zuNQv
Awx7bonVys1X1M5o0m+Jois80cZhID86ry8cjg0+UvC+2M7+nUgrxvPwG+6Vi6YihAZ73L8bQvBK
6ydrk5e+4gLW7SmtZT/2Fj4x7z2PvqHGiu0L6CFUj7AaiJgtMWxKoGcZ0XQ8SqewKc+SKCulBlxi
RcZOQQ/HmoS++W/f0V9ZaVJ7Bv2S+zZ2F+4Hz3r0z2l4ZcwTHAQNHd4yCROnkJ+Md1ZPmUyjdQqb
8mzNJ8gG0Nj6fAu2SuRVXZ95US1Ua9K0RjzVpFkh/qpUX6DG1BFDSTEEn1p3mot+IoTO0xQre8hG
GMZWWI4QIPZ7zS+yJPEx94lwv06K9ybuU/yc2y99aHP6vfpIaMOOauHqEIYlvdpop8nElQAEeuSg
v0zV1o1cd6PS/IwaI9qSHVYVxuwAD1mP2Yjd4VHwGiERsGpoXl6dNtFCLmhqTGF/I40BPdMjbrE3
uBiXqC5MBjEmLaT2JgIbXR6kSudbSjBuw7iuRZjLNig4ul2EnmcYo9B6Fi5STDKn+bsDH835Xygk
cw84UVpOwDEtKw9sNG0y5hkI27zWYcgNCRNZRpxuDBvDKAgxFthsruXPTRH5oD0fBr0zqDX1C58W
bwNOgUsgrA8LKYPhPlBZBaQEncnTCbiFAwGl6bbnsQoZIuxHxa6wlGDXMw/rk6R+47Is82WSrAtg
fSVqLOuqh3X7LchGVSPAW8QP+5nI4wtlUyL1wPEhAqNN/2vD0/KEBDfS1XR5E1bzbpXaEsJuLX/Y
GmKsXrpuCj77oDPT3UbX1/wZ4nh9ZtWHH31Ulx23mVVODCN0bPN4faeM2FP+qlv0dG1zAxBQS+V7
5AG3uShfoHui/bOvON4R34EvEIhhQEJVWHSlF/B8Axpsf8XOADhIGrRg6kyMtsmHLyTyYuvEQ7zM
R8KBSHdENSx0cxRP9P29R7Q7T47pAPapvmNc5PcnQOS9oViSNPVi8R+M9bRrxR30BT9L9GlAP0wB
evCAdDXD4Z5qz4+a9wdNZi2gTQrgbSuJjihx0dEK8UA1XXxS8jqNaJi8NpG+PWUc84gNtqiWFRwP
UK1M2kCWQggrOmcBHXk7kp4sWbhGk3flkNlU59LX4qdSbAkXtaECQ7w8B/du6U2tVJnUXkyVIcEC
5zO3006TtJdRB/s/9Dpys0vA4COyME14BG41ijiMFrvVtNqnuzpwyaIPv5hg6bjSYqikqBB0YI/9
jHf+7NTL3Af/7+rXUPyCET0eUHrGx17x6M+gSqedfeoWJOs5D+Lk6nBe7mTUjofnx1WOWl6qZerY
oEaehki4w9dwL4GFMpgC63/SKgx4ul0Bvi1qg86+vhXbiN/EN1hkRMg6nhg6jr9+YuV+N7+ICf84
C3LqvhWvdUjc1Ss3Mx8cOXeqPMv0OQ8EGAGIDqVCwXFsujh7yQuMcGgfkjtD948e+F3XiiwlQvrG
RYqmqRV3TJPYkq6qnhe+10XowcIHfpE2inUjV3QlBn/Jl0JKtstzCqZpzkQBcCbLOzndWe686QwE
E3Reutl1N7HBVRGQgaPpQyYpo5N8GgUYkn+ifLf51Llj9UxZ7urQjO+8EKPavEd6iVZE0TiDa7jG
DbQo8Xx9MBkEc3n/AcR+zO88+lK7A9y1yuXBEAjZx69YvPa/UFJE2DbS3COW3IuE1XprGOdijx9v
E5vHE+EyEpNJVwZnch9GuJGFZLeLVOzLp+Jfjnbmn+q1at0fmwiPfnAD9k4j7a4JkXYs5wNl79Yh
+2N1/1KFUB3lxwqPz4n+BiZ9HKYzkHCwkr8/bFg/qlzcNfOAyxfJQxYta/BLOoT+/bCqjO50HLC1
yYGn4aED9AfLixB68TYZ4xWeFK3xYRuOVv+xy3HhdKtweeCoBc2uZGSqtj0pgN7i+rNMy6284fvr
yNh77tiRHFuJ8uS5zfmOtvpxh2d6lJCAquxuh4kdTIb//j4Dyy95jMkDliRbB4Srz5u/gr3yM9vt
fPHmsVZDhHB6dyrAadEZOTgkMhMBMDY7M3zAnJLh5RyFv3kIkMP9/t02NCj6aUlzLhjudh+/imT5
hFStgOysPr2EGLh1uijTjgAQYbNsiyMo4Ux6ezAzdJiUYE6FUNv+F5tpvzUDmiizd2vDcG9csj5J
h6A9tOwMD98nIPgvX7T527Uhqm5RiWEirQJykhMvnTbEN0zyLwLxFkKcxyZsuDIEylNlyu7jDYM0
+wVyvmVmNw3S80c8L+VElayFAXM1dFNwz/0Of2yDxg8QH8DLQzH3do+wu0rKOpbdcC48mvDqotMA
Sn4zfQlnvQ7JrBp2ip1hOektX2C0H/8gOFKRLtcHNqaYFy64ILmKGJCrwqvAfHdeDw4aC2Iz20mr
CByXfNkyKNXMo6CwIhgb4/YODyv9qBETgX+aSHlPpp9ajyYKK/a0eUrBhJM40QPoy6ajQNL1B0NE
K3BkGpPP2lC/8KxfnSNW+XnJfKsnUckW0vIBgjxCapKHEhEMGvGCGToprbG1Kaon0eAnSZQGBxGa
MBy9h7sD0umNhh+M5eKG6+2J12voLZeJp9Lps1qBxnyTmr7H9ILeX2RgnVJ6bUA3/KNinFn5huVC
kSq9zaklkoWHdfgQBNO1RGIZEIkdoB513JzlrT5LNuVz+dJJbd5czG83IkVcbTl021ZAp3NKxuI4
fliDlfClUAb1eCSxfYo6sPPMqZem8UA9zd9JmKRF/8zvNifkzGB2XBrSm0k4Kt7q/jvyA+dXY0sv
5uZju25eVZBMtDncRUUpf+YA3TgUFWNTlilJUs3ugSTY65TuBtgfId0cVzEblhae0j+difl5ERea
B4T/C6ObEUwqsHVl9/2+zqtA4pNUrgC8ekvotlQfyW+usFMkocd9LwDbWYLLW6KR2/N+h0MpXBcC
lx24ihsoqke0gJg/6XC6ppCCcqoEjWw+zAPzlJTvzvN7iOF8NQWHtHwFTixzUj3nZblDQWOusp1C
VqJZmzgo0/vdXm5tAxYU2gBNaCbYn3ARuaDnl7WNqw244S529lEpM+4Q2X+t47Dd/mK3v6WvgQ4i
gGZmTQILKM6srwU7Csykqc8Eu4IkeR6MJmxo5kG/JCiYiCMryH9JZhE087Q9yM37b4iEddljzOgj
MPnbfvOYhZ36LN39ucLuMs9+RH7eKRND+XpvDARDtCIELZa7uvuVCvu5XfrHdxXYMmwbYMSAWD0G
3cXggVD05QJFlCj/3pVkhcphV0MLmulNrRWFzfKoApR/R0YFlHZY70gkHMCzu51Aw0GTfGof6jCH
sS51t0f3src9sQ2z2hFQEivJ88AbLKykZkitoQWjSSSBbvzeORqN3cWI9wuy8XNbxlSUvklujV0+
G3vDWQNi0oMm45EVSm0JQNfp8brXetbtKXc0eu0z6aq+JbJJp8jA48BzQvTuzuUm275WaXwDTw0d
/7F0ihUZONPLZjCKgfTcxHEQGK1drpY1raF9TDxx92LoPKOGD1NNyhdZlewfG3AVgNTIgwT8w0OR
a0jAlEth6DHrKW4D5R2K+GIR3je1z6TVxtj1kBg/d2RupmAhKBrUqG+3OpTJjNZf7ar6mhQslEoh
0+nyN9tJYXuPbFsbs9cZhwKmsZSptNRM87bPSt2xyJJ/v3rhtENM1gq/iIfGWzVZKUmNRP09v4SJ
J8zrQh5H2KsYfhyLVwbyzMqf2PPnG66mfu80ITdwtTqQmOAQZY/c0pkAy7U8MAGkoaz+kuhOrMaT
cT+ApuJxsp1+IQD3f7qTwWPvbRxhLNEhuNiUXG9NFgEApot6yVUDX7DR5iCBB3faucZkeJWwReqg
CQql3jibz1oZhYtl+2D1xfG4LtS29+91QCZZR4jtMXBdOEL3Q6vSvDhmpraMjn0ZbgvieGvxI+2I
m9dotsjNVD8pdOYf53KnaH8+RnSbqM98wKLlVVvw7TnI1u9M5KdoYXnQ7RhuGZP96oHltxc7T+gz
am6iN8Dnd20HOZhXku/N2cJz7r6Io+5jQOfIvocyXFV0q/ucMrWBuGTDNMs6vFgK+dzCzLsreTOn
hqjePwnHUmnf1SuPFde2FLDa6hbql7XeVzJtS7gDpiUGY96ucMZ2gXAPJo5K/IpnACgeCPVDyIsb
Jg6dd6UieP5vSNxHO0tnpoBDzya5uJ15Cgj/PIFKlobSdkK36wCrnUuX71gra6d60BQCzcvvQYid
r3EXnFjHlFa0j5TeJKbUdZIMT3xGUDIea0sN9xA38imOAY954k4EsmNlPaE/X1yH9uBZ/dQKOpPZ
ZxLdwm6n/HpoY30rtJiSRmDY27OmlJeoCXzUfEynF8H/gKczgP6eFGqQ596SpXsZx6Gu5iJsNNQD
mfGlzm5FM+2d537ruJ8fq2JRnu1QgZEoy04BfkOUWdVmreQakgJNUIUhMvkQgoACRyaMehUSM8Ig
6RGe5VPw0w7qdE5fpsFXOtqCslvr2IyuKcfZqHoVRxPpR8iaCkBAxI1WTMuWSOox1aejVCh/A5Tt
rMX9Asckp4JvqNaWhob8sUs1eWpSzoofJWmLTpoSk2fiAPiz/YtI1b53QS+1n9T7JSfPxfAWxi2/
xGxXItNa3426CzpRz8x7ZO5uxkPy4bQXPpo+ciRFTY9jmvBijtK28LsOxEisIp8eD+9GSOpCDaq/
8TrkijhwoAqxDiezsG0kfmXBDQ6ypzryHwuCycA/Kr3EaHiZXpRIq4ZWGNhZE0PrftvyL4mA5ep0
DhjI9glOPiRtWS8ItNFP/wVzqiYIcJgsyhIZ7Hi7yyeQlgkhAlmTFgLIJuN/FXEwN3yJp7RS4hJ9
2VB4hFk/1KJS83X9KBcd62/aAD6UCW5V/hE0cMUs2PPHCL+4rq6iNA0YZvewYI9zB8CGRa/VGyig
v+OVpiGZOUmAqjLwVeKnMyoqFLOoOTUTwF7791Z2dA/2Rdwj1L9+taY5KbvfzERbqXHQQiWCH7wE
HVtm6fyUdSW8DgD1Ogjp9RNht3sI8XiqUtKlBoftE8a6004nmKct9R/C3jji76LedRlPl2n0UEXG
ml/OCJ55Twbb22g/ZLLht0dbunviCJoVoV++3pXxXyQMw0/gzKuiNW8v2bFgSM7RUq91X5yJMwqa
BJSpMAM1BPCaWJjlGn7fLqR0Uhm85YLoalpUzrHHru9LP7Y9iWxesbTFlk/cgN3WitSaT1WfnZ9t
PwncDCa1DZwYrHi3yfpvHafLpV5XFQlEg1u/8ga69wI349NcL4fngJAmIBZ0AcszNAfQf1GW+X2R
D7mxGYhWVvZlZ4gyI0TL2HQE8jpojHShZ11djJjqdEWHbY65/SbJWTc2XNQyBa0CcKN8VG3YizjZ
IwMYn9Eru8XYj3qWkKoLD8nU95XXYRf0D1h8gOyAu8YnqU+tmBGBWBEN+v/om1rUMGs4lKkZ3rEO
mE8nm9B/tX9KW9ES0zJydhVpQHmQgY4z7yIhoixcz2lNMzJ7Ph3DaCC4Vyl2vPxTw9kyS+pxI+/W
w4lQb6GUGSq1idBZ/hsG4e+2ZYbqL/sWtSRvjfeKEqQdckHKnxXj9kYEe8lmd+VuwYynI6268if4
ETGrgx0bVxzMq9b17tJ59l5varE5/t++RUgwVTJq7yg+bJvvs5fAG104SgYXr4jXslo4hBKpIngr
11nYEfBdQKvgOcjW6fNC0tgBsotyaO0W8wlqRT66NUV+c0KRzfMbUo7hxwl4neRip7Waw2q8jtmZ
vl//SLedeevz77JgWVpmEE/0LGQ91ZDVegx5O3vvEdSPW0VKswaWwuQpIOIa9dfC8RHz5G4X4Vpg
o/IHDg2sWIy/5tEZb3nHQWcjc3emjtpA50H+YJHrhaBmxLWWLKq9RJdHWO02UANAQby+jIQ5Q5CH
sQv6el0Yo1UClffwxJMmziACaNDh0ck8RSSuKLFyhOoT4t1nqo4qsHEtalyVnVDRzl+y4YU0T5pZ
il05VpWz5p6YGWwQ1uhrebztz8sWX5BIoeGPJTbsRvznOF4NoW8GCCrNSkUzV+XPv52O3uCLvOEU
tktqhX2m1ZWsynUoxB00DlVI+ebxfukCzYAISS+ahH35SbRLrYg5Ng+cuDKS8+2rvRvWvdrHF7Zp
ACDpoRCTEC9e4ucqunBUhIFrHCQto4u1YRMxIrBTXR26Lc6Zh3AsT6qhqAjTxOWcuS6M7+MCVl1Y
SQYtBlQ1HDfWBLnpt9p98YHmR2Gcu70SH+x6n6F1EC8SaSIW6ZKoia4CHYvtbxwWBMGH14NzvqAJ
GmR8SP5bzc+g1lDXmtrxDOQWNJL1B3EeM+Jfu+rz8JJZkcopxSs2a1Bhfqeq4/cPUcVmdje9RhGQ
Aly0aaqDZst3N8Yzs7S2fMukGuHlei2RepYdp3MmHPkGEUUW8GVAt1HWANwk1MLRsNkaQR/fYynS
TlQU2nWWudyRpFiUblKCMHDOhJygD5ih006bjOQHKa5cFkFPLtf3/uvbfBHSHNBdkcrflM8cYicI
APTpvvS+ZODEmhdkEsdqGqVm7EoLDlLeiBn4BC2LiJ/N05wJSe9RmXnUL33eo3Hs5t8BujY2DbMC
H4TIRbKL58f0Or0HFfZ5TSphWUFCPQTMbJQ6dhkmleU/QLNH/HkLJ4fFqrmi463WIekEufzVMJBr
RxuhcksxhAqVPvLRWjg31+JHPeu+VXpv8mn7scmjeOQQWTxgp/dDAADEspaUPbBHpRhAVYtpZcWh
r96zXZm78Uzn7so/Hi8hEvwI/tisoo/owuk/pY17B+NiC/I6F2dNAE6E6NUL2FBGl/EcoeQTp1lj
os+712Y58uJmwToWCDDK2/Jaj5K0JlhhAh46/ddQkyQqTKDMgon1eoBMKdrvqJ2ydPwoKDVzTYoL
N7OlEu1T0CLEFMAgndhsglfA4mQYaChl64yjG9fxoHbvMvmPerAo472/qe1qoROFywmXKglAbYpD
Dno0r5NS+99lD8OEkDKF6UkprtUh25uc3Y34wdsn4K4eQzWcDQ4asg4IF1nK9PdePmuSn/ZeQ7fD
ljiMoN72I3hAFGeMq4fQ6S64X8dnw3Kd1AfwvvYX6TpkoMhq11MtFZqJf+AcsE0zGAUOqUPmTTum
ZM6f1prnRURyFB6v73ed//YKblszagkwTkfNNFKIiPmuuANQ72R0yZVDB9sheGSFCqYHuPWRx+Wy
AIpthl5zpHhSqiu1PhON5CanYsq5dWavDzhw7yvw4ihTlqwSO0bcPjJzXWof2360fD8aexP9EqGF
eoXn0Dn4iu4ORMLkEuBtUmo4E9SZwCBuP7hB8gHopAK5zCLhCsxIMJuzQNZDACgd3r/9d7dqE0JT
tKGowubBUIexxX3NiLpaIZ6Tj3pXPtjsF/dGP+yVLHrYbAzH5drQ+yzNgSsIJdVrHHxfl5A5/Y7M
X2ZSLg1WvuZY7u/rweZNg26ALDsJTjQ0uicBo0wOwnRAy7w2vTeS7yqAczuhbgsuKHDLOzqSpun6
4BW5/DOHWyjYZF/2acNZh11XWWronZU5sSd03Qjo4Qa9zmeXYYHGIeZkk/UJtVyUa3ZtNHg8D3ON
Dw2ZBLfkgOOL0W8U+S5pYUql8k4jSSE52N4mGeTUbTOKklp2FbevCxaxCULBl4g/ZrjhnXumTq22
8df6abyljUXKeMZfEaoDltcionS+VO6VhbiRmarHRk8kfc3fc64eZtsojSmASsaIdoluGSAS3Phf
9i01FipOMJ+m6gWbo191vqTqrJRvxamLDVFvM3yl20CNezFskpC/DQQmQZf3ErzcSiIdzozn8ld6
P5hLySZVv/2ZgFtbmAC/32pPyvCi/W3kzgIEUB/hSMWRGioVhTF8xcavPGAbRwmWrTXTQ9GNMOo4
0Ktd9FycyPCvZZ1bgi5Dn3d58Q4c94dHZQj7m0WycECsFROMXKf6Jc8Kaq67Bkbvt5hO5/mM4swf
i5DjTtGaL9j5+qH0YYvw0cK0DXlT1xO5IViSPWzFDB320WBJfxG9j/1aHcRdZ8AvVQSEIhGf8b28
QTwxUg2Vj3Df6lX+A7e/C9IUAXff/r5Ic5vnkCx/WPnjEr70+oOxlWvMLVMS5nlzdpqjADKgo6q6
ZGr7T3QXoePKYgM8F0/KzXHoD0HMtoC9UFIGJIEiegoLOigFbIZmTUb+kiXAlUM/TnjHMevHQBsT
VCB499rVvdtk0aS4Sc7BrblE4v45CTGUPVSgOU6le44yTeV1458WFEuCpM7G768bH0GRwQt9rZBF
TpBgZTjuz0ZLRWhvGaKc87jUSNPTPsruKaG9iXLPLhZcgeb7kWs11nRhaaaFAIno9CNK0tIYCKQY
wyPgRUwJDMFD40gSI+6CFsaNFV9w11x6GPbpZ2CUEUafqgilAEymO/ZvW01ixLP8V7lanfEnmrxY
/KhzSHfGDB83/c7+TAunsjIVhZ1K6AWXH71GNjJDE9XXh0SQLF9siFBU0fcV93HdulcGGO6tllx2
UAkwgU2xF3A01bFBREl8XFOhOPD9DWGz7gyzfqAq5nE6u+8Aeh3dBiPb3LOF2cmV2WXdfPd1+lGq
PO3xtMj9oUXFxM0ZMg2AvUwl6wC2Fkj5xZ5zBLoQG+RDO/4x2IyWWP3z/qVseR7q83rcU35LHprL
SQa9O6aV5uC8We+xj7PgjgyxMGLUbOqUbkkt7G8yjWz3iezyH3JMy879KHshjeZMW83KVOTTYEeV
7xhPn4kf24NjTywLHSfC6T/CC8B3ij3mZ9zh6wbspaoiat/Ct9z2nzChXGDCaByADFaUThTK/qZ9
TSZpd73fIL6v2yob07YY+IK1CM8y+0+oCHyDZGPOqLnqWWc34hmM9KBvKxhUDI+PV1OLYoInlx1G
QDNUjML7xW/2bVWEg5khP8RthEwbbExbpG2wdAynL+jQ50i5jmsWOAXnzpDvlE/t/qjU8YXOUCaM
HxdWWKZ0mXwH7o6EVOcThuPKHT1pLyfqv8j4endKyyyKioMXRKrYqlqfT5RiHpEHDXDKIUVQIgah
kuckKZXEU7S4C5d2DT2a4A8fTBVmHK5Ge6Ok1netHK72MS+s/EDHyc0Y1N3Gh9jmq9FbHHkx8h8D
5dkMpCpRXHQpt/fR+DGbivoXbpp6vz7NZP4mpzZ1fmUC4toSIM4M1ZrIkrp+Icto8tp21Aqni+CI
K6g26rrmxEpHzEPDrfOycOJkDFBoDo1kiEDTHKqhVKaotVBwI5k+tbCN5ftoNT4BaVeh6A1AneMF
sSNmKsqG4F1XldXMSy8LSf9Q1l55g6hUIxAv1smpsweMnwGAUHBYVn0j9OF/V4kWQdjPaXitMTHh
YaGKRnQVJtqLMoT7LC9E3okqK+aSGAfhkjZ9cTHI/mrxu9Tg664+rG+6azlAHZ4aIawDntImB/y5
17QkTGlDO1p+CbWHJpX/rVwkat1pWuN53xwUyFWa5elRUhhE0nfcMxLNNOFpbqxMWO1Iska9vPPX
IrNcjjWPsi2yGJhGgZxpzpoSvVxfd8dMgKpBXgdy8MEBZAvtqb1YJiPHP+TtOnnTJfdj/wBeZxLq
zzWFuZQi+5CrF0RgDcLrsqk6vlZvWrjn5NeXbX6mU4Qj0KGSTx7K1IB1ktNvBpi6sEeFJw4g+Fg0
WIzBrwL9cMW4Xu36FjUVtJxQfC490Fy+4OPmvTWa8aJjAoykU3SdeQI+/6rOIXHZBHjaruvF+8Cy
w9SgJpa1QuTr0tyfj1RADy7CSwCv93XiyvAmfOA847nIGwE8+7WGzDVoDc6dbHQ60Trm07qFrIr9
//QFKiWyhgkJbWeBOwwLYQaOWAHhVWdDYxTm69J1LQr1vktZv+4FeHmKbUjvVDryK7RLbIDbJVv8
VAPo2EEufB613ywuFwN/Cm3acUBhRg7C6hTBwHwITlqB7Arv0IcOXdZLPEm5TkR0EplvuJ62fJmn
p4AzFEFnc3rzX+cL5535WZVTCeJQ9oOAURMSLDX9PGRaj39p96B6PUd0GiLV4jn3AeWCCh7Tm704
IrwLtSXiBqCBRdVr49W30WG76+i+62tbPRGk0ok3lvb22VDySzVqHYquWvkbQIFXSkVtvkTAciaa
Lbi2xPpVEAnez+53Odb/5B0iC/PPYGDKFxwGLmGglEujmmWSjCdJ/5BRVaGCDzkVCquzxw2Dm2Hq
9QczAUoVATDKKAj6JiQ/4jPKxseteHK8Ajtfh1VzSLVYt/rTet5L00lK93jbSAZpwMjT2MATGV6+
EJdc5HnsInbu8e6aGaN4GWTQYkzuRta7fbAvFz3uvjaE+nFqYlbfOhiSezBuSxuLcl1RmWjApQy9
bZEq3nWY27AWPOxZZZn4QoCb1AQbH5r+HDJ9ezGCCDKFZKIV1zNLh/O/wnmq7mwBAfqyXVJhoy/k
yf8v/PwBrlW4qAhaFlLWiT90KLW9w8q16VnPVPfqZM26kfoYy523/DApd77pkKAxj1H2cqlu2g7b
v4uxeLjHlpQfoR2gD8NCpxhRrS/UD+fOnxpb15b/kg2UqQ8HSgJsZzuZfgLQN50JYVpzOz+d1+1/
bO9OCspmjhKhan9YatjbzH5MVIggvaBzGLRemJxkk+TGuCm9gDMEJnpKit6UK0Tftz8shBgsCgyq
8+KqiLORAOtf5M6txK5G00UpDznTLEnssEf+WDFgKqUR1wX8R2fno2+hAR5mdyt5jgl1Vm+ymbMq
vBXCEYhFzofxpSJvGA4TUFHFjzAyMoT86zf0SbezXzhzhuQZrququKAHMVjL0tAaeTQeQblN1Q7A
0uB+OJE+HTX+F4sKxYe11+YYNo7SYelwXJp+d0/yJ7uv3Ybbd4q0qJ4vEI/HeUJOvwILmXtV4+yd
gZmOSRjGBAFbJl1T46olZ6HLpkZIM8VpVveuW4mzv9c8snCSDtBHWUjYzZ1Td7Xs2MOdfUewoA+E
rBsmkGKAbZQDNvU66Du5sCKDGcVW0SZ+1MOuQNlclMtaRUQFAB8Isbxs0X/6JinDcLuqxBETRnwu
lVP0aKrWDw8RRLN/uFoGS8aQOph+uxLyDH6R3mvHPzqqcJo4paqFRFbffwOCWQrfkgp4nwTt/I1K
olZFy6pRd4iMF1eMfQA+8uA55NCfGDxxE90Cd1k6HZx+nS3aDmAV/6gWd5Rz/4kH0XBYS00Tuuqf
3ks7xOEhNnEMjdboya8P55Ww4ruOXajs7QqPJ2phUOC7v1JAdpVIz9p5lqROQt0PfdVvdm8MZIeT
S/r9m2ZHXqDpQxJFC4k9Plx3nx6/ei1ARVEfHpIyMCNu8COXd4zdxVH5lp0UYMYsfL3eYPS50tjo
JQFwM67LptvPxAaKtslEueQhnvsJ2jo8GDYA4DwlYLnTbWKiB7Q5/aTOM9fKAeznBiezbUKCsS3W
lqrDeYopA6OUTBZPVvDjPmruWmyVqQOW0s3LlvvTNHbkwXFqHRGtcmja0UAdhgtSU6kYWEMD2xTC
EfqcXiSpiWAQrHQLFPvr0Q/GnRMXPmyuL27S/s7PhTZfMu3Ak+5c9UUFYFb65QmZ7dVPuW3F95MD
x/GDnL6BH2uCL/rkhCAbThSfiEev+8L5JPZSAC3lkwW4AUoYu7rsb9ga5sFtqsr4PX9jt0IfTUkp
1CM3O6m5dNgn9/PTd6BeN0X0PMKHlAVu9aLrORQLR7KQCQ80AGykYrsUtbi3FEK+LvxXOdteLo36
j3vlq4EevFNQ9zrEoc5z0GuGwkn7kA06pXXWTF31l5Ud+hPX4tu/qL4o0nEL/9VG3ODGLyOUInZ/
BHhIisP7iIVZlb82nLSwLhNNOOd60hNq6lodTTnYi84Mdi1gypVXki7T9B7GU/8br0yUgiWNnlqo
pMDbYroxdNbc8mwtNXUoH9nugj7ZKiPQnLNAOcfV+aUy7jsF3tBMmHiOPuX0sLyA0YQE38R6LiHZ
MxixG1+VGLuCdN+SYBlIwT7c39J3En2n2tfRqaehsmomyeUPXIca64pezi1IHPmV6ktheoRAeZ2c
I6lGafXTsa4H/m2VbK3emUyjPMQBJsX7Zd5pFrMm0oiQGsSklgc2bokmOdbHXmiE5HtO44JCCXOE
vAdbUUsRM18/5g7R+TFs6BwvsqkcOV5wL+POO6yCQlfY857CPrTcwYyvpV8TPi6MOsCHeTFk9fSO
PcE2n26Fvq+VW3DDvd9Mm0Q700if3dbFmqhC8VSid8XWhjJJRkq2x8ude1v94iMKlHbz9a2M3uLk
Z/Tx+x7kgulNVurgfPPTpjgHSyr6Bd+3lDuDe7QO2BSwDPNFHAO6DZiFf9Cg9Os5xkv1pYNuWoDD
eMA2NFGdPicTUL/c5TnX9CXjzPy02tFFvEJlC2jGz8R+aLei4Djlz1UR8nuGm6a0qwN9ZwRdd5j9
FrMLa97a1qa5v7+zunHw6McwgeINZQ6WM4mEfLexOf2t4IhttgO3AoOHZWAaLrWSB+ic2MmT2MYq
4aM0s5PI5p++6vWks7gz1+mew/rwvih1s+11iAAj0J7KJIEbFQy/SzTnUPzL0MUtxDaAD9Jg0Bw/
gsA6FI9CLHvGlz7w38bzMYX5W1HDYRVH3guFTVCpsxovpsLSOZdARXf3KbL0O65AjkkWGPCLmnAA
loEzabfNtYNtVGmHwX8hQFbyMRT5u2T87fBBQl/X5qa8amNYkKnPOQ/Dp40aTeY2dBlsFcUg2xpt
HI4uRaW5ug2rekTtMzDWUTuAdYPv7QOE3v9r/pirxe9OCZKX3CZSK7AZLmypst4sj4+vDFRm5/0P
6VfOx1VrufF11iAtjgmIlCOfFDEF6pI4a+xDIubcM+lZhrFkcuCJzzMo2orgAaboVWqv2NgBvbFS
ZmEQdw0rxoT8sVO0mIZL6G1Y1ZNXYB5OAUYrJ4Qtp7zPQDLO4qs5/vMidCHP1MFBpJ47GnId8vCW
wMfWgWefXkLiD0Ew/zYufCwDBtXAZe3TxVg1zZAKytGZZaZoZstO5oUzCteeuB0ti4/IKUyUxra4
3lYjlTzLxaYjS/8xX9AobWcgT5Zh/VefXhiXYVOSwHerzXtCrRetmvr4rq1zTyzYbZq6y2t8ZIBO
7E2cVArLKsY4xGfRtRiumWYmqrLqNJX9TdCNTPGGVg7VS1CIdcHievkjlHumaW7zYTzMSzq5ESpj
OuahQzkjhJzvQBjuNhl8632+5sFVPksdIyN58oFo6BVNfjIOOFmiJ4iUrbKOs341CNzAUpMbQ99s
0Hibk/iW/3pxt8KH3eN2+cWc13KqwUylPEyrLnkLyYOruX84fwBhNAQ0fXhnoCQ37URQpxgnehX2
SkqqMlWHTwJj8qz9+jzPyAQ5SoLRRkZsL8/N1ZWTzvnzC6nArRFhc1MtlkTS20mxRm1JyZJWpZ5m
rRJJInt7cWJfLi+Hw1kKfw4nlfVkJSQjB5SckhBk59+qXk7RLa136RkkjVoZm3l6bquoJaEZuIZu
thzAuV96zm4dJomqwKqqG2YUXNWAwHxlZzWioGPIFFMlTb3xKfXmPFnBlfDuXalZtV5J9J88qgcO
UpsM6mmatwLNxLbPwS8wQsHkAl8h+2CvRsvJWjwcIzaBEFsi9rSQhzyWWnPCUuLCzUekI8+n1Jst
jhZH/4zpjKMvE97DOrNCn7bjXtG8MWIa6sISazattyULQBtVct2viCgxuwv3cKVsXhb71wlX4mZw
jwRyzGIYrawMLaXlRjtVb5dnnxCb8SLXc5Gdpj0ln9Cr+dPWC9bAoAVEYFIrAb+gwXO+NX5fPE+i
Ycd/y4AF1SsFflrVdm/myehyWkJ8yxWIN2S0jGvTwrPOT4t8DLVE89RArGFguCp9ROGnoKIy9x8t
4fNcbPyPBAmDYoLgAuCEDV0gMXyxUyO3TZtAYBr2sDFcxunKNYQlOmFeMQ2OGQJrgS22Eb0rtkny
C1rO27t0Lr4q3ueTLJCUsWn+qckWIrPhrej7wR8Zn9Dbe1h1NeUz/M/ZmDp1wUDnQhHA03ZbpDmc
WahUqb6Mjss/VpwKQ9f4H5PNmBzhTMrS+/a87ZG7FgZNht5KiHIBBtoTF2xTQUIi83doGHqTxRJN
E88gvc7gFCrJnzoiQb6Wt/VtZpJRojnLfmldvzCIH1dQ7Y9HCON9NEySso4DUroBFmurHrZLrG0R
orAzekGwHS55UGobHSMeHis+U7EfP5MBFRHy8mlrqlT4SLPiQvn8jn6RpxiZS8oBZaS52+NxNsmS
5GyIoMurh9L0f63okHM/Fz2WhPczai+33iQjYUts5jiVf00Vit6rAKIxHWWEe0VdcHlJJiRChI/l
MKhgLM3Jo8T/swVEky/CQ25Jniim7URMB/BTqq8qKrVCc+TtSSvxYPf3EK9Adr+KXf3guYqOLyQd
MRYqH2NEoD6VxmYscU3Q3Y7AcP+GNYUKuLoa2F4lwnMoURgif2K2d1ACAqwzSIyoGw+NLdMJKJIB
lyjHhhz2PJIZidwna2BQesD4lM89QAifH/+SVlcz8Sw0TBovIHMWsXagzrFe8ohUlZmUEjm4lvu9
v0ziAwX9MVzEaiXIGzti17lr4oOYCxO6A6ohaarYW/rC4PD3vxIHPUGIvH/Xlqy1vOK1OUBP8/3E
Cd5JxclRUuo6/DHabnVy3u1dbr8Rtqi1BKS5nVsILW+/ASIVr4f/SIUDIwIlzkZmjqvG0sYt4uoK
yBqRmWQ9FCbjZMSaIV1NaegiMWXnlaSmowOU+bMRi/ClGJJ+P3C+cG7NErAvc2aztsPy7ZZhkmeA
5tnSvkgEMXp/kKqf4PLXN5XRfTfabYmeT8et5v0bEe34xyw3ZZ2FqvMN0WVaaQOAMgysoZCV1UzF
0yk=
`protect end_protected
