--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
M0mHrBCusukwBu5WhS44qeBn28rR4FoBB8c629DS0B0KGa2TnMJu0lAN/2ShbeBtL7UaxBSQluLg
Wc0NXXBUQ+oojjQwooVq5oIP2HHhnD1e5k+nNQOo4Fhyimu+8DhhdXkz+qOFWWOB4S2xeo4XmCul
VVep6LORaLlkthCPHaMGEgBBnIeZpNVIjDbcjQ7MbJQsOUN6GmoTAdjqo9hRz+997Jn+sTYnRD97
c4uHYZ0lHoGFlShVA2LkbwpsRlgKSMD/UASSR91zfmjwsErx+PH+iWcKRupkhgjJFkHp392MuTRY
lpvejybBeaxLmmyzW/O/D0/aA4EdOGycZOLPpw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="/Kr9JdfoOLh1q5c5Ow9dmHJtVbrYGrroZN5+K4b82W0="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
o4uvBeOPZnusBcpn/ORvtAdZ+o6jNBdeeIMv/kz6weJ2geRSrySQpcBYgQjrNCeutISbeznR/Nil
UTOOtSzOJ+eiabb6vqFvl9KPtp8yweWog7dTKjJUvIkVRfgFgyD5AMVryDmvDpMqRd4iKEMFNc1P
j9WOoAbcMyti8Pd5x3hKhLvcAOmcSQ3Istzgg2lok+rVKtfLO1tkLDCJSjykIjQB9bK8jyrLbY2T
sMZd6n76NKeYojiip9qYc9EDo/+/6+QgGwVbKd7wsPAHSVhYj/LjWbfAIpT4xw3rMY4Ugasuj0e4
Y4nH/4qM5iiVD6NvGQwYpRXkTNZHLBtkVWy/Cw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="W9mbNj2sQARow+r3UbX8ovD+hMXVC6VLbZaSZctx/oI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15504)
`protect data_block
pvd/4ghCxFfgOJpc5BSjNmB9hG1CEkGre//YRZ3NFaxpeS/OKZqXQPNCZiUlWJ4b7GtEkHRGoxlJ
0VwZy2/wLQm7yqvKZ938MuwwzAKylCofxc2+TRAMyPL5qp+OGZzLk991Ft8lkxi09fdTzGuipocA
f3vC175xFqvE+Yj36CdCuASg7cQVoSBbRYRksphngt4NlebVbML7utnAwNQtbnOpffprLxaJnQTm
t1SWvAqpJowsmNTPy2K55BNBj7GI302IX2XW1gJqvrneYyk1NGYFuBE3wEMdD+qVaVo1ezuyEYaE
isWjyAD9CtaiIG9qI56jmbBDL6eqApByFmwZYR6yiivSJLkJr5pH5IWS+RQmXkH3tEszYsBLAdPD
O+q3qIb7dN/ctYgQznvygGY2/EI9EvfYAZbwFqnsc+1cmyB1plU1/7mosDLdk1rVpgA/YJZ4/G6V
jYRyWD2uuOxhVO0rVIiVpAt/Xl/OewoTcEcMrX61Jyyk6k4DQkCs7v9bsM7RHWolkFN5rSzLd9P9
OktnsTzRMqUTUYCrfQACU0vxdQWuD8IgKVu+EdgVXdHKbW1Sq1o05dySUGoIVzC21Y+T9JecuTHl
KtjcPTwC8iAekx/NkmaXHzAqMOL5V8Zo9GA1j1axN0/kW9RsmhfxXar6+lfSYA2ApygM15Bwd6cL
tdwu9VTLAu7kpRem7MMMgsyQlcyymF8lOqg8usVEVf0wlMfUUcVHSX9Aq+ANiofvcMSzBTz7cgS9
XYyJwaWkMgWNHkjNI4svvCyPf5D5e7rAMvHjfecfVt9T3JriBEk+/4fGFV5fjTJC4CYxo7MGddKd
LojEbVJGleiRqdIoD3EX3IQi6FGG+tS9PH981fdPBSdoVPhTC7ExHAoutyaT53IoqHAwKEGBbLUq
D54KG4khFgnkQQE5cCO/PkIbZt2V5v2CXCzFxh7RrJ+249jmD/nh2DFQYsDB1eG5crA3jUVdDxeZ
3eau9LMoIbm3mEEIS2O/HXgrzDoS/8RUH+o2WqhGRy2jhebdNou0aK6V76NacaxBLL2/ucegI1Sh
ARsYNmYW3sO1AIMjDS43INAS26VvRuHwqpcnV+RzUkJy0fG0EiZNZAVzrIgC4NoSJQcN58E/DxJ+
ECVJ9Y8xZsPVS4pHHOi9jfVTPDoIDc3LtoRdFIDlEkZBDZlhdiiOAZr9tr0w6kUaH4wswwaU8nyq
qzufuxG8FkubUAv/WHJa+HKAMBiGPlhHSkdL8r5kyui9W27LQDYfRchH43FaQy/Y4g+zq75b8lX2
XOVOfgFmvJsdpzRIXuN+uIDyG8nWVDCWUdSZGVvaffdr6Fv0MKqOZF2L/uqTGbl81wohVgz/2EBO
ovc4supMQo/9e2uwOG7BxVIDNrQH50Pr+WnwgPM+0nuQhDKdlAyMMnbmyhT2kK06FAtpbdQO/Xrf
M3ytdQW0a2vzJ01FoKNs4qgJsreSbrDgfJXaWri2qm4eohIm6AYehgeMbVs8Vb7j/rlFmldSBtuX
a5BorSlTFr4jKfMY5SW/TwrIOfo3Ze/+Ts97w5G/gvDfG3vT8K+TtgVhd7jJk3E54nPldEaFhdGl
rhzTKlI6fZrvunpT+w9qyHj866ma2uc7j8BiTowrLwgtRrQW148BODceBGpWrOvngCNwEKkAhk89
fZCBklBAth8XVWB/haa+xUFYDNehiE8NLwmqmKfqR5a4podRYJnTdzuMkqRmgcIyBo2rQxhczsVR
CiMVrdSDnO7m6zL9ct+a/GdbkvirSIlTk9ZEYtDmYqqT0qk89EW0kZj6roBJSegxkhJB/pWwrqHE
gEJ4gFo3AeyEUefCEsgUU67sm55Di6+GzIU5plsofg2kLz0guqX6+vHX21CtgIUkO57tlAtVt7o0
hkJlXhsx9HZ7RKPV9Jj1/CeETVqJ/IF3j1/TeHM8zFuWdhmZ47j8wsj/dMhJv7AitxCJNxXaT/Zy
9AuCrRXupN6HHOoNZH4EI5E7ELIzyZKiB9SzutHG+XmSJ9NzuGc5k79HfZNmdC9f4wNypd5lm+kL
N0hOFqHZeFezvISG64FEXQqTnsZyufaZuu1kuSx2rQmltaBBtNI2uV5ExwQFsSTuiiSEk7eqpqyg
WF2WKxDZphzqhLS+VR8Ta8jEIb3aK8Q4HDOr03cdQ5yKFJuHXzCXHPHOaBLhXzUUulJ1zijwfYEj
l0pRooRzrykl8URRC1r6ikQTi1cn+bLgZQdewHH4mBBxsMrJRJSVlahp5SI+xdxQ80EITFQdwG0c
g9KqTMcXhyy6NOYdgt1cML1qxgIF8BkCkSKBio44LXTvJ6qtz6xE+Wqs6Wg1hG0UMz/hMC27vALb
gNKoqH59dmVVJ5lin2cD5NxDDkCloqrw3kXeYv3WekX1LEcZu3l+FZV56wR6KP024mNOi0i1W5uU
q7o5CmeXeqc70AXqAdCFj0h1/Iuo3VHP+qvKgRM9ITXLCDevgVZcWLdAIGyiZhxaAGZJWsF0ROmX
ZmuZxqiG/yceAGtGfWRN5Bxz3Xe0e3o0jt9AI7IFnhdJRksWCbqc1zmeP6Z+pgzYhbnFy3D8jve2
4uPMF9qy6uOzcQQOu24AoNzVb8B+ygiumrzF3gqyNRQVPZKwpgwai+nUQORF+JlSVt03xl/fw6JW
voG8SVBEN+EhhqYibAuvYM59Et6mXX6LRPVgZD5AA2TsWc25grkDx1KYnkRCOk4a+MyLNR5HxE8F
h+w+EJqnQW5+N2Oi9sSc0sixdEFMlVdYS86dRMe7XMWV6yLeuZjgia4L3YknpbaVYo7M2e9gUiqf
Yk5FfkDlSBaeJBLT1MlPsuxq3mauFrAyp1D3yOeapl1mJOm/8ZOsv7z/rDk+rDpTgKlnijICNXS/
PLYNqwGHukZrUXebl2TrJWubm6iPFCEgFZjD0ks59Hmb3cCx6nyqR9f9EVmu+SjXkvMZb5LNcSiK
HAlVxRmlGL9GchDG4vl+nKcS7ZMSGMXJfqRNP7b/SgEPGFMlkfrGiN49+8MW9XGIZqoQNqUqPLtg
PiUHpqN1guzZXmNJLddPy8Rg918GtEDppcY2bEMtk2xr9cksbRNdVUm9G/sQlNxKOM75ec4jWzo3
BSpBeVsNJlS5M8vCGzxmd1t3cSyPF7nDYfwxkVzLgQnf9NYzthBiREVHtyFCF8VCprpTGxcftczT
kmfsD79gwK6D7V0fq+tD65a75DQf5oRTpMghWqZIDqiVzkddXgRKl710ZFlPrc/xdHl7gfDHKnf0
fq6+sixveNmgvhLtwcmzWg3jucsPvj/rPx8mGk7etdT+6yNBEE+/giPjapaDOavtLcXeEq4UkegY
h9PLUIMZoc8PMCe/UNGNzDB9K4g0VW+AdL7lewczpG0tGPv/vz1cw7VmxKiDILxuovOGWLblQ3wC
FQO4UJ+dGcarzHK+PKDWXhiabkY1+jWBD6+Zv33C4HwKlu1rzszZSLt288pSdkkfPXYZ4HAm5OLM
uVLrCBgcRBdrBaXJK6/elFd66MrznuC6/rGog2B/4El6/fDva2eg6CjMWmtfIaWF8MrWXz2wDO3H
uV4fVhU7X9uOEUYx+PKH7NapKzvWHgTK61GegRJtsnvir9TbItG8IpXUJzoB1Nsr4D/YmASe5gJx
08eJe99lixN1UxcULHP87104iQOCbEgT3BTy5MNF3UI7Px6/MW79YCHpsl2rMowqKfUP6fkgw+yq
SR8PmiaaRDLwPZYEu6WraedzcWW1qaRmkT5fc/SddGTqQ0izNcjJ+tA8IHEQb5keEb2yk3h8NDsj
rGDQs9rP+ex6GSrVrfmIOUI6eSf8qGxjeSycrpMFlFBjTYCvfUvupimO+UHpfJzG8ChdjJpCmK7t
Jre8HEhzE2UYd6ISF+3dpVEWd1sQhwRPwYHOmpzX3JqJQOAqnyoAgS+L1dFraYym86Ra36H/gG8V
/VqHWTmBCau8ETyGhZlH4TCdZJCZiKILZ4K28EH2S6zYkzLS2gSqUTv0OemOBWzg+UDFRQ0bUq3n
AbRWIPckMTVB9QUUKueZDc6DeZGjf4iazsIQAkkanfcWyFSawapppMaOJlg4RT128NdXb6IRw9EN
dU6foGX740DYDSVW5zpI1us9C5fkftLX9TnPmI1bAIQf8fDqad+oyw9SBLUDVaIfOiMsAn9bFmD7
V6xjIO1zh4Ljo7Nmq1NNh7OEkIdRJwxVg5jKGxiwcQcMiGYI+LmipSLRh6ODmewNCaEornGUeY7s
JXYVFfmGZv9qssB++7+Sr9vN6HUfhS29MAips/v4NNaFiRDtUMFK2Sl3pwDj0abyEVR9eMi3NwnA
acuD8Mu/y7/G2lw0Im+OCP7MSZynpejCW/0+5y7YQmFj64caQWxp5OfmEhF6ErdavIUIx9n8C+fN
caONtS+0GAurtEJhanZi7frtwKbvPJ7N3gjic3GQ0BG7pUJiRUzhiMKe0z+2ZbHMOxzfzZztqfKK
2ylolv8vlvZhNGQUES8I4g6MWylgJpcEXaKfQC0x7G8uutBXrHkcA//FuZAt6Z2qjanRVtz1/ZGj
aH1gGyBXGiQ43wJmgAJvW/EHEXM9wmzc2AzhrBQPSvfR1Eglr4jNG7BXZjExQea05IoNUTBCaElp
tnlFOJF6OyEYSpp4Dzc3is6ge7a58OrUuXiPEiVeu1akYuRW9NViWZ4EtnZ56QTyBg+ouJC7Aowu
9AvFZQDMl1ZEvsTclobQFNIcHrNBRkKTnI4KBGyPOHzPV+hNR6SG5u/F3vBBjYIu2QuLRDygsGSq
7jNhVZDUf28rV7pmqh8aYHw087AkLHAuqEhXoNomxWojAm/YOQQyhL5n7ElCdJ2/DUpdwX75Bai0
+x0zdECnBDh1CahpH/U0EE5hh+x8fje4VLPOWdUwau5dyKn9BZIbaCbQ4Wd6Pp4xlh7u0KFiXLjM
P94KgpngwF6KpDcLUwltG1+Rn+C8L6/Upy+NcxvTbbqdcjHzrqv7ht4bNJZ4PAPTIiDzJkbCCfg5
o23hUxpgoiKcbPEFDRo9VguFBRHoq1h/4PSXy0kiwLDs0EH06IY5N7fsPNwbzQohP8lzFi3wjHOG
YHdKySC1F3mGWlBpK3JyZ/Xb9TtICJVaJR3TxaR4/OXotj+aOOEV8DTNAtGzMK+WOxaaFN0vlCq3
QPFdwgTCDX4JrkodanN7W1/1WJW7VNp1/yu1MUGm3HraegB9zpTVaHdm0fssxwrf+B2+gcQqvlxi
SR6auGGHU2sUk1ddKHTOxgM0Eyz29XHMf4Omk/b4tiAOp1eycoMGBkejimmiwvQMpUIhcl4marpw
5nnNysa22R/pXucVd4DhGkXdP+QeKXW8qtnP2IHOLmU14NntvtYVpdECT5BpSLU7sn7Me+NkT7HD
RN0NDsHwjrqYlvLh5+prx4UfNhyFeHUA+Mkfx5zH8apbzIlJci5auvZlS1XgbpI63CK1nCmQjp5Z
F+8uFVIMw9ZPUqoJR+ZbFm0pdqG8UvWk8iqTSbyYpf/nneDLEGuJ0kirH/7MpOpImfOTGn/bvsZ+
A3ajhHOafdsLfVQBhC/wE2EBurMmWIyj6xi8/7ddpu3Y45Uky57/PE7offm1Zi35A57FSq/t8a5u
m+g6Lvxl0b4upqBlVWYjRSxh5cyDaSrl1DdOehNgcEANih++Zb41RvseYfzM3/1OEAB+aFkZjggk
z072zZvrQJX76BlbtQIYF9u28aH6vKhklXBUxWxf/XZesZpqqW3XtD8f35NzFXrooVqW1FQoYZZw
3NZwCYQxXH/dxhXKMkNu3F0qG/hNhxVPigZTWe3UTlSrvCay5HwG8w4WCXZP4v9Vb/TVjHHKu8WK
Wj3jmHoRe66dQswddmx3FULSozTLmVC0+hlX6gSB4UBDUoFquoyE9HDJqVSwALSm1MjMpKSo/T03
xb15qkMZLghlPPbAaXf9A2Ht7dpXSdIORmRNyTVoK1qOx4/zN9Hqv1ApCxReXxowWUJTG9SgO6cZ
S5qyrEcvFcYXBlTzRnaydiFzfGuK2ttE0OA0184gYPVJ4TA7BRmXlkTfXe2i6NH44njKHMHiVh6u
g31WEaEJhJk1dLxm+1UgnKNotumAgG1rO8fSz4gFef+CXk5qTMpUyV7Tb5FN1Myc04ob1ckUy2lj
KU1Be2oK+UEaSumyC+O1Pnb8NzvttTkj9b6wPKI9iW7r2kGrGnpQyfe42LAdGrhV88MCpn43yRUE
Gxc8xre4rgRULBfz1+Wgxr1iQsgxUYYS/0XlNVrXyIuzwJXYH4qtmbdql4sZ8TN5/Ll4o599J8I+
T0mwWHlpvxliTdF+FWbeGBkULDmUGxsWoO2zO3DZD3AIXeMdrhvGih7HNY4zXqstAdAShkE0Q1U1
Hma3UwBgkoCfSDkn5Nk08QxJdveWtLcdh94eKrQVPBVL+QufSnee6My13328YmWTFNMb9kg/sSO5
+qKJy1evRwhZ/GO8cJwjTBSTVA+DwxssdUN4yiPucyIG/GZ8k/Y84/dg6Hs0wfkPEmuRTxV4opDk
f9N4Nzx66hOOnznhXTQUV/Npa9H5j9AWlc5qXF0iS7ZfF9WSmJNf4V0RAOW5Er2+I1PA7Yh9Z7Kj
W8Vs9aQGjW0EfmT3bDZPDVq1soa2MxqlDrE3ptjhH8YEHWMlbqYG12qlHnikxlM5TOKIqYH3DiWI
NBmNzxfHIA9TMewrKh7uLb/pj4Y6Ksw1WwifaFruSW9Ydyfu4CQBy5zfoaPFzOSs37WVqXEMKAC6
ZO1wyNbw0jGRrHoJDnhyMcU9bIoL9GotNDQ/1RQKYtIjebmYblXQ+S/xCIZgc77yUkw3P3uA2qrQ
Ia4a2RhiKGvI3OWoeSu4uAbI8C2V3Dqt2BPCrR50oN127Tw8FxUZ21dQipIeA6W6V4ESgMTw4EoB
4glu415t8bqUtfCJAN1YYsNHjvI3nYYW0tPu28+ME4peQAv7Hbb8TYxh/3w6FhZ4PnVWMJ08Xphy
HZ4+wRDV9kjVMxRLjAjsev/Vcn0V/ptDMqM+EWGQ8dGUiB0/TVpju9pOoWHKSTyAKWZJqn08C6Xk
Qhg4rtdsl25f4o1hAX+Tk1pO/Zyak7nbDbzdqEe3l58ZT73F8EXl7K/uMNyKbe5joErBgZPUoOXN
3Htu7ttLJFtZ2bg9XBlsJDxplCc2iqWT/LBjQEoomobaF0m+TyHTlj5DzOjAj6fEjVMZLUMuuqie
76vijA4RcC7Pja8ATxQlGiaYSc/WAWQERHhBO/DsMjxg/dkSbHZju8IuIvHYV4ChU7xLTrVIApcW
8lVqV1T6LssetS5P+qz3EMnURywlS/A1rirwOzQFjoxOPVrCYAVMibpKpNrRwUru4GRkGx7+eC58
TkWvPPpog4Zah715vg2QCF9PPcZhExGStW4S6u3OC+Ry5bBuF1gOt0kOSZlIkTvdphNzgA2Cl/6A
wf6QWpyDMA3WJUrUSVKZy5BdTNnruxLJ5EfUhE2A+CaWqqcK+CDKgokZA2dIkD1+HV7639y64767
Kc+7PPuTn1XLop/VjjcDGWGV82Bbyr7PkP0nGqVOJ5VoqwgZwE1+7i7945s//RWVWmwCmzH1gsqL
Gpj5GPvjm8ZmS6VN57TJAoyCKfIsAoh8o2LGEQdpXoePKnP+QwSPsgAlWHSoGZCPEEQqHa/Ec5Ea
jqZZD0hmCLIpj7AYfeZEZBxv+SZMFfTE+7jhsY1EE8p4hbpCrQBARlxw+hr4Wpu5XtTjHeegWIId
K5gou6IAVQK/vIvS64q0cZaKkRLENlnsqFy6OR/gOkUmCHf5rAK0rB6EcOJ58iaBWGHy4xhL+dtB
JxfglR+7YbCD3kc21PJrqyRMMv+aI9aqXmaDpZ6ItEvaSUravIkOEKp9FYZH/u6duGF4J/83Gg21
Mi3jO7ZKl+4StLh5N8Scb165ryPYccNQj3ruVNSwyiZmfJRoxBjcS8BfKoUM85OFAGVAIFiCJ7qa
Ky4nlT/Not1cAgnil/Xa86yzFw2lDAjHGfXRv10IL9RGNM+WVkgCba3xfjd4G/Npv8V4AzDKe/Mu
PYisSr8Kn/oPyntViD+vglJZDCDfQzYeE3NwpvkgtseGxohW76K4XZN/FvAFyobNXq79KA5O2zjg
e1mR4grGqbTAXeZnehv6l1hQtAadtzpr8dL/pEy5H+r31Zts2SzyKJ+J4gpjXJh8ViyOoclBLSac
tWYpuWCPW9hjZe/neumx26A/2Wm3VHlx1shOcErmekg+ytJYZ7gBdrSoEEEjxUxCHVXxS3MwtbSc
Wo9k3JMS/x+MtUbz0Ose/AFnY/T2ZWPIdEckI34w0heJNnZ/kpEwwg/6dnWjQwoIZ+AsiLki6XMA
nbveFfyfv24lH350r9sscpAFs3gQdT8EqrhIL8s5sZdne+z/qDtzaJcTSYOzYagjRdG1SaQF2/Bw
FpmEppfbsqnSIpf1O0vfr6AYAa0ALpGHtltipvQuN3fL1IzfTQFN6SxH8k00oHQFTMN/enNCbQa9
uWAiFnVvGlYICxnmvaoZGhHL5HFcKc1XxxsIsqy7/2EcxC5HoO/bqhrtllU+UKSfVUyrHa6wtYqB
tbnfPxccy3g4cjyghZKm5P4AWTEo2/uaqvivFA/xCmS7V4I3rJsxLKPTdvAVzufjZNyF19qdyWRP
OYuBX5PIRP4SXMqoKF+qlufy9dlWCc0RMJ5xiOniTtUt6ArRhRU7ru7RkB6yDhcfPyq0dyUBeuB3
3g9afaK52m4kFfhZJPFjx4Q1Cq65ErtHY/TaHc5zC0GAly19ZlqrXEtfGpcDxP41gXKVn+FI+/jp
SmmEmmXS1mqYYUot/EX/oDl7dwqxHijpR+4b3IIGERRjNDgQFQp7sZlZ5IPupr/u5lGaVZpIs9a1
34XZxz3wZmu6RK2fiC3rZqaqNbCUM3bMEVfOagKKRgSt6FpcDqK4tXlfdhMe2K31s2K2wfDPBlBf
rbM9TOKg601a2OYWUML68jsedFspEk+8+cEQhBnH2NrDyxRw5hyNcsMMOyzBARbeNjhPD5RqBE/8
Bc/0tecL0drVIF6XrVOpVso5ZmNydu123UaoCYPLdEJ0W1/WVEwABT5l9yfFmajQJp0eKz8qxkve
XNO0b4Qi2OCVY7ty/HIlO+f+GR9EzCLVpvE5k72JuY7Bofktc53i9yIqiEjpSFs4Lac9I0/K7Td4
xIx9WMjD7s3o/9KQrId2O8zI7BLRsG04B/u3uO3YE0lzoIk7VpXOk7zE1FJzc81tIxPcOTPUS7yP
IGolu4huG8XC2gR45UdY4g35acLjdY8KIiydc+IwSNBB4GvaVLCNMoq7OCmtfcaAseceGsaSQjJ8
btbQgQZIkDlHT8Vmsjfjq/bi/pe1MDR0AHOngZzkZ/NkOS7R9TnnH+QIPyjTnhzGIRb3VHFAFkWu
78se7ORKCdFh/yz02TZD6m1JpVNZdpJMELbyLRxYV09XfSmlz8KnvpAqueJ2SOYW+OF7iD74fHod
IhXIcCV1tUgQFfQwzJQHJPNLhxbwbmt55dQsIj8rNsb9JXY50BjusixkU5crjOFRZQSEz/Etzk+P
0z9ZO49tKykMQDn3LhzRWWt0xAQ8mN5048L/5yL5suPeFz5ppAOVxCjItzjcRSUISpVmLobZwFkf
I+17w7gI5mUJuL1qknHGWAbn+z5vAhoHUBMUMzF7YDNKwaPNzW/CDD8tA/jhnCkBSDSFthXJTHb9
D/6YIW7vXuarExyqS4gucFbu7hv9zTtthNaHTbqLFlllNclMj5RI0r+brnQBMzk+yvkxSQ1SkcBP
K67nzY41k6dEObNvk5ewsYfGcQt4rg37TvFCbo62FDU0xEaT+e5kMKHPU3OUEUIbXjGTs/eQ/HhV
mLqNHvcHA/6uzfYeTFjA3JKvkwGEJsRFDaOp+LRrvVWVFnT+jKjsTPB1B4BgZLYXHJtfctLfwZxz
zzLcPoNwMMAWRHWBWgywvKV3GdxTADSTE0oafPidW8aNFiDqxPs3LG83qykKtAKbiGNCVHaJGCoG
uPi1rtKv+q3yIZlJIorhvpnlSRxAhByf4kzfGp7BWqkmyXOqcUx+8+DeKxAoZWylpmjmGbFFFf+b
i8hVJ0jPGIXSDG895HUWZNW01mGqIlGckfuiTHOtr201dveS9aOKUTIitu/B3ZpyfPfedta/7S0y
QfIOPZvz9jB8EK4hImPIyrd47Ox4E8g/Ik6pN9H2w8mAOpu0Fm+05MRvFzSG25qgxTuJDNYANN5s
xUcehfpqNVyRI8VO7+pv1wTiMgOtnViAIz4lDH2QeK25yXQLAP9Sw7/PzRhcdW05kWb1xSENTOKP
ypGGs2THLnT5ZQEKgALM2IcP5bqLgJbdfTwvroom/BStdCvw5pR3C+10UISeQmjhXj+GwyFP8rBQ
ItVS+IJWx1wZFfa0XTwHLkESOLrJqnv2ZpjqCMnTqymDGoNu5V8T/2solDYCvIYqt5ieELWdG7Tt
h773OTGVAa2uQbJnWzVcVwrplzUfZfKQ/40nKHDNV6rjsg/nZ8f76j60Q5oPN6GIMh5yfkjmkpRq
uoYHj84BilUK6CGH3IjEZecaWYhPoW2U4I7WIrQDngAxAoDaFinps56LUSagD+rkijg5QVn+OUGx
NmiSCwxbdNQwEj0HMl42AJy6Uc1qfc9YWsScFx4wp/WV8yvmtdhXNoy59Q787pk0u+7fU0BUaQPU
XZJycg8tdiuFkJVYEJL3VNhWbjsRfKVAGCehVyA3y4Gf5wHaZt8JfoK1NjWUdCeDmakNy3/EHMfP
sVWKjNY1AX28Cgd5V+ikVeZaIdbKsPyYGhtxs+OMYEZga+xgKwZ71E1EsCX0oH6N8bB/7JDPJcm5
R8P4LDIVnyP47db025cHpc571zogqs6YKGp7b66TXcMImDmdkv8hUaC+Y6mrGcMUXD1pg/pKeEvJ
DRHgaD208GYlYvbSq1bMrCmjl/lj2OLSu8xvIEZVcByMqqr6Bz9bkhizaQ2oOuX5mhI+/U9Fkco2
dMyJwZOadBA1y0hMYClvBJZRdc64wHp5t2pFPgtn+HeT4zD/HJCMn1axjlpqoW7Y4sE3ZiPr+Nyq
Nh57SH/7jrsHkNxpJ6oShvmve0tvvG+YBFJPlOqwvCNbdq2S1SC7CydiBCLBRaouymIkYa1K9WGx
+SJuG4JNsKRhwLUiuweF3Iq2WM0gBH6139CIKA9PoTBX0p7KNVoN2llmN3QI1eb+wMize4Zu9CsE
WdnO0dMMXpFPN49mRJEj0nFesgQ9PcrLXNIQ47AoZk9ZQ1cXBZDG3iuU/kssRBunp1SWc7B4mshK
oEpMrFjcU7+tNsHpMNDc0Ya3I0IR+dpgMENVKA9tgPEwOp26lYvFgOcpRXpN0EvbX/+KpyPAn4bl
BuESPZUL+irrxx+0kgUSixhq+Dpycc8H6+BnylffPbSvUAuSXE839EduEySP6gom/nMe/YqZXUSD
gf69MmUTiX1C8hYpnMJ+kctEk0dTqzuztEylbqT5eoA9gi9z4fJzPG65i36cihm+AIKe1q26KJs5
BdzVmjXqJAGjP5fdco03mWwGhcj888XZnj42fyRx9NujuJBdBLC9ndCndAr2N/E+yyVcBPoVxdd2
qp1fLVYKfvijCX0Cf8Robv5ro9hf32sgjlII4J1DIcyuAAWhO4A5RyNtHnUCgobHZ+6zY1vNRQkQ
pTXeeTTKRIirk6QT1q2oCCk3a985REvFsJaGC8jfmzvn8x9mneDGROyVPAtHs9HyZQTCEQmnt2n9
nzY9NDgHiGlZUhMPhtKh9p4bFOrrR89uCs2sAjDyzG5KFS1hfV15avX9WoQm6SHqbm42k7q3sNls
brEZG3slYjriY2wEwYO8iqJaC1HgaI2iXcHteRPdfJffUwKn1WRKYWc1LpwDi+kD81qvzgDiNL4F
+rkfRSXm14qbZ+gz1NNLT+8OleVnl1fE8hHf6vwi5fHids++vwpTt0zUFvJdDNPxrxjr/96QB1Y9
7OsY1ud/XZ8SJkIOfwjHYOeSM2UG8WHSjqfFa1P4NEputslFwm6MCtlAtwuHAdbIe/2eLeSE6ne6
KWkDP/ZoCBg9WyVfnEeAlxjFWLP14MXL7t0uHxy0YBBniuHjSxdmpSDM+IFDXcjJ9IWq60oWtAOu
I2bHjwOHvbATDlzg1WJiscJyYzYPoK366m6ydvtWncQinsZq0EIacn2SOEN2ynaw03bPvyR48U70
XxKvMjKdft0fkEPAwRTP491LFiX4gdwj7XgjHp4opmTuHEs6i3wTYBLt3hn3wJpn0NHubMX3tHPH
hXJYT6/iH/qioZu94AmTx6rQcR0t/RpyywE0ypsdPoTFp1VdPpUKYTLyMZdmtS374wojRkbgWtJ1
G2k2Vo17DRGgCQ7kM4hIh2YEeBuV10kEwrigc9aZlDQc3dkdtJqIK7w9FmcFE7PV2dKRM2AfM2/r
mLm1siwpymEroGjK2kr7D7hccNIamUzHeQi6ER6M7QrIrVXb/Q5RCIwa4huXgiHWZzekqqo/vCEn
Zn0dgFkBJtjRzUYtcPVSmoaZzQe35WC+BkARUMP/6rPpBdAeUzmcopdxCeN5Y281zBU+BDXe6NzI
nPn/6tCkXsV8Oy9TyOvXXwJMViN2/x4OkvMZ+M0MzHSsTEeVZJKXPifHf2RTV0qJNNCRDVwYroBl
CuJVN2bn4pjD4jKevhabaN2caoBw5drrKp8AkxgYBR6eUVv/tALIhOHGu7Ajj9mK+2+Vld4ISGTv
kTpVDRUMTxRG0NPtoRhOmckBlSRN3rEhaxyHPM1OG0yXCgJD3nnvos1Ff6RtAKHKi4fvATCD7Y6z
WeRerJZCekWt4U/p3Zf00UEuA40gyVF5lqZTx7e9/DtajwJYIW24iIv9CIdgX3jGlGM22c8qI52s
xLcu5r6ioG1+PzlGqHTr/EhyTkINjS4rk5y8+b/Wfo6EkXiIa8vkhgYzTW+fufDJ27hjDf1QLpY6
QyCJGdFoA4xzndD8lBs7cFtQE72RpJxC52P9JqDzQMnhMcUPHNtvbpTv3OviqhmsrBTT9/fhl/iw
A0EFbdOC9F4KKea84eKqNSx8rotLmlKR5LnmLUr4H3dWhgVaGRwxCqLPXmQy/nxDHOP0t+81IL7C
hMOPtmUbSeyjhIm7n+H5+/Pj2Up+QYbcJoNOrbytwxvBo9hP+Wz57vrIRbOHLIcCuSAICQpu+Rsr
LhpbPm3Ih5vq3IuVZk0IG7vgV7HCfcKlBS6NOwNIM+L5i81v5pSvH2DZibjL82wr2cLTLAOET03v
GwJzjv5ho101vVacAwN+p+u9E9s8PzbsUODMd+EITANWUmGPXQkoMTeIg8iHhmBC4FJ2mfOI05eH
98XmvhUobp3/mhqHIJllmegpkyMVBJjavJpKpriMmHzUQa0WY5855tubxWDHd3GlCEP+c6aO/4YH
EOAAxezTtX5a10BPgDfMIeFezoxOrjZLpU5jMzbOrgBv9x+ze5GVNcNriVIBWgCBxFWFh3O/ZVr9
vkwAzO8KjrPqGymPUaR2UM73ofk6ybhiNoCdNMTM8x01575m9QzeTAatDd0SaXXLdlH9tEM4vmzF
sfQkROF4D0lIuABbSbxKVs+13wQtNCB+E7GlFAAxq7L+GcQVizpkg2vVuC2zU1XtexK5nSIkSBCs
48l3fqAFYc8bTcHWgX+So8Aj7VzVSnz9BUA6r/OOCXCtKzCSLKevkBEMOrv47B88t3PQGZ1joAZw
u0Kk7yUZ2KEka+01OrUjVOqzBlX27AAnpb7eTlzzHE+EHP6dF3/UBdJaxFtve8XpzIyosEL9ilTj
yREKbUdiAyBES4EStTdoAR5uYsm1YlxsXx6r7vjCGySkIYQPJfF5RnemOi4BAJqErBUstnB7aX+5
Ng98itJHpcqqTG4XE/Q+5AHZIieI7411Ch7wfJf51lCDWqa0Av7ZAvjUOmtRfQsGycsgjY487+h1
RSo8x2re0k8ca2o/sY4Z6tXVxlEx2s14BK+ml58N0wAX8jIVko04A0mztDPvNTcJhXwsYBiCLLGY
e9ORK9K1Yyxv+5PuqXiovKrWz5oP8EO/hlaCU33JyPKV9LiMbz95oOfVEKN1wlPOIzwae2GSD9uT
sGpmphLB2hKB5bzjw2ig6q5Tt0Kk/7dGwT+wvjdZyPam07Mcbg6MihQtGdU28o9piBZjAWG45ymW
pt4EIaXZrifScPH/89LjgwTg7ogxYTwhhPgS+air3RSgT9TpnFv2INO/WUTTRO3F0MuAb0oZHuTg
PAtuJQccT/AyHMf2CrDpE+FERQEVsUByngCW3wTxszXafIJCPKhf5fvMKn+3Sy1ycHvblGztBehM
FEngps3rm7pXVinaCTBSlYAvHRIebEdxGBEtydA+maMtYKdFoOJbIVuw2oW97/oFjQyrIurBETSR
CMbaAbFb9APdaOkO/lznaUzdssy586RpvFQw9B/FBa7adULTfZLxnxWbml935golWbBJ0kz45Rit
sECmxHCW/dyKWs1yJD1us8f88HqTyCirBkETr/m41NxizMX5AxanguybqiWT1De2sFMP1xHkXSa+
bh2JXqj/RCBrD1mpW6dveC7Gf3VMAwhE/ET0Nln0NSX7fcyLAfqyk4vrNTK51TyphYipvxtUgEq2
gOQd5lf4hvpNgE7uGrJOBA8lLi1Evu6Ab3dHtQaKLQ0mQ4X5kK4ZJ6MRv24s3XJSGIAzswnVFdY0
db7jxKKj4W9ZOeaU634A1yfJ4XBjViMX4cAl+BeEz7QatFlhoVUJqN+4epng5KStuY6DE/Q67nYL
0FDRzGtvHB/89ruF/VLg7Lme7O+kAZeHvpG/CFZKtI7Xxw5t1fQHcUJC7SFREZ0duDaEIW5p08qW
5LAFOwC5OmofIktaX0E7Vb1CzoSg+s/e9A3ktjMwxpz4kKHWc1VzDBErkJV4oBHfM9W9KgXdbFVx
vUKImViFIbQGP69g6SlWw6Z9o0o3tAp2XIhP6SLxpUWpPnCDEUHpxEotQqhtldz3QmIzFy3k8NRX
pIetbn1hZ887xbAx+emrW3AHJeeVfktKcNZk/ANT2knWBB+o1sgTE6naVUgFO4AeUx/22YUkVjSe
RbkG3zcFbsKEM13Z8V5zwCRTfsAc74KO3F0FDv65z3eP02+MFLj5my5Hsw+QDy/6zR7I/ZHHPXT5
sdZ2KA+WIh43LW7sHfqxKCiusA6scnLFCkeW6ow8A7HKu9XIIKsus/QINgNy8QY9TOGFNCCo0Hl0
In/M/4uuv17mu8hz64QZLNr7smInvV1+MCCsjf3xCuMCgmACXF9kCHMC2GoT7OFXwR37qV7RdpBD
I+0HHWOnzN7MNqbKd1f+Ustd0YFC32DPDHLt6ugpBnZzXdabiA6c3xRg2A15VmsPAbocJJOcHVFt
IOvqxnRTukswOZMcNdZkDVuXIh0hvZWAKQzNjUntLFsw1QtimWFbwDnsaQ3JNlCG9bgcogYEvBDN
wBkAhNqaE5paTMLmeOaE8oq1cTnLajVXsM0Fv/hYZxQPIy1TA8/pVZXqAIkusgANxZMlpnW3esJq
8BVQt4gmDH16zuLA4zLVZ6fRZL+NNhDj5qsKNcl27bBwQEbDOZtgCmb5GC4TBHKwOOZHlvdxa66i
zxoqHMCp2uPmGHb6tYRfGr9r0OEkYtdDDo6dSqZnGAxp+135sJbgMjvR/frVD+TjnHUvCfdcUVDp
BMC0IZ0S43mTu02W9vUXjtTiT5QTw3d78Wq3TlQzZhoXhpwXdjj9+p5VrL3bDirp7kE6EfqXCR4w
gUqMiIAM4KLRBhFy1qJ+4T2ZA5ZsEHGo5ecC28EnC/zvcjMRRTeaLwG84CYYI6vbPsqgXtsxeEvs
TiuwV40+yniaHwQG1oYIyvXXcy7kxxICLeBsXVrJ75QUjb2Wfv0syCw9KRiM0MO8fu3g1Y2vCRPc
FrPZ/3rSLtGgWu82jjfKiJqY10UxZ/ZQeF35JIPqqrMqqb9I5jJ674PYpG+7BYsDuntleARLRAqh
PtVSWyiSL8LjlpXdcrKP9NjF0AhzYA0Rz3MC3IWQd4ErbUNu/3RnWXmwhkyjVuecyNLEJM7P3bhN
xxyh+uxZt7mbTOzWoX3N+ACNzy1pUgjofUcLnmB0MjhtBEfOuJDhEgAgKz2XNUQOFUkUbKB2twHy
tkcGIt8FQp57h747pn2H2LrQaAIsOmVzlgD3DI8PBFP6mhizOEj3zR2uTeDzsqJt3qILliCuKV9f
ffas+CQhNz8/jnewC4y9Qn1BkzCz5+I07qe9QyBFhdQLEz0x9H40N44KhL0gDQVPj8wrqeDmcPXi
wVhzeXQVLAm+OPOD9X3J9P6Urd/OiUE2xVv7dqNBsdjfB3bLMfvqFKTuQxzNREtPTRF+6ib/HpxO
yh3UxivPK04SIWWuf5lEwgZuVejCdOcbouSkPTKFpq/2OQ/UnNiH1DuBZFcsDma8INmkEez+F9oW
16FbMRQMDzyKqvnR06Fua4GkBFKuRYW6jL30oOkfKsXfeG3SkWwWrMZw/pbbxbJ47F3Hlo1ZaSJb
gS+gj3xzfFUhWAyniJ01sq/elULCb6XgzCiDgmUHOHzhRUC6q6cJrVWUKq5SYboovku44tYXEq2c
frsZqND8Nva/fgBxHF5JjeapgH1v1X2eIut+YviJ/OTPI0Ks4cOAoLwY86NIf4aRXjd0QpHupH7e
NPCvuxvjFoNlGmZrKPA5bVU2fw7pAy+Fkwd6tlgc9xsXiI+ZD7N8KGsF7BYpvGlzP+6rrPn1Y/c0
mQTMiOIE5brimcnZJgdmRXB8+6xTCPZJ79npY5Za2YByOl0WUKZG7aJbF2kyGQTtJypWghVZKGfC
auFEhFIzyR0Ytm3jEvppvtfhd923l/+mTJvAmfKTACOzYsiXU31oJirstzvOxi92YRcu2cOOfgAW
+UXHkiyFvWnU+VzGinRIdc1bl/rOwZomzEv7DA2TA7uChPCcEizAO/CJznhqVsx6dvbhJMx0fhJh
je6cBkXOOgq+dUYvoLmd85Ek3alqmvkfyvC5U/SrMAJ8BHBzECYr7p1bDgNjdC+ddPYws7sSmqJn
lFnvwnU6ArzsO411nUacTT2YoBnL0TJUJKbhRJa2H0BDpGOHnHtWJvbJR/8whAdK0BLL9jDp1fDI
ThPJaE1j24pBdrajjwSjzxa7wK6bHsQTTFmnvT0rdkRqm6AAjOTO8ZTVU/Ne6xHRlrp4m3bH3xob
EuLhPCkDh9O/s+e7FAUBJSMdJe93cR/N0hFR1MWEjVyZxrP2jJ1rEFrMVfs5KacU5soU7fC23IPO
NGuFlzIpIl3XNygKOAj5pJtWOPeVHv/vKkb/FW4jVZ9/Zur+j9LQQQWo/pPetZycuARhBtVl5GO5
l1iSsYAYPIZuxBI0vivq9IRflNMEc/ByrPUs8FzcpnIEkLkr+uozrnvlfV6KH2geU8lP9nhz0hsz
BKvib+TOdIaRfj2y+7GY4NBFUrBBwATiST0VdVBUnuGUW9pZf4zTGZPRjv5dUoUQimSKa9I0OWzK
Abj5SiExBf7XvmQYV499Zi/o+4UtB8ab2Ok7kQY8rGcCGX9NzkarrnyYiic5tlJcEcT4MFR+RpSc
IJK1/sFggs2qo+R5uckeZQNkAinhT3A5edYrFD3JHxGq/T+Hrcmlw+RbGkVD2AYr790ERPFJMz2m
Y9hxo590c2Kx56C+s6R17J4YBj1s7/6yMU9Pik/C2MZ0ckQ2JfNx9nBzTeX4CPcwP+SRQaSIVPtj
HwMQKdS+JIWjpEiuz6r0eOg4Q/SvZKMJ3h25zvW0KOevfO4JpoMY52FeS6OSuAS9NvpwR7B1iegJ
jnhOiMyxbYRDdIldjUuYCj64M2gcR0RRytZqtejL07gtxWevWSV5LOAJLp+RAUknfMB6sr2Spbpc
wY6fa3TGQ1TvWOo+R/IAy1Ivi0qr5cR3iy/qdxPd7mbbGxfslpCBAqzAPGPC8FojXCZOHSBg7Uam
pOKqZuzrArEIdPYliEZJ8b1QVEtETAyB9lDCDMw3BuEKY46V8aH0uA9n7qrR4VhzFqRQAaouSIsv
ONHx4FDB/TSlHzXl8mvvEcgBJnYhaV8NmbAj7aQDg2LVWjhCOi1YoVRXO7U8daftPisAuSbLqY4m
ZB7YQUUerpyFnHxBbR0Aa14C8rIBTpfYkGbU6fUEGK5jLJM0JJHO9CD37N5wYCGsImIe44BizZRD
8DfvGWkRc5LzkBSZkpV5osKt4xvMQOOVfp+KO6gPfnY+IcILm3feL6Ojn+e5CWUBtT4JX14YW6+e
axMoY1Hht1mL0qqNMHC4SRmGhBe2vW/OCX7K9GUnf5XnycKFuccctpBls82VLkza7o2gWzt2FoFO
UeFdZGH4EY+UWf3kocBePIar3V5nHj2g4Mi/fkUUfKvW3eTipOHnbEYjuTVxmHjqzoQtozctcupj
X8PLVZErAosMoLAE1pLsSwQo5OmDSFqqZgTodvrbt1S2Vc5DvywI9Pc2M7oUwLeZ4d1ZXnMM6J78
8sObRB/ZKZeWFbOvwLSJ/eIzYSZ1XH9kZHjTPHgp6b3URPhjs2n7s1lGH4zPCLne3t9KIPjeY+wk
MhcXwonyKaHwm6QmOO1mX+AS8UsNkBp2HSvQ42uZBT9BqKb8aJdbgp/OUcbt9NPlrgnulmwmZ2UL
7YanjTAfzDgnFUTECi2v/VfXTexLsLS8yIDKrkxKx46zh9Fd7/JpX4AdvNuljtC1LrFTYYjbPDDa
O+t1XOsB/UV9Ya8B3by6opHAAZpU7q71uBm7dwUHgYS0dM7+qWt4q9LnO9KuUr5uipf1TViMOvFl
wWz+J+tU7NRfkqnbC6Dc4oLDa01nd8GfYPYjkz8rCLtjMp7/em/yTS4+aoDl/6iCZKgZDGceviZy
jj8lgoYLeDyyU91oHiey0RKsWhgRVSfc6ZcL1ChdsD0JBkFpSjwdxlVpOquENMPYfGu1baB9EkaR
aIsDIhpxIY5bgiodq5RJoiHylqKLbyNVtBdQwKaha7tmcl4jBaToy9DCNqMXFeWAs0XD1bESurD+
ODqglzCRbPADzHG67uedKwjQQUqFgSNcZtb4PWiERZ6bTximaqyjJ8CjXlcU56dqTn/et8j3h6JI
Dbnl/HK/LgK0rYnOjnjhROCagCdX9n45m2nnpGDIyr/S4rjM4wvxm1jey5DQ4xynXmkSK0QTT/ev
apPD2FZCFSqiSTsKlkrlm3TILrDT1T6bbR2vNljm/qoXccWLeGCuU3crOwSkwZ6oijD+CYEbrSdC
akLbPWmPeZK75O873ZlqdByS9H3KJBBQNIQ8jf6Bqf4B57j4VIf52OL7DAWyGiT8H9TgYzvqT4iP
R5MUlWXkxTfjQB8VuXGvkR0IgB2d/P91HnsZ0ZfTJR5dqhbQCixqy9EN+pif6H6XNgMCsVcbrg5+
ODb1z8Iu++uUGpbR7S9rzGVJMDEwQUXr0IPHuLNjOaRmv5XadBrl7KGdF806fUuiS4C7SMPaE4hc
JLEj2OuHtmTC9MI4SlIKYmfIaVt7OSbHJAGVhzra/oomF+Jn+djZTryX+qmUknD6MVQOIxgto9GP
CiuAydXZFVuiRYhfVaqnAYh9XWS3O7nsraxl+0PlXkPDGnsfikn6szW3X1gXa9dshvL7sS76GEUP
77grIlK5bmK3wyRYLiB7E5v7ZFAzuWINrRI0Qt9zmSQi4hf0afpSxqNNVmGD82YOM3NFVo36jTrV
vEe40cypIM1MjktzOheTpBdR5p7jRrNTaJVvVjrWvWvXTRFjkB14YABnPir+hXHlggiWASUS9zM7
ih2lesJ0pCnbM4bHDhc57+2tD9D3hRxxJbgPiqw92U71RHKOlok2bsT90HmZEkbiRbYk8YCXxUvm
/w8Hcxd0//3vQcE5kiUOXmnxnrvlYO+jH3MoNFBLJMnDrM0NxPF5/XH98wa3v6lTJ3GXKPlMTgjI
Ykcy7CeFfcBO45L85Pty5kpugcjgsZuy4mFSpuTSQn0CKSRKNdnLmxyfUMkDITo3rBcqpScx3jLN
JHkgafu3he1Z8bRHbeWvR8ZlLlhWeuu3LxM62adt2Nzs2eYjiXjrOkp2rc8cJpvCbTsWoLn5bHLe
k7DUf6NYjAlCijdc7lSr67PNR7GRm6XQSyaZYbUI2+pfUdEhj4a/c28ZJOfQLIQBynFHKvF3OJTX
XdNSvnQstM/TEKI6XE2zCBa7NuOuUNmVaLQIYC7W8Dd69DQbTVh502YUEIjuvGHidwRmyHhq6WZp
2c4lvNhXajm4QnupoToyvUBe4ZI5oqSsHKaL5jipgA0ks+iTBoBCH0PdWUc0/pyDZfnsLLG2gKRb
kwKndLBeZnSBa1lq5MDinsEwdLV/TuVH2PHuaOtoXcoM2abOxVguEjTeovjQBMkZ2Y2KId242xr5
EOdHwrTL7EcAi6jlUDuj6KdBVcKrGqfMmChRVvNPhBoe5i7SVZIa61oRBGs5OLj7I0VTV1zoD1LY
GHNqkmHcFKkv/B3vxQDyftGBjmHfIDj2dHIFzXKjLB23HQgC3B2e2pUXDTx0aJfRvSJxfj4AQI8/
w818hMQfumhT2yg6hdvz8ryvmfWgD42vHcr9gNN4UlySIlolsNmApY7QX6GMDjwjJCB3b37pZ6i1
`protect end_protected
