--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
R+EjBuaAZwNT2SbOdACpWvILPcmfQlBPxZkHskrTjsMR6Eyvn+dQSQ2Got46x/JLm6bzQ0zMZlHk
1O8krPrVQoi23tPACigzkeAIZTZw/lDvAbbDhhzXn6nmXhW6LMiGmu/BTPEdM1iyKXtBpXZKpkWc
kMiQk4at3YaMrl52LA32ndwV9VfI41L6pz691lIWkKpQQkPqP/FXNN7bpLIGurvKf2C9odoYvzxc
qTRBS/04a8QlQx8ttF6jf/SfEndyafM1UMf+e8HvN1XlMsOO7kJLCTWa7ZbuCpL0Egj6oZ1w3mrZ
mz9NRQCm+LSiYXE4JBGXD5DpU5TPC/g4lfjkkg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="/mNUt83PMMfNicOJgb9JFlatBfnIX+GdOMmFIBXBkTM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
MaerLpzRwV1RoxojIKl8a0sTX4kvtSFPg2/ni9KO6IktwyKsPYGUF6bSH+yn2vhDc4Knc8Y0yNyw
6Bazd1dZiX/IBnB+ZSazyN1cJ/gEJYNCgPMJCfg3Y9GT9XjclnoPcKxaBc6Qz2DspxIyNqFh9fLa
+d67kMLe/OvcnIV0XeAb3RguRxARFiSt8+UysJscQQTKu80ZHGh33IQOACUKLCCt9CNbkFdvLWyc
bVannjdrDe5G+D5aFsEhh9lQIk+IwfwgAUl8Aw0dA98mj7CICGn2jvG4OMUiUwavuslPP9P09nUa
4NhC2FZzXetCnnWTJ5KqfFOo+O6uakksre0xOg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="2GrkFdAk64cSQFwOKNtMMi1MCdes8sgUJwAfdh7rowM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40016)
`protect data_block
2mwKFFMLF3EnMh9NhJdpXjIwJzkPA99MLSrzLZm0b9NrwlvfDEApkPFeQKuDUOiPoh4zhcZEyEQ4
XAHr5OtabiQ8i7nyPRHbs3DHssjBHfLwgEGj27aYazllGcc18VAn6BeYhuJt6ZRQlkKM5CH2lG7k
E/Qf6f2mvLrzfqsl36xNLzXJ0sRRlLeFFpJ16PDtVq0G9nBBYA6TM7Gwyjeau5O0N0g88ZQ6/sBB
t5SHGwoEDxkoxnX4btZs5YRwgxqSIj9kuZEI5TbUIzf08wodZMVVpQ1JaNGKxC6NSM9IL+49k238
7BSNihY7r9v7v106snsgEHj8SXO32XD81ZofD4t3TMHrjm9t2s3tFDu6i19gfg4/DOMvKrX0+zDa
EpD370jrIgvPoSzEd6Mfuh3VvWFuINRsn91YsKDIOUGoCIPUhgnvNPq1NIsGR7SczYHM+CQXg9H2
xOPdIYmqZ+rm8Y5NYWy2dHEruCfp3bgQk/LJ2AUSEy2XQK/IToycN8pEyooi2ad6nscmXXoM19V5
MaBvRkt2AbtanGSeP1H2giDw5dscngjSdi9WbnFYN/gJN53z7bDxeMWn43Xncu1RiXxSigJXFc2Z
pDPZg4vTpHyZm1N3RSytVaG+0Zp07h7BCtObLjmNWvBcAyLide2LJbqfmY1+KlQ4+YsjsC7+DVr0
9lXFhoa+3rRM9MyQyNsydxnmTRruHpQlJmQLJFIDLJmfq2xTNzi5ocQph/rQycSTRlWNkk3aGlYI
ZpRML0BKOLmWTVlP33dtx7LT9mjSPAGGfsTXN+TkWIdaivnZ/8BvAAlpcTQ8lgjGz/T5yBSMSA1B
5+zWRWTYOYYF1kBtA0u1Osg4xGw2/BTCK9ge15gP04MTGqtUw/ZqGW2ylY2JpIFS9ieGbsMDrClD
/PsGtAMNyPnkQIrhdssI+W0S3zYZoPKI1zbt97sN7qkBzc4Emxr5RYA7KKd5IXZU5esJPmYdjqtG
nidMIFY1e5D6cK9lWbOdUL/PxBoGmDfPXFThPlstCFghvRw+KrIp/dLN4F85rhe4dnZ64xrwhQAD
hXV48O0ItBsREVHLaPUPwIc36OsJ7FGDJCKyEp0ebXgM21XkLAnX1Uc8eKv+sA7uF3UrkoT3NIkF
sqls8mVNJ7eGu7Oqe9Qr4uRNg5aASIMdm6Ix40JwiMwvtg2+R1W/fQufzt2WDnDC2Z2he4DfBJcA
J0c3Cy9A9SvY11tKORBizpuHWk/H6dYTPPNGx79lp3npEqcypoUVy1k55iTmUBbve+MGLW9j6XFY
Xm44nuvxljfRYifFFpzjjsDeXRgw2FApYHlp+9+RnPM777dvMat9A8D/Mho7gcsh/D1Zqqc4uLbQ
LR0U/WXDGiDFVNuRqei+tJqxxwvTYamw7XaO1NQbpgXF63wJ/OEgiJ3GEXUJTQHd+pA9vOKo0Xr+
8ZaS8mmQ3mNn5N09hVhunjkN04jjZEU/olDtx7enEDGJYDi7q/9B/xIy8+459if+Hxn13QWEt+oI
W8ssIdYCgXN4n2uIKp8apYLbCqXcqKhDjd65DMfz01V1dC+Z/ebajTuen1LHAbaoKVnY8/usAfNt
aavVQdfQ8rebH6/Akkt7oQJU+yUCDMGbT8OxwdT0wjbWLuG5XKMbiyedE2DMRxXBqUV9tUbTcZO6
KX7NWTlkpTXwqHuyKyN4gAJ/mD4tCD9+u40JuPxFpbkZyAsNAeUINhqa27dEQ7yB4TihjLBdOBiX
L0KCaU7g6250xk5ZlwYGiT5LJ6OO9+cG5GJ28EpdkWqXTHqVNjWpsrqlE9sU192cAqSm7WAz/4La
EG4v9mQOe9r9LZjyU5/u9ToLlkNWJQYhbr+BDh3mtgA52aM9Zj5Aq6uB7IVObaD8ViM5LCmtWJ6O
3lgZ1wdY0WUOnm/Y/zkNZ/T7OO89GlOMOoLtFp4n+aPoTX/u2h9B6vy8sEGSJlJReZqAI3/aRueV
9lfAUvhyyHgGAZBKImv4aQPXaZI1OZRc/eGaem76LSfKUli6gVGTjgyKCKccY6Ib+2UlfCMWPxbg
tuR/Z1FA+d5xnZq2hP0TADLQlXjHL/4DhkCi5FUQLZVpHGXxzqJF9/CkXM4XnytlOYqiDj5u5Ceg
VzNH3nR9iiu551pK36Ep2oL8XQj/IAA70wM5d+JEuHPcJMpC1Lv1PSq9Y6Vvfz16SZbCtI8GGHdT
NCEc0Bm5uf8uXqxcf8qZhYRoqyy//DAvIhq8E8n67WfWL2yLdpIf+A4ct+QHq5r/oiVDuwFUM/w3
OqLzK3vvMTVqXNrtVgZpx98kMAuy15JHpd/h0PkYj+Fn1uR93SnLoQzLO3RV71xPRH7a/VaAfsMz
KhMNN/QSfW3KsXemJVHgJpeQThHh99z3GGhta4dYgvEothZsjFqkjOD3H9QIO0XmUCG1UOcAdeQ9
OMbHhYwSiWVlXA6lDRrg8X1LWhJzFXl/v+rCIUY6kMpGNJc5xU2SaCZXMs+3e4r8kieMHSxvoM3+
yZ7MRVELG7KsJiNZWHV5GdclBBkRhpI/xz+SFX+paSoUdSe6/FJVmPscEAxegRETq5tRX012pszG
TVLmacg9UwKabShbSPgMsY39zyiWoEnY8MJOllMX3GVgF8L7md9RNjV1LtoknN1CPRq+MuvPri57
vud5xIAVgghLcHuNly5+JFZBPH7nIbtGM9PL+rqfdBP1XY11ddudv09uHkj5hnLOA6RJWb6S3zB3
UqXhox2HfuI4ksakiWbss4X6gJQkGHTcwDDfrxpgfxX2URfBQVKsXIBzus/EdLqMC1ZMKXY0WPhH
RiXFxz0hiEDowTGXZRT7gkQ16I3U22hAIcXc8wQV9hkDABQLJFASRB2f+0EORBIvHFEu1sUx8pek
noGQ52sxbl4k/pYWsFiRRH/C4VLo8VGQfGHmSiVJOozksUf8o10rhGE+HjB1fPXHNBecfLraKdFE
VnTtBx6QEIzLI/9G/eboSV890ZGTzU4JpXTuQYrnLJJFN27ofBAiDbYiN9t0ydIDzdNgQEHyXsid
1X5KKzxmoplHg1I4tw8LOc5/A0ELde91fEAV9wORmpSO/1b5xgVvYLdvi0UfJLdh4MuZSBTAa584
al/TygxTTmpR80QHr9nv3no2w+hL2uw1qsXsCzgG/uVyCdoC4T/i/mxXbkFmih7azQX06SutWnR9
D75SnGKyaJUFRrq0xQNM0//DA6NdFKgXth8slpxLIMCLNT6PLYwUlOLTsWku+gZOfifDTHGhspaK
AUXaJanN7lhVkIaYPzFzuL2iExJE6vwIyp+LL6EkIEwHtRWwlwusxFc1qadsL/P+5CSBIyvlI2KI
XFHn0zOs60EHgn+gh9Co6QXRsJ1V76ZGl+uwK8l1HVw4RMzBVrQL/K6MdXMwAX2VEVSNRgGOWIGp
cGBbm/x/BxjcMaEo+YuVgM5zn206YYo8sb5NpOaLO0Z4h8q/rSAHeEedFXY49dzA4Cg9TjLGJxv6
vNoyEi1NdysI7JrXoRJvAld7CCEg54hdknOFKVprqGD66SN1Zmq1b4SwEoF6JHdwNd2bfoa/zKmW
kijqI9W8RwcjBMUEoWEAbp+URX2GUIl7iC2IP86d6TqcMdmEmWA05t/VGBXxwZbDI/fEQj4QQQj+
jE/FylGK2J1v7ukcMUYXOqxZs3QTRon9fdlgnhvpX2p3w8NLFALxkQy+zrRhH/OL9YOY987VJANQ
a5KABw25RkrZvlpUfWhhIdEcwMxivq61VvML0aPZpe39XrmBytVfhITyOw+EC1NZoRnw6OVzVQI/
p1dnZDoyFHeEeLiDVEJURKxYod/Prlbqa/hROhePHJ0MWVT5UInTPv4MUW4ENLLJ068y8ZKpdj1B
dYhOHjsNPhu4c+2NPwKkH1RhuE8Da7BzthZ3AqDiOea3bDA8WhsEHAxNnlXTXRztPyYF7yHgMGyF
bVu7O1HjWgZoemEjEOBqGuq37fABfUNAgP9ss60k900SnqC6wryaN+tYLHl/vVAgeu3KlqTn7R8g
cv7d81ozN2unZzK9WBziflK746M4UTjtAqwElaTJoE+CfoJnfBgFWy7PRtv3DoByzBYRwV8kSx35
RnUsG98Q/N6k2zrZIHzR0986XSyszwjR2DgJGZfnLoW+1N5ZCzvUXx0+tGynTx4WXadwu/PfKaDz
2h8evSV4PlKGGXTCN/QJQNY+ORXlRpxCLGrbOwWmI6yrSm6klml4oC+GebRxrunGGWfxUX0+RJj+
3SZyYszqopjzmxyj/Y/sn+aknU4XGmPSOQH2tXV2by58J4CU9I3UX5L54onEuGa8mUlFR98dE19o
fYwVpUD6RSUU1I+mWyGylBjgQZ2181gg6x7lzSecxKdS+qsdNdIxfmyYJU4vk3CsiSqz3q/thBsA
ZAYCcV1thsEJ3Z3sZ+tzeqiDV3u8jVTVOIkBLQ/W0xUHapy/+1w3XSDxZ1LbNX2DOisWCGZaVrIQ
JZ0yEVT9KsMLwacUpOfho8eiqXh9sTUHMFX7LgbTpifBfzKOICFGJVB3Zc4FsHPekTXK8WkkVu/u
CzbqfJfK/pNKGFAg+O6WMN+fHtGOBhSQOwL6kuITPLLAmThj0yYOwLqVZeJzY4vNrDb61hXF8Z7f
ACzjs4UK+/6F1Blte2cHv+swNnSHZaUOh3ala68oxGyRx4JMNr45Ex2tygI/xMnHmgSaU6VwkEFc
rZxLBrvL4tzBk0YZqg+9i0IHzXKBPU+zqmTF0Ol09QAhC9WDNeeeYj7wUw7Lns16uXqPTd0kFi6I
WfpiX9HHG/OV8korJ+UQwXIKatULl5QtKTypjs5mtqZhAGIW9sKyl+wrMbkwUABZdw/+qHtf7eX3
9/hcCZCCbLd404P9iBcFf1wDAXQLt10nafzICbeIMowBOVN6o83Z0gsbOT7obJIyFQliTDoIECLN
FFtPX0Kpn4BhaWx3LYLCWSCcIC2/QJndZ1h2mrNDYsghaJplhUSvuY+xT8CBM5+M3pg+Ktnu5wtN
dnwuALFyeEfEIq1Q6iHD2O9c0r8a5O7qg18y85KlIJ3n2rtZv1prRVC6l7wS4e5SbVWuwAnSWOUn
bZu/Qi+fkOsKl4Jb1Rt84KYoxXzqwzEJ6JUpjmYcs9CN4mM3AiqDG9uUY+4caM1ZHdLnQSrrBsHG
qd9LTamRVym964lNwlybM7UnSII+7yYwFc39pMR71mnF9JiPlnc7r0y6YcrmARwNp6Soiql2pvC9
K20cHtoQdbIsq2ditblSWDU4JAjB6rx0oeRe+7H+PIVdjoopsQaExvjzsW8nsvtPMDQlwqHbPpHN
W8g953zAML2VCVQgWZjAmouNBg2v3kUwfcUVGW2cqyt+gTfI0jDJu8EJhNr1syjcybj/IeP+T8fb
YW+uAygwgq1nq8UKJ7j3u2SrutjTrr2/osaIULy5s7o2fm91N8mvktFIKgevz8A2socJtc055VSS
wDy3DZ4rWEg1FIa6aGiW/gMH/5MUCc7LsU1OApfchqqJMkfNXSV1m6q5ZsEDhpjEAjiOVECKukcO
/rxIw6bqO9k7JcVNJ85TvV2hoUWOUS5e6b/TfvenJBnBRfWlOADlL6QESefJWzPiom9erpMFQHB4
EOwY9NjRtm14mv73CVhRcVF9FkWE2AfAETjayESlGPiE1FDyJjJ4Nhs6QXlqq1HReDysvNs6CwLx
s9Jtxw3OJJhq967dE+/WswnnlUxiBweFSc2oNWKSzPERDAXUYPoLd8qoJOxlZkRKDmH9VHldGUx3
GIXyE4qHxNoiw4wgpSGdRtsgITPpQQCDDxv9q8GCsl2sRXZLzeYM9RO0ASbe8ERTXKHH8L7RyjHL
TzyLL4waXEkrLmcHIfmFBxHHxWr6YD1dSlv95QFC0Y6BhobuV0fcqPk1LWJ0GYDz/emsPfzhIcea
fo56gmD6gZWhY50vvAfcQPq5EF18vICm2CUlMeJ9QAPRWOEnu9im4F2Jw62jRb+AnwZOF4vWn/Bs
+UYA2uz+OBW6EyA415L7YpvGCDG+Q50XNxK65H8VdBkMyz71GURX+77pO0XFFM2FTbwag7IhXD8b
36DrY66QPijGLn/KU0ohV+0pcQ9rVEUPN04+WSgzoZk3LR1sWmZUIMUUhV5do/IDHVqA30dWFP7j
RMxQ6MMYHl3BaIcw3aRsCiddWhrf1LrjkiljIftBOyZMGrmtRNHOPtEFLmFHjKmkT9kP/cBNOaEi
AVgCJyBhK/znchMV0dU6bqM1pUNFEhu0hsVP99L/30fGe2PW2wBGEkX+olyfllOSKtph7QkOzkMs
NjXPfKzjWgKq8zbn4I3i8Dixu2GYnmWeogNRco6H59hGCkve0WppbdFCPXF0b6Tzp2uUG1CAUvIA
b/ISb1F6ynDy8Nc34zgzaFl0Pcg/kxj5ftcKTFqeY7b3lKvbUcd9EgDUeIaus7PFcph4nXaK+VTr
+NLHR+9+nxD4sX0tycP8COT9F87cBgQSoKkND/BQuzGurtamFJQEVkeCY/mUlh1BIzttiWfvt5yx
Lew61SWitdTOwirb/B9MOWZpcSWP0RwTRX7/lgLSEDQy8MGD2izIVqoFKv5cRL5JCMSu4J0PdaS5
JjGwfyhpL/xrfY9OmC//z1jN9NLIK82NLCc9IhjVaZs0c4kJ+2F2/THdCelR7fSpWcCpnI1AbZhX
AEEhZ6JE5O7IDS8u3b8y4SCVBzLDRakvbug4Mz1tp8MLzZfuYau9mGZSH+AFJdcKCPPprcFJ+7yQ
/caR8HVbYSU5ype/FdejrptvqmZXyLgTyOwqpamIWkLTfYLlfxMLAi41+hZ/E0L49MxWkEbCyWO7
Y0ihkOzflUjEx+yKJpWjiLOQDZblOQ+RNj0ZDdolEHZGzjGFHkgW6gLEHTsO0jK95c3PqnV/5TEx
ro8tJ40mGBm9gpGScV/pgivIIV2TSKG1G4gYcBIBdnzNd3MamEszfIj7ZHuOs6SpkCNL49NwUwH3
C8IiCz0py/vOYIUNdxQp3W7unM8p9fKMi4R7GGFVSRRfuibDeT+PuqykK+VBoEo4owIVwYLetNfm
7YNg8pmU7gmN1f+k7Lp1J1qdG1uHg4WXfuBvCCiEKc9TWymCxTkSvj6IxjOSr+oAxp3f3ZsPAq4f
kP0GSRHCC4Eyc9PDCjZDwvUW23UULLbR1UdIQW+tM+h4zKyOtr/jyDxN4MELx0x/dx3pYs0COEed
6WsXGlS6hGC523YtB1IVr4Xb/pTGTmtRBDYFVoaYHkTo0RQZz5J3lfI5Oi1lW+ZRbhXaLEAA0p5R
9P0dwgpJgYl0aCOV5/p98IpdhL/71aemoR40hvUm9nb6BcwwDXtbz5z/OlyuRhOPVSwhm8b5CEHI
RMDF+05aZbGjHJtbqs/gbWAFMvTons+IEF6mU8Ni4nssN4tT26gf11p0Q9XNljwTF9z37FqIy3St
BM9fSkBGgUqoDFCL0k9zC7DFs1EMFFDfn24eFqvHa6SRPRQQdbBkIpuu5tDsuHpHldsyUajcKpMc
bApBHV9AORWQXWr2JOq8FISnfsFPluzFmREeX35qNK+It5Wmm8eff5Ppzh4C749jUSxdpuaUDOqY
hN+03b25pcNXu/YKNxBrgR62oQZk6uPtIwkQJV8ovATWGN+thnMQtkAOFRHVdbRRItySCFPWi5dQ
01OC7fvhV2zAQwxpMLGRAp9p2y3t7frwPA/Buw7no0l8PTFSEds35zeEoLPOlJ1WTP/AArOGBI4s
98KLCQpHoobEJRBriSH1ILewIuy+fXzIEOQN3tPq+B033gvnrmCEYRn9h8wdper8fNWzZ8/HSoz4
5DgWsdkKOZutsxI82EB6Nz0a/lvavSlROJ44+neufI6BmG9W5e8MXUGBxrafrkhhy4e17FBMVz6i
UWqxpwAQZrZMivWkKdqpuYHUKsL+C6sM/mE5eGOObyt0OCJcSlrB8JGLRuNJwO4+FuAqzEOgrL/g
W4PQE7zhpu6ApYTn1PSrBQAZSGN6fdHjql9zHQCMZY6zH1wHRE/oRfDMTkEyvX0pxmsYvQ5YF065
JJ3U3iV5cnCbsEU3r7F3YPRIS9E0DI3wQjKKyv5bIMXT/XMV1wLBlLGre7a3m4AWJ4yswGAZ0sK1
ZV9rI06cUjeTHiJ8l0ClTmk/A9Y4aQWn/a3U15mQThiFuq4I1sqivvuuUjQwv5b56sULrNu26gZH
BQXL4zUrjUEf292vcTHxDPxA7oF0D+Oh0mO4n8xAs9x4kfoegGncK6VEQZ1wKz5oxfDWS48XeHJ9
gNkp4BkRCj8ImfcBZxmos6BnnCxcabfAt9OokzLUodYySxBo4N+dmB2mobmQDP3VNF6YByXo93fi
aReWUn3f5PN1XpPJPo2Cy7Gp9EZWi4PgpUwkuTEbsP2hjQqXlBWcIxYhUUqsIR8HUSnZwf6XjUWl
qNJmrtB+G+rA5llV+LMpF9P1D1bqy7HPp78K0+jjFStdmXhX2DZLRTVJgHVaeXUQ8G2VmsnfqTmq
N6XKqqsnRRPIJgC2wQHvBcykl23pxA6LjaiIdouINzIW5XsDVfKVC2vnny8cw4/JJhwQ+j3eDfOt
TtRoOrjtbC9BzOww1X/NxhLknYLxcUELdpxLHZSR3diKxO9Fd6NHygcP9bs9g2tXxG8tutN5V/6D
T/A7W0nqmI335u89h6Zh3htKhVUlWQZqyJXlHNXzpwTeEKqAfw63eJNGCet0wNUd0V55x1vHXZN4
6Lod6mNN+xDvdSgLEc6LQZV1KyISN5wnzyzgiGErEesE3ukFpxUsvLOGMhcGwInxIMdXmPsiIN71
QJJiV+poBCfku5XjUw+VnAAXUF9xpk9DXx2QGB+YyLdaj+hThZo8oYCXnrVe0Jn82zaNomdUsmOy
P/ZB/fRWCJH68AIkZkbvUvJHn/VtRKypasZEfd3ssvaq83GU/8VaOnikBmQLpxKUvkQCL/qVyQ14
Lx0YnQDDjTjLc1q8BIPcZaifi/cwWfZyV2bsap71n1sjGDKUGPshGGsQ1k2NWIuinW6xwW2sOslm
hlrC83u5g+rzROFxME2y3zdVFmmo+zqLM8zw5Eki5uZM4cGW8mLsnlvrSdl/Rle/qeSVVZ68Jp8/
9Z6Pv+VM68noR5oYgVPYxSDm6hD/ImBJrOoCJCiDK9/sjYcj9S00oGFdZL7lRiaA7r+CQ65DAomd
qo7+qVS9zSfhMcW3v4dFIInGz2RGA+rTZ7tvXyQ8iuBFQgLoTJwbKEHx87ZgFBV1J2vEk/d4WBM1
KFY/giSZ5PkmpXUPf7Jdbz9T+PT5RZng6fiaFuhc7829+TaKYl3p2sVxLJYT5Bj3z7OHUhU9Nhve
mBD9CEkeblhgzZVHUEiC6G69ttzvRuBY4BXIhQXMEMcoMWdvlZhcD+cIexEns9mYC7GBlL2bx1YN
hNbWzFXk3P9nXeNvS3OlgPZOVZiW5sMpsZobCMTYGsTP5B6EJOKPWqgNbOgxG8IHOOmXss8qfl4o
isTGqSp1U/9EiN+C3xWF69tvGjI7pxhCWFxMp1B4AGS6ypxdaPuqEO95biikU/HPny/WO63OC5S8
rEV1xkFByNAMTXUw5PeyggEwE8WZ8uDF6Q1ouN6DHEtlGZwnnT/0sUw+645di0nqmz/FSKznXGr1
PGWGMJSQd5lTmav4csFBU06bVhn8a5bxy4gRtPHsz4UzFk7kl7RdOvkePdOk0Vv5M8uZ45YeSIPA
H3tuCYSuFQjaPkiYOu6b9UTphrz/rOKBFZfKxA9bTtxZGC7E7zcvf+Bw2okTsYHnktyOtOeEXP2B
YCh6hSCmJdO9m2lnYq1ZE8uLtFxezN9UOlwNQqDd2XGDASCBZseRh3CYRpvF5hiZ7vKm14Rjgm5M
ZrCpbks45v42E8BKMXVwBhe9aKgTcU9X5CJHTQH+lLfC85LfJBAfac267qMBoTMfN9gzxKTRgYAn
arc69IoIAm/UkLILUPC04HuYkhkRYNT9ekQX0lTfgI4s/v+d9UTPFuj2RV7wiLXkvNOcfCuHgdOB
ZPuaTfm8OnH6JngBStm0Qi1zl9dqs5N5chZ8rKu3GfLxN66MACh7Fgdzz00/3c+6cDf+CfVT/w3b
vuQPMUHbILuZSQ28UeUXNL55dWcqfv65AU301poBsQljOWEAFnXWwpP9arAz9aLXCjXfoPddOpQv
EGAa0JNu5wMKlFpHqIq0ceFiwe8v1/YLQ9PUkSIcNqFylkcce5PoIsphAp4HK5G+aR8XcMacKug2
YmtffEjA6euU7ONIJzlmONXAie0JCodnqCCVRXdZPZmwsJ8YAq0hM0TZQAh3r1MTBeJfGThSxhsI
CRSERGm3SUaNSQGyVYjgtR+IAb/TKJbwqKazAYK2igvT45PA8QLVMEHlmwQZwY0Gy4/NPP8v28u6
xZ3QkGP/xc2UWy+o1dVbkhlaTnK5O/m92BXKOHEqh0MfOWtJhExXUh+FkphV2+3mhSaOJkmUs25c
P5R99JZXzMVQkNfkEsoQRKZEebbfdApBe+VOtByAHP3x0EWNiFcPv7foj/qa9c4iu39P28Nsyg1p
hp/4SmalbaIyXtuKZ9A0/vcf/GxmrfATYCJo7jhUzyNy7LKRWgb4rn3XQARORKcEfNYU05w8E2ze
Y7oX4jM8ASmFma6pjvp3qECQOKoUXdmYyixZo82FDpVJAVmnDfzZrucyq+NCBVAJJVBaW8QdVrPQ
3idh79zV25mh5iTzY/onvBrvWc77SypUKxNjykpBDNZuc6zuRqz6g+M20NtNZZ4aeIbNuP7W7Mn3
0JLeN5/5j0kb+cy5gHcWKy4tAwA9NEUK2VVBKwPPGDYYtPGPeF0B30OkeoRLk/gq1iaQSOwHYO+D
KTdwHVqPCOTvDLp/Q714vh0swAXjMbklmBtkdMwyqGg5Uwr6Fe1wcq4jlCkPHe1GdWWtTcVZpo5D
WyzkAqQFODMU6fefqtZgC/ZF1qeprnj1YKVb74Vm6+CnEoRQimyB7Plyg+muixX49q1vXTuGrBGF
tSZruMvTCodDaRbudEYBlHtIwp8TL87GmFKThmgPGULBJi8ee2P8zSNy9Ek/ea1+eRSYEoayOEMt
fQC65fltvw4rt+bYGYJrbFSixbrX2bxBWAW9b5xzooT3SdL/ZwDa1BxIb6LJlZvrWkEzaLguh7ha
4Bt9Wfo3KedbyZoqgq/jeM2S1GNFfH1ez9htrTg7nHCw2cuxBvWsGPlkl2JaDTYZ2Vf2eVpkRCFW
ZInq7QVtDeKYesvfpSfiaOg76srnDF7W5NLwVcAYF1Hxz+8HImXvnrdyAAs4TMoJUW6wtIjYoq2H
5GyyD0BrzEJVGmSCHEMpqCnXjzNrXzuYcztvIkpV+T6P5uzufmV3oHVH3FnuXsskuYq9028ikMgN
MfINRRDV6OqL8zuyPK8qE87koFZaE9+Wbz9lvmBEXSnExcx2HPM4MG+YRCfmSOGN5ZOxvWIS248z
4ZwcJAqyBP2NddeLjitD3YddefKGEQBKmpR9XDSRU6EmDcBaJjtczgUbnHzxNSPIAlo9aYyc2TtB
kzpFoK7mjD3o1LNj7CA6J5AoVYYezx/pK3lZlVPWm3oZS2iavzJKmZJ0LN24Ni3zlkuJKD6PzZNY
BAY30P9kiC4+gcC4CGtux/jYU6AuZmUq54/o8rUwfYGYZSMaVNzet36Dug3s5eOUnQ39ScyOMeRA
/W8iWhDyIwgr3V8X5BAMc0O3cPLkAjoIWzBKOEfAeQaxNp4U/0JFwh+P68hr7MInT9mvCAwS2COb
HsfSi8CdN0dgPSv0/mDGJyCzMPqoInVMuAAdjRzCE1CJa1KjS41AllqAhC27Erj2jkc/0fWpNkDs
1oi32S7Np+ErN8Tfm7J/16awLaqOwTUwO4vyq+DRRBj1/fvrUSTKFm6FQwGBObpIPA96YBIUuEp4
u5RQO9Rvxaxm3UIn99vjIVfYP4va4BNHB+u0TBWDqzYkTwzHJT9tEF2tAUQaNcy7YQ2scNvnrO5u
vQ4QAY12/5HINTHFnUaGXCv3qtXt8o16rPjjihy2iQ96rlGo+e5RyfrQps5s3vqYvcIqYmwmpXhw
Dz8JOOPC6naBaW4Qn2lF1kSsu9FJEzCFW9cOBEViZpWG+oNONg8dKLHiXVNlyQRIP52v/+wxGp7F
PPIc7DUn8CQlazRaNMToeuES3KSOEdRKSKLrEiriKQyhqDpWygQ5sCH0x8JBeYO177fov2EfUuxY
hOv8xVZYZAwu1cYuQSWPrDJoM6zZNVK39dT7z+EF4eYi6slINrA1QuLzJ7qpdt4ggDmsMpAotU2I
P2zo+PaGsqkmWC6zly9aaZZbo7MwJBk0tvpsZuLAytO1lAazjSOBO6v0K6k0OMVbve1zwT1ABxe3
lASNx0k7QTx5VAsetktBm0//UcWQ8CwPlNe9ZOWr0bWTM/w1Go2WOB9ffpJjzrgilwOymdNqW9vn
Va2Bdk9V1sY/VK8IRpO61VFyrYJB9Kkepbt3iU83fwGDTPmHakyuEB0ydPevjFvP8PEC4xHQsgbt
gNo3tBp6uExYr/Eo2gAV4dLsJTWppxQHdDKTjpkI8/3zJVvbsGXHCVjxvRF5RIi5RrZmiW+eFWkf
OTJb4yCiA7Ti6t1tnqPnqfDZ7rqfkvuQ03O3pU7e5Vkb6nfCyN4ZR8c8fwu7ZzWlQ5la+yDCee3x
X62CLpgm3KLa7PcF4uVcQ2pm+0Vu29m7ZuNdwJXx31wSpHF6sxRbGOBUpmNAh/5ij/zphzKWq2+W
Smu4KztDhfBO1acsSd7Muql3ZwZm2I5gSpHlgi+K76ACcFvpPyu9BOapnBldz3RvOMGMpx75i4NK
ctVQGguKCIYo0o0dVHYJgJnzyPYe6CCSG1qIh1KZMT9IHCAOuKJNO+fVFziXf5p+EzPsBIde6eKc
3AtqK5s2xsmHmayaxUrpGJdJ6Bx36xzkv1Ne5d6KaVcDnHfM855OfodiGqpWvfg8mIJI23ff6dle
HZfTd8VyAdsmOgA0wDOD0CRohIEeSQIEPVXRwAmy4OsesS7IxtKTdq1HlI429rEFOqR1EbT9RAGU
mOsWSkRLoFfVnDa/mLWX6tLT5FvK+UTbIikHUXSTb3yBFDndFIwhod/nmJOLa6iGoQUirtJGOP8U
ak+lxExuxGFSL7/5/wj1p9joyoPEO5PJdPtQO55GKhajInCMZTVhx/fIohPgdMfXTPLQa6E8Y363
Uw+WBWMcpPNJZQg/a/M4YmQhl5m7BFIrFOGa7GqNA68eJNjJUEbYt7rBEPjvSXwQMtd1VzBVoyY1
gj1VNXXrWSUzVRmtQq6cIKZnM3Sl4CsSCJiV8/XLJ4m8rcXYO9ufOBTd1tWi0hmK/OnwRkKq6Hcc
vPyGGArsEAYTS+JzpGQLpPOSfwcHSdvYtTl2HF8MI+tznFm5YPlaEseS2pkbkyOe2tXs06sEu+an
ABMVkoLEJOZNhoBk+/WXUPDfJmksP6CpNbaMhce4nqfKXctbujrlz41W+5xywgQRQcg1XgPpWkjp
tqlyDgPeg3fcQ0tU1EqURpt8mUbZrZEPFOlQ/CDL9bfBHu1cMZEa7y3HpHmWV+ugBP42qmdz3J1v
TRs4Qa9IXOP34f16Q2tmVHq1Xfo6/mj44xhdnnxC9BgbS+qJDJEfoE3kZH/4IqfVlaApoqjSgjD5
lzkmuy+6Skz6eafDUjUcemKDrVPPhtePp6+6N05fmIOexpsavrla9wo5LiMDDT4wg/l2JObmuo1I
q24OuyHvplLvIjEB0l7FQukTuby48UVEGSaH2K3RBkWiSWB81Pq7XZ4Ribnsqw3uKa3se0u0Wub2
A05z9tx/H1wRJodPByFb191bs4bAMZvtunN0Fr4fnkcVsmoh5XwzkJmtVGs3RzJyMLbyea+cdD/L
COQxBC1iZMGbNBRzf+u8t5ZShAIFO4Nfgoa5cI4dXdjhCF7ydO0CYmRVrJ9WBTotK+M7EI+YN6pK
ISxHfnbCiNXWQZEIEx0WEI0UPpFEGuflDpdzO4yaFLnEYyAL6bDhZ24oWhYOmZxMU8s2Lq7LlCBe
MfPm3E37hbFyc3NNwZ96YdcIZMkaYX+qDILr6c7kaAhTzsyQ8A8o/Ne0SZUwDOCsXzToDbGIbPNS
ur8IQ4o/Y0yShHZv1UkBqK79B3JIzMV5S+99fCH/i17Yv0tU3U7N6zfN7++HcCRbabp/50x7ahrz
fJ2RVikWKQUgyNEdvU8pWOKJNFqHcOS8S8B+t8ZUEbemeee1iK2ioRIpSa3ELWB2xKmt1XUOlMNO
0Jz7ji3KFRvfPFQF37X2/1FurwVGYA8dCsAqpwQuKw94+WSaJI+riUjtw7Xlq6qm5xqdtkm/x7Yb
UELvyPCbfQfvax9qATIWglo2hcFCH1gl4wzafNSB4FHuMZvnZ34vqD21elZv6yvhLP38hRSu4MHS
nQsvhLwSnv+F1O75zvOu2+5KA+fbxEiYrX4Tjey5tu0/Mi8uIyUvnXwDa/DwnJ/Slqh2N8wC3mZv
pg+HdFO4swdeR7oQHPyd/iLdhgx1/g9R8nSTbVshayGnzIkUNJ6Q4xWxq3t/ORMux3pnaxsNp8OS
CqZ9cGwCCVHJMGhat5mJJmGk9UfSvGu3izG0OR5ZT9e8mDEe66YzJGTDlkTjk/+4+BenoffZ7SIa
jluG5uoOOj1PcLkGJyWdJdkdu5hZvMdDveqY4VZtXL/2PpY6Y+16dNP0xLtpIdhVUtJszlcNDBJW
XUpb/mLxT4py70FKDX3SpM/4ZJGrtsM29iWM7FdZDS4HrIt4YR+rS28Olj+XJD/oWzGxCi9BQ0UO
8R14w6IhvoqGzeEg4MCJSjirbL+HkspCCnGay752kfhLRqzCRHl0yk5MndYGEh8kVS6VPtjOGHA8
25+5AXXkiz8mgfw02qsSfpH4vQ9zausCCvFYqBEIUzFVuaZeq6NTLvrWxcG5t5q3UjiQinyS0CGS
UmAgtwB328uFZDjqyAXC91URbq/b8UnoBsjMAmF75COgkN9140lh0e/ORWWPBdDMJDMvsZR2X5fv
5eh1u/ZjPQAP+LmtYw2dULpVTDht3QWQ4MUZxatWD1C07k+dlWHLPvKM7xIYM/yRDRtuuEq5+reE
GSkYRSfPcWuyAi3wydWbrSYQueFgppbDq4+epyfu52hbOgr3V2uIb4443KmuDjyBKkXf2XaMdVnD
gyDL46lDUxNPKDF8YLNr1d8JMsMId5hmWmKB6Df14sL5AsH6GonZHJLcjL2gTW9WJ9qeKCpQxtPQ
nUX6qbWbjWS4FkQPFtXm9FqWB8CeDgbSD1jG8HnTxxzdVcjTyDfMTE2Zvrqlpzbr21mSi61NmKiv
p3lWzC4Zz9xUyGF4h/9Xb22R5VNB5iCcQs3Z4SoKXJnGpBM7YEXB5yJmn2xm/3tqMrtOG+GYSC6z
vEVfWFFU8kif3IoTCyLg8EdzQiLk4f0iJ+W6EU47EhWNgkiMYpKMIKRY9rhtYAKzdbsholOT8TMv
nqJbQugVBCzo1S5bhhjMD8VOaLTND+Sfka43Ng8N4Ip39am7Wk16r/mpUNALIeVVthagy3tCt7/r
/qmUMZPAiTn4oo8Q/xyorM5QoS3qh8fGwdm3k0s7VgTYrgpcYuGMpZlBuak5nLl3Gc/cdHIP7CnQ
hQSGhzSUq5wYb0u4yi6vWZQAw5bQvf/SgVfAC1/t4ILNnrUUvi+IET9dzi1qAZEob/AUaEGzCSrH
5SGnPsVXsSPtwgcFq0oksv03EA0drtz5gXA4DmLvuqi8Kgd34S99Vld0OiCda6tcQs2+YulBT1Mv
MP1/J3nZeSk/lDF4MqHCQlqDnjkYgzhOx4zWOVqb57knpNKT1h/HspVA0JDqfFjzOFYyxwvjN9b1
IKERQ0NjxRIQN34GUdjpAldt8u4cqfRycMiRI6mn1ui/4k+X+HfK2Hy7K/qBGmXSN5HB6Zcet0IZ
QSwGuoZL86iu3u7Mx8d97Qx3IUQjJbTQ5igtFBv7nMyjpXc/0YmGwgQP03oyK7wenzdh32TpD/aC
jm4EOYWFKVvgO4wOgHlqUit7g7caa5Z5oipsQQUeq6O3c5K8mVt+8xojXxTSPLAFNLXojIQWFfOX
4bopF3Du8DcBRWjDcaByUDpMj/cXtzc3GZ/YFHItcm5rzZg/jae/e+Raa7xDJm05CUsBBTyEgx/y
NRO2ZmFQ1Cd6panvpnWQwOkYU+RdetQAff0t00Rje3yvfd1x7Y1njS8FwHEWderyzVsRqtl+3EXT
tIsT7TftOVDSModqQZFW4m12q+mTDClikCbIN+CvR2BV3hwU5rio+p7DEAk/nPcxTXJdNoM4oUek
+eMlphZpNw3JBn6kioo6HfvEuFCzyK7doAhJRNqaayiT4bienk7H8bQdrgc2tSikpgZCYe7W0kFd
SXx+yBzI2iH7A4PXsRFtVJrZ+k/W+B3jrsGJMc2s88V23jMEK+oNxUr6iKH0BUwCKtRtloK2CbMc
/ekLdgCYwO2jlmaTRbSKADeGXIrntjq3s3jTdURXMs3Xi477J88/YfqRtCebHXNOIun8WPSCEq/2
ifyzg7ddkYET9uV13Zj4AkgRflOdujmysJ+d+YCQNjsF1hRiVyZ3RAFhri0mllrSbqN6uy1OkMof
dUWLBo+vDtAwLt5qfY/jD0DWtEyZUYjvTyCbdMdlECXwvXkBmajqZdmOGzvufADc7dDSwsmUXaAj
XqFbcpatrqeKINXt0qFCCjGyiUtFibtiyjNBQN9f+UNEJSBfcbDfF+QqNufrNgiDR/Ff7yK0/Jwe
S8NpU6tN/f1HkRcI0Uk2UWQLeX1r6jT+RHkeZ/iW5etuhvwizOosLoa54XO9tEZnaKcUSL6s3u2X
TdyhmnJXVUPYiJT/2NOgm96xsJ6vDc9+9CM7YpOjLc07BExhc5cEVlgTeOObdLG+BYcuPYnxMH0b
+x7l2ZXE29HU5qiXvqDfpbipNF/pQH1zC1S9a6FkCeRm1SiLAB3bjOQjpWHdlcSg5IgxOFOOQQZV
ZWzrSMtqxclXuLC5Ix91JIAmNMydQmw2gtOVl4AHnb02PwHcBtGnsZrumsXxbzm/+86hNEbIxqnC
adRTQw/aiVKMxEhY3962u6bMlQXq+bEwNKKwAQlJ3u+6TZnnIpZ/CmDmVFN+ttgVOSOC/udjWSCt
w3sl6IsjlIbWcNjC0SUrabSxobiBshSYcBcEODSD9cpJd10wbzkNPyuQWJP4g+ulrgDS7XX6kvOS
9ilUnWeE1O3JC53x94v6M0iZ0kB4O5WuegeZOIXcTnOMp862rtKlc1wJtNWctnEev8Y78hYais6/
cWPMNsoLHm806As0m1D02D+9ym76Mc7NzYqA+g1XEGI0J6pxevHEAysTDBBawgqbFIhxS+eWRMqw
63618zpOJuM7bagWaDeZROlMsajGzI3bRA8P0NeXD+2FiRNpW0RODxOUHQvv8KrKVKmy+M3/enU8
QcSJ8tKcpS9xEV2dEt6Z8MWhqc0br0NltefN3iyd21lzLGV0mXUhbiiTPWF/mWMQUSgRqWXeyCce
775M3pmpXJsKAzSw0CFu55rDMVsYjiQUN7RQGCNHuM/icPLr+all9SCj3wWyYPxuq3MGmJ2XHPFm
Tmv03ybMX+4BoHWnSUjHm55ya7z5952POuXkjognoc1Fl+kA47n3CeB55Xf3K2OjF+ObV/DTsJPd
tEc1DEHP6RZygT2mNQgBuFhOwZYtbMGhvoqOr6Z7KLJ1uBTGwuYJk/747H4FkRR2pUNhp0ea3awA
WKKRdvUk45GX723cgwdyTwOHp4LDgexr9M7Q3eufn7up+karG6yEEYGeuihJujc/YZkoj2fhF6p+
/6oUGSS+xEEku9Lf9idB1vCL0wdsBfuBS3azm0KwK4DDfwPHN+/FyNhfqXZcDipy1aErdC0/RYdd
yzx5pj6jSztFBrXOFjdAIoVefZoKJET9Kuy//gbNLcIML9evkJqLVezwkg8SSxyCi1V+QSRRGklU
otamNLnZewfZu8VZSX1e3ccVtBxPu68PVhlLJ4jPaBVeu6rDfmoFsE92nVhTyak3cr0E0KLaKVfv
CR83fUMyhSeWMsEtZlPXgbuxHVCgvGEDBarTIkW2dpZqRa+uFes10bY7Ui0a0dM4sWiHS674grfc
olJ8ESF19LDN0HAnoGfXxdzWmUiMF3LeSrxNK0DDKimrtEwhNiAYWSKpzqDW61OBdInHrouxPzu4
D19kBZLWas68XduZXEKrfiCRFuL+h2ROu62/0mK4PgLT/c/pqqONgXHrU91pb7tInY82Yzquw9/a
On4EzCMm3hncWr1Hj7GVM462WEnXpANnjVhN6xNQHNGH6sT47KOEGOiW8JrxaQWArIXFug0A106h
5wgedzDkmYHoWwLvdQaBJYoKSiDNQH2FdQVeQV/Z2s4cnWXBz3mBIqjdvXTkfQ2xEWoNCZbmL9K6
71UpOXT99tAO08sjU1aJe/mSqLmRV++S8wiS9gWjGb3DAZ5wOk/cwuJbRck8Ma86MaAYKWfb/1Lp
rX6OFd2/HuNvKfJVl+z/ztPFjcHUr4IG2PnpWY82byk/UedMJ+S/9PajhLKjDsg3jZMr6D4nKQ/Z
osbA4EzX7bR6nkyjBsW2dftEq2TblPSCJMAxBnjW2u3SrPpVjeUvBbFvUxPNBpNIiNdjNmfjdiUZ
5aUbsh6HEsLTYSQDNtsUUNx0C1W5lkLRNuD/vhoyX8fWWCa9zk3ToUJUQM/mqWTqcAc/lMQZkJsI
CIuW8OuOWNj/P/j875RwTMH1UPpEJ3GqPIDSpeWenI765iJyt5vrw8ByqXIxDqmaflkt6Q++NMom
P9Fc7K+BJK8nxq0gU7BT7OOkAMwYRqxCYOUBQ/7q6dj+1/V/JetqXDBa6KdAzzqJMCp4bHhSYrvg
Qs1+VwSE1R5NXuKEOJnjSwO7QZ+SuIsBn2rdekm7mPS7ubWNjbIw8kdPyOwV6KmwX95fzGTYaCVu
LKBoyJKqQGYjh3IwXblqHKsUWqkdrCpGGYQVi9r3KXQ4cZ1w7EJxz0PocV7P7CuK7qQnuLBAERt/
Hz+j/bbYk+qU6jbbtF9dfc6tgJeF+YuJhdwUf5QFHrvmq+spB/y+ulggYp/b18MnXz922m8A7Zn2
2n+/HbnPmsOh+mNFePc+nUJ26tKo2xUIy8Vv6JChXQc0O5t6wusotzZy3OYsimnYVh3gKLhz7Fk4
FgMaKFhzBf6s5DfRuwrrJUFU2qWPTL/i3N9aewZ+pedddRr4fHQ5Zeln6tBbYrm0RzOl6MTRHxec
odMln7s5hrAIgEcRNI8b5s1n6d1OL8x7bZx3Rr+/1WHTGUeKbISSzZXTqfRcoEzwBtxjtLorc7G+
CEf4S7NFhj63yBWROqClJ1zD67BATl37ISwJAloWCZmK2fKI9Xw4mMoJ8Rexgm3StOXY3zYeVEy3
kRQ367cUzAQ3TJxJz3TFv6wo6BntzPb+fdrZObaiGsiw40Qy0s8Mb/EhYqVo/VRb1fNCQhkjvD0+
RMrpdX4AI6DA8I/u/g9kpb8ikQOvK2xumCRVTdRzgNbvKdJ9BfLTqqOusJc8MO2ZSCrHcyBWpqMg
Y5c0b8Btuq+qZj+0k3hEyzMp5HXpNoCZkiDz+oYneyh4jU9448jfvgN3PmozxLFDeaROs9v2qaqi
Ust74Q50XN2s9TnAhtiw+LqaYIVL4uIUCn0kQaKDq3uFwAzYoTTEkOzig8blKyzxvmUN+FongfDo
IWFPYDRvSb7xrITwW2zaMMXRKmTXLLw/j0gYnCqpF71jJl6va7PExEjlSWOeKCHF4eDAPjRUB4IZ
CPYqmZ0/ZnCaI9pQm+pvyDvQk1UEfekDoonaCtcCnA6LeLCatdXhXwmV5FC7nN2ysE8tZC+V8CLi
uj2lcRTCAC/5TbCaWzLiGSjRuFpgIFjFSWsYXR214jP45g+fTEYHs/6Ga78QOrgsaYJvV4trPg4F
CS5VJZ05lr/ngy20XhHy88Kk6+fbguGbzIcs/lDTZhdFciV46kcLhBzi3mOAZU+jOkPy06WFIsMi
xF8WEmhFp7c+5RjyqVR80iHon9WeKMVAivrsu75/RuD5/C5OGORwazTz9NYIYo66BYcffmdIYp7N
w68ZOdn8wNC3FonBtgMrxbf8/FLhz8GdVYB/CLzBQBrhq2g2EGoyzMn1iLJV5xMzqfxWegqUHxPl
2lcAzlqqNn+MwBvWf6sLIXyckRsHe+aMLD4YbVcmgwAAeDqcWW8Kwyuhu+hGPgs3hp6iv63fJu/n
+QzO0IZadD/8FUI+EnjzTE49RbRDlcTEvpJY7SKb6S02wNY5/KZ8sevWm3XWFeY+HGnJG0vVSmPr
X1HDajvP3ycwTKkPCB4Qud+JX0O63qnKOYp0N/h0jKb8jNiLwERiZYNx+wTPDOvCvxdYry+VHG55
87LUWJ1Syh6Lgs0XPMg7vrLEtaBEdfkjBPpJsn6wWUrm91rWM9rOmEBoad3NpBcbZ+odIephrWSS
r8Ni6FGHcI76ufDUku4cPALw2ktLQ1faGgxVQ0iaRBotHAziZ9T6b8+YCUYD5jIX7oomrO4whbSx
cgQ8o4uO1KGat69xkEKQTJ2LID1SRdSHcFWDxvKDIJi22B5rUe6KMaKZ31vTjUcPATjLQvgl298K
fdufo5wHcQQPNZass+ENq+IcRi4cIJ91Cht8eLcuLQVQd/N5CNeQaqjROsKfKs1JJt7jgz0oCTQx
B55T7Ns0HYfFllTSjxvLZfdYK61csQlf0vQz5mWFko3yTl6sZibRz6gtF8Er1orinVPVfvuszuQT
4Uy9GbH7B0Kiu2Xvc3Sj4j0gS6YqwmzMCbW3Ha8Tp8ARNx3RwoM2EYaVkslnCftthM7rwW8xwCTk
xEZBQDmeQc22uLz4qvxoq4PqEIUobHF+rOYZuDcO9/DmR6DS8wc9vxEnpFMZf69H60qA1ug5XYEj
Mj9CajHEaiLXzX0/FiE3jIpuzrS8DCzvJoku7UaJHGrR+UiNDYgWRqQlauPOKTi62pzCq1d/o0D0
Qp/yOynhLwDt89okT/jGKegrc7/WASxnKeXsziEcPXFnDQ/I8cjrh2vA2ztCGEByAxHNJKIx+eRv
aoxEuCzEbjui4R6e6nddHvEs8U/TjV1WjTLjH5+qmyne09r1ZjdC859hPagCpwOERznYIqpRHACK
3IhdbLXfmP/irkyRoW0lkJ3JuEImuNF15cAbbk9rckFEeSYP4IqPI8KN0LsYeVNBxanBVaRLJ2Ah
K8lfIr0ioRREyDTcaHtXebhhHXhkJMOf9J3mQ8EMIoFUyT6kQJjhFiT1sonXDaaJYyM/lp0Zj1jx
/5koirtlsz5hXdBoHeMQds9JWJU3iLjIobCf42so9AerS+K41g3hus1OTcvFKbf2mqpTQFBj/Ekr
kXeR8KY4FAC82bzXDf+O35FU9A35wiOElgjiPEJWD5Lm5np0pWYd/LW8KT8dvOmFYzmUHIFyzIp4
pGt8wyKEb/pywyrPHScOrC9oNUspW0sCsHlzmTI3ELM16m7gw7O76bKVGeOdefLm4XS7fV3ySK+J
5LrqMEeW9fypnZl7sulUx9qreyZVOMWOkrz9d3buM9rZOnSIoA3hOKnu9Zi/q6RQpr+682MebMi/
O4Srpvq1dFwHev6T8U97fSTJSt61WB55HHUhpcQluVdjYffO/f2rjydtDH6KkHqzSH0yPF0cbKYC
aEZ5EHcpbl62euSA6HTb2mtm9eNLttjTcogEja6E06kAP9QuIl5mRdJimCvqXcVO6ZXTWUbf46sE
zmEs7TwvsT9VCCX/9kIivNCHJDc7jXpotqbOSHw9IFyLrU8h41LPPItuk3tRKLhTWOZDjBNwfnhf
fxhF3xDiOoD6ZEYIMnF/zcXu6HGY9oLmu1VWGLlrlMXyK66EFeWoBr0Az401iMoqp8UDeUiStwro
JeYVnDiW1BuPxtAUHULL2RUQXaY6WDMkijh1cIlomri/yFai4h0mOqrq0YXL8hEDgeIe44cdhnK1
7/gye3uRwxKOxUTXOzVNum9KYEB3fFX+b8FVN7LwBIJE2/KTxe9gYW87R3raXYb/NhjtnwHTniNw
ohcsfKSj/wh7DxZME0oibuSOiqgdO4hhKU2vBqnH3X5dAfjQUWeClU9MY7qM+69Qa5N8JHJ3UDzJ
UA+R4aYIz93SzWnR4CW1UVYT4k60XKeKFmcE4dA5ZKSm2uQQ1uxicU8uFYfUZRAe+WFGjt0MmfnF
WGIXq9FAdqFE1BRmGxNbDVQe3/shQ6iZ+cc/TnnL73CW2wBNkKXWE/Cdps2UinECxvXgGG8svwny
UKhQxGNiaN/nZk24pXxrUtinK86SdRQ3GS1DpKR8uKD1uGaA6pZk2oWtqhS5vTGuDUE80UVOaYU6
FaCU+E0kZNsKvNSW0EipG+mi9TWSxsQ3L/9qlqMB0Uk4dY6zUbmS7Kx9ixuOTL59hlwftSfF/676
UTDJJDeASiK1K0qAtsvkWD0x7WZWy2R7qvWWbEi7cI/YjVWr7pqu27PmqpWSR1uC+Ab6OmPaqxv2
0hLuLMTu2aPhtJ7bDJKWvaZ/Gr1XH6peovod85e10nGPtgGpJJk64qEKlxIThP/T4zCFzabhgH+a
t69AQ+4SdoGjlp8QfoxUVK1uw+R+v9x1a05oB2+V0RKgXXEdp9gYS7bZx4wMHbMVpJ4m8SE8PjIB
Eej5NKib9BsKnga3h6K22PdgSUe35U5o424UWnFgDWt4NwJi8rc8I7P9b3Zx0tL33KKdmImtERpN
b82nk+nTZF9Wa12L/C2fn7excP4Kl1xz1VED47G2c1bKojDFP62RRi87NtGOQ+a6RZYD6JBMV1eo
2QlF8G+jL/V4SVfxM6Cb15uQrVl9dNywHVGguClDomWGcff4jkTUuR2XG8aqvZDeUACBCPYqLAWx
4amMIaa/t9oBxuAavaVdTxsWgBXbAz+Iq+juz2Wn5FjrAMJ7TryvPsBYDz0/XmSqf60RCxbpHfam
6ajMjI25rTK38Y37/5Rw/snJhqzZUI+9siRO1dpjGX7rTBZPUKuZEu9/D+CPvAfYLhVc98jjRgWh
8MKmXkX+LZe6S+Y25ZTgnHEjN6zB9ZnsMNg54nlOY/zXxdYSESETBdqcjKIUyHZhKEgd9LZ1ZQMD
HWOia9OJ0o4ZGyOlqnG5UJkQCUJSNpZwcXwKE6Jg2O10C39LgGzG2aj/lEr2BV3P/pjmfgkz3a8q
GoPhE8bm9PL3Jplt0r96egExohuo6FLyu5YL8Yb4aZP2EExOpU1PdmxJ3sEbgIuG/5evKfvg4OD5
M3bj4GU0UNyQ4TmkR1oFsefJhW5Kdz8GXur+OHh2Od0gmUl25JsT22m1aCRe0WAxwtxTdtddsYJ/
FZ3bk0Dio967XxnBmmBN41mhW6J9JcyUGMlqrPjdTPV1F01glOBDuGd+jiw1bo7XrRuHdSeHJoB6
l7NOoHczv7HTCEJpoErb7AvmjkVOEpfYqShIvzbKm5JB5FpOZE7qRwIh4PvdqiH6p1BPQfnheS/m
HTRuC5xXKu9YEH1klwrZ0NvWpgXVRXQW4ILkTQvWalCDLeBG5F9gvCgYrG+o7VBEnJjYcEw3P8HX
MIe2Ku3AjKOJu+TQphwhKHMRlO3zbYN5Nc3wpJk318b1WhxMG4rDc9SAAKHuBQ8F1dl2JdRNiNQu
gS+O9arIGJ0Cd+37/l1IfZLYrRq0CRaGZUXy8aKQBFXsjIJG4I3ckTHx1f/XLvCf2x9i+A+3sxdY
HzRZEojmB3sWNsxbTOpLhSNUc0e/BXF7nRSGltTN9yXvDLDOuj0hDs6IVbGUGPWA3QFtgmqkHf0c
I4Gs1G3CMUsbNf0vR8BlN55KqBUOpThU4b28tdcKV1zvlQjpoyUnhWubQkNrPgbsZDx9Y7bnPOq+
MA/c129QzVj3nR1ySlLuxtSPcXwzWh1h4iUDCchVaS3xCar1YkFyo7QPE/g/UxnseFF5f2Aacin0
kHf99WFsmuQXtT6ZfJGQI+j9j4ppuGFOmpDararN2dtU3yCSTVXUfGSn6B3dA0XXXrWoamEmVZEy
qo8TpkUQuvlN5BnHL/7DUBccqJhH9O+VzcPocmZo5dn9QgGxfLG8KH24t4KsoSyKBKewJvPM6EC9
dDZNKtHmXEVQPdZurhnaPycwa0g5lvOc3PdFLFhT09P7P0R301A13tJsKrmwiFU3+RlSGfoORHIp
84aclDSeDI1aKDuCOzPLVd1zOFXT783v0ABzuJFSfYWIu4nFMRKYRUzcJOp7H+I9WsCM5uShvbWz
x8SoWa5phyhoOXtKsq2BjwTEPKXS6crsXsL34beJNvi2eRXFVt5Ydk6IbP0CZnP3Qy9LvUMnz4ip
IM1YkS3kuwaTVca9+yRdpsSSjXRXyYj1RwMPxkbEvHW6B2GiGH5cYmnFWFj2taCyJR5FdaGMg4rf
PkiURhRAqpPD2mCzwGLpNKG+7zpDNnmPZaOtFsEJ2gEgvK0HuHzGqVqNX3/irVKFuTyOKvnAIaR6
nnzHdXY/WeVdkQYutdNFKD9j04dKW59fghPviW32LpnlDbgvkHce5hIMg5FRaNLayMfzON8HCjSk
28DjDWvxfMU/AjlSl04UBIL+mOjB94rx9NiyN85cfjLtigzLys3N5RfWvQ931WAtKvLmZG1QlrD7
x7uVAst0dU924yZ8ppcGcE6YFBgaVvtRI28zu7O85huWxyig15r1bzIGZTUDo+CQZ/vxRgBlC+1x
k3WTI3kxkFR6DC9JCtDGcICPpCgpPBlvtyO6sPnNr9rDF5pwSf5YrOLcGEDRyGSjLaU01ZKUtnKC
Zijn9bdR4Jw/3OdLw9HaHQKqR2uOWqwB9vaungRlH8J/k6f5d+oWjAAdADet1yo17BQqGDBnXt9T
fTwnLHYs7KNclOZykXGX9AeNuCymnuCQ0y5DPx5sTaERk7DnH40hdB5tRSwoBzvI5ureRKp8p23a
uccIRKS3r2WG9ePaYZ5LLQrTY9/MLEu2TeKdFszg9Yhy42tssv72dk4TZVyi7RN8stHBfabUxC9u
Jt81YvpIMdIAjMXaZ2el2Noc+cAcikzHB2UM8Xugl+bquj97BZ38o77gBoBMdt/tKz2BTz7/nfWj
G0OLqEyDslDDEJUPTPOGNiiGH9LVDUpOhLaHLTYYZd40A2Atk9kxnOoh1mQRPqShqpMqgKuoo3E1
hdfgNTcPgo0q4p4dGN56xuHnMApEOei/DBCIUl3YIsjaApX1gVLtxtnmm2fsq+L6OB4E9hk7B142
m6iGI6l4/Ph7PhKKu7HVTjCVUWaB8cdq/ATd8MHADi9JilghGa0ozIGBgjkDbYcYsvNqT25qbQ01
zd8HNDDFIY1MKbZqHYkLrUQGHzinRIXUAdyEg31/5H+L/wgWLAPZ4N31SBbM2fkQC1996MvZNA+U
DgM3MyKNPqohEhSeu011driz8Xxe6ZCXf0jxUTF6xswf8NpXQd+8ZVjQ8j4RNQ3fbylO/jvyPEoB
7nI9jmHDhGwnf1RTqn6HxhiUGly/h9BJ6xnVlJUWyfo+Sryhk40MukUCEFADtRontLPobNa7F2ao
sB+Uwbqk9plPlScXkvZ1j/jhe405p5r7LRLFr61ERCt4SgJ5WlPu3xemY3CRREMq4Q/9V63AtZQt
Lk3qsLheo7qPE13sFO+g6Jf0c6JNsDjSkr5uJD4Kb/6/kkWq5KVjwjpl+syvXAsfCbG52JA2mQMl
nxydLpjV0UWhwSCkwjNMGIrec1WcIOxdc4uUAyguVqWXMVAqJEfiux3EejBknKCNS91JRpHyjSoZ
tndf4IkAddAF3mu0TPRHCCIF7p82kPyLX1+gAOKTI+PTVpq5d7JHRh5UTVezdzaXNsZZcOpME0t/
JS6YmQRaJkMhLNoLv5Iwmd0OZuWqncM/cPl+piDkyFbm5QCUpylEuHAmwZGvK0O9bZAuTU9xGtIZ
L0SzxX5a76Ci1cmz2Se6AEgiO7/CNiisS3+umSP9qnIT+AblP8h7nhvPhqotAkPHZKNKKDP3FIhj
hr9J/SVpBdvNMpsRHnYuQGJJ8MohtPclCiTKXXmLYl2VbC7x5Dl1vt7sP5XHy9lrlWJBzpz4parg
aDyOr8Dk1beyY7j2Uf0fKld3gf+uKPdJ1jJR0R2CaVvDwOcNrP8SjWIDpmaStK4HyebgJXuruTFh
xdu7hWPsaAiDI70I6zSGivaAeZR0E0RHg4PswtdXmayMxb3rlrKMUySL1Gb57aX3GMYqRlCBj357
TWejqSVDH4WpaMUVOZUd0hWZ0/W8AMV61kHj7CtwkyvBJSAaGoYxwoFZ7b7+RRC25romRFubNtNJ
U++ZN25XfPlxLwGOg2884w3AtwlAiAhJ9Vu92g+gLmXD6FUUMoMQsZBsdY+5qqFLqaJJD7MFgflB
w7F2FWSbou4QFJW/A6iHIDfyQGtl01PPnUIQRiDF9F6qPwC5y2BiEjn2yH4j8QHL03CCw1COCVCv
zt+SC7DxO8hvBs03pI+SAAcOQU3xfPoVc+7iRohoWyZJdM4iOGLQy2QnyPESZ/wG148+2+SuXa8K
yTKHpuQZUfHhAjuj6BUHHrWzvcmWqd7/djhkV8Y+VtwHzZwH2HaV2f4W0NEXIdn1NIqzQCRCjLFq
tmNvOyKeZyzXvvp1OMtrndIaIZNldGmFl7TNRr6znpmGB/xDqACOIWEMJiCJPEMb3he3WvDaiam3
KmPTuR2np8JcLZS8IkLAfCbf3KyV45dKwSuysphnXe3spOAWHpGPzbV5X1wp8FIaAIMRJEPixfBf
L5a6x4ZQ4RPDojAYK9EH3BOIY7EsnCKqYs3GB8HRSaN6BE81zzZTF6OgKzL8YkIvT11FvEuYqLzM
vKzXgJsIPGkhWNRd83sF9xHMufYWItPKfVzTrAsx31nLYU2VkmAAUn8XWHwx1LFK43g3mhfG2ref
7PPS/jAIyIsLc+sgqe4u5wWV8yEzImqHlsZPfeyVksCTnktXYVbnetffT+gTEt+ILy9TJLJqtA53
a0YuvxnlYzfnvq0w1nvzCgDhfWz9zQoZZ1MljAAR+7pr8rovNwDm66tHrM0MyytmZhOztXeWSJoD
h0F7uaDjKbdCbiycQj9VML0fARIzeGkJtffamXFGG5zb7+Jqt3ItwWShph+xK+NAga7VTSegR8+9
KYoGXhMZuTupONdF4AVJ/vfivccNBJmYYRYvsdAGQAs4GI6XHMDrCtn+nayXn53bodwcYs+6KTUt
JujBSmOzm708quUQeXiHayM4/wqGeHEdN6nKPsWGNrIqApKo+NI7St/M4fBXUpIkm+4loYZo3Wow
8UTXsPLbp/n4CJUwvK+UZTo5X7nGsEZNuU6hDePnqb2DPvQGWECISDD2sxVv8q6BrcLqF+O/HbUR
vi9RJIDGaCrCXXx/cUf+/GDCEzunZWM53h1/q9PLDx4nH7PKme6eZepL2v1fjQ9VPYE78fLeoBNX
fbMgRC4IFK/YHVQDNKXKb0AnqVZ84yX6HKPNQAJ01Gn5+7JKqnuCaO3lpSxAoiwevSIr7nQ7jh6A
PeLALrG/ovypMOzg3CsdWclpZRwcFifEbGRf38uOrveOfvL5D2hU8uJgGizguFjvqviZUWGDCZcp
v2W2J5tnveiHtWmnTjvGWdDTmM083qYmUNXe20LE7pD9lMMsAON4AfBP1FFc7meROcMZEF0wqHn6
ZbIEnfCRjjA5r6furBeuFUo/B3czHocefuakVTbpqZSy+Hr8GqE217QwdBm3Py3Rv0/sAIISpOuY
hSGabGoTXMSD0WhtPTnWbzupKZeOzapAywpXN2FU9c4pdNoSMD3xIJVFwLO4KtVQ4MWLWHK48sPe
Dl7pSHPE16SbF+yWwJ27OBeYVdUG4x60qp68otCnDAsNMitkqXKbqc+SJqlIIcOI9j6NVqe2bPW0
Lv3QNCqZsR3XMggEQOTw25Gc7ItLBfrEvgTglHvO2kV2DQTnIHKnznNnq+vgXDJdlemS6E73hXV/
hKOiisfpcAOtOzH49dlXdZtTC4yQ2y4Si6sjs/1eqtd+IkTYwNA0dzYbkkSSjVcxxKJ0oqEMsHYn
WYo48FAAHCXYX/sqlQEGFm1fSuUrbIZB/Yn+PS3yJqFUwyiO+5jue69E7a+2nxkN1whRSbm6jJz+
GD9I1c6mhiH4qXuuhIg9tN4BqGT46z+dEmUFk4rcblKQ3UgtFbK0Q5jRJpBQC5nkmKtjqyKC8P+h
P92h+W0fMYGTtAA8EKylBhZFaPKej+sTRRGuGf6llvdoZpD+LdXvgBvEk4E2k3AZTzeXnBc/WMWV
1lsOP+MUxVv99UAxpCp7ADxfP9oPxXGadxH90vf3XH0rjC8OpCXnVrp/QvSOsY7HCtSiCaWzJurz
xNhBf3RkIK+ibsKslbF7SoiI9ONghYhjyKUbYcYjESRrpDXomA2z72s6gLsIrjNsKj4wvZ46m8H1
UZYV6tMVOU298LGeBoTcjtucvjypmxb5IbioM8Ea8PPzsa6sEoTusXYosU3Eu6KRqZmTf+7EC+/T
Glr2SdtEZm13YfyjGZQSC8y2zA/qjOhAxQGJoQpPPx52zDKDvIEaWAt8t/CAlNSziqoEVScK0nr1
RNvE1FVdA93OKrpsAWU3Jjn1+KtGtTKdQEnJbLxIMtIvCeZVtwqlzCzOV/ai+YW3g84zwrejrA4k
v8dotjzIx293G6mo6Aea0tFBnn2dAeWFgbDFO3vGgIVl2fjnSUBz520qMxiHrVnKax3wgFGlak99
p8cZGIou0+qzWk5saVPzDhEWC/QNuWf1NI35nVjsGjJ51JCGUSOubYdNyZrEbhJPuc3YI+HwVLeK
WzsqhJUzjHBexsVqnzB+/F39LoCDXyXWbZwhMnDtFo26j8u4Tm4a61OQP+1QZzMqFkRa9y9g5217
gWUhZL4GEmEaqAb5m14tUDWQo4sgbiop7XyMz5H0nxLSHUCRxadrKjuNs655MOK9FQio1naVJCwx
4KzA4QdchoY5DK5nEoHUZtYtYWfOYlzNfREtS+SCHjrqSG0QJWWSBkwYrR5iskXQ6XlpAs9+B3Zr
Xjo9cQ/MSf1Q/qNAO5EkbyfVV9f+KrR4gHeTBGfbElJ+jK6V9jiQ/e6ULXB39KOGjG0hTppe0aSc
ccvST//iF70Ds3mmYh/EkDw+YytDeC2M0XLvS71jwQR/ALUYWdDj+1aCxkn0gbahGnYsL/73e4Ni
rvi4+dhqyQamqOE0eIqmXDnzI0VMkPDuiskH0tY7IsKa0mTnbmwuIb6SRFh1FcrYmVk5Ha1cPE8W
mxfT8soIltTfXbZrzNB8htK0wHu6/yUy043lXmJgkrT6eD9AmYJkFWVHqaeN/4MfRU5fItWUYe9Y
WyCp2Hf18rkBHoP+wqXhhOuUH1EBLK4te+vYz3P2Q5y8WXnFO7NbUqChiXp1djAlRTCkl5WW8i6s
HOLxwedatBlvKWJgDSzW1RlCKuYrCCRNkwW6f8Hs6Qj74uEnmoo4PU0Ir0Zb9MwvzUekQlmptEqr
deaVm7rP1CexJDgzB+1bGk0wg4GoCk7A6FOHfGQsPYBMfgkkYS2ThmChj5HxRrobZDOxbwBBRL1s
FlmXqEL7JTe6PHk+LNrfnQ2e33HtUB+Yzi6w+49evuswd27cl8UGso34G+Q/26JoFLZc+cYFLyxC
030R5QSj44HOzZAwaOOBJZJimawkIHzusjXmojDyNzbCmPBCMSRsqCKckQWZnobmAlOGTGZZWWjN
y9hHpiJwgyWQ4p/Ip0UUPUS24Z7niYpm+yJ68raAwxOLbmkD1Gf7wpqTpLql62zWGGck4Qc4vkjE
botyTVsjcTAIUiV391ROb8Pa4hhUrrHIt7mn7T1YgiXNvwaUFnoX8/Yk3wAKztqfgGTpX5IgopJk
gY2b7D8IxCZBqmtCRWLP7Ti/7SVlLAJDQYT99TX1x56TObnv/GemkX2JeQygYR+dFslitrWBgE6f
ne1ekI3BAAGdgl9ziDWhFfnp5aTyxuZkoFOBikZXYbP6LXJ8AdLO1+PAQ1ovcLU8K9KONNkF3JnO
H8QNKo8pFIhTg8AIR2rf2lGjTfwmEnVtzharrCfB0SEN1NWnRAtzMtBjszEYgesAU9iS/5VstiQO
tyNJ0rwEljgJmkdrg/Efy9lo7HFdZRVnYhzVkzsewKRVyHvdFdr+2DOwyoo+sV3GMa/vxEOx5zEK
PXU1KaDbhuEls7Ne/hEYV/T5lWCmmyoMH6aV9vTH+catopNaPYhYlvZE6IkohSEC3yPtJx71YUnp
qNiLCqalYQis/kguNpME+dwlwJb56CMdl0vZpS6by76GGI2HrWJyiRWZZ/0R9gdHwwm2DPhRyIjJ
AX4zD7F9zn/fBkXuii2jQ1PgvR9kJ8UaBYOZ7QzoldvLMrr6N/pwX5vuA3Hl26kVTB8LhjS2hA/u
uS1GhTZGy9BBDR9pJ4me8Tx6dYFvZ1m6DHBmfvTu52nazOz2kAPkN9LJyiOKX7A49ZubbWBf3MP8
U+9gFQm59MqcKxFht2c25M+c7yRqWvEuupcHQrMe8/cIS+vVpz+m8pV7xiX2+sXBwvvQYb1pivKr
ykCabqbXCPeGHil5p8Pfsodbu6RljkX/S0Z5xlgZmI/bJlTQb4vSE57I42bxPHdQAmKk8nHrSold
KVlJtNOSoXiO9nL9mvoumX8/pzcwV+muAfozXW8inDtfxV2bwXIfnuzHD1rkyiltjPG2laC6Qahq
ul7MgmbWq3z3Wfdt78p1HqEA/2gTeB+sk9KUTBZRcFw/JNllZsA256r7HDhkezpmRsIoRk5LpyS4
8Pw/3tH0Xe+/4E+hVkTthQRpR8aYjvkxk33fvKiis3QdjWECyJxVymr7GnsnYU8WOIO4TJ/Xjm80
UuXLUNbO5lsGhMEIO7wJo1A7mVjuTLuwnKmNX7UeYBIChrBz2bwI21Ir5L/Yjw83hI0DbLSW6kuO
M+c8ddZcI2z2IsP38NcpoHlcO3MAQQnZTun2zQ7pBun7uhSUy3EKBjuBl4ejUU5x5kzq8ZMwKHyE
xnlmOfCa+Wpmrzb1oKhdLh58bknarrUy7ohDZX/zsZtX+Qx/3vRCN42B93SaQEBvLo3F61XvLQbY
mgbjnjpvpJbWfazv9jiSEDMueXXjf3yJXDuKtMTX0TM1zHJwpVGnvynnQq8BTks//45KoUTzXOTA
RPWGIugEhL6CPwvvZGXlL+je7R2yrjyKVxOZdrJKeCr5yZI+wZZhbeDHw5MsZB3+txec9tfulQ/e
x34dR6DuTxDiwO5NR1g63jsmHxb6PbqmrZU6ROLcRIhdyjU3zrLch5ul8EnGk1RWK3T6yofQ7sIn
BtvTUbjsI7CLd4uuejjZCPL7YjG0VA7d5FgYtJ+qVzXqz+GlbtNev0T0iWd7OfjLUl3tZa7I8eoW
y0HmDVUT6Fl0MeK6QFWU0SwnyG9YuD5gdBxTDJ4Kx4Pm+etBdYaxP8wK+JFtAFoMYPqDSlwDcqiB
+ao++ve7y8YW0P4HRWuu7IKtoFD30lHgHja/uYMa7fICQS8uzuS/pVzQhHiUY1PO5ADkcMLZ34wQ
NxOXPAkq2mjqbonmBv3d9rVO44bojz5vuQq0LquvpYfhvB6mgn121t3XqqK6OSLDQE8XH/1Sqad1
RQJjFEjZcqROh7u4OzKZsJQ1aVFOEVZKI7TdghFG2hGf9PGAQfiHNfHSVog+7GQlsKA7eBY7HGau
lTV7YE2Yy9obrJmVc1hX95tnKiehouwSHxRxwfu68+1t4jZRxNOctSYmlMFqpVG1EA6qX36O7swV
YhEdXw/U7yOYjOOhdzZOk/zKZk6zCOLRIjQy4w/RRiXZ8qluhwmrFiqAosvT61130bg4s1iz5xOu
L3xG6SIZTRoNhT4p+Fl/zQ2NuMxKVj+sFzfpDxd8wWqEqqa80rGS42MJkbZgO4FCdO6UAe7lw+Gr
zBPGWFwG/D6PosA3Js067r3xE05l7i8u2aUNzKLnr5VV6uhwLH6dfLxSeMdts9XTiTFEoQy9oItA
D6jjNXHSWE8inpu0xlNzquRFn0pgDUKOTSjFjam+jdiAFqZkdsWk3IfzRr9dNobw3FccKfSPHrtN
7AyrmxjwrFF0d68t2IN8CYpp+lMZj0X6ZtTRayBZ6prrpIN6MkTM0V0d6zdYgii30FVqz6y1Y5wD
f4ANT0op7vawKBgGsruf/2U+2W6hvBMnUH21KO6X6KGxaIOMfDwf9xjjl1jRubK4cCUhx78mbQm2
Druro+kLqXiG72q+oRbxGeOkk5+jkC4JIWwBdGDup/+Xfwu0yF+f1sZWtZb/Hu6mdyaPK5y75RQ+
oGhX3zHtVChci0A1QuI0COVjOQeenOxcAhwV5Tj6VTcX1C+1WLVCJf05rp2TmTsBLGBf3syl63ON
vI5EKW/z+WJEpHHMdrI68zoBNSAJkIlxUkRDGgSXvoKodEgC2obzUP0bpC5yu259caVWMy+6tNzO
Ui4fFdDflCYVW3pC+RcVLjYpXZoGF95wieNF4x5H5VtlbWn0oh78bED4WzLposePHYEfnqGWTPXE
+9y3wF682fnxldop4B/vhdE7o5CqckUd15SQR8sMBTGBrxbIjH2vhIEH/YT7n8Z+1DGxz2pqppha
rHBcdMR7DnYWxu9H2jgMqYa1I6V7ejjj0Pxp5njOMYXqS5p+bmNO49wrOFqS0L2p41/4pXvy3n6h
lRV1zbx5lvxEJpRk3aWXXKC9rV0H/XJzFy0SfP7te0YQwNQqaYKHIkqC1pSaCjnFYJUZjG9JeQhJ
lapYRpIcoTOc61l/nlLETmylYfKqVAJegfuImdmow1/NUwBMJm42/E2v1ZobwWUtW31RtH+m6x+V
X+YbnHWQFqZOJs42WS0MS5AxUZDCfpuaf9V3Q/SCT7znbkG1fmQBluwUBo7S9IiakdFXai+UXivp
ms4jWhG0Mp3cOsTm/LT/lwiJgn4ZBxuZSkY9ngSxfyrq88gcj33gqzOAn4uwBDevHSuNoSdwEvnJ
W0yGgstAPrpAvl92IpzumCJbssR2+g2zcJd7O/l6HWto+x6S2im6FCb+kq+V5sxacT0ZxI7gwwHe
Hu8k4+50sQHtS2tAOWVxrYhvmArV8WhFqwTaTvEqUwSFEODNOFAp7vlFw4ejUcVjDVw8uhuZes79
JhZvMxH8G77Z6eTMwd5fKs/Cq2bOl3bN2+Mzs9WRFGNxSnhzBS5sV5/xITxcCboYxgGMeBX+s/Ae
fadrFhO6iwWH71EgiqwvikKK97NTsong5HGhW+cyRyu8bLuBGAt5mKRfo9HrIVNb4EvyV5m+Kmz1
DiT3F5wVK29pF9+wMOq4+MeioKu+iuGJvdC/hQMYHtWmXtsgGx5PG/XDymjrNS7PfMVEvpgBRxGd
qGDZXsFM0XGE1N84VbKM9CQfKdYQRCRhvorG0Saw3Uop8YjG6M7cTQCDo/RP0Co+7RPn8IOhEssE
7PgJ+ncZsTehyhPv2S0hEGwMSBWyuEEhcw2cgRAVX52ThTVL1WVriXQ1q851eJRx/a/VK8niNQ5A
npP7MQvyUkLXJ2su3FfKYTnPeLdrjtF6YzxDrTXdxrW4KS89Cv58JgTRF29eK/PGPJ3Rd5H093nd
6NgJuw1IgysYclwiIgc7o45KKNtK+ooteb1jrOBhhRzMoYI6kyfYHo5YnM/x8yextiHOVeTtLOii
nqP3UBvuXg7RCsk/hLCNTATlJCyFIyBqlG0tjxjyPRxWmUlH3136S372h5JADGpUx9g4pmvjUmfe
FLuiTrXlhg0YaSg821zoxq/bktreY0Ff5m04ODZTcQAHRhpKuCn40pIjAtdGVYyLepM75JUW2Hgq
dboeJf26K3y54QCIbrzGyx2O6cmylQlR4YvlxHZZpFri5OQKtNr+Atpa/PiFaQTEVVcwEQ/L4Kce
WNUQ027IJgnWRQ+mn5JEDtf4BTyp5T/WarlDEkOlthg3GxryBrY0BNniWHggUTx7Y9OhUaahjSoj
lXbbA3Pcuk0HK80Z8VYlnezvfRh9ddHiFgdawwUQxcRYoXL1VOsC9WL/DDZ7VErxXFgv9xI/b/sT
ftWjf0FbCk2lO+QQUpIwVuyW2sK3XvO5lg2HPMuEcA7BDNvkHA69rwzvRLwphvwTunQHWSTODdEr
UA1mq2KdmWhrG9j0gc1iKkjdzSUyLw3gdcEe6MynWQWujSpCQcLbI/RrC0ocYrf3o4GxAaybTQ9G
up5J6Uj5bcCNVJhlr/dhKmp0NmzPu+PFvmwTK2JSflxErKOKjda7zrkK/DIDdSWBXIPNPrOQdEiq
5kQm+/Y6vFoOHInLTZPXZodKzSlWaYD60eRLkm26/EkAOzVjdXf//UTpk1iOUryEDml9T0rf5RdE
qYj08WAPncIBN1khp+FE2HbgNtCw20jVh0R5WzcltIlF2jSnPRIhZBnhHee0w7AZJF9pw57iuGwC
IWIOWv9C3CmZqUVvLpnw9nYGnzhRBKNFvwBjHQpEpmtjkH9PvYGL5BuSi1ATkk6+lPcP77jXzWvX
PUjFGQE8KAKDT17aRCJj0txOIyZbM2CRtTvK/T+vZqPTGQirMrWWFC2VXrtREmmi1xuWXO2tCaGC
SUErUQn+6xzklpNuJiWZfONItfwc3+EpYOG6sGXhjDdXjuFgauQtpsv9I8sDd/aNNIhfZwxyyegr
ai70r85Xl/w+P1aIUksHveU06On7pDBmOrh0YJmjpfL6AXPJJ3veRah+AP5l2Ggd5KByH+oLDn6m
L8CGRRN4ch+kmUSONIm4upPPFeYUCJlTPnuVkgw1Pm2Sy15q9b1F8fGFlt5Z9EAhrKxGX/D4tj6N
6W4NdRxEnFv/Wdb/Jcr5MPv7YXKqAC1QHnNTgRMRNg9odPGXKoM/gnwzdcWy0AjhEVZv6gzOhY39
WE3Cm8qSNOfmLSvOugLFc6ushxQddIi7cV11EFzNWfo0g1gWQy31Rsi4IS5ZgZKa9VQ8JxuDGjzm
nE/u1GLjNL8k3hyIdToymGJhWHzguw67j8/Js8qZHUsKUsZ1LSVluMG0NrwzIbdZx7eoySM4BQWC
PoFSC1MqpJNfMyl9jrzoT3X7yPn9UIX2lZxPxW9/RyP5fpewLgNHqAzshvoFOEzvYX5EVKEIGa6y
gz4OEh6JYPV2erJW14vspummNlWg07iIAza7li1QBPMVXIyaUBoXrrtx2R+xOGJEhZBsgYR567bg
UDsabvqhRt1RASBSIApZjldoHT0QLI65nSRvz2/gGDC8xoLzIQpXWEI0EgQMh7gXbSELUjjNWGNY
3vfYYfD63xdQrAsIW0pMNK/yZoNx7QLh6esdAMlAeHmc29osqWlAeVk9M8jER0PQQzh/En8Sim+S
Dn3k/IfEvmIKWReP3tSwthSudgsmZa/gJuxdcv7qJBXI9JKZ300xBXSWsVlPqw7j4GQ6OSk1z8aP
GOtmhSuXyS5OyBV0apt1zFffm2WxtsBfWZvM2KAifjj8czAegLUTQy2QtYAlKzhAO4Xd5/12EfH6
zdxn87gmnDzNxsN9Yl1zKUwWPuaTuzGSZ5vmkmoH0ccorVo3uFzEFStjiUb0Hgczbx8kPox7/Cox
u0GYuO/VS7Pgx0pv6BECkQcFJdmLU5A3fyu1I/NxqomPcXDcIiABRkvactUW9qB5Kps85uAjqFwe
tJxHzqvGHUGzuChSZnXVF2LDs1texmfX7oLzVyScjA5jSKQakTw7GxcUJgX5SHFjfAwId3ImXYHG
BJpOKiLzW8hvahN1OA3y5xAYQRRRHoAdcX0xWttGWRJfHFyYtHdPIIySTuCnY2pKjJpHeS0Nt14t
oy0EeYzKts3NWOvgKPEiG9AnieLqa6pJNVDgHS8onSOGjsmS92hkVxZyUgly+UvlCm12Yhv6U6HY
B2hjOK792DLIzSzd0JAwRrcMPzVuJhjVU9Ks5OkRBVmPZlDnYK5gtjACFK6guZFMycY/zMdj/6gb
BXGT+Pa4ih2xOe0y7xm4+3FiqMj6c53av3Mj/3SuIAPFCg18i0PuH74kvWY1y4DKpN0GxyreSA4g
MXqcoZo2wu4oYeURbeoWzKRFY3e/vNahAC7Ujx2lahOFMPMLcvdQQwXvZ/xDKH+pF9FwSF2+NxqN
rrkdUORRQWF2H0JoLX1SBkzQqmwDTNM+d8svz+1uQkK5pdPi5lnKJ2IMUCqhjBVQUpYGKPLyceN6
cr8Wv5UiPxyl5yn8JXvWnlQmkbCg0AeeuoUe7kuyXeLM/93IPxiUOK0FjghPN7YjP4arFv+yI2Iz
LDRRrkYGD/lSli+vKGTG5BLTKQmueDRvaNxJL9MF9QSpL8/lDM2481M2NLdd1jbIzUmaBqJBn2Xx
K6uPgkeaykbPdQ+tiVkssCbOtPnV5HgMebu0XYL9dgaQn8tlCruyPkX2GYkqPc8fBxpZoxHaXEw6
abgW3DIBmdGMES1QMSXPW6ynwueozLKKnrlZugHY399cgQxQkj+v/AGUjsMOPMJydtDibe3eaJSW
1ZpYlh9UYjLTdsdqFzuPP7qZrtGWH1IaVxYSSQBHV6+oAqmyHPXe+Oj/3Mx8JmLc3kfu+0iBO03e
sGqzuPNKBC5iKDxir0sJZK7kE/XLZEBLJVsSYyxm4QeGhrZ9VgCNBuX3kydMlpm+IYyU3HEjDTQ9
xpAsK9hjydZKOSubuiSTZsSaeXfr30fffSwkhYt43mCdSXhBfLsXv9H31icuLgohh8+Z/jm0IIZ9
xAPU90TvwP0RiLxXm/Ajf28CjlTnGklDSj8ULtQ5VLNsLhLIjI+SD1R4iT4Ep2d69PwgmAAnvuL4
7wTbVgUrLY9RIiq3bZYoLx7od9gQ2B/2Dxh0KS+kQUWl7BLRDM3CM6Ox4UEOTiKWRP6szrN5RNgh
0wH3rMtjYlBrhhDL76a1ojE4gLtyY1bI4wRMnH44rp3GH792Qo/tUTT+lHLjXpxtS8RsEqXeOIjN
+Es+fjZThxq4PI1N+33vwLYKqHSFq58OjI4+Blfu7pOr29nR4eS/59Ny1s/lSCrI9v3Kp22rgDjG
vDcBUrDHKGNIttGSojdJk1ezUIG8g488oov6od/OOutCXSqDtpxXucESwyq08Bsm3Xq+iFaW4XDR
ALQIFv8KU2b7Pvb85HQuDhbn/HD3XAh4KTvaZ6VWvnxj/QG+HPj79v81XDtjrhrQOkRumlvayma/
4VnOkwIYxqJMQXnSvzsYaL8Bcu7m8K3MAkPihQ7FcaWQA62NZKjaXpvgk869UL3IgU6GT9Be5XSx
g5xaYUA3GK2WXqhVVTn5kSS+954eY2Bb85EqFWF4PYp9Ly+3UX0Bf8pl1bAMp1SWQc+sjrYt+C/c
7sNN4M5/HnhrJFcDFS09VZURZywU0lmo50PeAxNiwzSZHePyPRO5OmnT0A16AQdZIcwgjtD+/XLz
8em1xSD0hw6XLw3J/I+CfHHXqy9UWZw303Aba0l4xlozJZJQuu9ar+ALrphBoe9V2v5m28L36AkZ
1XJ5rAc3gqKCJUYGQmo0umroDeWYuoXz3T2sPXowjJSj0op5DjiZ0xzcW4lDIniEOEiBIO2Pfpi0
+g2mYelZjQlg6m/AS7ghXFvm+Ok6OjAHlGnFuJ5LczelSLCtWh7F1/yUKlbNCpfIC/lL/k2/P1a1
qVlDHM++RupoWlJCK/lKEPFWaBmnK2ZEGUopDyubbRZpfIYKjurs89ytzR2djXYwqyOAq3xzmVi0
3oBnrS17Z6HARESL7kW3ee1bIQMfpYIc610X/PhCpEJgytYxnQbi/YuJnUIvRpZIGU22BvhhMuIS
qeENCWfqKJfYQpah8YvRcx3q+aaNNPBPcp1gowIM9W+xz4S1r76Cn552O9q1lW9VmDpv6E05X9+W
lF0lgbwX0cRd1hpeIWSTVpzD+pupqiOXqJ0aoJ2OlFespU1Rd7vwFSAmXyEn3izy8H4oNl/ba9ft
ztPY8AJdZVFpUfHPCw82lMyCXanJ2mp+HMBDl4JiCutksrR1f6JOQXxk3OimGDHt5Tu3a7P/GcBG
rQ+n4HNy4CkGx8M3A+JCip5JSZ8kzYWDVaBNtNaQK6i44VbS8nT1AIBgBLM3geEV3jmlw2ZQF/x4
WJi22RB0OQpori0w5PhOkpDJiKfd62pkXCBFi8AdL26G1hACyVIZLnew2kjRYctwZFWNS+ZiQtg/
jWl2Q4HMFJULjtAgJiHdAwPDQ+wIw/x4Rm5Qqe71oAJPErQkFBn/jk8VovF/3kemckMm7p6KeMVz
tJWLYyBLJ4vfRw7ucWfQUcdNexkFSEg2CbiJk/GvyoXSG6tk7Y3H7mEM3r59cNnwYX85rxJO3A7m
d0xAVxwwoTBt+cRU6E4l4KepIam0m/RI+e6Yiebo1pMZogj2YiCQXjcxR0KVGeUBmP1x9GnuqNn1
PXN+qJBJCysNlDBQ08gqxvyVgAElZEYrfrq3DGmmFozx4XozdHgoWmsWfu/+Bkb9izuSjiWoutda
uoQRZJsIHAToWLTMq2oBf1cOlIYrOiO7DYc8LDUbOiE5BXHtmNGBZDqGba8QN7MBBWBwbhM4e4R3
v2spojwzus3l/aqh0PX+/Tz6hyyvNG5vUfIG8CJGzlBrFoxqPrKBW0w03aQI8EsGqS50p5WU/UQ3
6jQFBHwGYXo7PRL23MmTrBSNFOqvDJAtCBLV69Ms/yZwa+d7UEPShPh9nHLxUgDfD+MAZ2DtvUTK
PJIQOIMqyLwrPUv3X68gXSQFHfZVHsfGSIFyGBsMMvwZKGu+ULndzd4jqWT3HJeYo2rdZX3mG5Dn
k+gvci2o5ei9wVUFIZi8jRjMzAVkUinrWjZACUNRqX4tUueqvT0ioBP9SB5I0hox+xxaLFKAUhZ0
4fQxzsYTFkscUT56I31qhfF2NrfjVtyrYZMiai2SVxAMioVO34eBca2gw3+IziSCjGRfu/e/hB7K
6U89VEADEYYgQVbWh4FEaqZVPQ46f09XYvwpr3hwOBhc3ZeL08AG17b7mT6a2WCiaoB6+HSfeSpz
pUfT5QkWGu8Hb8gV+yId6qXWdPBnPR+cgaYvMbgIVtdZIWoj0mar/y6iGLHScycOXSzR0RB5u+dy
UFQpY5VuqPtEclyeV6+1EU0gTr7onghUg0jvzM/k41obf9+uZPPAc+TcM1NRLiZSf/HNuWjD2je2
VyBaYJLw791EEF0ALGmofdj8i6ZcsEr6hTCj8YVEdZgWOY9fuKf3/8sq+b4wpYTOExMCTwiq336B
hlPZrPVUcThLnSU6XHtRSzXhMfwYRRDt5QS36TkvIAdcduSmi5xT6QU9r9uTdhy6bQFl57/iZHcx
v8XmmPOdJvygLMSfrsrDGsSbv/6aVU/KqPjfZvNaPEjTalnUi3kcl9KGQ8ybhjyEEGtrkSHMELAY
Fi0rcyz7YSJwKSHKWh0b0b22Ofm2e6GivkaC/qo2or5rPO9MWKbkjvuHxid8XQJ09MxDTHVQIpO/
G/at3aJBLUGLKlvU7Ty5ZHP8Xy/sZbcVBsOqaybJNU98Bh8Ll+q+pX2LRhf36PshMi5wtlpPbIqE
qEQ2hyhiwljPZG8l4h7oubfinJQugrQ4QJqxIhGFfh3jG8v44K87sQoIRL07jMjOGvn+sFlSLeWI
IDpWeqwtaA8Q9l9njI4/AEbuFkpjAAsk57tm4SXoh3t840zxnZCSerjIMppq1oDNTsBvgxtQ+Ih+
5mmGN9/sJGYou2ooN7jjUgqaUIWueGC+hgGjN0nUK30tify8RvRtRBeD8VFHCod7hj3ZgqLj6iO9
Gt+/Okpq/YwtpJ/uR3AikcZkazxTV4bLY/KnmIMgO05jAFbhmQb0YZgTJvOUBKTmF/qsLDbdtP9Y
wQf8yq6xmOaTAyMAjr7SR06ervnmn/bbjf2A3vBAJ6fyBz3J2+GxkNFux84exXlwXR6oO/NhXy+o
ltgVGTaSKBpEcUSRFNLON0bDdIZraFmi5ICuD6nek3R3uj0rhghPC/1VJ9CqhpuQ1D0VbENQ0MQl
9q86TykmCNU7zTQUZXc68AAK9NOv6LKrQ9Q28132ZreGJfgpcEZWjsIrjkUlgetTpBp2iwxFNFDM
lLjFGfnj1MWe/f6qinrtsLaU2Iis/X9PqJ2WOOp3K5xa8m85xu/u9LK/sd7PE8dfn7yODZEhJxK4
jUgkM6mZmxT7htdhda+x0rabwSr3Be0MdNvaglIccVRsW1fGWfY7GgN7Xz2rI/zZF2MJioQhgL+T
VD5MJYmF4urnNKXDz62T1mg3MQ+gVXe6d9SVqCXRCcnTnH8THpbUlj9dwge8f5hlvfySDCqWl2wP
9V2+ihITpHapfj5cTSIhqh254sCOrLi+YoW4fHB2rqL55mpBBIE0eQ9k/95iybCcGKngyfhoKSUM
LuiQPZ/M/VcIvyHehgVQCjF8blPC/Olk4v9kfolcxD/SK4oGmVvxw8FGr02WmlNbeSvSm7PUL7VM
d/muxpk9YaKSBZf4D0sxgnhMd4A1YkqGOGNcCcaKes8YV2b4wwaeRXGqNfYRQtV0mFmOfiXC+aiO
kbSkepI2GQY0hJPwTtBb4AobMhybcT+hSGNQHg+W2MYsfOq2qwirOUb8Y+bqoebi6uVHciIrvWCo
CGUGODZTRbTFLl7uld939hmmGlvOL5QycqABUNK+dAsn9MrDwOvZChfdZGY/sEQt3g1F7YOiAY0Y
jZdPkmrSjuR0l1x5bYYE5zhn5lX3E56lrfbtn5Gq/emN8oFGVmphITlPW37dve9dq+l00SyMW70F
+cWhdJ2VswNWYMwb+MOEcqk5N6Eoip/ldQmfAt2qJk8SKh0SplH1Xkm2oU7UdenGP2d77ThedfL4
kzPZLQDe/tz5SRfI463wDo6FiQSdm/7QuPxWerFNoQsJWhrEVf8V4fQu+j+mb5ySPgBAJSQv7vbY
jNhjqimjsOcevVUWk2CNAqNLsyX4aMgFt2+P4xPadIXu/tsKYLmCsQs7h/E1AG7dEK4BgvoXD5zw
Nr5lvpER7vXD/wwk8dC6zF6lCJPcGer7fwcLFcvlJZNZI/4PV1ire9WUfK5KnZ4Ikfo9AcoW9px5
QT61U7mK/+323SOYu+0PGi+kcyUuDZdBGJRslr0DqPu2l8ZJMvGLaCQH6hi3c4g9LZVnpB0IxFcQ
B2JdlxZxDNVC7hV7yFZxg+pGgHIS3lpuQ5Iw7BZbeSt3+iNH3eFy3SJXwST2F7ArYr86M5+SXk0v
J4KvdMnqLvZMTwDf2IjeWxARYUrrMUnF8hWhzrbOOjM6OVFPF2t8gj3zty6CTEV7muXfofJamT+p
mEtL6SymYTSeNBu6vrPXtWIwTVJ00GJIg9UmO2N6qkBKnFqOq4pOD3K8G+BxGWCCIMT/bSv79xum
PwKsmUwjpNKPlVLGPJ+4tljVbNfMagcvBSSbxvzcvdc7BkqrjQi09+QeqYvhGYBXFjF4FXyHUsDh
55M9xGkc51S64anFs8iqf3yF6XZKyehrcR0PYWhzXEy/qVv0dUj03tEx98n5tjjloU+MzL2Mc+qm
xtU2QcawGv/7x0JujFLlfhW/Viaco8yCThAlWf8VzKBTVIgfHzTNTsEHKKCx+/4uz9RFl1E2Y3Hp
iOtzZTMC7zX/whaaEOrqS1Nc+87IZJKwhZk8KzYX+zxu5wwqk9KbyoMYOwsK55EthGaFklgmSSxL
u5+4Fw81JYNFqU8FEfH9vKeMRSg9FJCqlGL15HxEdjugqmWE7vTvtoC3xYA0BYo8wVgA7/5h8v03
UVk3f7aXEEBBZcjpGWjz0CT/9nNxKl2y9BRrPDRzJUb1zx3nxFrVCJ0fRfDSKuLEP9GVD00PxQM3
2EZtn3AQMAK+czuesvEzvgOS4mM332hR3n7pA/NchbLQWysNM3bwWVMeXEz+ji76Lxgj37FP3WRT
xauew7bhTagzb9ciBAnGi5IYa6P4xyC4X96d1BLXhSPcbufLd/kaSd2JR7h4BDISpKwtmZUGRzWg
Lv/q9zfrEx2I7yAa+eT0D89dld03Gh3+kBk4ux4O0R9bNdISSn2YQMcus+Idjx2tcwWjbCgJ5cIH
LL2+1Su1yYV8Rv0YA/ZoupsGAkyxHVvEEg8LNagTrbVM1XbYohzRWZwUDHoApjhyJoP9tBHsk1yK
IikSIxBxaRZj93Q72WhhfNoO7OiT2tmthaSHtqIS0rWCXCjn+FrgaRbpvbLEawhkgwiiG98KpKlY
U/3mxdLjLp6oHj2jZnPqFiCWeeHtLC4eWl+ah+fze4vcKXi0RjzdlZEUmZqLB7dI4oEiE7PnuMcT
3T+LPq/rY4OoatK+ZDjg0uN0e4Xlf65Xzkmeogzy517qqaZXgETHufgKaTOlT5Yhlk1L0qOYcK3l
sc0SQS+kLwDmZBnuYdgM4g2fmL3MiOkMNzqDc47rbaQ6QAVIRDAgegEB/wcdItD4qokKbqoBTr2l
yxZbmf5nd3R6oVw8SvulLCPMesCAxtWKZHxPLMDmV3kT5DFlYf6dbF8kY6Cz+vLEr1gOTUzQeJZh
7vTGXb0JGzHfq9B1Ykoocj8HaRlMBc8VtfcRZ1SKLswBWBKYPxgFQ6lSED8Zzo056XAkbYuO3LEA
P2qxhgPhfvwLt2jMqN60Fg8TqgiSrxzUUIy6XbGG7Wirek64y+yVtcmlXWGjE7QlNrVTW/bCtuht
xhedoVG7viLBxIdHu0MPrFR/T2xym7LtIMfV/7CsIx+cK067GsRxkRpjqJBfiz3A4XeQz9S+tCI3
1HnE7GvTXro7PK7Hxn+8SBDYGA6LD0duuce0Rhx30aO+SdhU9ZSU+ORdi+3K8/TqzW9OTNd2fgTj
/uaqXyTLVQ1YUwa6vIDdCVXT+U0pv/tWMLYT+xU6SzIBFO8EPWDKa6fBfqsRmXgzTvGcdn3Q64Y6
+D9UjmRKG2CasOcgisKc2LESHiigQh290AwdTOPDsP580fhxrKB5P/ct1lYV9oEg5N7ZI3JTt4ES
8FThcYtMwTQDpesE43SLHWLQedZOvV9f089hHW7yx3cxprafb85Lq1F94Ow1w8fw5ih3vXaQ/SM8
TBnYJu5tyXMQFgXK+rBVGOuVMYy+onSZBnCwuxfc24uxGinIXbBT5umabN6lKUPjNfS7cHczgtRy
NW4zcQ5PcceMON1qMqBO1sPNzzSTQEDMgqzaABlUcJOI1Aoh3yeQuoQueL1KncmDuLCy+wfyEg9+
UW8T+jR0ZERJ7CmHqvKPhi4NNRNnnROQB/o5LIgLqnuZBdZ+ZH9JBIHuOfw/aDPwQ9mMPni7Uh5s
zjVI0xJhnoyV81dD4ayQ6zD14fw2t+M0zJdtWysgkdXTYtV90EKP1mNCREf4egg9oggrDr2nbnt6
+XW2x5eXw6MpvT3gEl0HGZSTcH9iRfVzBqw6xGTtmrcssckfrYy17kM3fYi/e9L1YqjkXb5kgKqD
B5gJiuB96cF5/MPb5U7DrfxmR1UOEVXdGfT+vjcVcFUcbNANBn4W5d31xOaUlJZ749wUV+rOSK5F
HYceag2Y9wOAmiv5DEl8ra8GH5Rvjs28A/ZftKW0JrDzK4wtysWpjqwxuN+jbhzKnDG8p7zYMFQw
EJw78PJw9w0uQyVkLt0C/k1vpWhKjpIMOchP5ly/w4gnEKU/EFpbL6avU8E2mHvQuEBDuKdtQQ52
rT++h/AKArK1eAH3RTrxA1nlUTNtF+Nr/OD2J4wjcchyna4LtGzhOP78oZ8V/x9x3vUu15kKwMwl
zHM5gb9q3UokJIHNrsT6yRQr3ssaq9Wl/cdf342+Ra27ucZqx0zgXuIX594nPEH7FxpvGICjPAzQ
xgEQzFXq6DZHHeh17P/RmI+c77AbWdhUP/Nu9HhMXUaAWqd8gg4dTe2MBIDX1XYQhilrHtxY+Nym
664XpyxYpRgKc27OTZaTo9mooQ7vl+a5xl3nrztQ24Lhnx0q7CYfygD2m6XurqNgYcZ0C9G3JfaT
LnaHLHOa2u0uWDW/mYof7pJZgOeTcXSPmo9IA+b4ytGGPstoCEAkPtq0Al6gTHa6s2WPUYmFe7cI
4K5rnhQ/XG8a6O8mGbXZJ1k4sVS6l0OtJGvJg8x4GKMR7DllYj5oMkekt3Txv8Tc5wsZOi1eOKyk
1JmJFh+SvSmHVw8XZHghFmR/l6ol6+Fc0+R2ppOqBApUJpfGLNvc5U1ASxnYUoSsTh4nMnAXgXKJ
8jCq/Sybkrt2SKptoXOFs+jDIKkd/V1ncpbGCA/+ozPg9/ipd+lF8Jo5tOz7NgAdEYJZrz91E9g4
1QoZadPLs11k8SvN20NMCY2uc1kSKRJv0d41i//hTvjr/Rn4hPbAdYXl2r6IjPZKwC0IKd4JMuZB
1wVs2poTY+IeRs+UP5Xszmm+Wc//dzKvgp85a0uBLFaxOsimrpjjTy2+Sw4i0ksZA3vUaT0yEdwL
I7BNYFTWUZwYazNPRCrDBHW57OiRvRXTMSbDZB3uX7gsUgpdE6QeubDZmT0MjZFDuxZI+kwOwwT5
R5tgQsS3YsChsKiHIRLSSmin5lb5vwdgpwmC6xBTKi8eP4Dhi90Ilg87MSN54JPrufV1hBcnthq5
PrTxtWpMEhp0n6UKC3JkDnkEE7JyS10tVfIEByANE1/uZvak7qupxhLLr6RGa13bX8J4yPxXqxeN
ayhbAMrmGVD05cBXDT5zPPrmOGGV3gL0VCghGouHJ2OpLbxugn91vQIHFG5sTqy7LEsC+88PsRfC
hfx3UBNBzhygx3EU7V6yYz57Meoyp8BQGTjv21A3dsO7IRcrqPz7AAopxPdDbANqyMgFr6kkjIEZ
h0CcKSmMrEKxMIGqmjjqrjfVpVhnvx8qy0fmzARwvqmsDrGdWwQQhOHeHPtU79P+n3N/MQxi90L0
hAgGBzG5S7MwaUqQ1sMN1+Z14zIbCbJZt8oovW25dgQtmkuxhAzb10C9yjKD33zUZJUGs72wtBfg
vy9CCI2nDkyO9kGUuuSBPlfdsv7vy9vQqpgxc8HfA+gZ0A9jjHB1MyBzK+8Ezm2kmuZpOT1O9FYf
xRXdA95J/al9KJfhKG7nI0jd6xiFkchT1C+X1F39w7Su3zUODgxsIVP0VoAmMI4AJsW0uhY8jSJI
h4VL07gSnwsuB/wb0RrFp2Vk07yUNgT1fSTQDiGAwAJtDVJ3Q/eUV3Pj9F3QlwoYKG44lT13pVTU
ek0c/A0I2VgNhO5/Kf0FIrYnq7PNe0jqj/V81DrZ9+8tVsLZmKU/2SxM2yE1FMmARhnjGoIAF4J6
VJwcfGHYHpqt8W8nm3GPn17i2Rt6yywe35iEEP/Sf5uCAt/1nAVTiqXOfIJ2rqP+bgZR9ZaMaBod
ICsSLp6ywFgxvBYgXpCbwDMh1cq+hdVE7GyOk+7ScG8wQVboJ0H1BpXZSh5Ki4jdrbTiC21+XMNA
hYeY+niaB7V7g8ap8qN2tHeE6XxdBlBcLNO39cjomzc0quLSpFmOe9N2iKeg3aaetEdG7oMCsbmD
xF7UInnx/PhVZgJR8E6J/4bR5sGLTrfwF5BASr2177nI1ihoareIFLTgVcaO8XFSnFxMxZ/uAa7I
gzPwM/hukz9bvZvsFZ3wCt8ErDnyVTnxsgE+w4x0wOCbjG38zmjH47ru9iUlhA9lgbh3e42TmZUu
fRuqc5th3kZbs3R9qTzlqAjKrRpHneixfxZlOtMJI3UvOiT5+0gTvgWCMzkUJbEvw9vSUnqCenAZ
On72n0pp5vvW6sgVmkVMtQT2wf+8/3dHNG33hr04/+9UamilmqULwk3jTnonp1h4N5AVgESXSGHP
A00HRoQd09LYWpqeTUWV7ELb2i4y5tvTl9nc9mb36pKxmKlOFZGSgP1aIvfUz96ADy7kwLdlpzX2
/Y68nVXrqivsFVXeaIFVmhIWxxkAEkRDsKWPvuCjywOiYBHZ/qEZj6XPx+GHDULMA5ZHrZg1EZMz
oZ47kQv9G0Ox2Td5BBatHUz1oz3JS6cBM2jG3piyLfAW6EqdPSnkUihxY4e6wWm6ZjkFzlilXriB
k/wMRvA7Nljy55mZWePIKgNw88ISPeWQpaDrqXuCX2xcLi+50RCn1nr1g0UEOk3cfMtr2qbEsxjW
ZN/ydWCI6/xVytPoLtdzFZnitHSrJarsHRMX6XWdE8NSH8z+7ssqjcWkseMcsJI2pyGjBu0Cj7vk
1R4nrpnkgVPr7w/0kGNmJF+G1shL1Bcg7jTlSb+NSBjVcrblYTliooUzcok/uoTB5CXAmvUuISfL
9ZwaKHBWvSe2o831Lkboi2NalhpfYUsiESTyVEkxOOMzFy5VraGFiZFLwOeufNonpirU22rfJBMg
33UGiNl4ZfMpXlgzsWLVZkp4MUMmmQC7ect9faps45yqLUi5tHfsdMpMzuKIMR4q+FJXyg4Y5nxE
OqNm2zMgAj5ycimrVpIGzoRzWUdqYZko3yCvlyuPUPrJn44OzuNHnsrioqV9kAgSn4NS73I4K9HM
4tehdfMTHnc/FKXO4djX9rIyEYjOc+4wPHAjVc3OwxwhwwvlUQK30Gu3dAEunWRSE7/lUZcl8NGG
ttwdMAV/vIh4iHZoUC22K2bE9N0qiUB3LZvODK0iUkKyV6vkWAJrHJoqk4R4aeFalB8QeHmZuyx4
9R1W0CAr9oGoppQmKys6KvVo1Vf/yWAF03/Rl6U0GwNqEWwlgenme6oxYKfdgnt2tjA7kwXvljJ7
dekJhYm1VLdL4r/IcUjOwWjr5N1lgOCPVJFhVjHDkvvxZN1ssGrGCIGfckrjmXQvxpcunMPTH7uV
lTHFaReYYycslhz8jEqHD4++lROj8AxZORxp6S+QFq/P/XmScJ6fVCNizfw32ylzVwt7cL8sS3u1
X076p99bkwXRfw1b1YAYIC8E1Le+KBFs+czCeNCTRKKj9bZAlgOSn28V4+qxKY5Wl05rc2gxeRV0
CsCJsEJ2e9wDCvH+umHYrZzqWJgbOGun2ehtdbatlw/GfgKM0IM62iIpDwPWWNwE4LNF8fbwTVcU
VQ63enGzm+mitPEf9ET1kZ380oErxZMk2SXhjxL2ww1Typhq14AVqyyJsLMhJiL8X+o8XPasp/A9
cpVIzU3VFd8NgAQ6ybiXHdxXhW9/QTgVeobVXVBfEoc4Aa1oasGzUYcffi07fJMpwjH075bDE6Vh
8NGa9pnKiq8JTM7y3FqWw3uvkVXcu2dZrUjFrufPYGyl6goZtc5cZFj2mCSvtS66gajjzTgCi4bv
UlfCldv9BrlDGFm9ohIkvhfjGWyAnwSVq/78ow1gP9NDjvjiHit9SwAFYxFulB5k6RgPKa/w+VCg
zPVuNclJwybKUbmFiBAYnX2W7Zj5hv+6mQ0ZUI72LikpkIpf+BbiP6NxNDN8/lJDnWVXQdj7HRBp
D2txT0buY2Qh/73SImFwDirYXjkb1A8Z/2HoQw7qKg0v+1Ihppr0rkuS6cnM3BjmpP7wQPooB9H4
2nYY9jnS3W4bx8Ga+MwuNtuRzrZhiC8Qn7G8bcOrwaekUkrI7IsHhSb6bK71GzyhT+SV+YVtvTsu
VznXPwjOPC+7tqTN5qEpNFqQbfzAm3i5chtSSzWF5Lxpg0PwFTyS34kRQ9YYjnSbCkX6VTm82ROE
kUY72+Qm1kwom20TySilNiFZNmP1v3JuEwdc/m3x3QlKTtzkhEXhDinSOnE9Np2E+7P+01G1NZJA
bPFbWSCn1ZjDs00GTpGUP0Am0padfORKrWZKfx1AxjM3I5RUe5LqXu7RmiFqjgsuldCPL8Grm9gk
y/3H4c84C+htflNHRIJcGatm96LBil5uBsKgbW7iHLzygZrenrI8NMDoedpNL1OcxYgedAbYgp8c
qehJGMJGMGDccyCzA6nyIp+jyCbxHFG4B3JtRHVNDtBO3RoCqYzu7p0LyFNFAw7fHs3br3l/mHBZ
efIMMYGJcubKOsHRY3MiXq0AQx/IXgA/qZc5EpkDJQU8LvKq1WSbM8hKUuPyJmfdx/9c/nDUAJOL
dtBfNNgoHjFBBDOq0ryfoY7F9suJGzL5gNc6VrL5jP2aDyWRK8bJrrXsUfuS/1vDxWrH1ixN8bMR
ImPEI4Vt0FmWZB6M4JycJhIzGmmITE1l2ocmXAXpDpI3frOJiipLQl81HCAHO5kWQRxj44cBxHtz
MWqm3CtcAdiEJJpF0Q5COon+3LKzzS5Bt4jkLRM0EKBAch6/JvueGVp9Vdtv0jpnGPmnJx3sOM0O
kNy29VZ1n5F467xPBm7nwl1kTYTkgpYIeImLgNrQhvffnfnWuHcgREKzLRaVkAhgvy0VVIIP3nJA
LsfPBDWUidZtn5KK8G2D/X9+Wc82c87KYaOgXbN68wr7p0zaxOKNS73oEVG0+ocoS9bLRD0+F0sY
NQMU33Ydh7KCTIQ4gJUO+YwJOhHwWHPRnj/EppZyl0SXYm7bjNK0FZuQcRyxfItrUNk7Kw96CaGW
aW4PnZEcmhjJeyN3vmIgfftPwA5upKgvK18iFoKjYkJvHiC/6nwnYfzE1ILgjLRsJjz6l/oW/eyc
M3/xfy1PXv4gEyEZ4Ofa66tWHQ2yVLP+vUL23+URjNJqIX4H5dOWW8c3B4KZw+vMhJHV+CnsqkZb
2pyBGYY02krG9kbyhW2H4PcesAGIFdNQrLLV4HwUx42GCZAUo6YLVTixeC4AFrYvWZJ2rHu63uod
tZSyEvSMOPNFid+Vy1S+CNJ/o7k68pZIHE3Up3TnX1AEj9ZXzCvoAA+OZebS/bBBTN/4L7G01qZh
2jsmEq3V2tMd4OeRz0Z9qrVYjCgbJ3oDFLfBP8iMbMUuNM7HyWHkmSJ+75qAGLYe6lY83zeM/dkY
hrlRptwily5sHvB6MeI4RaHZJ6pjU6lHuHsbSuJt9QoV4y2lmT7MrFWVduyYmemAbtPSUL6Eca0C
o4q0/XlHnAy0Bu8FhI0KhdGB39ONVL+1en7oDTRolKelOjz1J8b2i/demjHag2Z1uUmLk1WKjRAm
lzjMbVrueVcm6DoxLJOFhsqvIwttgNhjty9Iou32m/E+F691x92luHb87dlX/Jgxma9uclsAiiA1
MxSv/Sh/GyRoCe4ltP0KSWLV4S0Lola9VIjjGr1YP0Rvr++j/FsZBituJpSTBEi8HR0YB7mMsJcM
f6Xw0D0Q0RENfl/VA0e3DC+/wDsSyMY1w0TIrK1pg9Jy2ZxnrJQhwp7rty4dnnUOkzM8oCpv/JPu
Z3EbnuDTcyf2MiZ0KD+Kw1Sf9VzLSu+tvdSYQrLI5hwlCSEa3K+lbDaYfyhN7LWbukYg/hy8kGqf
zQcxT3fktvoPAiFzimsoLGL3e7Z9kbAxdx3mRRsFMhr5U+mUrO3qNsUwmMshqQ8lYZ7XSz9TXbik
rpFbUxioAi+Lv6LWsDadD+n1gBeRD+1y4DMdXlJ/537fe7+hVLKSvJig9xIAQQrFUevkHlBkt0sO
1eQgTFQobiuZmRZjHTG/WgF4qHWeBYd3IWk5wXXKzvy7KSjwbQ/pZeskcflV06PxD4vhrOkElewe
IRIhLvlDtr4/yy+5keADns5c9isaPFGSsY1AYkk1h7sJLE2MPI0N4TxZ657npz0dU3/BKPYNGiX9
f7PXwlAeGeace95shLRFLsm1u915OtjLTuYz3gYDhWPukTACdSHCKwfe8aGzLeoeuEVbvjI8ZZZl
rlmoKwq7w1umpeB7uoWyaGPjIUJhCEYFnNrUNO72HfV6a5IYp0n7BKHBPCkkjX6VzS73b67pA06Q
lB3X7mRwrVxljkTxxs2YzuFtlEgaXTN8bc5SOAsabwKnfXzIYArfVcKyEqmZGkQuy10Wa2iUC4iZ
Gk8yz338kmlnylQGPjqXi5n445PUPXGa3CL9s5TI9iwmnNh6pYNT1KyiT6M28JS4+XrU1G3mIP+h
ZZ4nRVGmVzkk5lVG4ucnAzC4laseBO7Fz0v7ZkKOi65+H86uov5EilFT86LU5Y6/U/P2QVco5z08
pcTp3sG3RIx/M+bbH+eHfnnWlfEzl8NwwTgR+iImhGn6dpBKgqHKix4jh0k65NlCiPZgIKoYX2c1
3iRK/2J4ODfEMLqKpRgFCpdFFjKqOWYebGY9G7tAU5cS4VX+aTtztA9KwYxdEn9wgqLaN1/3UPz8
Cs3fOyZHL1qlfSj1sg2GTW0edH6sy45MiMwTOGkBpCL5wstIW+VVqpUZO4ZjAqOMfnJSK4qL10tq
vgqJZWujEvdKdpMZqNI7okm6fNjPIXEzaRQr1nmzu6ecweThFCKii/aQ0OEUM/kAdWj5lYLgvtlo
+BGbPZVLTKNSqzehfwKfxKeXuzCi8Eb6rxzOPBg83YT6nQqSoZCTaaFvjbGya9SF0xGucuvQ+6WJ
w5ef132cOU3vtJUHve43wEupiOQJ3s7AjDdczHSSSN+QfAWo0+ACH4kbu9gjq1ovZlBK24D0LGMb
O6CtbZMhoOYRJQpuivR11t5BtH7R5xd99JqZeArmuKxppV6Dl3pfcW1AD5FpK9RYz4Z441BbTKFy
mJot4eG62ycGjX/vL97TXU+IlyNFDqrpR38yFHj//jB9KcrMZfkTdoK2BswsZSKJzNJVMvi86XBy
95gXTJxbazWMHi0okj9kzwnav2NoQbAT05yEtqC2dCwRw+onJ7xvW6kO9lX2Ymwc9LtatAjNxkA0
94jgkCjqHdHb7ciWh0qjhbSszen17uKMU6UjCu83ksa2xZ2mqQsL5mvn4hZbik9gwlwo97MFdXcl
homgd7T20aG/vYQtuw5wztpQIdinlBsTfCu2xYr2w5lvYCreQDIjYxKvPdLXW5Icm+3TPXtZM3FB
0BUZcWhDYJ7oZSB2PD2+HHSGOwWwUi5H1xpLbMDDjjNtycHf13cFi2YLkjfzQP4VEFOhIIqYsZLN
DTitbt9BGDQGSxerJ92e9rFTjnqKm7qivh0lctKmPJ3w8jkKiNKSEGoemlkW7LZ3YlJe8bqwneP/
xA3eogFmjA9B3Oces4WQEjIDcanYWvJUa1oSGyJ0xgNhUzCeuwjjrXzYq6QLWsmYw0erz/PXrASe
Ua1xeHhfTzC9m3xIxP0g6gKQay2opk5DiVj+BIvcWVpoIlHiPPIfQ6tpsO9PUCq08si04h2vEtHs
L6dGGNT8vUKujnS+W3lTaDbE9vNV/A8/rcqh8wwkmH82tmRkYukNx/jrIc/mlfl6xaIlYeRvwb/N
XifM+n3niwl4DGlf2UfPeYLfSqjsNTNRVR7HbMQtOKnD7IBoizktIQ8+28VpfxhqVBJ6+Dlbb1b9
ZFsOfcE638tJzHJw9lg3oJEHjDpKznTy21X6GWXkJRP1MXz0RbmC9ulaLM1CECM0Wa6/YL4dX7lC
Z/0L/OGdb9pQCXIWGDo7td1bQ9cBf310INBsrBDvA9V7yaTac1mFvxYmezZNEBQ5zbUc+m5nfbxV
M0sJOXuAcN5aC/HdaRmtH81VY7IEhWQASLRcdsdxUwyRiWz23V3eYzn45++ga5PQFUo6szdtvFkO
rYmVc8YNi186RwKGj3c9o/G0eWpKS99wHZpODGTkxGJIocVNcjjrjqJfdjhQ/iiHNlXrV0g5jcQo
Zrg2nXJyri9UHu3HWRPyQU3yhDgoMRntmfHlpJfAaBzE2mg3Vy+E5qpV3vvCRc1o4Igx0/nnhIky
KzbzCbrBy+jOu6lKhfN+lIkig9Q9xj6wOBTOxAMfZGdK8zeBKVzYJ1ge87t7BD8Cn6XILQaZPM5N
51/N54rqKYuQiY+y91A/cVAizQPwIndHdPcAP1izp3UymI2YsQ41W1qePAyLkyoSW9UKsVE2YCgr
MzaLkZF30hi0+HhxKsl+MsCSoChsBD5NdKSvkip1dkP3HVNsGRmyMqqmUeb6MyDZ63CSCGPmNKoX
Di5TZ6zRXVIshv7v7kUSI4WoxBZ311+u67mnpPzgrrtv1EloKYPbvY+pj72t7+aUy4qYzobUAAsS
UdgZTlHw0B88cItlKqqGCFu2P4ISzgZ2JuE2mAjs0SQuXnDUKWKFigLGBEHJcurvq/9mBwX3527J
GJ89O5unlMKfkMYkU/M8dpk3qdVDxHoGKLrD7iJsWpR8T6DTpWksBm5OD/sHSDWprRU9llssnDL8
+/OmK9UkJOmva9F2HIMBH8wXvs7QjxzazIJG2FHSOm5IaeNIP4xJHeNFfqDSMdtQnimVs+TnavxF
DHgoYJQzTf8qnnxp5qO7gSI+klZJpRIbAQ8OsEPJQzexaobpRBsiI+DPk8HUfp2X5/LtuRjxto+m
5mVg6FExCv144ZW67OXvKT2yBjJI0ol8xPbniGvRRS3sB3I9k+oTSxjafEEw+U30Xs+lrn21QklG
B9X27GHWVE8K42NGocqnCIHkqjlng39Q/w75DH1qhY8GXfpvIR+fIrgXzjBjTizuPCbw/HeGUebM
Iqbf3bl3ttEd8t9ZjhgDrGSO+fMJHqSV1VfYZj4p3tatl67gpPLJkPqZvxH3mQyD6YtD4Ot+qmpT
a4ULsbf/3ZkTu3Bc4Wzz/9I9yXr4Zr5KFuI5c0GVq9zFNACWitZgspbrkEJsVwNM7AaBzhJeKTX3
1YR2oieF/W+JPdYq3Zubue15R62MaO3qf7k7mtYJpBPMhfHarmdygQH4rnlCl56hal2D7fyze+jK
jv1bUOKHkSO19rAmbiVNKUiD3zWEud6l+c2LewfWVYdZosLDS/KGeziJDlRdIonghCJC15irVGbO
DNYBnoVoPrdz4hus/EoOJHgaQAgFMmdSwB++9sLbjFwOW9Jl8i8JbCUR8rRBcS2bTToLlB2V86XS
1WaUu+us0RoijYucV8CR9HWqjbPY48hqDT8BzFUEmenZaAlHlD1F7DBjVHMDdzpHr8tqjTWvP8PK
4E9kbNYxn/+jP2YE6Bcjum5nvzJSBYSI7SRsD0XUGjbj9LEibAIlNFu1nOj7w4cSr2Fj8P8L6BPs
Uz7wbNdee1phthV1q2bfvd9h5xuOBSaDo+PgkOSuar62b5Gu6fE+E6eu7OyMli1Qt0JagBlHg8PF
ijkR2gEFixv42vTs6M/aZDnVJFSEXAZUa5q83SIjG04aa2i668YONdbXUxR1cUdNSAGuFUI3oTYh
hixGuXe6dNvcvH9xnIEkW8chr5Gy5CJuvGY/UIzhIxq7dTXknc1Mq1KNnwCObnMA0qSmx7P4m2/T
Pfc/ZZdGcQC2twoyTa3yndEeKpAjf5RWXAhgC3om5Rgk6eJAOKiHnw3I87OmzPtp7Qf6B+Rt+QQN
Q2xg0k2o+B6gCLw+jrqJSi4F9TvEMv6Acd/PBjDtohip7LjFmJsiu0FTTbpm6ZvAzFgVVuAEVbhL
12k=
`protect end_protected
