--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
igglUdxqGJffuI3/xmwxdIJgxckUPUvwotweP/ZsoB37CMwqegpM2G8oUlsjTfovUes8iNjxkbtt
kJyvgPKVGcZllXUGIeWPmrdhXS9ijBUXuG8zDDEFfFqCH3uAyXPqE3RpbNFVYssUgAT4nf8M1PYA
kJa5F3MGOXUtt8Q1a4efPo1BbaK+6QOecp8eWeHMrfZj/DzKZdRIQ+xspac5MGj5tfGZJwV59LPl
G6xX5iFZIPtX+ILSmnpxS7GDYmH0RLrkuyePK9ox6/G4WHScYbG2YxM3koWQWLmlgRSOrEyNfIOT
x+C9PlIqhUZGFRJ7f0iaqUxsbt/NaBVnJ6uSqQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="DQ7o/PuHjRbzhDAuiML5lngtBXVmZhLDs4kwOoO0ZT4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
JsOjvQXQcralKQMAmqY6fLlW8qvQZuCZggxMBNr3uI4YT23bnqeRCAGNUc4aKL+/dqueJ6ObrkcN
ObXGa/is6p9hvked4djowcMf1I72oatcc2yJWYZ4/QVZT9/KCJLuJDzLCBH8n7AY5OQ+Js6lNBrn
5m++jBOLZ+z92b/9qpW7Po1AJsNYkivu8sgk0mXomLAwDMLWVS132BXaSQxderqcBh6Dl+qwjCcf
8o4HjsMOVKBon0eohtF+gursQ7oHPtd2mLrM+SdsiDTPO79BqLa2vtRmYdbOiOVits9BoFT4Vj8q
MccJB1uWNOFNK3bMbvSgZeCId35yqqyVxoYxTA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="mV0vogSL+T+HYDOnuShgItoo7uj0yQPWxojryODyYJY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4480)
`protect data_block
t6bygUYJIaKS40D1nENnlXR3q+ZtB6nruiB9qcchIJFy+DvYlEUe45+QjZbbtk7uo8cHj7eh/aUt
7RlF9yA5JcUbtnBb+Tafx/XJsGkNVvVsb9ZYV/Z5zIvp/HDDeCdnfpbKTp+fM4JX0x2TGCWdZNqU
WsD+W1i8VZRmr51OvjZyyE66MHclqJ0x6vQws4IUDTSH+Rny81YHMTVA8zfINYIOvghsHCmwyjC/
1MzorYMfYJvu3bkWO0QcJYtU2g393g24N8XL+reJR7+Fi2OZmjA7HlPXe86aKgPXvnvULtG7JTyz
xxGM5RqWslV50U+sJuY1W2ns+zrLjeoqAwUCx46BdHq2y8MgzfCSE9OIg6uuPhQatmxDGdiUNtm5
PefRPNUOOKlEeW4j24rJxR/hp5mSynzGQzxWPJmW314HkhcZnraWGEadsCKmn/Nbk9ton8pVDEPa
bNytCQJN7kT/wg0V2VgevHUGJe8PPwNuZULhdAFZR5C3FZHlkEHZkeI8QXMdy37SJ36FP/jLNr77
CZn2l5o4HKHuHa93bTQ5jIapnAw1/ZxmrBqyAeKtqQgUgYLGGvyoopKzYmy/aaj+qoNKZUxw0YIB
ZBZJxrmS+xT5PLPyhfH//+Fryx1j39pDmRPcLb1QQxoxF8c/RQ1DSvoKsiUoEPOVC1Q8vWkR60qE
vo/5r/nhr+PSBki1U8if0AvJuyBSHzrnVYZPeQeJ3cV0QbVJqsAX7EPBmTq/BohWsz3ekJCA08wf
n1lNZLEs+fczoNYSqHFI7aFnVHjwg9Xlo9Y9cATUiNqO/RCNJ2Bo81yh0ymu8EYIJf99Lc4AU/Z0
BStCuAGPmOb8EMhfLVteeY0PNvgMynyGNQjW43M+Eqo0ccFi85M19f5dR4x7uh2wK7Nytl24TH8A
kTMd3XGQ0bLjH4lAHudhq5A7Ym8yUzmbQ+2vS0+0E2ONIFj+1z3oVpB7no8NIufiEScr554GZjcE
xOSLgb60fvsjPDxtBna5HB/w7BIIT6QC2Y/bShl/7z0+JDDXFkixaCUD0V2xdsitr9MMaAxHEneX
ZDnvxuXRW/FAFZEiYpW2ilcVJww2llXqC8huoPxm6lX4w7hCycwobGyaIdJmsEPSQ3Rv9o4rcL6N
vJyxPHD8t/pn0H7i0cRz++u4TNtC9OasupI2bDASVu+fQwwU8TmvZ6mz53GwDBEimQjaub6W2h7v
2ytjubjNXkMak/NApwGTy5Grbio2XbEvewCpSvTdPF+Op6hpzONoZnxiOKQ8NuwvvMX1Y9mQSXxd
nqfPqmzD+hRlvY1pDfNSn33phNfGlg/4vhBdeZy1FgOkSFh60bk3GDmLZCyL9XULdpolwF/YAgLh
Yc39Z0Ogsmk8Y2EVr6fCZneIQRoiLz5QAph8GnDleWQJjmklU8HUD9iydpIkqnQPjkNyn159/DO4
OovIe7WqItEn3uTUwU5XEzfHXM/ok7UKJoLo5362D+bEg1brFuOHIwXc3LRlUa2hOQntRhZ8PCrA
VQ7RcSnUJzPnqP51uCFfTj3YreSDpTtN/tlC2DL9oVDElydt13i6dwYokqnYccSkaf+Q+9QXwOEd
w+Hmjem7wm1vDP/qsVcZnVRCFL5Qmwef6R5vi1aL8HOEkezrosKSetljBZcH+47hzw3GNULjC7YL
yoN5rOdPQZvAQQA9YIZ6qOFaBcuiVSP9tLPurn3JnVkU72f9ISfN03zXpOFFi2TzswGE8LSBVEC7
Ms1+jpnM/xum7/E+SOGZrUv/H2BihiKD3nGrLqQpttzZ1fTgD1Jhb5UeWSxQahrWig/k5MeytxYU
12ZLvLuaSRwO9/ksQ+O3m4F1vuNSIqza5wCr08kO22ve6WTV3VFi8vPrSYHV3nov4xbNJLa7pd6d
pD+YqLidbnMwAJDStdQ2z/yXa07VRK2f+grZjmG/wiNBpBN8tZYogyW01dp0HLUK9yBR4Hq9Zzhh
/PkGVovx1VuCm/wWKE3//nXns98a+4hYJXJa9H2ewJykoi42+An2jgB27fYOyEbXi00oIg8MlQNI
uyxEByPdbwizHcbyNah9R9sANwMLkV3rfYCnIz0EbrQjsTyXyrg8NUwaKHrIZd0W4wYQr5K7CApP
zlPrk5ufsBgdbpF5mEqVgCzuY+Suz3SBJWvQC3gL9YUy7r/5UC1lYSUDvatc7EzAvV5VnK6Jo85x
Ak36jjP1LSupwsQRsTuOCjlJn37UUbk/dtcgquIg1AIJTGueJNQq3YvrfL6ys4jWDqnmChdhN571
0DX80jGPyasAaDDSQvLS+D/pxOPhKKJxbk0xVGXWiII0uJGpv/wzMx8Eot+LBpUGWMNtgB+J/wUi
iOwGsHHv26cb63C+IRa4Ela3jb94/RSEc1hWESetqL1YeqZQ8rHpO3Fx7xx6ukjDnWEjrzWUjoQH
1bHwRRbAP4yj4wF5FAwufAQK64tG/Lueq5aT4NPFtXSIqG4X5AcechgaNa7s87F1NEa/LzCZe7Z0
xfYUetB9ZuwS2orPDRvv24WgRHHLzb0z69ixwV+J+GxOa8aZkhEWECAMQm/hQGGPCMwPhAnc8Mhc
WgnO6yF5CMwRyT11PXR+ttjJ89526M+zruXDn3G3kJIKYZFv/eKq4qenilihxAqpIhozmUGYnJCY
ixR9xd4G6tzyV3JJnwN7KOX5oF7yR3gUcusapgk66e9URLyHz1IDkCBYbTXUhF6EGrvnfxzzztEB
n4uhMX9D+GkgvzB59VdIyOdVjx/iNBMyUiv2G0gQZD22R4e71dMjvWym02u+DegP8OwjNZYeLo8v
P0UEjK6WFQ5kFVd8ZRUpcBEw8cVIQ8kzJMwa4+BVJK5Gi7n1s503lPNT8o/xgQeD6jLY8CQmtsud
dFPg0dprRLvkpLIGPwpEkpztimRuAN/4Sri+tGkGw6Evc8kSph8fEKXAvNQK9rdqUbxaUHoRZooB
BgP0fKRugskqQfUiD6aHhLPqPTw0CpKhVobJV5vOwH4Ai/WE9lF1ZRNc2jqc11k2+9JKEI+c9rIi
uabXlP/yYjRH5KOPihhPNRQy8xajIxbpAVyyKX4TIBBVIO1x9bHvCfZAjjWYBIRF25WJPeDlHJRl
jX6F1I6LjOKB0pzxQ00J1nMQzU+XscjXMKTXpllbwZFy9nC8FKephRBmMB5di2RyUsnZ0QnVX3OW
0BGhyjscq01QtzNnuK19Dp6KbmzmP6ujcHTf+7U7BkhBuBG2xhYkd8b9DjrUwzJuW9rC817D1fQk
0s/mbU3XQPe5oHLdt8esfg6T7VDVr6f8ag0+Zxphf/oIQoPnwCgIBG2ZzUht8cZ9ExaN7B6CZslJ
aTOa3JApzOgPg3YeR6V6y94CRSb1UZShCw/Rcm3Mtn4pykDcoR3gcheWTetGp9WzqvVBp+DtWAAB
z6bwsgX5AFviFZ+Y4GRoTXonSLac8F34c5LwmBkXIQ15k+yQr2PszwQzC7FuvzSkiZalorg2UjsD
XJFxg07x22I8TiFpVY4LOWVge5eUD6rSdjBc46UpFWAc+8B+9GYCj/CKvbwgANqRu2ZV+hV2Nybo
oYHVbusTXjCRbuSXkA48CdDZGhkz80BN0mtCVHvEofTWvg09ohI7LJU2Ghv+iP+iv2V2Lwn3XGoA
79OdrNDrd6X0zvfWSMHTF70VF2yGiUMxgJ7HTxZCFieYJNUYruijuWF+nZ39hbIYmG0KtiglYWFt
Yx+WS2mxFofuF+WSdm/+CMH5c0UhnJoQ6vOMYuT9+D2nzZQMCjgk3mXlyFuNEmBURbfhqv/L30fo
VRl+4G9ts5LUZ97gBsSgvU0DNhByXPLfxVVjLYNCIKgaqet7CESrh/xsueOTtAqN7KqWVn3FSpQ6
zc1hiLxnwBFJLAs1+y+EPb5rWera3av34jNKOeWllID/OFaWYDvHQcUjMa12pB6dHLekTGfQESQ5
qEP9yO7N8L5XNK0Xx0x3pSizCqA6GVkjBECOfKOhl1A/RWEBM1fCfF66xssBPtsCYdzAGhSK1xcD
usl9lCqZE3n6pxLLgQlwBRpwj7jqeK4OpaHiRn0YOz17z2mgWJ86holKIZ8x/p3we86U6AyHeyXl
yLdhQGasL4MlxtVU43wFInO3Ww3qoFP9mH2ENIfG5ui3CxFx8/g8g7gir2bAn5Trr9xT/ras6nYK
Do4B6doAsKT5+dNSdh2EgoCYy7qjHJxCS5oTlq3CT6QjR5YKG9yeU7xclKYNwSbYFxl9k46zarWD
aXp2Q8swAlIobss9JtU7t65v/7j417vtgeKGCrnQ4zMTravwe9Mr9iXAAZfx7qsw5Jn+97C1diyV
zK7sH19eNAaU633LPv7aIwPr/aelnb7Tg6f8Xz5ETUSPc7XCL1YS2HskTo43Aum3BcU72Up8NwMH
0lGC3PMzTD9awHzON+yLKLxBS6zqGI4fSOsJjpHmO8HezBRPVdkj/SGysw343jJEy4mqbEz9q5h5
hHOVTBSNeJWJ8NtriZ9PzvtAbd5mJgdvMtoiqzyxGfAKRXsJ2XYtfBXbb4aYePf5eZLGMkv/5Kne
TQ4nUqzyV+u67FOYPzcPQ9TGOYgMLmgAtDb2SvzOPiMUBCA69hFa7l0sjXEAsisWovUcKxmGcmvK
UeanBVjXwCGFoIJebuEIvvvyZ5YVGQeSRNNoEpfhprtQ6TMRoy5yaQiEYE3Xop3+6Csqh9mmUfPf
uKe/W7UadU+ahgNCFl/Fs4PdW2pzFyLKdoBbv0ethngkBYfWQK2dIm3DX1GW6GqXAN9Xm2hkZWr0
n0q2b4DPCwW029Pn4s+HWlOiKF+gU+vOHN3lPDT9LMPkJ/BomuQ+mCq2I4q51E1kAwiEBs7qu208
Rr9m8xoY2fg+dpMJxxvbycubGP7zO5ZWd7XEp4dOW4TBxQkUyxmgqkLqDdGVGQj9pCiueiXz3vQ8
CEZarY/OB7spVdrVSuHKXRpD0focQFu93uqWfOkXBIqACh7mWF87pSyuuX9bqMFhlquPNLGc2+RX
ZVhF4A6sDf2vnOnAq2oURPkao9rib2nZsc2FzDMDQ15thB+jix10JFHRcX3sBizXdxabx8Qn6WPI
3wmPqTdjWc8XScS/GEgRBVzhKgHj+Udq8wOE529fig3wqpfJ4rcjDhyI7xJYY1q0CUXhNv12tsm8
m4i9V2oDMQb6bnkYNft7IfBKVAcHJI3wIv/4qCxNfrFwl4PiU1yhR3EUwMQPnbcxTsPCRzHkcUJZ
FWKwFnhNx5I9ORQ0HAFeSlWUHV16qCNcTmU1HXKa5KpihtA7FnNm5V0tbS3IMYYSlOrDyYsmdB88
cc8tLc0y4fe57C6NcJ7ouk7fd0ieXUwafHXp1jNbkP2CgpwK2JYXj0Bo/G1KVCjBuvNOWoqU51em
3agF7isHkcNS7jwcJs0VXdx4uFPr+6gOG8oU3RzFia8oZoG+CmjwKFp2AxhLtvIZAIE2ovZLpEQk
O1imz7GftBIBCuy3BV6tWAaxRQs3i5ATHpNOochZdnfz1ws+p+gdfPa8JW5pK9PdzTAwSvoXkcT8
bfXZejFeBTuzTbeAphdh7LiKk7Z1IiE0NDWlkn+FleB/e99ROLNKTTG/SqspL5EDVFqfc13/fH2k
vlS3/adJzZ4pbzcnACxPyt4r5yLa49g7mYcz2bkVlWXW/k8wcJ8fiikpz33iXBVUcyju+Zhdd70i
+RVzP2qVo4EMEmK05YmbSi3F+VnHbLV54q/5moPUiJqEXTym0q21UvVDstPTCbm3stdWaDax8P+d
9Dov+S96aFepZBEEp+xlkePSJhoXJoDCve8sJIAcrKa6uX0Qb9Zv9QIQ1YIbPWmDQMER48wepbZp
W/2zF5ctR/w0Z9s2+zvCSE87rpHodrg41HVrRKw/quls/+v+E/JO8uFvIWqV63r4fsESt1VeTEVK
Wb1nonjZ4CUS0TZEHpkWiTszDO1TwXhOItouLzPTCZN9aA==
`protect end_protected
