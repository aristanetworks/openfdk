--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
PkeGR0dpQfaswTpOEtbfDwilHLbuWmwyt5wRMHC39ONjBFhIU52cnFNr3Mvp/CHKcVk+4GVFXIDt
edD8Pn5Yzjf0TB7nnHr8DSL2mirR/TJK8xS6eDkgC8OezM7jnw0TN4Yf3nqC3wHmMBxv4SBaP+ke
/wJS7PYG7l/8Kv7+7iLQR8D2mOmo3mGXCG4V0eeiwrVUoYG6HH+a3KtankPbeY21piOT6/owPYhB
aHyN8B9UqXxrMCl/7JBIYAqepgJZkViCGqLCTVgC3Kjqbwr9slZ8GqZ+0DonqU48514BqAizRZ35
twU2pFmkY1vLXHnxgdPsmlcny6sH0kwtNBYMlg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="COQVz7u8+Y/WdWORK0nZlp3SDOpvS1aGCd60F+n2Ifc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
h709jbLApX58tK5mfc79tPEVvrAoQyKN13PA1DfWLCSorLxz+b4qoxbiFrNFdSlHAxr/8YLmiKTX
Xv4FS69fKL/yGg3kJjxVPzUCOKL2UwzMJNCA9D2iCNfE5Jh7MdelDB2guo7f+mUfoeZYysn7NLYE
tjUyGVBCUpXSHTyXnMzq3hg7imcq/ZV6LRfm46pG5GW8wvVld+5T9/4jj0Z11iLo8llH6IxWO1w8
SZhYcxVA2IucRnGZDr58+w6BqULcqWQckKMZKIK2jFg5JaZ6BmHRpuA/evuupzHgNkyf4+NPJAot
zza0MtpmLz102cbVHe1lqZAiVw1WQKJ+v46toA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="5thYgXG3Gab1dXXJkTXqGyIUdUnR83ZaeD5ZAYMukis="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34928)
`protect data_block
tsv6bPs7skjU+VNUDFMqzURoXa3eDYXxsIPq7dB5GeUkmt4MJcIFj5PdiRyjo+tpOt8REqAageoV
WGqtByS4GdE8+HvLqomD4yuabFsRycI1ErvxDq9k9TNJoCbVZ3a/Dx+nvUZfbCKDqPSZ7zawtcas
leNL4c3F1PoZ2NJena7Ee4+yLoPjo8jEEID3OkyGXtmaJxo3+Rv0TdO8NZfPjJH+8h8RvR513C04
8cuRlnPM3z/O345x9pQmg8PBmgOdo45krtYYWuw9TgMTRTdUODt5SueFPdcsy9kgbqWhPvE64iWe
tAoMjJ+O5VrbSiorkiJayz5AAfuTYJzLA0PP2uXo0Jjs6EpzTTqlEULQDmXxwn975241v0O7bs9s
W3lu3p5izerw5EJdAvmk0qpA/igfW7MUKcRGK+0hOux1sUCvUwX5vcvu7fvB+qdTtZQSVy23Ub2Z
4WpjT1wQGTANDepvWLc32TcYNl0nEot+UxFubUbhuUaBZ70fP65Xmb81mGD9U45bPoVnIqbcNQGg
D+IrUxcFcXnuDgpQ4mrR0DuePuH7Qqm2L6VdaW4ZiJ2ou6mOKhwIeAc/edFL628CQIsFTZ9He39N
BvIZUChuC9DFUZ+6HhmXD2VSQ9sobPTcufN6CPK/XPz0BxBt3S8PIHlqbqHZD1deejaoYNJc0w+h
rJiUVMGMnlYP12zXHkgVAOtT2YdkZdKJBRKuWx2y+cUYjFhTLZKlnXGEq1V6IqG9EXPXoT1XlVG6
E22mY66e5k/b3mmeq+yr0vYUjba39CNThZ/McnKpK8noy+EdFUsP35kFPKAZ6sLRKa2rwhXmwyWI
x14mFMBbqQbnpaVVcf1NNEgHjJEq/PbcNkVUj3CG6oIs+UxgiHfN5mlTfm7aaVAKpiFuxfDNlPk/
2tQ7tnXC1QI5NUsjDYjxxSYSoiRpAK6CjIk/KcnfMBPRGzVj8irCs9fhsK+xhoSJcMY9p7otG0EW
39jpk9W5q1/Toi6/c8s6BlqdDV9d0lTuSJgxHXyKppKbmnvuyMGLyl8IRKRxdzayyRpLMT6cWK7F
TYFqS2ewNeiTIJ9S9piZiCmaiZA6UJvz2VnZdLhFn4ZpjW43l8GW5Gmew2NEI+OnoSvgFthEHv0A
xUxQVR908MFq9hiDJDtA+AoD6g3QGeNm+e+sPm+oyJ/l4gFHm0fexlyGMRn8AtSvEO6AdMQYs4uj
b2FDEOBd10TCA6oGh2li4l9QWqKFIcXz+kjeKD2HhY0YKKOpBLaAaXEdhu6uQ3f/n1nIi0vZ4SfI
kv19ZfhYPRXgvwgMr7XztSWYb3KsP14r+FRnH2qk3HLMe+WlPaJKrByfPdWeuiCxlR5t1FQ7FtkP
NShFQyMF4NP3Eg0Akgl5/oFP60NzfvXuI34Yg7bLgXRqeBS3OWgwfY5u0Vo40TAFjtIO+aucM49x
HgTjACfjXyFxoDZbzxG6xiQnWYEabdtS+s0GIP7UO4IGXJfR24uyauhKxRiBD3M+96ZAvzQ1LE2W
ZB2g/yqbig8q13+GZakWwXwJAoIxy1xNC0lQhYbmWLwMLeFdoOSq3vBF+Wq5rwTz2GeK3Vz1Ulpx
XbAKqrx7PXZtjVG90UDUqHES3W5nHPSz+76siNC07H5lrqlr1FaLwO8Vw+NOJrb0X5hmd9lWra33
zWbXL77LtROoy+jvS2Yc9/gs2FJKEdOZqEMI1TeNDuHLuhJG6unpMj7nB8F/8lPp1bnxjsRMeU/I
cMYIFSQ0mqQnRY2nkQdphfZccDF23mGI1bl3p8Va3vwxhZ+mAfjSEAAYYuojwyif8LHtoD++NrBp
Rfr9FdabkkVUL2YErZXLn/vy9pkp3DnWqt4lxtDKMBlQ7gqEFckp0aEGt/UC0CH17eLsmYz9Crib
Dl4TymREjJk6QZxj0Y7Y7QWm3QUZanuZXZImlmDriYSO7lPlcXt9pgk7yS1oLRUXUylCSdVR27ym
Su3GGwDqmfic58PgOz52J64P+Qn7MzurHDKF1kf22bhZb9DU4qM6UaHJcQgHpQSRogQimIzfg0TF
PQZWD3J9SEAWHMOaxxBqOVgaX8ebfCEFprKFg7+CbfSJpxt+lH7RoFAbrOL9VIXrcEePb/2Uts5m
PULgC6INdznMPG2x97v1u26n0yyQ2ZGY/bhEJeRyGcJPbkynR3IKkUoYy/2NiKrQY9kOhuvGOEg2
EjW0lJqgCJtpf52S0RwxJck36lAkDgyvNzEGx5crk+qd1JVj904dZHBn428AbYAuTvRPrW/5YYlC
UIln+6cz/QYgJ3TLSBJ+C6QeQFeNp2J1I3ITiKoRDhhG2SS1TlDauV6UsxglEYiUYFH+0z15SNRz
euyMNsmK+GXuYOyDkhflRBH3+P7CsT5ytZh5kL+H/zEYFL6yXw8TiCj1p6DM+EjE9qHc0nJ/03M+
V3LncGNFVo4dOjZkUoK54JRRlvOs9tkffjALousw+f9cVoWp7kWaKtNfQwo0FKIEnhMCDoS2lF3H
a2Yp2d8HdmJCmVmGH//faIQjCNu1HizhWoJOOKMVu3d3A5g8A2pNIObemasI4DNMjYYh6F/W1Y/Z
5hLAJzFl6sNo+ag5/AOYrCVs4YXADz57+Y5CsAmexDCU+EtRmljldXrf+n9CIlEu6Dd1e+m6ZdiZ
2mD28ngfIJq4CEA3f7lGWjHjE/S0uEQluhqv9EtNtb3sg6Z96fM4Ou9/0TNbI8JpwY7WGS4imUEs
uzCvzYitx0Q/KULbNxJpeyaoZlSeyHMHsHnll6FXw1KeImvc6WKXpNOdowizHne0l3him6eCQ2Lj
/LmX1O/NWzoOt6nAsMdc+BUbLNfeD7KyQ80snl71AvZomHhgS5BmdJmoAzuD97wsFXRvmxMlqkGc
JT7ijnU/oBD4xXLrUdBUQ7fPwMyJxjnkaSm1Ek0RlSIzpG/kG/VZZo7oKmvpuBgyyplD/l4ZPgx4
+kH+Eo/0+mFYaQDYyW7oZGmL97O2WNYwige/zleY5hMJEvPw7CoIAwUY+ggy4BRZ0XDVKjOmb0CZ
hIEQiV7ughVJZZJKCKq/a3RPnbtGQDtPecc3kkTTNHmN8lpYhqrXnGEdYZoKZAofTwWk6EdmAw/I
58veZcFJDAcpUuCiDvw0mDSEMpP2YF0ZwU4zGNxTmNB27WfqazGuv18y22p0Mrv+nD3pCRk0XjUK
yjobl/ei9eiS97wn1eQBJikFhK09dLn0B9m/V5chwDDUKpmY2LNrWrfiABvcFq/CXTp49Zp+PolE
L4WEJvG7kBvx7b0uQENkMKJmhn2AS4BB7M4nXVWSoV0T4scWg/5dYSq4S17lYKVGX+h2dW8uNxe2
OoZrpmDdyqeudhylaKW8Ft1eDNLdpgcQ+eed6F8gk5p8mQT9h8z9ydvO1SlBWcCbE+CHkW1901hb
rt90GtbUjLIHo1cr2c/Hry4n4eE0+ZgwYnFnev/em/VAnIKfDTwgJ+BhMN85IbUddNeDUfOeJ4FF
sgp/BMj0gb76JDMTMdjYlZiAt2h+SE7/5uOZDnW3R3KSnJAilOup6AmbQzN6njF9k+eEInDlQEPQ
potPligT3jlb0emwpbRDOTjpYH77n6YG2l8VuTJyzCEXXVBVCrcxgvPGqL//7+hKFcHMG3IoAm6W
R14dcQxWQg7m9BPPrdcZV16qxZiHuDS3eRKnhDaGugzCAireon1gv/6Afu/VJceGFdSBpWtSQq1T
tLVVn/DYRv7rD890ESHRfL6gejki4O2rMiUvmc70RsemARd1/IvR+h7QZrAnIO9daG3e+DfzE1an
lC6KJj79wwDVzbvbqeGvmMZfAZlu7RKQXB/WkttuZq3Qetn5EMHMmo+aBxxAP5ptGu4jE4296wKS
s1nU8euByU7vCYgmvqEaobquNzptj5NKL4c2RSZJdQrYXDxV7Bebz+ZGYOg+mSYckwPAl7qhSRM5
sl9MtMZCkT59qWTvdoMPiDik5/aEI3oWHMYcgiqA5JHpSpjiWcOlVBvr7qhoonr/a9bB4iyIqZ5M
+yJP9aloD7YKuVyKo38/Bh+oEaTWqgcpJpgA0jZvAcMhkwdzDavJ+qR61LmItEmHEWpZNIdnFzBi
nS+SZBuVVc/1oYj+hxHo+KJ2jEpEKhmww1UQ4eZuAcOz26Bao5ik2Q5AvoNlE4kgRyY/eoGaFTYs
XQrg9yPHIhAzKY/uX9ygjickG3K1+5enlF5521/3gcNVcVwHok/0TjLEGGRUWg8Kh8+CM9G+Tlkj
EpL3fIerFYNQgFqngiRQ+qtiwGGVzYY3bus/xoEusSpCEK3eRNaXrD9je65UwACha9zASSWgIUaP
B/YPteTXE4hLsPI7AiTY1HAv5EVLevl3WZCuxEs//6Mp5cDLBtsJ/Wpxq1HOt/F36lzX4gOnGceP
UOMeyNjiGUPBgaM2IXFbbX3ZcaBQqe3Hs+8DMSe+/gOTYTcF7kSH1ZIDpqhMPjjLMfGH1+Eypjn6
35XI4e94qSgmZcxMGOb5xBZn6ee3IEbK2V2oBCipsXuV9dIl4oiW8x4LqYqjWSdkHjz2p8b5Kq+9
R7jZOtwjTRfofyHNhHxhTS0Nfn4rHLqIdRFC1bTXGgnZzcDHM+mWRbkcNdgzflIkyXxGJ+H/giiO
3pQ471A5zNGXgUfjDwcfppy69FXo2hk3WftQJg1PqbGqPPc7BG5jbuufq8qS6TOeZ8ObJz+SuPY3
fhX5SfYA7H3cf8fZQg4I9OyY6Y9fS0wHagKyP8pOkWxoEGktmMI/xfQEbLKh0zCkHJrFa87tZPUL
wsqav4B9QMHwMLomPFo5eepe2f5G5TuP6YFBHjz39FgNs4MbTDhen6L0dOBWA7gCraSqC2L8yc1J
K2wvcuD4JWGdtLLParaMAevoJzjoUzWv3doqMD6jB66itghCu4Zz43ZGTCxD8QofHN8LJrfvFr4e
z5HK17I+/iPhn1fqAeTbY+7hiPTLVtXeqM69A1LTGQACw6++ocl6UkxZAjOMoX/omO54KeIORziV
gsCf6yqPOcGKt+xZUVDz65nnr+NxQ20ggxGdeH3mL22sUR0GG7q0gHKOVBkPHoBYSw0dh816/2Zz
qH+LeSCm1GI0ilxEjAI3W4+Bs+4aRxgcfjVjanI8gR8K+o7jS9/Cc+0peWY/dzUPDNLQ46FwFXM0
1anf3X1mPCwGt+f02PzQdazDe4QtBTyuswKrJeXii2+Jr0MJlc8wbYg6eiJDIeS/Zi77xHN/t4IK
H+JDnJ4z7uadQQo1tej6URKlvnWK/jMML1Sasl9nl6hMqPyVhoz9wF4jBKetmSr9RfL2C2RQdKf8
zjrvglHgELkA504Jf3o1WzTpGpm7dIRb43QKThTFLi9XZh+bA3tkYxRiQWD8LmkFUhpIzVWvwPnA
bh55SKln9a/GDHUytZ8lQ88KPK9sQwqkFRBpHfkn0wtoXAyVMAlr0nVlha5zdRBnigmieJ+NyXAl
bU1l6yzOj7jK77tiGr37UgRriQmQeskX1+rCUPIQRZnLetua8FQN9YvGCERv8Pv1287RpPDtPP7p
vLtcp5cfIt89t2ah48zPAShbQf5YkHleQrrwUuqKpcUB/aCbAcbmtlKxCbKc94yS4aBp4rZ6GcAh
MXfqgeEjIwOMy4+6L8Zu43JHjr7s6ajccLcD1TD0E3sqNa6W9rN4bopt8QL289ipmK9aY01vFkDq
S2GN6daJw7aoFb31Y5P0v7jN8bJKPz56cJ7zqPCFpo1DwCcQYGbgYrXNYNXwOFzj6N7FpWip0Z3b
VEtZUsnoBQIoXGgihS27I+6Z/A7afPJSEz7zLNG6co27TvQoDYtBZH6ScEVh0WeigftmCAYBgUOH
0MSHQ3HhwsA2TmjJj4X9CH2/dlWPgQt+g85oDDH6aDhEIrHX67J/iGIWboWGxBqxjrpZShQ/26TL
k5pmN7hutZuGTWUuw/nKWVsaTu+j6+Aq0v8C/MXBZantRqkRmi+yRKHaiiRRifhSFvWLxR9jeaCe
W56kPqlm1vkuv4ekxfRls+JihCiJbHIUnKapNgIuzHTHJU+nxnEnmoYTNEHwrclw+vkw5fe9bLQN
xRe3VYhQyRFM2l8q6aXLpvc7fJUGDIwWtHK3Fagf/WiVWvaGxRoj7VFufUbUzCssUXbrtN7a3tbS
rsR6tLbQD2VcN/iGUDscnixqvs0j5JvkiUsbdfKXJHK36w77l4EOnu+4JETfD22cD0SmhrgiMrVP
ECKLSwlYH4AnOoBkzUEfsz/4qSwntHofqwDM1NdaQJFqvMHMopy2VWUsU1hkmr979nqVlvK3/anc
T9ywqt+BFJEd6EcBypMEjtOPqTFWGYf+zIpVS3QZVna8HvteJPPZYu/MteOeMkQzx7KhWCqwJjar
7UXlRd6YFg+17EZFUOr7SkjM+vWTgnVTF3Y22ltMgy/rxZvp7xZhEEBulJ41e3H4ciJahKpSeGdE
VGSLu+buVu4DgiIWBoV28kvZO13ylR4iopHSBY3BI7XzSicJ/xNf4+dDDS93PwFRkZD0CfPB8bEs
toMJi0TjPXKuvTbUJ1575kNVwyYLYUdWeo2ToYZnfSW+HMeK8WzjFY0uYahLegk6CE5/ZHemFg/F
vNOVOlUA+8cL+b3S+ZANcKOy8rATWN1str9zzXZXWRqXcO8ps5GhWQ01H4mQqjS4obtgaHc4vdC+
uB4dOhMm1DR6oS+3Uhp7JScrv0S1y4Y8cM5D6Bx0AwbJ4c1vPKlB9vb+ODZZY+EDB+xib29zTO5D
AIculcSOSlpdNqKQjJN089eGzWZ6kvB47uutqEs+G6GyxW0/Vmahe73ibqtaVd9vM/AErbQRYC+w
zmjc3bps4ef+Cq+1vjU9jA8RWSanr3medYuekNCk4v/q62Ek+htqordj1PzlLbcFce3H7AQ4ssuh
iqxjjYPdJm81QYBHBrGaQejzhTGS7Xy8giHNK7rv6HP/3/irfFxC577A664dKiQP0bQ41mh5J9Cw
aKGOj111DoTtKWF9Cns0cDFS+tC2JPyfb2U9mOXx1dzlOxqDnE0UcynaH5sFWnDTqXnnrraVpZE2
tDg8Nifb/N3smUGr/R+/oEUfjJzU6NGb5F5jR7bX/HCnWBOdLvC6o6IchFsNcohtRQTrf6y2kifX
Y7GUC9xSd9gVCeO9kcQ2+x2yQe/dpZIDgbG9uZoJNy1KHbz13dwmWtzrVwEwHXK0Qyp366mv3dgO
c2ODA/RWAWCWQk9kEnUcdeH89rSn+CLU+DCuIf5ZUjWXoQrFi0ZRsc/ldI1ulbpP3q9vdFbty1yt
K5lUpyiwuftI7Nzy5iaZLJkuJe53VjaAOVCwpZXBifs4IvIsritX5pBaUaJJ9AG5Fu6V87B74Icm
M9camdb0K4T0oFjTBED4LAmA4GN/d8wuMILYTX8FLl6qpmpfI5jnJUS6qA/21cWAbk675ueNY+/0
9PYfa4NEwJ5JFc7sGvBKMCMmmlOAC2a0gJ86I/Jeu68vbrZyx1FHR+BAAU0edlpA37Q2A60uqw0l
uApwVWK5fZkyFkRbVxZsdxbS1jeJmX8CHDF5JGQyNAIAaLf4w8YPWPhrIJ9EJ+pmOZ/ANuqXqXfn
kHroPQwpScFdY5VvVNLsg0hBKZlELvY2+OjPp12E7YhHCTpMqFnIWM1eQ0CQs+oGIsyP3rky5HSk
x7T4U+Sh60gTvPmAFHDchAabFuTjFyjDc3VRh4IRXHZ4QgzVl6bZ4M7yODidAsVt0ABgB/aA6N6r
9ngnRELau6VNyoYiryCQaOOExg7TDKhJI3erPuFfpDpEdzwuW2ejWim8Fs49mU8ry9Bdpn+mcRvt
r9VKSgKE/SRoZBeCXryxxu5YB+3LrfHOJhxdwfGx9u8B6Yc2cITRFoox2HopLRiQAiWbSmc93s6i
CsfMgohoEeAfwzjt0TTBThBPSg5mT6EBgnD0sV8IM0T+LFtxcy4rCOAvtehbQywHo81FcJOxRfBw
Yzhqzc/2LTJmurklGf9IEzB99GeeUMwpqf7vidcoGO2gGctHqxnJA0mwvU33XhdRnKfRiZAx6yOo
CkJnErbTamyJbk3mQ/HyyEfzS2gXmSSy5G1wl83SsuBhFI0xJVoAVKcaMEBFklX8KPF6B9JPY6iI
BIXNP2cKO4oFp0/aweX2TCEy/pRx7est+Eh69qgylsGMczPw7n4r1kboVJsuJQEPVvEy1iBSv9fB
XO7cV9nGMw7wm18hHVQvzgoIwNGDvCAtsAtb4GnPwkotiNP35A+zgp3axrLehxl5U3nMvgbNvEwm
+6T1MK3iWTM5vUi/rcEKmeoE3XbdxLMHTJilr1cfvQN7B6B9e54Q8OHy6S1G767sJAf/+a4wRsjp
VP770HBRCTNvevgjp4H0eG+EVb1LjQcqmz2qECG7F2oLwfuZ1UeiE2xyAvfvbUdIt49lhQvtlVYN
kcY70TYSqILZTYK3rduZ+zQc073bD4MeMwNxNXJpgfd36023vQM9k4pm7GU7YXc9SPNs3XtGi3AY
yI3CYkbZQYaSZF+WjY/fbpZ37ouOM/ZPU5Fva4kq8XKbYlxEIIrF2olL85Yecp7zEKQRtmXUV7Da
bJ0x1fTqGRDgPofHljT8PFPuKeZWgZX5/mTEQcb/s1Dfm+sZ/bpvOWz6eHlOExaM6z+7a1Nr5A4i
qpyICJxzDa1fgRBj26Wne29DFON5FygJVpp627bls8pXyqLJo0he5U1+CHkTLsWbOSt9EsZAjmLB
7NocZvt2dATHLAdADP9qIYu6gR+povgKq4SXwseQyyyOtIr03l0aF8XdZi83w7sZH8IBe/h9wUJC
fiCS7Inz59NW/f38L9sQWmGYC5O6+ovNO9rQTQVnSmYoa0o80bwUWCclRP4t6IWAD670JuDMYq84
WKSaZjkHKO59XrzTF9QZjRDyJKljUWMmLNJp2nL1+G3U0TDuG/UgJ3GTm4gRCH6S6dIcbvxKmSz5
fcMhrpcKzQEfJ1MnS+DYX0Few0st+/6YCbsurh6wE2gsMmn1KmUXk7crRUY1K5vsbqRHsWy4+19S
sZ3Hl8FFqMVkeQw4rVw6FW9tFATPFs6HI1GRKYZerY3xoVdS6rCgvAqgIggQOkexWM9rE5CC8/Iq
6MrjeHlJhZJj8a4UZomrBNSwj7O3g3jvsX0cFWz/ppArxWEZLZr71f8OE88kjvzrK81HJkh76uA1
Z3+cz8AORbmMqM2O8ZlFppUqf2Aqpg078xDbSgyq3fxygNSV5KS/kmOOizNf3AGwraCajk5MVjZG
dkmGFf1WAcgEqEXGpdGyi9kOGnHykaLnKMntE1YiMhGkuIwM0Jes06LlapnjfyNi0X3pq5qEoJew
gS5TDhfu2PJm2zd8KeElb//2hemvfjsbfhrmgpo/KzP3QveawSS4ewV7zo5QQuwKG3fRZvCoCARd
YtDAziFS/7CWwfrCN5X6FEISg4KVT8okJcPCOQGG6HFHzumTPDxvzI6w28luzonldlvdqj6Q7ewK
tvzB04OqVvNUZu8bteDler5JHAwCrtJvJKn3u90zOxoaUXFVdQFQsdVKxKLooG46xV2ISHN13W1m
gZzJMUPzhi0cKLNbfaiA4PAbEMV1IDHKCfzu3FT1tUQ14+R423d272kUAakiQjV5S7/H/PrhxPJK
qMfGL2hnHBV6pH4Wa7MforDXKDxcoj2SycpXAqjl+bnfSo3luybZUnKJhtWo/UEbXQdyhmc3TYZU
cNnT9vPR9SQkiav1mHDxiR+OPfNkgtPodvbGARbCXQFTGfcSRy4JD/MP3s+a8nElqd3HRfIjxiNl
ueudn8xFmi2b7lhPJW4XefILDOmdWAnuvAK5/p9U7sVtvdZH4NjeWttqueLT72alMzpw3gGhnMCW
Rz9NDSjkVXTaRaJ1aqORY8xzP10FEsEmF6YZFQfiwlyqLo4F/C/K2yGPAuXqqtUcJQwg+2lac0VQ
aAQZ6blyXxHfm40aBrTavJBYNxMB/SEhvAWncBQ7vRNwJ2//SB90YfyxVQ2zRWBi5insUjH62Plx
ceXnDFFoR5IYz6GUnGiTuiwCH7M3/KrvuSgA6f97yuN+smrTpMgr3fk81G2lnM17tjnDncWKMxhJ
8bpYFKfyuIMTuwxQ2+ZDxs8sG3kZNHcIf3kTPr7WCEcV3XkUGnfxEAkz9jBorkkLq8/1/jEjaC5k
gkO46axfPPmZ6zQqOaHb3S1gwGJ2jPvwVANZMxzjPUdWgunac6wkndRAN5moSc9uSrrGB8QFsdnP
ae/8HCAqj/XjVBlq/CAv6wUvO2DEBWkm2aKfEZBiYVHzsyEtFw61HE3ode1UMEKscCPIRSCNgA0v
USxQQOYjcfnEutA8+k/aqdAwjBDb1REGNo0jICRD44lfnouPk6+J4PRsnxCSKjKOJkDqJBR5dZHG
pKGnsmbvP8edw/fhLIbbOAa8u7dJ7d3aS1J5skfkZRHMR7TGyY+/6fWZNPDj63uXjSs8xWkXdZWR
a2iGg5GlhYaOAV6kskyrwrRpfVjI/SBXW+geMRzVg7OA7amZNX8uaJj9X+uga07QcU0Ds9BbPJR/
VxzD5CR0Ur13PVTsp+DlUVuHwp6cC4rCkysjC7/Cr4EJfOJDJlgbWOiSPdY7omM4+s6qCOMy3rQ4
qtHE7BzDqUI8fhy+C+9QqLZjIx1AVO0Elx1pY7tDNYI1D/s8M3zsmx5S+VFVA6jEU+PX+W9OqnZS
bfjWvCN13m9rM3p7aNhTEnh7J3FLzGSrUnSHWYCjOtL0lF7oqd+Bs9BUR5cpdfk5EJSHeC8lEJw/
QLP7por0v+NiBjFXSamoUMqG5Z5UZ0Z1d1mvICgTle5w6pvKuJACi/HWII2ADFxJPsVH3r3ZO2Y4
7FBqi4VXAmeBsSyftmJKYsd+yA4F9/Cmg99RyUW1kdNEXLV2dZhL40QuHt/DeSTZ8caotGlpxRl3
4GUbwJ0DvWBy1zSDAcld0DmTY2AJ9DuV1muNaGpNpCBSWBaZrtUpg857ivvHymY28/Olth6dbmn4
GWyOvT77uiruMuxb8+dxtzNaT0gJA+gbN9Q19M+g9JvaKI4yPCAyiMaIoZzkYIkVPtWnO+TCZ7NA
COcOzoFqwCBjSADMBV0WaI/xn+jwTXyeIz16RJNaIjzj19rpmUy42YZ1IOBHRCLn/KLXzxZRrkGu
QiI/PiU8P4Jb5seIH5p8pi3kVb+MwZCJiTqvfFZFOx9iTARxlNLmRPn5DbNN14OekgK+vRlvSYBF
eLvPDTMxk6Kzdc7dZhp64b80XiPsj5uIUiTe8HM9flrs3G08CHffV6X8srAghJPS82Fu4y2CKUTG
6UAZsyjh2V7PQFKmm35TDNzuNEzY8faWOupIcXlNQWIW1K9PoxS6dOc6s8UMfRDlAQi8yuSgKjNK
bTMZ+bjzqtaHePdzkEq1jFIIv16NedMloLE0tiOZIAM1aqf+Q0hmqlKuQbsoY9fWjJfmCQK10OAG
cSdD8jSLkTIXESw5LP5CtMv39QAZ3+czBR1LxC7oSekiVKYLW8pchBes2Da6AQL8wmLmSUPf04iF
Y4LkUyO+vaepd3ju6p1P4crsYJvqt+OUejSReFRbtIsWTILtLbtrPuDzE+QdqjsfkhMq1+vUF7La
iRzQm+9Kt6KyG2OV//86Ek1US7afI37eXrdDvIaEfiE567sYiCdLkYzlzWqUG7o3/gTVBWxKp9xM
VHxItxeV4W8X6UuaPaXBnhRqiJnjBYzbPUkM4awkpENkgLkmn2sTbVBH6sKC8ORTTk9G3Q8Vp56w
aJRq2IVoP9eGUZMtNAAEONzDmw71YC0v5LAJL+Xrf59GrtEuwEvnYUX1fzENsZhMhshf5jt/blxN
+yUXj2AcejlluQISMlYJ4NPFeb5hFm99paj+PLEhgcXCZ82X7iQTL/2rP6HImD6VSdXH2dklJLAm
+Xovq2yFWiTp2ssRXThUt4byP3v6WQvCOvwn/OFcX4U0q1E7f+fSsFAI9TuLTyDAA37cCjB5GMpL
5fFbpRV+3l6OIgkX5Mgex+a1usdcFFi5cQ5YJLgeB+lOMgNBYCLwxltSaGTQjHBk8D3I1mpbdGXq
rfpMXOQi8fKjjIjrv2sfZVVP7FAWBWfuPV6TYOB0Wf62W63agSD8+mIwAqhxqBFpd1X/42mB5IRz
8ghp5tF/iTc7aqLlH3bhQ6Mv5GgABTdZRLhDUVqFq8wcBTkO0dq2msAHXg4WhTzb88jgzuAg4hCs
tGasWSljrWnUdZ+M5DZvCfzE0JHXN8PMmzWOM0DRC+u1BjcXGDLSVdSYJcm5iGkmQ9xx7A4h6N0e
2Vl9H4QXtqrASUBECTunvL3TImEW8ZU6wKM01Q7b3fSfbyxyYzeF3MsUXzF0fv9n6r7MvPUfzEKi
zrHbd6q63PHpR6fYGubEsYf8ICpk5jDahpot7q4DnxcLIq+Shw6Vcb6nR4psOI9xdhaa3dmvxgtR
QASrm+Jz6l9GbwpDxCHLh2KrAMzD6UEduHh/+6KOX9QVzdwXWp1KZebFpZIooJPdt/x2d30FzfnB
3BRec49SIzPRDt5mGt9Tnd8xznLhZk/lToaEXt3JrI280fGDasvPCaQn99tsawEfL/t9z5ycqeCZ
D1vwYQJVDFbGTx057ENSXop5doffT2k/oxfY+nIbvZFn4jJMOd4JNGmROGn2+DVf4U4UFW22Q+E8
QgGsQ1t02H47hcybGohheZoE7b+kRnsIHevxbuSRSSfkehFhWDg2aVsNob0eVpstdpoUF+4Mbrjo
inKIs5O1p6o0alkjTYqO0qAQTkPhgTfuSvEYSZWEzTbeGHUDJuttVM9Z8GxvR3cCo/cmqQV7eYKy
bg19lnMmPxlsemr4oQn9Ub0a+kNRyz6KwjLKHU+3fHAW15nEkGstZXsMFf8e2d9zCdbKpTvt0+0r
2uslQud4WdhD2I/KQz2UPd1chTl99s39tVF8hQNXq26OGf+qTJg0U3k2C3JmN94mKrOR2MmVpM6B
r9Y4gB21zm+ZkZefjOjchQZVk4Miz6+JdNZmMZ2j0vWdluCz3Gge+ttQSPEGUJb1FVbDI+d2/tnU
KZ6N8VPGb2D/YDY6iAYw1/6+MXPEqAihiC6K29QWHH8HsmsNXUJjaZH6Klzyrx/7w+LMXkDRvwnn
Tnes0cEXiyMcEbvM7VmhxeQs+i9Ky6wQU47bgZB10Q3bh9mU1pPYZ5MOfwC9sqJl0VsYjzqc8GjP
PPNEqvB7nhSURPSIp+lf8yaLNrJy/zoX7GCiXpcGN+dCRKogCZ0woqA7dklGhiRvTvDD3igqXSZL
ttis6NPX0NPhJA+pZiNqru3XMkwrMJM/ibN1QeyyWMWIUeh5VxK+vkn6VVQghYuA7TwOiM9SNGro
eQsfOmKcswyHCk4QbqLBzrDGcxurw91xvW6pdCu2Az4K4WtSkkndB2h82iJWiBm2ZEuUkZ/GSH02
tBM+hUclF35M7eFHW3LuQpNZvssg1D7x7MNvR8Wj4whXZ8hHDeZtoNgj7jETBSO9aZZJFNzb3qnw
QDd4azZjEYdQAihJaRFvRFXjsoz4VuZcKBX2q8J/G5+fG6Luqr9/3CIwhTzZJoQkj4HuNszKYv6v
rPvJhbpmLfWVNQv4akvkpbMvt3LsOoEchWQ3GGsFdFxQXOPdPGBZ8u4PPJAwQSzWEfXTwNZMcpKw
321s5wOtHZ7hPB2ywTjF10wAoWEUpAKHQWy05co/usqNaNnyL2KKkBJpMfR1hCcSIeXpgsOXDJuf
J4UVttsCUmQC7DQDJIj1Q42hFMb1QP5soNU9o1CMvoLQ/11VNlN/vFIyUF99XSise34QypWwiEO7
aj9ws4azHMln9rEXoE2CKdAYxwRrVrInmGlRkTWs9CGmeMjzffwYSzEiqKjQQUU+zKRA0VjBrkgU
ifxj428ALSauRD0UJGX8Nmw9R2iwLac7rXaxnjiA2Jl+q3kLBD5yy+vGjo8B39AVmybw4sHNCouc
9sQ3Z+uJhZW9/NtTbNlNY+CzCmPBdz5l9tpNorUDWywTIlWizGqP/x9MRVS3R9yCTF13XYSsKzRg
TLlWJTUsrVn3ewdtys1TckLGg3ZLY8h77pZY/IC5oZlIR1lk1hEApsdj9aDtpLNfdbes8h9Ou83k
zHocPhFAgMyoFUMWj9lTr3fN0oqbSofWQVV367ckLKMun4GYeqtA2uw/Bc+JxQD0h/SyiF1aHwJr
gQh+u5hRMpI6sVcDuH47cyH99SHmwOV4wrzUASh8YoS/82uoIyEXuKdfCprSVJxAwSOCvFMQbJYu
ST1/RKj3nErgiY2MP0mJuuJQvbr5i/4uY3Tk8xT7jLdplvLA1nP9EdkwLBQLjTpMQF1Yr+r4B8sb
6PJEbiLXBsPQnr/uXtWdlyiLoCLBWxFggdXp+fR2/lnc7UytkHapUNL+aVoJ/vGFaYZ1ca1N7i3v
bvCt/8PmyeFwgkYuoE1/M+p6t4QHCR7WeGkJnRW/Dn4pJUwL11M6luFQhQE0/AgTTc6XTjtfgJ7Y
rofe2MRSk79w2hUyCfMb91q5v19Gc3GN8hz4k2p5VJlq+/BEhd3L4mB9i8FMc3hCLPwX6AwQSnma
XdunXza0OLrAaW3mBI2/zx5CcYUH9LVFjuhOqwlycImMd9KuTUS/e3ePDrn1UrAJ6uEn5szDtHp/
Mfwsct0GcCXJMVogeCjyI/bKC5D5+CoGaym5OmQLAlzDS3VV+0wkjaVeIWXa5AF/sqvoOlOWvE2A
/6hjoDAxFHob3hj6aL465XeXkmj7sG3qQcG+koqSHj5Oi0/GrOuVytNzF91b1GlsA+rsKVn2fBka
vXKTY0KMUsx+kYymAoOEcQhNUyG4TFNTO+imh49i05ku+w7FwkN4LTqCxzuQWJAY/cXALSlssq4e
YeypHgho/3Bvfj0sUAM+Pjg6oPFKwshETAI65zRerhSMbHo3UIf7KkoI5eEXxOU0uz96byXEdyqh
S6kKLcrzB/j+bSjRZRnVI1d7+0ykJ9LHz7rJHdYT3a0HQnh2lzech02gR45jZOqpKWhtnswygLXu
CjkXjptSkwxzwyMXInx9Rn+5tz/kr/JQ769aR9C6zoT0xoSynUyoHzEZdYdfYj62KU5SMIzTbJMN
sRJn4iZG3eCqpdo8EJhaGIbG7cPVezzAOqNskWiI2Gc8mTRCFcnFFTGmyhpQT2XhbSqAxzGtvS4w
j1loMs1NZ84gn2VheA7qr72k+BF7oBwp8lcfAozXDG+V20dHkVKYtNHlxTdav0ue6oBHZr0m6VMF
lkO/qHsP0mZmth/3cCD5TeJUTzoMSFskD1cX4OcbZ8eQFHOXaItBbIhhg/rl8CCok3fQ93arSc5h
Y7nfFK0RZ1ylQmNUN55YBTl+V3liY04aepYGrEVdRB3RmsccFFAUMEG8isfItU+xf2xSC1t85JQk
EIWP/GKKnKKqJAteXylEhCEmiYzUOH6QlqooWHrBIWLwlLkG65ycJPpHNfcw/Xj36TkgZcNt1d/g
ajVTLJM+oBdl2+jMjN2R8bmHsHs4IPEIxFFQgVn8iwJMHrugkmiQ26ETbh4uIQaPssQVB/JYAneM
cUIrtMbnIV1Id9kF3VMyI/nJt4sBTw2nFBO4d0Eo6u2/VVN/goGoJBnIxChx3LCE4Ct3bR/qJYyA
+IS6Vrbelrtv8catn9ygOrMM8N8fmbm48YCDe1xopm5lLKR7ZWwwWL1M/CAZ1W3vxk5aRL7MwBD2
7rPd7ExVSGqISSV0pOw9aC8xhmR7yk6KmPFaUNKmpgNvR8TsFmGbs+W4BOu2jl9ZDIE0quC5McUX
yQNvVhjGXHXrSYIcguOhCd81deKS5YsYlw4sDl2M8B2yNrl5sBacI2iyC+FPnJWsInaxB5uEOSlN
jzrOzCPNjzjwVaYMiuMPN+c1SdNBAJdrZ+ukag4SefD2WP4p+C6zdDjZqM2qX4UeSiJAmy6DQwzH
hzHZmQQj7n3GDFu6WZBnhPukfm4dyCqTo0Kfph2mHcwSxaxWmTNX8jhFnJHWw6TVY7IEXe5L6gtp
FyCONkAqUBRbGWHdb8CZSoGFwSsgUCrDDBNMFpYrdMv6xf17vZNk46EzTipQbgxZvyVkwjX2v0Qu
3jW4tHmxt7QbXQTBPJGOueecJuyBPS6E4cI4KCp50oD95vQHlBxtZUyuAHLosVbXPpOOV/n3kMnm
PovTAFP0fXdN4PDT7QijNIDE3uUbmmoF+yKCISOMXaCGqk9l1KWTXOxldMKHCOVMfONCRsx4XaeJ
RzDd4o5ExHPUF6s/31koPbguTPMyjjDQvXNAHdH+gqgRPdnuSp1kujIthOJZWSeZeLApOk3yiE67
90BZl+iyvB6urGVDCgPYnRX5GqqOEOe+D6J8vN1nOdAx0W3OWc3mCCGuacRbXSoHZNvOPfVzsipV
YWDLMr2Irh34KNRGAQKn3RwaWYuhXLAXTFRYkYpNHYZaVSH/sUJYkco+DbSJHxVj0P4e4ydWZvBz
0SriWLZQ4C/IakLOZxJCu/nYdE+utQ1XrQgCaaQgMQ9LQ1wDgs/5XM4sRhb3qZZ5F6VU4KvHUCQ6
uha5cOMJtMPq+j3lJl2rRGpUH8lixlO++YaJxMaQOb/Bh3xojmGaktUnJdTrHeIvsSrppF+acj0Y
UKZmx352vB2359FvyobpPlw0vNhPFeKcK4RsgoV14sjKLFf1TLR7OAgxL7efNtjEeOtBksffQ8kW
xoJhQREJH1iNy2Wmex2POUU9i5OnIGhuLb3pdf/7qrmokdhD32gyRpOH3CBldS1kd1qYNQnqolQV
JNgVuhvWCxd5/F6p3l2Agr+0DLLQWobqem3r9bRNbjUUp3w3LBTgfXb5KRTsS9Bm682SQ0olb6+n
YBBbrS7wPwpXy73ULIL8+f7QhWpFTp3rPql4nQA5TfmE91bKVnXr8/FkAKVvo5a1Wmq/l6lC3JIC
NX+OysLwNYslVejHPVGpDmW27qlbhWmvE6cWlaIUpaMsFux3ePsVg01VVWIBPQilSo0FYjrdmum2
kGa5Mym7S7Hzh4jKgUd2+n0BFeRG/ptHUWFo6iROUh3Yd8u2VIhpJQpjqtOxL7VwHT2zbt4PskN5
qITcGiTjmPNJ6zc/fa+LYlJZGo57fHz9a+mdupXPoYGgQ73twP/hijPNxbIZc16i9D+zPHIktdpo
/3YaC6G/TpAiWkmZ1BuS49rlqPUvwV8bbpCLj/Dzhxjo0ntiSDiZ6uUQm+RbN8cCsK5kyk0/js3P
Njlwm/Goee7Vl9AwieMi3b7yOFmRCc8h27B0OpZz5VTMr431wwiEndzz5/ow5j4KTHx1U0AazcvD
uYV0D6KmmPaStB+2AmulsWrVGxLs5JfuOqtx+Yef6XxtSIYU5JNL21MPU0txTAx7CUnRIGc55xfd
OxaqrIDq+Ju8H1EsRFyynJR4gOyi6pp47XgWHZs0IHRNFS7yAyVZQaMaCGMSGbX59dMztC3KpJ5R
jlJTMWSmb5tSxRHix0o02zmib9S4SRHmAY0PS3Qa1fLyPT/26CGI618ojJOlKJluikgwcizJ4CNF
O+VRK2YT0etaoXok0NBcMbsPwik+jrvSvjzADfqJs3ZXTCfJ+bw0aRR4tSVKQcM1//I+INQgGfht
KxGpOcEh5/pCjGcozY4I1GjRrCuopa1Pt/KxtF6e+LY3vk0aU+IlkpplU2R/KFq3OriOFNUq/j4c
RrYgiNva+QfKMrcw61TzntxgKmS1zTashK1Mkr2jH5yrOWsOJHkTaJ4kbyGY8jz4pgN15PZblF5Y
i3VLin+kpHKfhzP0zd02dUrgQcPjkCP8vRrUvRvwN4gKkWo0SJv3bRWbszhhybLTPCMH2w1wsxgg
dKN/293XQD2Q6ad7YfCqVmZKJtqh9FYHrFZus8J4izBayK5aqiMwypz2IZHxv+PPRmW2HjtYljM3
PY6CHgQDnr6NhDEazm9+S4gzD7AUIzVFypc4Zwd5ZNbJYzb/PyxfF9lZ/Wewp67e4df6jAB90n1s
+i3Gi6Wa/6NOaNKuk9Zn0aWUnmFldwUu2wiLaTU4/1RFmQd+LUcdtSB0nTypGw7bSofLQ5G2Xvh+
0/5xed56f53yV+ukg7+jW6J8ShGwX79qes04yIZphHVWvWaJQnB/aCGaIgaUR6rtfVv1pIAAR63r
1gj9Tf27uiKasin8CPkOGAMlxTEh6BlcwXOQGR4nAN3RSdPxC+PNaVfxWlxiV4xXVB3KKq+R37VT
Di6lQPtc9/w2rDeW+GAQsX2AZjH/ZwQizvoj53T52snmAx+CeBZN/eWN1/tfbrMGKMxu/+pINGb2
30b/RpNfW75KJSRaUDkdHI0eoXrFDrLO6Jq61GuGxwI2uya+bfb4rpWGzddXVDsuz3b0ZU1s9Soy
DeA2hlkWBxCBBcZj3TPi2hf6kzoTGxEPuRQ4wvmogxf6+A8xe2GcATrZiIvmFj0rMzHFMLJlmFAC
ufg3VOBXcCst9z4rdipLClrDwbJRV0xy/iI7lFPD1R8jckQYyi03DD4JibQhcthl1NdsXsc0iUH/
W5EYH8raqBh37k/4nK4+Upenz84/6Xags2/1+o3WVacEGa3vVATsOQImMcpdMNs6ZHITSdmWGErQ
Jf6jXyZNS+F/5ZbAuMe4BwRMAs1DJbenAeE1hgbb+GYi3zqMMtnEan98kH1eiyCG6uYA3mlq8rlL
2S9PZg8vWfDnx8tsO9bFC5A5qrvLPx9Y/xR0RtAQPC+QAQmNasJJwboVl+NzMabc4vTKg/hsrd0V
WTz6Xrih7UZ4QOyQFJO9NImDPdrJc8fPsYxeblYZhBwMMubnTd21exb8Rn+6NXXS14rUJuErYKv2
yjuK+ApnoD51gRlhByTjM3E4Ch1FTYlseGDWM5EbRBgrNknTZZNu7Ai0/R92nd3LZyzkE3Dn5cVV
V/Eu/kKq4El7DhKEU+hi+cUbzs+LZqX/8Ebrz5XmIyiBpP/7LOVCfL/vfWmzVIdA6E1BWwlbhJ5H
PnwHi8sUWEp8KVk8KySGp26DrL138dFhtdelTjSGpy3UrA5cW2PAsCKp/6uzzPdW4HwtD+otAE9s
xIY0gFnihMiiG3rCiSoaMEW7Ju4SsE3gfCBjazwHk1EqVYT18h+yZaTT/X4q0+zEkfDp3zw81YFH
T8WA+t53UM0u4H+FX6ZefcMGDnLc6N/aMf+up9ZUju2u7lGDEV4wkBp3hp/khNmC2YskBJrhfuI4
TE/PoO+58pe41EZx8K2ai6ACTo4mWWpk1X9/HVu/A4mmMjw+YmeLL13uD/sH/hJuBx6qFRKb+77s
ld2fLgyb26V2SzJV4b+LN7r+SryTSaa0CUtaWfPdZMk9oALRuf1AsqN14acr8MEWWLB5IIHnxHIu
EKcUmQ2bwIvjXqEUfNFeR3Jm+gGXk8W/21wU80CCTAQtLNWNcBpCfsFdIqH3dMHdqyVPKOpWmNxG
7Y5ZMlsphbHRwXQjuggvSlNWruHP5P6uSalo8JiD83lytM/jXpZw/K5mW9utStLVO/FizYGsQ5HA
yjYPo0o5mUUgF6CEyeIPycOXEHhfTpgetCNuTlONT6SWXZ3bZUoQi02DY525UETR9jAAKNnx+thD
eKrvDUPjKkzEB/7sx2e21n/d65PD04j0Dxr0EzrD0CEUUetJfT4BWzwJtGGM60MaLifDO1+neeVS
ff+x/g/03UeXRrxi6EkV02iEU89PmnyB8DHz7ahBN55pDf0mgkAgF4CWsX22CqYZPCMA1ToYhIs/
QZGf3CHFkH/CXlgmVHE8sMgUgPfGV8sMdF3avVPcxL+A8JxgM32l+un10RSFBZlouw0knobodh1d
sHtb38hRiARfccoo/jQabFrMrihv9tN0EAssKiSLBPfaspW8sMZ8xMyGJ7b0m/MBiJK9xkZZHaq4
PwwWMWbaOdtwsIy0tDhdKmby0itaQass3GpJWPq9zTwIoQNW6kSlWCpCSLiNfGIJPfYMql3xQRZW
9Vwu5p8lvwZ0YLDbkwqDYh2vwqTwGUI6s1iYMMbK1kEw09005Aor5ZN98/P3D04O/XQUMJG1BJHN
dcAqOxg8RaQE7nN58h4K7sxSFEjHsSh5smmZ9bW6ueEQ4xmnFn4TRKfzOZMQnZByQMQrrpsfh6WK
EgCZDQxWArofnYz9mzgxeU092fU0nN0OPJnnTLXRZsKD9wu9EA0F2Y5gwjvBkLUjlMlKXgYPWvRD
X9PA2lH1dc0qQVxjJSNrGzmiRG2xpByTWGoJw6Rr7dpt6b33P0uZjP10gAcZvh5uurn007n8v7+u
7fJQ5st/cpdlwJjPJSUDEz2xmPg8rcaHsUnE8JAuuohBH0PPXrW2V+T5v1SDGP9UWN1H0CEthofe
tq7ZLMNAR08B233ALuhHub5J87RQqcQm0JWhyZ2btKOoKmQW5h26KU/vm4039Q1KtgirRz1FdYK6
O2F8Qn2h8YVN52eGjo0FagbsT2tXF9oTGy707Rgj1IADWr7qnBaH/4r53YFPSaArMd8oAmh189P5
QPPVOEXH/Ljee25Pq0Zi41Gerivu9+wB3aNxIIJm2fNH+oZ7RwxCl2Bdong1Dvut7GdwzilFAquT
KY1fFvnHb6w4rOHasQQM9r63JEUg4xhn++5B99kCrhGiCnHWBrIfkp0BUCE8N0/xgmvnCgPTzMhd
U/RGlptbAEmjasvdvrs3bIDPn4NO/eN1PCPtHGHC5AFAQBr8J/viKaza3BW+2WuLoe2FLl5pamDz
EEIO164oVwPYgCCGGPcWM5ulPMgmXRaH6DTNjVDQmLb/vYI7j2lJkJwlmGM1wJxDLrwlR0V+2AhZ
r5C+b1xT28SntsZ/93DKzWB6e85XIw3zr8JZFKC3sFSF5m3lbu3adtR+rnMIYc3nFcuUQdDDefw1
zC6kcQqhTUwFdlqVq28VgZqXhkyWwdEPduO3rM7sTFCW+I3toflLWmIxc5nLL3CnAnBjmXl4+iLa
T2hrtDf+VCOoONyjd1yRMMlpxilWdJJvpDTA/jUCuiQf9OQNNcDugH9Mf1QsyowCadHxyA6IgEJ+
nymMedd2eYtxFT6mtZjMip4FgRDthKukvD78NK6SJPBgq3MoTWsf4+HOC3uWpsandnPbxKHzWrEE
GlB8d8BhpHtfk1Op/PHBv3hodORCOmpF5/SDww5WuA3kp2tUCS5NlUXVVtZhyrsl/wNR/OvJeXO0
4hEB6hIXOFT1vt8YJMSpq7sPYr0pAPG1WO9xSlGD2WYo9g3YvlSitRYmXo0kHnvotbcXa5qmXAgO
U3l0u/CeI1NCK53qLZFWdUvyQ+Hhsix4P31pF9PxUUb/gfLbx9EEckkxGTf3R0Ys9Yya9nhDYYPw
9cIgIRH53CNoOjD0GSlvjIXQ0/S+RmZriv0JjmcpTdb0MukxNdDwmB+gwtzvFIZ0CwJfJEgUVJBQ
Qyq/lGAEwOX10XQucoik3NKzwlpIkU35yLwSK4YSv9u0G4SLzLQQ6AhTzglTsriDnmS13U2SEj0M
d7uA40/MxIspyh6KP7JffeGUu8GM46KGdyHNCIxql/TaCAB2CkBLjAaJXEPIxtTvuk/TPz73pfNQ
DNuwKEBk97+5czlgpkoj4jlZdarU0+Ml7I6KiKvrvG0OAW39mjuhJEZlqJgDjEXsaVVVtVxjpUAC
Q3kVvO+abkp4f6aA2t+LO6XHMNnQoIW8LR2tq4yWN4UszcwqoZoU0r8dIFSACQS6c4OHglQ6Vg4T
0knOHLOlU+ZDWEqbS6Q2piFcSU6sat9RZkXBdfR4NK+hl5LCdXf1vvlxmxzUMbrt+Myb7Vm+xW+C
Vl3JfxU2aP7gtl5HNfCWeI/JBtFMe2I4KSaSktqRBPFgEx2qJAEdOS3VlV7vJdv7fK3Y0eR1X1DQ
QnmlwYcZGijH1+j1JnkLSieXqCe15UsenV9PlFe/ygn3JHD/unDrsExyw/PbcIbd9IvLet/Phu6Z
Rmo9PGNwsfiz3VJn8rtAIIUd+q5KQjP6cpkPCk5pcOBRlHg8VHNeCrEdGjIWMRxs9Y6wKaz2WM3z
fERRJQ/4ptSQAO1+lTvJTWJs++cHrA8wm0AXbn7M353yOdG9BmzVM0OfRM9zgUs0AJfCM1rIMoIj
cAjXhePTyyCX81C+hvdnqFFCdPPy3MH/2/MWaHL3qyM1iBp3+DiRGTeX+KEopNn2iGf72rP0PJIj
06tvpmjsh/jOP6BIwzEjg2q3n9azvYbQi059Os2TFAoYqSBADllWYfCvWrli1RAhVJMJURSJ1t9w
MxwKKoG2Essp8bGVEt2hNdzQdb0S9pDjzeexkScGZlQnRi8n+KhvFdpMi+PiA6tg7Rmt4iuK9Koz
BdUwf5zDFTr5IiS4ePHqAzD0EfFbJPo6GvxbHkeO5ksh4xE9EZl/J8jPi0FxCePhzdWliQNFn7ws
ulIiW+tz91xajaUgnfTCHU5FucutMqEMeKN68Ae+CsepBwskEA2OSBwp/Yt0KbUlcle8/qL+Vba+
fA6oXEG1YuXliitXECb+BE6W64Hf1bRuB2cu6EtpQWInAisplTY0XM+8wp3/VRxV2slz6BUQAcEV
BrhLL5hAx2yRqcepIkg6Rvno5Oy0YdFSQardCEzzmnChnNUdvjjkrIjVu8uaUs6lwqgEFZBAdQrk
UIRee238Rbaf9BVclv4G1zS0FMvOhNQXnD2pu485r7JOBzONOf3mYDSSPtpGdjLBM7WUmWFSt2+W
+01ONRPkPNCxcFid76OTX2+TQOPRfZK3qUiCKpT2B4zJ4dcXpZRpi8x7Pgv6LEHHyh1WU3v3tlXb
PFiiQuqWQ3AubWoiTt6YfiYVaGyIjIF6T1+GZQcbGOe2K1yKyaeppnCDMDLswxjXgnUn5ZReqOJZ
jbkE464dNinV0R926/ZNaAKTfm6T/8EdyEcBpIrvD6Gi+rQB0JLstPxbpLliUncI8my7Cyz4O5tY
LG4CN5VU3Zsp1PjT897VFFJm7Jp1w2ATfw2h5yRdB1OLJqJY2MJsG/BSPYMb0Cb6BR46AZnOBxA7
I3SsbtpLCrqAYkBfgcXHh3NQ+QI628vNmB8QS5DMEsnY71lflmigHMSemaxpiFiX8uW+ZNHMJW8x
C83Os6V7479hwZsNkNzuUmrhPkO++GqMeKH1GCnw4v9EUqtO2AjW9ZSb3yAm3fNDWJB17sOsYJce
ScTgYOjAWq+KyE797Us1z1EGSUcbdvOrF6tyom0068AaLT3BpUaw4FZipzOZ1cJKgUaZF3WqNe1k
ZQqApVooMRq/v32f0x4EWcYXZnwqfVl4HZR9OmDkgbkhJWOKU4fk7+9fNFtzybxM4uJxYOVmnw2/
M+v+uMLwHRDWk86vk20FUyIHwSYyFxTJeebFjq0k3F7CdwUskGJ9r/TWuDhJUg1SITZ0Z0Gv1sYq
E+T9QYgPf7Ig9PhgowibYOL8m1DTS4yAX8MrUN5QET9rxejXzPmDaXFN4SNgeS41Bp0Vqzfn/YJM
RcZ5DcpfjqBLemHydA99GmRTPfTq2O7nv6aBAevTwHytu7G8bn2u+TIU1cpo7gnpFwbRVhUEj2Fh
zedWpgoPcs95yY2VFS9/xLWgjp62PoWwy3SXz3LHvTpcQo057+GRVho8Em3Fq5Pse34HJzMOcOAm
xIhV6L9GHvXeXMjS4zqEpf4YYMIgTXfcx0skDFZAYjEvic4dqZbQ8iUcDxHrk3BDIrGZJnNLNOZn
Si6Vkv6IzyQiZwaVgE8TuZV+/F9fev23uGsCen4v6u+4+kEe5I3XIffqVJ655z1efsMVIonxlj6y
PNdFI/bENy1VsWInbSBtpNq48a6LiEUowYTbjX14OnY7Q+XxjCxoliRl2SMITAcBei+aajY82UU7
ziGZ+kAMO0CF3A08Qn9I23s6M+Hr7PmtgKjEuP0evwBm675+HvkoOrCRJ/6x3qK6g0uvDbxsM2n3
7kOGpbqiOXrqEpPT3LQBIkyMa2nHvqr3Nldnu0UcZ4XSmqK4ZB9e9yz98CCs5x8PqddtDsJ6QuLU
//GM8SqHwFLMoZHWPkTLTjJ5OOcYwsguJrdkflsxbAuB+VTOy6Cg5FqVAgdSCPMJy4IMivrrsIoZ
WsJjYquEXqAC/ijy8/JUqG3M0+Sl2Dz+i07xqBpU963Ex/LMjRU+Ww0BRfN7kB7LI02CIaHhvFD0
aLBIc7qXcUkm0Bjozl4utGZ5VJyG98g7Lkx4WFFNXOuIahYLhslEo+Kv2gUoc2d4mRoigXSbbfok
DCf82pt1hjt4c1HJyTelK2ZEZnywzLWeQ9vV436F04B3PAhTRyitR8QC0XlmKkwNIP705+avIF6/
7WBpMEd7kU/fwPq5+HDVJ6od4ojzrKRSiUXee+gJNyZI5ebyr6M58H7/e3NR0UOj3FMstCJcn+jp
57cv907TpMNAuUDv63pzZeDoxZvG8ClOgwz2od+nuT+usDxaOc0HD/qkAf6aVhjHsvqdcuCFcUVu
Rz3kl5BSTZmCU2Quo9uU/I37NZRz+SThAu0PRgm0q9ikSST9qum9gV61ufRXjsP67NHHOE9UgBaz
XhG0Q7O+NTGquJxd7qh+UNEY4T16Y135iYILYqXPLeYoj8KhUhkHuUmG7GVAOfVOLgwfv0Fuj1O3
yhSLGrxX0Gi5W+X7GnXHXR3OWF7s10s88EFADo0XYv32jMgZ2hOo8ZgUHrePELHXF0SzQNUOmEKG
aGYpew6PYmYrROVIQgqY//5bmyOtDrp1T3KEfQ7V+LL03puDhVJcQoVLBC0mO+CJOfYSX8HINVKR
+Zim34zgwI01tuR77Qg39ap2LyvOIgpx+Y0ESSJko1xG8I0K00M+8BjK1PPRGpze6QwLIAsDZ/au
MHM++MVdgqozAE9/o4HckjrJgeWCTvnzeVHrZUAHoYb28YV55abGjcMymThIUd2zfw+bwtbCYN5H
UHcaGQNCLNWXY3ttaGUOcBNRhOCojriW2bZk8RQDHmY9/5LWu61wxTlzsuMyrbJ8SFgF5R59zCZe
qpTeGuq1lRxPTMjoz3ZVU13cNA0+JMzZ0x9aCduJhjitnxcSthOBuKc+dKrwqGQ4K5Y4KL/rjw9u
ZHnq6I2E6X8yNEJtTrLPbZwX+b/OT7wHBFiSB7MYH92vHtjCYfWMV/xuYAOlvIll4A5+IVWfRi2K
P2Z8DeDy8BrpcRIQQkuEt0HcGiwMspMYYcEXEaTvwQZjuXYYkfA5CUz759JQyu1LcCxNvwIStzqU
Y58GWiY5V1Vtq8gFJFLMTkoWeI7LXM6vu5E4NV8BypI540NbP9pwNq1vyB8ashYj8sH5HDU32Q8Z
kWTDfowfbBCiN8CV1v62/mAaQKX+OgzD62nKBwJWu1ydnAyJkP2C14yhdX0Izh6wfxQg8EBm3G53
DFnJxsXwaYXrJ61in9G8fwqVKn712lZmpIf5IjXq4CXMOCIZarpsnh4FyWxP9aCEn6X65CX+YVTM
NoHttFA9BRPA9MxQIRlBhEa1AXc/a3NylUYLtel+q5c6aZ9GTDtEbXz3pDWJcstru/UrwukXjqgm
u2gr6DI9c5k84k8FHhCbDYKHKDGpI7p2LygKwIsnUUMBephfFNqF2sAvqB1T39zryZHqV+a+Q0u+
MEUd5MPfMWAmY8rrvY8dbpY1ASp94I5mXoyYHKRz+/tIiS7D5B/Jq+sKoowUGYdu6duOao2G1xqL
bA86q91tJX137pU0MsVKQtaYP9RMHuMphtJ6J1j8yeYbOmOrC1bJRxX+bwV7cUOd3b1RLqXTb1Vl
36dujk+GEXCTsNrFvHk7gdFwLfKH+60gGqzkg8Qq1j9gr0cTIUFEy0IZ+agjuGNmY1R6rJy5elzM
z5m5DRdE4fgvEVHw7uM35lZs+2B1YyU3p9363+9arC07cVF7L6yqoI5DqHo5KIIst1Dhh0ojH2K9
LWDHEFlbeCPkq1b8NVpTYEhu2oSW/U/hnX1VrUaAJyq3YETqiJJSpqNkTCkvxSOCWKa6Bgmn8yBl
/HyfOXV4rLTCLaE6udJ2OxZYplS5ZH3gl67Jvn2VC44m7yzd87BbvzDxl6dBh4lQpIHkZ/F4W/Cc
q+yN//0huENevph/i3kNJmv757Z4kfvns2+8ClRTydfyHa1IvJA4Oho135JG/94TSV9aViKIGJYi
InoKswLnAd39EXfOg5dk1AHjjCjzquiZndDld+yq9Dkb4juVcem1AMaIgPaYIziuQT9iFFWV1/d3
dfybQLPnqqf8TVV5O086CYX0n572AL+oXbeXXsYivhjmPx16UMikMFnSO2hb49jurKJkxry+LSYh
DpqpqV4i/BVmQa2rn8Wakr/Q5sgP6Ka962iJ3LkWX0vKs7diErWF/+5ikxIMWFvat3Wh28oGrZVj
s+8HuV/8U92fQPhQBQcjhyy1P8f4FD+3jA1QE7yc1XBgiena8MGawqIqxps5p8FjHQxsGp/h1lKH
/uoxd3wi2j+G/EyunK4BOxmm8DPyjXW8A7pTPh6Kjr8OPvq77U1rvmvhM8P0kQ8yN4DlJVq8kxQ/
tjpqI1H2uiSIPy+nKZXdziwyBFOIHRV/f5Lp9KdFckznCPanqnH6vp9DLRbBThiPO2gO2wUGQ6cN
buH0BtixxJX9oTdN1MWyoH2gH4TR8KfTfAt1PFD+5+oPwxp0xHXIBaOIdVxIGg3UkEW/r1d9eRyX
hByYlqS5cp+4f0KPZW+8gWyIkMx33F6B08zbx6N8JDjrJoSUQtBU+erFovYeDzUfb+0DISZm9GFZ
Vq6xbUWv6xBpoVcX0l7ixZ6MMSdSPlUaKVTMzAIt77fCvnns4gQrQFBaZysnjjn1n1j8z3qZIkkF
Q2CwDYoRFuaAFlyXQpEYmReOhjJZzoEHS16ZjGcKPkg3DlMZQ08i2Ou5Gn1ZG4SEUy2ok9jxjq3+
gFN1IYmC4TLSdiV0L/t4NC/GKi3Hum9yF1Ww1Ge6AsWwEe6lR+aRNqoX19V4RjiYooleiPE2w8aL
iAwJ9bGEUD/4zyi86bk3gvkeutZcyXGUg5QHzRLit7+bTyL3g8fyXWsEJ4iLB7qsY2GGEnDugHJ/
t9DhevPe3g+7BxUphe1pI5f0qrwoQN//tx1vpNNZBGlm55BH7Y8Q835HCTi3QfpCdzpIVtlnR+1v
hvVGBmLyVPZSs9t7OFKeZCoeRTN+7rBpG7YAARLeecFnGzDbiTcqCXDWz0P/pKbJv4i6VgkpDt6k
DTyTbcLnXqLXFHoqKY4rrjwhRP3Spms5FKsvAFSmixcZ8KPBQuWUhstkarfLi1Ohd3dBSzE8Qfgl
ZzRyK4OAM44fot6ty+YEw8xGHfFuxbGAH2JxrxXUn3TzikDaAnp/Gd+jYHiLPdmkH+rGKFShKPIF
b7XnzBUkIOPxD/Ns31JPwtjxf6qFhjDrTYMF2/YWfOy738KX7x2zzLuwwtxbeb38iMJswj0630tO
quaUKiEs4aYElC9RR7pCu+A1vL6SEky+Nj53xPSbQ2XKJfmhD2kh6wyfPnbGFJ+CDhjpWCE93mVP
37f3rBz6rKcbKuBWTka24noWmI7haLgdbesNQa4MbFoWfugJ+YJok9w8LNwiY138f2eAZ1Qv40JC
HuJq9n/pG3W7f3i7zvozMuzsWEbhLCablxgmjtvc4UykBru3b9tRalpJU0GJ8qilRxhR+Rx39L/y
Yb9CBkaboW+hMPsaMz0+EEsA5sovkreFWa7IrLYR15faw7m5GwpNJKT+2pZIy+i+4HglwX9Tj4/J
PlkpniKaJ7hS5DVxGoOcWpaC7ssNfmtTZS3tTdXN+Fv1O1Be8SwXbNppqjqxbBpf+2+Hlw9zZPkA
fF0W5rXG5aysyB48dKCRP/koVFaHusXm2m7ydb7FadgFDMKi4qRx/+Q3t3Kw4KyrGeZi88nZqvbl
5D9zjiAOjjfQ0zZAphmzCdpbiJ0aGSdG31tcY1Hbr/nksMPkXKORmdow/Af2YB9G6ZgNnBYM//Gr
NlQir2F6WxYXmETcVMyGP0NTXlAU7cbEx1nxHN8zlkqXtJ+sw+tCUJ6LMkNsEMETQrgaS4u1WkG+
C757k55UnuQlolotWAc4YNBUp6/VzYnJHoTemGkD7Y6rvhlyJP3cq6GciXBHPIJ82PkDOO5i0nea
HQ7BJZnYoDquMvOteD8KHf8wcZA+A8bcrMgKyF7yYpbjejg0evNqZpeHMxy504c9SyM2o+OAY98k
3Q9UBg43/WmwK71D0+Mcabt5GX2bE45yBHZemoYhfyFM9YPIKGQIbnB6HKjislZqlFbElxF0gcEk
7IKGaURe/G+tp28VeL3TJQdLMqmvgU9MedMAtGgBMyiwFbTD5DdCKyyfkRqnper69235v9THMVoW
hgNX6s0BQsGVsMW5zSAHp3+MFO3iAWogBxiRbca0OeZ47xukCdRaGDMOXBmnoTxSmxuODl2zmogd
gD+2wJHLaZ6r3NSWqdVnVdAR41BHG+Irr7bRMQNwGo4uyoNUIf/EcbqpFGHJufaNpNC8rYxHwnjS
SobpkFOXky/UEmXv7MnMmLzoArEVSeiWm+F2RsTYKtSK7aNHVAx6ZihTJtlXHCf58D2Vkr6yqgNq
pkP4u9lcsBC4ZhQcdx2de5WztnpvWO+0dPzTuYCB1JkWeXUbqNPXQm4oXcILZSQxFJQPajai+H6X
t4lVzIugSsCaysLQCV+rId5QcFKNT5Zny+CXtaAJuE0Jbb8cBZ4KDY0EfYaOb/xYUrMyQSK+4GRn
CLDN9fuxdxmqL3n37kI/DKlFqfL2jzHePd7Fd1GVU54jxDJ8DjTpUDaI4jvJNVxkJNw6iwiBtqOV
fhV+Uf30Ouf2OtH+t+tes72XrsjnpIfP/rz6oPgVfKYhHzxKL3bb5KBAvgxadrACYjj6cVaTHeYi
YxrXW0ncm5LmiRCd5FMLjAbOAlexVhT7WdZHUFIWSXXXjR0Onklc58D8fP38IV2+8WcM+OmUOpTx
lgJwyMtq1W5HqQvDKW4R6A08T1YNbKkEE9cnWoEIIm5/5JFmYQdRT9EpmMbq5iao1/C4tnGFp6cH
4hfOQj7VqRhOMx/h6Lqi+MR3EqOIoQj1XQKXcfrCoosgKI/CQIq7owIsh+QsYgw7IJLXtVIYnEWY
GLwUyeVZ0ImZ+SgQzgf4TCiirqmw9igTlIGWRzQaV6yXF5LkC2Zv9HooTTRv2oCk82LDX75w5TD2
IhfeH++3RM+HDH2Xh77h9imsemViFxb7awoo01+H6RPVhNxhWuD4bFZ38uhTslR+Ngb/6cfDptOx
u4rHLprdFJ7Sc2hiYEmLR+Y0rMU7bJg2Q9iXSVdnVGpdaFjJw5bdbJV332d+ZpzUCnURp4nrp4R7
UPXEtrjqyFwgVPLjzpoaoO8slti+iWh7EQpuFIlZ1n0wX8cTuf8Pzjk3grT0oAkEK6uPoDqnZmYb
zjQpDTLFNMKBv16OrWRoLYKF3u5MaBMz9qkkMctUBNN6kJrXmy8RVH/PQJ1Y/QMwpOt4bg+at7zP
0QfCZrqqL+7hoJtFNL541J9O49SW9XMQfq+yA2EolLWPlHnv7rDerSFr8uf8bZ0ssqf7e9YGX4r3
63fCrmIEpcN2Xy72oW/PkLRcLQ3xUEQP3df1AcguyNJeQ7zbwNd+zt1vC261RG+YneeUCcVlt1r3
5kqFRU1NzmoZjsoW5H68HhZoLdQ+8T3pWDnh+a29+dq/hPQh3UP3lFQPXnFVzbOW4EqtSlflrFSJ
Wdh8mfsMK7DhOIENVfrxn69VmcRy15gZgfRjubfE450Uv1UC9S16nRNDtZDOP6cRZ012KqEwS1Oy
Stb6e+GG4BIpG7t7lxik/gVvvZrONJlPYwlT919apMVJNc7k/XHZP1yLA9Lnoq0i9q2U0fAlL636
nWcsLe4PFZHLEFBHqpMt3+RUAldvQaFV43+Ap5WmHBeAcQSNtLeHEQHpMb2UhDOgsO/Hjw4oU6iv
pXn5XSiVnH/blA5DvSeu3yK3n7pI8FPGfciKqDV9NRLl/y2AJfntCfQ1SxrfXejMI6fAnTOifh3Z
oTH5P5yLgswJHdzYbm8T+oRA0WhSFp+nLxZoneZGxZuhfw9VhwgmZKFkG1K194r3zpgQQwJdskW5
OshmwXv6u5vbdZjfdJ2Ylz8lpnjldBlPJzCBIpGOkVoHSXS1Waw7JPYTt2CaeII6zrnqYzrGSKhJ
wK0FV7Lz2kQm8NA3I/BZX8YVymGClMCZgq65CoIWD5yZRRntvTnZ/8Ll1atI6mw+RG12DVKOBTkK
heGRT3XWkKEzoyax93ORBDTFbD0oiqsyzj5SSVF6nGyDYfsBckQx8doVOLe12w2HQgIDDiBRBeeI
m1haBJWxDg18WmgKNyNNtHHTkOPzblP0K7K694d3FDfSj5yTXwObYuHiS0M4t9OJ0aZ/7u2J/x5B
O2rY/q13Z9d9j9r2vRXImu9Gx5DzLUH1omPsT5Cyh11pLJRgMEvLNJZjQRGmpNdpwzUDX5t/fj1b
at2BzAem22+CO3Wu4Ag2rUMwHN8CWIjXHV/y0ppgJs6yhOa03+pqq00VGz+by420nP6Q7qSW5hHC
pAW129lnXKUBfALB69ZF6yvwKYqdsBBMma+S86HS4O/jYA031wI6YOFmWbpqJXGMUW+xbGDCfwqd
xQaAlme+SY/viOHTY5Ncuf6wTorVZonyW7dALDoVb/g6VlDJD8DxqL7OlGhNNGbkD+Fo1PwnT/am
mnWagUHKYs/BQO7Moc3Yy5InJv5fr0TdTBmVhE392kRm7ecVMssrdeC2iKcIdSXTez4fYs7eqvLb
pFIQEGiXuYhUnc3kKjBDFcPW5LdMAHdVw95e0RwI+bi6FLNEDrRiYsSduv9n8efRvTYQJoFE1BWz
8R0cplrx24dWtrbMMlDBPG4im55br7VnoLhqneziQD6aMJ95ebqwFqUJBclShq1uF8y4y/z1s9aX
iXp6UFR5EM1KIOfn1Z0HDngTc5MmZOn8hPAHKNpTQ7RdBG82CezvZW/VQmu1Kwk31ocQKij4+8vS
ywmkZ5Nb6Q9UiUhzEaDKMaid6a0omodLO/Fbh3T3rc7mM/59aRkAYjx0Z0v9TpmZ9ew4k035aDOv
5kk7DfwaGxWIXBBOnE7cUoJVJKPM32S+WySzML3mbgzbjO+kawXbWaDn21raP9NUUP8eEUwdCCgy
W1bj3IssJNSAYuu63pgWLVm5S64mbVn4nGySVz+4IXLRKFP7GAqYQQ/ZRzP8diGb+hR3HO0HNZEb
zXbcQAIRXEFPy4go81yH+qecVF+C07o0vzP3NsHG9GvCIHm8vdtxiC90hj8Jt60IAMut/9fbQtVu
eEqsblUcVtGcinum0EyUmmrozERMYbudZqg+KpL1jfTOLHDrFT8Q7xUUBYs/tW2qjW38NH+ZavvO
VlVS+YuhScXfg974NA4ouVPNoNnnuCjxAtJmc0YILnZ4PXGEr6bx5aNFb8aDb9GbTNGr9lsUmPhQ
HXGtUrO4/7LRlFPwgGa0PNgEB06QJbSkp8sTs54rTiC4mIMfZ+pk9pSCVVwbv6YC8pxxtGsaZtwd
aOIjPVLgxqIhiJlP/xXqMf25S5V5Tcfj2lUA9fJ9mkzSZ9yvQqo1gzg8W7LDwWPZ+K5UX1aN+G7R
MIaqN8Hd/7njHaLZerUshpQhlOr+mIg9BJHRoeRHZJYfoyLhIg4dHniPkwR7AlnfSG0kuep3Wf2L
qSrbTu7Fp9lqehFdpGma/3dSf2ixRoDieuE0YNJmjTDnWH9srBQFu8vHVdArE+odqZ71z/ezsYxJ
T+bZL1a15YgYVvmIV3auJbAFAfWIIdkhBS8aOPItBZhLjpMAqiodv1Tvb1RNt5H8+9lDA+oAzt90
muVVITVWE9yJ0ba/dv3acqc+olpmONFpLFrpKxIlqAhsvHzl2qiITYExrUniNtLlLaFSWgyxdiqG
2hTZ6SrWpJTotTVJXsu1rF39nmfkoZ6mcmTnNOb10GWBq6aHHSS2wb9IKfT+s0fJjoa5FlxqCRu/
OdiPeQACLEHq41aghErTx7dPyWbyZB9WVwQqx+E1M0WnOCF7JRiv0Dirgy0G+kq6n3Sb5EgO/7RX
lkQJZT6MKiuAmvqHW8WOBrUQkQGFueMlI6B0WqyGC8gHHxqgO8oXqReXYOoZ7CtwHJxQMfAqRQu1
xRGPH4t4lK1xS6L89Za272NqNT0rpFknIUzhG2pYmuRqZoK9KKgNOXLGTwBcE4SnX9e1szS4KXJ7
fi85eRj7JwhgWWX+9NXg6fDsRJnwdkxKCBIEXkHscbXJInEh11mMImuh1qtIv1sLn+cXNRDIO40S
YOyuvxABGMdQNsfNiD+jv04VnwUIiwwI3P5S3W2h8VirgsQmPqNdzwaKFvt5nr+ZYdPSIqAjBLgU
AO4fodWpL5u59pK/8k7Drt3Ohr3O5yFZvpRN1mUpqcYLZ99w4adkbByBXHx5SDqjh3NTAUobAEgy
P1qZfEwGc9dGdqb62RFpvs9CoUptOCm/CeWy5MIRsUGE3FlJd4m3L6i4820H1ANL9FIuEflYsnlj
LTS7lWt5jWE06EaHblOP/3UHNXKmwTdQwj4Wag1xoJZ1z1o44SOdyaN2bVTK5+gpXvQ4xKLfeeJo
64PkLdwpdakHpEh2jHPGoxeAZflZpz7d9BGkOQwUVV1T7egm6z+/AC1cXZaYGcBWpVy/ffD6BXQK
HQHwflmXUEU82G7GaI2G6sbcq4Vd65d8hAvp+Jz2ZHGUF+vcZN6pW/tH/Kr6V1IJIRDSAEGZazuy
V4LyQtj2JQjPXBuqifq0XdkwwtBwBm6aTdJH0HxuSQ7uuQX6WezCHD+H0CWgIVjcvjQAO/VHq4rH
1BzhrKMD7QQ4xt1dUpF+aZPkT3JkJwYmZ5eUs0+fIFZzmAvxdU7iP7M+2B9yESegddB0ayLxxkCs
zqeMzqiHABylpd0fQWW2/+MyFKe/C7/YhMYd4Wfa32BzcCMP8ok0mE/MjBNx/BCJ/P9ZzSuRD3YE
9mLzcIsP38IhJtcmPPPKg4N9vrSlUvsl7riN3A/Z1NbBpSt1+gd9KLsQXz0sW/e8ko8vl8oPgOii
1Oij9s7dB8rWLrWnIR1p1nsGOnqLgBRsDPjUkaAH0axb1Og0iKIs8kafLFU4xCEs3UF30/1CPQqi
eW+bsq63xBHxJBvgX5J8hieiUSZeNdwY075mEov6ydfwkOg3U/Mmx25d4Wuj0yTmedj6u0PFpqxG
N7AsZX1+J2mCxJFNJ39e+LZJIgDCpmYAKHY92QdpqZDpkAE+0CkYnGZZq0KFBMfNmTT2ajxooKma
6+hAPOr29N7Bsq4MHGt0EKIIqkmCXcvDIPwPa/NxcG05fHWwsyGAd5OE1DG6c+FHQRAVNUpZzeVT
xHgerdpyjNzAEVAwbdf/+u+LIIJ1ExjI8olM6c3OPR0fkcyZkP3HaTI9LRu7624+SKm4mHVtuOHk
ZyMTAgDIs2iaFi9csI80Xp4c2lzCJJ8SJyrccoa2ElDuFDw4E8tXMt0VGXv4RZDRCJw7d5zR4uWs
VRDPD26lYfGaTceGFxKdEOEx9GjT/SyUEJF0h5ABAISy7voKQZYnzFoA3Ydb1Zg1R7PsR8/zCsby
07WfcvChDqgCJjelpAtR5+3taMZ7gg0lUhDj5Pqj2R5wxoOAIECPuPgCBJKb9BP2d7lAbqbv06TZ
a88DhVj9pYb0thAHmWewKJOz3ZyLnYO8aCTo6ZHHMGdaPaXo46GPMLf1Wms46Om/t9FrmIGXT6DH
uNBReNLcHzyxS/ZsVF+SCzF6xk5g0UY2cvQqA/hD3/EVGSZ6FaIgCQLLFpz0BBQeA+AwWXgPnOsa
P6Ju0vSG9i6RrQsbgUAbwoEfRJTFwTMUbmbwL76ke+1r0wk33TyyAscxFIJRG8hylhrs+Oewx9qj
wkWnX0omsSi5DYULqocdKaM81Zmh2EJ528OPsxLxU4GhS/6dAxB88cVJfuvPCLsu+UhLqKQXbP9D
M5bjepuxPnwAE3jchXma1St/LGxJiRUS5xDlBb3UV0swQCCeLDSTuVrMEoM8cw+bkjVDHBXvkMKx
fTZgz9HNWzEvzrnfylpc80n5cyxLIDHA9eeXPN2GuuVSeu+e9pwnTOiojKAgJfpF4RUYAsj54k2f
ZqO5ZgwCwCqIUMTVtPYsc3LMF8o5+keP2PXitD1Uti1sKHEsxEy7/cvXJPvd3ZuCro8C+CMKHC2B
Uhy3e1NHL/ji3AngjF3lGa0viGU+WkxZ0dlD2hYatDZPPSRq+s7jpP6OacQt/8h4BekeClSfkQuH
EbLCOkDa2QS1vkhBgg0MFpDpqtOrPZVq70RswX0R5+adgzUvKHuU8sn46FbzHFPKQoz1Kzrr2ab2
m5wKBpQyJ2Ht6xwWz8o5jPEH5GYkw0EU54A9839sK95dxVLRnNX/LblTeVQM4XlUM1gc3DOi0GbG
SvIvnjI2Yz+uMnnU29ZBZ6fwqQzUfe0JCTEPJC/dLeivoBlXv5vMhJanaxgbokvvAKpWaqoBaRcI
9FiTPq+IDWlNLMmLLVTnQ++J3qNivqMgyf7zPs14NXh6r8xlJYpJ7wvd/02gJLPxdOaBBqPlRXdk
Ezg7Wqq3dAhdlTuaUKCpQPaLTI28YDN0GbNYkRmBiLEY/3vxONr+gysKjwnbrfeo6QXW0fU0FLAW
Q4ktB4Dn2a5k8JMkOxM5b0jdhjjrPU2V6OSOUBEYqaehERvQzBQ5vTew9uUOWoosmu7kYid0t69n
JpHNKxTiM4RRs8P4jCGS/X/y9fQ4fNP7oi69QQH/Hb3/gPEsdfcLAtSAVlnrRzcXBVsVW5bR3FD3
28wWJG4YIJkwU/wzSq4cLx+88pJzctt5BdwtU1efkY2ehnqXdfbsAu1dUaQkW+CZHa1vV7ll+w60
g3rzfhZf0wDomLVnBb3ZexneUQJmOTcpXKOYR+6Ta5J0C7UpoyF2gwSCrnATr2elZr7qONq10qaS
pA9bhumYVZCdv+9bupFpjRyHeS7IEbDoYOTHz+Aw83Ilj9M72zZtJ/MAM9tA2NNx9VoJJhHoQ71n
nnnmlKbSzYHoQt/+5L4PtDBOZxqy/Vr95BVP36weNdd+8/hwk7ILjDDjgpbVU25A7BR8P5bymMUj
Y1a49GO3NiQi8X1w2IFiij6se5cIj+mKmE+YSSKSVNLZyho7rc5fvz68YTHjNKGsMjuZQC7eeITe
qAT3mae/QIgI0kEbO/KO9k4tpS0TlOL2qGsvAw1vTn6lr3Il2aNVlRutnClGMWznrrdV3ajxtKKD
zs9bly0/MHTVCO8m+7NzB/cANKsdh/iC6PDfJ/xvCR75kPvf4fR3+VYATsoMZl/4fqCUOXH0NoDS
DuAs5orCwTPuuGU8DwXCY8n4uMwJJG5Ehh76yR0jMKSYvIKVaxnFC8iEbVGn67HO7Ijr24SM3T62
filymhq1TaAEFuPXBV69I5URK3yUCcFAqgf0+TTO4shZuRCGU1kDVEwG7yCUExnvoKD8zJRqZN/8
k4HJBIukhtyIJWgxRVGP98Xwlfeb2OhgNRSWSf8WFJM8duJigXUqiVa5fLMGHACC6D0/2xaDqSpF
d3MZ3HVYmU8XAltULEqj2ssAwCQ9ynKabkML5MpeU2ATHEsR5tcQ3QLnlewa7jOTbN0uY6uXbcFS
AVrZA1dAFjAMJtTGcHqMxSbJmy5JHrpGL0xiUjrrB2k67Bd0xevL2iXxVb1mlnTnBM9jsd0FNq8m
vkjMrZwwblIBS9UNr3cIeUX154dSaAzrWm0ajOBypJuV1o8qO3aDIa6iQIjv/nS+RSd8epgKm3UY
CMt9E5iLGw7vWaBfQuuSytJB47vmbmRlzBVKvo78kb69n5hgo0jGUCo0WOcktR3hQ8eCWCJnq5+e
hfG4Gcg3wPqer1x9VxzSquo2qLTMzLyuATcd0Ix62Im716SXF/Rr46s1c3jHDJ8jMXUwM93yvQ+c
bVysLA6x5BYjZ6yDKHrnJ0NLUubHjIa2Ar+SsOd6f/puvM6hG4oa6O4tDlbPMbFQfvTvENpCFoXb
S9wKLnUkb/d6rU5jJ5rRHNarXVaYiQ0n3b6NLNkwEC0SkAjD5x+Avbdt5YBd5iTpINNijGwTwxQc
V9SbkI7sdcxmFdo3NazmCkD2IZzUHByn6n6EFsz6MzmTnS3cNNQQ6KxaxgPWfwfEMl/tCx1omPLX
AP2w0DMRCuolG31z4Utya4aH+w+YiQDazb+D8M0TSRjw0STS5zYjUbDkf+5wzxHiHtiFj5DG5Og0
X9/p1HqfFPQkTcOHICC1lvZq51KRBUlTnxpqObzpQeR9/Y64MMXZ9uRGRgaAiPoW8ds/GXE7qgSv
POPjel5gxX64CSe2T9EfQt4FZnT9Mdgerqf51MdddLd3JYCQKtyLml5U1iu9NhNgdXd01fQS3Wwy
WFN6nM4GiIqmzJoPidmDRFIMxKkW3ZhjTKcvarlAgqPmtqdjurM1mbT75qrFSXQYVT+kbU4x8wC6
pzGxghYbcIq3He3hgObOrrCih+G/YYJeknGIZBDR/myrRmqZH7ANQAJtYQgU7M4V7vOGQCp5UDwM
XI9GxssNuO0z9bGjAxB9RNGpVRoAbHL3QRlx2rY5q18kNWI2agrRVxG7MY3wvsjnae1XmpwAGXYF
o8LAnWAwtGPNJThDLmQ1mlkPmcIvpU1blHim/ts0ICcXVaicEoL+ajkbMtmpmbumFjRB/XzNwDIv
Iyk3JRX3svryOvSYsw2D+45+6qofFqt3RPkM0SfVY6hF2Gd3Yko8jmDUErejIYNDppY1QzumlNsG
tdcPj5K/JGFYmLziEWYjzFKuX0Qj2kC8+or+Bsr14I8YXgtV7jmeizLqyxSmETv6KJVpN+MJUML2
cUqvznLF4Ijx0gD2t/1sE3HGbR64cFKy0Tq/4RAhn2A+9PuK73SdW0+7xYGnefdjeZLDgYC5PUPk
mQN7+C1XIVcS7oFTSB3vsC2IRDqX7cKzA0j1i5doPnXm4+SlKtP1Cag0I+Je7H9xWr9kJv58vyfd
r6I2iDXiCzPQJxKOD9cIRJ7VVR59qOAjN/wqVxrRPGx3OPgyd1lTUhlrZIkImTbYBH+0qPMCfrQa
5i9AzCAUTd+uyo0YmYnTq4DuImmvZ62Y5fKR4k8J8Ya9UWurpppAJHT0UOUDcqcTX2OB/6WCJVAI
kEb4d+fj/NEMf0f5O38V76sBLtSmADG/JqvbL9R2X/39gM/caQEel7aPS+aVAvQV6a7vcA3dNXXp
vY8JFbo5U6cDGOiKJEsMhnk7EE7/U0qmXWvWOVWxPoBCUEcp7HrPjjYq+lKX0B6wZGj8akFDdAZp
fPPYOfNFvWBrJqp2ngIAz2WcZ5SecSUR4Cbi2liWz2dp31NTIuUIFamhm3Ql+vkRXGx02fG+QYOE
B8+zQ233sWubZQha5RdtWJTV/DIRPx0QZN9878veLYeS5cugAxSMOYe1wJTsVhqhLLscWBlPsnMS
Wws0m8wqB8zfi5Xr3vLTeUIZApgR57R7A2FQ/eZCoCPJZNNMcBOg0sxLN1P+1lGbBG7ZMKn1KQgR
YDMuqsy860zNL5495tujYa8MF+QfyYUdUZc274GZrqDEKOUTiWN5y9FCjeRnDCeXHhM3Eo8nSowe
boQjrqIayhv08i5ZvVpaeLFc/EtVg/5MINhAPqaCPWI8UFYpdCGhl6uVIvMUsEudxb4OvzdQiUEt
UpUq2By3SydH8DIQ4FksN/wO9DFH7hZuozn9K9oY0ms1K6zwh/5qR1rPePsjhGbYhoaHNsV/HabC
VOd5aSMumvcrfw0ZNs1KAgMM2h/C1UUaE+97uHNiSa2rIjmUf5D28dv7YgqvgUiBUi5r99RlE4vv
Wbr7lmSlA7TzzNA0BRllGrT10PFk57BGd7VYYtuw0jMx9VY57HLsFHQVF34PjjgRgR2zidL0DYta
DzSzPIx+Np9zUim3bYakB1d32b69GqWiZR+kItduqzMhplwNHLD3n5hZzK4c8rRuNt5G3zXPkBbs
avMHsfl9xfuSqrk8W87uCjTApQbCSVOUwW371JJlmjbb2P6XV/fSXKxVgQ2mLb8l069trJEfHZQX
ZvW7B4Y+mX4NpJTxCHklq+9lUJU/DoxwweeZqlNLwAH+U6fVjwSx/f7cKc0HUw2UZzYybeTU0eA2
hQWgzcvCPPxjyFREQCD9rHFFdedP+uT9MVRuz5aTTO9/n2tCu9mtLJN9FphZHpshJH1QoG+Oz8aX
a3Bp8Hnhvy0tR2UXdpX48eA42Ou4TO+jQPXSr/2/EuRM5IUr0XwKmCpF1qhqOEJuD8wn0XaKwUJD
qhaZFcdAuRobrfJYsYSyCvQiqljxucwsuFUAIZgemC60z+WhTSZx2wy9cnkBLdP2smKebiktogqt
gnp4pBc3Laz9/zGXGVbJg2Bt/xAaTmNCdu7jUdMszwsJX/sVKGUtOFB8IHYuYYiMoTQXOK3jU2+G
ygLi9W7peGnAm8zQHStJJq4hzIoiGqThwzWxST6MJpy1+v7w9KZfS1WedDYPZByekwqWU0LaOa/7
oRSg6BjlOiyBeMq/USLGiEmRUpeYF5S3Z1tAX5bHNSm2Ijzy3S7gK9cEyI5dSbzWjV/1TH+6L4cT
vyTnABTBG5Wy5tvFVWbAvvdLcd+c9ccR2INDxTOubasIl41YcMdMFKz89tjy6yWIKMPVgeuvyoiI
Skn2OHxnlmUw7yCRVrvWLT5Ffs09RgUrq+aSoJtxP03lOYjOnWNVigia0u9R2q71gg1rs1v1aMd6
2yzga9WCx0WBJ+4/shLpozwRlTZv+8rSQy1aZv/jLHcIc6js2p0v7544TTCksGppAPEaolOLvixW
Ii1fMSHFI9UqVU0pjFyhrQfqqOn8HvB6UrTEgav/oAaidS56R20Kz1jS1ZLp+AGValYRVHTvM7wF
Lk4bHMDGnhpkN8eRFxCgYaUcD/T7SNT1r8VC4dLQxgF+3MnSvXIqcWzZ8TX15Ge3nrokp6FzXMOV
uXdFEw003oErx3ta9e/kH9CI/6KlroyVIXPLsU8aUajey/uKTzaQcF5xuOnRfOtEdZm6wa7dq6CR
94CjGegH8eBz2LWR7BkvMk+oQLIUsTnbugfO0l3Z3L+l6YusgYNyxt0l3/LPhykTKoM7FmA+/6eT
b1O2CGDLc0ZarfVpkK1HpIxxkIxe8d9IGTe2QGcOG7nnyiHa7UNjxk3TYLROfmY/fBy/BcpRmGpP
8sePShxo7UNtfDlLYxE9RwoM/hFSG0cA1K/ujvxEpo8dpeI7Y0zajvleoSbD74DC+Ce3kg6cI0jI
gGIAu5Zcn1f7vJh/2gxv3oXV5iacZdXdtt1wFcX6IJ/JALXs4VcgGQk/RlhW6cy9iizAXrYbwx6H
lDN2LsPWzmrl553YgLAR26k7Bq6SKfhPbjr3+FObKezpEtfEYXwMd/Caz9Txleql2Cm/T2cyFApN
hznKGslDaVeUM1QFy2qyifRPPC2vKV4jvVIbXWbWMH9Hkbp1+dmYUYIB+6tDwzlx+HhyLjdzuKOT
5xTbSqPVd0MNcBCEbKmE4MWAvX2wS71pqpsz+5R/D4iVcYZNm1UdUS1iqygibHz4ahHc5YstROq4
R8GYrAK2pkFpwox+fF8dvRkteGw2nGhXbcZQhv4U3mbMGvEZgc1rSNIAkKRmsmpI+LI+gHi6Xqom
QkMjlh38ESwtdPf6cues8CDIuW/Oc24Z3sGRQ7NKRD8dxxjXtACshy+4CSBLAghr/f9tChCVeb8s
icoDpWDNDuerbvJJzhXCqjV2yGmPzG+RD//rl96j1KqqvMBhbvxxB/GlScrn6wLoYNAHKxoOxDiG
tb5IryEEKYP3sN01At8q5MVmhTvjwJLlg+qGSr0D480OzgpCYiYZXacsUSerxL5eMJNDJT2zORlk
Sf75Sy0OiBTitooILZI4m4Ej5TkUoPS2EmgpviKMpc6ZosLhojsrgwGwrnrMJU8pBw3JLpgftioC
EWkBplRxb7vq11yfpredotEdvO+Ex5UukHo7IaAHTqo0yxOwYfPTRouxySJFB6Z1GZl7a06lKU8T
HaouGU6XsNMg6GSY8ESG0lCJ0iZ6EurtNLRrRteuM7UwWWRBp1PWwxnBr3Ej/2Wzb57lMWkkefY7
hpYMxu2GZ2BG/JlX3G71llbgvsTTUNPt3bkYHRHTOsCBhX018MAmt5BvsnCP2jyeYEsKeGA2yPUq
vVbKKXk0Ujwp0Ax4+DfCon43iZtUok4PDu8U2X0sehDx3AeHiM1PUH8L9Vg6QQV9GNfNH6WrfilK
9lZpOmPZXOso4Y7p/fTJoaoqf/ucqPlE3a96ZS1lAroaL8/EUf20zi4avOUigPB5TIzTKjKg+Eea
WwqpmA9bmDtFuEHtCtqnMo1ULDjo2vUqjYqTMCUMpsXiVx2n5/eevc6WDeqjFi7vCTKtFVtBnxOR
EIAE9Jr6K2GgI9L5L4WIGFix7LC1FZVaHgpwa64VlG4hWjE8xeMLcuoayrqT6Vj0mudD5SUWmFUm
Mo7kLqx96KZMvvT4nfo98+//tnf31AsK2cLN9FhsvkGb2LwAIGSMPMMEDjH8CXNumDXzzXSrtCDe
kAk7tbTjRyerd/zGPUWBWNKdfyVMGWCoTZrK+tOqg2BxgiLfUYZ2pyJCzSRi6cOgKnr//oIo1h95
oskgBdS+ZNqjgCbmzwJGPaneolL5+G4R0vZwh4rkVnzcf6hB05e3NftDMvCOV6MtJJwBN0e/HuPc
/5yKsgid0nM0S8hgm6R4RKcV2vHcSJg+m/7SU8bYttmcux8VV21dLy/PEHShtVPV+iymwJpvrCiU
lxRkn++acvLeWOxkipkipsNB+Jd2NNiTwswnOk562PZwzQ7ZjMfSgRkWXUE5GXRKrO6ISlvAjYWL
2/2plXuPYGdF7mhCCcDOKBj9i9ITjGXN1d4qbE1xGsgMvnx3BxEkNhWfRBtIpExqQ4BVUZEi3LzR
mdgB3fDTXFtu+JVazV3ULYNGD9tBJfJMpLjbPOXLSwcAA6J6BAI+KSz4MWB4I9Y7Rhlxe6OtKdSl
AYC6wfLeVCP9ixQQQ9Zy4Z3ShoD1rIqpJWNX52tvWBnK6nOlpxMnNvnGC+mgQ8DNWNilEXHeLnQ/
whhNtRR12SxMeHHyOVsW1ONjJVWZ354dPVQsSFRxjOHW59r1dcu6vlyev4wu1MSEoKeLuchxYjBp
LJ84xBGYGJ9ITlrgDDbwx5YJhd3jJ7lzmGrIicZQ4jGsrQ8kDMIOydu3wK62vfj5Dj5ceZQpvL0G
Ws55oehwTj7ekD1Y9XwxKwduXc4/wKf7GEsJcsKBgrilTV1jQr5+qbMlvcsxPNhA2bR2XmGPcWwT
CvSo+CI2a5gojP8Lu6uORQsnQfEHMdYfRBUrtL8hATi4MM1hIvhiEj1a4Fjb4lmVxWtiooTznfxJ
vz4A38R++QiF3nIpzZVilv77QcyMgPlOdE96oTqQ/qjstbkg7sb6jB0AcS+Zm9LxM+v+bViIb9lP
YggNtVxMezTIQPkKiYjK9v2XAIQXlKsSazpTXeauDv7cMMrET5SA34hDHzsXaM1uxPFxU80zrS1f
U5voWKZLxZQdwfUGqETMn/F3hlga72quo6ttuOEJOo1BV5465LJcDP7H4ZpdxSPnZGI6+pJPAXAt
BMdaw5CIO+762vThjxbcOKok570BGcBhuQaBnkWzgVsbiVnnOcKyVm/oy9NR9k26iueYFzNC/zEq
KACFiF342LnPWpwxMjWSK212wVcIHErS9nR2peIgmTjVXJY0xXyKkvdposniVTModuWAGZp1Zk7i
zll/OSmCbWk9q07Bm8L9GwI5lBll1S41m1kdDruXEsHv1sNpP8zx6QiUSUQMX4/HE06dtbj/n2ER
MsjwvMUehsE3tTZmkUBnBQqCC8ChO25skQu60Sswy0/aCtz989seHXAhtvZFlvQufW6N2JT/4VGu
EL5b9dnqxCbSvDYCiOBcQgP4Kgwb6VaMSy48CbhpUpKq/bhrnVkGBBOwQxwK8ly8KklpPK6IofYm
gh8gFKvW28SPptjD6d4s0iUO3BBTEOk41FUPTB60GoeNWB+JR8N9D1LgT5K4wuSVNiPe8au3SgJB
EL9C9mxgqFiGsjPKproszXeBNIsjDRHMGgwA7S0E9c7NV7oVGwaqHnpFFDqgVYVO6ezd3tVOLsx+
TCYjEhaFWUaTL9qAS+H1LD7ZyAgOeiyoeuVG7Sji63LxrVqpRohC2knPDDbKc5pVXW6atMHuoZyA
jtLTnNqnM2Z2Wp0DzQmS8hZzfBN6O1oscuzo0a338rAGYpGbGhblnxEUHKkKw7pGhwpIamHyDYSS
aLHNOD27YYxeptl7TzB+K2Qa+HtfdDwt22HJO1xOv4O4dSsWW9RZEMVXLcsyAN3pdD1WsWBRjDbA
ayrk3mqIlyzhHb5/SgszjtjB1Zf63GuYh/ubB+RQTZKWz0VrKq+Jsl2muzyswrazMHIGE8jqulnq
2UbjY2CkQMBf2tZZOCtsGFR04RcDg2uT0tMiYsPe4GKpuQtPRG5NvwwP7qUIK8g1AZ6tXN6fs4EK
BF2rAofuEKxXfYojFEtPE2WRQI9ytOyUdAoNQOf2w7OfNHyGBIOnGu3mE5bdOW6dD/lap0NclXD+
cfeE1N7k4mluANntIy4lwBMJih70UdZlBrGIaqQF02eCSlJyFiBRKJUms4cpl/MlCRdONv7wpbrm
1PWNPjNxVP/vY01guDjWCUOk25fK+olJt7teXMSH9t3ysMygJYzOHQM3cQvzKK4qop4+mzht3iJM
h9G5iQ3PFdbfBgoPkXipiHWX6MgZx1C4qcdB6txHI2jkVJDEfzHc2zKpBcVc9FZU7aI4oIDt+eGq
AzuDUC9OLIdoJOmRfswHz2PtKw5nusGH/uCBNLgCnhFoNXqmp7nmg/l9wB/1EC7Uua4TeduT0ENY
Dm1kzL/o8ia3kyEVCiiivu7XA69KiXSaUWzU9D+wlX1Lq17gWO2R/5EnTdKHF5KNk12v7+jHVwxc
HO3BnP7n2T8Vm6aanpX5jHqKOicZR0LYiI5mzhWG87Yjevh6LGuGSjgOm26EJTOCeA8QqN++qYmJ
GcE93XXXdZTXf40BfFlChzsanJ1lZdgjBRTl3EaRe6AOC4DjM5gd17lr6ryLXSxZ+CBB8pOZF/CL
S2V6XDSY+wPVcJ30H+X3voW6/At6Ke42GWuWpzaf5lOJla8QHTgLr8HjxN9uzfEUv0lB6siI0o4Y
9bfoe5uj2BcZ9Uskb5ZC04afVLEZZqHf1XXIzI0jsY0PIXGs8aJsPLHRe+Oed7LJceVsTe2fjeOO
ib1gsOj/BnfLXgcmVeFJR7L+QDKftdF7dNjMQOydHDLKb/HYs7Exhc0Ii7Z+JsA9zkX1UHR/PpM/
86x9YsrArMCzt63bZ6qJmmubUfV/NyJMpVf70BTLU3uaKlwGyZtmPP4K8JT2uoGu8hqQjbB5MtOQ
1AWt3avxfUe5ClXhETeHqvzaRk6r49MdkYCQR9C0G+yE7NS0ay7eib43TPaoLdJHJ8RFowjJnk32
Ux86Nc5k3w4RHqFYDOv61aNeYbh6rG9Hlo+jYqLZUM2pXzNxK7U7m4vNwhXmwg4iOgjNyqPMqgMI
TDvyo4kxIUiwbnlLweQn3145dFG7bJ/VL4Hw44WeTtoJKG2IJEaDQXA5FTV1bG0VliqwE3yqf7Ju
DkbcYNLWeIRTPFRB6dmPB/ObwwZSSzOwwL05fsTO1b7d/Q78mqfbQE6seM03fCE4xkhrtSD8YJdt
2hdWPabrtv4DQyS7K+avA6kGOLjDHBzzpm9Ftx67PkllfKSguwllpR0QIjv/qd+8tTz+cLR6LPDq
z2hfo5sG7pousGhaxqwgRlgD2v5il+NTmN9QVrbVlaEtD+5BPc/3n+fVQbMjws3n2OpJ7pbiMUa/
0LQtRqIWihJ6JRI7vdo2Yn3q9DhORyhpltl8HCPhNYCpSpfRpX+BUEnn0c2imxy833RwZRL77rID
7fOQTUsXbsd7x2tejmsa6yV2A8GNoduylnpNeyirKskLJiPIF7eEYfB85g/Us1l43iv20CxDGqbY
iomF5EhjxbFDRGdu7kinjkm6O7f5T5f7pa47WtKeouWA2J6boUmnEt+pKKz4to+FN4HXEK7pXtxs
j1WOBQcN0RSndZHLdrDKtoanFHuplaj15d8NWTmoup0mW8isea0tt8A/nrkXAfIA0VxWGO1DCQgF
noKqcvCgNEUc/0HY/C3AAADvkmgdwDLEtEHSQBkzipyAL4j1Ab7euixotifELtxrY8K8kj2eMb6f
A7cXYWbcvhwwJle4jOcluEnkupAzt55dUEsJCjiaG0Ek9fTc85ENPJeefHPzKlCDNlYha0WRGep8
9EhHUerdiVcvVC6+sLwJp0nsKUw+iXAO8fI6ksjbVgCmPccPtD+Z1yd3iumpSwxQ6+s+hIgMq0F9
wXe5dqFIkek6Sfpt5cpW4bxf3Uw0rDWcuVFOEivk3sig7KOXRezJ8XQcAhWPeWFjo1amoV3jAPdM
jk86zejmsWIZ6O9Z3Ddur3UJpTAMUsiUzInCnxTbL4T5VsWX0qRu2cWLBjU2IGrEElqA37RiVBtE
U/xTp1dL9rfv8uoZ69n3/qmzQTPhVcxIbUAkitg0X6ZxhipAnQMyCYe1w2OLuHeTLq1YvNFOdUUy
LN75FWrecVioz0mvLoti5FhYr3IdMm0a47PQ6J1p/wDVfjERXVC0bqZNdgHAbMC8nGePzh6i4pOX
RoQl6AZH067avBPxdaFrlpoKR5jrN9l3lFz/GiVZMrWdP8xJUYVarbqdBqqSYnq4yA5RJ0uA80fm
LevJ6m+EQhszA1YyNbd9RsG2MOEKVVLZS+ux++ZAegt+BXbwlDgoVyfDOPeB84wLnyE/ZV+UyHHW
EBh7w7XAMOOusiV5cK5qNtmYVwDrSAWybO9TLe2af94zoafoLJJfnV0ff7bkjWhUNGWhY3OjrvBB
QKBUnUc5fwoGVymG0QLH+G3u7C5ewLcmbilNgMBeohteiDvsIMtvgEjfIYLMxWr2HrZukbdJopkJ
XElBo+qlHBqrmljIOq17UPYvKXo/l+0eyEVMcSOC9CkHle+59Kvig1vDUBXJHHFEHorzuSThbj95
fIa0uAEbExbUkky65xEC4am1PI3XBMiDb1u0BLgM0+OPYvO7xYXgn9uW++WmTkTQtFwCT6+kg5YY
+mWPMyhit+LBuzE64OYma7aPC2iv12flz5kdqhP4vQvuhZ9Uax+V1O4eT8nEk/o24Z30ZHX+8WyC
qZR34vMmvqQknxG2Pt1z4D2++bZF44hSExehmiXmTfMDVPWgwmPwSnZTGGZyAiCc1JJ3X/HsdZsE
mlHKdfpvO0TlNDZvOyeVrHPQUnB09cIeaarnGVu0oKWyGOqxRC+5s2VkiB28jK13RQ171SYwwf0L
UVvF5sKXsZeM3QP+MHRdEAc+CET9QOpltvSft+GxbkR1wUV8In6OAu9QIJmoJvoom/aL/iyrYN1q
WZSSAKo2z5fvbeT2gfbBOcURUh8ubp0Y3DVUgTNsbGwmupqm+cSSTUcJ4m4J9HQKMm/H+9j13ir6
NXKgb7g7sBj4V1+J/xAd5OocNs5S6pWqyOUpWONPW4F+rW2lYS/u4e0h/PFU2imXqGqnXLeVc4ZX
BfELwi+zr15Fmw5jLFnBPTHvBZBgHPtiftYk2fZQXKRmpp9XwYjRYGQEdG9AlhY+F5im2rQ6QH46
l5gQOe806UNbgkyH/PrgQCSO3q3HpUxomTwIxBEhtDzBkGJ6ReLZp4U6dTKTIbcatGzZHHhOGo7j
8uGgC8CvokTComC687Q1YNsIG8/nVygPSNimTTROYlKd8is3TvaHeDbJQirW/skZsOu4aULoyd+Z
Rpi6vK14PRIosiqn6AIXZSM9i42UdFx8XFt+hlzqyiyTTCSa0sAsz4PfE1a0I+jRcFTdugqTihO4
fxBZ2zRClcIqO4wPoZVl1EOW2xreRsVKwDcATtR7rEu5+q+Hmvk+NelhTVbejjm7Nagvj5aLqfDj
198yRA5YJXKKfQuqeUUyjWBJuLjGasFVLaaFMeebltJFjJ7L7fQ21BpOHYU3eb5CxawJaQtHfler
dh3NpuK20gUha8w6tKI0howzlcRF/IMafbdwhTf0x+jKxK4lLR+7vzT5vVH+xCCitUAwLM91zX+3
Rdv4q2iH6aGknilo9Nh1XW5BJxFh30EiOSDevwneBs/dZUsKIxYN/UqsLIAZT9IrXgM0cDyU/KdO
3nxbICD/OP/AjgaAmsqiVwImvDwndnwmcVYYRQ9NA73eenh8Ao7qVQ0Pkxxl+5ZGDXKBllaUU58u
zKBzL2F+NNlPdGOVpSZc2vXhpfZBTLXXb33XWP7BhoQ9B7GnReMwe41JLp5E+sYW+r79xYm8qDIW
mTM6Mkvz8sW5il4GFXkj6psB2ibSefyPGSGzPhma4RtP94DqzFghD0bhXh6kbKB6CkkNtzi7FW+m
EY27Y1CZjch7rRVR6MO9mP8oS0V5ltweiiBXuxBknyG2FnS/jZtnt3Ok/go=
`protect end_protected
