--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
GlUAkJttLHLROZ0b/fJ1ygjQAdeiSz5u4Gkb7uirCexj60dadY/eJeSx8QGGx9r4ssEAZiH0TJEQ
LAkK7F3IS8e/9PlbQGteZS8OYKvbVIbGyMrarVJ8CH22xO3hgeQK8wptpaocK/SvyuV4CrWPof9A
aO/khdzjrpX8am8h3A1Yd68nrvHKBDIz8u7FAtFiUxqxDpgUdvX2SaRQ9HyUAs+QKZnxx1v3rNZ/
xmixQC80NWM7+JsPO802yEHlUvRh8pMuafNPakIaFAlQqpAXeMOQGZGkUA7CdT67sRaUmMl3vIPc
fJuXRmfTaZm58exHXIUmD346LArlJyV69oxUyw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Oj8q2RnzpJCcGPdqiXkVdwEbN4gduG1qWeCS2D4m90s="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
sABPto/O2NFWBuRSmvBp3JMa0rRZbapYsh73Mx+hK3t34YeSDQCFUCWcSJNXVtSw4CUYIWpPAyMW
kvF+eAkaIukSWh2Mbx1ydzosDQnNG4Cfyv0cR/HBw00JTrFnTIxS2F8NKtZLQfJqXEqSE7Os/c5K
qCZhfd7Gp9h6E/vU34p03hsEWhXmlfxN62NSIxE9ZPsG5U8SWccxmV0cKn+pxstYLVODwkIEZsxN
qnw/l8Eb1DDfvBMPrB1Vy4sJgsi402iw7H0DfrfLrwdbvvRFxYiUAsnexIcu/HjMqaaSaUtTKVrA
g75gaq1hLwH2YfSQcqjedPznuyCB0/EVvOa/gA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="imZx1Y91N9n6FeiQ212UV0F9rQsyki/mvqkVqcitARQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3888)
`protect data_block
Mdi6o4qSe5+mrD5FnCvqdNZ3xLGHKrTd5LdHq1r8E0ZLDkSD9LiUq8MjP5Q+a1WfZGCE0pgewcE0
bomHT7MMP/Wy0OBZh0aC0k1s03d1qwJJqlU8YykMifslbFIqMEdxkSfROQ+Vo98Kj9NxM2utckyR
v7TmDtL4lhmgxP0EubBkfVq1PM2gr20Ydv0eXwvywFYDAFH3RJACmIXKAIeod1ClKnh7s2dqO5Tc
cXQVm8OLupiNDVHk/FYoTEOgVPDN1cR0CsZ8VpZpg7/xA6ZsjgA+u6SSIDJiQFdEPbBn+5PoLS+R
8tYWrvo7Okc7N9rRZ094bayHtEeL/HSSLN2J0CNHiouO0a68vfmKgf6ggb9kTPR/BQ10XLJn+eRa
XQOqS5Lj2u3W5qc/Nr2U62GqQmwscB0XQFPa3rJPFqSKb92zXIVKACja+yKsecfjk/ZqKvBG5AvH
Jc8fA8KzPXe/BJTQYWq+L9budznfEC92We3Mhl2D9I3fm+6V8HzfGhtVFEYkWfQ2aVTIp6JYD0zM
ZBFyEKXGxa6CJta8wJv88+iZYCzqflTYjfFMH6lAGeR763w9As1TNuBVu+8XoXrR37tUARdbuMa0
LpEpfAcbYpw5HGoI7Jwbz0S386KSI0sSK0+IZPHy1HZFOYD6CtKX63vgUlH0TYDZL5BJPsUX2dT3
qMfxGdD8RwQMJ8flpAZsBudv5tGfvOFKwqUaNx1VQ54Kc/cet+MIJiXlUN46gMh11eFa6ApyCVcC
3ExGARjc04ykzXI/OR7/YaKiqiGIubtVCNwEnCrRqt/2AwwafX4LfXzombfRVEiQhx/iiDGkL3F+
hN+n6/qsRZ9pIloFO8pSj8ZKklVpOO/sr/KxoTSCF/wdZEGCYHorqr99Ml06rDz/BiUpHmx6eVwC
ma0oqFu7m08X3TDjlHFQTTcI0jEHFV3C3D94AGG9oNUbSdiWx/rMLxElb8NTWgQpamUHLFzCPO+S
ZqM1WTMhqt7vsjwgkYIg1aOJqXJpq0mSELs/Wllf3ABEgeCFx4NBIuzFWLmefOzb5WNpsI7jthnf
ERUB3EJSkf9BGzahTaK+krCpu8ItpU6i2+RcZbuYALAQ56NZdNpM01Vp0UYHNaGPMqCTIG8Q1x0D
Kc0nWycFHmjl1mDe3s/kNSjbBdCJSXWfgx52CDcS1Ykav8S/lrTOLflqXi9KVCDJye2E+394ldY9
CiZg4tEOq6S86h9aBvgac/rG1xfCr0yK0mtRFUukFPZ0Z/Usrmn7b9A1wWS5VJE6G1f2sE3DLqSV
dWYC6JlX/hokWt5/LhUrRw5Z5w+99Uebh9eb1zfQC2P+L1iPgOvewcgIR87ZXHgDjQFX/GTxiB+O
QM0jW+Wsb4q6d7yZiIvlRk/8IGmDEmK6KSeahqSenaDQD9Y1xg3/gVsI70OgurBoPZ/KWdpza6K2
gxClJ8t7RwiDIRYOzY5PsnDA9ArtC3TCpdKSc38wvaP6qB4ffpfg6fE6i/XuQq6l/zXoLP37Br4c
0X0+zqmsGy4RLZiGrJpNc0H9RahLj3sc/aJh4IHNho3Z1zLXX0MX/HfUnA6dQAa1sohpg/L7MUKw
ZMzQZtZPzO483M5dFiNVxYQRWRSqLNNj1pvr3oqBPivmvM29Gh7oCtg4Og2f98KDliw2u/LhcB/w
7NV2rvhibxu3/apBxisyDOHHzpTwhiG6SCmiutxcvFM3dIYji8Fpx66kWnwVtyI4rQc1rHBEUI4c
+3A66dPXp49OBpmJ/cdVUGV9KfUQ/GqFoSfRtTDNLg468KPHOE7KX97ucDqoJid27XZ8IqNFNbH+
oPj0ygDe8GRJhj1GBPuplMig03q32DNPDtDuSeHXpPJLAp/kYtRU845xNoVsxK0rPjSUAMcXckN6
6PsRVS45PN7dEDVw3BkBgnf7BlmlvS/uROYLlzxdYip2Xcz4mkNolq6Gp4W+bsPFxPT2M8n6Rjvb
aYlSy8CFphWDFfFZMJ3h8bw1po5QBddvIEv+EHggbow/ItEqz5dvJOWcWOioiyQ+S+kXq5+m3fa1
cQ5Oz1HyOENq6NE/CfBw7hE8ZUSVy0fGHwvmej4o2R9ZDJ2zr+UgKwIh1zjJuDoNhoWL7HjfDSYU
CGlEUXuLsVRnaRUX1j8VsyRRhdUZE5kpOb5cdcYYx4Ytnb1V6G9Xk4FohgKuZbLJmNUYcYqgV1ui
Fi4/kZCBOCq/aDIGo5mQqTl2/GLhjVklHgMjRzWv/w0w3X1knd7btKVEcXNgAcVFjiLZii5IDlA2
c4JmE6TcGVkJ+5552ztrq4xketw/w8SyKIIcS1jvvxUPHRimhRNrEpSemZl2DaxO41YOJphHBWzM
3Gg2YbWyaH3bR/HruhtCqRlwidTTv8wEscQobDTVQgjHqqE4cNwjgw6HYa8T9ti5tMiQsc+o+pZi
Jhw/NtFi2n3TlC8q2VZNJ0OhpRLblwvsDfzhaoIjNg/evL7Vvb2oo38E5Gy/agU0teMYkSu5SJJL
D1kiWBMDX4dtMwjtVR9ryhd89F/Got0pWvQhNAwoOAxTRhWU/R1u0u4B2BuAQ/lFne1kALDxrUQA
f+60c25rDG3oJzzTEEeRiJIeQjgCYOppvKXaAM6GKrxG8MXr8AAnEjR2xKN9+ERfTgf9cWg5peYR
jqeknsGSPQX0jQvmJwfgjj4E5zgDu94eFqqFf4VlK0Pvdnlfln94neqLDFJWYb7/fRfWjy1PYgRf
CRK8LBLpB7by5B7fSrC8xwY48a56JzJR72eYpQnsPAKx9Kz/QlY8Q0SPgooDZuV4HZ2jzOL87yfI
61EkHoatVlEwEwBBDOuE4ljTXZFgT+lL59i4hHb+GyfiyazaViRaTEbtnDfnnioDECAAqN+tJV9I
yifa9Ra0vr5Rv9NUMHFUzYYhDO7btiGToJrDW5k8mz2KpNXk+i+2eD9c1F/ufb1/qikAqkEpJJER
G6RqtXQ7jb2sCzoifSAcqufpzLQgnYiltpSgLRQpWkjEXhBSTVbTV8WdZt4Je80U0rXILdD7LIfi
848GyRUBM5R3lAg+6nv2IjIdG8JpQS+gYxtBuhbRUS9cvfkJBiHgXSup5HnZvVS29BZQQV12EhNH
jr3yyXISNhPnu7sMkCqOCi3OfFmUSw9VlOWqDVzq5bvOhih5kZ1DyiWYglq0pWrhCJjaxMCMxEQc
Vgs3smOVmsfPL9ijoEijCCnIbdkGDRdmsSBrej6JyiQr424NzX7qQQSPTCqFs0YYsIsJdyLzSVTK
aNEz6ctjnx+ATYrQJMjQC48NE3PG51iDZKo/78WA6hiSXnfzPT2D4d4qWfE3Bj5dCtpi98yUY6vZ
AD5qHob8dDTamWS0DspmwEU2yZnarj+yQYljVbQAK2WFTF87LjGdMFi31IX+c+QGlQamAEiErGyL
+Av2ULvSZP9qufY7e8kRbKc8ieK69j2NfJ5zgDKAK5W0NE5CKdaT/cnCb3GJ4YbRmQ3m9IKAHPju
pat0olkOTi6wG9W0DGiVYYh8XjTCLkYeaeJhYpbSAXS6tsDh1JgaWXlzPeAdfZ34MIFVHIZeUVIu
QacQfO8rcwDcKNhfOKWtjTpy5fTly2kujS5dM4KLXjv/FUHsaccdx20fv2mcN9HDvSp7M5fBX27o
3EF0kMitlCvATVmA5mqC0KRIMIhThLCjajcNnEhhd3K4g4KdWzZw0AC4d3gqzcBrVFqTcTk8MxAy
1efpP7Qo+6YYiaTgmZQoVwDHywwjagC6YVD0uv/kOz6X9roLmResKleXzzGnXRZsEn/OKvR1JxMs
18NQ7uCb/NxcHy4fN6LcgrsWt10C+I6V9h571/JXobB8XG31ZB8xdrmr/g2ewZQyn5xwKKeR7yk5
MUhUA1wn8PO+88NyHQ4XugISWHlY1jAyZdF0swfWBDaXFLUAWorJ5QOkdat8//cRE2wS1CkZ9x8L
b8l74HhOQQHyaGtzd12kWJhhKt+wUQx1ON4CLjY4tLAT2yBnSrJJestqK1EpbKeAvxi313QWlD7r
+ufunMmFpxsT5G7/sN3nGKyfcurZ62d5xozjZw+ztCyL/hg4yjUyUTezlvLe0nmQ2SnVEDtpbPUI
g/efpo/5SzuwnSs/KwXcew+4edyGSnwJYYqyyNSinsGawfhOd7QM36YsKmSd3RAvscatqhnIdjdC
OuNBNm5CKS6LznDvF2y1hhG+ebW2w5OBNH34igkqzcdIeR05wH7/AfMwGeatyS4HiSNF8T0skKgQ
VRY4BpljqMhzPIxm9XgR84B5YKMXw4AC9iumt0zKh1ctNReCvQ/KuFhNy7rQeymuWXLqjuBgKbqQ
Zq54e3l2f2FYC2C1u5th2TnUXLSlHDSI4a4oVol0ysrbTP9M1uV5cFsx4xoBNV2WcV6uIuRd7AbB
Po0OzKqF1E6+qTtKOpAEE1V/W9ft+zQXumA7P2EW8miV5NFiY56ul0sBX8UNJpYUGIpFI8ogg6xZ
zh2iTyJqV4ZyivSeRUAV7jc2V5ZsWvSTAwoyX7Oq537sl9n6xaNuOv+sXn04WkexAJn8vlbjYEqq
Bb2EI3eV9Ccbq8HoxyseOKRMVPizv+EcMIkdk3zWw377IYUAzsB2zd8syvCixaIlvJxESzL/Jh9b
QKzPo6j/81jkgtEQ/4dLcUjf5r3ZfvoGXJntR4K7K/VhVs0KCb5DS/FQ5q/sE4JQYTkE5pattuLR
90w9wLuF6Y3snah+5JjCLMAxipnPtVas6l2KemCpGPcUZAEukT6uqAKqwXL4qfVSbIAKrzwdkm7z
WNM+W/ehzTFw6MQxUQMVGYPfrOugtqhYavE7A1BQH6lxFwlgxKuUmMEIPY/Qr2pjqZSZC/ElQP1Z
rXzBp9S2OIlGFTa10VfRNpAx1APDdF9pW+17eqPGPeWiejo2u8a3nhaPIpatRkx3XMWuZepAtYrI
NaoiTfViDMLoh37aj6haMR7lrNcofY495eGtvNOxNetYb54IjI32WYTZUX1UFe+Bm9qWvMWCRvAb
OPu0GmyvG2EByoEWr//RoF5VdJ4Wq9m42GkYRfjhVmY41eWLjbYeqqAkY4F5yolCmj0HRTjaVbPk
M+40Pe+Pm7lHF5zXYJvwg0Reoe8S++47cs+y40cHWxDhFJYSVvvAfGmoOI+WN6E0CZ8sjUj0gMvg
JeZvQtIIxoYLV9+h
`protect end_protected
