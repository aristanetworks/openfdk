--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
fIniJquc1baLa1tk3WgFZyo3/cIQDRjTJicSNoKLXFGfHchOfd0uRk9UFLSyNEzK/cLZOb/OgE+M
yQbHywODkc8JedWWDLabtBo9Sq0esWa0JepCrtR+SP8PWsKHGVZ7tX+dXKWr9mnaNRLo+9vmqWwH
6+YrwvkevClCwG3aq2fd8vVQMKO6zEnyG8+gTTiRFo/5Tf9lLtxxVxxvjDcdGTSRMwlOethJQOVb
4kwIsx2aRpDflvHk/3UW1KdTuhx8ujkVGr26QvyRFxq6i1cHpQ9sAsIi0Yk7oa2iWV2cXf2P5a+R
sOAY76itwQ+UEEuhKmICAYysIEgXRRyxWzW1pw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="UIeQBPZSn76U2diQY9FPigQ+u3kYssg3wYXwtOGD3Aw="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
NcHTIbQhLXqNc2XCj0wM+cfsBVYl44CGxjHy4EzBR0envG9/5zHC0M992QLAoYnmGgEuIU8vwJKa
XIvc8YBPqTIEk3Ed99SWiYnmmVv45w3bsVy2QFQ4kR26Y5EUL5JD6RQz4GPfwUQ3BjRgKqZooSFU
v55Q2JYqXte+QpF6ZJn30DJi6M7j2CfjF482puH5cRK7TOKezRERya5ZLlWV5ELgWxCXXux3RH6M
mxIa+dsxJGNvyGG2ygKfsBOrGb04TvGaBpe6yLxAd50dYdW1RAvlnyGt0hZu2TVa7kqqc/hcTaZz
wIeIlSR4W39elQG00DQoQGxKR7f9Mic0qyBzlw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="DgnWnyAQTGHGHpeVqErfRNDyoAqdln/DX7hE2xX1Ynk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3888)
`protect data_block
8SXDBGoImFgyJKaAkQ7F8C3rYHUEk37hMLoJPSGtDGNy1zgH5gmvGMmugdLyUdLrc3hIsyzcP1Hn
3P8GrQc8+O47glZAPlhui+eclIIBJZJpS3Mmw1XjGomzn4NVIXLNCQlVC8RlN/sm2BxpwHOYnjyh
5Twg/Qi85PgJD2JNEttkF9YKotxe9nZ81iSz4hLnQzDn/qpZNzPTawCxbE6q7KtvivU+y7q/qWEm
XSQw7Gviig3Vby+kVvXJqfVD5NFM3zc9KVlMhhOYY0VmliN+13NpIjQMNstm55ZPRUS90FXiXM6H
b0Vh8YiDbg5+lA4Q4njgt2+PXEdVp7DjzcCZ+ifoVyVDYrDu1ygHfT5SlNNl0S1A/s0HhXFvgjbZ
FHbxyRMYdmtKNstxUy6kX5aq0t9rzvZu2PLSNfli2Nbxvo1q0t4bNqTN/Sq2hK8du+2Ko8CM35zH
V2scVbva36xHfeNrd6o67HOGG4zJ9J/kqa3VMQEO5Q6YmJdj+Y7PDTNztBZTavLETi3ztXJgtN5K
YsNeSDnRd3CzzXtXSN6yaa2rs14LJSRkZkGSwXrjJUvZ9udunjxqdrfziSFUOmKxLiyYp+z/4lA6
8h/bQ7KgvinzZH/XZgbIRwuBBHqSPorpfKYr5ERCoDg9oK8B520HB4yMy6B8z4n6jKRIVysD+k2s
nI0K0WmXTBsOVh48s2ZSQzEldjwgluOz0BdKiiazUjt6Ibx+UdOXgIBuc/7Q4rr4Km6CRJVajnRP
RLpQuRoT4XXxzk0aFEwvHqBTUfExY3nEwmfjLPXK8VyjgwR5YZjHEyB+CZacBWcYWdO7Q9aMfVN1
qsx/glBdl8yr7Oe335BRdGEZ3VBfYn8PXJWHohksOGVYvfpPIwvwQR7iwjWm1+7eU8m8BqmaAvt6
MLtzW1meDXGFN8zMJWywWjL1eesjD6pGFVOFfsToZqcyHls1jy6S46Ix3Xvuw/3IQxlkxHU1BP7O
8zcRQv9mmtDmEimBmF9Wk3/cHn2Rq+ziP0A3WI5W9BhH7l9ndKqtbvDTzywIOWY6ccnw0HiTex0b
Sznrk7YZsb5ca6/v0qXTHKkzCBmuZM13AX/Ia5zxr0WEYaG+YbZ8g20Oc9VMgfS/xZpMJlbYb4C6
2GgBUITkU2Fix902PltiTg0vnfEc7Xcob1CDCvCl1ghnlNL8ml3WraLtUM0M/2d8Us9KPLwKNsaL
CJP8F+gLs6U2kILzg2FTkTg/79jAxWCwsjRx0piS+LY+wGaRzx+CHibC4kXi0UQQjV8I6mDJt7Wo
6o91oK59OHU7F79zdQO14j/Zw6Rtw7FAqWHLldXrUeSSYGENoasSTD3LIHzg5vAbZmdHHPpA0Uex
LpFS7wzlg98HVP6rYkLZU/wUI1fKKfwUidIzGepw+Jlv67DBQY383+PIDhaL0Eydh7YB1svfhB9W
AuIEe9gVjWKxfqsEclaxDQbh5j2yn9xMjK/XbE7RcWe1BNtc07G7SX6jHiTjTq7z0SQ4KQ33NW90
lWH3XyADLkYMSkZoByGF9Gfct2bL/LJKOY6hpPqxN312gN0F3dvhx5l1Ud+Ra/g3cqfKpfhBPjAn
Qj77nqY4jShUMrEUu9i1SDD6I35Ei+W3WZLaiZf75Rdq9vnbatFb6jRT6oGGq9dGJ8Ch9FF95xcM
BSo/4SF38zJjQoV/y2AU4d16hcufVi/XkhMeo5Y27ANnnPi42AsCJeg+1NZxqOXjB+d8Sck9dINF
J/LCWe4b1qse6aHXRLgTHvz0XJVV4JXqvbrelUyhctm9Inh2F05QbCepqj7qHflzgjnUdKFdJSnq
UTiV5ua9wmoXh/jaIEze0VlwqY8pR2oVuY2wSsJeQV9CJXQW2EYfUWJLuX8f8yN/itbENUFV6pIF
7zkBtZ+z/9pY2sy6bi0NTNdFsHeFGqbkC9ezxUSkFEiv4zzbPXHAb4lZgZOgkOVfYsjyecfdfmNP
11Yx7stUA41VXs9zklGIVk5cLqnq/B0wc/a4kV/OeHgieoNwH5f8fbBg1qIZk2QwH0oVJM97hyyp
JFe1NgtFKgDBn35s4t5Fn6lGSEVHFXXMvs+mXsfuJ3k7N5qyPf5L+JCBo9rci9Yvq4/pltOOpurK
05i7upAJiwXrg3fJ8ReksIXnMfI5oUFI+j967llbNReE14GO7y4dkeQeGSmnZyI2UGh46UqnRHto
UM/6BhnbMPwsUN43FG5hHYTT+2+sGp/8lyr6zPrLgXr6JiWflAAxI6ovfz1FYV+b6FOFiKmRPKgS
iHcMsJnRr7vFqVJIWGaEdGxHI3+nBDKttlMVreyaNGvQx4GldE5iE59ahWDHP+Rkp1c0MvRIkVbz
8ZrfDuktmn0bYAGEgLFUy/B7ULlbzsEFgYHjh/1vHziea/Cg+G9jerodlzjjdMuAi2HpjgJ8+VFQ
e4MzdJrDEArv6I+xK2AOQN/QVzKEHDQqThe50EfIEfRLRinX9b7XlGzC9JdaMzjzxA3PPoQcDIvZ
xR7aag8w52xizMhpdrQiopwAv/ce7+kvPiiRYGQZAVMTOBMoLipIkIYnKesjHj7EtLu23AkLgsw5
KWIFOhIipSTwVQXnyxCqzk8XQzXB3u6vzElgpWR4L8kCULeBuR0o3BsT/pzs1IC0nOjLJwG7kSJl
mr9FwTRjsTAwx2K9aPsCeOYbFjKtJKt89ffrXuwrDMo2bM+rzfjk/4XTHVJWYNsZ7QdJMXvZlLTu
4dUfMky5m3aaXUctF0MQdXVuY4pxL5SWK1tfQPM4LAGyhwOW6vZK+jOd91m9ON/9GoNtXgMngZRW
VJempMku8UN1HvGVFOUm8nx1gAmnoI+N/ucrRfBO0ETuniKFsf0jAa6Zft3TxXZOUCCkv3Ouhtgm
cCC7kJhOrM2XCPHU6QUQ9dsjscbiC10/CAzu8r3AixF3pDyYkGWzx9riNv/Rg6nqnD63ogIq8QmK
HapmUPDv270UdFpuOQ1AF7/bk4k3vXK3plzWj4/DZ7LaR/hWlRbj2DJA0/FU9kqYLmvu3uyX1A4k
3Wq5k6t8UX9wSssmaNW6l4ugKEbcdPtbC/mKR8L/L/QkamCYl4L/jOSkkmjZ7RCHmLs9PcACcB/G
l6DMZsI2gSyDn0y7KtlRjyU1dZUz8MZBJxYghibHh4t0BIzeTf0tNnIZH4MGm5lNcUCne2WKdV4p
89Vin9B5/cx4kfPu8ub4n5Z0R+yJis34RJJmSghnYkdv8Vdnjj692H3TwOD9FVpOMekFavP55siz
3jvAuQgQixiqoheoF8spyU4jdu2u7D1cWsn8aynVh8W7DKe4kZiKRTA/aPi0BmQmXo3FfBIMsZ2h
SO5KXV3w1l4xIHcJqUqEZfkEWgO9LkaDp6v101PaigzEdwUSV3CD2qpHSpQr0xw1NAdrTsbhar0a
Nt/xCX4gJE7pmm46UE4aQMADTJ5BpRAwz1SKZ0TSpibcGf3KrA6RCpXMjxz8cFzH/kdHREs3yP7T
O3WKZfRbSPp+WKjpOSuMe3BSFdwxVeyS2tAzQcf93y7n6UpIEHbl8WuEO1ZchVoG16sARZL3szxk
ZppfiFtd6rZRXUto/oDYiWMarMl6L++CgOKi7auE3HWczQcBsRD2kK3rixB8zpre+IhhOyKgiVXc
zR5B1xuLmkjtSRZtZ+NQaXvr/lVvlvxYY7utDRT9DM+BiAguIVBRCY3efWcr4xLFKMDLN/Lz3LaK
FWIZImKk2F+rbMAcQH06vNP+vmsZM7ZX7JOTchBMBBtvVZdRHrPhAWNfSzHJiwNYlhtRcaZ1t1mI
14dbCwvQ+CIQCxtm85bfVJ7qo81Y5EAcbQf4Dvahl27X1ogEJIkPUMSiDHA4TMinpcz3xGPIzipv
UVWBnMecUNBw/7y+YbZdcbUCK//GeQ+ZRJLhERKG2WbIPt2TjH9MC3fFFZkR/DX2sdTf6O0/s2lW
i7NswHGvFZWXfkLb4nDu59NtOr7YUfbBHkeSVJXquTQ2rMSuxwazBOOM8sxJFyZMXsgQtF0Wf2JU
+Qxeod/0tPNwlxGEghFNbonE/GiFvuDUcFVdiea0HpgVHTYLPXnH2Y2i5rGLjjGJT5U5HdpU24nT
2p2ybSJyHGrWe5kWL7RREzSmVOl5/IhxOh/cOclGDNvWAuuEIUTQfRDpUn1YhFyjlZPfIdZQmBnZ
wl0/C908mimSAJckXpAK8tZM9DNgTYISSPhP1dN+gbScp5VAeOejyfOktMk22Dr3ZG5LV6KkN91l
K9JUaZ0z6kyLOFXPIk5KSQUaUR5OnNAP5dQDJUCZVePwo0vOEWiU4/yXP4NABnHxFjV3wwpMapvV
d0Ob+QjbDR5n6bXABPh8QbBw5hdOAzNzQ1jk15rNpi9IKoBqXg6aU4fHlqRwhH1vSX5HGBuyX3Kw
exTaR3H0ZM5opga2ZwcqpiFMaic9Yu4g9/Aeo6XjvcnzsPtUg5o4JhL01U6Ho4VRN5/+YYyCw4yS
VcHwqV5PE1OsylBaC2ORQUgbr7nE893UWlL2DynIfQ7bNs+uMitHqaM31b72GtF+BctFowBWP/Ce
LobbuAekg5/ZokeL/6+EvNGMjAqrgL6+/Rek2s0GLsGeXzDOokWRde3t/Wf03wR9LW+RFkW7RD1r
qZMCKD3VEXeYal8BJhpVRUOSKIS4N3v+kwAw4pb2Vs7Nps6tTo70wihTIZMnijmW5ez7tJn59WeI
WRsfU2/XM8ZtQqkdKnc1n0reikHGM9SIRnzcSJovLew0yHQS0eL+qCt17+LrR4jeF/g6mZ5fbfUg
5MR4u2wX//87RdVi7aMMlkCaJLJfvoofuFZWRN3EXg6+Ks37cumIZapQXavHp77h/+PgzgZa0FvK
WG0AUJFnPTrgHYr0/GIciNlBnZ7Y7+A43HcqhLxgnW78VWWPQxCtZ+wxS6HGURAX5whs3fgsn1q5
13oMMZsIEKI+6LcCO0FRm+G/Hz64tHuD7BykpxCAw+3EFBRtLsgHayyD7UjpTrr23sBxjP8/Xn3q
iPn9SVqf9y/YILkOsDpnIc4+jj8PVKEl11+74xXYsBzqRmbXiQGs357pM7gI/U9H1w2drDBCup8G
f2wg6fnuIEDCfHylc8deU/NCODupwHSNyDOiIe5ImaIS477O0gLwvVQ7pCW0vdRMZg/N9HKBBHFA
ZbEtTl0ryIWwygN2
`protect end_protected
