--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
PN67V7bnS2NmC078nt9vqmr2nP79uJLe0jJu2BqCoJlBttrlnf/eo2nePwPWHv7NUlAOMC1AKb6g
B4B/94uDNuy8fZZUzoh+Mu1hVP1guv5fq9+pQuk95SmdMrhX8Mp8LkhB62c0tzpxPNGM2SiBo+0D
II8nzjw5AFGvNRoReKvRu8dxazIvstJ1UdmkJ453NtCRMebf3C1bey3rLmD7Qi/bWdium9IG1pYL
2lvgvhCeuslp3uXo4Tk9goWoLQXJBfFnEOYeygQ1/gEYkV6znoxIEpFY7Q+ZNovo6FKwvElDe0ZO
fFiP0giRESXQH13EIkaO0poHS+qHA2tF+lT1ow==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="BQoLPIWkZP4DuAsP8CBldDLQyCM4aeILhAIG8RkJxtk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
qI0FR1ViCBujQwCRrA48BQt7Z3ezYhb6DpvLA2tp3LvKE06ugRCcD/NpmH0ur4cTsH2rCDaZw3kS
oYKeJDcR0QYpRD2sLyJ3zjtTQn0f0V+CAG5pwn/fGCwrD92zi2h5VPn04LMY3tQhWQpFgAN3wuUd
ni/EuL93Vo3BSi/R+KIhk4UOr5tb6ywJuGMgDtVtC8ZuvhXeljlY732JL5A8G3VJi6C4H1Bq2dAz
T1S6nawOMNoG+VFl6Hqt1SsO6iJIi9tWbdpDwUMWZPp5IRaIJiOMuX69f8DBTyoIQCXvDNcgdxZG
q849m/n6WZY7syloU65pQpQAdUJQQ8Rxi6glGQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="ZVvCGnVukWdgpiqiowKXdGLKW9vbr08Qx3pBjqfRCJg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21840)
`protect data_block
MdbCGClX0QEJek/2ED4Q2ihV0yVWFbXNsWB5c7sM4Yj1/QFF5nPR6B5KZkYYdReCoY6fCh82BzLK
lJzAwpsVBjBOFAl1ZPSrRCNs2ka6xRhYoo5HsSFmb8iTq7ORNNwog+vsIEu/nGiuTpUJqGJo5pFR
r4eH122mwmXz6gOuEBZ+ec4uS+JH6SXjaycrjTTFPAgcnwWWznJCVyaNoQ0Ua/L141nWGiXt+fAs
3F7OkDlgg7+fdRCxjVYp5djg5BTlVhXqNlWKe1sCLK6wJzoi5Ecq6BfLqApTcbqha6cHQNAq4WT0
CdsBVsKz0EQ5/hOvRi2smX0kI3kNn0Sf+Qr/wluOK3JmFBAbrRDXIS6NMOrbpxJYjzjx8B61mM3J
86imn66/K8DrXnOm50be5q5B26eg6M7s1bAYhNwxht6EbxgRTIwLN+3HXjDlu55WMQo/y1OtbgRX
cnTCAGSaJBR+MbUtfaNfR0NkUFP4ODyvb2yBQaBbkOh6F4R0TPBLd2kCdMnoUqAjmqmHeoEUT5t2
FbJV6EYP3veCHMviCz3DJM/YjZs8gBpoOBRGGkwgC5MTIJCQhIUyLE3OUEwbOLvVtkn0/aoN8LV/
eXoyVLlcVXaMkGlC5+YsfgNQv3gB5Wzt4Om+/AEUYCFCgOcKVGc2YAejxeyjao6DraSAzpv6NDfe
3dlroB4TEGfa02ELJ4nmCG1znooIJ6SGIKI/S0JRx6nqqajfVWPIzKX/kDBY6/zsPMgssWFoWlW6
cp2/pdAeY1t/gN7fqiwMKPGRF3XC0eP02o+v/0BFW2PTuUZ39xbj6uBKmSaTUsUMLpVsP9dx/Kbh
SL6hIkt66+NgZWs5v/+kVEmMsC04pW6BXzaaAvYJtrM3+6ug0b6Moz4/Uj1h3+zKqLlBm8DeLru2
UtREl0NLh1obJ2QAG1zLi7RGiIHepKl3jFhh7AqIJhRFeagnwpuvPvV+5tCltAi+AnHcRyh6T6Zi
FtDv5LakPN039/ZR1IBNVWytY9+HzbUyHL84OKYrAlyMEqgLgwp/+N7gZHpKfaNq602M8L8ULQzv
j3vI/oFb8eBHxWikXeK+F0iZf8dWqgPfc06wtfWQcQ4jSyp4pDulh62tdCbtVsja6E7ITqnAGsPJ
3cGoNyZ8lbFFxqWUbBz+iroACdUbaIhgSUSgzH0P5xtQ/8zjjD+jQPLI+95vG358Kyjpcxrrrbz3
gDwDxqCT/EazfdckUlYfYjwykTsQDExfxuvD2/Rnqs2EvL6jye9nne5woRLVN3svzxmug25C857Z
2Ie8d47LIKwu9jnsCCoin63Xa1dJS3Xv0By0SvBbPfTW0E+Cs7df8rAWbTznc0Ni2J+ZJtnZuyib
/bAPUJA/Aa0rRihDwxKnK8rTlaDJjlx19A7ctGv1rdRCjVCl0JH71bQG01BaubTmjJSAjs0rcPKN
agzwmr3VJBBFdJfEHfht7W9P+BBjghzH1r6uo84yUyGXfyDMUT5toveqACUDwK+wtTkB2r5uDxMF
CbwxmpO68IS1JE1P3b1t/S15qQQTRCAwQIg82toSx7S0x80ShF2dBoPjTXSnETvtQ1849uKxGwBJ
GNnj6p+JajTrFAU1HhigHjsA/28QfAL4pYbB9EHZw6t+lzBIvstXF/sierIDoP1VImuGclCuFd9L
kjeiDq19OAyiLDzDz89/V7gcFLVnmdS5rXiiOA2N6gqyXUSogLWYo7ZOd7V9Kc5mulFLBBoHaxK1
X3fqc8Nli1Ia7UyETYVpSxi3kQ4WI3knl9PdNGtvtVYNXR0OnvnU3wKDbo6iiGvpq3AjvMxP0FP1
b+W0PhBAv5UvlH/0+qUGu8Uj41HBAIx/WIbKuBKhWxLm7pzMtHqARud/xicwfg3edxfuj2KhKMRC
2jPBjo+WBlCYkYk+epK7i0yERXy0Yr5fMm3SDdpwZ1zBaZdKty58M5FQyNUPsS1p9THkMUZY0udL
vEeIT4E+FpRBSN+AcQUFo46skPT9N7yWpfP4eBYCFyqRj/FhyFHpg4Fnmq6TxyAA+g7Ee/Jl5iZz
bN/KFCAFjTj75ObT1bi6tFZ0HYdHxjomOQ3G3tT03Ctm3x6q2ybBjVhIFMS0go/8n7iMJ77/n/tp
/ORPEBKE3N+oBcgq7wiDi+JDBAwdb+1GWrSpibkjAVZL1GX+j6zV2Gz5Tb+9iTGJCkIvbgyd995r
ao+xVqszvxW5rci/9n8oK0PGRDmDwqdSKb6M28tD3jvb+8XtarkK6NTPmG7gre4TPBM16P5eQtoq
iRhX5uibSboJ+M2lNKsvsyetq43FCcF+8h95z8cYBABqCxOc+wd751jb8rADbkfLynpgt5yJi1aO
noJtHpiAO3mK2/yWtkSlKh8ec3nBW2MXSo58q+EW5wf+4bL+iJRgVFBqADWAyibyLRsBvC4zXIDN
HwQpqJUUAj6nQDrN8+tyFDSgf1AZyJ4i4GwQZnxz7oR4inhig3KVFOaZLGGid4Pdym6Gv7gOr5xD
sX6Q2g+HHwPBo2ZSvGV/ou1XNtn8UoqK0ELUVH1Cs1SBu9Bs5kTL0JFz1ViUAzBavvktDp5Vp9Mh
tw6WrrFvrvzYTtRhpI9yb8KL/gnIQ+icGn7S8+d8nC5TLu29dts69mN9RD7xaB7m0b7LTMGW+RSy
s6bGTgq4Gw7Ljk8ItNlW4dx9nc/j37j+6cYr5CEXHTWW/wEtAZ49cpT9kvzI5EcXBzdktPt+Jqn+
hPoQHNHaLKiRA3Deiapk0oK8Psv8EP2S01vPzWEAEOSeX41Ad33glDlHT1CoR2UaiijwzR1qbhrN
GOVECBLpcvzGcqG5NhjATxdWW1vhdLsyENgzGfMIIIL6Lr221kK3wss+CjWz6Ov7doJ2wV90mgdZ
W9CHspQpPa3K3CasQ/b6E02aSzrz4/JoaGy5hJAgvsec/W4TtG4Wk4CTqaFigfv8CeDj7ZK/nxGr
KAz5cNWQAAGdCg1g/v/AnEjDBh/JbpOeahWVFqRR1eRzUkS5Zd0uclOff3n4dPboB+6C2be/QZ+0
knODrX8zEJHKgluo8heCbbuKXweqZ7XvRMFFgwYjTM4rhTVSHI7MtsbtueGhfvw30egDzf22GgZP
mcknAef8F0bnGLFRLu9+3NMrFSNxP46HIZTBVFlhWsQjoCmASvskwctIzVrdyzNVPYB+kXpkBg5d
7HbdjTwh6oDW4Q5wfsPPwRa/Sn6iAfzcwZtExewvxrzsTvzRO+5/YJ4i09Tx+90dKU/oDKfy2KpB
CrtDv5rF7X+ALe9QEPytc997rrxXUhIriLErD2M101farjePSz7VvWBW5fp3oYY11m5V+fG0YIzx
yz/KYGaDC9fvfC8ZLUI5p8z0ZxDVzxukDFR6/h2QYhfFaQ3vioGyFXFVTXx0JXmDVOHfavxuo/0a
3Jmo0o0DP5i9d73jPJK+JL2EnexVQaOsT7v2Wd4SFTx4LRJmdTKHAJrSc7S9XyQ+s24PZt/Qmn1q
XxMwCgMPbzXsM5uSDe7zRXgSzbnqaVstri4fkvxbZ/xVPOI/kdI3O/06JwG7obYuRdO2rKuIL/nQ
dv/ZXhhXCU2szFcCxiNBFNPl7/EwCjMm7qVQNBx9aIxBoy5AYCLWReif4R1JPTJHbHgJekOXFtbh
fyCkA9wkM0Vb9nu1LKk8SBXT+hRugv1VGqNJ+0BK4y6eqDJFkkiAzz//iQED7q22I9ZO+NU6Nqon
yGz6efz7T9mhbJDChTuuxFODcEmxMcrfrMKb/kEZQs6I77pm/stnBR70Ilq1BbBYCvAriMlFKKgV
TOy8l+OQmPamI2RmEDkyGy/Wa8sPIKuWu2pB257567keqYrvHl7tZ1Vct/vXkXhKzUIgYh5zIvq6
DbbaDDGx2C+ZwxS1TAXzyKWwD0lRtXDEH4uO7hkGk6zQM3gFxDTrVlz4S6sDidQS2JyQqvDUXmXN
qDj61gsEcxA/eLtOZoTay3FHaDZ/066XN1nOQ61M4xU8wNVoAxJ/mOw2aPbJk9aakYC1wmIcwLRj
sxZNLjnBoofw8MRwx5HUgdeSzqC4o6QOE9hJM595GKK4BNCXOwgOK3ZFOJHsKuphg4aS6/2nwB1a
GIsMTurrUbJ4/6FKProhnrAC8u3FwJXBzxFVLdOJledem/rjCSuQFgdL1t6/H2/GBuiyVeqWOw06
DL9uGT2N8iXcDP/PQ80S7PZzdzJWRQF++KCnC7S21BkOTPaDcOaOlyNw1Hc+lGZqNVP6iKL9HTuT
SzdqO3XGDYEnn5Q2C8Z/NyU27oHdzHW64FQ9YpFNf4HpPzqw6PcYxwuwcheyWk97oLRiRdcNLh5b
ZIyiRqgBFjPXqChUeB4BJZmNGE2LJkyDpqg1O4+886Dpzo9WVYM/7g/3WOs6vdyLAA9fOB6Sdhg7
0dEF6QtKrfAnkliv5Bz0PV7Vkbt41s2f33BjbLkKOao7b020aM4A3dHJjrFLJcBGmymaX7VFEvK0
6NlB9Xnz57caxzWmOeHffsMQcXl+EKeRM/U/UP4KAUu6x3N6ZSMaqPsagCz3UvJ+hfN45pfHOmpc
SawPEpe3HATbFM95K7o4+anTp/hkRSu7OBReBiOzAlw/HiV0EOkl3eZ7eEfqH8BWw1CUyN7oiwzN
QlrmJw5tqznWu8m5HequozPgp1ACnSSk89l+z4iyhImG0ZyxNrjB5NLJaenkcvYy82hpb5mjTOhW
WsjjbWOchGnPTKRO+FXSaRGWEFRx4Q8bgG2LAWvyGS+L01tljVaorFNSNPdTW7m/o+EMqBz2Nzg6
0jY6MG/PDeeP8C19YBcYsSsiLgwdLZ0/n/edbijgjhoQJ3ZA+obd+4xynnLDuPsa5BoA+4coT4ZZ
nbcgV4WQDZ/jRzBh3j6ELH4cIikiUabRJl0FIyBt5Q1mgB+bzWEM8agyW+CjIPoUrXQIo77AEUBg
HtiltmAS1zZ4+qYvKa/PW9tkjz6YhQKITgYWSldEAN+8azz5bhV+Nn8HCugrqf8sXOX0d7PfP36e
komtTLtIWBi+BG4M1VowByBXqRVIjChdZucfBlVxGH77cGn4YNjpxRbshsY68erAPAshJxQSyuC/
7/9HMbcfAvHpItL5eIMWpz+eG0zOJ9Vbdeo68R1HiSKDAwEonROUXxc73mdoI+2YynOTml5KcNIN
Sr9s0ketaDzz+wzptVVqaBNuNNMeltFaRlA5YWW2/TNLo1SK/AeMhM5JjP017kBgjnMpz+WEGD4j
gKRXvLv1PO54QiYGm+cpZC/6Ledu5u7SzIsZSiolsYWkMXA6Cs+GwktDb9qxkLbZcjzoByDuI2wb
YusMstX6pNDRiTN+viHQA0NUv7ZS30gFEV2DuwSwnZJ02j5R33Sa/v2BTjE1WhHobJ6oGsjezj8+
+SSAVhjtzsrF9fPs8hzQUvW/Eb3l/zOpi1lTbUfgRk8I+rLWXpaEuiXjukgeEotXq/U2JOoaXcLh
cDnqDrz2i9S/fsAE0BCbMVgeL6+FbiEe50mFTwco+exkMFSXTjpE/oNr5W3prkjtIXY7yXc+g+/b
BgbSkGFAqFw0STM55N1kRV+wMqBgUMkRBm8bvKei/qd8lmgWvvJlbBbOWs1qBfbjA6yknEeRSAmW
V+idU43KnYvNRqmVcfLvv1J6B4zr7GTeiPmnp5rOj/qkenj99ttl4uWukkz5VbtihXCf4fWW7X0t
f7vwpqdZPWBt00W2o3kFKwQA75C1iyfGc2FSENQiz8rNf7mrkOneBcZPB8UqlIu8ZeF97aEygxVC
Y9iGWkFPslU+Du4EqfP4xOCZ4VvytIcGp92+2SSZk8OggXAoUG3OABaiB0hzZW2RVifAKqrEf3vV
O7rpKqWyIYSGtwvTwNwoINY3Dw5eWlFgTzmTVp98KouYGP18Mx8tzbZvdqpbb3Adljcw/nBMeGue
V5V+EKUVL4qaMCnXHgRYaZH8mqaS/2a9OLaMNYfbQPMfcO82Md8YuZw3icevcvmgoHzZR0oywqYU
gWehKtWrij0Ktw8PPtEE1pH6kzfXRZVhDi03py0cjYng/SVjpmqrRbzjXcc+hV9i1WcSnZNa1ghe
v29m8eE1pbpoyOS4Hls5NL3sTWbYY9T6XiLjp987dvNQ0mdjpfSxwxM8QZeM4pDGTlWT40tYIxbB
yup46IwuO+H3cRB/FbAb1NmdoFZwqo9G3VPtFHrBrtcIqOAyqr4hYRSzmNb1d4zrwXD8BjJW5ekr
VVfAqqEGHiRW0ojkLfMvYBfPaLv6l+qi36Xeaj7kg9hbkJw9n7i9qADoWaO027QNeihx9tUL9kLi
dNaNvL8efTruF2o5kHfq9dS0555lr8ySjLteMQ9EAL4iLBWj2emKIjEmU8FAPoHzfvSSimjIVCJv
oiGMKKyRM2a9A9ruh+5wcj6gAMhXr8GNHfjHyz7HYkejiheo8QT8TsJ68dfBIjmrJ/5LKLoEGeN1
4TnAwZ/4GeuI+PmpCW+lvI024iutpY4yKoCJszrZJG/ql1FL48uQdqkmOCMoroeMzmzza6zgx5HS
GI/0Jmdudk8j44bkKlYQ4NnKkawmsms2vWUncq+vOmlY6AKlsKZaJA+BYCNvFFHixIHiqlwBHWkr
b/zr0y873JiGidmY+Ce1Vm7rnarvW1K0CC9XHz0nIylFEBAInwl9kwxsX1kEaXvXg7GN1ufcsx9B
KFs2hcFrhg+152lEiRj+LIOJF8TfpSzxSu1mOgDltqY1Xawj6Menkre5VBwohToV20w0Fu1n1knJ
r7P37wfZ1EeSvdoow+RdEJYQP7SWIQ6BZqYh+eSGI+ac2ZuWfAFVOXYH9CghsgzVgUgyphrBIoK6
ADC4hrQJ1/aAk5FaKqoHVWhwc4U62sv4zllp2mi1LP0yLNJMiKKHn2jsdkU23Yfk0nrkER4P8cOH
qxaai/TEYTUDoQUECuulWF0J/SuQZDqpunk1EOoHfkV73AG5k3+eN/7Or83FllkAPXNof/Tz5iv6
qKAbYBmo+j+J8mgbArudn7SVuDn80XHuEraeUDfEN/nxMqciLL6KQHnfFXr+4gsTJZCs3y5pSmch
vR9EQjxc1QE5x8mzbuO0aQZCuDAMDO5b3YWr66t/58C8Is4wCq0c2LwfXg+6/YxMMMXQUcyOjK8z
NwO/W6RERSMCBXX7wcPwFcylafvFc0Rk64iY7Kw6NwXg8ME5NKTHIRgsPIKAuQJoyjlqULSskAOd
A1sI0WiGpBRAnwaFGVKgyjQNro+6B+X3pMVtbYiNuycl10p9rUiQZpiMbFMk8kM85IKHyt4Ol+ij
NdxlkJsld1ZBMHXBthPeb/jezl7sdufpuR6rAy2rNoa0/N9nzb38TSfdgbrze8qRj8VbWannLvvc
N9jTUr4tkQYdFzN+mKN8ucUhO5kwsDDzCIx97EtAcpoqxsoqkeyiutrEEhBZacxGtlcTKGTu4E2u
IAhj4QdtC5kN8lXsZUmNVue8C8CyAUGCfXWzVEtziq4V2uskuezUhIg6mbEc9Cm6yX91DxRToNhB
VQEZrVcA9ZVVZu87i5JPCq1rdC4FLYRFwA1VmOXFfR3vkdRRbBDyNBj0eRnr++2B09TrcQt2V/jp
RVRQCIbseWytgUwJnS/cvu0rLzMqR0mDewdRBvPAUcQzw67dQ7tOKtyv3F/ssoW8Q2Gl/LFMX16H
2LKPcR0OhEIkYuvPXBUpyc7C41ewrTaRpld+hpMJ65HncXNMrNYsYCVbeVfbPY758aZ54g+SD4Sb
O3y27o4JrbYbGPo/HcH4LY342HczYLhLmDxyid19NhaBsw8JszUcoEMLgEUPK1H1CyDVGWwaBF9j
rs46/PkB82uSdNU/JFgqt5m/AEQVsMNSzgQDszmrfivB3R5lVPQG8TP/WWI1PA5rEjYF9UTAZXVM
G/IytptFFme566KlW+hJ8xIDmzaLdgHNGFMGLjPIUQCagQvHF1SB5rq9wqENhgNa9RvQbMcql7NG
Rmeyt+WC/I3ZcMElDu0Ic0ISITumwLMCxdUOgbWU3cqyuDVlna/tW95jp+iTvVtKb2YlS6hLp2lT
T76+pTeKqmh5D8SMjU/LGYc0R/bFtDZp9GTUC4z4ahoTthqYO/5gVh3Rt/yfIPcvBEdZ+ma6CN4A
0EnRvVdxxvFeQ1saklJ3wIOs7WQT38jONpuV5unWIYYEfZmKBbWTH+IlGl6YM1ssxHB/IT5cp6n6
suzf2wd7naAEkxp4AwT4hIfQ5lBYb5C90+MpJf/IHEmOfR5bkaqEH3Uq9vtlhCSugG24SNUAyNAF
j4jWCeFhD2STmqGBgyV2EtnbC+VYV6a7P0NiG+B1BYo0Kf7MclA2sL8D/XLp2qHqtz2BwU/aFuLf
6wvPW2A7vaExH0n6WwQrQqOABcoiygRrNvEAW9vnTPcksDOPpkhmMBhcJYKXdVSAEEP83otTv2/M
xqnLkvu+KL51zJkqRWd/YSqOQpdCjjmxZ5kykG4rt+C61FVdt+VeZWgqKUzIlvxrkdU6s41Rjfkx
4GPevH/87F3/wwq0Bx+rzc20bEgcIHyFK/Vl+vUzdOltCg8Iiuqeni9BrTaNzVoRNlQrjEnt4Nd0
JqT2zwD8SH7Ys7ergoFX3htW9kv0ZXz17TP9WvkaImiGNh4zxNinkGf17Vctx65c1uLec3wfHzxW
kdq/tVQkbMx4DrHz5Gw6ffVqKJ3lO05vnNVAejJOGPh6gqFE6JX8rTDeMspUYBNJhyV0Y8fTD8rV
oO02gUgZYoyN9RpRtw8dVzW4vc43W20Tx2LbVrVrpg1HTA2ktBHAv/mPMxrqsRY23Dv9Oht3hU7D
YHgmdfSuP31PZQfdU/OJpHT5yzFI+PY49QEbeVG82MNJlHkHHsq9UOwji87PK7xw8aL/AQhNNfDk
/UJiBuKng3Apo2ngFf5VtbCsKpcGSX6rcAAGC8w8GeuYiL4Lt3ldMz6MRSkLxqvL2bPtv9eB8T/c
hpey72S27vDlkSW/5X+TrB4oTSrPZfoZi73bLtdhMPAg7U9aO36c+lmD15pAHH1XF8ZjSoxAeJH/
81RstSqNQEoOuMlzDcvanrgjtpJ2oX3NgXTNpSyLP58YDw2TnLV+IZnhtIcxKwTNqhwLzccF40vq
L1YkhJs8WPOzm24LsWFSz3q7vrl9JnjVcm5w69RhGJBr67Zs6z3g5YW6D1fdFcQUju8tUgKtAm68
Lv607E4X29Qz5wORnyyxlQNNDnHbSqnHsc571f3fdv2NL/E+49UYGC7tT19UOp7kQgiBk3exs/jN
5nl1reyjXl+QuK5QvIeSJHpyYuklamQC4YqzbYW/pA7WU4FO1i8rOP47ycYH/r7C/dPLfLOSqpz7
+xIZxbJ1IjAm+/o433wZKndjzHSrP/gJSyrfYJ+6AhJ9oFVRWG2kbqwDkileN0hDEo9Uulj6CSPf
EIf7Q0Us9z3Zn+EQAL6k6hOpdW/3AyJcew6JCLpYsGX4nbjlYaHUDV7Qjlsw77eHCYgoUQ1iIoxF
OqwUYq5VBfxmDsjFszcXHUz0GoejF0DOncWN7On+/Y1vj+LGH+Akbvl7LV0g9RIj4CUIRKawe/oa
B/PLxOpZ3K1FmlnhdWeCPIT2GUtU1CpHAM5xpzDh9zpVMF6pjBcijdJiCufYRxL+MmqXelwhWH3V
KKiIVwXLPp3wNNE0joqXfsEf12jddrIgEkQV0yswQgHiKL3e2GjEBG+u+fvgeMJHdrF58EUiI4AA
tVlMXZErrMyEpIT7hH1LTUX+8dpzy0J3wiSNwf9sCfhN0P4QOPEffVUAvD9E8pw8zWe+7M1Ayel9
cgSgn6wpuWr/CyrsnhwTZZe3UWdfE1udY7QFINJkgkmie7PiXlXoj6iQSu4zUQLGkvgcAmtIoeTu
o6Pry+JMqCuGOHk14Yd09ZFhBx7Wwew/mqzAXho9uBRIn6ghBPF8ojnEvdS2zhsKofbzefGoEg4w
dD/vQFmvBtvjZNuwIZ9WLl9sOLJiYNTGK/EPoZxhwN1FKUuLY1m+VUcnp2jppVWLltDdYkqvL8PR
jpDHtpJdrRKuBUldXmNvLUfhNoVQp6S4BpoSWS5BKqLpl3pLAO42vAlEEvnnC0wrtJrvPLLoGdLF
wqmoOQeOS3vKhZh4brbKwsYhLItbjrnGlPuX8ksLXRS+EHbBxJDYT/7uQ/xGAkyPYAmSdOFohr33
QD6JblTBknIrSlKykSsaGvpA5kjUdH4oEAh2SdqmFY/sWwhaCGXZC82vM3c42979On1bJvEZzDqg
2aTll2HwkyLK9a1Cd+ABL9WbaxzbD4pfvW4gms5iUdn5QO3YRGjFHA9Ku3HJoFrLCFsvRrgqhn2a
qQAn5Ycln1lBvftdDRIGboclk59rzKQU6PqApj7G54BBgESvEvyPfHT4rpthY5FDVjDo9nTY0rOe
1SgJc3naoXTKW/Fv0RYY8zalZd0BwmUSMmQDZhtQYcSzI831X/gdiA88Wusfqc7Kpwn2Sr2XkDBg
Q6yICgy1yImlDr3xn4PEn59plJs7l/OB6NpuykJ/Hai9VYiJMHU2tQUSYp/NAcwqSgfX7Ag8vj1E
X8zpvUMtofa4AcDClhXwiqHKZODU/0NHvejxq3V4eQdvWXEjdG7+EY8xhSRgqsz0jzb+7Fq/COVr
tYBPVQqQBerek/oHRipvY5CaRDCm5Luzs9AG36btVmWVmAfWq5wohLHVn0wzhkU2wvd9AesdeV8Q
fj24iAoE6uNvYoCZesNImvz3EaakNqEAL0+HMpq63oQ42vvii5/YMGvosvlz4EvAGJdGAOgEMjxt
Yp7mriBemJEzzeN2pMjUQItKHxrido2TBoMgMIPTteE0AgpQFSf3JOHbJkPC8JX9iKP5mXTbXMas
MGTEU91zF+3DYevLdHYvyNGcoiizF+/UgjRsrVp4PLJIq+Rz6aFuli6+gjE0yN7kwjlIDjsh5nZN
CZ3dNA52agrf2/z2QGMG06oTRHxiTcQWxCWPpe+yUS3mJ0bURAe51/eCDFd1oJGUCpyosbhIgrdB
MY5CTLu0pXJGul+zJC/NnVPP/w4doGRrF2w02k3djgDJYhRo4UmoqLa8vHER+g35u+hC9v9obHN4
ad1lvTOYdmwRuzP7C4vZMSTNqdOCi2auLDgRAQouH+AbhKG598DkT9h/8YOjOXB225skbhqvyPYW
Fp3zhXlwAgufmVZoBkn0eXqyHgvxAH++yBny10nNZOZspLPynbUgCeJ3Z9Sj4dONUUB+Uf+GkTy+
OQL7eI+GG1tqvvLZJGL2gcgatOEjaOQGP3vcEFeFTRQg5ZZXP6V0ZJsjKL/rdl1bAIx0uzu+aPTd
ETUryOLUHHgbY3lzpG6TqwJ8ef875nOVcn+ayOYaYlLBAWS0EkcXNE+fOeUSpPBRbOfftPKo6uck
2fDOGzU49x25gB0AjxQoz7PJmLPDx/l90dbWwDI+0f8cDCgvFuKqP6HsoGdmyO1U+dt/RdxT1WXH
Zx7RhgegJQ1Mr034Z7Qb7Qzq9A4igLyQzECS29OcCSdg8udYSr3xxCODCgIx909HYXTPdv4hpQ9z
ltE7UEQWgczh6Bo410uP2dDQpnu1Nqlwe8bJ8pUc6+ref6GsRT/tja5WGuwLHjh79+nnZH3nZWH0
f4VlVoRE7573/oqR07TFeR77UyVlYCjPzO1mkIYhSW9bohLZ1nIcvAaNUTJpelOkIX4bM11X8Qy5
Z3NiS87Ccwo1StUD04UvIILZ4Sxt0yNEhXFp6dyk6LN89tPRLJiL8PWqLk98R4vmLD1xon3IqgZG
UgWBWEjKgg+zLW4vSNxmx6TwqMuusbPsD69TpFRagUD7DQjsSlVUiqLyGZowlUxUjKheCU1V5aff
KuwXuSyhGs2NOs+hkeMduDn7SGA2Tz6ehQAYTRoJviQUOWSPTG/WUuj5T/IeYa/ML+kS5o8xjyH6
4B3zH4cmy7pMJaJ9IjkNvTBVldaLn8K48uVRGO6JoUonFZvN8q02xUEHlIY79x1WVFEvRma2F7aa
pRxwOVutCZgFrDLqoqaizekPdiesCKXWFSDMg454cca8Ry4efLWLVtYSEn2so9/2Dj6pxS5n/HG6
BuiuwhEoSZSqRZ+aTltoz+DKko1EMUG6VCvyi5kNbeVPf1AHQO1WqjJYYCdrDzyZgVBMpxmIEOCo
aF6NtS9gniJMvZnx1yCtONitsG2D8DoeYw1+Ihtq3IucEngAtaLfZ1QM4NDz3WoZerMMXz71ebUy
d8xPerXOwylGYiyhIz92Ixk5Uo0gz5WW9Cr84ANBjPmgl6ipIhMfUXawTeEwZIPiyMNgFvZvwkxh
y5XeDj/3z/sflmEhWN4trcMbWaSaLh5aCC2A7DsNNqdTJeFAPGzaTt+b21M/H9spD9c3J6pWHrav
sK3jCMwW7JujRln6guH/EznOyMtHiwXvzls5ImGLrvHsxNy93flZ0ftHltv+ZzztNlf2XEQzu9jP
WhtBCjNR9IxIp+ukkBeAezqfcQJKLn/yGFoLcTaMyRMvcIHH25+7iUyLf258czu1ON3RNtNg7LHm
inwEX+MMYT6wgK7iX7VGGuAc/fmcGOSm9AQQUM+bbpP9qJIeTMSO4U2TAG1OgUBqUOsgJMWd5T4A
1fux/uThi/W2z5cWNdU/WGOwvEBTVYeNyYQlOwNOtRqHmuE3JKqRvgiRNbYhncA/nBY6o1GDwC2g
osHG2q6U9+HOVAZqftGgfLjcOds4oqkIhewsTUTE0wSwZdwnCzVtyXfXXlTdlH4vEbyoskL53R+n
ncPxUhfMUBEHAjp7hKmgP/TOG+CBc92yLjMWXLtXzY/wsxnnUunY8lkmwB/PcoaEK6N6wjBdOmcW
y06GpvxT8LGLbyFBR3GmX8Ux3KJKuvJkhyYJNkCNoDS3ZF6URf1OiFxGhCqDqKDY19TnWw0NefOq
uSVput1kHhdWqJrUl9aInMQyKScpjZuRLbVsOOXYjYxXmeH81RAwSyGxv8b+ARh2pzc72KcyDPKN
dqq+3wqQuaLlPPTHjeI+OvC5cMSVsyDaMUqkmqiv/J9pbNs1/fz+Lku3sM94GSBClZVw42kL5p2w
0hDZ//BoSUKMU9D2Po96K08FT/5XJuEibb+bhqh+wFVK/6oh4gHaKn4Mwyg0e1zxnkXzb5S5dOCn
X1dVOQ+eWev1dsq4KOLQX95ffuqu8wItE3/CeUYEXnmB5GASPiE/8OxWLjgIbVF5FkafJb5g8rcw
emI6TyEb1dZOAuox5f0dWqP3xDoYabysfySWXCQQRNASnJ3yUswdmDP67YB7o0A0j8ScTsedE5U9
ZVr1cZ3uxu6QaZllAEithRGYkFOpMRTrDEsdoJw+p+S/AsaVQUyVgr+/ZooadVFZC09uUQp0j+2n
3G7tRcQuewx7ksE7f7yyrGnbOK6E6Ax8GHJngPld+gs24/rRVrj+9UuuLFUZkHsjmXHtDZMwRTJw
YK6LuyU6Z/NziKiCGK6CsmUbISiZR09c9CpaQZiSvsokRXZscI0tssVPfMntSf1YMVZf1+GNSBJ7
y5kbozpayy4Cf+VTPX5v8dadnztNpqXrluGDj5LAxc6sSRkgiHPCfzFfTiiUmbyqu1p3m6zPtZYN
GXlxGADulrtDiuaNWojl7uliepvngfaOjLWJJ9Oxcai5FCPiRBz0wzJc/bGfc3ArgY/GXNCGEJb1
8cmkerDTtETN+WWYo3M4xpMO7P6RjrDaq8OLnbNVXMMuszLQSth5iD1d5YiYE24zD1F2Ih2m6mto
eYAkV5PhpbZO2X41iVEDRbqAFbJrAUu5UrDR92Ms3IWFKKO6rw64fQ1JCn1qB+D5jMhVh0zH9Tzh
yt39aYymsZQQwsmn/ui4GGTqS0ZMvkiaA9Z8u0YgEf1LJAzJzPnP46LqZ0qcY7gcHF9Tj4VUC9RY
4r2SeMDBZAdhTvTV7Nj5b/FRa9e3EvOQ1Fm1hFXcTp8mEW29xvj2F1uZ2GkOrSmr7FvzmuBCEOqj
WrgjwWk1LV1xXcO6sUkXDk1/4VvFckx05/TpCYJ06UX9oi48I/BnePdYKjiIJG2TjULgr4tTAPgm
5/xAG/EcwKWzNDcroWND5gY0kJ29B2D8oSgzHPr9Nddq1f3hoIR7a3Wxp/AdxXblQFUdizhlthfK
YUlMAHnJAVIWBLQkp36qe0GIbkMJY11xaI1aXfaLK6W36M3+dGL3gaNzoaRwf6RaY1oM5Hx90Ntt
19nxMY6C5uvNHKrG6XoDDh/+yjWDAAXVUX9jNxtt2tBKnReoTOLWaafMwakO8rcWR6e2EN32qYIP
J1z69kMEtge1OBsv0oSdjUZMArVISymB0r7UwOce2/JsTZKU6y3STZP01MCUVKEWe/6UMLECMN0s
hIq8KehwQLNBp7NZ6wIAQt1htopVnTqTt5a0jzxNDZcRjCyqSQRSd5WMchnwmDSPfqZlhfTAKm9c
jz7/PWzo311n0qSacg7/qdumpoSitJsdSUzLkYlaGBhKbd/S9qy+IFBr1pT/dWfpValNx410ftdN
ikOvUpFj0bm7dKVfSc1YwArqtDRtUoWm6H3imaOr5QpZHIij+Ecv7eA6Z23lXxstsIaNgBfD5t9t
cQBhoMey1MkN/aUY1nyAsYbFHNsCi6sg1TnWvl38Jp29XIeM/tzJtCRdUGlB472PEzrnwyRi3v9j
Bnn/hiHNpXHO8+GOX+5XO1N8aAo5hp3gbHr+B1hD2xwwFK32rTllue60NtSat4TDY2fTTwsOCIMd
iX+FAB444e6yoHVmZ0keGSP8ovEEEwqdIevnFBnpcWIces7uq3q1HOMymAiHkDsehZc37rzhNlPm
IZlVnk8KcsK81KTz7indfZfPL08Wq383VC78jHWCkCh/3wvWicWZLS+kWF5MKCabdUu27W+JNGsC
1yQSJwGcrjYlEDXdHYtKb0nqAil1jFvr+OarOScxi3VtpLaJHQmeccLXwLp1Vh66S5PWt5xpJBqL
set/bIXIZtYtGStuUCnAZOus0BHObxzc30noPKrGLfzIF74duFSNcuUwS1zHUcXsebrIUYefF5wZ
vtvSNsicFldUwcoDCkAW78kpkwhX+uBfkPkx5dbpJnIKGCNxiZEB0mX+1L+zRx9YyYa9l89H8qST
3XejA8qG61335RylBKWUuz83uJOP3Oo4/TsTJvpGA+YSSTJdPGEEAaJuF7XKt+Iq1RqYQXiSprYL
o/RcoZ60LyLpxwvjsL12jhfhIO98oMKfw9edkJRTPYxhq74EsR2gplYa5vWzaiIf/gN3A+2/+ZnZ
K88jCg5D7ZtksAec1qL+1BPwlPakxbA+ik6YBfoN8nD5c0Vk/oy1VAkxVZM4A04pZOHuvTPB/FWA
7zG9BdIFInylpqcPslgz7lU5ZwEvcploxAxA0XVJB5U/+S7eerp58e7enWflVL+RaCjsXJL+9jfY
M6uxed/hZbomXuWVOjV5xm8brkhxutt6Vye4voOGOBHa62TRk52YnzHWt6w4dFgfrTHLXPJhDPm9
y6y1lsBhB6HMolJbsv80jK6EzHEnLTK9EZzAYXzewxj7WGau7lFm0EPSbHkxwp/2lBxlBsy81I3N
iT+ejoMBtRKgkAh65dr8YpkHjYTRqoxYotrQsSBzOMg9xo4clc0M49fFYZKLdQazBlON2gbPu51D
pneVDm5/JGZdK1ltnGkg0dW7h7woktLr2ls0XARb5LENFJzzNsMIFEFn+enxM/7N8T5Z1ccR1XoD
vbYfTX2cqheMTPlcaGw0QFnn5tvL5Jf4Nsn5bMSA3GM/2lMbeVCn5VaJJ3XsrhIg+pIgwxOlN/yL
T3mSm2tLjHqDM6h+eDBiV9W9g5IY7Z4kg+zxKX00KGqvchTBl8zx0QHRlgkU/7psE9j/m3wt4EG5
aih0U7PNF5cB+Pfv/IXr9FiY8wuU0ljlhRFP5c3KeQfMvh5YWMVIWLYLODi+RBKVo6XVNqYyqlYL
+YzCZWmsTpMcreLerv8+JbQLebuIY7QLvA5CNc7X00mDQp9pQJbAQgSGT+j8hByGWyBJ3NdbFIHQ
cX8c5TOKst2yVGJrdNAnWVorDWr+aei0qeKBSnp6g2c5N7uCxRP5PNZarjAimGbbhFCrQ4mvc5mb
hp6pG95iakZSW2N8/n6DWGRBqe7LcZ0g90iS0+KNm0WGMMQtTgnwxHNnuUYNg3jngskxw7ncNtGk
eFwB0U/67DdEirVltGH8wkv3Ozuq7OqXsstDVFgYHu1q3VWi+6+GOAhW1qYfXJNX3upw343COnN1
n31aConwFmdaDUbn2bVwP9BN1Cbi9R8cJl5FQq6grZ7IiFfxPZ1IiHkidPi9Bwt38yzIrxFb8+0S
3bhtRP5Iys5GW0kh88HILEwzeqSR37AG06y5czq5t/m/k7PilOlCkEMAA0Y3IN9Lx9g8tbGUShpI
lQ/tM9dY5LKniGHaGMK8BIuQvgLIdf0+jaX8btERchwlC0O16saF4bdUyLur7GVUV02uFYT6kBp+
4A6XoXMtuiOMRKMpVwL5umnsqircB4wDHY5Je/0NFiXi2Snqq9pvwjdTMnS2D8B8j+Np12L7UJxi
UxL7UfQtxQEX6wIfCn983wGwfZJVDNe1kZaMYJmzL8pT3QxBGKxcFN3VVdmr9eEUfGu55jwzixSW
CRRxkvZaXsKRnMXsU/qGzXtASl26N9p8YaSKrbfohXqxlH++wOPUX71Iu1O8IbrwrPWSol1YwIjk
C7B/M3XTo8/kGqwkw7T4R3octbuB2LHRpvAl5G0QzTl4TxaiCTzwbfc4krVDFoGeR8EEyCn/d8F0
2K65ioi6u/ZppU9NgeHUzRrcpfFFIWNYJHT9fVGOtaotSOerkSlyq3RgwGfRXrQnj/1IaWvXLpq2
TNZSmsulecfCJqvOkhN1v3vXMstTUVUOEQ6MuK/Qfsf1X4k849Bimr4HurNZFy/dVPZOSwElFug3
uh/O+xyqJIFy2+2mC3LdgtrLCxZ0NOewUx8DgUv5smm3Td5Pw6z6iSIKUm4d6Ph4aJDhXfvMKe6X
P3QthKeUXzFHIyRWNcgX1jVBlNnmVYE3XExHQ1ZgcfFex9bopMjrKwVGXJ6mjMf8u69IleaDYSsn
i6KawRh9p20YGw1PyOxw68C1gLH9yfR21IGM/Au2wIkveBLcYzIo0HQbhZdA+rjfF8qMPfu1JE2j
Mh73aq6q5tJiERS+fs6JsLD3v3QiTgHBDRpj8VLGi5+zY9FVeeCkLeWx5cyk53U7EWl4umf51RIi
czaHPX5erS4N57vUWApIT0xuoYF7arRdbLRR5INEXPZSByYxA9m6EV7Kr05mGuv2Q5N5rpZAtXcZ
NioZKO4Iased8dnVXgf2PriOe564tXGp+zZ4AfG0wZSHFvW+X13araVP0eiNwGcqKuWSOK733SKt
LwVyl+xWDb1ULInDxBgZfEX4Q+pkjLn2HU8u1raIIjlZ9E9ug6BP84AwTtDN9thi0gQuL6iD97IR
0+e7jNJxKBp7gB67KaCXGgyPO/FBtLXrh4Kp88MCalBxDTdUClonCKuKHPpqRD12C5XcZ+EC+6dU
TVkmJ/Rt0R4e1HFXNm5Uq3gNQZ8EXOGBW92ZBapG390+dq7UWygzDHDSa2XDquT7SCY8FkendmhE
rSuUsk1TpCi6ZTDF+u8zZFN1P3oWZ6v77uO4fvQzv8blBejyVmq+0LhrA4Hn9+2ml8WNY5JfIu+Z
WwjTgeIBzs5UH2c3Ci9IdFePS8Tk8aji/stReo75S1oWLKe3ZAdPzWbLX1L9HNW/63rAVBIrutEv
9aN/5HgE0SHGqTGuIMagKyuZ51AlbkKc3Zfxh1z+CLqY4fQ8tCzQjFoompPCotobhNnrZMQa09py
/owoDcxPRio+hAQuFyVB+KQeDtdUgBTqCOBH3AAhvKQvn/HvhfzozHsrukP5DDN3ZrQ8Er54AXev
atZMFkfN4T3gTdb3Z+xdY9WPGalxAamfvjozb8dTC9OY3YJvruOQG+CSZrBX6saOymsOdXUx5lbs
DwKqfp9DXtaDTHBcVzrz0MI8IxMernvT8Ka+ZkBBf7x4LbChg+DCwfYf9aJZ2dJy4JL2YWshdNaN
bGAnnJD4MnKH19A1v0w1xTYYecQSNzl1ecl6DEVKyvEIytm7UBijgzuYaizW4DD02vM0/vNQ/kvW
FZ9Ztlczaw4InGR7vBpktc6g2SjIEHeUMEOnBZ7eiVKalV54HZ7fhMLiNDXrjIw8yPHP1B+QBl1Z
vT8SiDmxolGaP1PtsWpVYAkEyehvFTV7zKyAK3UOEtUvrKulnwpDwHIf2gH1tPOWlbMX48e1YbNx
FXpa8iZUQZrWaMD9pN16api4BCoWgwWIBimfEI1UDFmIDq52MJLMKdDYSuWOk/vLH5JhGPG95uRn
qHwxFBnl0a2oXv7sukO2EvZW9FLzmBjKx62weOztztEEJymrzrwesrZRfmzrog/69WpuMgLUeqex
J6v4OzqpPQjtwYqlgc+Z2eGdxtrIBH5xpgvgpxaf4W9DUjTyDR3wpmDWZiFfYHN6MHcQqqfvJ4TU
qDzG6zYLJn1m6cH61tQtBMb2iAoC47F0+g7/055Xzul45EZmS9wLLObuMx1TGaraK/FD6rD1WHoa
XznK5OdUume1JKxzFFKPsnPByyYOT5BG0M9woiXoCxbr1KrqY43aAhtUwBq7hOgX0O5tl4ZmCAAJ
wBqa9+KzFZ2w+kdGNIGWGQxyJplFbbUHF12hgxITxFlJ/gRu90sS1mbxNesNjirmM+axmYICtc06
VVdB6CfMK60dlWBx1ccVRg8R/sabNYQytfHK8N5RvdLkCEWzsuc/JEPNvzUVgBvZbVb8srtBSZ+n
tahxy5R2FK1z2YR9clYgOfp2f72xPZdKLN9exQi2fn0xx5xVGcUwf44htZpfGKOXHpk54Semvbw8
EbjatxoS3ScMD+DK9peTQEGPZFBT88zAD/zowh/zisHmlo376GAHuZNyihbv1lVu1AYHfb5vIXn5
8vn5DiowRA162kOiXUuP6gkGMf8yrNSk5ZKc0tgWaZPMhAghIa7aydKqCad7k53ZaBhytxD1O5xt
a6Uw6gM8y2X8dvGoxdFNvOaZ/DlVKYBQljHc0Sxk/yazonrTBQqeTHRw1XBaR1ew85w844S6Sdab
cmXsOar2zlNFZgfKMVs1ThABpnS2ByANAiDHK66yIktB1+IgHLEGhY3LNLdwaGnOf9pzjZUC028b
ZNxGhBt9HeiPTumThXrtIdchRkuY1xEVBZKWXF+Uag82HQRX63SvkRARF5RKZlWbXbzFj4Y+19/i
2ctFuhaPjGvuxI7Fl9PO82Ig1lz/Tj943kp5j+V6HpXwBWQWfh0BqgDz9BVRgAGnSNv2VbnPn2Xw
9HQx/9Pq6uOvNhiNQ3e5CemfjjJW2x8oMVPGm2wBugZHvM59n8m79ywJyZrdtPb0ZkgjEmedUjBY
k0rhmJfX3CwPs+Z8+U0/sncObWT6bJ9yF5hai+IP/E7wYx9N7nRQu50+6vdDswAStnmgwO0ddJxY
uylS3OOoGbEn+GPqzzRiyKB8yJ+fF0ToRfMYSmOdmpD0ETIrzg+OOsU/0JEs0vTOQzEL8yxbCEjG
yufmjHoFu4QpdP/saWang1oEklYqzPA2TMymd/rEysSRHtQFVVXbHvgHdZQiPz0YKflz5RlLEfAQ
sxmYikLjmFiJCCFaF5d76Go/s5YCq5PdBSd5NHC/pPz90GNhOJVuaMUUwn98adQJqyme0PhxErjh
OXzlKfoLG4VTZN2428fFcVHvuHRgGRI8kRmPN2c3xHkWxtHKTaQJggYW8+1x8P35I92lAlw46oy4
6aAHDxHGw8IDkOsYj5yWFAa4kJHOjgYt0FJwY/E/oTdEaD7OOQdnGRIubN9GoA25vSQJRmXfikE5
Ba6mLZ208iPiC7a8b0LKTqlWoS/oXeZSZD6euFG0uHbiy7MFsh++HXcH+i0qfDmypbtlDz7DWUfC
E4XiT9JudwU7WJix1xxQXiXi+ma1xBCbY5X5Nk6E8AH+RspSnkD7gvHWgqJE3Rb+R8DzelkudgvI
YGfnS6n7WHckUkR9OINBK+2Q+zyQQgig+Fyh/N9JoN3HeHAUmMJQRfUg53o72f4fePFt/jJvCDwf
DV625Fq01sn5kYNA5pnjCMYrjW+pb8Vufz+J9mBjpGTGxB6j5YjhwNdnz7ay0afy1c6FNklROM75
Nzj0+BXAx80vRzau3Hifo7+2N2ktKdtFGcR1B3dsD/UoQ0wAtOV7uJvle2zchnpfNCcy0u5neKMv
yatLjlYQat2IfNfA/fn40YTIaU824gzz631jKUFytPn/3T+ObGrYISRurKA17Ttl3Wv9IlFGvRGo
gExdNJQZ328spZxi9LcH07Kg6i8onTsz558iTsm00cogYSTRlAqtOqE1LbtqNyIcX9JQ76B5B9Gn
lZ/ehxLBPsJ9jhSxbpwrCqq7T1GyI72Zjt8Cx7SaiT2kt4e9IA7g1U0s8LnQ50NAKAnNPJlkz5WY
F7LpekFa8FhJIqsm3JHeifrB0XVFs7fjS+OfakC21C8Pbfm+ALU+vFiEHEyphE07l87+XvOJYcpg
yCTmAwrSl8qaKvgjm0vxd373vEo1aMhuQ0uQtJwurWK2LLv2CBEThFrF1ZUvy4AKL2Nut7zet/ye
JIVwiexTo91itoIgA3Tx7ZFgKknCnewvNb0GB01efn0bU0K6/GwRYKZmQOdDniOvuOUUUuQRp3Sq
2gRcDBm9LfgWcKJIzkJSI4pBh2m4scuV5T8h+wH3gs7GmCbxa4AGALAdsA8oEWw4I7A/Li9HDj9J
quF5pPBNukqz8uZYL9e0+//67nzVgkrfsWDiuPcKJtLpj5KvuMg6C1oR5TkIBbVZ83TcKBQJ/ONh
RfALX9Liy5j+AkutnJfp+cJiLkkfvrkw9lvP/qrXKXf/hgvrx7126WPEyFcae6mui19KXp2L20io
7VwX4LJBMHmZCrss65Ao0wscPaJkH9IPShi9UxWzjM1Qeuk62M/ZFxiDbxYwg+No7Ml9ruTzJfGg
35Bl3fCjmbhCkgP98wpwOHubtb1qsx1utTCGDgXnOUyHUN1l+6XF+1CwVB8JTiMyJlmxXu+MFXlE
4gLY9RSKbxAEXTqhHnZ/+vn5pRMKz6HYzUnCqg2eD1SZohrYu332LBw2DhBa+vmelgxMpIOQ2wux
8NRarRmbUa0dq/MQ6ke0G7cXZJ3dUg2k+xTYlzQcxduzWg5upGUgjrjaLLpg/XJZ9JZhGTu1e4F7
ewm1REf22AbCpFKEuUNZf3ClAVqPU0LEqoc4CjdBxb4T1GYMgal2Ep0G/pGS/+eX6jL13fQ2CHgi
cfCKQLFfDFDc1R823OnPUCTRsSj9aS3uIeJgY2EnA0oa3E5A5qItfqmw4jxpHF7gWJ6XopAJZT5v
pGpW86u2mb6Vqpdl1epQOPcC09OkQrP9yCBZF8l1fip7IbGvf5gHuRynZnyF82FgNwsbMgwaUki6
/F9JdFm+MzeDfDw/Ep+bfRrmTabnwTClJj/61+pfLtJA72hmJ+CK3g3TuTlBqCiyBnwObtn28rSL
9bgae9fe/uXqvpsU4j1yUoPjaFaNRDKnWTFGHF8q8/NoUQL4aSnQ1/uE6yE0AkxlB2AzXVtZtNUU
zMh+Jz41bdILOpUaQJENEz647WrCd/LIQkyOpafaEQH6xm0Q2VelACAFlJxMUkggR/uvqQc4zunW
iTQe7rTc/tqntM2bklJInJCa7wF29kqGTNBQArQVpKSiZmV8K2yQxniAC0WYjaeTJ+p4hqOPBHOC
cC8ChTV6Ch9K5wqSR8GIcMJhvqKLwA30O8yUSs3JCqRcbCy10ptCraVf/f2Ymx2wzxfh8pqcOfki
Bf9fEc6wCS7xb7T2KZNyNCqr2x/hRwtY5lZ1ygQvDnSmz3ErO7FULMq9AN8x6ejJ+kQIN8hBH0jO
cItoOFeBqNFqFQTLHiGrv9QB0X+XNxQqHDlOMVxWIXCafYox2+IUiZd1YGWoyGgr97HghroiFZit
d4j36vmVaz7rXZXqZe1X1RPdaDnHg6DcRmJVXKLlZDPIP/dzWLDc1FeG5sereY7Gty8hr2STeeBJ
hQO0KRh7LuWWokjluLWfzXsfqrBNjT4kF9zTbTvpCIeIim/P8ZQA1jR48UWBCSxR4LQ7Be8SbY73
UMkzRl5qJiqnz231ScQAn5lJq22pOm9H01Wyl/RTHU2GfVMQQ49RZPTnE736UbWo74B4RO8msTsE
XPIURwGOlJG65WT5K0+kK6PFT3dqKGdn+vDbCoM5YqbrJjZHGAt3cP/Y/ZiRI9jKqkEF579BKqkF
m53h4rxhB1I+NMbvWE5MfRupTkJXhjlZA/HNyNMHM45q8XM/9KWzakf28ulugsYQ1vNfpuih8Yf+
QjRfVRpybFsdqAHY5kt1NBIOetxcpWDsY9gXuIEKBv6NVWFgUA7KDQ4q847H22wtMnCrOHQ1l2Su
HqGks5YEevA74NOe9Y6altLDo3fmO7Bi0IDfdRzKpD/gBEGHer7Z/MxUfDPZZ9AeagRpLPfGrjTF
yISyPCWxlhPaYeLQjumHIiGkIbHv1QgHN1tQsDUkBd5mLvLEjKN7QSFgy7SOG9n9vBDGC9ddf0mp
o7eGj/JBNYe3WKIzF0LbhBi7qUuEHLlkFOImUJRYYhiaaXHZ1CZD99oM+wX9waFmAlr7fz3/4v7T
NHj3VgQHq41MpEi7GQSwLwH8wxChZVt8GCNqu4FKHE616TSQeqZb5QP2X9DYptvY8n1qq5Z+FRB5
MbXWYMC1Q1v+2ubnx8VMmvpkRaNapH/smwpz4IIRLif0ZoaRWlf7KgLxHeZz1EUm+bqhmQfVPuCJ
ok2raVKvQZ8GYV4VQFy/+xjxec3/HVq1Jnu5u/0O2h6j6ed7ccSUFI7FW0ATXdlnL/o6yt8b+qlY
BULRAhhKSw/ThriNtHHnvmqrZ2QGsSy3aB+UI7kqWNM2yEGM281ees7Cx8lFzqGRau9PKhXEoIYC
Dmd0E7UKk62mvVJ+Bw63BJdmi/E5D0IdfLPUB/DGbj1VZyfmFDOze0ZI2+JuWxkIrnLhaGrVjH2n
8GcyQF+17TWgTYyXzWxDRngKA7mUYaQSn5Xlt3w0XhE99xhbtUh/nKoh77/chRwT/pkgQCqK9om7
Objvw8UyX7jF4Alw+2n+gCjL6T43RaTETuO5kcwGXobQ0NEBJ2BAExc0QMM1APGbj29sUYqvysbD
+UllsfOiHaGgFyKGS4yoHDyR42P8ud5HyolEyH8WCExAnHwWLnCv0Ho4i9DKjnGMMHymd7Ld6EZR
I6f9BZk4CoVHk3ukuhaDTF7g1iuGHp2nhqcqHu80Sa70QDz4OEfBOlflgH/cV5oBcuseXNNeahKm
98xgmOemVKDZ/bLUBa7t90iDEGebQQAYCKnpUYedNxPH5UFBIEkYLEIEFbA6byu2LjX1OltGyUrV
TClaet4sATj39FNuL2G+MkLwLtP2QOpwIFlnE/pZBV/ZrcQoFgz/NyGIMUqoSLgyZuodK8Cql0nU
nw4Rl02+cG6Ijj/IlPDtyW38HSvdxWeL6Q8AOaI0zPEcxqC8cvNyOxJN8oNO9w6duitAESzi8AJx
r/ARTgXZb0mFcPor8LoyVVa9LnfxFIp3RZNp6VbdWQxwll0EqWl5+7u3iBgdqaJW4h6fiUIwn8ju
BZW0T/gEbqCBLJk573hvwnIDFNQeSWCDpWPf01okecshKO/dhIAdLhIJAb/NQKXuCXq5ieuul8mP
dCWMvVMb4j2JZjjFY0ZpscQSFKwfDzhZxUr1SqG4mctP2HsUFFwV/hYsAGyDqRfGg/iiBP4Ua+3f
MaIt9Lf88kfsHo/k3IisVMcFVHYIgOPumThLtY8Pp9o7a+7Dc8d6EFpbwl7AIOW0Y7XST1A1e2Vv
B6i2SIS4mObF/dqQO+FSA5hbjCXh28hF0HkbW0R/sorWz7NncSSYloQfiSRVXe20b8bciOf8y3Nb
ctDsTslhY8Z2LBeWbvvmBBlDkN59ig+gRtRD0y9+7MzRyo7+ZdEZ5gwVZ+x074ogWYIM1lih6aEb
csxlmzsHAuVsn4LL4ClYxY6t+a6bSLn9U1lZ/MBeukdss5HeVu2ptJrZYmwThHt3nCxrrvUk2A3V
lapPtBdRWWnFEzn33esk0X0EaOhZTg/RDVmNqJPqYkCVqeSDth0DHXqh/4EzblVIDvFuBbar8ejS
XLwnTOywPHeE+HE2qxUX38oyzDYoC9eI22CcbLUCuG7ufGUPQBp8Pu5ayZri+DdNXza+ZbVZH/11
Crzjq+1TTSjo+6U57G3JkKDmKW2XRaDArjsyAb1fhg8tTqJweygfmRIP+5FiOnfMsws/itW53cru
X9joNBtSAUkG4tKmV95No6xtkkufIH910DWJ5PcjWD/Gm5sLVR+dx9V5SZ0BUzc9stQ+YSowAVo5
YaKhplRvT1662d+LZq0WejS3cmGVQhoxLCmOCTW5KMfZv8MDSdCrTwQnLTXh2CZsiJHvYjqu6fcP
d/P+BXXNEeWGMD40RJZtMamppGPDxIAFvQF+bINrjEzgpgXUzvv2XpsMtCohJvx7Kow0vQT8jIgE
5BdfbtPhMpt0NIv0uqk8TZoEtUF2jxJSqp+mCsxETPCwoBZ+hiV1wsN7npG/v6duGaApF8s8JGFo
yAgOoI4BkI9kAxVdQi8Bx2A57gQf8/bT42DxGSq1Jk89l3NaM1RMauGtyz/hYSTW+EYbs7dB/l1E
Udj68jHjzjiXVMVGsXB3SjE54TWX2tNPGAa8rv+lPCUQfrXQAtrD48zwdIzjZzQr1T/VLX7N4pv/
3OAg+JzOvCm4j/GO+TQ9fDqv7B1de/nxXSrS29L4uXvdXkp9vp7x2EWU+ldGe7Xcg0cCoA5ZT7VH
TGixICFXTaBVgRMBnPJe/P+dBWb2+jrOVWtQxuDxoOMfilB4iW6L88aoHwdeabEli0jQlykKnULY
SIXEIDn3MgXKBtapjtD17BpvaBMgCP20t57Wh3N2iNbhCMtbSMpNEFp9yCSzUH2mCG4xZYFS1gbV
wTgA3qZ1sAFLhIZ7vwyKhjXJ0kL8boNKnsm+lPyFvu3BYx7P9akjFxkdjH2dTS8oFhhp0R5ddxIk
lt2La2KnKfKkn8DZOIAU4NMaium5MSqf49F+gXjGPmeVA/8OdennGVkQk9LTqV4QmYmMAtiPbl7Z
5WS6B5yYTZDyO7yAeRSAg3PWa6DlRX6hiUSrMFU5FycuaAwA9DeJe7S/dqxXo1Lw3f8LqFQO8TTg
j64Yc9rjtZ4ejRWqxEfaQ+fGZ+txmr5YFuRgIzQ1wP1awL14cpbt20YZ76glHBz21VW7ch2suxUj
yp4QYMN1lkwQ47a+5v6x+S1Ew8Z2dSlo/kmtIF7i2Jc6TY5WNqgjhgSNuJYXeqbofyqzd1ySS3ow
hmxT+RyMtSQ4Y+o0GYYBRNGCkdCribiyv5C1iPyHj3TOiQ6VzZA2mqbwxxIGszZ54YQRVwmFqLvL
0lutYS8m2d04PzzHnjdA9y0G+bS8bRBnyRWj2lHiwWwKmQMllrKe+OI7eA63i+EcF7bbwGzs7ggM
pqxgURvDLZBlpLuFMK9D5DzbypBRvIaIauVajUrrCa7aMO0JpLEn55IKcfIplQ85m+xAZTPSv4wZ
rLBtalCcELGcJa79gdK3eT2zGhvyJiWLHm+zWT/FLRv/BClpGjsoLm5ckHOo3q88Td2HgPMxmem9
IjRWalPH/n3/M0FT3X9trxqs1SkoqfzjnylPrL6iEbWiRhFOvmJcNKzyX1gT0511RxxG1jvd/bTd
c0ZpM9a1CS4sVBnq+ObMwPaPgtjCnGJknbU+unVodXc3bTXCRQXKedT5jzTxLo+zbsWjn40m/6pE
09Tvg85IX3c+3Yk6f5EJIG/Pr7vQBYYj0/iHKk1s3OhSb//6khXgSqrG8fyFEJTEYzb9tRb3hEWA
9+ttZ8Kll8/YmM4fHIlflzLsHuZROcNwpHczCHYQ4C5m0sk4E9VpJm0a77IEDykDFR8CW67zFvO/
gQ/rqAKF3htUOsbHcS/Xvu1YakSbGsFYtsdOkXAxUq5W/dY5Cg9JbL70l5IokJ39eU4rI1IUvz67
SxsP4il2l0X2EMOpFwvzHowpymUxv4opyE+8SuOCvw6nDyr1cCDul5Qw/iXfYdAE2fNBOk8CwpE/
V8OLh82B3ZTAPTV1f0YI/suBSLKxXY8uGhdgYgG4VqtE46cIeovTGg1UlvAfhQf21Z4TqphKSmNd
qcFiqRy49FAM2SJzOwqakZhdYVqyfgJlSfMP9LULiN4bz68HJwhXuhkodZLIGJene4JdLU5IA3CM
tO0sE6Mc5r+R4FgFcZzAQWITtt5coDxMeSDmEGVQgJpho5nujb/sg5oO/VOPng3jvPUXijVZpZEX
kIOYdAvH12HONF95r2TVbm/Q0ple3Hm1hWWGce/Q3YgB+9JZEg45zFuGvBfE2K2Fag06I1JJjXN+
UaP81loTIgHwhTaxMiMEXz3K5YMtxogzEkKBQnVH4UBnBsYbJTc/9ShVKBC165pFFZFFCjQG8y05
oINEi6+/6ryCDs7ZyriWWabzgT/sJtJfVoNTJAp/NkbBtFEZ3WlNkLqDmgQzvmGgkLIpAN6iy6lw
0L+om389POFaVQqKPTWLOrR3wVrhT6hGjaLCAvBI0/JpolCCEtfVMwT6MV56Ga7FyVic8hbHd8eS
3PS0NdxbsUVWr1sH0/A1OtqtToiNA65/g9gVk8aMOJ2lHy8A7m2lE/sSVc6y169lhAMwwKlp3BGf
Fd4k6ixzOsV1OcrvJ2jfZRINQg8daHufgpwgln4T+yvAJh7zEM/KJkW0REdPrRE67kI47qLQaVGd
E4n9Fywzl8/dn/pHWlMepam6S4c7Ps3Wy9l2m8SOM9BHzEeXRnH12s9XFB0anzqo7HjAqhB7wiTV
0lZqJHbFqwXV6V9vO9dEZQ9WFWwRhdPs/16z2rWZK4ILZcGGD5opqhucblw4SiddG3Mq2ndyyB2f
L17r3CCLJb5/GeTCgaC/21KPomPOaw11iMSCDzF+NoFheLKpCVdtpMaD0gNnspXD7ZxdiV9NWz2I
NhCckR4hZ0mejJSICofnbQOtbLw+zwDo4HucbxttOJhuR+6gSm96f3ZFemz6yyIEyCnXt69gKByH
gs55U8OpAviPPZaM/iuNcH0Ir3tFJnDNPzUIBL2tZSnjoZ5Vv2YX0ktRaML0NoK/5Upd/DmbJzT+
duAcJtLJM+5RLPcJ74VYgLrhHG3rOKyLbCUddmQoZBPL9oYs1biljYWv2Z1El3C4D9Ro54y64VFI
uUQy8BrKz7g6tYVse0rtoudBFRRCyKTcCWF/rtgFfkZmk9x5SHLpr2fUZn35RAC9Lr2D96ljJFu2
uOLlgh7T1WJxWA3MJkaIJlQocsTvkHQHDtQOd5siQyQFoRlNILujg0OEci8FYeow1szytohSFyX9
yFO23wVELE+5RevYMGBXnK7BPrcad90TH7pPFqlbwpCYkEEOwVgYZ/NpSr0VRq6SY5L4G9pk8ImU
VSvfVdNCJlxhwTouZZA1VPOrOsm/WP+M7mGChR2OO3oyGx/hcPUkyMQ+PpWqygw2rYB6fR9btGgK
IQQk8OQ4BNDZrwvkRJyHJZQWRr/wouJ0guA8dV6eOnV8ZDIXFzeK1OyFo07hTS5ruS2nIYzHmYBb
0cmk4ZynjzdZqklCAQK/GfYWSKt51j4dl/5fu74tGc0dHtXjgi2Wybr4a7hPJ0hMpZRl8emkVO4C
LXT64MZLL7lrAkzQ+MqF9AtJ/EnzP6wMcKhYBoQfFbKjHh9BVL4i2hy/rsS4BLHQKAWvZSLjxBDG
6gb3S04yKe2LP1edBhyh79TT+vKU/YtKZCz2sovoPZG+pVgY4+pkg7UXIY6h+1R5zU6qjyUdwh6/
kpw60KB4nlPgNX+09ylcRYGm1t49rARhIrwG3NqIsPVJuNZLunV8gyBQl2agEgd2VXEe1LiXHVHz
lyQMLEHkiyYwOH49LFCdrJVLXEgkRKoKj5DqBnYiVI2v05O5DdORXpJnW6ds2Dt4TwwATK69q9lT
abcthkcl/YZzJc7Iv/ZMFtG+hMidOg5vk+AklDwY2zOCfcd3VYlAssEGx0rXguEnsl64RWqh+1Ht
Aca3il6/rJiKTOfN248SvIYME9DBLC0jdnkevpvxnJL2IRd3C8jlzastb7bgb1PLoE+aXSC96ecg
ORvkPqzyeiG//a9ZDvivsaAI+gQIyo4M5oyw1SDQRCZEOkvThMagEcyrxqj9a6Lc56q2luA2ddmK
NUdJn4i2kDkU+YeRMHG+E7/8UgQIycIHSXKnTzW0sHVMHv4TcNJhF5Nvmy/igQd0HGxnWUR2jbYP
Bzp4llKstvZFZfAFVLM5SLdCqiUacoJt4FmkOG/g756EF44y/kAbymr6B6S3txFslU0rt21ucscD
ofxwf+RojBBJ3QJwed+F+vw6t39S+OUmc3BW8BbtIAl14i7zAZZqZ4b3P764NxMps62c8za8Rc0d
dpEOjGPDXgn4zhrWnI4SdqxgjFSdeuSDNdeDJVdGTmHTMWgPJroVYyW99fN0U1kb10UqrXZAJ65e
EMa9A8iQ+u2Augidwf4m/ZhJxLM4j7fDEkPnzELuN8fyPREN9eGtkymL1K7benAnh48gf0rmVcDg
mfnajtU55yhGNcEMPR+NkBB794bQsTI7l+MS4BRvMkOGfjsHBY+i0NGHbAPEn6JQ0EfStcCz9Iis
L8nRmTDZaFDtSxyGT+h3+qwsa945eiGxwOiQJiFEXTtb9/jeO7LUv1XmItoFMr0uWyhxtO9tI241
LbzjbFXZbit0izw1q46KgpvTAb4UZczNvFHPniwMaLU+9gUxJItUIPRau5VWgbfXp3UATk4cG4y5
eEpvL8AABUVvuQwHH6f5qqNL4qMr5yFJyoPezkL7UWEwFbEpRAClEMLquZBi2Ip7i4WIdaVoR7Z7
4LZw5BYC8bgzNb63sEkWyJ3wXuR+Vl0T22TB02d07DtgmZh1YEJw7T891sEyQopnp2/nl7cFjQET
QuJ/pmwUD3WU
`protect end_protected
