--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
QSRw+GrdyqjtBpvNNOgJwXW2r4GwNEhXWCuPsK4ErR0QjvTLSLZqtBCneVn2u61hCbB9fRRjclk2
Rv16nnW2hlb09P8KvtEEwRRdcihZV783Sf9ebkpEZULoJPAoGHrtjGRVbcf/HZwKz3x3/EMVDISt
ejMAf3eqpUwvGA4M0MbQdjYEuVpBEOq7bvQsxnDSQREWoVZBvRB5g4t09zKtfEoqT8h+Fk/p+Trr
umx/DBoOkGHxDUlgBPpw9VD+cn8Ie8ox6c6UJ2vU+rbytEvJjOs3iq+Dq3kpTxuIOmxBIKU4tW7C
J33XyLeM5sXtNT98qQKMDGZ+vGHPlPDag+JjEg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="RRi6CWL7DBCZ+nt34bB1HdJbfAh6a19+eHi3oG0ErCU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
JgmuHWpIhAFnm2/OPTHJQKYHl0vWXvBbb+8s5BX7SNn8X1ii8jepFMFcBGHHEoJKfUDxdYY9aCd+
XHwr/Fp5rSk9RXXyaorkKCBsp0+sd/vpWyhV+lgIcO49oIhhfuT4vAxp0gbLTWhqd3fYnrKZbsnt
l0zrlVnxs47g39tW+Nw5utdk1K5qhjmQrBg9uM0qaNMDtfPVJm81PFSL3pbuq1jFF7+5/7Pp6mI/
NjezW00Hpwkddan9s92+hbsI/R7h/7QzM9v0t62Ia++Bq89kMKkhUTokpoiDRVqbCU4T21ihQB6O
hc4C2SXIE8YcHjyJO4UVibWqiLTBr7t+Qyh7YA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="K8oNtDmhbQqUxacn0TR5LnK68cDU0ziLlZCNlnqObjI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10368)
`protect data_block
9LbSsJkjJX99iN4SmgTSZWc5GHIDs8gkXLv9NUwzXTa0plwv7NwNAC7IVmya4DbVJTpH4BlbpVZ8
EpZ91r/P1F+neSE4lSAUbXRnrwRBUpkvh7oLd9Akooq6U0Lu+yxrNJcx5JBFibgiCesgmoZ36g5P
xVw232z9dpTaSN+umwfQzMVx7JArQjlL/s6x//eU7Gyv+qdLGbJDnstPfd4yjpzDVEnxZdjk1qIa
V3qze2QwXXCfB0Amvf0m/L+Ndv1bIhGsEXRDE5rvBBLOeXOCDNLBJPJWndGgDVTE5tDIUwRyYMrh
EEyzsjcMuj+T8gejd2MbTaxxlP41UOO1co+UrDkpD6YsrlCcnRGKZ5ImUHc8gYeA1mGg3mUwTb4J
16X2EEptAazv6r4OGrUdhbnKIUu2rXIkKN+Ei3wZ7K3Keai6Rx2DpsM2LcaYhYyAow0inq8KH3vW
a8kZ515ky4JoNA3ewZO0EXmGgwt2py+a75LfAe2TZ49WOmkiVyaGNv6rhmpjdCJPtl74As+8MWFF
/shgxGy8vFjKbSrwlaXHIqwT4XMSn6AZN/SvjQPUcg10kIS91JWSJB+AeG6diW5scgrCYDM+QHch
SAOn4jXogFvdFgB73jnX4PErUns5YJ4HyuO/qf3AjWEqd5mpvJsw3t3hKNY3fufAos2eWrWMx6Ff
1Jk0VwJBEZ7Z/xsAvPbFfdVj9qKAc7i35Yif6+RZjXdBxzRaurcJkce5jMXq1VDf0bdHrEhdVy52
B4WX9Yg0oTE49ic8CL8ugkJ9nQuJVobs6sPluJaz2S/hqAE3nw2zCHXrwjxXHSW1Udvyx47bzUrC
G6nYxfMaYxFwX8RCabgq+gQTfME0kjyw70wNUN4UU5VMsqGODTC4rWQ4bBR5D5jAAH/rQwEInwIg
y3XBkJoA02GyOkqDGT0gXVTUbE/oymp95ZERHTGk4s3FVGDgpSYFeU7LI5xF6MkseZLjg3EQmOpk
rgYhmyOFcgdGzb071L8utR/R9lP11Pg0hJ36mrQCyuw053RXoZ0BQamo9uUd2pHkFNWehEYiSvRE
KxEesZuusEzy9vQWt63F6jifpDUvdc+0sD5QXN35z+OG+CbVkr8oCh9pP9fpfAx+8xAn9TC8VDYl
UblhyZ04fh6Yu5timmN8sS3R6uMF9vpR44CxD3XGbH1BTRpcr4M83REDwEiMGvKOTdqMuRwISGkj
/oCaHfAhVFc0JjthbYkuqPkz1bNToTq7C7DZdtOtyu/AEbDCZuSto8mJ0IfEYe46AOJRXeO9SquL
NOvwi3unoUA5gOdIIq50KF8RsvZuJxTDg09ie8p0U5RrPotL9WrhNu/mucXHdJZsMcoXkxMKbIpn
VFoR1T4ffp5gAsj754XOxBmRBv9ZgJjaw3b4x29CgioI5QzOvRtrXty+i0KaCBTsKKuNkqy0QbZr
8NVDH9BcZWIta2w109WRnNQge2JQtWKbCBS8zxIvb1fShFlQs4QSOrJYm9K6dpoDZW2oX5pdhTYM
3QYrxQCuicjchb8OKQXMLKXur2utBUTKE2+tdERJFMIQha+hFO8Pd3sW6d/n/6AH4gWETVFnpovq
aVYxoki2Khl90+RgPDpCzYTtmDrbFGIJLlR4IvnW/U6uRjTECDD9gWyJKmjz6EegoedggHSWXfIH
wQyXAj0NUTCFORVj/9XUL+JcVSMmGGdVMHmmr50ul7rHo2JcZVwxNLm/k95sYmuBVFtj352PaoK0
BA8O5ntH1hx3PmLr6EsMlgAfPayMDUb0mJb0urVAVnkQyYott6IP8uY+CwXEZFj6inF422aoNOgs
6xt1fvHrK4fP66RJnpzz5TMLmKd1sD5ZV2nwNXuXlWyY/OrdnkN9kAA/pZV3LaIkGEnsrCaV1cVa
rw1drz0dNPR8kT/PqrIWKxbk9euMMNMuFbi1QVOL550WNM3afnOqS6p+4LTHl/4LKMSaWAlNK4p6
mcNTaTP3fn5Lk1gbC5gP/7jM/s+NdZmKQuh3fWzthJjqteRSOieldfDoldEJ+QJD6lG+C8Ug62ww
FPUHeVK6UFxBegpivNES8MlUnqZh8mkorIb2MkXR+u9IeH2Kjcl+KM4so9O/BFPaapgB1V7RtkoI
AE+UIj2QsNE7F11BCqsv6Smx27heGpkVnMATfVs6KyfaYZKxw9GQBpQHzj4QJtOKhuUUSEYaN8GZ
oxWZMWAlA98lf23MxUP4xg9vis7JWy3OJ3f7K+rq9FgdI4Yy6765SQawa8TT/T15qt0u1AUHqFKz
L05EGuvylD6+0lF0UBse8HGVospA+R/GLXg2YBS/4cYZ/j8n8Vg+X0YO4JvhhwR6EW5oQYSob4gy
WlPFVeUFRAR5fiZI6U7OY00jxzPzc2KJh5f+p8zxXDGjceYh+jVSuwAgzqOIoPeZu/9Stah94W5r
/EU14jgJ+3Xpj7RNsc+mYySetwFjHuy2UdB6lJgiOmg3M/7qLsEbPNvljOUDBeL6Ru0WlQUbdzU6
qUvKrBwHbVJ/b7wT/NnHIjBHlmULEFsi79vi0VCy2IcszIw3vhBR9fQpzS/XC8s3hDu1V1hPzbzD
9msPCE85/1m3tQAUVOMGShBLbE/2+9cOD968Ye5yOEsrdNlQye0hcpJfarZ+symRfDPj7S7rbDT7
ZsFAk6HPrdVF94G4r/ubhu+biUmyPxShStEYY4He8cUmk9uvh1amYopFvknUm7iFS8kKrEuU6vlg
9R9FiiC27Np5pA2ntX9xwhA2r2ldHHbmmIa2JWRm8Ikm3hA2SykwyvvjvALPUGeu5NuBmyH4yMwK
7rOUPg0nXF3e6aPipG38lsiVyF10qHaizybYOr7OJFbITIku1gpwixbR6ywkyVajvpFEvqILb8JE
+qYLDhaFtGYuuNcqUY+1NeUOPjKuzL6Ib/pbuH7QHf+idkGRq22nig7vXcmx8/TxoZT6H9jM2VSD
/7vNmwaatilYYsh+sQ/Wz4sFo0fb0LqOnvIvIwuhL9j1zF8usz50fFyLUOSEWQwCDecB9yzSzmTT
Lz30BkZ17FwBYXKL4XO3p3XaOcqrX01Id5TKe18F3lZdkHY73KTb5QfLu5kFiCJtXQijlqdyNXcK
0FaLP7NCSQ9Xp6c8WdQq7/v9VCpzm0Kb7XqIg85xDaXoyRXZ9z1wlzUjGQdiOKQhYWtPbFi1iZi9
ioTTHJN1Fh5jOH5QWbjpx1w/8+D9xwBpVKe+ZfExb3PNSNhrUfA5zuxQ9xrGKxg6scwTn89bHqLt
Xkhm75L9YcHHzLeHhsPAVL8sCTiYhCdjLh8OPwPjC6lTNE0zA1jsnr+U8UeIGjtGPG83wLvdow3n
dqYarWyTIWrotduEwQVOApRUzwSj65PDWLxBw/RDni1ih8Dj4Hl3vSVDKNg7QTLvEy3z06wmzLv5
/6SPHv0XUx/13FJOIDufjRf2Ub70SFMq6XJvJpgAGXpSqBgIDnI+aCjLTVNVEd7TWML6eIlbOx+a
xO6/bUsLpZr1hF5TP9vJdnbjiSFaeZq7mrB4R0h5AaZudTPJY8Pr5cfLzZipLrZHJxsPFFm2psb4
HMdl8wHyd4nNpTRTAAKSzSI2gIAXunqY5jmzN4ArrWf19JSz27m3nsUPJioxgOqnIvyBGo8HEcCx
stPDB+iwPo97ChFemfYCcFagPnI3AGWLpTPrUQotqpSUK1PWK3Fa0BpJnDzo/11X7NVfnaKhRFSy
nDovzBzZZp/fQScNzVPvDOjIVF/TI0Atq3iEB4b1Z5SPvD7c9eEIwxkEwKQAphNll/29FXUr8gCw
AypbtMZoQqBzVvS7DNquvj8y4Wb3HvDecbMbYk/9DVxBfLv8OX8CTNzhfzlYS2F4H/mXZONTC0Y6
AEp0bti/KtJhYCv3Xu4uT7Cz79Niq1kKGmSwjTujmCfKHycSJBXfE6vTHEDnV8n1rdf837CWmBTZ
EkHCESPBWFaJZWJmhPf2RXQbH15QMZecYRG9FGQinrG3J7cBXsjaoMsfY8Ny/6lFTD7fcInTecJE
31tMY1MMYQgk+Hpw0C7qRky2B9xWJJ51ZFbf6rlTmGF/+XYznrojg9M6ea4ePtF++JBMKIpASayO
6tvNfRVczs8IxJkGc4qedNY0Y+BlK4EK7a3OMHz3u+/GQc5Cec8hpTlNAWPVqgxoSQR+geZbURSz
vcUPVOC3C3Sb8rg56qHhEpwVHc3cnugZfiNHJvx6/nxz4xzi+/5EUZsnOLrwCY3c1Wxlrg8bEkUQ
dE2SgDlbKnaoWorxkCwhYfQW4bmsVDb5Ftu5Z98rN/NtdkAtfYEVdnm6WfCorQdCyfhVOr4KfPYg
6MSTNTsDJXAafin80H+vlVfMV4d2TCiGs4g0G8XeHZzELHTIJfjiebTwzNQ8t82n3Ul7PofnwFGV
/ZwjUQMYFY9wMzAbWZwXt857bg0x8UilCduu1wHvp5vTNaGRT5GGuMSKqKcyLCdHj/M9H6lV6vPJ
sW8yDan1K4qxQypysJpZFlG2LKs00OGxGlN996RfYcZedKUEJql4uo9R2m5JwbsJTdB2goYSHOdf
R8Xh1Ca3sPbhvQ42nSTh1WR/0O/DUznr/Ok76ayTHpQHrkymmuThevdzZtW1Yv7ClYivFhSZWHeG
VY4/iWOe5OATjXWIwu9bkseg1uglQ7X8p979cLreUIKgnfXwuzy8W7VaZkqHl2AHoqbUUiCoa0s0
rqdZ9GkO6BRKH35e60HmwzBkLRNVXx7yZgmazdh1OdXOG7MZ6xwMJlKpz1X9mrHgOUxyj02QSEXD
QM1i8bA1qaUFh7r9NtYKcsB7/ZNGXTUb4PMgLWxEGGmwW9Kejw9yka/JZcdyHTAVvmNfzsk2yxx6
vUajlWLmKekxy4okxFgh7mq7SPtDSsaAiCG3k2gC6JnCweQfbyEkVQvh+SQ35AQFEC/B/af8e/8A
Afllj1X26wDShXmoV6ysWVUAU4k3S2LgIKUNLQFD36ENMTOlzgV/CuS1hnWh6LbIsrEsHYMByld5
SpJ96Nhl8ZspkfXtNxcsW0gZo9u8v61BFGhEr78WLCXxtiJHWX3kijqx+WKXi/7oq7Sc3j1U71LK
u/u8kqiPQvgh4YZfHS2VSjF4X4lHliRySq7BsKrO0eWTtY7LtDUyBrXYjheKGpJArDD+w/kCtcdN
hbGshUssV73UY0NrSh0BV49OvraKjyhEmy6IATmi0s+PHTOvNtWJH7zNPZE+MsmulcVyeG13jAci
SObSibMeH1DCLbkC2BKOTFmyymuGYP4DfBPKrZTdAiCDeKBT8i+36zKQqPc+sC8Px0469+Z4GUAy
V2SUSUohPyR0gG61VW23poRtrdpm62z58G70YaMSvWDkOh0NAa+oYEyUEFKu6qnPaOwQdflCbgbw
/axSAGET0XCctjWOflF/O2Hgx3NZCVuJuLpjz5HJBtqU9GQFCWcxnOqhlFECdRtaoYi/C2TDYC2e
1hycVIk++LwD3BjlokBdr7Jr3uWL/uRjHFp6np6OaYfI+AswWJ9auAGTxrdXy7USVEeLpkEH+NvG
mG0k0u8+yBnGiEsd+218DtBwuKVADJomeojw7wzA8IbElulhCTPbP2pJQbMeaeIIMn5RI/jxILUE
Ff0zc7QH4q69HjHx/5sFZYKNKNcz5JGaYW3iMtbLzkv9cWicqA2X8jSPqr7C38HSS24Lx0s6ZJXV
4rhra9LbiOThWenvvDg1VoMF5KprZkU2Dkc0I0W56xaaGc5brRFdv5nalcF9jKN510Qhb5zMJ2jd
16MFnNd223sjxhLzuuYamHpeT+z8Ul4ycF598vI76Cn9Rs0g2KqGguFdCUMMLXz99cZ5/g9sYEfJ
jyZ9HcgsATSQcHuWx1AXfKuW1psn+hp7jx/Yep4TXznbnXWbdjwReSQRdbr1nbL3sbZqye21YrE9
/WuUBl5sEWZtmqIfDbQQRr1jOIsH3REgAE0kDxIIy/wK7ByZAkqxmOrVbhpDZgCXmRusVeOccyHX
8R9lhyhMFxHT37ImvsHX+xFWVzTgkes7jDHomPgFoFnhVi80YzJmFXhkodasUhVooXOt/+IQlBU1
6tdvDCwrJWppcz6vUMlqH5bdfMHXztbhn8EccjeW/qeWoARY4o+h5MdWYUcZBjfQ6RSaJxQX7ThD
l/EINZvuPNBH1e9IY9LTY+Ur3BrG9vYPTPCAQKHrQmH0L3b8t5yAaOAAmlNDYuyUsua792upopCF
SQTPLZjbSQ7bCcyVV84503CTV6pD26bwMt8V3m7uFqcCjy3Vpf6kmtCMxIFz2IIzReqe4/phcFK+
TzeWG+IQRb7EAFQvojglC6Gjsiu3CmBLy4en1g3WYJ3PYEAr9W8vS2ZZ7fmyoVji9cij1EVrL0Zj
vfCRPSFfSUE5Nj6FCwkrm7z++4OG7kOn7hLXOuQp/AxxpLXb+y0OUx+6lkuR0CiezFreGLPkWZoI
ldrHoaqMu2vSJOFefaYf4pQGjyzOtRDao5rNkgoYgs+LuAtXqECXv9EYp3qY3RlDewf/dxY1tSZT
dY62M5hdCfTyk0K5iPkKzoCFqunLdVNeSZVIa6MDd7WCqW1fW8kPuE5eaaAOJOMValcTV57CNOzA
dxGn5SG2RUsmq6MesCK7wV++DMuPU/D74oH1Ul3j2HqpFyEkHk1wvAKU7YSofGukQ1DTPNXIJaHl
v9SLc/lPMe1aePVfqzcRn9IIHp35LlSqFz+jgyBSBFxQ0PVJV1eeKg9y3iduYh/nkMbFho/UvZ2c
JSSp3JFeLcIyzC1tbtLGnFcf2lrPnPimJh10FtliXpP5wJMIARQGKkjQlR64tm7PC1u1m8TLCLsR
UMFW3A4tuhjqCsZCHEbnyNCDVoLWqTsIhQ9iDP5NGgBKr8giY6WzQgZGvhl187pfpqfUa+1Cm8yr
VbhHOuk2nP1oKCv3+tAlmAztjJWe4R9vvcuOu0gcJ3M7HnT7Xlh0G2TgeIfINldYtXrOVfBbyTCa
xpDeMVJXwX1A3qbPpB77FH5LOQla6jyB3Fu6bAvcrrkoi88fsi3gSUNLdbOcYauqkOjUdFWIjx35
M4BVFvOGFplMDusHbVT0RS5ELUtDXp7aS3VEMhLAvILi3L7VFhpo3/QpdyLH9XZXBd4Jtnx+XXek
/h1kZExa7N3eEmyIQUPKczgziMr7/BMWQaeuY+czH1Eo4PXjIeU5ZglNAaY9+H6OAig04W1u60LG
qTTZGWxQB/Iho68iV/bNk8aSH64hlsfNM1OaUW2athWoJ8RtJ2/c+5BHMEhFt8mmHfbl8p7YVgI4
LriEF94qRe6lwCOeoHZbKlzdeBr2kuHD1j4sH2Y+npB5CDnNqPwalSRRdgrEBnIaUu8aY4/0317M
YD/S+P4SccpNeOcAceIfMDSqdNMjdwqJL86XfEtan2CnBN9I2yCvnolQ54cc07V7+fiGVy0RQhKT
aVMtB3U2cn/xcluM3q1V+B0/vMkmJVpUqyFAKsQW57xfkJ42YSnVuwiMoORNBLH0mahuMep1d4+k
erBcBEXh3/anvCLyZCjLCScdHDrIijsvT1obVOKgarnkv27KupZEIe5VRMH5LfsZEs2HbeavhRJ3
jvqerpBtN+JPCClsONmq2pV9ydNFBhFvYUHp3BqUSjWZOm5mv0b+HcPolmTB7LEiibWrtV+ZfLA7
7KVYiM687OtPNwo5NT+Psy2SneHWJBYsom5Ggv29TIToIL7Ps0OrNeFLvp5ITId5sahe3hb6ws/I
VwWHnxo+JKsz9OOLnuMKVF5U/+Hn98SsZ14mAm9zz6YDmYM5iM1yWJJ1qanh0mjIhKtYhPLeiqPn
lYz2lwNrfA6bcx2o/l8TC8wot+vgg2sNWAWfya0qVNrGAoIVaXespEJ75k202uC/fwmI0ddovxy1
fF56iuXxHL3YdFCGifX4gPxgz1CbeuxeBRafyLklHzYZp3QT5PmRz7xP8TWM2NQhrS5JtLMYWGWd
pWxKAIAg39aTHhku2B3xY4eu1sZ1r+6Xk4KRHVsgmdfWwHHvp08TaYUsyXwSqqS7UUe9zdKvocK6
sWtqxekeylmqsnCrZ8q4oSW020zHS/0zeTM5x/ccu7QkXBrOP3aenndg47eWw+4PyDDE+2MQOQpc
7aa+GmpMPPD7ddaRNW51VunubybHzynsgTHniGPwqSVe+1qoQ1WmoYIq5oECI+JnvCmRN58Znaym
O8VX77kXqHVFp6MvuQ6+NLjmbQhaYBldQXI6PJB4D+NdEZkrqu0RFgqjVfO+5kK4WzYrmQ97rJWL
2dVsdqeSYcDQ/4keT93BuCHRy9jGz0YKkbLP4ITTJ/7+RMIrGO3kOeBa0nzomya7P462Kfstf6q1
wMCMaOS4otGpY7hwE58bZHGC5AqQa5fm8MOa+eFwLZk7jcCrKxS6Oeg/E4J3yvV7jwkfeA3bLNth
QA+WhlEt7LhZzBXgCzkZnILzRNbZkuZzabyK1YsWj4aqvqM2b8E/Jwfpy+VGi0ZqHkaA5FLS2kh2
0ZGsK/r8s1BOANpV0dQ2ehcQ4gFufYANaHlFDsJ2254oFbRX6yeJkXXAKoSjenKz4pvjS23oPOMO
p2hskIx4ikGyLLy9L2ZHFJ86UuUQ8KAtrh2WuRv8OnSSa7BFXd39i75AhuvCs5lm8Ukp4H+bfw9u
JSPqzTKC4RPR3s/n8ALUz2im8kzg9oPPmVlObA3t4fJcB5wOzCyX1VKFDfkPIOFmD6ZwCe7rdLax
9CxGrOv4zvns3hLZZ4RLMGF00gvfU8ufGY4hg7LuaXgxXAP4Q3PiZp3lDs5K2sj4v9ZReSe4NU1o
bt1BJPw27o2xGX1o+DbXJGvEwtSPwnJcAIgCOxvXz4HP8ouOChogTj+xzMijeyLW5vopyxEi3T4G
1whEOxzBgDMGocLZrLFBm6/KsBGyXwRiFNok6QvgfAXV50mMcANS011gI81txYM23VZ0lACh6P96
RhVNqYTSFeRNn4rBX525j+ddrzcN96x1s3feUUbTkkWMbTQ+OFsZyGNsei2x5xJ84azI9gNzHkxn
p/hySkn49o4EiZzEybM7nE8a7v9NVsriLpQazaQKp4+IrWKwOBkcf/OiDhp7txT+i4M/+Z9eZhwg
gmFAd1qz2kXFtE0nhh5CjsnqZayxYmhOjYxs/tK8yXsa1qC6crShJm3kDExONTzftEn/E395gATp
cyDyh2kIf3nMN+++kSPuzqq5x7SimzeAYatvPvPNK9gwaaVzJxy5ZTu4ov82eYQZhAwiSW6W3PM7
5sUaIg+aGP68noXwGmzXhcR04O6S7XJqZ1AwzE9zDxudaOh5ciCUvN073zYgGYvOuvSum5GpUhj0
oUwksewrrTi/oF+s7ckNVU5PIxP+BbtwfD9KYpILxmipO9l22IUmM2KO65tSvu1anQw+PWjj8DJ/
vGuIu9MRHbjM8KD3rWHW9oFGWYOmLDorMdxq7sDkPc04dYFl8ZDQomOK3yNhS67Uih4jlooU3UgO
ZYCjr/ZFNR4PGD/97lRYtMsRfhcVWfPyetTdc3V1DNlpUdz8X5jmam9YHnHAwPE3JLCflMQQtVO1
Yv+DMBrV3ioAm2WhogS/tpecsCg6cfxsbMbuIbknbQALozGP0czrWzp+Bp75XTIj3izId3JXC9FW
iClRuIzsmWETqJqrjPo3WOobW+oXk3neXsHMiagRXcOE+spOzuwYHOjKkK4x+Kk0oZIpLu4TbS8F
9T58U5t2eRGDSzhE9Cbl6qqJINyzfA9fK8B9TYZMnqjFVPthgMTAq+BY+0gzk5abhyNuU/vxPAy2
bV+2UgkNRoazWk7XGYZT0PIHrugwO2Gkn6eaSP6YWIgCk1NMpcrXtaRDEVBbgz9qfRMI2a0vokdj
UblDnKM9EyddDIkRssWO29j2hwwXU/4oFnzGSzBgc5k02intBp6j5xgIYYP/89K8kXFOnYJae7mZ
P/pOOMasHKziloR35oTBUxjpczPumjPVr/rcbmIdyB3y+I1NxpZ/sfi0AJQfvTQ942D9a6u8Pmcx
6oObvUqazm40bJbGtpHBsHHBmKtdjK7tW0ZC3KEeG5mCrRMXf8+/SwVeRcDHXuzkph8PcQKEDWCX
b0qnJPEvkYpDh0MSw+VEYFyCwH4IIPkDXN0fNqOvuzby13XUVs6axUbNM0IUiBD3UhVwBVRQ10PB
7QI8vLAZAwlwev36hxEVEJJPYhhD8GivDBMA1zdFv5HEb89GZMaJOM+qJox2qmekzgHciaNh7NRb
5AMCevQAWDC6zSdbFssaENoOuh/AGXuUg1OfXnkPhM7t2pbd6YIsYYEvZ/+Y13sSkrILSZVZCz7A
74nlHRZYUTi2tHoNEEA5H3y7LQzmpGSb9BO4WJBqaAPDQM59EOFCM5FpLEA8/qa59C7zLDVZwpRl
37jGYJtwVcQfGyNIySpy87U6/WlYyOEtWPOsfaZDqd9LiXSge3mbCavwOO4Pk9SF/sqHAWGJgZqV
3QG/0kxn+4jP+dL+2IbtCHWl3WykVbMpIWOJ9vZmmU5+hr3WjU9sW+xlhT7u2hX1WtRfYnZiANaS
OLJAZ4cnc+IxWctwhYmlky7rCKg0dvP5QVW1YEblBcUYzRf/g5fnnrDD3l46QLLhtEvhRqZYX/I2
fpbR5e71X7s4HFlonkGyGnHuoES5ZkPZQXApuokAxjNLMnHtwMIxfyJqzYzuPs3NHUx2NIL2WTdH
J+ATffWbccqub970Zfs18OHkTmBabgszh5lPjVWqzA+EHC9AhpgHbrqTe2RBHGRPREc9F/wZWOaF
excubVdEjwPPgD5LnRm/Iea7v1rCVuHARQAv+GSNNHd/vV1Pwbb62SdI5dJE6Fo1b/8+7JhGyf4I
A6FF+FWT3LjBeXP15oNVQ1XVoW5ok2HvIGdSVuFUeQ6OqCt8VjmX8JoHjg0mJxtPkju33ytGZwo8
W7OEXttcE5IMDJMwA618nGwhCAoU+XbKMzlbO1s6eE98wpsF4XXGoQfkRkWKj+PzdHgMSO7jG4YG
zAZ6h+djuYZzt4WggGJ+yg14On+LNUZbl8ceeVyGSLhY+uKLGbtubFePEKtBXj1mLAUUPxuoN2Mj
1fWFabm1DmNcHPdLf7gU+/9Tt/BfXA4IIXWh85Ll7HpLV9557RDOOuX51GPz3QGqmF3lEcKVOOdG
1fQ/ilSw1YGAnbJopr7nTov0rEZ/3OF29ufm5ew1x/BkWFcZrTBR+6opMpRKCZnuK+U3qMvlxher
Rx3EKn5Cj5nz/myS2UUdMAScx2Gq/NFkfAjjbfw3QY3y5dAUQvc6Bpj2H9tunmxjgpDdRJV8QNFi
c6+nl2Q2qduW2Sbg6Z713DVMpCU+xwsbI8HUHVnjXrqGjteTtNf8f/S7W/abpTeNqHf9EXZkLZ2e
QyNiu9rCQJ1FSseZexntqQ5wM3cSYC0LlSL5ir1U0HG0oLfswIotcUweKMyWS+bLqfHt7tcL9CwG
9XI7bnIXdh9C+zZ/eoeilbOa4zOGfL/M6Ix31aX2tFA1raC7ttL64lpF6GeItqAEdiChP3NJSggz
MrwXnilT6/aaFVVBtBBPUsA5nyA6eWuv+dyZHR6kIhKdbvV8GbKD12mBSMYlPf3V6YoNq7JcAx16
jz/MpJvDerBMT1ueiYoRvb6gTO9zZwdJZTHJySN32QaZ+m3G7eugMUN/ZikPXIUfVr/eoS9bMSzb
HTaBfDtK8xgWJPCBtvbYri8dL14sj3G2UzNuTsS+RKbXXLu9Nz/gOuRGORNA9s3ItolrPOT9u7BH
xenEJLv43zZ1eCxP1uvp86/xvYsOaYbpOJwtXuMUfYq9/4hc/kqRFf61DQESk44qRxBH3oBhVxBI
lR3w/6f9Rs73w0M5BNsL2i3n66R0V05aCX6oTvzdDM0oVwGeptVykEvzBaPkVlbHeiVMobLmH+VW
7+Jib7MidJuPDAQjxJ99ZXq5WP8M9k2O6KREUWHoOQ38DB7NrYwMTCepmzi3rBkS3ZqBUAnEzDUs
zWvoEmN2Vqjpqh7ti1ijp5tJ22YWcDaWdlknU2o1lIXYCocx9yVgs4Y0pMCkkW+IGUM+DnRqYRS0
sMf6YlI7bZ/cujLOajUHpK49Gw0gNXkfspzliKclJL8Ihn/qWs/Q/QJHq4NHKkkmt0f3ZDXbVsaB
IyJL1YlqhyDosKphkiFpmwXIkBmSh64EpF7TrQQc/Kmddb1cwrVuDi6dKrQnZhEaqXznFV2C+Jfs
qn6pK1pmBnLF07mEOsO3yH0nKbWQeHUzFWcYPb0XlO4McXC+Z3Vbe8m78DHITFBh30nxzxrQWJLo
EhaEC1zuFJXYa4in2dPnaekBAddtnRBBUBZPcgrQU3w8U21Iu0uZTfiTxlZn2uqs4YIB6AyOiv2T
LPlmbmxE4gH6tCfHqJT+4qEZT7EeHfhmBkGltMHTb0JgysezA0Xc4m0bu5xjQQxSF6qE2WegB9vp
CuS1DwQetBn1a2Fn+pV8n85eeGFGxbUE/6sELXrIOFhdgKiopQ9XF0c4Kg/SNewFLleVOoUzszJJ
b5Rv4+oE+ZjA/wP5dTQcHuN63+paieycGBBF+xsYT5h7M8NxgkeKgeR4YzNKf2gJuUFCGuJ8J14R
MbKNGYlD7lroYEoTIORS04cyZcvxV//X8Mnms5o+XyMzNbB9yG/HgA45K+gjWrKXNCab5GQ4kZ1H
e1dI9eqPSKCcJAT+v8s9HP9+bLUPBEhgLSD0t4fck9OtzreKHPJbukPCXmR7vawuRf4vrsdwVsSp
jknEbwIyaVVCUV748c0gI+MNteJkq6S5bnLWiZYKl4ii6rw4Krk8jbBKr1j8X9Atk6vu9ePi55DT
grxlpPwQq0SxG0E7Em2OnFgx17YiJAnDSGQDT4A7BllvRWNUM7isXLCJKglHmwHBvWc1QKQIQjTs
JO6XtC3jouz+R/vMUnqSKEQGYmzP2c9sriypRwEdItdLgM0VlCvvFKzBXcqs7RzuIiq2HDww/Guk
8OhLb/q1Eb15sOD9LuKZo848UWqd//yKdTinhgd9uN+AZ8z3EB+HSUAIhe+O9l3dO3rG52o3Ga/o
URShBaO3c6ZcOG+e0+BwjHo7pJWitBDtSmxtB2l9hoQWIFd90kvEmzAoviW9ZSY4bK9RZ6LSVxFG
mvombu6iZDAFOi2LGGAbJ+DGUZUqkq8/j9lNK18Xg1Z3N/RqT/ZNrJtD83PABIJ18lzQpP9cwafU
30VeGPAuXORXI0SZjcW78DSCL9MHA73ZsIUj1tq44yS8W5THzFZCphkuQLFwASmisYALocDSNZs/
PVfsd4LZ28TCHe3a4AfepYGp2lMKJNUEcjrwrxQSK+aQ8yiA0Cg4QhASSoKG00QlHbKCWKhsvGzk
CClmcc/g7jzOo/Z4vnKA4jS6lhWPXJ9O7gKqU6c9X2jSiuubQvSI9YOHiyEepZQdRZnV+FerLVvx
lrhWRcQk3lywLTgJxMgs7V4JoOgBPJQRX3I3WdJHhFiXpJEe3T+gUAu8KWx8yXcEwqz+vQAKyCOu
edmHwYYaA4Vz0gsfNQtessg+b0w9jqjRqLNPnL4mq/4m14SKJZJXjuA2pwvjwEsurtvdKY/njzzr
8l+Js+rr67Z9FGBqlgRfxsfu4StQm5O/35rQDLXu/2wa9QsfkoP1r4+vxyccZW+GqjweBqtyCAnb
TB4L+nJyUsn0/ep8tjTn0a9ZoSmOnBOXxc9pDu/a0lmVKZW5spd/2NxcDoYtYLr850G65GELKeam
FOggX4tohubjsCwrMp965Lz7YImwGwEhvY+kKK90P4iAGcg6Z26c+cVlAtFwGzNsOxcN
`protect end_protected
