--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
axVSrMrfx6nznYpXga2sRWA6s9eggfrLS0fooV2YE92z9wejxlCdMnrSYOtTBxtR7kdx6SoXq2qs
nQR6F7XD85535TXGZXnkfWi87oWS9LveSK+Pd9Wq8eBPYiO4FVNjIcM4LD+sGdFQ8kSKmDn0/vOV
pY8ZcylKYwnyqQGCVfHQx4Bc6B1r7A/mwlN8roDSywC23x/10SGI8rJflmqaMUM8s/9HrZh1PSKb
w45ObWqY4v46gJ6Mbo0v8qCrKjw4zli4vypugNlNpaaExGV4OgEGeEBvhIjF40jNqLhajj23t4bt
l9jWjEx+pMZFrDqXKy59vV/iLowwBmo7dAkTkA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="pxR41uNY9PpkYepmsNAfXtzgfdPPMZull0Bm9i9Xnrk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
PH1eNtC7TYT+J2UtPf2fr8RmJrPCzc/5ZN1Hh4VRjMuhzT9lr4l/IYEY7QTkh2wFWfnsgpfVNlEq
Xavpo2iXPYIwduTwPyWTdSbEMc657fF4cdUasTbrLWz1SyREx6EcyZgQfpqgvZ7v0woAMiAu7nc0
WogeAO3CFKKhZBLzhjI5WYw+6sUBgrHHyh/Brh1Z/g+wUri9PDZf8B4otXcSeepUm4UtQAh/I49j
DSm79joiFLE6nYoTvdHuAzzXadsryTn27SpFcBH0/dUQq7hvRxr33EEmMVs9Py2XJ/Gy+9wB2rse
QQlKPGXN3KhuxGsK+7iMx+jsbErWHTYFB9rxHw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="cr/bh0pBTWrJ98Ptqum4nvqmJBkPUInAybjRPm4Gtes="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22816)
`protect data_block
6Skd0S3N77+8FQkg64xLZrDXZdOVbnos24XD4DJgUdPDLhCQPS1jvInJHi6CLjHeN0SQDAVUj4dG
ULAni5Gg+smjg27ZdJKBmKW+4jqhfQvMNVtR6hGJYD2BJvWl+Auw0p4x/9bcFvhHe2zaDWQ64SgB
zyXp3NxT8049ZGr1VUd/XY0zhgomUOQzQudlmntspMfBavh7buV+Z4c5FgW2Ri6Ya6zUvJU89XCu
KGx9/ooDu4abVgcTueY6afUqv1E/0GygkgvXBBBp/GEf1SEtm+sRMz2ws3FM5dVu1CWxIW0B6bKz
/SaFxey7gRfdN9yNFp+CpOOeSV3TPec13kbiZ7bvbgQ/GxaAEeebzhDuAkPHyIKVJoW77Md9VDSL
5M6WqOaiqTAxF+WsXz2u8GaoCErzXUTfHTo9POI6LLDTlp0SOHkykGTg9RjdVAoVA9oy7mYd5Wy/
vR8aoG9M7aeCQtgI7gIIOhQpiqOweoIXo8LGmjxOt+qD9lbHOLu5x/vMv7UoDLVrIKxjVCY9FU9J
2E06Su0UWrvFt0WQq0iAPG5i+Ibq4WZwu7m2XQ5mEK74j5u7y2S0KnxGIFOE1mjkPj0hl/ftKYih
SeKoKzKj5lUt68Ysc0xf1lmr09WcqTpYhn/M+uIwHSIxSnoEHl4ecw/KBgR0QIO8To8SgQ78WSAQ
BQIILdxH0D73RB6+wrg09VrLMKn5elakW/eFOhatMOajgMJ4BgKCvyYnYtetJiOcWfuLtheSE8DU
CAIhMf+VDpqb3RAeGsza1TVuCllwJfhD/urDdY7L6CXRR8JgwEKALgqfcUSlT9CitU2Af6JJ6x3z
5L/nVQhNmP4IiBG47J2mHuUxVl7q7S9HP1mBSKWBsCgu2qPBzDOKX7r/fXp2cqr601/Xiy6Y6R7D
obymZLOLZ9YJcRmwLMvACbCqkcR7ldL4rZIiaIxfI2zlllpwm4gMkdIepSX8yw6Aep0mEEuGxVMk
V6s0L+X7PPusQjjA4RqoKXn0ISVgu7HFS/MClw/7NlF173RvWBlitfzySQU2VNLQPrXJRdrmCepD
34wc6w0mEmfV61F0h0eJSPjr7u4UBNh2A13R8Syf79sav+8WwlkYXqg7OWu1zAq8vJfkUead3Epg
JXEiWMALiBdpuTKRm4yLtLch3NNQDMBaD1m/MlOSFSjXNGi95O+s+CFogdvw9Tp4KXqeZu3Pq7t4
UftEq/BzP6pC3F0a9q1GuHXPreupOfTTgUOoJGF37zbwXonkxzl33tXLp4JumFckYDK0g/Sl9qB4
PYKvv12+TOzh30sXGWsbjKYbrbjvjX0gUA+HeYpTxvemzUaMdufh09Ws+lfsFKMZ4+5m+fAFRUcm
sCIawArqIQXJ56MWiKcIemjYIuEUJ++sW9O3Lr1bTp3D4D6JUSZSXxBhg8kbAXdWJQ/dIhf+nWOW
HNT4GiHBcvYAccTZkhjew8XHwOgmduvlR4V5WEaxLVnuAEnVdliCptObqjD+xDfL5F9GTC6xhFWu
tIWQniBum5dwYJUeJjbiGJagbvUn9KOh6W7kjH/wFWhEZ/udgA4FslivM252g+UM5HimedvqdATZ
BEuM5nc7uub0RvONS1Pi0KdoKRanbf/TEn33vyhlZpNno+xOf0ZmD+NRm/zDja7D0v1PfsMZMCZ0
FSEJtbh+o/BBSMMjk3AjFb/t1KCPEjqp+djgcuA7j65riQyG9QsjLTdr9QhS8KfjvHBffjQFG7Xl
nuKRPelzBAVhuFHVrPmDLRGLSYj1wEO4WTJ+63Gktne1KEjOxKhcAo0kvNrRXnIYwbaVpg/k+oZa
9aoK5see58BcyZ3NVCYtQA1ZfiWkWPTL90qTVVAg16CRIRtaqD+bz0QHXXFLal5ba0t+QEC5R+Nk
5MQZnvDPyGHKVUh438MmJSnLAdJnzde7J1uYhFC7i++3lFtt3geFHqqGU8O/1vvsP6UTSy7GovaQ
FoYGbPbqNK408ptbHamGw5/rNwx1evZIeuhUt7xVQRMh93Ufo4lS2vXLd/mV1ZxAqikIZB1GGA+h
ZTIsYMDiTOhtH8d1G80hMC8szrA1AJhF0CiAsLB4gMO8ekkFcl5U4We2L1ld64mH9V9Hqs/UNv/Q
yM2vJmkprq9eDlZJd+DWt5ml4yLzR9f2QeU/rYjkuM7N4toTLPgN0wjFmwIP89RKyKey9JphpdTA
6vMT3Q0LiCgiHYflNrmBoh1UfSadArG8vOvPT4WGJTfb8Ob6/tQe3l4ijHwxYirjNIh/+Ek5HHwt
7LzTvSkZt42aYuYRKlv5A5c+WEabjTpy4QLGCjPdtPYMDFJW1ndtFpGvpoZ9fExkr/g96fiuABnr
m7WN7MXc4rtdYiCOikQJL9TbB4Oym4uy7M9A7WIUoIRd6ebA07lftXl38nFrdsP/ZhxgmMBuVBlQ
P5mP2O/gyQZ/ybcmE3lNoOx2aqnX3UUxBZ5cSX4BnRzcwK+AXgT8I2Is6g9gyNF/snULHn5xDIsO
qz9po0cN5+wAQJ6EkMHh4K1qHXkCh2PpJ+Og/lvo+RYbIcfyVh4lktGTSLFGKYaegFA4G4S63LRJ
eNelItNw6UJDd5n0UN3CLw2sdGYaYE3lxXHqfSW9AXVv6ApzCMyplTpz9CRKX3Rpm6bPC525ax1W
OCNtJ+MaVuVcWqcSv13PifPXLhBCCp/xM7w15KF+86lFstcuKcidkthT3KXddQOwhbrCoJRkYOhP
SBXIe8LiRqR4C3VHJdeOgTJmAzAILin8TF05OSKDza7nkE7ShENpswkrxiERBaKauzLYYWoZ5IaJ
dCsTvZPOOCOgVegcpH1jd8ZNQcJ9S590sxJ7nD6fohDj7S1eQxJa0dJml3hwfMvPlsORdvLl+Qkl
HAaYKog+LUv4BKWN/JfqS7nvur9eYGKVylFc189vOHlndz2q7+eDanMTUUxg6Wetuh76HC+GVs+t
3V6U/r+iwRTPJfN72ml+9HkkmeCcj/DIuUQE8jh1yteb3TW2QJLfBEo4Z5iptKb05hmwR8Pw2Ghh
MdtNP0oBZJUWkks1nnTzFe3JvFuvVWT4Jen2xcZmx2J9mkfBjUd14QZNplOVPUjCoHic/aQKMH23
Cw3bfhGntK+A/LeIza1UzNbd0rlhnBuVPrq8e1G2OY9wmb8ojYQJ2Sw0UBPkS2rCdAfDNoogQAKw
hc21q09GcMsesPM3TZH3sPKQ6XNkzu2iU9TkSubcZDTtflrOup/tOS1FDV3o7GR97AMCqiACnQo2
uXCPQlEjl667xdfb0T857TAfPstF4g6NlCkXtQyhrswutDmj+uYX8zJqHP5udWy5zrQX1RrIRMGS
GhpI0PN9nP1Qmxuyj7GO+X7cpHzTV+hbu5z9CasCmyEUqwPQ19XDurWUk+IQmLvA5aoFQZ9uY8Xe
prFzYitCKFTD65W/wCobMboruQ1U7T4FQQnEMkdGv16z8CeI42sW1dGBgGm2+NTtKDClVPzecUD9
NmrTmN3u0hOst9hYCwPEADP0pyqZqkh8tTA2s4PHC8TErfteJoI2X3+rxoaWs/7MmZGkQsSaRHuN
U63xaORicogcBaQZaf24hx+q+lp/rVfkEvABPAYqFJYjs3Cf5CzjXHDaHmQs7svdDMaPNV7smFJ7
6W72xKkRyb1Dyq2wo3VCchC+0a2sKSRB0XhCnZhVy+vt5nIJsrd5A9kIBMbvjGRUmb9CWhjLJthw
5vTaMvWkEbq8ckOKk128t6x8t3K/ORGmJrSW9qDHYo3qaYH0X74byX3R9shcwVu04PjWAqFvf427
F+eLNQ5DpNgA38hC5ms764LJOKSu9rcpZFOoope+e2zt6yTRfDmVj92hn706zCwgi0890AQb4W2n
/2Oi4UWJKgbRVLSteuomgG4QY+Kxx2lY7HSgm92KGY8pZf1o4uOz5fFEaLEIQdqy/YJ+94B+VzLV
6ISTHlQ8Itq/fL9qoPY9bx/aJf78vdZNskGhy3njDI6yTl91/9/eokjqB/PffwEt5bKKZmXSBH5d
kec5bC9i7vRIoTbQm0lQjPkl5qwI0PpS9h24mTuK9nmNVxKLHAkX+MSCV6GaxcnkPp+MFvPXlfDK
q0SgaV0cMAzxZaFGLasLXTSH4dXOggkAs/ltYRbwEs25exxisuO7IA76VREPINZWXCyYP9GRMkA+
U1WRiI/bEVsBjLKuAcAlwsOBL4qyi/FBRwCwlg7wl79YmhuXfENhxfm44nyoDTU6r5sS2cJGbfEH
B9euufVqFTU5V4V60W/5t1f4UcybFkNLE3XFxyZ++lO2fg9hEs6WSViCcn91Ik+loAca+7lQ7ozx
qAwbVbwZqi3SkaXl+K65xAz15xMAl17cF6nDxn2BX5FuBLtL4eYnolLw7bAfGA9BRw2XnwOs736T
8SV/L+sJnyqAqRpA51O6nf5pCBbvwYGgHCzVY5J1Xroi5k5QT3ZPBYJPY90Wjrsth4H5agEY353n
ha/OcfNBI3oLcF9td48VTDxkdgvt3pq4mS43LrXm7yVYa9P1rCpJHjzwjTImypyUiSvGAE36/hhn
GqvXbgjGP2llvasZp6cRnEv1ORaW1gqs3s0EmHbW8bkv1gpFkcJil7HhlNBF0+1QnADA4NYXc8Gy
idWtR5w6AQJLwbSFBGUGbtcZfx+9yvvo6OnUbPABDGMW6O4tLOPtvGs0kpEXnC7HEftOb+DwdJbx
JktX6hBvF+1+SI79pBpZfPohbtGxyECTA/iuiRG5Wt4CRPSfiF2fPjm9BOZOJqgIkAXRLl/756tB
8pYZm84HAJvyCaC22JrlgNg0VM+F60NaKRoHXoCg8lDCxsL3R4WummaE+1kcYx1vHVvCWjO52OcB
paVJmLU3XGhXTn5MSA2ySZkLJql9e1vYqjVWILLbdtVjoFC/+H+WMC8vYFQeLK+3tYNeqBqtQyCh
+vWswtwoFHgXvgpjx484QWIVAYd6rEXXZXQCpbSS/jW4hyPfatJ2lfy7uzPCBiV2inPvZ4vT1pPG
dmgdr3L0LvLplVvQ2AlfPjpNmOQhHBN0RJcBI0vtVtlAuBk0hxzBHD3bDHo4xNciEWQ4x8fF2X3l
e1+QM1/hm2bvyaGW1fJFyhz2lbLKMsThIDESCp81JwgieAcl2RCgIdHp5cLJ36l02J/+RCJNhUVq
5lXe0q8l+thscxgKW8iAw99yV1XIkOc1jV2rPb1RS2o4SsOBssSYrGgWdoBTLqUyYB4YxtLO2nTs
YwUF7cgPDByQRUgKsanqnRwkyq4q5cJAxKSwMkBwNVbIrcxdj9C5yDelMpMbxUVQ5iH6gIQ8jaqm
bng1xMUrX5zqNYjvDM1k6n6cKYBStF6dP9VDytWvkVM+42u3LqVam0T2265FwbcYUMhoHwDjHsXD
90SQg+SNtZtg+O68+CaYfNewHY/eTedm/3uUq4T4thCzm2VFwQLDaI1cKQWjsuAr7Ar5kbpDEZeP
E6yEjch17iRdo2aU65smazuQRjOvp8OXLxX332g5/d1doalXCsZTMGPCkqul52a1+wpMTpUAM1gP
qMeP0TkMCTq/O2jaZNEE1+X2ZZnVTX5gtKB2QJDnOOvEMe1L6ERMdaGxTjWAPw5O4/3TSJOlprYB
cOPmeJgSrh1TeG2x1MgWiAsfGK0K6gYe0CUzyQGPFBWNIsgrkJddJ+dkFcNIw03/ULiUQhg2l3r9
JpfLYfp5DTN5Un0vS0HtEDzEi4ZfAxIpCHK3kilQ/vRljCodpzEmMEUquZEytvLivFdjFs5tks+9
K9q7qdhE+AA1KIRhvi65rMci46DwMLtuRxapfp3S0QDN3DQvklQ/XLEZrrUrR1qy25x0dqZilQwP
oHnIqANJNmtthTB3yrycnxyJRaIQAo3qt7FsZMnN8RHGb0AI4TYJH5yCe0vhAFrHAAbOKf5ei1Cp
it+bU009TpU/PoXzVrYahxN9iBSdZqqx7yHS5GDJ8GEangDJ2DzrB7Uu2CmrQX7GgVjz2NINX1Zb
TFV7tFqij+Pe5dGrfVweN6APL9WEcGDqGu4lXAD+FidUYnRAVbyOpybo0DXDpzURgeFHk8uhWO2D
YKrCPUXXwg5EuJQX5JX01yM+IP1O1dQThQKsH7nZ6Y7e0KRD0hS94QVD/MCPtaD2vhTGfBwGrmq0
X+xqfij6GXawWSdfOuR1M5hj4f+evAC+N9w+pK99msEdDsr7yYrN7xxJqxT8qWJtdBSd0xnUU9fk
PTLbRBEQcW2vvktx9MnnrmVB1zfSfdu4LdsLFlAnCcKt9zmf1FBZ9gsxB+N8GpYk0XEe4UaPpBhr
agm+IyqsGRGKlSQgfJfgfRSYzwA2tZveRXguP34f06cQTTEUBJQ1ArlLNh7R0yCNiyYK9Xcqf2JN
XNbsSY+6ufVTDTzr+qN8r8n6jNknwIQzxByHmr7P49OcWSMgWBHaJRZhllykTfHmX33V4wmEP9JM
7GJrydgZ8WpSWY2fTwbDMbwRfcg14nFrFEBlpohZaF12dvDTNk6rNXnKfy0BAFSMT1IHEBvqNMlW
Nt62ZoTkCa47fgcCm3oQxukS8OMHvJEvsQtGLMpUm+56cVrCh0iokiwUXPYjfsplvtwxw1mStwAx
5ocv2+xqPG5EmsEzFZHTzBAjfNTRQCHm1q3OroiG/zEJzyacSkjfBo6+POse1Fd2ZphzOAbrgQ1c
DUMeXJUqBEtK1C1X7sp4YL32mXVALpkS7IrB26Ud5iutuF1Ek6+YNR2KXin9h3oSJ82OdxVeGPhv
Q74cXxuutb9Y4zEGjZaEkKVxS/fYlpnAPBmZ16UGoe/zk5IkcQ1Kg30DC/M2+s8ucCJK0mWcegWT
1A0DbMbnwX4gdbt6JdvLL2t0C7Hx/x87FswKcvNuM2d1eCDslCXu/FHbPQEeU3v5EEukjZ81/OIs
plzwwtE5Ei7IZkZmew9CW/U92ow+A53r264HP0AIxfDIU2YmCMLSar3eXhbdbWpA5+OCdgBHBTtw
PvgYwjCdtVxmS0o72Ub4DbXU41g3jD8kUL4h8f1hagQGcX0MgST1yykKPJ+ydnLHhj9NGxtC5Exf
7imUElmlUfXNoEcACxS5ajjOLub6os10KfQGTd5IJSknbwRoO0siuaupoN2dDRxbzob2gt8Rkodt
z8g85djEB6jN7OofYSyKD7lL3BexGGUvFsfEJgxoBHg/tSMHxR83/fSjksqxxINcaK1qCE31W24I
jNVaVGbrBVO30jLRb37I0ki3TLAAvxBgwdfx9rlCQyiIiNWJL+QrJC7BSMsFadjHsgxfbjkzGcmV
Q//8kjfJXXSrKb/tzlRGf59KuK5SPHz5QCYinYONEHlw9bhSs2NEqXzOyUiG39EVHj9k3Fnw2Dta
rUHE5hjNszfgPXB5xDafYtIWletT3ywUCkyhm1BjU/B9xAMYK3J1N6ttV+z18FxjtvKw0lEFsDzl
wDuOnwhT+NT1V3NmK5bL2iX3N9CYWhdq+g4pJK9P79AzMkTPzFKYkz7WR6zok2DPYWe3s1aFgTID
LzHKxRGJ5w4hzlprkdZeYaItYxhYL6mUzrydbTZhjBhQhuX1RbQ9O3ntIJwzfurgfKkXSYrv1+BE
HCr04mpqTMaBY1AUOHcox/hmtG98P5CegSoO2xp14oHnGI+7YoaUt8s8SbhnwQp+QuXX4fITwOtj
3xXu1S4tgQzy3C8eZomXbR+FR4M2KAdVUbnUE40o3qi2dwNKecA8BZJwFS+Xia3Pdc79uEq7adDt
hjfoONBkXjNBqNL5xMtkyPGswyh6LTWhM8Adg8lafpyMoomuQZE6XooK2XoIVvc48yITXKb+n3Jn
wOo9rmPiFT6PPnOKOJRyIEirdn8EHDegtUumfiG9huflU207KDiwe5IjIWi6EvJC67qqkCp0QPsm
sG/RwPY7R27AEYEdxmL/8Ls31qpXH8szYUOxz3i50vhudctgKLRpZMcJGrAE68Suk/rRGwK2JE8D
abSfvChtzlnuF+QsEmL+w3A3C1nvrl9qypXoxque3qRHC1fNB1cCjMCT4Rcv1XQ/NeWMXijxxvYK
6mbeEs7CUztrm23XFGFmN6PyHRKDoySfIpJfvm+Lva+qHX044ZgXbVuDxggjeOyPYt2gH1Cm4n35
jOk7e88VZbqguSjhs2V6d7THqUbm1JKQBL2z1ir/fvbWJBWxXWSn7huwj7I6MqVFRltHgxCRq57o
LuiXuir5OQFSKn9XuaQGe+M87Za4qcmUFQIiGCh5/WeplA1fJYGPC/7jhZd+kpgMz6Anr4MM+a9m
BE8wUVIj5bMSD+/egPmS516H5sJtsrbXeHeAqv12MlT8XjSxuFJBH/j9gYb07djx+M/O+/3xkG8h
D8pR8Vun/XdnB9ignuieQqQDK3hu5qiW9FJzcz9lM5axnzmTbY7XxtkDX31y68YiS3dqWFHzqZkk
Ldfmc2BCxrCP2eBfrdEt1I3ZQ+U1j5L9ByN+zAOaYNyKNpfFBQkLURQtiOLIFOFiEBMRJ9O78InS
BiQRh2OcNpiYeFi/2IJ8Cfg4FxeHqSK+DTArLZvT/KzFFAVKpFWtZyu42+iE9/sxWbeYi8dTEfhH
pXagg1DCnisjfGO3H4sSyfd+PJ95OP4RNuySi9A1JwlsrCHngcZolia0eQZuicCoOwvBI/u/0VNl
9T7JaEdXg9DC5NevhNWwj0D3Kx73yenFFKiKC+Qg/x7YMYgicNI75qAHIIeuWIMO2PpCQ3qtJaeR
8vLVj4/LOdrzTsW10w2CzSmLqA9sThWCMRFqMcmTp4BKIGnPKbp5P/6X0LLWBZtpTmozRj18iX+v
CtCBlmTLTGo3jmRSxyYrjVzv2L/io2uniYLw7qVjfChFfbm6sLrU4dcuwFjtUlL6o4x221LCFON9
ecy4YNyVEWxtinh7cTncAlAkmHSuIxdL+WPUMGp+UqVjzysEWWDsyzKJsi4RidaNmJK3Uf5dGmuP
iOA+UxUgVHDKlFo48SzDkLcCzmdhmXUFlZZcAaUvT0/RT4Txni4VW6gQms5clUhFeNlcFFQ1d6G0
6L3hB5hFmD2scNQvkaLJkNo2/bsuUTJLldvZ3XNhs/LEMX9l/OdM78MLh+/Fy6v+/6OeOu5pQ73J
Z0VFMsdAbBnB6OvNVxA8q+8A8YBiy0D8ePQOQa7Xci89Al8H21YxALpq/QDEyKV2InLl2pJr8tGn
FnuyuZhB4AtuEUk+8vxvADnroaTrVI0RxfnLBOlssNjTVcozMFSE1g7zGQehx/zRGC11senYRUqb
BMeMunZAmqUWI/Cghr6NM8TTFfKZ0IC1O9Sy/Iby71mU4iKlaZH9yBct61m7T52AGKP4KeMt7x3F
UTrtUcovVH9Xd8XSgf1WN5phdGgH+7z9Isei3OOaQs9DuVkkDhWSXBUFxYwufSuDLvzWHlLKgTzH
bWWpGLgkgcdy382xss9lYEoVUsi+gDHGo15oCR8h4fhDzU8MhWgzVmZhPFmok0W7+2Sf3wPAhb6f
Hec/Hcs6rKmwJAGKAt/nZ3pZ4OSsBgwSHvlnSCofcXyKe1+LLTqFvax/n6StqKnykn+Gih/5BKCf
nJcw9EIKUfJKUUnIz35kJHeEPcfxPh1pqMgrADKHQkHIP9YF/Howmgln4NjoEKztqcxV/NJ8d0MP
6VlAiLW3faE6UWzAA4JUVWNzSF9tZYuS6uxdICK7kGRD6l2VtK7Vf1FhHsLaonEh4fPl+gAr+WaT
UkwF1LZ18uTDPFiLFX4SVkMT/n7prc2ULMQ8zmXhRNHD4K5z0Fos5PMsWLzs0dfaP4erBjYxVhEj
nUitWKUlmk+7zC7rOveULTTTOzbpu9hETV0/Lxuchxy2TTvOvPnrZRGh5Oc8MjpBx7s7f7BbTCB0
aG7imMlutEEKI3Ovg6RYMc+PHU8kIzLUZQLWM6cRMuqm4YkDwyfO/OhtPBHHLV17NJ4rAj8cY7M5
mcqweO6fKj1rGOs78Xb3bugbr47n7HUl/3tsMk/DVqDdU5x37An9/8L56hzX/w588ovNNkwE1/XH
A624NiC5ZSIf9hIGalXzmFw/68k1n06U8FgiV10Fhx9zkCVtxhbiXUw8YqMWPtW/gzYgHW9QH3dL
GMM5mdX0KceofY/0ckEnGJs7BlG1FLgK21cnyQ/a84sInFfrI3ectWqOf4chIcYkokZcuHYzVDs4
Qxoo+XPUr2Bk0rSpmNSRYZmEcmzk7LXdmY9JrM0RE1NUEQfNdHpgHEB/4MyzqtoEEJ3tnBm7MEoK
OJBnFdwn6lbiMj1A6wyi286/5DH6wkKb+5NoBDRoJJyf8mbzIRiiQWpE/hySX2J+HWgWDkQA0xSW
GIFBTSLU1AJBYD4CmNrrUJnYD7wdFco7nbTahAhuj9ovgGoeP8G/M45D4LczoRKnYTFuX8VgfRtq
rtN2uzeZoWdLP9yq3ra4KJNfI/WwiziDxPoJTvA5uhjkFxN/yPLiaDfjYcKPljCFLqya99zcmy2F
1hxgp+rKLSZYiD2YC5ua2XMfDg/CgxU52vz0YF0c5QXWSISSJKYAiJn0JmT5EABTfHHdq5p9rwRG
VyDCK5uQvVJ9QhKduFh9/30MDPgY/T/9cs1xaIdhW+UAL8d0Nu420DXwzGnJXUTv9GmEI8CuLKQ4
xPeB+ch/4OmpZLz8mleBjfMb33vU0nuhvbLFw/6/cT8Yt1ytl/4eQ7JOU3kxmwplqxoeKGE1ywxU
JSpVIE+fpiKzKyGhaMgJuUQZd78UIFSCf5dWRhMW2IuA2Atw78W5OyU8ePXRwnGowGnwBW+M7rvJ
OSkYp4KBym6N/g5zR7swR1nfm/kk3f59ZgKVJl0yYz59OjOM5bbNqwLYZ6GOGEQQqF1qtPk3k/qG
/bup/PHHtUH+2zuSharzk3ya0SdhQBGh27n3Ry26ZfYrwqiPkvyycE536LAkI0/KMOJ4bbLpCONa
DEh26WfpD/EVlMIg6y/m9jZc/a6hrdIp7HWdc8qOhZ172zX562Xv+OuVUN5zPVV05A9F2yv6Edsf
z+xtjfSuSQGqfUdXvhwY6+4KqTGIOIVzRBZ6itGZl/4pXVyTna85pTTTYn2fdWFBJD2CRZt9sjaK
WAxROP99gmE6BCLEjFcCVsmoGY42Epo7vmcyM1bjSv1Lgqs0L2ctZwbutR+pg4O7/Mt3OdJ6dcOQ
e3F5qgEDz3QgUfKw64XXs+qAdXfpBuApuJ+l+2LxT8TLlk4eJrlD28tT2ilRUB8KFcGIeNQtfKRY
3HQb94YF4krw8nYhfJZhr+UsGTSfNfSYyHqII+YBo9zrSihDpSMj8J5c/JV56tpLiowiO1le3X6+
H5lZoRMzxUr4LTWtPsoa8WLC3fK+AVRrF72M0WSer4FsTL9kgXEXvvZoO40KGW7v3CjOvv6VKCN9
RCC8jrEAt4uu8ZzFzQsuR3x8tuTiJJVqZzWjo8bTE2aud04L3JOBCMKUtzQZ9beSbZZB2fU3qKKE
BnObwe+KP1/4j5Ix+qyids3RzOpy3KJeXrUWPyY3MWE2+wc8uSUC9BnXS+biG/lbe/6N6wiAPi9e
MPgcpvoMGKlH19JTF2hS3T1zlRK/Bbh+ZiDmjPIXsMFVDc1TxiMpyTsDeBnzEkHXt/IWmJT0vslM
22qVE2EiBpMWg+k/Q5wLKEBRoDBUdA9nWhFLY8OLgjegEFWVrmlIUBFszo26C8ja66GkaosXtxtM
Ha/3y/HpGfCT/LgaJGkO/GrMaAOv1olCh4ee4pEIj4R+bt0YhKbFzoj0WN5+IobjoMR5H4ugBLXo
hSJsvZnaTHdYNYsz/YGQDVJAyCxiMIkcl6SkbqRbNqmbPLQCOhal6g7ejaHI2bqFbpUwViRM4Bwm
60pa1hN1tqP6l/cO7DHDBypb8l3WjvKIpjWjmFjMvhsvCYQRRfU6bjbKjR6eIAyS58xj2kZWeHG6
N46JOYWlstpHufPoVPpIhSE8OLdD2UCnuRi41CBTwsEggwlFdHYkm6pf4T7pWCvHHH+OVUDIylJ+
TKstMP1kS+DGq8w/oXwqj4koTTM0toaaL6UlUm+7LzSCs0z8YyxBOKbW6uFoE1YHKSBoPOY5worL
K+4uC7Kp0r/dW8sFtd7GyNojCHB2J+5A6/9wjKQZt9UyD79549qQRgnKI8Hg7IgfhI1WJa/s1zUl
6cJ9fehCdb61sWJs4RhtZda7L96NQngldJxCSCtxWKZcTG84qG+YldCeQy5YW6c/cXoj+LPDLf4+
dw/jm2MO6zhX7mkVN2cGPHtnAd1EFGMb64+UNFk8acN8T4udW/8hgaGpG+lYnRWLQE2kspu1tBJ4
3hbdwmV0sORQ8nUdG9TFhoGqu4KFhLlBg0+YNqMwzt1uaAL9s6R2cKGKy3/9RA2LBqhyaL4VT7cn
AT5UmNu0DyFq92k7qyXUE+NQWhQgnhzs05eS42tZDFFLBMCFLw9g1RGG+vFwYFjCKwexHB5bbny1
JKx8jZ3Ja0tqrslipfDkkO6jby8yYV5iTfdie6BUMKoMwVlWH5d5a088XY2BKqIVGOSr+3VMN+me
Bg+T6UanPJmps018JPCYNhHuBl37nJ+GnP0Fcs9ManF4SVbquwSNbaUFXd2MTxOItJBoYrcYficW
an+IVUjdJRDSqg6ttBy361y6/EVwIhE20BgqXS98pq26g4dy0uO+fzHG2PzxlhOcDzvQo/eZp3NP
AQYfkeLjbtzmVdxJTJZO8H9xKezpXwaZyArRrpG63oTteXr0ps0AqqrXXhGXbd379IX3/cqvsn7E
c/rwKG71e70dICP4QQV+x/UBCXk3RJkn1fIQ+uVz2frMNIm1yobU+EMqdXKlxHsqfzJi9vTG0BvO
SKjS/mZtMO1LcbcwO6DOLryDEjrOtvgcdWydeFINApI01y6VYQmcY/GaLE5TZZPApMxdPbEl+8PB
PM+XZn5JUrFC4LBasWCyFoY82Iu9P8+8U3k/kl9guEep9IL3R4Blas00Hm8Qvgd7niCg5bubgdJf
3JA/G85OAmhocXu5ltieB95ap/+wlfvRCwjARYqPAmO9HXLwIKeDWv1sm0HNQW+lppVnJD+YwLSU
p8rPLKhkSkgmHemTYJ+tXkbFDOo/YoF7GTQvHTQwSfv4TyqSd/c0BMV9cckEE1V0N6urNiCF5mNZ
5iobrugIo8zPJoriiQ2zNwNxI+qc9D9VK4Ur8NptGl8VtzquJpx2ovhkl4cbKYqfJTdtJpJpK1V5
h2BigOpTSLchwctqYUz36NPMQT5HNK+V38x3O0qAgbVq0diL456r8cUjEsttCcMfBKUcKAh17ByA
YCrOSUoieTsCBtoq0acVo2EKmnf9V4zdTzF+UPjvF00xmfvsfc+Lro7ydFrwKyhAa6vRmw7JGLKs
uqB0QQmr58mO3aMpukak//e/p+F5M/6FYqmfSse6ksdDRvX2bl2KS1mFzZQaHyE9jb8/E/m8aNWc
DrPVSULB5vgLsLAhdpGDqKQmSV9h0YsQTJCKb5avfhioBSLv9kK+EA9tyH3WrR9xMBCJVuIJiXOQ
ZO/DjsClyLJJoP71x3i/2tjqcgFEAy9+wVn98Q8awXwqExxmiunFpQz9eWCWnLMMzUmp8n3lN5Wk
7icIcxklLmJpdgziq1jukAAPykb3DiumiyWH6AG8Xvts4GPUiwdqwUN6Qfts1xAvYFXAHQknqV3f
yZ6k1BKU2hKIYe53StukYUqWqk+mAutPLm2oungO24lNyvDOIeAgo3wgcgrKXEdEy+sDeKYbJW4E
GOGvxyDvhGZ6R5gVukcVsvU6CZcK732ckn4RPxawpFHpJcxBYaeh3Dluk2zC8jGY6NViazP0Jonw
4cX6AUlHcMbH0r7r/vM6f2OcyAPpOTfvW93QrQJe3OOAAq+/e1OI9W/ziCgBGXOZicFTDV73iBkp
B85hft09IWoadUoYFNeRHVDatguLHPd5lYuy7xfC6ohqcz7MbrIlJ9q9R8IXk7W6aQ+k3J/FUo6N
tfyn9YE6i9Xe1aXPyAVj5pjWpEPWUarJDz3Gkor7ATHmI2iTXZyxZNTqEs3Y7wwIi/uv2jOQxSSs
KbBiez4c8AHFbVW0Sn6Hvqs5YFK0wuSATfN78RimNYN78LMNZOAF0/MW5HLpfloyV/ihn6VlbC7N
SnlOUvJyap+1M5W7L1mZPvEHahLRQoi2jlemni8HaMVFi+4Vmpdktwey5hCu0cMmvewJ/tpxqaCm
0p7bB8/J2/4lp3m+7Mfiylw2PoY8SLX3KKnXbKRxGOsRiXkjQ2DJ3WrEfg4AhaaQoS/Rl9HH0dG/
yHV2mu6Q4tynb95AN/pQifYMWIA9ySVMXEjjcANu9ghOAZ5D/s/WUnTj2lD4roQZNx/gIx6o/0/c
Ju+dBVxat7ki/F1GqOA4PUgNcj8c3GJuAr5i8/mkwXURvARfn09JpA612sr7nnvfDHx4lTFMzawr
9K2kp+dtA8z38efSsRDX8T/R3toNNnnVozXMA7YuUplW9N3Rv4Wv2S+lKEMziE9lPboFIPXT5Fre
IcTFqYEeuDWUQ+zstwHwP8JY2WUX9vBlhX4cf9Sd/VvOQzzTTh9jFttdDSuf53Je6s+WTzDNySKb
3+3BJBi40oVEeQn+X9PIDKw/V7I7Nb2YzUWXYvno8/P9J5k8Ux8FlCB4CWtT5OJw1u7ZotD8vDNA
KUx54y4G8SCq/LjVxQvuh9uj2Kg0vQIEFceT0CBFNvlWH2FbtzZ/t/Kg8yRwxhpkaKx2bj+JljTL
8Q3Xn9IVei/gRMkaPXNGrVR3DUuYhBzitQnCITQQeNH5JswETvSt/8uKOKGxi2C68GTKPhlh4wJz
5S3V7zTxE9HLaJBcSVdCA4H4aCIKtiG131Cdgi4dyVMnNjY8xv4S08duyYCBYiKXuBkut6p+fyXX
++5z5EKeNfT56segjfPzDhiZjwKWJP4yvsbuPgMRmy3XM9pgyNSEd5vQt8w5R9NsG4wPnkcLfmBN
Cj8Jbui70heUHdZCspAW6TOE3e0n3JbsqO5XlFXw0kRf5Ik9yw2+G6et9JlF1s+ApqcSeTb+meNB
9dql4DaCgVWG7PWO2vC7dGOYM/99urmwKZDKJO1yuA2YtSrFkvV8hZ3wBNxc6g7diOD9f3lojy7j
JcOBPFikIAZ0JO/clgp8iBthu1DSVD7nBL5us9xURwXQrwjrjHxqK+98ACrkuaUXqRXofIC0ujF3
LF3iPBOr0zUuZVomSbsXPxef2i36Yo1iz4yJSQyz+WN2+NUvP5uynawS7D+hvhKm3NdDAQYFWZMi
yuvn5wnf3YkXsLNZ/ujqrw5y3bnSQ0eQrxJYlqyZDSq5oOJoVavBsvO/yjdRg1gCIH2E9qBrEeXh
0RYQ0N++9PCzrzHY9SbCmVsEqqVvbidjxLpaUmU+9X0KYf8iLE00Ub6xkdy2cJOm/POEYZfIC3W0
L5tQFxWuvymQSzXQCF8a8MmUvjHiU9A80iL8HxlwDBxaqCvTMwHsLr4pkly7tcxcxmq22/Af2M3t
QnCChiaqlKtBQiaV9+DzvGARhABNjardZRAQFlMxz2/yjf8lPoG3VpdCo+M2JtYH+Yeu/JBISM+b
+qEaXYJi9zIE37TR0gwnuP4dENR/jkicwgfNkncoOvKYqQKBqG1yczeUxJ7LQ3AoB+JNKa1m4vGa
6Kq1hDn0bLGj6Dsa25wAzrkErrUacTy0bMrTNQzD6uDxI5kWTqam4PNGHX2Y/0xc8zsAhzyNzY+k
e28WT1PC2du5DUAksW7Y9BLZcs4C+3zA697zrt0dtIc/lAnkjjkTw2Sk7ONhzynDV6JjVpSvW/11
rvWeAVMdL45cKkcYHXF+RW4ILkEBcHOPH1y5DTiQYH+WTCF8EFCjU39BUh+eAFozwt9JPri4XTMT
gy7LGiX/lxVGmW8p/SnuzN+He2vsvYJNMPPdsT6vQjQE0kOzB64kr3tRaiDaJ0hIVOfKJxc14BYm
7AJLb9ldduT+/1QfsXHjPKalbxuUBbJ1HbVIjfy6UxDRVfSQ+4TuB9V7409CawTCef0JrmM2A29P
zhpeNVG54+MTIm74gzp8xjoLhY8DrOf3PMxUBkBkexxJpIEV0UgR8tVPhWrnQarJ2vRP5Yqet48q
Deuj5fXekK6m9cKAkHpFbbISg3Vdd79bKUFvbOJzGmiVON0FMUr/MEkd9/GSjAHlqpgfhdF5dahM
oBi3zHBpZH8MEUQntu/PinBOtrQnYE4FUil/MMQEDOiWoAe0yGwMFmWumeR/jC+FtLwAlLtFIJBv
vdjXO48OW1hbe9Ghio6abAHilF4VJWuxsIHEGmEXgIedbelCMCCLdrSiIosXHnmU//pEvk/LxQsP
YePl/Kz2NJEw0u+PFuSHUBJdL1qHvTEHBcnkSE2t+aUD+omVPEnHle194Isc4qFs0+5jaKsJMJRu
B2aEKLvbnbVeUow69x45Bvl+Mw5tuDL7iQb5MWPgdNxkFLdoOqpPkRKPWqf3eucW75BSmS93iygA
eXNPfNwphdmUrGACk+pKE1NC4L7FeWQvVYS9ox7IlUKCq0FGuy5JAMgUC4W/CtdxfAFLDxvhgRC+
MCss+5xBkdMtfKG0qxXOR1CW9iyVaczpJXku3PL7NlY7dkZ0OI0UjaDCiGwoB4njCch73fDkspn/
AFQiRU+Edez+4VGOapJ6+ggMSn4b2AFK/2iJWb3qO0HU94S8GxNvwhzZyAj7yVEVdCiEdPyWIrK3
FpGzR7K/Hyyk6ySeSIifsxWih7quY3DMFT8QFD4X67xyOKH2IS8KH9AarySpaME28FVpznaBncZC
XrNpHU41HESYw00yCrAT2DQ/tM8uK+xk+XZpDM898iL2g5jZ80MVR02mLaSXa0KAOzFDDUZJiQ+a
2B73kaczXUKIl7mw4Xa27lTAu5JNnjz10c5hrfEFSZcJt5bNT50nqTJG03QknHIJr/nGfJQy5ENQ
VyrER1E/xhzpfFE7CJ5udg2tAJ7EM59N368H2gdDgb2DwYpjx9+4oaxAw2Hjo3WXE2U7aT/AXUlT
L2o1gDKdtJcrxWiYf0er9PjgRXPphUuNaSoT1Lrg1uttE1IvSAN5n6lf9r7+wJkA94tVYzNeDue4
07DjmD/eXx+I8GEcaX7UYQveZid5wCPHbG++hOEpKQcfuPnYmd0ap+dCmkb2zCku/NTw7b/gP1DG
hGitWANWqQ6B9U+5k9EJkBS6m/5I2k3SJLIGqcba0fPcyjhoowcFkZITsyIYEFd/1t6wzeMdWZYx
0N+788HpiBt1YnLGugXg+k5LFTIfjti/VytOA2pT9MUimQku6rOrGRbtZ+acKZyM8+zKmwrfFN4+
fMcHVr3Zgi2BbT9wbgV8oHDp2KR0yyc/C2IthPimdypG3hL5zxCoF+CC3dwhgFJ1y7GFAsNU87tb
n9JJ6ET/dDleBruTbaIJlBb0Wgk/W1ZoIcJRlJWwX8BTO+FoNXwkuvfBaCNdo0uJQLPQAqD8LOh1
5UawaxF5lcfjuH7+oEfmMWQQiMJ65GyyD25u1wP+K3QkClFeroBJGT1+dj2fHltyQ6VIilyocBDz
lyhbKz1kFkSM0QuLE0Jw624MQYpyhbsE4xHfLv9+hX7CqrmOgRGaxc8ZiLIbcUXGmDwtXnw2gZ5F
BHeFvWJ66VPIZRxgXcjcaCnIB1PL0zwha9ZllylX55WrcsseL/gG+5yYKS12ENjOICEaashUHHfl
KO16+nHKFctnZk/m22DZ2gAzjF20WHGvVUhZOO5hRh1jqAORte+tY64woXl9yVVmv1P0mPhljVGX
c7f62NZIHnoQin/xSpARecwV7peYlcHmixSExI7Gkv4HnADzGs1WBonx4M/dv694S1W+Gc90N/KA
eBMmODivt4ND9/8NSeQ7vG2ttUp1EAmljFUSRhXtPK+ZUzVfAWkwYffgL/tU2ZPVTrVgt8cq8a5Q
A25Db0TlcicbchqrNO1bvfrABMCY7OaJ3Oc8JCE7gPW6+XguMfcC0LIJizpT0HSdixSFvtbx6gH2
Q8mUWn+CaEdSham7WAHzCUdXPkYMSPMkkDX9+SwHOTaxy1vHu0iQphYk+cSsZk9pnMISUHe9PgT9
F9QaxjMtQp3pkDr29dYf3evWTfiKlsN0DgJyOAPVR+4bz/cnxHOOXeuiNrs4Nn+gh5ZYCLtowc+y
7PWQPD9WHWefcDByT8TAKKHT//6uDI8EqKbxcq1N6noFU2CIl06AtBexFSzekhOtjodSwCwJ/pqM
ubN8Yx7DxGosgz1st62uKmBjav+1d93iafoKWH4tH6aasMy/k6TG89Kl4SsdWpqwBANUZssD1mZn
c0scpNAxD7AjXPPhSDhFHcShZ1dO0x0X5qc3VSdKUkNUhmMFjfwF8LrrI9h4+dr0GjJ9nWmgXBm3
QQ+NXdf9/8SELMETgCIvXCIXVESlWPC2hRn0LmDN9Au2MPQyhUM+i8UKAM0Rm5Aj2ftyXfnYAZU3
toehfpRTAPnSkhD0QLSGv/TIVU2wrLocoRJXJviBhckRATGas3xMV3W+A6eEVCXpyiFWA+DCFlV5
Qpf4QJk6mbMVFW5LgpVu56eGbS/u/Irc7HADuKtP8UJOJL79MkvI69qAKaJQ3S+EnB+N4jW5wiPG
6RuMk/crfGaiz6CRXm7Vi60GaWVBTfetwbJ8Vtjow1eRZGlgtiPAqhNPpBoDKfuKWTNywX8IascG
GnjiL+apXBoCHrCDAK6xms91xeG67m7vYgWlrlv1cTmEd50UNyXnf6ThcvGOsSg+WQ1FJsbGTchH
7x/nz04C7Qmq1BZXj2DCp1icLh4jyYp7/yGrOrwgAHAx6B0F7i3fKW9gZ2nI4qLj0MuRTYkQRIh8
uK3cvQjNnDPl/dJvJQ1Pu0KsaLmIewFaHQY8/81p/AC6gotDupev7+sgUHbzQAZOHQU8LyInRV5q
Bj5APp6kwVu6Bj82dOYSOvAt0kF787PAjx3SdHUwFopF9BR1D01ehsK/QCbR84Pcz1HyWyVc6H3Z
hAi1QFRWcf5wEpwJJn3sCOl/1ITGdAr5JAHaxQ5/3etp3S53q3VchiaNcNfqSUT5/VCdHaV8aqaw
HGeDOnB30ACQFIGNqNzhwWNtOPHjTo1RCGnQ4vJyo/+SHKKw7QygE/BfyxscL6DrVbNYLi9+uQmU
ZU3j+qhalDSeziswMIwcYRu9oyEX7ZqLN1wbilcX1WLTqVQV4rIouO9x7tX9ckaa5qRNlvda7O6T
E6iYFwFMnD9SYqfS1HmATP48uCatEIeJxTwC2BF2Dj05BAfkXN7ChTdAg6kY09qpNmw0y8q4SxSy
0ztwnAsuhYCwk5KT1schrYUffXr04Iq4nmC7JDQJGZZG9QQIl1Hmt+aCvQ54zdF7yFy80hkZvzjy
QTA5ajtXXbvFlFuBjpXxb2C8vaEAr734YVsWEK0wA5iLnZqCa0rYYDvGmAm5J2/wjbs0u4VUZzGy
6buCG28efjFI8oss0sJ5MxPFGN8yP6F1Ep5CXC/a8515xaQlKQTR80yO9LKdbWgZEZKkx6h3lz47
WuCsQugKoraAKynOhyGvpP3+NW1iVjL56r3z5WAUESoArOz84CgY1bPNtQfcwdIrh0J64Ewd2KyY
6TKtPe1XH9L7FpK7kGpHIX8Q/Q8ipwDUngyrZChOdrbV8aQ6tfznCmnWKsXjJoB/pcghcdUGy1Ni
lbBdIwiRV+KoI1lbQup4kqhdq+Vu6OrjsLVYleCJiSr8x4EONFQ8xYx0LtcnqC8lqTWhTIY04rJ8
7JanxaI3LwDF+TCI/NtLJ+maT5Qa2DJJBdaY8woxl+SMZS1P6PuiBnZ0GZrBnrhXhHIk81iwzdil
hdl+maSpSitZjBlzmHKX4z6lYts84YbeIsxkJaQR+yYAdRg7+2h801eB5G001D9nCH7rJqkQ8ei8
nk6xXbO2E5ltQpZIi27oX56f//R0gWU/WJUAAvJjptFTxe6VxBmZ/nAMJWGMuVhHWJQJIkylY0UM
qQm/oiUpJQ8cWQVwHnCb8fi9iSGU9lQencu+5QShcT9oLuPws6QY/fMb1lLJBQrb58sB2VcLFz23
JLgYcJj2VgD/pwYptrH+zCNaIRXyddPAp6k7Qfpwxb0tKlI/RWXvd16KZAK1b9Iqf4SBLfRvdcKZ
6D066A7t+kIcz7Lo3mxhRiXcl4ndesv4eZ6/pJUya7W5FqR7kiLSXc698z9iWWo/NinYjroLa2Pb
khaCt7nwMiNxsX06zHGZW/W7GWblbIFU9opRlnmOuj9bIuMRazIxqqc5bToYYoHL1v22cc0jo4Yg
fgoOo1eaTQLjhWlbgSAZZrhDum8NqC6WZSk69sbZfz/WcumkY9x+x+rVYrx/gE4jiqxTkKpkmBVt
KYyz9LRXENfjt8EKIqE2yQII715Tm03eBz/5j0yS2sEfupmap6vYmQk4WLmRq2BU5T4p4qEqWoey
7ZqCN/b42FmMzK9PMkR+kiIVcx1u7vuMOHO8iM84zR49dT9QPXaIwOEOKmb9o/tqNebIWpgj+HB9
L/CfdSruDw9x0XDtOM7zyNNB1mCuwf5UMl7rob9I/Jrx+WosXKeRLTgmvFfB1N0PY5MtYtk/BaVU
e7rd0c5wkbyVypgIyJgPLQQGOvXswkJddZAJbhSEkvRK/iUzA8jcSYS7uEs511TV/PbAlCy2EKei
eVcKErbeP8S2RajZqPZEJO/t80O4+HR6FXsNt6atRF+jHrHSyR4lbH7qfdn4UhDJ85Gq87yb3kuD
/ExpzTfP5Q6KaMY/xqKHxflVBWn5R2h+EzlsDryB953c/cpu3wbx9molXHpP6zwGVqDuR2NkzHXx
iqF2/O/BntcxCNqbNMD32Kixq9NMXprjAVVcs6SrhOaQJD9h/TTMSRl71kPseA5htM/QM+mh2GaQ
zLokNg9rHa8xjeNxTORA9bCJEGz0N2/1fCyKAJ/TIAo6kx9790HK4ok0aZnGzlQdSQtbyv3qpiMx
C+NdX9JH2Hm7KH0JAMnPjFX5OsQgVBPwSQu3/1TpdcZ0Y0cIMj75goeuOHviv8g60mFS7HI2zEWi
G5hdPbsTy33+C57ANcv/iBWGvuo8x+pNJGShsILndMP9z9CULxZlw1z2i1vjedT9Nuwqqz+0tCtn
i2mqBmg0vH4g4vQLao0w2ssbAkOUtAbwaQaw/TrYNgxth3wDPmfmuI/KSWd8e0q1AsvLbty4zj7n
85KBh0g+ib+4Z8Nq6nU0UEzaf4gHuNjGDbkZrpc+F3PqWkhTVYpY4FE0xXikSVUgOkTAqCJcUs0e
lPKWznIP4kM3EfhE2rpFVIkqh4QeYmtUm9BEnQxsaW64I9lVHVSy++wWuDKwd9MoYR8a4mFQK+1N
vjWRfRO27CFKSrByS+SsKda49YSkEs9injlbluPHZVGnTbntUh9gvg4FmTnyNeJXCjoK1nVkconT
p1E/DfwDvdj7jal7O/yIRy5r2BI18bC364QJU+fr8P9Wh0x60fq59vO97QZyaWmIgPA51bg3RVjp
n4KVsflxEpEAtCyhAiI7ylPXEA4bUGbHlqvvk34HgBmjew+dnn673BJEJnppXNJHwNs0Aogc/mv4
P9drIoeDj2KXtwACtq/qvUH7bhfP2/FXAbAoRf86U07Bf14wd8Nn9rQGvJ0lN3RLwbK/4b7Fo8kh
ODhxt/z8Bjvg4HWhNP2hpAFqbEnkOYvoL1uWf3uDagy7hSPAxU0n4QcPNDxr/TEDIEJbpSZJbtUv
3CCFVTEtoIhriZLXYWGd2kicAF0Lzfp6uPQr2G+LI5AMG9p6NNjWDAa74qbb3DmEIF38zVBBgeRe
86iTXQ/WbdE8ES/wm8dCcE9vTdfmJbZotjp1sUmnFEbcVCEntlm0gpT+cgxU+lFC/uvOQh8mDP+N
HhMze9hG2HNy3dMWS9L+mRExWRz8EhI7sDJ9U1z0qLCbjFZ2WOvhs8eCobd+6T2xkJ0DLzKgwsk6
LcpyIY9sq4rxof6xbhUCVvKyunLSJ/36ZGD7vg5Jkth9dFgRGAy15tkJ5BxdUdpgLCgJMrfBqZiX
AF+9MpJwE7O764GiZLNEIq9Vp4yus19OBoSsR0VI4Bu9+bvGdlOYpxpJCnkDrRY3b0yt5CbuktoA
Q7bJ4nU2uChrZDW3u9+zEA4iiGBifJQxOC4jrAQbgg3QU21I5uibOLQSdLO37ymLtHCv1X66Ib94
2yMpF3emi4Pdh9JOZZ6ZL1NjOTrAKT1yQEAuwhNMuVuazkbML4ImGT2WBJhtsDRL7NZW2f58cpWY
340Q09ckbQmSnekb86u3E8VQYRyiHya15WHEG3trhaOxrG8rDrAJVH3eRLSo4HncEvbB2J/fwqwf
t+ihY9shylfC2wgSTut1Io5dCJyehToO4/TcqCwJGN9hrywD2s5H5n8jRYY5aqUG77DbFcp1Sn+C
3rohnNCtDbxI/os7uZCdvovWZIYcLq8mWkvXppNdL4CfJqbJADuortdlhEXdqsHT8Vgm0P7vqNIK
tq+/257siEfQymZmSm5lj+k3aNA6ZMeMO4BtVrbdlG1EpVSsJOnI4BqVSvaX6Cnj1lhSX/m+9zja
f37Ni/lX51Zl5jbQiHB1o0SV17knYCavgH+9f86LLN3Y5qiWg3YW31KEmW5tAj/aKxu4XpC0fJdI
yms2q/cd9OvxpLax4ZEpBhzQAJIHTVN7kwEqRsdC7xhILvW9Kq9dgxG23jarnc+MkCnbNuM8jRMz
VMFgR7Nf+9RUH4NSXLVXSyfYNp6ZjBsE+1wVoXvTdld5ujNkVspHI0FHooA8XSg0gcotBNek6Scy
0KsYU2+JfS8N0476CDfQBtLorcVw9GMs6LZmJaHrFyiP7ob7o4H4938a0v0sSD89M/7S1hVW1crR
ovN7l6//pxGFNcbQ9R40DZBA59+3id+YDxBJCkBzYIPdCMB5gcS2iIWdK5gjGsCj1MVShT8Cp/to
FR5EJ+jrV8s35BJyipBALXtNqCYGakQQ/Bf8tLs941V/7Vn6fQiNG2OY2/zFvlgX3huFm8BzOFmf
QxHY03MOl+ASzmLTvz6026S4W5RmcUB1+HCeiJSZVaptY7AQf57+bd2G8BxZUpzJopMLW7AsIxPV
Pz+Sp+Rbimoax1xAmBqgDPDQwUs9jd4HLX3Dj5hQl9GbsSv3Tq4gO9f/A+s/IgoH7/k1V/hq/ERo
IqweEZtPg2lrM7KciTWGsd3qy11QKdPoPFZfpK16XqJGs3OBxKkotg8YaIq0AyYZT8BRxJerzsfQ
9kYZQVRYRBjc1+wSraC2LlvXLbFko+UWFf2cZJ1HC/AbNJjv3Ko19D+rO2WYckGRyjso5mU+UgKz
4HxwrD6oX16/xFOnz8ay8vEK5nPpMRC/F/m/hQtwJ/DzOWsWuxjlAtaXiEvReoyALhGJ14K9CKou
iPm/qbH+okzpJgM1QQDvK2XqOhXLlwX1RcNeW9fy2BbQhiYaTaFSQY/CqCOaiNsu4ETmX80TxoxL
04YP8phter+sOe0iRX3WahLz4toGdizBK2PxuaxAumsO7hcsCSLF+vSEF4albNwm0Nyu5zeCV4nT
jp0C6E9CHZdga+U/Np0vz33Iz5PhrFgD3Ox1+4LE6nq8EiKqOOBikBN/GRTxfledHdofAYVGRY1B
yeGnx6K/vd5P+bzT0vUZgRRtstxWKjf3anHnYcOUC+tLV4r2e0A+/YQcEXNa/6DG/v+j8j7VFDS0
CAaFRjFjte3tiuECaM+N2DS/zIk++KI8q9z3d21SmU+Ci51W5NUrAQ9N1psD8SyV1+rIkjxLeUi3
BG2yZTSXX3x7JfQ2Sm/2WN9DmGB9fw1d90bNKd3NBHnUO7iVYaGxISQJ9w+WIJCZkiIX1TPfoWIU
VBvZkc0AjTmeQ+7yj1dDI5TRW4tUDf9F7+XJPQfxhVydlCsx08r73KLXjxKx7+NyeqsO6IoSM1kz
q20MNAmbs7bx/b7u50OHVYKTRgbEUzHFxcATsiIc/unuF3tTlfNyXEWPkG/vSAELevGq9PJmnryy
LdmuAr37JCzNZwzkWTpo/caOgXIVyKd4cNDNyzDNxlkQPHwQHX5fOxBFv/2tAw9kMbTUS39zVsv4
BZCL0dz1fvhJOnijI0/gMtU+Jsk5uzgu0zo3YmkzOTGLVD5LMq5kF6Gxyjy0ZB5s/Gl9clP4uMyM
RRrBP5rUB9V4Hj4MYkivOlMkgph0D9Wjse7eFaUCqiuoGN7e+Vf8cChMZTQwiYPjTyS83FdStJDg
28DuNMP3IYVTjhN3xobzBMNAXelSdUO9rGcxrxHk0SxmlTlGPYZ7/IcsKMiinGrK2w96r2xZJqOO
c3X8j615FuruWpYQxs8qJC0yGPF4wBuGY+tgUINnx13gptpExV86GzIRzA5leE4v+YeFo/OZaxDr
V0R++V36FZjQtZu+PjjdT9Ikc1SKXvvCgYitrDvH92zliNridcXAhpZyHihYlBzxRrQxhkK52TvV
YTRNdUADDWB/dP1e2eVaSkCZvtROM01AZgnvVDcjcpsbP6+rkM1rzNzARrsLqMKeozAnwC3FLK05
OOUHW1u/AU1bl8kqjyx97qVmJ86CSofcAsWyd/lrEi9wkv+jLp6padrHp9z+TwPYjOSqzm+IFPzB
E0Xmc0FWH1Pi2GjP0Q48zNjz7NLtyytxqeI3mNHawn2dllze3uhp5m4/7VZw3fjgfE7LcX46moum
+4cTse5hPFCxj/ahjqGxrq4A5+fvQaJSHAoHPU0Ph2ie3TEF3zz9kq8SSCnuX8KkOt/634vlSs7d
2a1cf7sZ7zfOSXcMW9THw183l66XG2oxIyNF1BmMt02BqVVGz8/jhCKeU3+UNEIfiUl2L42rcRnK
FGCB5BYcGlpjB5iINdftjbo0Ffu7fohgy6xUL3jKqqZY2YHmGTqQo/11XzrbYWkUNGVrELEqYHWl
zcomY8NV9MxJ5a8BSDFRi9mjKe0q0YNLcVCFYQbfVWkfMgpG2iU2dVG6tHI9VLyjfJghQPI4mtbT
vnIKvUS1c2lVZVsPWw0ppptk0cq171mirtWEJZiLEt9OJYEvKp2PY0eyOJGPtWTuvINg+0y3Z3gB
O3B5569uuEILVMXIWIL3OLuvdsjvXXHG3w0jgFzy1YhTXHKbGYU9F+vGJ55ke8QycbwHL3qxQlSA
uKkYTbGg2x4Tf+0ilxZ2imxHU5nUAE/y1Np6wTQgrzQLgpPHciPAscLEiWPFJI/tQe/3tDOE2hK4
TxYyD3vEzjnaChHugmYTtYz6vCCUvLJ39MFcVRSbZ6hsKiB12gEo10ttgaSLJrkFZMFhgExHEeI7
XPO2jjiYN8aGCIsghxVE+2WuWv01xnV7aCdA7xggRVpNiPJUY+rLefg2VVUmIgxCVi3Y2ii/vDhU
PO8ysaPw6108jMWxsD5ITOq1nPpZ6up8t8cgREi3DamcwFmpyG5F/bucjhgUHxfByWBjEMnQoEsw
5jxigpjfX2JDmmcnyg0KZCaqazC+wAekp1/VmxS6q9+JaQQl7cg+Jlx+jSipODvGVZYNQDNC5jYn
YKEJ/F8oCXUVQkmeDiqQbc/W+zwm8Yb0eo6tIlKarJRc9R2SUqeTm8EdWqSitXea/onLpst56m0z
wXpkLNYsgE2z7Ls3iOgUF2MhGMcheWZZtjkzUWDRUms1WkdVvY3ZAtveomyfglkETewVnT0zL2LM
Ad9QxAXVSaWIY1fAJNDEMOctmxQz9QkVUM0CpAfCOpmWw/eY9v2xLdo1YUx0V6ePOfdYco3pf+UM
oSxLpx1cg8TLYqalArAby89ic4XvWORIh5OUuI5ZQSwlq0gwQU+Ebn4N/cB+Xe1hylt4pf/taR3w
ARg/NGc09zEYyd3/Nzg+kMQ53ozE+f8phFAXnGv2Hl1q0BpK4nN0xjVo3sTAuwj3bxfSXbcG2O6I
EbvBRgjXyj5lrrR412BKYREGXwn0lURoXVNv/kPTuXa1qWAfPGKfLQtzjQGhtvwqRZJ2u2F3xgMO
gIeK8miBI5fH44mqnSYERR8J0f5yrmK2ILYsOjzjUn1pyMIJ2BDY+5Lg8ZatwdqIrFMVa539Pa+w
oWHhRi6EY+tGheVhHEkjhJVks1yHKXu7Ym6WTYSVU0SlReYHmwTrvVFzNzezfkalrKBC3h5tpLxo
Zm2DDcH2qydoU8OEg0HaqmEatwfV1jCeXSAwD7MDwe5p/aRCPwJ4MOKz3xGZKTOQQ2moTbpJMrA4
cWdfYj2JC+ygBSqI2n+DwAFmx5WgFm/XR8E9oKMyWYCzgxhVusU8zP2IxzvCbfh3sD0xOT2+FWrh
UJLa+U3hC3HFXBSCeJ2LeE51dwCWM1OnrBZ+utHS9/5UO/M8s5O9e7LFFYerj39/gdI38ckT7egJ
EUHRWCNCCZUPfL5NwpvT1AtdoySBobjYq3vRzdNWhkxyUWPIQ+jJI92kA1Dfz5ghmYey4iUcTJ4k
WXj1oOnAFqDlG28lu/19lT/1MI2D3qeTMpH4xG8c7W7XW3+2dTBIZbq+ECyJv/0RhX8L4bcq7XtH
szXJz2FBdxnuI04hLfggtjECVNEFHAXR68sqCt1ipLHC+cMZZ7OwlmGrWEU1ExwdfTeQHXQrLk6W
xxPnMfaPbeZMDuQfW7HcFUiIqNpkSRprJgVHt2BI4ZvLjCaJ0U0Y8FhhpCDwp1xG38bl5H+0A8qK
am78fXm1zzDfQ5tDMnEQVpg8Iog+ZxxuzZxX/8PWjjvDDtJP09H/n2PUL0b0nPDJ9CmkzG4fJbr9
x83RAZ+KCJRH4Qg/BoAKdj+Y1bgs+kc5JK///ZLsKWN+82eX7ONuRKSjm5YJ2195OrQK6pYqhk8g
GHuu1Xjf3EIi8cNPBWx/hURpR7tKuy6vPtyRnnvPhWX6FTKZg7tI71A4REMDuzOEQ2gACxXNEjYs
Fjv91Ru2jbL8l+5m/EodXDanJ1uyZFYSbykSuWGTIxJq/v91b2UX3c2w8F4lz9Vfkfb5Na33JZPD
dU6cLV4s8cMzVkN7ciY7sqEZG//1Lq2cBHb7tbCfOH0C9QSidZ/MucbIMjTs3J4f//MvASOZoDdO
KeE0Lbfeh0zPWU7ZG0pckrLC+Ev7sqfTyAJTYxi2i4OJwd2kDV2TpwZg39LsJkEm5m359tCgpPSw
oXJNsxh1E89BIse1ZxggLknYH9yJ7WhJZ+SC51SzT8fK759RuEE7wBdPdmU4NQdqUspfHdPqEwBW
lR+VKC5WivVrbdqKW7ePcft7JobMSuvLbF3EQAWSsW3LWQkOan/L+dbCgaDMUI9ns04nd4XwGJ4D
NSOt0m8vpi/Y0PKdGWbbj3L+Zthgshdx8Ts7MKTN5CgWkkdCtWpBlD+o82YncgEyZeBLVUnpi53/
JhZKCPFEaLj1Fvp4WZcm7bLUIoB+lISLIAukOu/t4FWRWanBbIzZ/8nab3wOqdYeNMt4t5pYbLzg
7OtcMmPOQ5h136HntwyAggDbBJ4eYrIDM0hAoCljSfEr9VQ7HK/JDCY2wl5KozPUy0nPS3oOgosc
IPilYDXEniTXe0AqIQ0W+tUTSoGZHxwgzV4ThV+CYpddJpbcRNyhha1qP+8OEOUmwkZaVDJV0d2o
2Y55gNiHhrXrKjGHfd1l/k0DSKkOXLB26MDsjxiP6Ib2vFGHeWwKACEc/xfATgYBaIES6UQjFkyz
cZ1gZasl2z0C3dR7o/6g1vZrpxgtkYd3Zn5m/VJYskNj9DcOGWukeJPRS6VV7cIKSKzvIaA2T9mL
+8KnLEyn6wJrEEgjJ4WI3jeqq0iATRur3jDODpwmHo2ZpC8RBW5GOk4EujfX5sNkajf7Zjsmmn0Q
d/SFLGLPe3DoPYbTwOZKfxW0uDV8bbz5v80EPN4Od0f3NN+F+4R3LulnQqcQp/rNuHxCQ5YPZBJZ
FotPYMLxI/4vTE0em1MxzLlK/ikm7l4UcJyS+gRYdtsu08n/K3bn/tfxZ4yWsqoiHnhn74PzCr3w
exPmMJmzJ4CuoR44hvb8uTxLRU2Vqi9CWTObgAJ6urZJIQ9pcOcZE+4C81nYFK7gmsZZll5zBzPp
US0itcyqR5Uur1IPU/CDd+rc+4xXAX8VByiXsgjClUZoe0BAfv1+CPUjYKxrjdBA2noU2Ud8zlKO
+/k5pX4T8ckDXnMjWpSW1UZAh+8sAoGN7JMRzu4rZ3TBYv5JieIqKNRwqt/81eEc29iNwxvECv41
mFATGXcNvkuaxMSa2omT3ULko290mEUuRasJuk9PMkgS8SkLR4YlPf/PkvIyuULyA/TCgqwFy6YJ
bidAw0AQ+9p29jnJoTRVgUy+HlcX1mLcfU78QWX0BS0JMsGgWxiCv0pbOU7nCnGJOpOZa1DgfZh5
Xq0ts/nCngLTKPjiaTI0PIJJBhYfs8mTOKFJVQIS9sEcMntOftvBNKgProfmWx5TMp7niAt6QD7z
2ecml4X3X7iq+UqYRoOvxY7buWzHuauzg0jSWyiz2DadQuWY7fw2XpVV+LrH8vbqrIRB6jZCBK9Q
c1Ni0ZETQqmiVidGxV1l0wmUmGrBGt/bAmQppVh3oX2UK9IRETq5uenHKt821XyyrcQwsWzbA/Eu
ZW9BgI3RftOm4rukxG2bDCix/WQKifl2M79XMBUesMPhezgI7uwG/dhvuwu60yZSsPtOAbPete9r
r+DsB8lznyR2RR+OV4MCVX/ik/zavcCBYCkXVe/pihN3Bk7Nlh3IutN3EsKn0R1n42WoR6MmPjJW
Hiouh06lG8TD3bn0n0T+ddjKfsGixCWiixoBGXUrKxlUASHex0rrwlkzRQivnerSBey/We0XdB8u
s8ScEaQqQ3/WH+7LnoK9BeQkjcJmEbfK1tZhMJlgbZME8t/PNisxZgACqPQLGxlk3P/7E65Lhoxa
fl90X9tI18F+c3cCIyGvHWOxzDAr/ddsaV7pSe803PzyggFFjuZ8xb9FYjyOW3JVsyBapVWVT+PF
1ykv+w8Hdd9vER/Bs9ML5CC5GIm4bm2k3Gj1z+KIXPqje682zLhtafykrEnWdkiDVDUxewLnus/o
u9Z3OeNoe/8YyKOgL8ccxdwarBVq/HQggXGQerXVbxZJbTLaLv8Lq5hvEvA2tlPtwm8LGQhcwB0+
t8VCYwWNt/lQ1IHggAzxVjzKZcl4vXSUKKCR9449fKTIMWxYkeAM9z086hJabIl65ahyse/lF2rl
KPhjxDVygU4u6apiAS+1STE7oe46+bhCydeKMLcnBo2BtDctw8PAtnqSkehasJDNY7pPrmiw97pz
Q34uODXmlgVY3j/2kGbdxZJmkBvNDDTzpKl4MWGSZTIDofEEIDlOkJLNzSH2V7WQI4i2WeiHCkht
sHkg+qwM5QbXou3iwsBSAnXVSBdMBs6a1ZqYXV5YZYz147AU1XsJRqhT+v3c8zdBrd3eID4CvRji
A6JLsP6ptVyIfcOo4J0SB2INF3gUMLKstDOCOHnBpVNYwG/7bu1NlD8G6HJTGliInXumXr7ypr+r
i7107oZ4za/saUvK2vXIwIM1dPSTK6vqloha0iioYLPn4e8uV4UWOpYaDkEZIQzBhkPe0bni+NC5
HJiZzVk/FhAJGy0tSmx9VfKm50Iq92/3pFRfhn1PibOXecQT81iPVJvI+njeNzUSbqOJlZ1IzlSR
1y8SJI1QDW6Sqg/TiBB4YXl4A/hYTIPvyZ8PDYLHrPGW+PqOCwMZOmnJ2yQolbTKZRSDTj337M8o
BIKJ0JMhSE9dK0yA4hSrC5ISTpBNSXCwxhVIRQ4ic1m+HYrk+B8yAoDnWWW/+W+i6riFnsshOozn
Ezf/4KWvNNft4WsRSj63iyTuZvb9M+xqlN4HdY8Q/akNx/T/XyKV/jfYVm1Lq/iusAPJLCtZeyX3
T5tqTxXPXiM7hzcK5IngyD8B0YBT7GGhzJObX9ofdkkRdGFFd0L3Aq7BVDDOVIi/ZyqwpGjxLcls
pT/U/VgehelPgemroqMS4P9nLk5uq0pUAHmsyfeDBCXN6BkvoS3EqnKaILqIim8s0K9eBCoL8bVU
7s4m2K3tN7I7r1mHZcl7P4asnhgS599iMen4rsOGVC7MbiWvsbu8bPp60R7kkvQK1071Yw1n1Wa3
85sdYiYgeRb3eZlyvzOTyIwzMB8FmN6d/KwPnOcpkY5OTyCGNOTgQrXM5U9uSzziJkLAaDI5lJrf
mpyyELxxeXJU8nK/8Yk/rW5UwnNWsRd8jMcfoEzYqfv7Iizhb8DnFxld4KD5vJYo0dDIm0a/9shM
VYLhh1kUaDZ5Z9gwpOo8DqvPid6nLKXWSCmxh+34BszTJ2+sIGIERHimPfRkCzs6vUchYbwcktR2
FLZejvdd8LDQuq7IaOabOz9odlvo2+PSF35V/cSU3Whtq18sXNV99n1X/sGk4Fb2RPetDLAS+lvq
2jZA4aH8DczA5dLuA2MuCQ==
`protect end_protected
