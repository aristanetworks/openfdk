--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
DCs9phVty2cxdDwMiRYM/0GQvMglLbs45rb8e22yflpO+C0cMVxouudGhJyfknQfoPCpLnBi9C6a
nw8/yg3M63JdplwyPsWZpYJAyd4OGDCqSsNrHZQNPpZVUrcP+J8X7EYOpF5qZ+jV59tBApvbhC5r
wEpSCuAAtR68KQvyB0OVNydPmu6MPw7dsSrch2RXOw2V7smRC/G+aw5QBZqINCMEs0oHNn7i6RZR
5R08CBWkTHxww7FhfDDwBjLIgk8SaQ/bB6+75XPqqrJxBotDSugl00dP2tg9MGTdsUBY6fkicDvh
Whdgu3eD9h8tb/RozKOZ+ZwOKbRr01g8pOpUhg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="iGz2G4PbIXq0G02YXdXG+KJwLKe536MeigfBjRIUwZQ="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
SXCvhJ1D2ov89tsqnEm3q6oo3FnLq18gSQkleDbiFiPG9BB6aZSD66kFa23dxlJCNVT5bMi9uIkB
iSHXXSIc3hI7pfopA4wzNeQ+eHemwXvOq/mL7a1YWfH56RgS48Y3pWcqNIRI8FfyiuKvyLFiz9Nn
MHmoa1e+QSx3wH8YOLCAESHOdzAkRnt6UoT1CrfMm4NiPn4QvyxmBH83iFZALbQIVUFFKEp4Mm4G
QjQujcTS8UtiBYxe+hQoTZpxh8TIEjssMCZ+IZDibMusGIOmHgvMlrJac28swvLS5pgbBTORX/pq
MQUvbYzvgkNhsNlUziv2HmY/70gSPb89rw+fEw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="vR8wdD5ppCTssrXbjYXQX0MDaLGl2+Nm3tUn5SxYU9o="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5040)
`protect data_block
0e6aVUcbYXlbTQyLm9bb30RZWpT5aOrJUDJErdNKKVZbayFUIIy0yUoVydJAv2UgIYfRzruFVzPH
TGBO++DUXmpnHr6ImDl3qPPJhMPN+utcZGfpfoYTp4K0ibYZJSBeBaSwFUTnHNbT1Vve5tLDqmFg
7fyjqapemx1Chu/AQJOwxhKImQtoqGeJ80t7NTQbWnJX8MlsPuGTfrzZ8/exqov759TtDFa7DF0n
eCxsWKv3VTfLDt/sM6GOXYrqrimihhV6ByPywNb/L9uaHkf4VYptM3/JGuJeYhQtxacMa+SMh8dj
pOxt5fhmg/sCgO5SilNwFy48Jy7SN/VN8L8o8I8UZz3JB0vDTACPsGYP7kUgZTHxmJd7QbHqSObE
uRXiAOmq0gKKya+7wdqJ7SyHUbLa72A9x7adU6zOwaaTRTWfX6IjLvwDIJPyqBMYyBBpnsoPlD8U
VzjBD+IzVXNHml7uUdF5qoZk7qZQ52j5YcGbjt9PB5GczUQCsIDy1hQiT1SiUrw/hmBQshRaoOxK
4+eLlPKKi0ixIC/5pDs/lYdf0RN/Yh9+6c3Mq+rTMIRFs+wJaicdJYChmHblNswjVnfPtAJBXeTt
BNP2dfoQ5hgcYls7eaisk1et0DrLyiwQmyV1WijkQmOcFfe/yoVF1i5Q7NvW8X7NF2pqCrURO+LR
W+kfQZ3HWsVPchNBG3/Zhyb2zD2QlJfH5tCQSXecqv3jMjPd7RF+ZgOoGj9NYc9kdAI3SiOobLR2
5fvgrX+wcaXUuU9Yj4V4Vfvk29ZRaWhwwEwhAPPmTe/+nfcd8D1viCEGFXUGtEcdfgg6qfs3UEWz
3cB2X+epgguKohjQfXYx0XRnYreJ4YNFoWw7y/56LDN6VtJUIqBtCHli+1UuvBIpbrkvdiLh7vfE
7rNEJNQ0L3oW8orsQr35hFSvopOeyLkIbdnEoq49nXOKH04F8r7iiKGNdmQN/51G4tS1mp/xsP57
cw8iJqr1TIbz1HO677FKSUysYEs+oUlMzSHuLRGF1b6Rb4Nvp1W8+mF/q39HP+c5uijCP/uPb2RN
t7goSo1nUYiC1Wu275GJMQHc8OZpHmyEYKy8xfsU/T9fl4II/GLflturgChtEtgX/PJWKhGo80qy
hxoph/mfRVfOzq93Sr4KNq59i6kuJirbSd/U8EhFMBRektyBTxZ1HSFAHh8tIFsHNMqVQfmlsJOF
fr15itcDDNLamPr3ZLJcPMXkIAJ2wuRMD6kOZCX7+F9OOMJMt55r9DPBZItaNi+7obTtCOOkX2p9
yOkVAWHodYPRVFhZ9jCuZ6HrMER0NEzGVAsgiP/BYlN0+fIhF7rHHjhjOezeuORhL65MZUX8840Z
eoi4Rxb7rtSqnFkQsv6IgUNQfYmmCo+ZDkpFNosCAoqfwSKdxsMHut8rY1H4QvNDFIAa2i0hVyFP
tvtI/OqkvqY5lDsyMjjRKiCWToTlv3ETcuBxIc5Yuq4tbibH22gFZ+mjmr35q2qjLLfrHBcirn2o
aNescd7h10IModhkiCJ/GwLWFhTAB8JcT5l8eCqINLz7q3vBRMVZZD3qm60pcPSYhd0hHy5Ksn49
lFabtdW5V0NNGKR4Ny187CTitc29aMKWze9AaJqSAHMfjAxnMtyyI7CH/e1lWqaSv0lbdtVkkRWv
035uLbn08AsGMeZhNkjm8pHok6uZp9t2c6Mg+Rzbp6Qq8Q2U85KwL/RCChthGIFpFq4Qk2t6lUkA
EENljFTkSqNAXxjTPHbWYcfjsWyWm5z3+YPEYJ5eIBAA26nPSqo6/t2TzysXhbpcdYmlIavAEmdT
KEqL5j/ECjz4RUvt43oKv1+xiJWZUIq+DPUwFAPp94nK8c5IsogBNJL/FRbXZ4Yy2DxUaVViU0NA
bljT3p4NjTI/FIUO3ekEXNBI94UJOAot7TOCbuJByTUkKcQxU6K+c4rWzvPrmCAXdd4pgpd4OLwv
81sQfwALwnDRYEkGRVh5YJQdEPxkPS/iI4gFlibcoH5WhCSfFfWzfbIEY42ZrWOfW5UT2enCg8K3
gIMi4mzPKaK0m031P+Lmq49HDIqeSTGzahhxawchkpUscjh23Szv1uIlSp0gE7bHvzWSkSYmBNmU
+SOYnjrbsdjlpeh0EROE7Erd3wTJBwiDhqJ+5DjfwsA6YKxqZNre9kXR/JJ4l17NXCDJiretJT/n
6o85nsra3hW3BR3sNtE5mUlLtm+dpL5PFQ9XIh27Rs8biYNDzmacPyG80HK01cRiFcFXR/paczAI
DGZft6yIyvuqgwASdMuEYvI0gINCx/YbKICwHgvRK8WGEZBvpRmyzCaSlmVVcv6V5tRXa9fyDDoY
aaWUZJQlJCrBr9pFSjzDmVhZqdZiZ1vV/7v0S/gxxLQLSAGnSI55KiUw0elBt4vOkNXebycbSYbv
/2cvWj2t6ZQRMLlea3CFS6JViB0MSCxJSX19iJ+ncDqVrnd5joWQiYER3i5htDfvbyshH9eb7Bv+
DSQsqT1g6DdcVOdkR5I1FEWOBSrsJVmedgrcioVFAG6SfMwmGlAO717RRIUEYMiFaAPGDnLvT1/x
qb9AsCltVYyZ1qJwyjRiMgWULmLJP2o6OGcCQth4l58uAbQWZauU5dhxs65AwOOLvAW8p929C0xk
lCtm0r3RFkDaV6RUVEQvFuE5A70CbPDKo/4DVeTkKEsdJFSAa/440Pzt+FqQDrXvYsbnooWWZ/gr
XmzaLIA/yyIb8RmDuSGVX4dIiX+ixW271mUpPpVLAe1LPHXX/2TegbCAj6euQAUwNQDD5smTdak6
TN3gA6vNSy93SPYfvtk9J+LBs8kHsvYqwEs3HTbIVXzhm0AQBjCEBRWbqRx+vm8m7Db1DkZ5QWbk
zzkW7rH1lmsctGOaOCuzgcn93F5l0UCDcOZRTSaebfXofgg0e8SN2/6n1PnOYdRrq7aGatOzIuAS
M1bB+YexxU1v6mfbvdcYYGRLWEJXzrsQ3KUUOXnvqcCXrfpCdvHc32CxqZcWBKaWuw/STCQMgOHy
yYBCDLLaDoiUDv9gNxDc7n64qLIvokhPwSFsCF3dc+jZ09vw/x2pwJX547PcmBLSgSJKuvCP0fO0
prQozGpprm7Db+2tQGog1eis2xuRJvaEMWneMB2rzEXlDMKRV6Y+njLLburHaPzr29feElm6WEW2
ZQhMGswWM1nA8Emky6ZQ/8hEPVXEM8cCiDOnJc4kfjFLR2f9TD/ojdSbrmgHMwg4w7iAumvx04/1
eB7XJKXXtO+mJBZHDEwtqQ0L863jw+2n6QdZw/0MSLTPBVThmYx9GEshfQSVKBPt7Rv+URUr03d7
7k0OYmnAi7Tg/WJaNbGsR0zaJ0lLQ5y+P8Jjzx/QUcplxDHJZb3aIIOLeNpk4ZSqhQaHL/K3ovI0
sftA7QS8HfnRxjSAfyAJWGA1ha6stDxplbTNPEeM2IU1jqlFGugr60/EyOr+Dq5PqyCD34c9guvI
KwmdrFrSFsRJ+6JuLm8U8IQjJEpOXumQx04hcJ36nPdzbt/1c4nuW0NbIKq0Z9bnrRfgfZsZ8XZ7
GMLBtWRAjRx+ELDtmzqLBpo0KxaIyDjApMXv415XjRqNDl/1YnApztFBXiiJVvYRib1y0NIT3vCb
PUZ3bWyka3U+zmym3wcQcV0vjGReN+jUo7NB+LSRlQbUbp4S41/az9pIsGazIEs91CunzuNpN1Sy
81l0Row+g0uCpqhoRo+TC9MwXDeab5cPr/mkgpxMsAV58DQG4o6hhbHbq5JHFrQOwwtOAwqjSEG7
TRb9DxSljYj/uFMMKyB6sBvtRlwT5I5CC0ywL9eiJ/jTI4ZdZogbet46GpkS60+7dAswCQLXwhld
Xolnn1PjwhyUE6cdR3+Mmf1koXLvDhqmixFyMAHnYomfFDIm3zSELeniCBCo9N1LFR/4OkhEmNSA
9dtdoiHqy/mWJp5XZ8wxLzUkPv+5jWNQbG4xDpTnLkeUlCMiu0LbzyZJXgZOMgpW5ID64iZ5jjJN
SXp16SGKDlcrYJCO6Ohczm3h0R3OdlhUt/VKXX1fJLZHdejEF/CscR1PFWh1215MkCLsFp70bymc
ucry5PdSDlvDJ9NkyPEYloJUT8lO0/15idvvJgzD8HLs8zk+q2R0F/fpX2juxik4tQV2QIm63lYf
VRfSmbLTUZU6bIfPVAjUoMUUtu/TqP6YdctvCKt5KJ/UWKPAL1Ddtd0aIRudtgHfD25a72jp+qpu
ep2+9+plPTz3xs1iSGWeyBA9wdXq3StsPzCvg49ICG/8Wn49ov1EOpdGQD3jWgVmYOS0S0QCwi4l
DCNL3uDF9whvIn1+VnR8vMvCkAzuE74QynKktx224m4ljXKPWXtzJuzotKxrU8VFr0Pxxfeb2Vnj
Xn9Qvtr4xtnWTMqBho1X5PuokO/Lk4GqsMpteQYDX3LSVXAbXbleH/s5J+E4D07Lasur02PZju1b
WtHHoj2/gwn9DW0VxLJcHLRrhJLBcsULsp/V91Hq8fjswRYYA4WeXoP7oo23pZ9ljS0Owf1y1pKt
1m/IECDeRyK/oRhjMfBeoJv1lQloWf+SNh0iKvMkZL6NLZ/sptRvb2mtD8U5DZ56uu1D+qZfchw1
zxsGxBI1FkdrBqx3+05XZuIRtZf7X3ekRW9927KZwtt8uvzuDlNXxtcF3598OgJ4yNIfzlVLdIkO
gY04ssIB7TeGUAm5hefGeBNJHA9NZpwJz3mKINuFJAHEWbU6LlanS5+756rwIh27XWZJDGNEU2d6
4fMr28wEbJBRhuvX3CfQB8guw57Yo5OUzBkR+TqkQa+nyOXZSzh3UTly8YN8UA8/TqbehqHKpgkW
7lTVD1SSvnZkYzZT+VD8wNBRsOzyKRBtIusEYt4toayl6yeEZ8QWFnvdj5jo5BYkrbUFop/axLDZ
Kdum/sMbgUobKHVBd4YShEoaDa1d/HFFpMtVYcFwjj6su+p/honfWFVdp0nzwhbYx9H3sLtyDbsG
z7QnO4tmy32+TUnYRMMaRYu6KdJAm9vZCJEMTv/CkamdJtiLax2yinxM3lBYNCF347jSoqlzZE8P
EH2z12c0M1sGUWajNIMLXEEaGxMA4KjZAHyUel0gLkLKtxrn65fZhmB1tkq5XAMyARa0Vn1GCwW7
+u93cihtJ+TqJWTngzO8CCfnPpePHOigGzyn0ch73NrXN4EeTo6If0xP11yMk18q0OTnj2CNlDyE
Z50lds20iclkJgrPBg1CdXLH8cFBvxbqmJgiPm6g2J48hAxcydbem4Tl9M3yLPn0reMCvA6ph3Ap
d1pdYEqGe6jBR9bYyxQt1PNtg9abZ/IIfmtzCIhD53o+k7fDm5jYiBoEJpwvr3AS39ijKC7j9qqq
uyic1LI5uze8gRKc6SDlqvFHSRhLHDI31INwffsMX4SuvnHodvqOj81jnZ0rnVfl/tBpuu9eqRTS
ABDvjGpp+wYaSbcgBlW0pm9t0NOQg4f2P2II6bDnjQmqDcHx/aPIAmB0/We2HaLldH9f9NmfEmqB
77jVAJDi3LqMKCGmbBrFQj2vznMsGqVhpWMvHRAkPPQfBKTiehUCsHbmfnPtGsiOKQYhYV6trnZ2
7OQj0bCu6Tz4FJqhS0jcUdsdMUgshrsG0W+4Yt9lgEDqFVnkMAm1BcK3DgBKMec5GJ6ZhTSBDOt/
D/FhS/EbD4Ku3OKlRcx/rz3X08tyA0g8oXdJeu3BG8oIb0Nqc+lSuwCw8d78aqKHY4vp/0b76tNQ
RHBU1blLpTyLA3JdR3H8Tby4z4rb18yiSo3UjHWWdfJQuD3KfpOM/URR/rO61HfWEoUoBQ3Y2Uf1
+xe/2S78YE/1CX+wdlKAopYcpSZPE0cUfWseT8/hXDG8Ujjh6kk3/IOY/durTG5sgrtHP3YLOKQW
R/fa3B12u36ou9ArxXksCbFsjPjHymZkdk0X/eGsNQx7gHcEJ6y6rjh47+jaLBu8MlSGhcDmUQe0
X1HE9WISteiQTH59SKt2nrpxis1xx82Dry4NJQpySf4r1P8+sYqlTKVG1G1NxuZ9GzlPBrHRUBqW
VTG8nkEfyx9k9hzSopq4YEdqZ4FnmK6nRyF8aUxXV4WJ7Sa1Hs8CYcf9+tm2W/5UH/WXPf8pdaI+
c0rpSqbX8MKCFlrISddKUAUvJjFD+VdQ3db0P18/U2GVS+nbqpb70X86Nxii7gsNEVf+c50m+ltL
McZyQm//p/lhW8xs1a1GosvgYOaruJLPSRQepOA2JJO7UGu1ClNbH34Pf8W/yqy65mipE4ysTiTs
N+kgiIiPqzvomFXHL7iLneYqJPIHOjx3cmqgj+8vJewbDkccoK7VNTfRELRxmA9Ot8KxPCF8faba
aLx4k35BqXfDcgaZI28HvNpMHqDBIC4LW6GJ1LCMqWMiHB/X5qaZPPhR97KWyEP0KUFjw85CIv3L
wWmlOuTaqGCN3Qqtn53IHTWTodjPU2XNFeloTnOWFvQ95713aODkW3VSTLmuPHoyMSNvUQ5fSReO
BREmfzxpkLg3Ql/ajyY/PCSnbbRm54rAv2/x7wPf1ROcpBjKLJCnUOZEbKbsrUy4qS90M6qNBBAy
qnEJUnnEMrlm1OfwTY6dVhZayXtKoFp0fIAR/wUXDnNwcZVxFL/zr+GW66biIuCZqXvGe61WDJI5
1ycgWFy/7kkcsmmqpO3mVBoWGckb6afg
`protect end_protected
