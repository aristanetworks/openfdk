--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
LRty1FR646uLEWNZlqI4rPEpX0lsQN+/b152bmBZEAlTGzcaGOF1jWdGUeQvHUloDXHOm9xTDpQK
XQgLsO0fj1VeifF+ROFZplfxNeYQQdOd/tgMJfLmpQ6B1eXBYJ4meCPgbqKmMnx7MuV9ZYxultLk
mpkh8rf1j2Rs9KZbgKoaq1l2ryqEjNhTxLcfv8tQ8gJaDQ9o+8xw54NJjV8q8FuBxpB0Nh2pQbny
s8FQmkmhDHiJx+wJ1ZMQGhDsPmO7i9ASH/5ek5fwGYaAngP5k+XCyND4VlGO3iO8SBg1E5JG5dfe
qwuKeEYA/HsN8hNUqVu5qpg1jRgF1rTCdpS3qw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="kl0KGz59bGT1mQVKtWY9wq4z4LdDMgjXfGFXzrkRFig="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
ig8Op2lDYhzjVcOnAecFm+PTxUosDmKuNLQ9OtA0NrCbjxboDVavt7PZBQWMxpv33aYoygsqErt7
ZgZt5wIrRL5tPW5KdUEzw2zjOANbuoIGX+6+4PpWflKuorJ61Hjig3Jpvb+QRPmrH8dGrw7L8WrE
iSzfLI687lXtDuAsotwmSPT3wiozHI56itvZ0jWIZZ6By/5p1+0l71zSajmz7Ujxhc8mq+3C48F7
0P0kcke1yu/rN3I30KYYHyO/Sv5TV/j6ERAGnuYk+6GZ0TlrWX2aj2KxVhUKIJ8J2AbFQy6QbH8r
aWvZPdpC3iVt33oqBHWWYsGuvTOg/vOivRuQ7g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="bQekKJAVD72YJVEoX93uUgDz8LPmhpIS48XVDy2VSKQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17888)
`protect data_block
hEb3YqDsq128jUuzPdgxbJk0Eyruk2Ag0qm0zV9GETymThYDVAuAEZsBjcQOFf9i2WZCQZSn+58g
kLz48rjYRgcPK9sFROwKPvOES31E/O1RfDA5FIhLskMy2lwOfelC0/fKYuKJIwzmTIPXpxcAwq0m
01OXXaclhS4G95NVD5QjkcJldlUW2ZTnXiKByYS/JZyQ+qnMa7BBey8wAtm/77C8DuRC0TRriIso
//nY1Bt4ZZ/M5ZfYPhDgTrVfDBkZXBqCilkOIQteIGxlW0xgUw2+Si3XGanIsAG9nElGeOWa5Ni7
y+sreQBiznzB9UDuSEW5qZCH7UB05w2On7HzsIofFORSDZl4K3dsA1Aflk3BLhtE8LfzgcaMJDoF
Jye5Q4y9Vhn9j5HShhzoYuLguwm9GKhgOuODK8bvJzEU3Tc6071lBRrsc3k4ezbCOwdsYgjzCM5D
/I2Pu8A5UBYrz+CFEI8mxav7/SsVCGJ63NhTAFlm1peDB2isqZDhNe96T5LQ4ROv/RoIqv47emjJ
LFfRlxY2qrUQrpraReKnzcfjEVlT8reWHLJUqez2A8/NDn2OeC1w9bmAnkp5Md5QZv3MVrUJZbdP
nmPHIWiUJPLDUpo7kJtjRVGl2yy382lwj8Js377EpTMgs1P3h8wO1R8KYmuOmIY5mcMl14Q05AwF
ZeF+4+/PeZw+gs1KeAiR+zbIiEUZhoubyFUkDAQGOIBukztTfX+ijQffInnn2lV/9M8GedRM/0LU
DZg4a4sXHPl5sGeG/2LEJpZUG2HWocZsg2316TQOIxvM6rjKtkH+zcNhQFCP4/8Frq3Aw+x/xTXj
msQJeYbpbI8puZgldRtCqrk4JwhiHd9D/CmqHz5xEGPb6WkA2GkHWcz5gYs1AzzpC7y1w0zJd+L6
kBpNVvQvnphl2uz27ba6EbjYpy1KrnuE+krE780nV6FKVgeeakXul46QQh4tnN7o9L0iGPDaDNl5
BvLid5mzXuqpQPpmSVZAAmSIGE0uiuRCphuC12WtinkFyUpYWLD683k1jM+oGeHfRHscMSKXkE67
oTuP4z91M54sPXYdLQt+EF+O9JaqMqn3ZASsc4PltIjRMEDER3IyQKbGISZlnze93YqEiNNiwBap
Ur2geOKS5FUY/su75P5k+ii37gIKUJ1cky5VxwXLjzQiNJo6U4+MQE/x94hb4Pkqr7ELqDyt4CPo
j7c+vxiEKaJYHNWZHw6Hsa/J07kNnky4yqqx9YMGfePh2wTlfThi20IQxT7cSBrcu4iLI5dY10mt
04FdvLGlTbu+pA5OiMwgS8HIx9Q9kWC2B0MOx0YlItTodYcG4VZEyMzVp44/n0yH/JMcrGVAygRj
501mlpePwl1/iqs6UQohotAGqX47RKZOhmLhfvabs4eDTITaC+4DTL7+hyG9vK2Iig7s9RgWELGH
Him7GvpT6qx9c1MeBG/1zi5JEeCP4zGgjfJbaQO/J25OqU2WdwGooUCkNyETl2HHdyN9oYh6Fid5
COu2BEl23rmjUBfLE9ZQ6yh/1xjZFhSek1CQQHyI6+hkgel6o5UuzAtSFGGIeKqm8CfIvqeoXlKq
pWFVeV7Kg9Dd0i8mtn6PFrTEitD9QsA3FHVd6vwkcGqcIWWEakhjZYQMALX/2att5snUjaqZa5nG
jQA12MY3IWGSYPXHR1coWWPghY0cQSJqxwpFVAXOozcUpm0iiljkpUl0kTjQ7EKiyyFiwIi4hTuO
U8ty6oaoMtzvsKObNsbEpkbUevCXltlbWG+hQbzcKy8wDfNshKjgU59wm/jF9EeZa+5Lf7cbXXFO
jFJUkiFG0EUej+1Se8EhUkgZBBBmM04iZsU1KF0nptMsE8P5mSnM6cAnkcK3vhwVIX4ESdPuId7g
dvXQFG8f+Pbdbdhu1CRL0fz7RpiTWMpp8kHrrK8G6XUaee8JfhwBqeuXweR4aR8Ch2jZJQ5dLS2g
1Cf6bGszguS5VsGmiyUsdUq47qo3YnlJdalsmdOmqZiNR0uaXcig9yWsRABFTM/LqUKMwUctR8oD
xbuGMnQi3qt1V30DMxKd6nolXOvbCHOY2IDhCyZAFWVkb1TCTQPVi39/GAMyU4vqFCB8SyGhb4IM
P7lODhSe6G4sgCtrRtiTELRrWT1zUWGSxtncsXc2iC59ao4uAp9ZBiBKuA7qohSs2jDKQ9WE69jV
uZCm32sNu32NeBqoaj/daV3QEuS8ZcioXlbcDlTiCfQBkX6g3MuoUKe9yNHCrC5nVAvBdP/q2ZzU
Awi6FTvSXElXPdVVZ238MGpqLWt0O+7bH5XNct3zneqT2Zv6fArp9eV94faXDU+XpKse5gKO6Xyl
FKhD03akHJIOY52F7y3xMhNS95YFfRKcztiEQlorKtQ4+MDeic5harB7pT3nDiroiFZPOej0LQ1k
I4oQtV1QRdDGTzZSLL2HBykMSrMgNA7hIltEQj9UGFQvLVFT3MEZXo84+qhA2xha2SI5noONn4c0
gmTzlB/fGNekzyUUXp/QR4jWrIgRjjMdRZm9sQjz4jVyt2Rf7vLL/bfR8odTioQjtX0SdDGLc18J
7lpFOnhuO4xafkhsOFScXmOs9e5xoS2liVOMIhfShiZqymmYYP4WWkign/TtMnF1bnH/yJH7b5e4
4uCbfEIeS5FB+oodoLW6d/lQGk3unEgu2i+Xaeijd5dkCz0Tzi3asAAycw05R6Lrync8LV712HZL
2zFz1+9PG8reKWMP9vBLZESOHV8oIFTdHccS3TqJRKeuDEUVESsJQg7rzlblGPErk0YixaoNjaG2
Z2PVATVU8VNxYWzw73r2siJ2E6Ev4ModoFGz6eEECHcWEd9dt6RCBEj8MFEsdXISo8Ir/U1es9lx
BGK2Us/Xi/OQJeY1BM+DvpxpYP0cD59ixj7+oPEuVGONb+Ro8n8IPt9Eo867K9oOJiaP7joJ+9Ie
fs9kWY4zzDZ8MMMYmyQTykqHd+ogpOLmFXWOBD5CJ51zNHMsArXWpkeCOgPCsLg9BV+OjkUZXNc0
bzZI1DTjTtqSVWUqBithLKfEes0TI4U6UM01ifS7CGGag8xmP3TTZ5w5Uy9M7JjmF9cHHF9pgs+Z
RNeplTTFPMG3J1qXL5dYNxo7FMYsmM05vwys7DoLgejqjikx0KohhbBV0aHScSEYsFkTGrhDjjAO
yCvg6IH0oGidi+wO50Z1TXuJNR2Zx/akMK361Tk3EAb5O2kBdFzmYhNvGcEA5JMAboA4iMxy+zHz
ohsGCTFF1FPqErkbLIUtcMEbmUajvSEVBliNj/oKc/uggx8aVydjRQJaqBvHIj6o8kA7AshKK4j/
IsnrJgox2ekEkoLMB+FaNpHN1P5Z3C8sfxtDNiekELaNezNFhdwuHTwdl4IOJERFPFo66X+DRI05
kdNvT1UuDMk0T+Kcuk6jrcccj3AjRbAwCOwTT2nBYFu1QoaMgpWFMNz2HOkqA2BA+mE1yj3e6KcD
3qtWlOQzi3jh/Dy7pF5UoxUMPGBs7JE7G0OTnfvaRC9JNC8pTavYcjAIQ6sJ1cj30T57WprCWtwr
qJq+AEFM6SvW6UfktGH3EOV1LTb0ewM0HMKcrpAVYzK4QlB+b7lAxsdTpNycpLa/Z2YruzUoFAwx
lQbl5J+PXQhy5SjnrIac5u8/IRCVcAfL+3ydoZyTjoJiDrCAIjPfzqqoJBSlQ5PikmFHBfJaKZP/
A08K+HzDHdoshp0ZuGcdIYamjhQesiCovvrKVVHs4B1xZ4RwQV7AQQIRlB0Pb61UBSBKj6JAD/CO
BQPRfvckHwtH8V/bDngXwlBozk+xhyU78ShbFbneTAB5JAdSS4sV3sD003Zcn6fBl0WiuxxO7R1x
67Vbrdxe3eiPdXBctikOSFttd/YNmgB6/1nOEbhDRd/ZnyyhdLsniGHs2AY+kFi/BklZpQLz3s89
0f4hShulM5PjVKnivaE0ZsvaneUSQECHvgCQiPQ+RhhobfjjZHw0MHHlSYetD3eGlC6pEa987gBl
IB96CLu5WZHVMmIq6wib0AWtyxY12dQsSI+ouQSCsP+ms7zAdRBWFq7foDvEZLDN6xDBkqMCibf5
QzMQIMcCgSi1r0eSOyMVdWyv218SMCWJ9WH3YaD3hWoqCW74l0Y+RzfOww0hOK4SE82aOrd1pO8d
FkjdZ8KUfxPVGG5787hbEYnxXLBSRivXbjOo7eqdJljzxXVG32g2MtOmiDFZxbeOpQ2iUggL2dON
fW4VUaky0wkzomvjJP+n5AShUrGphjoWT56yNl93O5G3TqqNUi1qGLIYRxSDq4hwnYXkVehsChsH
Kqj4a7rYWjQZ3efMQKShLxNOxFIF5Z39dSyqG2L1pmRmjPidNlvdjl20eRJGTy7Rwbi5beR4qT7X
XdKkbakbJ+wK/K8P/d8ZfvKTVnrC9PPBOzgqnJzGM1Jn01RlSLZKiO9qE/1nTnpjcqHGpxNQhvM+
1K87JLWImQWleElR1RwV3Vg6mj1M6z3FBid+jf/jyghniVg/MaEZWkkglkLVgw7Qafha9jZ895B4
i+IhM8fFzncPWloXCs61leyIWUqdBjcoytOujEwqXt4NH1wsnP7jGjXeurVssue05zdl4GQn9Mjv
vH65EGDSmyCBAotLHDU+RBpwO2vDSL3pXJBm9t1i964/laa2dTVHWEjOpQyvNnUHtp+N+elx1/jg
goJIwD4FZt0OHDPRJtmJVqWAG/93GvyAtGKvkTJO+EWMMdrTP2PB2aHyufT4dNj+Nvq4af0pqpV0
Hf4tezcBnuHj3gv/1Ui+aQHi+6JGBJfuXj2xUQ1MCg7EeiGavQky6L13o97fsIfm59sGLOWouerR
xrXenHH7A7oeF+/QPxHe81x4jNBBCPi7/JfhDXo0XqlM+qvlg9C0j99sXKSnOHsVXHUmOnMxoylK
9efSDMyiRGGQBolBbZuCPbY0UkPHYYGgzziq0HnOANP9wiHZ7TRn9dmebipfG0te0L5xYUCaJVnr
uyW75KM+JrIqQgzh4rRSwFLbd187qLwm035pHJYrJteuqMcRYczJRRORa34veamrgh/prGmM2DbV
p+Mll7Xw49X85XArFNtzPlHxvo78TDFT+mwWQ18tA88GGSjjDBxu01grWY88RjSQCi79B4UjpUOA
qvKME8gufkY8bAnuscI1OW6ycZPrSMY5MpfwbK0Zk6id2j6ZY+ueL0l2bq1FVDian9Z2n/mPrntC
VSyfC/F+q8skQH7gcTMyoKtANZPDnmOSsx+9d99ZpiAk8TdlBD9OsWwc3iAiugunB5/1abJwNvBx
awAhprJ99Z5TzFu36tpDxkfTaJragJE+6GAEDFNoD63UhJ203juAwfZKBPZ9ie4Q2TFxBwoVRJbN
CNFGkH2MCG1tXxiUth6/oAP1btx/J7hqsXO3LbJOZQkZFqxDUK9+ww0i0KOfag0vgJ7c8CyMd4zV
ReT/qhgiWyVL/NhZSiIBFfz8RIOpUBxivf9WTdaLZyl4Wkjp4seS+eypYkkEzGbdqN42XhuY4Dq1
Y/3XUMshq9GCJ1R4mkmxn/AR7V7gwtVjSaRdHBg2nz9Tcnb/5ZTTs/IOAkEjBuaMd58yFDlJDY+E
BWLv30vkBLJcmwTWsgfeUIWk+LWWZgoIgcME7kGE72FAYBqLfkh2ikYGdq0Kuv9gBksVpdYfBHed
Qeh2cxgNRmacsioBhh8OIhaowVRb87GP7jC2fKf8F7KKRN3ZAaJWSAt8WReTBsjob9fMox7C2Yb5
TvZdew1/A+mKzYliFTphMIdCSuu6n7UeZNmV/7UaYkyY8a9WFPROtHREcaribcZ2/srO7J4sI4q9
HjABXpneSurEP+ROzEUxdASiE4vsBT/CWkhccBCY+g6lD5sRcTTInDL35HMV0ymedq2Uzu9Lnmq7
GL9f8kANkJ0vAu1NrJZXspDzZ2x4GPBJv+1NHXx+g/vY1dTt9UqDT7HV7o2klxzvUdqzXOUdHUke
V8nz39yi2Rz4OI7IsHlziwPhBIZlI1YVp+2aKYNYq2xi69Rs5BdxAl+lQji25mDZl4h2dTb/aG7A
UCuh3zNmSIU8pyWybqPmuQDdRjw+o2IjpZHj4qMlrBsAWk+A1wzzy9HXhycRMON+KhvtCa6XBk/w
CcqtJSY+vu2F560iRVU7zHS8HHr1Q8efTZ+9o/vFo2MvhwGhmiFZBNJd57x2fTTed1mhZmFJgSnv
OtVrg3/WYQPS47PDyY3r8/cgFA6ie70sIXfbVSnbHp5ccWHMdbHc1l4jzml/5OxNkXgDZdQzwV3c
YVH6R6zhXpEpqgYbtFL/thP/wqZjMBcW5JIf3hE+fFKShdt38QJSLCoI4FQXnaIV7qlJK91HyHfr
HYA1/JSkIHlsKlZ+2J1LrlUqC4aBQc9iE9r5BC83qcRwTb0hI6eDYbv5JZzcVN/lgRfxlrV+3kDh
00gdM/kALuRDpWqiWndxZRtCBQXP6GrUG+ul/n3cou9IEYXQeX6hRSRuJTKzuih26CAN2KVIJUR5
nwIUXsY26dbSB/pMujg8PBfPA3jXjUBkh6kBFnDkozi71+OMR/b40vkGUfIv+FdU645nEguLLxjt
gUgarA+PuruVKpe6DdrxJdNv8wKx7sYeaCGH0v1vl8taS1UHH3ehcc+GzgyS5kX2PoAYR7MHnfuO
rMmKrbdcyFgUcpgrVlL0zC/2UaSV8caTueyr0UbNM/i47wcvyBSt7/VdZwlw3VZ8UQujU6yJYbtH
RgWRMFmMeL/2M1u0OFnNNA8QVZ4S4n6DzS6JsFJJx89P4CZl+kRpGREX6V4f+sGDJ2CvkFY9nyNV
is1b9JmTkvDxRTNltjv155lvtcC/XGZLCZ1oSm9GajumNOAxGacmyZo4VDhmUXrDuP+ar935IGyO
tIzPXIcD7i4OBxnJaHlA8NY8uBCGgAWi7KJRiiFVt/ug79wuqwnNtmDSgCFLLkm02oWASZJCsRrK
9kIhqvipK4SQEpwXcHTpurbe8P9vGhbneuUgir4njyAe7wAo5wsEOl2IlqgIpkqfJPO02SXFMa0L
3lzENAex0l0RO6Ob2OEx7okaYNeaaQ+4UBm8wskonoi/Y0y9Gk5qm53Q828FJbdByQWv95Rbk8nK
d6g9UZDa36tWTslOogK20pqhJiroR0GdEyCutFAg73NqLxhMp9Hx83N8cBdr50roDHkz2n/6IPV7
B62LY0bu/rAAO9Qh80hqy2x4kAuEAqcVNzIpyQAOqFslQrnyzbJW/QN2BgY4yzaHJ2Y4sSWmRWQO
JCnW9M8yRC29G0e6MnkgHHNMDWYSlsW3TXWn1fm0pgRAz+6Dcp/+qeJSvTS/LjhYU7vc79ihNgdP
fDrdb82J3xNTcFhtydE0/ucu/8+YLO49vHeEfy8EXgLrZefDdSCortsd9YT6O9fi6NTcTtHQDZ75
7SCQbufVBAwbCb72VKUQhYfHJdUI4gCFlAcWM0f6hiZp6aJC5nnrqIeAHv52hADjb8nIuBs6hP+S
+1jklde83nYJbHLWkBI6vjus1E8D+MKEoD5yO6ljwBW6lpjNMHZKCM4OGC7dEp3ykFXAoVOr76Cz
G4Rj3X2ZX4trhA50fl/cjk95CUyQE+FTVjAB/NnUCm/j06N35HOBxuQjsjRWjFqRmY0UwuE6edj4
rdj2NvMcZFVyKAhRsRP5yQmQ7TelISlyBBGTesOMUqvIbdfodfNsErgR4lwMDBKqY2j4SxMQ4AAL
+u11JxKrbcY0NctwT7K+irtuzWHFPWXNnNOCSbPZLkq/CF3NOHtDL2BT8f+M5KSl6nbFL0Tka+xz
xldoZ0AnZoxdiFERhiXRcNzX1QCYVXvPnIJx05AJ2J1RnLe1v2YPdpqqPJMxaV8/Gm9BtqTEgorE
ldNYUQLo2ppuqBlovNhd/M5wJ68eofH5bzcmeyWBeSSzw6XhGHNscSpJhS7CReKV3JgGFReMkCSz
aQtH+Q2bjlr78z2k5tLxL3aXdf5lMqgWtM67NreyIh+MfyPq2JMlpH4XJ5LEYOoU4KP0rpN6zrWf
bP2I99eRtTzODMmpI45Ssb14BbEzR+Is0jgkFn156tDidpl5cQY4Tolg2q1pfYoBqcdt5a8ycCKr
akK3IwqszYVXt042fZUjXSUbIjgdgur4Uuv4tS49dFqDepXh2DxOrzvrUXr55+hmiu6XSk9GtwIL
knFhOS+OQJ1hzq9aJH3T/NuawI3DYOmCSKqdPn5pW31qZNE+bHSVr/WeEdjPwSVJ8IoCLEI0srp+
XlKXlQ9Y+M51Vd07IrBu9rDrXfaWZyoMSLFyfVvq7iUe+nTVyMNq3Bqn+fyePupBcx95jDF7fAV3
tgDb07c3QJaLP1Dq/vFeKn14iIedfZuuORoFmSRBqPYdmTsH/1J/mOjIvFt70OnrnIHCqOIQRF6F
QlyeLCg5HmF5j7zucROEQn5/EwkvJ5Yq5gd3yLJqx4L+HfQpxWxvXsp2TKxc+Jq/8p+20AcBTS1T
Z1FMxjAg9iPsrwDPXHZoeeaBL20WBFnNPBMv6+qqCv7gZM5+gTqtLy0cej0vhABg6rEMEnLiSV1H
MZ0OflTLY/quY92P5ufA13+ifnUm/Ql1yGdww3Ww5KtQqBykL/+9YgW8rMuMNI+R//CBPx2NLvbM
rM3+tGXE/AmOpYgM2p/CV/n/YNCnyZJ8Eh2dUNvPXG9mGvb6K1r+6QUmBrvwz1Of3dLrw6rSeIx8
7oecfykJKSTDL30+P4FLhdzzfshaRHyoQWjJolF2zN7whfpeay21JT8Un3Y5WPxL4j9hj8DSTDZ+
eXCvo+N03wT77UJJ+HVgs+ebNJemWRCO+CPsz/mzaKdEGi2N2xB/3/vQlQCUhSO9PSOpXtTa/hpt
viUi9bnOJ89yoP3BS3O08pj42GvPdRHLP4vHcj91PYZdzc7vecjgogkjc34o8TQsRNC34sXj6SQb
1o8vdBKk1kQMteqJRt3lIRwNmFdY/oK/gK0UfMu9+hAo4F+vv8cfRpSgd6oKiyXA05CnVPvspBgZ
qTijZnFEWGP/BzmpSm0WzDuSpg2IOlKxxlFC0nVrpi/skyiz7LY2mImxM31Ey+lLUnOCKsTeHbkC
C5rLF0Z+ObPDR6XEVrpL/1dPe67NCrhQ2UkQ2zPwphX4F4DmOiePbAQhD7k06/YqlV+WGtDC2oSe
hYctgWpjJAGbGZX8ZPOtsiv/Z/bf3hXFTkAsafQL2z28dBoUf20yQ0lQmQPHft31u1hjWE9Vy8TF
6K0sm6bgLkUM6T/iSSzDqEgTk+LclmSRRZYqZqR16YAOM0G8y0nD+VWPJSJQAwofw3daNKYWVWy6
h7bBHuimZwIxz4TNI7OYPvqZFp9hS9BMsBDaai5Ft4jPyV00AE9irQbDG9SXRQ1t7LKyq7d1SJvU
mf/cQvLW1V/a+nr2auIf35UrRepI9kFDqnW4+cI42ULSlCv3MzNuzSWeds7iEyKHhHDDJHFpRcbp
1NHRSfGVaPyPKJVfe8gr68s8hFYBt5od6A4F0JSnUiejS2WMwiL/+Oi7n6uCmDWB+np0Y2GG5IRx
8EBwM9NtXOfnyAoMPvNDqB0pnutIT55TNyzELCeSp+wXuqAcHV5PaP8AjAu5NLXoYP3FTenzBdrz
gfB0FyJ5rjoqOdwh8JgbUPIxkcg15f0HjKvXCIETQwM0+U192JtAbZPHj+VmplDk0LUerftlumMt
e+GfDR+tB+6azWtJOmwUAnyQuGXx5x0iEbI2W3yb5atCkZA0Z/iS/lyaCbeBQ4qBlNyMNEokgPwn
DDzLYKjpc9QZb5s5ZaQUx4Lif3nvd4PQyKxaOskgNNdTnjP736cOE2En8I4Id9p9MT827nnTl6Vv
4V21yfRldQw/Elf8KxS0I6UhMnBVBDeG2Q9PANugRWoLFKUT9AwSR0XWnpEpKQHgA8RF9+pEZRXJ
9UaGbCbSJRhDHCdsG0cmgluqobi5ky3h3LLKd1veNHYqay1TCWKZ/1ZCAT0dDJukk+NTCsIGtWRv
GTXHdzDaLeRfqQVBWORPPex1LVsfAlYX1SB5nu4rNQ5z77oztq6lcRSgNFYkYD9ZPlCvreTmfueJ
2T7BK8SjZoqkufLe3T8AE1yFr7+rEg27R6wPnmcWFsUY58NLim3ogvgJjASWQUD9pvOa1ku6fZFH
Lq+hKO+vErIp6hEYSnJ8RfqARtOFs7kSotrfvLRIXt4XcQXcdr92qJFTFefBfl/CAfTUiEaBA5Ih
kwH2O/61xa8oBpYt1SqLcVswNHyEANDvXqpRzuc8YSSs/dgmBN4INkqlynpgfRPYPSuqz4mDhff4
1rtOMKnvLvaF3KXmM0N/qg+vUrpYU5EvQlOa6lo+SP7BVKiIYDjB7xiwbG0fhA4qLS2/cwJ1GAjq
Rxwk96uLpP5f6+5kC0anu7kIgUjKTPnY4DM2B6Gmxd952W4bhwaV+FK96q1lOED4VHBHtql+aXcG
t8YUNRA52iJVLOc1NfHyoApl+zFedGD052G9H0H3CtO8Pm9RlUjWVCjnWcCNLYtdDus47JP+j267
koVASeVEBbEWHjPEjfAFODAox7jrW6etxULjcO3g2N97p6coM0yGjNpXQAPhQnhB4ov96JltJoRK
+uuyL4UViZqD91WInuzL8xMiP1gj8eeyyz3CQB38tCDFIP7pTAJPyXDtcDGHhbpAFWhoW9SQUUvx
3OqsB8GlO8N5UTYClUpgcROaRFgUc6YPPOZfyOTiIQi7NW1zXhXoivUTIQYwmF9a/Hbd7BGOcYjS
JYXKY2lZ6cvGJeKAyGyiuDUyfIWvnUmaM6YqiIg0UNqHasjbojkhJOagKHHZuHoIcim7QlJLqTey
DBgaMAUJ4ggSNyk+YWX8cUxMBbvrgDBMPtCQQH3ymbx0f6KLIy2Gxuyl7WfA1p9y0iFCND3Y4F10
PaaB3jvN8hFVw/bonm+wxDVo/OW/ztTYkKQ6GJEc142/6B467z/ckRLxWPxPCWRDcWxfuhny5ktq
zAXwCSPZk7UpCJLW0qHF8UpHnbpci8USOWFz52OpQS02k9AREtjKaxYJItgT52gMU3AzpKaA/yB2
d/myGBYAoVC2Qq3D1h6tJcGExXFDgU2V0Y0n20zQeQdeRKxyi9DS5XxhUuP13aa27D/nhOC4sPOF
DmiFX9E5aKtkaKNrrmUk6sNvQSM+0/eAoqXeuNbt58lerce4ffbnF2EY8ULta7wC5mkMf3ewSbfB
ZkPSJ6mGqQnlvDTYW3RVfyIGzgexBBLvXRddfcTs79GWuk3qR7EWBilEmosOtIsfJXg633dnwl8h
DtAS+tlz7Qx0LTbMT/t3SCwTqk+xkjB79AZ0XQMvCVtY8b4bYh05EDrYbOk4Csp60wec+7cAuaEM
B6zNrN37cpQkmX95T2dOwLervdmN5iU1zH0zI0Lqd4C9m33Yl6iR870T4Bda7rGHlsJBwvkZKbIa
oYO5ZVsO0qn/rtustta7hPys/O3OxaPqg9p/XSToJY0CMtwi8A3cN5PFdD19dXGxdeIjyaLgDGR/
7FMp/f7nwTmZGnIHtHaAjTUK73yTrQ/49q+HHlWk3CgB2Q38EHxdzVYuitBVzdq0dKhr7FuTt2xi
ijrm420xb+qt53RHs+RKXYV1FJrgK7xfSZvHK9YdaN9FjFLTn4HP00syvLuzOlvEWE+6meyvus5M
KRee5Gbn38KyBcCJNtUut1zusLAMnYXAttaveWk/3KsFl9g41JEJSgNBFKutH0xAo1Ak7d1LVVIF
1hic6bAAexkAVCnm+nbnhLfhRM5OHWh5w5eZ2Jn51MlREW4e2qd1W37qfmOQVdwCp5j4CGBH4kao
OaxYTR51onvNYONh0aEWEBb9LkQAgR2yjOAfINfAriStwbRs/mkMkjviiEtpB6104zyksPi/GtT7
Y4WVn/R6mRY9g7wYpnZjyNpoYAT8/RvpxIpdmQHKSZgMy4IVrzaIpM9upBTlPwY3n/NWH/gWRer7
8OAwfaP704rDZXbdz/re91y9rqx5Wl3gSPh1tZe82+y4GkXZo7lqVYKZnPzas12IsGf/IN3aXLRY
hExpS9Xf3wu94h7IUY+4qvggQvlcO5y+5cd+3Z3J2gtCOwtiQA4iZNZxy2ndaJKIHwVJq3W/V6OS
s1laWQbZyzpitkBKMNpspnmsIHydzCKCxhvPBr8L4wLKP3V8MDuA5RS0kDYxw6t74tGxYjzyCJlM
XxebL95EPLb7/Xe6x+dq90LFdFh4nftELIbmW8hH4cxlGDJW8Qw+5kMieuEpO0Y4MY8ocLsnjaHs
5CgFZzCuD9QGcvHbHdyRzeh3907xtSi9WhH6nc4b1dBquu8OqTm+mfkfHzB05EDT0NrYrGQOSR+d
Et3HBidaein1iH5O7bqtS7H9PyJ/q0TYLqqn+tFhGJFb7pTPYsIgShz00XfnBeGmN8SacRVVSu12
qxlF/WyG+9Qc+wK/91QknnnOrzhf2OptLmKawoKw0bTvl6+8Lg1+wuz69gY4IWqbgfmV2OZ/NHU0
AyOTA1kHF/WWh35yK/595TUuWqIZ9750n0Va4q4S59X0fFp1IhebrrnFRf2mUXxcUFgYfaRMNMuT
5kTHy656HDJdopmh8oWVo7RcEHTIu+ZScHhbYbaPP4bn8OOEJItMZ9uCBqQ8poA8IWgLMaYXCfRU
ltKAdKpfbpQSM3Bvx/a2Q2pFXMWUdB+l/Cp4MuJxYqknvc/7fEbYMstmNCYPZCpqXlHeiLxvPf/Z
+4mMPN1tdsyZc6sMYskDS+UeGgKNagdQNTX8rYPPK39he8GNk3TOOlP2wkF6CvGmR5/MNcU4knKM
mrc5QXE1Wr9Ba08ra+R9bkFgNuNfUHK/8nH/8QP4inzmlMb2hQRsm+Qf2rfB14x+FrUy+fJB5ccd
MQB/MPb8LCND0dY8s5ULrewNOYc5LXasnvhBlKZB67o5eawkyBZEqrA/870dVPocdtcTnfM72VBN
vrI1UVi+xvfbleivRokoy58zq+JlZ/+0Y5cQa20Igq5Wr1iIQIO1v5iFppXA9PUI7lIrZ92StcJ7
OQtHPPbivmdWySzxdi3HBgdZKgQynoZ+9JLmeM6ax5CCf8POM9eniiJkBRzmU+CtZnN+BhzPygX7
RGoD9L4OnYP0ZdbwTwnnxhInNxy47J/qK7v99c9maVqOD3aOjRb5Ob3Hlr45RSuThF8V1zPtnVQ2
j/ytI6VMNa3H8cOKLVDE5nVHNS4om6feg//VVWQTPnoiZWhySPdkj1VUyulZeXrDFu7byeZqUJDw
EK9E1BwWC9bw397CYIFsIki06VrTKt/HwW2YK6Dqd5cIBnsKqTBsk/+k+X8TD46yDjRl7fdoaG+x
9n4hoCozTu1qfS5wiml/Q582upDdjGnwEIkf0GVqeh2rIKtPkzGYJDAaNYCVmtd2EyQgXDmrsm1e
YLImurvtTt6Fb85qgDU7aF6SNyG4OnwOB/nd9YTTl8kn3NApO+IDMOMetZZzbZo4QPLUf2gkdxx2
+0n4va9lGs+iBCnLBEn7a+p4dVjkXdMqF7kmeOa18DXkK3CwRHykoSdu+C5j0U1fAc/Z3m4utJeO
as2kpFKPBCZ+e6kOq0BPmJF5pryEB2CCEzS4O0/ID4B7GKqKv5W2HLxwaeqQJ/gLzHY2YL7VwHes
jNpunN95kEoItPQt77FMv49kYa5PWSc+IW243CDS8muOCbOCkRObWzPiWF7ga42O0g+ExdaA5tw6
cSHoubEJJQHUWAwEvMAUmhL5z1eA1NrXhCBLVC7jCVNh/PVIsEtmH+eyeeeH74ClGkai1dXIgCyF
BLUTFm3hEwaxJcger9/VdqX58oIso72fkOJMQleVjIB4YnfoEaNITuq+dLIagNhPmJzrQY1NCVs/
P8WnWkl1Vewsfhhzpf+YGDquq9LewZAfJiZHplZg7yHhgR+hMQ3xWzcJXeXybf1MN29BZq2GFKBK
VGelgfI91XKNCcImjiUEnkc/9DXXWwcPYtU3c6xeG6KVQkFatUF6mSjTQXpDhi7xXkTWtjiqiL9E
9PEBPO+UtU5BTqJcVFpgOX4/7ChWP4NcTo4i8CZwXlJvFNzMde9B8YeCdVCEcgNnowNIE5biZ4H4
kIrVmoToW2plh3tCqxVs+EancOai+uGYs0jCnukjwbkMEUmnZmFR6q0rqsfExL/0CSHgfKkm8Swj
/gLflaQ2oS5OWn2Ngqy3AejnFD+v+dODBe4MS2LZI7G3XP/zdGewDAAtAS/gc9Zb6v2xe4YZ/2Uz
bTdNcvKCtB8nti121//O1SJfajeUmGqL6q4cGA1aZZ/+3QfZuMyFUJ6ZxXYTiEE1ADoTjYOtfgrj
cevVNd0mDqfMe3n5vy2c1cY5VWBAItEDGLWZ892PwZFs07rgcwz0GjT0Rh4fD+x+Q9V2nrjIUgGb
wcSlQZPZXiEBfl/k0W/jm8azRLHw94AMOn3uRwvXRqJxOaAzwEc7+afK1K4IksjI0kcOBvnF5uND
PQv2FHq3bTzpqfjb2AX3Nf3kA1LyS/cSqYZkGZOzYr0NgnGIXuALaIrlj7hIWYjykhXL/czOioRl
kb5o0m7ka6bwCCCuDVIjJ5R9xnrtd4Ha4kbd2XzmyBMFGVH81ufjc+0uZfmw9t1OsL9bH5otzysD
ruulkp4hBOEYM5A64niLOpCWaKm8CY2NopmDwR5pHrFLUgctb38QyogplwaUj/VHJdJKYkCSgwC2
Y0JYh+jOhSJRFb1RcV8VGy5/ba+tvPZlrXtAg67VZhP0bGPICrWAmCujWmXW2PrtLuP/8KKhpNYW
tWqSHPCIHoGf75CKEcApkba1R7AuWhn7x16GWIlWwGp5eJLNmWwL3r/fKKAdqlcdeSMa0gnN7+mW
8nRc8dNCKooDInCWkXtgwSBGzOycadvTY2Znt4hq0Zd+o830dtfyOSyk1vxSsxX82BEujFxNrmX2
xLQCs5hSCmvBhykiOGa+QGLPyzvcbgSdIVKhj1t9mR8sQBIKPnT/z65gYmn/lwlFK/0HtTEj7I0B
UfCNSZba45xI4DkSqqIDnrQStqliaepDW1Q7pTmLzbk+gTjCKwyfvIskRlYoOqrZNeWkXS/YgpEM
gcP6QS9BaxHI2iqp1efj8mKKbX5hxeFYc1ysEmFVUfA7xK9NUbVxu+4DeXj77npWB61vtKSYP68/
XGGxhQ7HC3DXSJUIM1a8oZAUCK3iu24IaQ0DPsMLTHY6Ql9dtlYCafJNZxy9+LcpzAr5xeOpOTCm
IubFfRLcqBuuszLcqIPBREhnx68169c5aTWBvUZ2P7yRkee4hwBNvG1HUnLYqhAjCAmUMVgBjGsT
1Z/OMGmnr6eMwXIeL/WCbm7bCwyKD8p+xai39LYGr3j53nTpRl+gELZiAlX0DWGBQ9B2+t8Yfb35
CyvfyYQwgMSv/pAiJ55NcDN9M5MnQIRcfCpcteBHS1/XLFw6KH3LjZYZKpfLtGgJlfGPumE5OMV/
L6NnVeYU4DB+6izfi+URrHU0vVIlra6Fh58IaDT14TdCJs8sq3XEj29RLpDZw9DMIXtsza4FnlEI
Te7gkelYL5S6HN5hshf+rsIk7N/TnMiiw6krcRCRRDClYKoBTwnvaBSXKXWCvZtMB/cj1sK5+BKz
rBr+LxfughvL9tIBde4YIJK8OVZO54Eow0QoQ3LoIh40I5x2/GKJAaJ9WiQfhjgkZD6X4ict7m5G
rLsO/EioP8Wxzk3NyXOV0xYIaaWzNp24ZXpr0zv8t/TWr9EVHzAsERcM0NXH8uKO2SI0Fgj2UnH/
MqmEzXoNvidwcNy4LIIgJFDyxJ6YeHxb9/+FXXl0wCucV/DPw9VmGMPmFM8Kk6EiunXiuY0z7nXa
ZZI6QljeAI1YHc3rH3CNa4TFc549iB4eGwbjsJ14ouIhoVIi4bIKNW9ZkzRhSotuHy/1DqqAczev
3j5Ce6w4lVFUQhxdjuqTPLfcC3WReoEY/HhZC2jp1ZfNJ0MEqMVmEe3MeP8OzznU7JmoHGk5vvnE
CcKiCpaGUimOYTYdrt6sNXl5ZMBHt7S1xnWkan1VvIf6dGvFjMkg2meGV3/R9a19GSV4fUMW7RNf
4gwFBd9yneSQF9ef4wYWY33kuyMK6qRUMZqkreorZFZOL1EdmXNT0CMtPRtPijBEYnW+l5+Zzjjh
AbNUAfQ6dxWLI507ldJ4wzkvd+Z8nDhAGk/2n4Yn2OErvDfMHZoZJfxC9f11HV0rxYeGHFRApTk+
D6JQ/F0K21nxV8Xw5Zo+EZSzShm9gVyQN04KHR3wi9d7mYkFCfaFMeFc2GOW8mXr3GW/b3zPMwY3
EF0vV4vcr9+szopOgDmicIN0s4ihBKyjvvRy4UX+xuN1PPHNm2LDZpifc8Gsf9XDqeciS0R3CsVt
jSjVSLu9TVmi48wsIOeExTKL9K54g1x8/PiBLlhi8TgwZ9pK6SSgVvDFrbl7QHfZANUB/nyhRowW
+fYpNsikaWKfj1UoK7KG7RTMc2Wzwrrgry9BIXxnamL4CYNtomJwcFNXpgm17g7OnDySAiz2wMAr
Z876j6YkdHt8/oyPsB8mgn/WIacXrWlnSVCw0+KDLH17ow2Lhr8zHHCMj1PSCr1YuLvpEMuUaf87
8DVct8vqWWUCWcCnqUQ2KW7WOUi27+7bXGFRmUKYCvMnfLsXxB/WO8PRDQPyrUU38DBiPNxRCMxW
i4ucxkEtyBY1kwqppmjxwqa/KgHGNoTGBRW1jjoMOdBkB30KqYB0/ESg9Q1CubT16ABcLvmkRO02
OusazjwHMXq9+wNbCpIwTMLUmuEuwoOnM7Rg/EHS44fktG8mys/lIvvVR7vrL6LBjZeWpZqIhSGd
qs8tyqOt9bgvb9OCX3sG9F1dwgaj57ERYkgNJ9eO8YRcYoci/3A9j+HHp+izqwoGBRPHLqDsOFLL
7EHqLZgASSwxAA20rI5baHHslaDwOmVCmssv0MvA+HBjTMPidhzOtsqZuWgFxKBk/NyDyxmTqljN
J8xXfZ1xGkz5IVBn01IUz6Fqcn0ibpvof/iZMibug0BMqf7DyAwzrbRP9v5809GV4o6YS+bkALoK
HKRm7wdmB3wMiKC4651kItsviFvl3EyahKIpoleYVv1FalblPhl1J9okS/6rPRYPO6CHmwWIhQwT
fpGWsVddJzyzg9f8UWhobg/+qxKqWZlWLHhhlphba9z6nGyZgJO7Lw/RiCcFweuTsmTQV1vE4DOo
NNssR+6LOdUmXgoPGLF0K3yUkjPzl/EsMOT/S0EJDYshMMkMMBx+tV30D3IREjkMKDad2QyUSr7U
9bjZbEs4QyEK6+V4p8QGzUPLA6zSWVOpYV3Gu3gBBenlHN/Gl2uB2ULLUWlIzAWtaWdkLDl71tmt
s2a0t3rybFuSRa8Z4LHJ0ShfS3n8/gGCo3nTp4+1FSA7sgFnyabyGeou6v2yjX+PTDr/EOAOZSl1
HVloCFUTmCdPtcqHFDiGUubou3TJHdIOBAnND03h7q7V7wtXP1g4M95Zqptu0tk501Rd7S25lyYa
d6vCr/61o7KSVLF1ZACnvNNn+SSQu+wWbXZqXPS2IvH5v7YPn63N0GUeBjCdZhnAaCzoMToB45ew
Mw66hWg9FkQCrzyUuy4ibpjBN1XME6bazS+GCKOvhpUzDIhaR7W8Tx7D2INQpN7tN6F34KM+0AFH
ZLs3Cs/P10jD4JGvmFc0l1AVb6dBYeB0jROgMf7wWpDm0FzNur02DzoKEXIqkbJQIyp9tCoLkFfC
P1RWXam8CyUaP85Q7R4z1MVYrZsRZhX/FN5up2rrYaQ8OvX4uNYlfpB8K8AZRwXnEEceawIrzLP8
P1DjIAgl++QIoh7NPn1Oe2g6/xhbcgVCRO9P5DnHTzyYzyM+CyO5GDw4dAHJOcTLnw9FM20GFKf+
CGnbETHeuYbVbO+6HdBK4RXv3wyUKDzoe0VNzb0cay43E86MJaWXOP+szsYF2q45KVka3BtZrWya
pQBijLiPt/P0Z3OkF9jd86hKKS0WBzNMUFBhfkXqNUKa8gtHWMmiVXEdGC1sqV796XyNnj/erXpw
IJ+hD02j6cBEiaoZ9xtrj8TiaeuKu0bEazEhpwwFS0XBAMXdPpKRQ2cqDnJcEYGvoiL88ySde8F8
WllBbvrKrCmrwwXS1vedYMZhnnMYt4CDWBccm3XdWCmELyQbgUT7XiZYs5b8BRjohVQ/xFfg6Orn
HvCKp2gbEGzV99DF353S1HdXfIlcYRra7TnnbazYIZqhzBU9KvMCoZOjGoPGCGW8o/5DtON7zGPb
FwXy+bsViAhPuDYb0Y1oHokBqkOp5WVQqv31jAX2blj3GY8D/Ns6hUMbsAoaOvCGUvKGEmoXs/OA
xTNMxxPWR2h0d7gqHdxBnvdXxCxrHCfB7Szqc9tEXT+llrRtYUSjWzE7wVliU4Qi+LX9eOe2Epxu
+CQtZNttL9Y3F6z5nKrMCCdetdf2GlsovGWUXJX8UwpZIaFLX+IjtQKq65oMFet2oHHJdVNH2wp8
2SfLfEpG63UzdQyXMA3i8yvGO519krwFFI+qqBOHnt+xvmcyafEUSp85wpLl97MxFthR4D6IQDOM
sTl7Fc4B/Sob63g5rQ//lIRhfnsKuAkbKAAb/I2TfE2F4R5GFJghAq9ygH0dPJglHTu8Sl8RaFLL
auFCtu0e9xh5tIlUBVDNHC5Z2IoGUK4OpY9hVZDvl8+ysnmzqzzm8Gay3gInu9WCTY5zSm/gLkkg
6l6lPrQd3xRvPE3k/wAoJFpFiZ/RRCZfdC/vlL3id2A1oB9cziBycy1DcjM+Ykt1QaSNp8QVXAUP
rH7X0q1PdG/4rv9Ogzz7hqTYIGSDmOVT3vu/SEq3XCgtnWGWB6mBzSv6/DaVGN+z1nTDuDW8b6/2
mtncBOtGXcFF6FGAPlH/dDTcNLF430SbFoAxGEvapyXltBsUHwhSBOnygiv4DtcO7buwG8SPtCx0
OgYkR6w08lfbaZfev1e3zDmCgAERfxEdkNAMqxEfBmkfzHLL64uKNQyVtmKBS6+3ZeUfij74c3Iu
yW2MOQXA5U+wfPgQG0i9lTaXide6FW2XkdSvHAvI1KeIqBsrG0GBSKbXGxRXCTtjVgaP67ugvSEC
EMln4hqllvwaTle5kD/3ZuUk8HAl48saewd8Aflqn0Fmkc85g53H6+PRAN73tS7nQReyfTO8XOGj
pd3gFRiAInWKYQLR8bItOnZX2xwl38WNiNEcdYxAl+erMW2KKeCGLyjAGoXAs0LGMfgkGj5x3VHC
QdjPRMvAgcDQrpZ/vnA4QKdx0ez9rBB/OPnxB9AYGfY/3L/tM/a9S9tQKoQukVfJoSPogL3Rme/F
5R2VNtR4B2p0oVTK4W3IKyZaHOdDf7l2suRSnnA0ctAolRv1po5wS5GmhOZH5Q/XsPZcaQT8W5ao
KH55AVPf6fYnIPcV3M8ndfRqzVOz6mHkn3xf1vHFXSbIyt+bwu1GtetOrmdk5x6yuKjADDvofgTQ
abuKly8sGWBnOWpN4fymqVZxNU8MXWx/PV+XnKNUWcak8RJInMLcybYjdL/6BanqCJqBO4VHJusK
ccpZf2jrHSFEenCMRGEPZnL4Kx13v2S2pA9+BTNiNNJHtOBF5q071jLktRDuMgUb2aOHkVhpYjtS
fgwAMP2q6lciuptJ2f8Eu1xyfjCK4YsJxVAgTpM4S4VwnZbpm2xo9HvqTLFYPjDUdyKs7ZRQnBIh
5/pem0ToVZHHj8Dru4bwFP5tuagPS0S59gNtOeToszkMxeRiaoxkwAmWiNaSBACt9KO/XuZOSMJm
yT8In8VWPwVLdlXtLQWL4gBbnA+Qf6CrFWJF/5LnPKTRlg8mmaFcec931p4dxjEKgLeaEJPNrfFP
3bDh+KBbof2Jgl0c8zczgHHf8c5nhP+eb/Dg/GrAv27E8qVpemILfgVkQDBJBiS358fNYArSSayW
kyFsqksVjoYVZ5geO7owopx0AqGra4iVmnv/x0G6oH0P3crMSr5PGqvDuPMiCwMVyafXq/GUf3Py
Q3D/oHfMTlnm8tVZqsAIfQYEuhYCegQHdEKOL5+i4RWo3XAH9us4xM51U/FuC5L/Eb+cSnvRHnFJ
ZWSFXKLnEEz5hue6FL23wM4HN55MZpuLMNSbKpbBVtxqUuSeu2okDo/66HAD3PdSEoLC4UW65qjh
26lT9HeV6U3RE9DnTjJX8yh8vNfwk4n3r3Aun7UYJ3is6NXAAPJvcJOfI7pgquTQttA3+W5M3z6M
NaPMEa5bu+YiKHidGOi3Usw3lWsFFeihOQszbTJ/L9NK2oiLP+HrG/yCMbr+z42jjfpMv7pMxnBE
+q9DkmAOe6B/jGsRlXquRkMCAtHD50eyUJiO0fGVYwwszY8RxJXycUAyuQwvMdIAQu0dIfqJ9OHE
brPs/gN8hY4x+UPT8Pc5LGCcu2oA8ptMK1n+Asi7XRjeoU14+kvxjg6sA7X+G/nam/e7+ujye1W0
WP/ND+Lpb8UX4WGLR9H4JPkxRyyQg5pZPqT1ElenmBv1AXDX+aRXkKoc632p1KRPPlwzxwLPirMl
fZf/ZLDWr2gi+WTZRDioVMVyCKnhW3ia5yM/dUp6eLQS/tjDhCYemZv8iPELZzfK1qo5KoMLk79i
d1yJj2S9z9UGO14Vppy70XPr/XfzPoVx1NOi/mp4gcaZUp7kUOuT8YaPkME9AKXA7x28sySgyNWV
Fl/1nMygVUYjPZmXyx2T+qarSNac7CxZHmIhnSXicysutXCaIlc7aL+G3l2WFhsou1EtXM+d2uJN
JBTEqTlb+40kWfRDFFjXVUctnWdAeBb74YBKyPdDz2bmzwiggoYEt6JdOTouonw/x2eefBrY5rHN
fMdrw0b97bGWhsg8AvJDS6jwwy7GkWtjiOKl1gAqSbY5jFCfyFglVvyd+A5G5zTLLF/gBrSCa8R+
tlun6qLKrSSxJcQSaHYinJoXVe8VtnRf/Nz3yezWxeDu/67MAX1xgnnLy5m3nkyGqj4OUJjZ60Jp
idWgtPb2y+laEReJLShuTKYCnM5Je50bo7dsJvZQxS5sHg5yHnSeDVF9uuqeOaFgTAYVtFveqvJP
5V7fT0xuyuGWiCKVP+NYHuQtB7Zb/x2zgkHABxdO3F4dvOLFYa+Z0slupuz3uWeKaUlng9xWsgWJ
i3z0RToI275mvjV8+16w5JZkJCoFnFNNGddNodzVSMMAqa6lWikSt2ywjtqNZeOhankBIOT6U0JY
ShwKYMiwwOszLE77guCR2c1KHz3zgDU3etCVwxMp8Fnx4g+/EtewEP5b8WC+xp/w3EqCKxxslEjd
P0WEcqBNXnm11s++9S/O/SnV7cC4R4f3g7m3mwu3EjwjaWRJqG+VSK5TCPTNBBS5uZESQnDFv8UO
Gw7WaPpFNxHyf7rqojSEMDSqMMFf4E9TNkZcYjbzw6V6kDQg4LxlUR2ZjPd41ft99HTRhyAWv/bc
G7HzwyyCYCAdpwgxauu4T/RXuYu9JOKeog3SzK3RDS7JvwBn4Nk29YoLUNPP8gE0sBrCw3pW+FYK
VCVFgr2bgXn492X0mpulwn6fqG7cr6RZT1DK3o/CXUd8mThyQ/3v0RVc1mTtOz20gc4AXNYnJj5x
umc7gQGRhBgrXhZAmWOheW5EGL/1tZxjqQu7ySXbIgWmdomSuMOqJWMrS4vDG+EOnpGJWeJMZycA
+QWX/gHaQgHLzuQN2JsHhICxHVobWA2QiD2L2znIzuyIkCruBLKV+oOG+RGufwBnz1PHnaqNcWJd
kYY2pj88iO05NApcwbwX1VcHJnsXDpBjip7Y2nr6RacJnauAlB14DcUTgeU57HcN15IxXes4Rab+
JbxKq9gr3R3nSBz0Mj1l0kZonSaOCRXCllFKC8Z5qqXLyVziIk2paUSCFLS7HILIFlAQYbl8eRM1
WzQcIum9leM/lQ70X3kyjuE5WTf22I2FI2cukSgwCqYhPzne+aEktxZMmYcfY1q7Xj1rI6NCk8NG
TwU1/fK7x98LjcaceNH537snSgrB/1QHpL+DzQbaHfGvaqDub/RaMpTZqKHq58/RzTC8awhwNqYp
z9T3kZGIgZyqmVr4/cEbLf5HUVlDBMZxRsMh64NMWE3qwJvDEk6F8TPeFPic5Yp6IGgX2w1GK6bu
EIYIeqn+taxNRxTLhZB/CaRsHG6xGhQwWFSSzBgMmxHuK1vw+fT6AK9Hemz+XgkES8/VUirIAP5+
bJEKmy4Lv+Rgf1a7L8w3wXFbeN3M+3jGJWP01X6bEwsD2+EfFrCi3yzLAiPjBEHVRsLQwz8nGh4I
+qs0DufCvwIYe/zYctMUIQ26UEnJhaTChjzwLkG1Nxdo8WqBuKtu69qniAfm1Fdx+WEwhQ8Iy9Na
dbtkQ4TPYTYPEPRZY7MjoVUFJBOGktpa3MmFXQyh8zpkvJjRY1dQ3VHtJvJsYu8g/igqLhGJtJjQ
UNa3dpD1KrD/ss7buM3bBd8ij+Ibx5SPMNgCbHVWqsc5BMkdXB13THIqnnA9V4B5u5k7xO9farHM
qxH3Fk2D9k+bT2EXiGmGwinOxv/ESJ5S/m4zqCAtU837IBGCFRRckJS7fjySsjVR6Plxijf7Ks6m
UubpkKqiG6hyf4o4xQpQcAhdyVLZHrZc0Nw5nOcwKpWU9gvUf5LjsUJ43SbW7Qt7x/iYi6b0TZpH
EXAvmsIWdeGXZ30ty3wPo6wKOD3mCEZjLd/u8IqNUe+2/P5hf1M2kGe3VICN+ovbNCR2JJYpwzqg
tqNv89gc106yS1BwIF0Rh8Vu6sZ6iQ9Jqf2u0n5yUY/8ZDqGbzn7Z0+jMsHB5g7V0TrptrHzc3Pd
vn3Kd4YzTBXEuzIk9gvvhAgjwzigndfdp+Wo/e5XNJgHJktji81b8r9aB8diEJunFEw+j6BemDdz
4KVSjwbRtia9yXhfpVu3Tw/keOt42iXFjHGC4LJmlrM885y5GuVh3xoR2VudBrodfLn+ij2+mIZb
AqDs6J5RFPV/mH8PqP5EH5+kYFP8v1cbKG5lPIXKcwnNfv8hEvtMAzRoRDsW6ddvFlVJRQF83u1J
LJ9+ANtr57nTzcdctbro0vcxY88zyn5zWe0FbKwlNBpHKXhlsobE9qiLuI2lx6VUFsz4eU9FlHOT
apyphW/1vQ9YdmXm6gXUN+myStcxn5gNwa2r1KmjcVKiXPXBNUf0AEdoC/34dnjRs+kpzQSVj4Ka
k8WV8RU94XqtIr9+1yqYmh8OvO3Z4Pit2EOk2Ln8ivhnNcT9b8g1AhQLyhc0ItDlbLomjk53BXV+
Q9f98i7kMDG341HNF9/epaNZUh1czkbGIZOzFJzAzBoJzVfvCdXeObsc87y6CoJdXr9Zb0clDj12
AfCxpRMEwVLrzIp7UYHYKNhZ3xdiShIX3sIDGPwtG4I8HSf1nrxEA0gpyb+k6kYwYXFOspLi+l2S
FuSsLHzsi/511dzHBRuS95w3uF/zVm6hWYNPfWmlLcRwi1wGIwbn1QRIzJccSWwNsYabts0dzNvD
PGhql2KOrL60NaudyZ8ux9ruhTiefWf3kG3/CmO8hd1xRhijifi/QRaHuIOAMAYmH9uJbX/pZl9a
fr01mCOOZYu9BDYoHdy+tRacLl+SbQouCJfZweDk2smXiMIL1DMa5gYFbn+DTrTBBbsDY5Tn49ja
eFzOyl682oanUvlwbt18BnWT75V2wLbUTKs3Vls1MrglCrC9efHBls91qJ5bXYf8dcoxLCNl/BWc
1xryp30CAsBRWomOLTprEqXiA7TPpzqtFKIJgAJBnNwuaDeLQAVKMCnhPQOiT6E=
`protect end_protected
