--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
GgrvRSM0dHJsdbRUthyQcL0Le5r1DhTMDLOojXRCZ3XhPKJsz+tksf6UwT0My7uC+HD5Aqvlmao8
5+mnmR0MbCIZVfkaQCpfpkyC6NNk3G4g9dAwUjNIoelST52iOYBdkjyvjwnW/h8Nx6pFEtCU9rcn
vZv/uhBhYtP7ivynzfdXdP3iD9h6acL/xZFIIzq6inO4gO1dLwZ3orAyyXtJxLgaYjCfyuNS4/Mx
WfidAKiEJaytmnvedTH/ePl8BHENzFRi3WFDV9/VDZyUgsNuO0fJhn3m5P8Z8j0TeeNF5ry68evd
USfEyA7QRhwODYeqQyyU2S8sBnns+UJZ/OnqeA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="VsDx0wxCPGMh+D09l5SYB/ae4vR7bcu49B3RexZjtjg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
PbAD7MaqU3Zab/BxABIkmvsMD84N7KFqvEt/Elv4umgKNmeeUZJL++8lsXhkHZCjJA7DS6k+RBKN
jyMOVBKc/EuHP2W3Z0Z6Ece2XwXJegoTi2XGenE80dFYUV8MUGp85gvY6fkRL0Q8KxPJR4QIhWxb
iB+/nIEOOq3ASzr1jxLOZOMltOixPkH/qZ4tFDIPEZ1G0YUuRrz03VjpP+qssminZal7SeMnexyu
KKM40WWcqv0Dyz/6dw998qHTKEUyO8WED6C2/6ERU2L1MsEfag8FHqqaaVPg6vfxQr7gecw3XV+6
TTKBXgOTOdE7E2LjNnJ4w79NjUP3uCKyC6OKag==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="UuDG50y5rrGisdcFGZrZbM49Z9zwHkciRqkLvGhwGDA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7632)
`protect data_block
iAZEEbM0BE4feoBnnYjNttcpapLkk9417S6xlNEGGyCunlFY1p0mxvxNNZEimKM1rSUBxwHF8do7
uXzlG/Y9QzlmTZ/Ht9Wt0pJTV9DFpMDa80N6vPI/dtFPgRbwmx+CXdQ1XGyue1PNm3yV6bZt4W5V
yy+8PdxZBYIi3nKF+Cve6hpRMAcXMrXVMtTcglxtNwTwJISFbVid2q97Vlc9mHGRIOS3uI8Fn8+W
zlAP7UKsL95Vjv7Gc54Su0swDosxIuhDCD9HAEVpzWP46rXtpCZ1r/fEvMQ47rbDws9O3KTvIdl+
sHol1HdmFeWqW/Rgxv83fc+XKVGNh65HAiH3B3EAgCNZxVugkGgWXmuuxACtu5xZXZA3OlRjKF6t
DJfbCE7DSt6WxiRxNdWkvF5HV9eCcSHIHmOZAlckdFdzyif6OUEI9E/ZnhZtu5RTqT7xVJ2JQ+xD
QI63jW2cf5GbK0sVpuOtbSCPDXRS/qQZdh2nDprgcTPgEZc3Yv5FQnJ8I/DGt4ueEHLhuymefwoj
EwOi9NH4GfsAo07fD+oj2KLhI9sTizUwClDstsWzIvgVREcL2Qc57SFYojC9spSc1NsdJVzmxoWV
ZT9itAemFwXopCE0EfnHJa4Qo5Hr49OzDjqFYVyXDH0nUoG/VPIA+ziLu+m4Ere6ag9gw/Ibik48
0/SKsBF0QWqJktHRfQk8szHGYFJAtQpyVevf6z463ZUIHqY9JCz4Tuhy0niXNsEb0j6P8qPK+z1D
WLOLcoqW0sNqJFMceWNIb9Kx/ZT8/V7lF182NJ7/MTt4Q+LnHeTaL0AS9p/jyXLMUa2v3NjT34Zx
IInomarIIe7glBLxKVTjtGO3538LJTEXPLEML6cm3uua6hDdqYpdWPdwXhIb6fntYXXh/AEkWH+a
e/4ODZDKZuExlzSYdDJq+sIkaqjhvreV9OERNfgyZLoMOqQnUaLUuXrwq0rSde4T7z/qe5j5JHWy
cIV5DMcY3vsvtbazRF12kt+yJZpNa8/D1F2P3FkmoFQ/tidVJ6TfknlLnwavoaoLwuJQzBqzWdeM
4Q+4usQ+IwhYhrsfhNRRh/jwYkqP+u6fna85VqGP/Lataswr+dqvYsdcQxEwtpizs3AoaSvtJwuN
wPYoUrONqtH2m90+MndZsEQmyvlORmIVzlFeoSZ93PqL3oPvcj0pMMHJBQAftfO17o/OvlQwaJPD
XiVTOz4wKIwWW8mEpSs1N+uaa5Bcd5o2AOh5kfdfjT0+ov5TlADUmoDGxUH/OR/Jm+jLggbFwIY8
k9JQwV9HLao2wfGHUShmqC3EaUpTX6ON2IOJelkF8pl0U9QXoqLfnBz8jhI4etJDC4thx56S2iS8
zuY0pLAm1K2kpKWPfT2fFZi1cmq5OJe8d91PhDqvtUqoflbk1wmrsCDfQ5r+F+RdJDy8r4sTN1q/
5gtvt/jGNt0jH/+e2g3rSKICyZmKkRzWAOneUuE64TUSod2r0utFIDx+UFzoK1SCl70QxtGdvgUs
Xmn9Xt8hMKVKxizEaj52HcnfMl+qWOuaDnxr26M9FPmExz0+niYIqrBPm9koi8B7Nzk4mtuDcNi4
otTmzV86fmdyOXoWxFwCDI60tPv8r9Bquh+QJYlPihbG5m6v/M7jqnl5zPzpedJVkrJ/dJB8/jVw
0vK5lK4qFg0wAxtFHyH7JfJLxGXeLiINXstdy22Q4CVyA5wcGmtlEayo+CB+lISfncNuqR0h93aJ
/hmdCIrMW5sQl8bMpNxuifkG4cJbKcnqgc6PUSIIZ3EG06/YZidtZmeb3KUF+m1qcLbH4mU/mhNi
Fyyl4ReQ/nWELD1dXkVkbe9si0++ZTKW1QsbH07PC38KdHNscvcX5BwYFh9FLmsSPzEeONgLjORW
yKzORFnYFXZgTkR7YKY7RECg620YlT+oP6+ta6pQuQj+wh3xRAQFrjvlp8aK+mA0+lzIpwr8NxXL
vMTrt77d5eYdMoGunrLVD9qe2RjX6zqosNlCJF0KCsVXoAOzZ9KJigJr/Zz7Kc5ikVIIT5tHslyM
P0Hh7cVnVEqm2HbYLsfGb6GW+18VhdEd9YyAPMXR0Lz5lBrpiv5mzD3uyXea3Tc83oT7rfKp+Lg9
va3yC3YscgWJvFophlFGLSIggYhbVzjPQSs2kO6Wrb0pIiwWZj5gKjt5ENJ+IMowmrVU/QxmYIOX
+Q1+gGkoZ/xs2StiuJKCjoAPWJLzvlguZZ2loGpKkTLK8EiUeI1Lk9oUu/Fek9WCgxZhoMZ19072
A/gUojXsGZ9L0fZJ5P2ShaL/VzuFswPFGupBiCsOQKnMT5l69i1ljo5R9qSsdsldU9URg0vDvqnx
ufmpJ17mGw11ao0nM0ScY2Fv0yxY6nVG/ygqlXcwlv9tXH/REc4QcpZw9fQ89B3vcIepRZvbZx9T
+TLDUuuYC3fh6qSv//f4e7isZDyRCjOLp5EN3Xq5zehkJw6/zbZLKCBYZMllTQKMv1/BnhQz1RX6
shGc4f6gOAyM5r7bdjZ/f6Mb8Azv91tPy4DHNjDqrTAZWFIj5wN2vInu65Bw7naqaI6sMr+j/U/i
uNG6HVdUzYFRZiE8NcFn9UAAa66F0m/OOA+z3EwQ8/W/dH8BwOv9ugpL38UPqrsas73Cpgqy7Reb
Vq2cPi/HdBwKcdo2dAPTero3YNJHm6S1vyDyBkz1kytA/kBbPC6bWv/lGhrCHh7IFh2bcSMjgrpU
AD5PhmFCzhpi3JOY2QxCSnk8fD094eIvDwr7xizj7RzTLXRs8imV+xUeKCLyrae44JNVDH6PetSt
de3UYFtncXp6gbGz/S7IhSyjxqZuhWqBcLWksa0rSEfE43tI/p8geMr2RkYhL1Bu27uY4sEkLIUC
wOChmxrAI8udVNtb52EotYbVSzGvg/ggqhnwdSyeino7u1gb1LLzmDVCKcjUfZkijjPbdn0PU83/
FFYEWb7x9Xd/EetDRyMRRmfMwMKIjwpFFLwQzfQKUOzQjkFdsnGltdq50JUYE61j/DwKMIeje7x3
ucQ4ZiN+N1+TFpPqbLHvkAxn75Bv+XRwOE8dUBQBX0Lu8eST7M7Dpk7gkC7FQ3p1nNY3leezr9dr
J8HG9dpDM483TnkJSwZDo7teXz3y+cXPoK/dBJAPqvA7RBorOBH5IPGf4Gv+O5wfduiR2r5kGTae
uFZ8bAveoPZX5BL5T73rZDnD3PLposOSkD+CWszqiXUqGfPY02DyTLWnSKNz7l+XhAVA3fc7ECOk
SbiG2g+C816tDW0Ep6vGoCu/8XgotfkQpyQfBroVhfYyOo4zkukgAm2RDD3j+5Jvi0KSAs47ULap
6+ZJSXRbTObOTD01EGnU2RYzd194On+UzvliCnHNtuRtdtufQIj7C7nQZD4mFlGbdVkYvsRHg0xE
amxZz//2yiqq83BYzVzS2p6yzAzf5BzU9uueXoOmiyZHqzk/fh/KVNvUmxyo/NOl+VYWde8QLx2S
IAZrFrjg+AiIsH/IWQZzbtOkbPd5CKfboewsqwanzXQW542An0dm1mbki8E1mnVUrICiQITiEEYi
hGHpHvajWyVC0ShZpFOYRsWuH+GF9cZPE26KH/WwV+j3G4FLKX86V+sy0mMx8WIXIOec645oE3wA
feGKdci+Imm67FjDHxGAGDjDTjUfcK+m3wju+DqHr1+nnSxTgIoUeRTnTUMKReHTPfjGyLlNORO0
HZAprVZgKEeKTg9TQw1qMIrsQizTLdpnEXkoeITBcho3jgLGgXr0Ldsf9O7+QU5NGzcu0a6nwZlD
BH8S3wN3WFsyNSxNnbV7RgTuhy+2iXQ6MaUxAKspolM91JIFnlQ7bAv6pmC/Mhf9/fJMA6FZ//Ti
6oHtqKURYRHKkQDbODPO3GxYla3ryBCgzKCP5gqYGi1hnGUf+AEFxmZ76UCbCRMg68doDZssFdTq
piSuR4i2Q2PnS7JYT97BOCOIVFE/dwyzgvuo95fiLqF5iGsc17/k4Y3YLV59ehFkenPAPCt7dAay
dhxjS5+jyQN+HEwlo8mBQxMywTCEIBKeyWxYaau7m/qcb/uR6juzj0GJnOn0Uzzt+iU7YSB/Wm3O
HQsX2uwfc0O+7ooGPjwcKE3fyrhAiX19y2htBHJdiK/Q45Qjz9HpZLa2bHpc4x2K6ux+ayqgMjBs
StUUhB948eMEacCXO6EXAr0pCJh/Vtyh4i3MiE1G0wP8XeyeHdY9ynIYNwr2GwEeY2stGYh0MCUF
yRXWy7MvACX76DTy5WB53dpSLufZLX/jFuQ33tf+OBHqnY3QVNu1yFrH4llyEMuBBgfMmiWjHcGM
4eu5K80EgSBPFFDEOIWPJ/DmmOWzehS2umGi/S7ocVDw+1OQ/RQBVi7I+X6Gu3W95mzNtA8nIXoo
iF9IipLfvL6Dol3zVzvIR3Ne5L8iEdeXHc3iSZ20+wCGJr4IvZR5nBrMYv/X6ZpaxulxUL6jFGIf
TH2By8e29E3b8u/9w0yidioga8TaNWXScayCSuXVGRPw4srWygrF8PfybNfFAIi34P29rr9cm1xy
Q08mOhISpkfXezNNP1mgntKBC91fQKXqL3RR5JXwYXCXcbFfeaiLotNoSZ4WjaiVNad7Ue2kandu
iWwKHiY4T6dwxXnwjZlyqjX0THHvLNdXulRPfVZ5vU9servd0qbS+BQfHb2uPPncDWcU5kbWSJ5F
YOPP6dSxW7F/7yRlQrJ0I5n3iMxiNqPAqN9Uq3ot6OTaRXz6DsooxyAP2MUn+79Y2tDOCrsNkf0a
Z1Lw8s0MAwvAlJeNgoO/7OPak2D3bv7Bvp4eYYNIuoFJctBE0MJzerK8ltzCbFQpiZrHki6wuAta
8ovbCODyvET2W7JBez9mz24/LvgKUC+SwZRQx1CAYB+e/mbVLo3tg8HOpvMTDIzesBkwHSZepTMu
9tqZNkdJuTKQHmHq4i9U9WSUtsYe+g5S6bG+o9owJK1D/9COCvi4ierdMIr5xHi/JhpbmERQz3a9
McDb8Ptmu6Xg1oIsRG8wo7tiBn82qxmcg6pmPrC0QDGXqi1pfnWGvMUeKmyOBtT44h2VI4p/Shuy
+vbiE/B6OAPtVeXA50d5s8jvl8M+aNkBj+sqNxoejmhp0Pt2GdfviaNC44YINXF69+ckyzjdpxCS
7xy8VbsvYT76vrywg+psDXp0f5oT8ZXltaN3oIoH88eFPUQvNijbVMv4fYoRg2TpJNFcqAEkdS6A
J3TeU2P2Dd+kApAIozHT/SkHjT7LWuQIxR73bjFXFBGU77zemWb7Ur1/fFIOOD7HB3S95IVeZTZs
tcoXJgKbA53tEjwJr9BejiLaLQi6XNljSp1e61UySGlv4ZlE/WlVySt72vjoExu/ztiA6Czg/89L
5z7CbOaxyHRTzCpQGhHRXmDE/7vpyZv0iH74ylmZ1m0PgEt8G4yr9Ogbg67zGyl0coRJ+k3vEUue
NCvJx2Kd6ZFfDRq+xePmrcCw0QZCau03hdzzIrK0kLcUUKjmrkMvhOPaNfsG7G0Z5KE0wbmjr2sc
QVWEuH54iHX2NM8VXKVKyyPCB8rVoRA1xo2Y7uYZHwOy+bR4lLqstV75F5DDJ4W8h+W1mpMKhI34
iif/OJNHiPI/eNWruwCArzNqn8xVWDBz0+aj5ZIoe0No65c4lwRXmhOmXJhSil5Gkuj2cJJrU6aS
DQ5xvJCYAN3IQ4P36PjFUJ7RMqDsYKQ1OFVQIYAgylb51to8I18RyNDm5SCvKpRQIjR7IOXXVXGS
dCJ1oMeFD8nk/CD9DSj0b3HuJHfj9MlVp2ppmfPsGNxLq+gJJHXFwgOgnXlYiEdjCWBaqLU/glic
isLgNb21Vgbm3mLjLyKXxMSD+Ql2e1RCjQbYCJIEiUM4aBkIyXrZEoObSgi3W+MYiF8FQRyncwHT
x86FZVAoxxa70N9c/bLyzJ+2YvRc4naWU6KtKYmy8ClTRRGMsk9Fqx+6asSByOj9PVYDu5QQi1mU
yfWZX41j/k2Y4PhjZ2uP6JKEBzjUYHoGQ7pc4eyLkqjEWq01Y0E5kAy3JRqMVc74OZY+zQlqWM6V
v5z/0qLbVr14lCfqSxnMp4ZoHuyfWQNZsN4yfUGx0FavHWmQ/nw2MtqKtUg2VugDGJ7o2P6KP/sz
w8ek4NvPE1PtMhKsHBQNNnzyJGzF4qGEgz5nH7Th+206aA9g8xDbSFM6NdbqeWY5NxL9IPAZavuV
tm4r78IPmxAuN5QUAIBUsqPvurJYbguQmKK2jpmLwp5rZWtOqiLbTDDvg6BreCz2W8zQk/YsXUIX
ZXn0mPXtK340e7yDiziOtmIQopvC4lXM2yd5LQ55KWVzrAihCVR63ujkRi77S6PyCQSw8jt5abFw
JkJcPqEf14Oc2v3b2OfWpvuGl684MvHqe8yP6nQ3xGJrH+4KXXqkwIkBfLeZM+1FSoVvB5RMxhSB
gBUYTCXbUH9jI4Bd9EsRFNQxN9SBegDzD/J7415hjj3aVYl74uchpuQ5i9vMk8XlFdHxCK1dFwIA
DkURryuQNVlAXi6Q8HOMJtQ2c4fW2ekPgZQPRwkiCeG+Y5UovIeLx2IocJuFNX0/PfG8m4vZfNUA
vge5SbxEGPwijY1D5t91VPROmbBYbJ4xWsvaKsCxyYQ94NCn22EJ3+PYNlDEkVsle92kfvzEXSd3
bN8f4dxTJbv/dTnoAfxomalWW7PW8rTRC2Igpzw7o/KG7j5FajGlJq2O6vgadn01uE4sKoyWUZb/
sxsjfrKKoeVuZKkgTTAXCsW1ucVNwj6fH8xSlrQxhP7lhiarXizXCV1SPZrCQpBQuLcfOtN3MZcw
hOd9YZebcNw5ENzPJG6rFu23l1/XU0+9PwD+surYMDIoaaEOk4rmCMver9I6UVECiO41jqIBKI6r
/QUHZC4PR/BUe7WRTHKeWryW0HHp19f/jHGkX5TL1bSGjoEJ0wVbfMK2RDjBxmz/7VEEx9IlCULj
SdFv3WWYr7/FgGR7AHbLD+oOzRtb3xSV7/JSbgrBjgdy0syRQvvCkZymERxmQJ0KDOmBcJqipvnI
nRrbSmhhDbRe0IYEdb9YS2M/C45VsfFaNQjuWipjIlZzL2TvmpSE7cyjS8KRPM20a0p8Fv9XYKzD
vVA4K8oqmrgy6MspQyrVD6r+4rZVphozIB5A4trSXk7L8v78YLZ3cI13f8sG+5H3ROTFz7BtUiGC
iKkLZHFnyxJJ5zK/xgrH32gOSLjKo3f6fmDH1gaWsHuSpf+xCWFm4E9DLQEvnM3h7e02gewk0rm+
9XEU7lhOGJ8ih5icJiXq1l8RVJmQxxsv1PzoGmyQ8bdd+x5ry8fiokiPL+crscJtKb7H3eNGp6dN
or4V+4GBU2HjqK8tpLtFwpFfLMXr5GYge6N5MGbHSfDkFC8zOIt35vqPFTPIPhknGGY9bPRt1g+c
wcPZq/2Y/lDB700aV+jQR516Q8IdQmK4nmZbOvDoXdv13K45gJYKKqPfr0bV1933atJaXz03+2Wd
8fd36i14zte2IwLMZKqRWCTjSik+kdaTAmKYfr3y6WIl1t0SEP5Dn9jLDhrrZNxJvO4popIehXm2
CGTFxbGPUJ2luS3l8k6uTrMUBThOAOzvVy1qYeVjo/KHHUrCQAJUD7MvZD6MHk5D3koLDRBGXMLs
uFmIgZcX/F6og8KMsyzpSo7nHi/Y+tywqqBGBb+/1WBdqPFO/BJk+UouZ3nGzEYvO5ukgiiVRNJ3
4K75tYNMnqztWrpqXThXdTGWtZm2DqR0ucVjRngliwaLNa7y52gc8JPk5yiUfGpX0EEjQrEyyg18
kaFAM+4T8SlESNRsrLoTw4Z5LQAtNvqrj4tISIQZShdEFVBlak4lxP/CgGIWhXYUOQtaL/KKUDu0
OzWCtrkHrAlXAxby8xBs62c493YY23mD7px1rGRdGuaJ+20FNlJzZD9tDFN/flvy96m64g9xdmtY
l+yZUARHaeD//ti4XqPCGQz0lrTTHI/JjCDZPV5g+xNg6aG/NYMXnnrmH2IPO5L+dILBWhk2RFl1
0noXyfTZrxM2fRSo00z3bocl9Sglfa9by3NO7e5QLpYZSqZQ/dRkDVq1VHcHp18sTrzsa5Kq9qsr
/lzeaXZuZ2hvnhleAEEDw0OHcRknNok+ptS5xrnIBHCFZmVYkBJjox9S8B9z9wHfZnyz3w1WPfBo
Xa2CWW37pvmYQNi0K5jm/jaEqM1RFjD+OvAHCYWpvj/rdlhbiJdgC55OkxbTkoSwENZHilQmSGJK
llQBmJbJcJO1j5SiNYFA4hlw9fbexTBsLydP5IhZ+bWUuqqIHinR4qyK7E6lkh/3HipVnF43S9sB
87zw8ND8xMa4b9qE3rB6a9boSTEa+x0GWRUoD6Rw2Tv4JmyfmfgxAf1y3TshIEC3TUBJoHv2C2Q8
K6iS9GgejB2CXikJT2vGrLx8m8CKES/HkAMig0CFD03uwWF2OQXkSXYY97bLslvV1hRXkBmEI6ql
PbE0BtW1S1svHZm0szoW/D8YoRjQUJAG1dhXIxNcu9PGnrlcSbmdwoh3TmrSVzyO9ZtLoO01dlmh
RDmHsrB8exqH4O0X3CTQarJEzCigj5p+ZMXpqZG9UtG60a02H8n1v7XZQN6L2+XJ/PLchjsSvayY
IgFD8HvA9v0biPiDQxtypdru5KidqynExzfIP72sMA+hZHLfOsffy21JPdrBINc/xX98bfoLkwDG
HgBJXR339s35zuEcP60YNECMnyLOHUY2vdmfubETrK4cJ1tnDmq4ZNhuw3mMqhGKORNpvNtAAlbQ
QtyJfIP8G+OrSnmwptI288KKSL5xDg13hjCT519NIKcWLoD/bzbwU3OoyFgrb8adyNyTesGP1RmE
Sb21lezRMqjSxppHig8GD966hFBzT/aqz/L8a2TDCYGRmKwexDgNiu0FTkR6kGS+YlOYbCMytZj7
AsoOO9uP//4Ugck8QS4CBeaxwZId8A3BQ6H5PP8Ff1o1zus3IUzvbdThwDb4uEf27MGIuFbz7jqM
x255YxLqA71nT8bAQ5d1hlh+cojI4+mxL4CqltGJ/xLHRufG19sBJ6n2S1G+vqqGDjm0oOe8g19g
2j0t0pUu+MXnkm2x5f7Hn2UAmQbU7HDh/tzRlzz6ncd4tRCAtFFX3hlEi5xQgqPrhMGfrOTxty9R
CIAnNml9CFdslGMNvHSLobU1crSpOFA5XMJl1LN5WOHlwc2Porxv1R9W6/a4WPqivbrBWuFSL9Js
KmVRL7HEaWcbOGAtURSnqXQ5lN7hnkplk0uljm5HhALmyTQxYlkDxph43G2VQOwcG7WYeDxJ9gtf
1L+m+zqjZBtpNevduqnKYCQ28Kkaai8ai6v4Kgvj5H4or7Tf8iYFFp/oTF2XnJlUEFG9H1Hp/La/
nIgC2op8ceHvzfehdSrtgf3nHed8B2iI8bNNe5InLzISCgsZQsM0fqwlgykrnpIqGCqX+YmhSrlV
FxJJB+awZHM3fxcsZi4Kx1eVfJaLSXcDaLKwEqlGU/gBtD2D7rhPj5lqMH2/RVMpcdqxZwhLjyut
BtmAwFxyAA4dCYb3T1o/rmE2I3OVwhztpQiCEkg/GAew4S4YQZ3rkh1usUW7z1gWYIMcb8ly1JAB
s3Fsi0sx4XWD1R2T4wI7eq8tVAPHhBy09h6Co4qJZzL3XNYtAVrVkPo4C5AZ34qFL9GlibeWEKrV
5XJvVA6La/Xz1IeuBImkAfIqTKb+bRS+gNvRLJ6s0F65HkfVh6H5ZR3Eux+bXyZX4IB5jLgGhj8x
vLdjhHwB+tDRPmyMXNCMsniKWj7vKCNFd5l7VtlcGm7GjfuwiBvawAF2Py3X2ttq7aTYzqUAphte
LXaQVzVKVa59SVJY4jTHw/R6CefnsOP+KDG0sjPFzvjOoUzSOH/bEQLC0j2n9K4VcnA+iIv/+yey
u8a8HQozua5SSj12+eyzQVpywG495I0omE4QrubmdOWJGAVHZZEC5+05qy0EpN8nh30bejlkrfgD
blm/klyuDhBf2sanQJNGHNIt87ZBscLx27itW516rvpj0FI4cVSyKv+qQHJdGSMkbDzVwm/ZqInG
eL2ICOkqE89C7xss9fePTh4JG8TrYf2I/tJZZbw6sRoFBjOaNZb1Fn6wzBMVRuirQQ6s
`protect end_protected
