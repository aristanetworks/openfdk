--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
as+jj5C+LU1P1Xexc7cyHdpL2BBGfJNtUS7mUjp5QH4D0EizE6x0uW1RNo8GJRLV1WJn753iMLae
2y5VgSB6a2Zolf40Rtp1EQOUKGp92IHalQId0ZSZYDEjUiGvzHPN+lzH8SjvVEWaS5dVA6XheJJf
zAjTotbfFuaUUpBP7YzgWM5lUWn4FB0/l0ZZdXPhERONsOvPUsJk7OHA9rImZhQcUBMam0jAN9ro
CKjBvc0kPRrIlbIw/kKJ407s1mcYn8+qg6S/on+VOqJeiskaNoqXBKnesCGhk5hHLYHbzIeROdqS
qIOH7EOMDAglpTRPSYWla7vb6LUiHmly1ijr8Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="YRuBTxpIHkQaArKtUMBy3fIhl0X2gxW7jde73f//oZU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
r0VGXFN04bpGxkUHE3gkHPJ5vXSK6/5JEXDaDUtaHa6VUynQwmLNh+pNkTRV08NFOYi/0y7z1c6U
NybgcXG742LGJ9bYkgP0Vvr6my/H+Oy1C8wfYj1/iK6ClFj5cc21xmYlvZ/dZokWozqG4BqecFoK
4yTETLgZPjqDW72wZzFDDYd6qSVs6X/712g/+VsU3RZMQhc7VDJ0KUJ37tBGBogiCO0jtt9Rvokg
qp2CSpG0XZD6WlxsOixS8dtw9b1Vu6JMj65imYyg06lfDVN7AS1BtvpbY5nY26QldXXB7c24Y02D
L4TpQremHL1awYTPlV7egJesbEjFvhYfFek9sg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="YHNeGNkSOd4TJyAZ9+HBA8zi0hRerErqxQlOSKjmsg4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6624)
`protect data_block
spfUuauvi26ajnRQyI2j7746f7xdKmTHm51O6fGkxT4/i1l7jxTZpFHo6cirPYIaHSVQ8QLIUGWN
vtfk5AMFnhkWalkMaDzLmykSYK7g4qbggD++w6yvCcGiCKUS2CDItNmSjw10te+gvmq2RD96Bzil
jNCngpGVXq7sCsUq47qBdIWAcKxj8T/3ecEwgRPTdF4DBBNaBYZJobaXGdjLjMWD3LQZuwqs653J
CLC55uK0W/plJlMU5h68hsFz1JAl6A9SgChTImSAUtEiPwZDr25d9KxhndyFkkn9BVcyKACwth8w
JVhnex8qhqL6TJ48+j4zwFJ7PzuPKbUZ0DYXU8dNExXz+RvtbSHrVqZTw7aSXvUHBJOOz4JQdkzh
9vRGVAe+tbCq7TyQnlhuHved0YKbsV6/ZjQzgr/uYT6WX9DRit8/MnDJB9T3SOsB/7Bh/AYmuoEw
KeNOD4PbHv++VRuGT3sKIXSQ11a01iOjFeZiRr6A30wsMCtu23RRZT7amcrY969AoJc8zODSzm8A
H5CTchFxNAY8wQNXfPk/y06fEdszMoCtQRXSnYGEDeW9OBWIwLtjUn0XUDvEGjrAX2xyLP/qwjvx
hzhRtUfojxViaZ7BB0T1gQrY4oPObkt4t3WEObRG+lQs8cKov448JLotQpNNqaSIe3erZB2dF8j9
VegKXrboIcZ5pUrP1bbXDeLTfURxarBhvfl20V59qjUCrpb/WBxs/hO7W9+r/XLDh5T8AN6hmKkl
PRMEruN5gVs63tOdfqB7Q6D+dVUqimXcbSosZhx9MBe4H376M4c9O4kTILWzeXWe2nzVoePG/A0T
R5v13W08tQ2QVW6sHjIQ0u1x8ZX+by4jYaBEcJNAMMxwMqiijp2S4GBZEQVjAMPhhREUjnmFZSR9
7Q3sxZGgAxIe4Owg+HC1853jz2Xd2wGS8hGFnEfCNXP/5xnHwNtRR45xpTNMCfJ8E8PagQoGHRfg
Q8EuTK5HeL53SuWy7Ko9N64KGZNroOBTrQurN+s4mhB/7Cae2Vm9HORqLg6NvHKaaG2Spp+FEz3F
9rg6cw0gxrGDx/4PDYZdIed07970Ea4YelYPg+XJqoFHnLPdIZEdM6v5lOc2CZBdZPvOL6PmP8gZ
+gvokwJjBj57Ck7hmG1A7YD4NSsS56JNdpXmQ/nP9xHTkZ6o+dHmLl8UQb5JqNEx76f8vD9xtx7n
fzVHrDb5tN4DGYP09nIbuU0Sd82rrKIZNjVi7ZHpZu1cEK9lAG3c6MaH1m3A1ZWSmkjGVSMRFdC7
2M0QwdAo7PG0spqEsIsFg1A3p119F1bI0f57uUh5ryhooFITZOvFHvFWHjyUtSeKFh1KwdsAeYo3
7yX+PUB+661Lw7m8k2DWuBMmLo+dzNK35JTTB3q7h2pIYcN8CmQUNXDJITnzfR8A7lgPecfPtUcw
E+pQOz7g+Z0DvaFGw3Ql1nIgtuFrrTwcV738dQmiGmASRn02oNwLzWfH4U3tO8Ga/voHcpDsJPJV
58xEzOiksN0eYNw0tj6jhO68CwOPID2giJOlInQ0EnFWkjMPOTbuXZIjkrLoiGgFmM2e61VhS88q
Kdgi2Lr0cZblk+uWb5l9WyWJ8Iag8jvzen1eE8Cj4RT5JL6Te4gkK2ahuCugwR9HoBj1gdDybpZF
bp/vQOQ7ZwJ0nKKhwhkHSebW/lSh/9SBEjkMHxM3ODTXIiZBDOsjmKFkR7Lk/x7Wfb633qo3q6lE
TnyCTptWxcm8rE8v4YKl8rV7XD/DV4CCoKav9TtOW0BOuexL7uD0wg3m1jbm7+ikrgKNssGwEivv
WjumXENAFuAHi4sravoPUP7Y7b5ef+H5TUTZm/OchRITP975LTt5/o5PWY9nztidRGmEKQV6Q525
G41SRjfmLnn6VCVPtcXaUt52myBWvuK6WG+vo5j/cML7E31bdY1OcwkCJjWJsYE0Gjqcrr/k6NiN
1jNjpkoehjcGLNzUxSeINjH7+25P3sti4uWH2o4LgXc8dWfto/KBorLerlKTiT+aa6EkhSp8UJN2
GUorjxNT6uz63vZG9BSfiOowoXkIJqOLdA0lCZ6C57/PtQ30BoxfW66qpZBnSCHRcd2U82Aew3X9
Z/iUFnA3s3oJDvViwtgdRNmGlL22JwrN+cVUdKdRJBYPqUmMZg/AnXmQ+KFKSK/iB3LXQSFJVi68
LddGW7cX02zFr9rWh2M5XfH7GxMzZw9k40qMU65dpfA5iv3FQxGv8P+9XV0FkYuVvHxX0dB+QD54
sWX2SNVdhVAdPwdOX83+wVE/3mu0OaS8alWJugz+6ZNu/SraIqDMD82i/Pw6pLdhj92JU5rU4iqI
iNyWn7/qcNfhqEssVGEbtblEWJJvSoIT6RnnNc9Gyq2RMjZDeiObgkHzILEhKQUiYJMogNY8t67/
NnY7V8oW7YcyeWXdGqox2EHAJ1ZvJz8fshJ28omM7Ksi7aKyYXed+HdDMATa6HSpbZ8f54ja0Iom
Pqlz8updW0WuvUIAYmzkoRAHocWP6jcoaQKxJ7acbxwAB2/BxQjNQw1FpuxyfsZ0/bmS/nhvPt99
VrWs+Z6Vgx1uqjOWwrOrfdKtmPDdgJmarB5gwdvEhqFfpeiBjpgKKRDPCS+rrIRohOmh//E3NTZ5
EVnoor5JqfPx1E/Vog2UD/rQH0DTryCdrqA8xRapfFDiz6tKHgFxGQaq6lnY1L2jOlPpIC27oI1B
M+FnnoY5FprB7POronIx2VytEZhRHvmy/bQlB0nNOvLGU9+e5CY4FfMNW80z5+35uUduWEitNG9a
4ucidVOntHRRqB3UfaVHJpnZmUdRa4kJ+MYR6DT+bF1hBRjizx+KhOrO7DV153Ww3rfF+AY6wyuZ
yB+v7WyMAnfsbxsLsdaYJ4W+01iFgITwwV9Hmrdznh+I6FgEGcFshbWqZa8yJLmHZ/UVOx7TxRLR
HptUk+WBboNofJ4A2j4ADvoOVDskFu0w+jtw4Mb1U81GBkmB5QQXHvM+zOdFlQ8k0xjytCrsSBCO
29PGqEEE6/S4OMkWR3W4ADsaPekS1sXnmSgQM7Xm5ySVm2PhowJ9/Udbx6wrNAWghf7hjfXRgdzz
ytcDaxdwbiXwP9C1p75UabziMb/ss7hGsuVt0a9Ioz+do9/Q5g+58e4bkYnxec4wbkK9HWWRFloL
nnMB0j1YZf0UymFWjoNdNK7nJYx2fBLsLeU1jlmRNlPr0dbREpoiDxZJgVx8O10B4sxOmzd3+Di4
pJQn8eXTS6r91QiusaneZzKq8lX8sMeCmDbGQWIAQeqhFGZCNLRD4jThiNLKmpcHq7OK3KzNraql
DEQqFy3hSN3mLGQRQXtYXQch27uLafNXXtMEV6Ygnp1firmN/mFrmBZ907UjqOAcJecC51HPNi+K
VORFkE0RNRv3u/GWwDqSXfx1ZU8Dt3hOMwtiD5CVf5dnQhDrQSDVGj3UCbBMOEsAQd2/q2gtiuEL
TzVpZpcYA+xG/3hVyTz048R2HDbS76KOO/dIvHbyY9N2p1Cg2ErTrlLDpEFfIYoZCOZl5tmZefJK
0LI4HMKKWItIY4BU3fVv/3r9s89LWbgVuUQqlRu6l+FP2mjH0me98iCyeqg9rA0kS22SWQbyY4Y+
9WEJlKBfBsV4aFixDRMqpETiz5PBGFKvdgHyvSBTW+lKOS5AY0sBF69XBS6LamtRVHdVL1dCFyz8
G12dwhK/JeobpjPhotZ/Z8S5ye9pJCErBFkcIxpE+t/2NpZWTuS8tn+sYBrAH06ZZfwQSh7jpDl6
lAnrfx7to8wT0ImGNaUWT2Nx2kPWzsrjGZHlYe8N9v88cfOD2nejh3fy+zlDPNYuzzurrPiUjCyU
rY0bH4IdbHCguAFAHwG3HVWITmSME5dehOx4WqLD2I8FTgiDTEAcL0TXva0GZtL4GSbeQIgeoX1L
khqEL2L3Nh6fAGKve98n14uVmx/Oj4I3AzIjALgXyMdGqWFh1ht+GXulQImqJrTvaTNJPUx/kYaF
vDuy75Td6HqeZVwYRdX8Fc7tQ3MYuQ2DJJaiDRSF1JWxy2AUFE+MZRD4udqSW77Hc4LwQqthEU/U
2oMOxi+BnVAOwq68Gq1gFI4jFWVAKUAfrce2Pjbxsfort40x7keO2WPcZbC2wUtXBw3gJUZTC3gS
x3hdx3dIshSf7pKWj8jOjgnwl+Ss/Zg4Su1JrRfL0ODU2lex/rRFzFRZhVqRspIzCLP3mmG7auEi
rQOw6J9NVYtgkOe8n/C6leoOK7uI5cmLxVtiabqoE/hn7cwmypLa9wbKgHS/2CUfLpNIEc8W3LNx
FLNVN0k9Ks/tnYUuK1JYIUEo0dcw4QfN4QcaA7eeeh3pWFAl5B3ckMqctT6MwIbA3IW3Oll1CIoO
VR7HWINLQZRQyiHEisz+6b5JyBXQO+VoEN9mkm38q/YEyPB6v9gHEVI3nxtYll7NadILb5QEqPuJ
Tow3qpL+E3CKne0hGPqBLzPwF3NaTaFkM58i/IgY4FUX1DT0a20jX1/39XGvkE1O8dd/TPm2nf3F
bdzl/nP9p6phIpvdnF8B9aGT8l0dR2NZCUzcqGvBcAquC9jBwOMY9x4pb5bqwEvIgUtIxS5aVxML
WEDVddCmBRVUgXKWYz5ypNvHyPI/E+MxvDo1274a0EhX0Kmhgr0bTqS17tdzenc+PXaKJWTMCOQF
iMed/HBasgsAJbsB1x8D01R7wwT/5CUAyhS//yAZtlqnordUi2GBhyMzNsGhZgMhc+ftrpyh8llt
r7tw7LKHVf2igRyDeJcylQ2Da7gMiw4bv87vqTkRM9Os/bVm4w2gBnMgZnIuqT2cXWIcqrQ5Y7DG
k6M/f+LWCeATY8P5BUf480iRYkLWeFURNaGwYQaFcm2OXv42wkLfoZe7c/kywbj5yPUcgoH8twrO
OBIp6YD8nxiBw6n9sK3OjBkxSga3qQDkicYCpzokN3BEG2jHIWDaVyQZe6s/flnE30nCul+U4TWc
Wlh4Apv/A2GTiTPG2Vumq9qwtAafKw7Bo1v1JsKtqlJ9jpKrz8H/u4howZniphupLZmb+TPSFnm8
GQL1Rl1WVqiQvDigrkhTfafSUqr2uScQJ8FTZPkiPYFdDvAumUrqdPs4bxaF8W08bpb7rnnqdDO1
hmrIjvc0VinM7UCMRTkck32Ci3L8X5v++056TarxNuoa/2KqXu9WVLwKk8vHeY9GoA1/giCBTGXk
X3f0xr0Z7avrOHh9+M751C8BsA9UbrxJAKv67pH0nLKKe9WFG85shvgiMn9okXXt6tLxVSIr0kPd
HOa5Eq66tMBdzRsX1GDzIYO5mng8lbfk9Imp8xtuBkgs6129mPRlKLmXun1TSzYazUpl6CDekyU8
RNcXewtErO/S5TiNSQdJfuSih2ApV4hmrIbz5+5ZTsV7lKlLPBWDTkV5uMkg9AQv6PnS8TOu+oWT
PwISGgTDMyw6jrLRTr5IvDEqc46cK0K5YufGXR2A1T+MvQNra51WQHlGM8PZJvrvCOk+KPT6by1j
jZZyVgBWyQvV50f4gjCsQVjv5pDIcumvGh8j5yA1oGjzMuhJzh/guC3l4Owrsn2esTSzPBROfxmr
gmWzftlkEPSpvRc+SnXxgaHrdf+nn13d0vQ7gQA3ziGsDMYQ9dAbuMNfb9wQ+QDQXagHFWj5ACpN
mTVZ4X76IRKWTO4FqVkYEyfl68mFeXvok8immEcwSbpGxBg2tZqC37WNYeWKaZ7mrhCeTSJGt6+9
I69CmHDLmF42ru/Fg3kiZhyQima4/mdYcWYtjz4tONCNbMtcFiPtw+S+AxWTmm9yF9NgabYC3IWY
WPwH+6q8rkD42DNMASF0opoeJmd5w9RBUdnNReGZcdDUStQv5X31h61fQzj9c6EmHdrVO4+rsYPC
clli6iEGf2l9ePsF87Uw3oDkFpUMbWN+6FlGGi+0x8qQqi2VlzdBfoLQvEl+nRiRyRxlxrDSeqWL
pMpeJwBHQgw/QC3zmJqvOaCwZFSKv5XEotCp3DPm75OQfsCvOPnzdrOfFAM0S+4bROlOG66DkiPp
/crmtc9aT/sQBf6a6Lm5YQLGJe07Ovyta1ZzSGCqo9buTSsTG8fhXf0vbfeEIL7EbeeQ2XyhBf/B
APsVt/p4FBqCCNI95KTmc4PaZhuCiMp9ctngzYZhUNeIW5tqPQBaDCPAev/wkF+Qks7A50cWl9nj
uldo0doY7LB32AAoXdT2DqKXvySypEGrl8uDcq3zYNvoetbEQTUGpE+z4JkWPz7Tk8TEMP6ImE/B
XMNdxCd9txCf3Tr12fFRS7UvfkJuiSCgH+YnlWmfjTsVUhuIDgf2rjvTfJUYKl1/W/+TXY2dt9kF
bvNcoT4J5MeP8GJTECgTjqjeJ6mh0kFK/WLY7dLlKOPc1gq5XNeXQwTI7bUy0gH5KhM7Uuq3CNIC
bdAgWrNILtbpCaMPlDB/DrANZDrU1xBaP2mf0dfDbyPG5It5UcAerhDEuHHdsA+pFSRGrZrTn4pY
03PAriSfxiuWmAxyaaFG4OjLdwg4RijrV4TUKpMnD9tcHGeDbWC7Lyz1EDb2pbvHoGlvIx/pqgeU
mI4rm+Os8LAELP15yQt4ejxczU+Rlg6y0iSS5ujdIVBRZik4pOalQFKQOEySGBQ4aAHCNjiEyPfs
wOEZESbJCBBttShpA0NhLQ4ZfGAAhlyzCWc5jnCbU20/+U+/P2PtYU/Wv6KqFdxjTKqyZREz6/zr
KxbEMfJwIcoXkdMcEPy0OKKFPyORFjR3IGMbozR2g6QZaQBnm3rNmkrQTc5/aDW44HQuOpWBMlTg
TLvMTyVC+oTzthSOTFtjhKNvOCLBnjewQoEBZuD8wdkpQAbXI74LiX5R/h70bIR4wjiC9GASPG8J
g3ecvWuTh/jCH+0VOiNMo/f3aUo0Vuz3DtKky9GMr6NMVqKJgqRzAuMbCS/g7H24oDhppUKuQkN+
bE1o5Lh4pUkXJmtra/y2vUDO6Rt3ik0WXgh6nxyk4WsRVcb+acK93D6plqanIfDCbiinbObG+/oR
XTmXXIlYlgvivJMxXMm8jB2zdGCqO9lcENtNHQSYoNfX9mjS7iV3xUNi9Ss/e5sFWZpmORKMBzoO
E0Hx2bgO0Yv8sjM0i44NzqKNhiArE16W1E4DK5r42n/gktvwsXp+3WTGCDvlGpuLzA0E5rggl867
DuG+DShvpTy0OHucbvB3lBN2YG5YrjiVGC7bHkXqAeZ2o7lFaht0ooPoYeCvf8OUP39WFkcu9nDo
qw4MuJB6h2pOfFq10LZ/soBzpuUhPeEnufSh6V6m/qCH0Fx3iI0mMxCtpg0f3tmVEsfRFdNkjp2q
Mbfmx1eIPI2/Da/9fNW8lb+0eYtLfP0GI3wBwJTkQHOaP8kJeE2/QktpOuSPxLFFf4qyWifGog2/
TvjdU+QmruhsnwO7RmITohddmvTavXbSuNWDml//WseUVWCA4Wr1BCci9sdZWAYaOb7fBdPIrzSw
5+gKj4BcNrs7KFTahJKlHCSmeT8tu/XW7/c6Y3lp58Or1wA0FasQRI6QPubHO+Gpuvy6Dnj6itCW
uhQ6mBRUqkhxKhgko6icjzBJv86nGNGu0sYUnyFnXMnF7Ueebd1d8DI3IWinCjMhoTAUwXKmT8P/
w9jhNrSD2rYdHswwr+pQgMuX736dmJ4SROTgx5YHsO1O0qCVMAXZVGhjw0OlEwZhppGfMOTh5xCT
JVT0D8z96rPQxph38t/eLpeYm1dzaCRsV+WiaV3VLVNXkvC7E8EjYaGS/7Q0mQfziDXE+B3cPEd9
7QTSLBbJAJDY+f04WyxrEtKb4DZfGqf68yUTM4qqfv7hjAc0mZLimC6Dz00HqQLcKAa9n9ed6tS/
BFedxbWTer7aJDWfzOl/pEodtzbYOtM/hpafYrbWRK6N0cEB122pls/hHEcxcqtGlczAsknc0leh
bu+0Zd56+f6wPC+hpC1w/L8YWHjnL9GRU5hBHc0NPEoQCqDRxhdh1aBTIGzRDkfhSA8dO4BHWIMO
OS+2y7ilMx7ti/Ut5V3wn0ql9nJ+JpfRy8Qsv/J5uEyoMmWBZRrSZHEUbLJbvf7+UVO+djT/f1KX
LHPoJ9oB1OUeCUb+4zbbe2opVbD406Mh+ElGHpcr8OIn2fLY3416IJgkv/vfM5NwmULsrSDcnMud
+c/r9/sN+P52rZrUdUmDG67gWi9JaLkNF/IQwXIicuczAbdfyI6ZHpXwWA9Q+EWNUYuGiWmfwodG
2AiwWHOe/Pp8EIiH1qH7K937lh6ruWJUi+Z2rJf3iLFFSHjAWBBaBKIJQfPYrd7l1NqulUSEGXnE
xXr/JZyokFYlv8X9659UUb6YkvUkdmXif+hGFRAWg7ywPGJ3Cn+Un5IrLjEk8kXj1dmpF/WB1cyN
WwgCgrps5T47poyTLSzUMx27L/Zyfq7ljC0KwbGdwA9X/MRnbo0wOz3PlGkR4IVriaaRjPYHKeM+
9/0AbGjSg6nPP2zVV8liHZbbmn73Swnb4z0+tkyTjiiFL+7kofvIVTi98Wz3oRE+F1gEf3O2/cbF
io9VsdEU/RlgQC2L1xWpjUQ9WJVbmtReIWqYb+itGciyQS2JC8M8u5+dXpk8EgSh6lzxmuM5wacX
tmPHV8l2xhgbHxwAWRPCshmHfnmtsquHG6Rhkma1lNEEjrctmfglrZaGo9g7/qOSVMNMFwoj36kI
oxANvVTFEUhLf733DtNWMLWLne9aoUx8e881IyA2SrfYuQOO/wPP0aWg/zMeSUKU0UD1CTVf0zth
zCccrLw1JPi4WFxy
`protect end_protected
