--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
mZ8OYxjEo2VfKB6mcTB9f3XkLBj4v55FJDOAcUO/GIBZlKuz5OHhtuNR4/zFQHh4nhDvRKG5zODB
MFlvLEDH2vWOJOgmUCZyaFUlRm7zEwAn54drvGN2WoiR+6ZQcbILb4T5xiG6q1wtq4rqcxuvI494
dq7sxZ02GsnWqmISjikR0D4AgLKFYjk3mPGw4rJEBGu4m/A5NRoQhVYfMwxp/UOaCrf99iKUt8bT
b2Bn081g3vNIa9xvPmjJKrHNNlSLl2aigi7ia9Ury8gj02GYhJfEIjK8ttA4gRgLQEABL5dStmrn
BQo8vKV9FM4ChvxS5wI4A2hlW4hMgJjd5uaM7g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="/FA/IZgn8zsfBTrk+Bu5HMfAHStx6+7nTkB93FN2Q74="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
EQJP9shg89hPffLfMgKKX0IAmHyrOE9Yw/SGdxfGaxrebCvYDD5H8kthgp+180enDyzQB8i8cmjI
rCtzu8X18QW2fxZp+weeIhlaU1ZCj0aaj7xAoupJv9+0/3A8fi2KHLyN+MTT9LWMpfm01ALUS0M4
DNh+obOkfUwo0HO/Im6SOm5nLtyWmjgAlJhdEOcK93iIoSeNnk8GZO9DYju9AXoKxhE346P0uxGP
A/LNTQaQa1DLaLllfc2emGGqaP6UeZf+c7oeu9PM6V3FqUgaeVmlgRvqkDdMe8YAOn4FSkIQFugq
CSpAAu1Irc64+8xd7xNItfHMDtb14tv6UxBXnw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="PdtAOO9U7eVUNr6XS8njM1N4xmTOsmifziMm7StdI8k="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10592)
`protect data_block
8yWNy5oZ5opf4v4kS9Y4VeOtXPATyWS7TNHWkt7OnItAp7IrjJTXztB+2qt+fby1b21I1JcIxUQG
95o54VlkbVBXbSiL+UYGnGJwfGkdj7eMzbnZNE8LqQbIMp2UNZ6J5E5O/64AdcSNqL0lnmDsZu6U
qpU4tB+LViwuEb3Ujre9Pj/EOdpMbUqQDYqcuOMUKwz3i67y0SxuZU6r6HdS659yidsq7tJUmlwu
WyGz1GD4c26mL0qt0dz/3z7wXP2QVhhYxFCqaeAs1knLmKJwZoghC7F3TI/6AbXX2Q03LASk8e+B
Nrm5YisThUlTI2u/HTNKvZ4pTyOiHxhi6HJzwtCWX/DIG3vJkWLNWu0BcN2o5BUne8za0OnqOW9u
LI/K3I8Xb7jWKcANRxYoH7AXgyflmBzD6ecceYDQ8m/zIjED6uKPdRe9ht1aINlDXNXVwd/Np68q
RgOpRPcKodrItUA658GhdZ+GKn3BFfbnnvnNcBn/ypZIF8v21VNR1dwPXZ0yYuKMLwP1idbWW195
fi2RmiwWFz8Y8ew9/dmjn48/zGIeY2cQsHokt7FeBe9eDuHiuoMwjHPgc6ak+uk8sxctTBf5oCTE
AlbuoMnHysErTHyptke1O9LlVRnKKLA5xWhVO56wxZYVM/TF3GRPUtGn1D2wCFsroJj8dxeFuG9b
zP2SBWmuGb2iMykM5UJN4ckffymyQFZrLAXahvq3vk+sH8Ht9mwQxnoMZxwYvCnCU6+uZmhYFevb
V1D3KnosOrxhJ66fSvGVhq1IZ5ANoh0M5qxuAzVU+M1DNPFFubWw7fCpf17Tm61JCY3LYV/VMQ4Z
VKOh610CBgo26OfIR4LMgDIhvzBeol8IHsF+N+m61k0O3uwl+Xjdd9X4II5DDFJNZNtEnnrIovDy
6aGDsuBaVDY5BKJeg2GeXb0t+x/zNUpZDrDzOIMHZ/mAMbGjgV4pdpi/qgh7kpjF7QMRVadyFpYO
sYoCUeOLDxnIqM5Cs6QcuUW+m6wYHn/ZwVLtkLAiT5mhzNkHbc67+mhULSEbJAKlDvTuurxSBSdr
yXwE8ZTqGCCaCaagO/psT2JcfqGONWpR8MZWAGtuAgxIC5SONjTeubtyythI9Fekmg3PiDkEWLzt
awlsDfTPWClE8Ep2jEwqWM7H2F+VRPf3Yj0cZK4JFV80wfvcoKkogPSLleXX8TMipcwOgT3m41Jr
V0CkV6LTNqjEFRCKb3xByIix4m95tM6HgMUvQo39DkFu32NELYAFLmqBrCmZilP2FlwkkIiDAejx
vjEdWZ2niOhk7gAd4ises0es961S9FRBJLKMoxo8EgG6+2bbKyiCOlCwqiFRV9TarbQv4Bh6WXox
ST+dkhyUQ1sY5SicsMzFNeCz5G4fLHYtd0glWQ7r+vag27JBZC8q3Tj3kz6EB6tioJwoy7zvTlSJ
71OcfblBDK4gimzmxRD1C/zTLyzTQa3mhPL9zrZRDb+PKHFcLAf4FbUcY2dUlsktMpcH3Rqvx/1s
Irn9RpjHBeRDH+g1xlE9hpm56A6z4PUT2J8kqgoI7GLERIeuPhIaRM33KxrEgffl+fS399xA72uF
E40tK3fE3r/RFTSCn5cMYGHjoXqlQniPWdkJbXA1v5O6bzy5iLeOpCQpFeM995Jo5MFXq/ZwZNj8
b153SgF2oygcoxP1pqooxDiSS+oJTeg+RHeR5IHP81RDvRldcew4n8H+S8I1fqrD1P2bCbHfHrzk
mQSYSi4kTpQLc8CBr4f7woYFiK9v/W7q5X1EFi2umMWoCLTYdxwOlc18YKaM05UcMXR/o0i8ey5T
8kPIs1BLgajqC2CTmuNKBLiyiIlUL+6vy9pb3H0nfAeY5XXzR9JPosTN38VGef+sHquiF6gQLPa2
N4xQl/Uko0XbbOf0bGzmvRu+UtNV4N3vtdZyTjHyq6h8fSTuTxMz3svW0T5NAoz10xnDQReJqC+y
UUXi8I1WSIjRtXa7MYMjjnbkcgtj7Vpw/OrtTiVbEz6FEpOaBR5reyuRcWxH3UrUt3doGFNX/3DK
Zv3IS2VDVlzQPty50+62x5aoJ178T8Njoyfpdce7K14c2kvaEvfIUoirqR7w+RiyinrPuOkqAPlY
+ibUkMEeCehZJzpooi4UyAyK9PEm5ft01rG/azIUwxLorKkn28u/N/iP1AUixM+UOfMGHeseSFx5
GQHpe6jusEU86qltz5EUsnXpud5OsK/2p/+JioHBnkmNo92e7y4+amPwEA0HYv1bscrbdb0KquLK
gD9S3hJBpypTJaCjtM6GvYusvhZ+Z31EQAWCTHKop5obgXxPy9xqOwu2LigvyJJ3BaDRYSHS0Utm
ETIKym+eu/4QYrBYwQpKoCR2QA8RehIL1gPdRQ5jxMCcchsvwMlomvVFgADPEYOXbYj+pWGWojZt
2nhA4dDrWkkGottDcbdbyy7hdGhIGxD8SBp/3UM+V9PxASmHFmroPtSWhvdlF7NbRMd6Rmdf5Jpo
gfDzmX8gnSgqHGFLPKOaC7lCDPk2KC7HIjDfEtbKn9uGHlTopkIreg0j6lOlBwPc7K0uHnzqzcKr
ET10ivH3EC8le8LV5QcFU0+BwA+W8NgvWdo8HzUvo9fbPdnaiqNqPVji0XrhEOp4PRuiImdRiQvi
LfploUlgfcVMCKKPVZ0FfbWYluJGaDmtwoaNpT6hCS4Avxl01UU2kgprmznYwwzZMOUUvTOnKlyd
utvgE+/eoV6iGLT+V1Pw3Jq6JeF3aRG5QADVH/DgvNUac/GyyzgVDkjpFosPR1EEO/IhqncULtOj
nlim/89DDfciuIsTDPM54WViWjejnDTD5wQsjlFB8s6QzpZjKf3zyOy1VJM8JXfBHxj/t7YRY/Ef
u42cwuxThm8Nw4ha0/DLZMsl4X/xpgRvXZbH2WWNFVNHgXWUKeLPF/I0lHhaxtdbgvMaJLbXgmpx
2+eEvQZ4PdFOvtID2R7gMj6wVLhUiqGzb3nFYXvc/OVBgFMi6grW9ehoXDtp4W0aEaKBh5evCS/y
oT45txjgXZ68L0JUZZQhYc+ToRsobXTI9LGUdYRSzbCt5TULgxY4uhAwHKurzDmIuycAoSqf8f2g
3qrm1X9K2GK4+n2TTekV2JvRPh/ThDZJWo1+B47dhZGwgB6l97Ft7F/8zoOvAFDoDk6TTCRzk9iC
sz/fpOsj4jm3sn0kQvL9VfhagP79KsRNA1mv2TjzPlu7/tI0RPldWuXY8gv+RALOVJiGLUjeyic1
8O2m9pkkDc+vU/hIXepmG7jWd9V5JwUNS2E4U94XZh9m8r0AEP2UWVKJvdr2x8lGH/NrDtK44WbA
Nbuqjr2v8rOlla+JFK4WNXQ2EEWqFbhoNSa51iHm34dgK6uJAAEVvcHLBBajA6rJ29jqODxNOvAu
FBqrwmLrgoU/ga0FAyDUrDV1oNU1lL4UaPJHB/igwwlEMW1dfrR5IZiSLrEvP8nV5a/GXqVOeCIR
KIgcmb0oVvKsuSVe5UEaSJmqlZfGw6gGmWSrZsD7ix06A/VCr54yCj6vWxJBY5PT3fwJROiXP5VW
fu7fY+WNE+atZu/QAxPs2gx2BFnIByd4opGYTtkHHCc9LMxa1DXemMkVIPSMsjOkLI+vXFZ8sWND
Oi7g2wd7RHltJ9JeEJ5iROwRhF0J5hsPGClcjNIR9wXV0+NAc7AusMjRTTAf9ecJgVQ2WR1bR8zi
zTBYBNcVaFDE3OkAx9KDorPo69njA5jJyDDGb3+b4Alb1oB/8FuV7f0E5BON03iosteTDE1hNVbP
/T3k1b4EIKFodzZHs1Y3kjtlD6PjOez8YwkBdIF2jfUmD/os/CVT/vj15sOO3TvWM4xkwRxU08Nf
Q61OGpoRoCoVZpcys4onNMjXyy+rCFmqqxnSAQ+8PpYtx+MefOsl0T9kNfMlnWfqHaqweybTimpN
bzHwdwjVrhopoMjzJFAHH801gUK4TAn+NqBTBftaak0jh7N+R5iCgvrO0gNcHrlLirhaLXLfqlEQ
iFv1zpaVjlIfLd6n53qz1eGhaXTID6vS+O61sU64aZI23rjXnCad4rvEPW4OuWp2DOnrF9XMXu7w
5vqR8UC7hBOv3l6CpVPx5ndmj2D+6/H1pFdWNbEj3gZ1+MBDNiUeZbgfXFgTECW7mgTPbByTNE+l
0EzhbYIRTumwJPiT9p2DArxZIeSr3erp7nSWgnWLT7Q/d4GFGxmB49pZC+IcKs/PxCnR8Jhx+bcG
1enzD536Y7GI/DRJSH/UkFH0KSWlhPUXroK/ly+jfUv8SGqz1gjtOJS5UPO28On7v28IqWTQCLvq
Hgp439FKQExidBsBsUToROzczhrUlPTfWFnzkGwyX8TOaOtk1cPDLYXPrQat56jilvOggC6oTVzY
kCyaHQ22hTiZs8Fcxt0esAP6UDSXl7Z8jkg3ELKDiz3UHt/4v5rKP9VzEC3Q9VoxtIXcneKajhZF
sRvdrt6YkLKDuaUFq29ESSYm8256RiEpBRHQ6A2Sh8fzQJps4HETnfctnZooIPA5szI/MZpOLRRH
obtVR3Fta2tjE8+wttVjftG0yNZsvGT+MGbemu0uCwZAZqAGo9CYnqjOh/cYjgWSMtFm9ErYJhy1
t6jXTMI6lVSm0RttfrGQyUC1LqfuGhjCo4lj+EI/gFjPZbqp26l5gxEHJj7p3crvNy3WFJsOJsH3
bOJzBlli3G8djZ5veHJ336pUaZvW4v9zeB4UrwQhKW5bBjVCcwIVQ7xk46n7NwJ5PC6a1g+S3+Lp
eJeNOZYOpVXbWHXioj1+1IBKOO+XkhWDW0dCWHw80GS5vk49f0TePNXIyJ7QpXFPfDGDh5ZmgvrH
5QejNduCfFcIA87NCDK6cOw6eqe5zdEYC/So7gcXAFL7lIX+qV38ETh4bi0Pa9jdufjWyKiYGtkt
q9aSOF2zwdR67uCffkeq16HMMS7vIH3BicSUdDTxvNurRiVK1kZ3kKSy4HKhI1QHeIGxxztzuho4
gt9QQwm02SUqHj2mLrsAAQXnHmhr3zZo6DxLksogDnBLeU3COJqQppR2dtfonUvRpPUIdNv8TP2h
QiPG5xpqWoGI3VnPNFsrYbdj1fTuw9f8VZRqSMd5qoNQCxuHvGKP792rKfFTVXD7DulBjUgdBROi
2RC8q4YJpPhXV2TtF9Z1Y67RT4upSSslPJno8wfF7xlPS0qhzuYfHrZiWuNP4v6OpBdgY7F90LWP
Oj83/DFBQ8nWn41xdAnFKCWfxxkG1CjtwGcmsWJXBEJufYUFsiWImM792ZNWvPOXnfbyVaA+IRdX
mLXTLWig1iSXHpaU23b3tRemkC5tkL5GmU07L+2CxLb3F9Zn0Ci0J5rqOPeyfa1VC4LIiinJ0Ic2
2d0/5NX4wZfXf4I5bFqk940jEOmqNCEVwBE0OSlXwb3WtEUOemXFa0TpiWLLGiEbfgCjWCx47II9
AD9+sVaRNLgJ1wj5NWBt9NNCPeLpWePF4rp2wty36DdEQzQLWSkX4vR+ZifQzCMr/19jpZB0v/kd
REKreBPptP15qg3KWuQYKfKXFaKONMHkeZ1FgJl6thZsmhuW/ZEGAQ6KzbY2A6h+tldy27YH2pe+
/MWng5wWp6R6z2cBMWAu5khoV1KT2PK2bY5CvcvF5YflJMm4Am/J6WIsZQ0czI1RJklCqJuzbLEH
/6+w4dC+Sisgx6LhK2aYJAPZIuXalmY/eCXuZK45f37s5NMBIqIpVKK1TsOky6cLCtxkRn4pU3Tv
+GFS7tMTmhqixzCkR4Nrefxn+EL5ncTn6mgUxUVAN9nWxLJ4Uv3DUWNrV4OLd2ZIrNW1eKhPDPCg
lvICQQU0mgUjsq45wAq3rrGmZbGApLmigAe3nHUTmZONKtv5KVm2bN06a7oM7OkMN2l8uExPAzuu
cF16MNl10hbL1t0pynv/ALVUTjRCJgN3TjRuOXV9vwGd1v5XNragYivybkntaxQvJnCRQFpD/YX5
6NGcluFtqjj0mup+qBVGqPytmdN7SFp428VovMppEU2myYUp1yDBDpL+aeVAKu1K+uXD110ExsQt
1uHuuFN84shSGrPkx0vZD8yojB5T/uLHEqEcrEBZById0Y2/3N4Sxpg6s6KW7vFdXB6Z32tsQI44
B6NXCSCyP+pcos5em53kbw4PCvWUwYOAy37Ao0x/TWOqL05ibt16x9qEndA7LlcPzR51AvoSww+I
3AqNc2lJMNbqw8g+0HFy16dqlQ4H5oWcs7KukVXlFlEM7oaIzVK/xE9ZoBqhQY9UAODveHp7GoJ5
+RjbGadH7DOx3ua559CYEayVjcoiAN36KpoLylpKBDcH6hADSeDDpdiP7U8ATuPttebJB8gv0xHx
xRIlubaq8I2Jm9VpNpefoEasQE6RX5+BchpKPUE0KMgL74+6Kzmjo6vSqI6xFBPzNIh7nXE+G8K+
xL956j7XSpRIc3TbAluKwkniazWDwlQPzPcqyl0apPOSITAcBs6Qcr9IaEF3VpsT2uLl7wOoYzha
g0PxjBORrax6ENWvDQLK/yi65wKDVi7jl/85bF161QMazddB5kIIe3zX2r8kL4+lWaeShyazzGY0
n1IZ2D0rq1Dl5EW4aSdDnXmD4eTTuz71yB9gPAKHudFhwefuwTz9otJ0HNLTJ9dmtcNTSc03366i
hQQOLma507+PIlSWDf/v6WZFiGLC0iYwetsoIgq/9e/z4a8joLterVZkl7ToDgibeu4paXOJVwsW
bjAeeTXSRSvxBVGFkyEAJo76zf+xuZqjgJqNRM6vKCPa92+6rRVnlkluvBnvauROq7xfhFFYbbqF
StRKAbOKohzlcPAe6IPN10T+2zcgvwui+4QNC/4RUv5ROgb3gWE2QVvW7XXPh/4246mj5v+BflPi
si9ox9l2C8k9dN2Elq9FTg3juY+u2Sux2r8o/xHSNuGJYMLBVkptnDAhByqu6ogJeLIxo/0uJJYH
5BHXi1fWMESiFqIsGw3vY9yNnSulZ8VqrWgN9HivrZkCKtSFnKUEk6kJsWP9nFxY3gquHpMlBtdd
lTis5aiZrjxRjBG128emrOgmLQ9Yq6jO3yk0XojUq8rAfw87EGjM+m9DLiFC3Xn5B6zh11NLFT6M
2GOOXY7HiRnBPxgPBQGrhxHs5zwooLXJ0J39MJwXGzpEBVfcbz3gwrRc5knY02PfTc1to2nfE4Ag
HOVi3wWuymFZJFUWOp9nrVzJn4qjRRNR7aMnWXR6tWc9eheMvTslRvbfdXTCZqrI8pom2Dl9Feor
Oqq8bs6FhqFn72yvDl3wgvvdnobriTkwT2SUIxx8+XE2V4lhAUhmNr7Avl1EbHGvOpjBD4g2XZqU
JneghoEixEEIypYPa0tzgLSDZhpkOM8Y+E1KrQDDofRJMyCSOldCy66XiWtn9sKowCEXAD9yNPto
hWjP2ngd9hFYJX1dwUCmLZz7GVsLAoAo45Gm6mws6e6p8HunniNBfObRxsDBuJBo5PFzvXe9mIaA
IqrLsSYJNQsKRROFy1MN+9kMfbkB+JdCMHGZLwGFJfXsEZLLJIUIqtrzQR+JF25oIZclgh9mj+R2
08HRXQiozmM4W9oXjNGMAMzN95pRC70y+G3KqNkThRxpr2RrSW1/Pw5cZR9CQn7nJ20+P6jFYyg4
n77qSjpi+s/8GHhyat6yqhU3qMQstUfN+SnPZjGQLC0XivkkTDdb8sP+F/f0XA5kF+JyhmO8rTHl
DVNmtVwx69+9JUd7rVkLSx1rVmGLwJ2nYnvMtvMtRna/VfewEx8sHTrPu7St7lg9Rl3JNXFiz4ou
hKGy3xJlKyIIc6sjQ4IHygnTNOtkHel8BgrnnS0ebYTGXkUnzZHldrHRCySxabSYFoYlkECb90Jy
CFlK3SPcBdrXkfK3A/l8lcEEmYgGJBwGw89YPPdby82bLXOINQUqmqIOTY2s/jQREr0FzY4eCXmC
Ii1yqt+5nKNL842tmIo/vMzADO4kZ6h4afsIons17omKS8JfkeIrgcxYZqyj8yASyDfNky+3yDQV
JZUwr2asPyYObr9EH82TWM5igZJa21dGybRXAkeoAizlcinDK3dT9ZjeYxslUhMk8Y4IploFXnj/
jcyr6HRvWBJxLR2MD4gzVi22OztuQ+Gr7sCSqSc3j4VH22sEvGwC12b09T/C1hBlgSblr1UNtKwY
ld8LrA5rKN3K3ic8PkyiDU/AqEwsQdXURqde6+hGZ7/lhcN8oJ63JMw8t8aMkFPld0pZVynAW1Ne
3ZM02Hld2uaGNFp5ieI2Zi+mAkIijS1OUihzJlxQswz7ropzs40ODz8VkrKa7/UDQLbmigewrQN4
FpL4g4i3ULcQOkssDBzInwx9GGxIc/s9kmcsH78iqBpNE1yw9YgYQi8clF2b8ISpHWoETmzIUHXl
PO/2rAnT2s0VtgSNzubSTDStz+tukYpyjxBE78+hAUOmBQzuIWPHfSmFNJUmvKXm4Nw+ZvI7gcO3
iJDXbI0iRlwt7mi/KaehD+auNbxvO8oymc7hmPmluH3G0CCiVoWeleIk6P4Gvwx51ZzY4plaAADU
oGUm3PKty0k8wm8x9QzPDGkqDchXfyJXYXEjnDrZig89FecqmWSeV0XkTR+38E+RquJMV0pbBVW4
9WcbKh3Y4N6pTKm96M1n2o8tP3CiCtDQIPKr+p/PCP4nI7hOM/AdU439MJEz8aHWH8nTTjQkdpY8
I0K6WfAPq07kpEkr+Bbs8bX0CSRwpNvGpaWSsx8Ns3JEr1RIG3syjAfKd04ikTWM1nrZHF7HKeO+
RUX2CQg1UvASvf33C0fK5I3NGPQVt+zptTGIEp8Qqut0jUtw23lbJet93e5JlE1zqyNk3/y/dkCx
UpCfaH3bWvAp4POTNlSeNZvZxweHKbU7sR6R+N6D4sG4CmrP0TVtD4/mVNlwXgUrPesicpr+NSNJ
9PwM0YfqDX1nhs71pbJzyeoVDF6SSM52rREQKzLHnE0lfU669b/0N7GfkWgTzUdyD07vAFrzHWX0
BZ+2ylOqdTyUbH9rOUk0Vb4LlR3ceY6oVFowNu03oILsLP9H+ivz60sSxNSKzQV2oj4zIw4ToPzE
Lp3Lmg0aUOjZGoDeZps7tE38+ZkfI0pRZvQlALiVzPEOdJiXLNqBNEXBDssqnvY5B8IErF9XELFe
o2IGPlso6CV59tFV9W5fRCmkzlN3JePsCjmH3jd3gSXYA6Mklqk7+PcLKAewZvbA5/9CkHF00cvF
qU4z6571fSnacaSpTkyaaunR+xZ8C7vlamAKJWXnKhH1w+83He7dkUf6DuVModw1Xa1N6kyt/Cdc
vje4/Tb95Ot63GpnBLSFfwkv0kPZNuMARN/SByJk5Pb4R5hgkMnmTF6ouMadHGwv8T2qKeyZR+uX
FH78fz50g++ttzlVQSNHUo2l0xeVe2DSb9MBfe9oIKxsgHObJGf3LLa6Pcdpibg0+rSH57MHY8zo
KH3xjMVZL8njtYr2rt8QaDnurVbXSuoyv+FS+spwsBRmV2s3jBpNZK0W+g8YB38dOe3yXTr2I3i1
Ai5BZ9jF0muG82AjSFbTDNldWGv8EB+X6wKmt6SguUKzwSZ/hhXHeg8IGM43KzGGHjoHWsBp+zQy
QR3JGZ1Ii6povQDS9fMvwT7CZz5dNTUs/WyryabCyPtDO9Z4XEsxNo8M8QstzxUCp83ju6WYGnOi
Z/AH/C5oZK22xYrN9f85WQHH+F6zPvvvsFkVjESJldw7b7yOO1f6omddFXTGFbRPWlUAhfeukzSk
LZ5zhZn+m9Fz5631nHb3TnOFe1MaZLF3aqqANbbBdYQFOFZE3KbWQvyyxKWjP3PxmOXdsx5igG+X
PeeuJxOGvH+KhHlUyYXvv/+1WcvRXBCtIwJCUEj+U2qs/IVgppZBnbEHoZxw/sr1pq7Cck1G0XhC
jsnC0wXLgjzMuZ90s9sP+vPS6TKFD2aDFmvvTVvIhL3Ag8EvjYqw9jhg5jGksIl+QVnEAgzvsaU5
uauJ/uXBpTq9rR/alxQoN/EQxFCSfpUV87x2k1GK2HBRMnjrjmY2MiRsV4XAIag8enPkfHFO2OdN
r8ZIpg3EzfHlG2aFxfHh3twoG0DUIst0vf9r+kQh22ZlogcHXLaHHKRX6wTdjDAljf1Ru3lqThUR
XBqDbk5/bnLbGmQq4bqIlf7KtSDNk7TmbDkbvMrbe/BKFyGJGVf24qCx4uV73qFsELStB0KcbW8i
hN+dM9FmtD8l8jsgpaMgIHsTF2V7ovN76XEK3t71kN5JS4WSzGLsYgG5blWrp/8069oMfr2R8GkR
ZKgmnKVdDgJ+5VYZk3Y/izErwCn03TYAeaPSu6UcnaiHLrcgccyH6NtHXg/SY51UnjhCQqN3FJOK
42TNU1Xrm2RQIst8+uKznnGD6cn4b5Hu0o7TBs+s8XHx1LlUUwd849+Zophxvk8bHvXJ4kFf9tkc
Pkc+lg1dlfgJbah60+T9/ufR5Gnvos4rqAYMle/J+fROFFt2t/gW7JMg2Aiop+0IyfkVIY3HWBvH
UEHLSytUOuPfitsmUMp7f5iEawMdRanFJkXenwU2145M76hBVcWgLm2Uq0AZAStTPQt7Vfq2Zfzv
v2XfNdqJqxw8uQtZ5VFjSyQ55e9C2yoqjyiep0ly5rxcffKOTm8yYCW4yGUt0HYwp1okOiB84nQ3
DL6641pM070rZXP/9AWBKx0jceSqYSjA5JzN9qOtefa5eG6TY1aQIewRplTIotN/IQP6fd1CysQP
fFMjqwu29Qz98kI/r/4mO6N/bFBhtW2XJ5wYxXjHJgot5VkD4YUNE5AmACzzxZZ6ZzzwV1Twd9XV
MTobLHOXrIIzUqyXx++z3g8cczEbXNOIQsFzWGtl4pKxwkv6T9KF1VOgPdvV/o1b21EshwbnN8Dq
kTJ2wvUxAVhBGAu87LHv/SZtIIgidBFLuUC6FizcaHTTgZ25l84TjYtFnXvFbfjdzU27z475QBww
q9NtW/h8rUpxUFSgKtsHJsebeqe6uO5ZbzJvQTt1NTUISKlUgVByvOSEmhD5QIDWZZ6mekg1Nta0
3Gbs+e0GgKwDrSZmxwjVWdyQ7Ez8hctFCQxjI+S3G53+3cR1J6+kkkmkA1/tVmo47RTQh7ISR22L
ClBsWrPe3dLoqM6EJ0a276X4qhg3w6UwA6+LdUptDG5mQj0ls55gzursMB612kEm61iqY5UR0+km
uCWf5nXFdWPtitTGTMT/A6PD4V3MrY2NjfPdbFiJxKPhEiNVKFpZJoWenCQjv/SPoHBnmAexsYYi
TOdnnR4QZKl7gHF6ZNprkHmh6h0jIjmZOEu+lGQOd6/zRltUQx2wLvor4okh1EHezwi6ptaJ9ET+
DscSHgbELkLys56HvmkoOgkibKqSZjDwhnT4tIgrGm8sd2NowMi+NL0QWBrh6EL1rKMpZNdf5tfD
6xsMOstok1ZaAmxOQLA+cTfqClaxGitVLOSbK365EVFOgBEw8VOsM/r52aJdRVnW4LjNOqGUFSyy
rmi6xvXESRmvHNo1v+MOd9GpHK9YvbUigSdEyqD5SPM566tDtjGAhyiL4j7HM7euKGjTQWYoDOWM
3W9ODsYrfap9DrBebgaawDp9iJrY2sDjEqCvQaIC5stidecyBYOgG0xuXMQlDdT8ZwN1BurvNR8f
AZMQo6RYTKIKAQHAzAzzEER5oYJIixNxy+DmsuBpD37erxd1oNBKHqgMHcuTyT8hdU0idhTs4PkA
toKqGmmvNoLIBzccWr4hI5C6rcYmUcPAhSDSi7/G6vEMoisUbDAXqZA2VCju9V6ioHpUyMH24J2p
MHW/g/iO7r+ipvoFGGg+ZILmTTggufyF9D/qbkZNNQrmSFCJtMei45+uC0nsbh4j98phqyFer1Kp
8tBw49vLTCLOWPcth9JKdAGPMGVDA5AxSYHWYjKn24zsBiztEuJIUXDybEJPrRk+dJAcIze7irxh
fcfB+/m2BYtERyWRELxhVCvoaiHs6FvrC9YBhIB2OK04MQtBt9CDRDrg25hSCCvQy6DVi08CD5bo
/PoZR/zAHYXpthHyNfoBbaCm7eW3OH6dOBIq/7Zbj3xRVEBvF0Nzf/bFq0N1YQMgFz/WYIknh39H
yxfDIHMaaW3rBN6luwwrfZ+vW3Lalx4xw2kRYJEqQnRgQ2no0P8YdxGCC6trZAseUXrC2io95EtB
s+2uHDq3/7da0cDtsSqrVeDX8DXcobaVItS4Emqxoyk3e17/vMciH/Ahrw71fsOTUdeMfYGTJ0Qe
VWWxjLOZlymadVLxLZvYsIHE4hMD+0zx5/axbghGnNfcOV+BqOo8MRsGQQHJj9O+YS8GPlNIGS60
4KB5lWleRIC2adtWw+cTLQ1JV5zpLnX4xnGwZUgpmmvLzToHUksIaQwofL0EhCNE/aH30flDtjR2
c91eII3hufb0vY8Dh9HQARMNFdEubjCRkVaQuojJInS3RCUAEQ3vjpOAA7oeDVUtYXB5GPl5oDPC
/+C+ca3HI4YTxXBpdccYrWDI5qAj5Hb+B9HjAnYSCP5dYiL0YEH2cZeI/3WLKjt0fHCx7A+ty+H0
SnUey/XUPjW2SW8xTr0evST9qmGanm0FXTQv4GuxUhZGgIuoCnh8CXQWP3q15pLNMwXVH7DUpGnT
dirCbWwa6jCt67VSTBdTxPnNZ3K+8LXk6xT+vlHrfGVlx0Wa4wFCKVSnYIwSMyVPDGWCjxjQWy/7
giG9ebupfXa87eBq6d1/UpY31sg+suz3ZYI4IzwVZEHYSrConiaZBDGFq18prNpCEI6INI/dCoCu
XyUuOpfaEencRSx12TsZH54uIR48+j2oKZCVfakHKe2zyOXwRsLKHwP8E5kJdDTBrdpM6eVFOD+a
NZF+g70R6o5sj+GmyS0Qqc5ev7gsb8WSO5bvCWDQ85a+MFAXHz88QFaTK68FXHE/xw5SSEwLzlSl
YwGiBDRbVe4ioGtnNsKLCGGR8TOBpswP+fgrbwPlc1vzp14R9ly7T+KtJ6+GnQEQI28NEf23vNB2
OvBltgpDE9LQvhFraEvku4JgxhU9w9o47xK20D6C6u0y7g3zhuuV5l+2E2BwfePI21dU46K1bS0c
9MODrVfWjEBXaXqtWvmQHxmFss5K1ASdo04DWTHvcDCIOd6Z4Ogbqxk04qxLEMZqFIJApYYd7foz
QJ2PPbcjAdxkZhonNEa/COzJRs7E7UM/qdx8I9z3xFww4DBsI2f7itIeIdf4ObDpQrcOW6S9S5xg
a8pylTEmefXMU671Biya+5/pdzwExgRS0IDPXpivRWL3hPfThFUStuQZX0aiPZ9qe38vlYMkHtVP
TKOeyfjQXwtSte7X5IUjHzjDHtA1nw36rmRJMtQV4kR9biLDPRqVsZVVFvjLD9JcnvULXhOhAzJk
jQt83wFtU+TsWkJ9T/jZOgwqme6lATBUWekEL9mJCBTa49EsAIUCJ/OAqvBZEhg6bfE0Vg2HM9Jx
31UUHO83UOcPM205J+hKAwDOZDNkaV9ELKuV8nxtkz6nkzJPKftWdaivV34hYqpNnas+2E9gXyRQ
+Zc1UUs8veNaAzHb2SOWP6izRTSf5j4Tl1drAB0Mpgw5ak7aT7XS5t08ZPI/vskhOJKXRhrxkIJg
KzL0rUNpy7/m2MZUmTeSxohBUKt0hV0WEjrjachyM7yT6Yje2sXaxUEY7toDSnkcjqCxD6Y8P46S
8mKHXazs2LxBVfJZBMz3Uu2d2D5KklnXZufuCqcJndMLV6w+h1vJyq8bU21Frr4IQDMG02zgTIdf
qzA0Jr2Xtc7bcf2Djl4+Gwjbi/YmBrli/ffkJz+OJ5PzjKokGxueRQks4BUK7QtWv7L10gcKsi/D
22wm3kWr7wWYRvA3QCyXqyOseBm2l2ppScHWGx3Ab5cstrDPz3pCG9geuu342JIVRplnY8LHQlNk
3ptpUlicvQbGhiYWrzHz/gPnmCf98VTGiZbyYQqaazlCzW8AcV9VUftTX4Va2ijb1SIipOb2AU5n
O/Ku/LxaE3qhbr1Etewcm/tH+xEjF63XxhbeGlY46j6YUwZqRw6T09BZ8WRK6lM=
`protect end_protected
