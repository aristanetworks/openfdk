--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Y1TaWFZ4JlI1GxmSMMKSILTp41TrzDB+cT1609KDOfja3X8bFZuZSzYuWWHQiRLTVj4ITx/SVh+Q
O0Hv4YOREbZAalm8ETecQp+pwy5n+b0kh9a0rx8SMRf+T28d6N9wG6NGkTreBA6zfIJ95/yPZlxI
WjbR8DMvqq0xkBKquVhakjAbLVsTXkYB3xv/FA9r/OCv1COjnS0cGFEQBT2MVSx8Lf90KNfetQ4n
Vux9F3VGK1mFpfCjLcOE3tT0tBRpRD7NrhAfdLKXV9QjyyP8eWYAUYUOV77RinGwDbH6ixiADZ2R
uuo+NjDSRUUWlsIeHKg15+1In4amBP6hWTfupA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="4MunXS8Ve+24mYpiL8Kt9p62cc3wNqmWXRzx2pimE7c="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
NORRe5NLCaARuZGu1t/R7BlOfJVtZsU+EK92wpJfGh6P0hXxi9nFF6z0PckvPZbG0xOSVSiPEINz
ZkdLj4lzgXGMMneGwpNjPErlSHHUaz2GUWA6AjYClZzf0SWQLc5ACXiZGtiSb8lxB9878l9TRvvG
l48V3IbCh+5FdBxEU8WPdv5bl0qEJ32WtvWrt3ahVks7ppRUeKEcQNRolFisCcuYhnmKHTOZ3LVc
QOLZeII/qTjCZiqRJuCnUunOW9pAQ4oA94XtqHcbK4gtwHpc46gU2jKQ7e/gSoLsK3yeczgkSJMm
X/poAAGarnZr/dZR8Br7xuodIWNSTPV5ApUfng==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="y0d0Wi8N6o9VRxtWJNNW/lcUH/wwVAIdkue/jI6Kpls="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4496)
`protect data_block
41dwzy5DSxMV0mqt2Qsw0Zp5HzCDEG9HRIWNMF9tULbh4lh2MVHGEdNwBLVe+XiQgvuwVE7tDbgH
bfrR44vHD6oRYM+dfg8JFrq8yjy/xcJHYjMIl/2l/EHfIPFzoqF54PJV+3bmKSZx62acDrN7KQCv
crP2m/+ah/VyNFgFI/EsXdLrh2Z1XEul1T7KPqV1X6Vm8uCO69s3T+WgSDTSymKenzELrINDFMwi
D6v/3Ofx5BoUTyNIRBkwsl1KJFSNMfDBX8uRnJY48hhQpm+wLSa8Yf2m/iQMYQ8sLU316npQ40qL
8sioS+dSaMPVpBlrFUO/yllKOrSZYEXrZ94iK9ofcrz0VqD7Z9b49USCV7QbppwYDd52i5CqBoUm
mhdYnfXriW8B4wi6os7fwyzi/woG7avjWmsM+ImBTpvuBPDAsSMsloRwhnKKwufVjK3LsZ3AqoP9
dmO65KDjPEmcx7VhhB54ov/Nf6x+KTeFsKzqzLmUtE3+Q6dvKNtlgRnVCEvLiOQ2p4eS4/W3S4rD
epHiFELjJvMhFkG3k2TldiRFJOjleV8f+s20vTFtmoXKvHQ1qZa4vIBAe0oBa4FTmHai0p8tiu0f
HXQfEA57EwdjncZ+96N2QezTqcQOprCxuzJBxaGdDkKqBRg03drOC4EFEUHoUEKBlhWCjFfPlkj0
5ErtHR5o0rlcQ0xeRUA2j3qsdiWWjK1VNc4admBc5sRigNusZAageAaiTRl1RjqRlwJ9zMeAtvcM
jD00XPhvA5Oc0OkJ2bH22OyJVr3MGR2C6JVtzWlUa+ttZzVHTIk8R6LcSsK5W0sfmfuJOP5i8Oxy
9EHvjqrwtr7wuIgF27HDB5MiulU/toxtPzaJPF6Z+GnnlvWoZ0WcykN2IDFWXD+1QU/X+wbKOCyE
Bzb73Pp89uC0LKZVl66G2kVptS36TakMkAtXPp2/lZCtjbbab/x/nB50HUpz9Ls/h9ULo9xWyTcy
f/59Q46QxEFgSCL6AZpk03meolM1tVFjK+9eyIfAiAA0CtshsmOYKKI08HK1d74Q3Yh3cMTFE4NX
Z68fBY+r7Mk2UfR8LjWAUuNS3OPCuNATcIMg7z8prwuEsbb81W6KjnB8LD8kJLrG7gunWzdjBWpE
FNSsHri+S+DXYE8KKypzMI4LRpOsnh3PxLqu/2pLaufQL5XzDj2tx2UmaH8zRy+5SBx6CV+VjlAJ
IXEuf7NYHkcYGbxq9CvpnQw+qz2GmxJB1BBGhox1cpwUjBN4WnYLA+GvZ9sHNynLC2NdspTVSlbl
dVVLBgdufYOAsXNXAnR30lL4tCa9F2n+11Qgy2DTBYNLoex26Ua2jMARbbzS/OrGZjL4xkIirlX0
S5LqJ12VIoHAzoVTDyFdzZRdDzx+1309QXElMhdJtBHx+4zuWZ3StjZ+JatdcPuGBPIqGm6cCWYW
KwtoSqOcZXqrIWS60zVQg8Bz4j4JRis+bNe3g0LB6bTSluHYqzyxe/qPLZUF3yG4dvaj/NT03K0s
kIvhYIjXHY0QqKZRe36iHISslYHwjqS4iwWIFh2M1RG7yQ266YeAheGcgqVOwaPVp2Lr1PY/1ESA
l7TrRt6WlRyIv7zFS2QXzH9zcSj34tjFhI380sHRzZqo1JJMDf0WF9e/2slsg4bebJC/nPIJzSLp
mT/Fo8+/+i8NWTIiSYhALYSXUnEYnxJKvtUd4hdb70bXP0S7saAuiTTwLZjI5e8+fhvhLYSENV8C
wdee7zQfB9QJT1ow4CUEmbk7TIr2SbeBU6t1k9iezROtQlYPO8v+qPOQ+c9GkmM+BYjwsjKNNaSn
y6oIZdG9+i14h4lGNX6seq9GVZ6XQAPay9wbbNqq0kTWZg0WzKsfoPEI/1b2cAmuAHETKlKTpEi8
EOdnrPtbHK8hOCQ11wJIknkCIyY67TTXiH/6QgDvxxitdt3sVD1RvOEi2vSM/Ef382kco/pvjzup
pz/xlofhmBphF/H8SpK8/8mzBHKrmwOq8EbI7IVsvJ+SqTJ/BUniqykY5mAtvZBCYvr6RzMuwfos
Djloz93o65YSAKaydfzonlb4nvpxi3jR29pX2dhAHmHQL0OyAYyUGWS6tFLYDug+MhuLopegRwKf
nwgvOjol35wg9M+d0wikse777MwMljV/JPAaVlubdE9h7TDNmfrxvboJXIbm7KduRPh3rlOI82PO
yKu/D608I4acwmmceX7nLLdBRlALf3RRIrPV4Ao79dBcS0h5Ta5EtUWDEyJiRAy6D5FdVOuAU49c
BR8qy4PH0GmHAgzAfsDXN13wYyJCyBqc2LXBEZ1RipOw7eO2pCbB//LA1aIzwGnwEae+8N6UIF8q
57foG8G84lOj90q8SW1BSQQnXjX+DXXD9/s/GL0dLXU5Im5Gt/WhASWJAizl50ykFzIrBRw3q15A
VLVpcxFj/H+EMBQ4H6uirgL7jW+Ba8TOrdNgWqNtJk3zNUIY9bkqelubkFCoZUmn+muU0MVh1A57
Ov7NqH+tr2Lc2RlPKX5FV06/MHhvM8zJjI0Ks5cMCsEnFpj09nBhXvo47+9URmj9bHoOB1qn/lT4
ITQ9ItbUdck1CZSdN1sJ3BeBYpMWSIYmYxdHHL0q2XjKep0tKXkQZ4PWEQUJnPifM+AqaW76BmNR
hiJSuKvBk72aAEAZb1Pvj+lfNV38lHS7/ZiUkhLiNthIV1U3rofYLmIRnA9FurtjsEaMWWUaFx1L
hogCe0cBfNXY4Xqc1i5Eic140nKTJmm84t8b62QntJC8CvYxkatFRYnF6as3Wny1S5AvNalaggc8
xzc4za25/unsUJWfAZyoyx0nU3qIMqDK5XYFnIA5OdyUY3Zd+Gm9FKoN7UvirhAjCycYxZvxDgbM
S4fCM9sTCBkd7cqKJCw11QBJF3Z7ojbJbYQZ2iZNrHFw9FiMrCcXaVrYfGMseeSGn4Ge/+W0u8Xh
SlVwVXy4WPby/JrzfRax9btjCu2ou3K82CLgM/7oAMj45pPrEroLFdcnB1+zLHHMmnRq+qGt48bY
m802Cv4ev4w1QZUZ7zW5Dj+XdXyWYVEMu8w0IEyHI0sfdRsJ8q7z+9W+U5IVCH1S2Urgj9QuwCfv
W08VsaBsmotTeMfoy7t54X9r12mD7P1VpjTSmmfFd1GzQXMinAa4rDh+VogAMEO8oQJK2wWf+05J
OfIkGOjh+QTvNSOyDUqB42m1Yg/z2fNxxFoBIC7CCRhAM/JMx6wYCZyzp/LTWF0sYIWDKWNocZ6u
tL6Q7xwcyGj9gI+3SzF4u/rflzunVx7cziEuc7ELLc2v9lkne3As/KzwT+aqggHPdsEK/CkN1gMr
OwFr+54l/SZlEc43zKWlKMZ2Y0vmo3XZQRD3GPvuGTuH1487LKb8BD/4woqesRvR81b3Oj6td/69
QCyz0ULUzHUKTp4BS0XdzJdQ0467bhtHXOR0ngVZIizrvfDv+Fhf3J8nvp9rr1l2ZK3iD+P6b9qV
tJ43AWcwtt2gkGdY8QkxstOTvbX4VXUv/d4yFm/SSeVMn3FCo3MxmZ1udnDkVlbvf+cgaCJwGMtB
CQvXOHcnqq7ot+cmmUXeG/jVyOPijXK5jwppAqhqIxoqgyNoCaPZGZVHsNIOXVEfeG+nX6ImfTbw
eeWHMuzYyCBOlvdNb38elgNNhBWytwgzlQzQoaUhlxGHLkeubgI42hROcpIWj5axsf1OUkB8aBUY
zG4+ktqmlcLRlpVWvtcY2LzdiszNBUKxPgNC9cIzF7NpM4tuFNB6uFDiZsXftMhovYzJszjWS710
KyYfMJJhYEtcSIx7v5amgL+z2G7ToUgn88Yhc9L+t4tZtQJKxVs01Bid+ManldKBARVPhFfzGdBG
xFXkfwvga/hNlfvjhDKE8JBTw35HGjekmQplovVtpX6DTWCw3xTnY0MhlCw9p+b9VrLyXfhoUPJ7
lLPP/wKpSkayKi/qf7PtRi04y2EdW//yA9VMgIC3w/EaNEvyOEJ70Wsq4kaZ8Q6xhOlMc+TWwWEh
5+eX4yFwTW+xPrMKoP68vner5TYX0PhUsBP/pIsMa/I+tuGpk6L+036YpCA0rSLn1aT+AHFLGrTV
XILlkS8QhyaYw0lPtaXTyHKFbSdQeT7mwaStYBgr9PpCSRz5oeCtYC7zHzSN0dXSD/6Ybm3iwZ+y
/83tP0ksU2n80AOYeLFE6a8ycuj0EmYMRJZKQOuWy0LVeCw8gWlWF+/+8IeRppCcNsfH/Y1eptjX
yWHpgCWsdjY656hJ50ml/ScnKRC/BdvaHwcyjvn/QL7W9JnbDOo7GHmOZEFXDtg+wKy6VAjubT/z
fyX0OOmWHtsmI9FxY+yKXEQ+l76+2pCU157wE4tBk8rttDriia6PFqoio5l08+dRJKbuyTJA41qn
IhvyqSv4BWXjHpB7JV5GIvceRBPYo075D4YIaILHOqWHHmUxakqxBGPcQqLfiEwRvTHSwuDZETEN
X41ZcwD0DBokr1FSzYVhX9roDml/lG2jeTnqcW8Buvc+8pWIlk0xab/t4gAEJe0C8d6wsYZd3vvY
/mMpCR5OOhZ/D2ANmILAHsYUxiILvOV6ewWAB1GVAfbhnDe70hmHtOW+9kI+JnyaYCodPImqDQ1k
YZYdn0TcAT5CwQCmbcmx5gjoFJ/F9vVeBiMkixKAnvQFxhOSFdET1+f/wvRUOkKvnNkv6wGslD/H
lOZ3ZnmEYmb+BgJnrtxJ86L4h8tltJbTL8RzyRRAa+op/Yr74cdhjGIso6jpzqmbDCnPYi3DN7mi
pq0jmMapQ/ZkAv6kMkEnXOjG+1/gMez85h+HZGUfNbv3HMnXgqFR3GHk6PQG2KWUwm4Xlwtr9goi
ckhcX/eVNwociiXMRPMGID6Wr/BBmH1Qh7XRsn0dxRT9mkC/z6GjL+v9Ffs6wrtHrwNSy0Icg+Cx
hWUlI/O+diR8MC8jLe/xWf0QbPu0wH941BSRG7FcyspxvLULo7qn1NLBvCzuSorAGQXzPVhJ5niK
/HsO7UD7B9Zo+mnH0ogGgBHjFw80s2GOWQIc+8UzYe7Fyjuxpa1EXKBws2uPnY5wMh9qjUYY47dJ
mGO+3ZDP4TqX+KJifuk696G+89RcsENJPuI4DRf1cwkHU8aVVQ60REuGb9rorWf7eLXKFAvDmuir
XzBcfumlsGQQnfYVVnpffJs/8RdjqNrkYA/0agLJ2YOZJ86D77NWDBVo1sSjd5gRm2ZasT0aZv4a
MPjOgcnKl5yMnEuxl4FE7/8D7XpiGw7QKuWDsSrHtGUfEl7bkb30dst3IWzk5C2deXPRw/2fKQnL
k2sDxDjKZzY8/LQ8g0Ummm1LFh1NQ+HWEISvLhkcrQXs1TgXo/eSGxrBjryVLOFSkOam/49TrKfm
gmUm6vz7OJDryHMfbivkmQH03FXsxIuJzwnwYWGPKM2PzrjieTfxg2JHehN4zd2Qp6wzxpjdXk4H
QUeP1waOyosALXFFYkSEbffoFDZ/3Qu3ZXBS6UZvAFocEVBHJdLNdHvCERp5bhwKCIIok7/jsKpu
Q915kXQFGSD20gXvpkZK6yTnyjzpGvVlTHitzRLrRezhGR+VvN7RTXEaY61HY55uZV5KwUPyyTOD
18+oYWyHY1TYDoYbAIFloV46DfXE9IICpjXNCEMzMCZoxQIwzUI45Md/NJpZNLuCTcUsR/C6fyPu
n2eUX0eOHOEcv17qMlcMXSn9x3EfpS7qwgwWfponVoMfp9UAxbdpWYXciGEEuRZCW6T+Esyq76+S
sqXW3fdbOiLphhU0cUB05x9gSL17kVYvkjFn79Hym/D7sb/6EaFETmeO0j+DlJDud1aNsOhwdc9G
FPwl9udg0RVJqdkTXeikp7iDSoep+hpVH8sHzIcCrgXLTNVoq6MqHfrETubAH+OiWDeeSvOUyKDf
mp4tu62Djx6Jhm5TOVDG59Ie7MWkZIyHqLOJaY3LTXOS0CJITwklqAXnmEhtaKO14FM=
`protect end_protected
