--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
bkZ0NncezlOp555yT3AOKJEmBN3dOKU6qH+7/GOpbIxdmKLJ/rpL/FmLmIzU4cmjBEZ1aaBBk4nV
Gu2VOGsNGRDz8TelNk8hlaCsDwceM+mVVu4E1FFcD4R3H4UrVd9q9YR97vgdsWTSqyANXsJzpJNh
4wo9xYRAiiAe7l04mg+Y+xPMtWJYkdnwBNzpnVGTX+t1u52IkPpr0ZEunQxw9xSegS4eSdEqqJJP
VNz0cY8FSG4UKEhx2lpgYaiekVNE+BgGYbGumKujEX06jBA1K46mds5eecGObAR0/aj6YLTK0pWA
KbS4TVCY0I73l0tb3gxFIUBwhJR8eqDyqEFTcw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="VUPxSmuHM/kRThxUq2awPG+efRBY0E0Ru/SQi7ZJiBU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
JgxDOpnRkJnQjlBSjgwguD7leKdjVvsjGolP4sbtx3X2M6jZUONr3zPWrGSiBXrOpeCmjFR8+WrE
EOwzs/BWaELMgGNxlruSqd7czlr4BXHnG2dwX/52XqhRJoWM0uv0UZdrc6P/Piio6N32gHTaYSIS
nZme/UEvWkPLUtJBj/qF7G6totC3Rq65IHein/aL8YlUUwOJOQoflKXsiyOWeO3zDgXp9TcVb5eV
0S64LPpNHJI1vrt7q0Do/hAYrHpLGZCLOQhNUMoUALhKYU1GKuhslDpZVBo8WYZvY1vfFjZEydAE
csuHRupof0xlF3pVlik+WNwbJ71qwDfDl+ELXg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="CRReox8PZl7eyEjbMA48vkiMa4kO/K1f3HCevwy6LLI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6048)
`protect data_block
STiQEYkQ7Z1HbQL/EZOVOXYNjGgsF+ivvRMqqlWZtVcwiqmN8w3hmi9YIRJbiELS844zIiwjuU4Q
CIELWEnrCVfeJ6yclMoa3CxWm2VbSS/BS6mSp6em2b7A4doplNEzxUPczexxHUBiJGDophqmln/t
Jki1WVrpISZFfLhuTtP8/beoj2xo/OGQsajKqLz/tlh+Q0p2mw7JW4llUurIt6P7WbeXnzmw0ECP
/UXI2RaVBU6hcRQlxG9hwEHEUL4P0b7HjwP495YeNPYgwq6zABW+r7a+cNcYzk5lAXabCHC/J+bj
YR/VW1NXVIb+hci3DG4mq5ug6iyci929+Py8NGJ8usXV2HANnRStCI0oBjxVM7cmeThv/9klRN4E
HQUdWN9gWuP6XClK75NijW+btXikSTCvfA80GNL3XkmePjGCjmrhaTa7+PEp10JyDq1vKbxkzQe1
BwE/46VIsCmtpKxQ0L2TP9MTwAPLaWTqdgvAcE7OiGwS5L0GZbEWEIYeTRGc2o4Yzf6XvaepOypA
XpNDQP5DM0uQhj2rhZN0A9ruhgw8pLvwMGegmLeZWOHxqP394mcxLo+4ctr0iWYnx+kgeTc7MnVS
8em5XFlUCiYp4ugqFwoZdEwdAuY5b/lEf7bq3QMk1C9Ehly6HFh5AGCWnPFEvkOWyav8k6a81pkd
UWvrwpPP3Ne76etJU/L/AQk+ZJCteNyp/WMq0xnqn8V2AGUx+Ft/4BwxUDZHcwG7K/KLmsWNn1jZ
BUcQ/BLTictZefvhEA+5sNm9Qw2+xnuXrLgGA/+NeTIl/zoQSwq3Iu6tTtffJzekSm/82BShbqOj
M/1v4SC49C+7OGkmHU/HpS7HI4CNaNGtH2IncShcxSdC/ATtg3QYJnAzb1riJSlkyd+QU+Cikkpc
o4z6Rd/FNdKDTzCv8+SX/h6buUA5nK/sKvmmNZHIb8Qse+4AyQ4qHHQbeRq/crg8rtMOrZwdvrpm
mYQHilCh19IDW4y9XiX+hmDiW7vItKTl5edfhJkMbkyjbS/6FfSxsscKd3lveLc8jnMeZC2JvNp3
Gj1U4lkIQThyJ6BH6XW53A2v06gV+kbNHNyWw57VKJiGxSL0h2LSGeA0DG678uUAUq9nR2rzHaSO
da115VE2e73NWiHfSp0xjFylaWH9+wIOT5/pecl91vbWBrQm6evYUnyzUR0JZ8WRAlAzqWbTNjQ/
u36riOTJH5ylJ1QnhBXMu4HrEaHBnhp9LQTqrBWobZTm8Hk3nUa3NP+f0RjPi7/+yqBlFC/e+Gjt
uGWkav6TTkmVB6EQjCOKTJWMFjLx/gWhBZOzgyBNdemzmJdcJB7kF9q8kd96WfL+9kZk9YgQA4U5
hWyGN4R3KT8CRHL7qmMila8/tqpTwf+6UA4IDaLHAM0Pd0Az9ZzzOZ9+QMhs0j7YpTc7bB61bENK
nc/fC4WCyUSeQnhwWbJOy9M0X//n12/yM62KwMF9F5xhtCNglSOHAZq21wJvmf3DjUIZxt+155+T
O8k9AALZOPxZtPfmaDd5U+YAtEEN6ZGut1onOgLzk2ZnxpKU4GEsxTvROJVkrH97Lmkps+uYYra0
QicOoSaeN4wWzGI4XUb5X8zJYXJwUmQVzE18m+dUvl0owVPJJKFDKYF96I+cbBw92GiZAkrxivby
ytbx9knjYp88jI/mDRaU0q49u+THonQeF34y1kvroiBWeFc53DgyTCBVUBqiVLlS05lCIqQD4oFZ
F3OVe6DXoWtsqGdrfc6efiI848YJa2xlA8pElyxMywYuf3vU4OeXRhWnLefSxlUs6+m9vCf0BcN3
Ns4ptNDTLellNGwpEZe92JAtO4o+yYd23YO+Owa71XmIVO6IZq59jzM3RnHA0+EoDbETh1Jnvv/f
MJDmd+llH1u0eamRd7WXoklhP8mjgi1Z4lGq67hdCBYm/HT2l7ZYPgXQoJwRv0APa5nkUxS62yJv
ZRL/AdkwiPktPkLHo4QhpmATkhsHOgOo1TFf76yGXEiPawKrA5JnuJQV4bVjnW1uoSkrsL/TSc26
BwJXAQmCXxp6m5x5imt4Qx1aMCB7q3dzMRrW/JzHltpzqz4O+dW3JDf7mMQVuVvwDw/CcFXx1I0M
l7p2AuEMEBpFAYqsrysdLUswyi1rWxZl0smWZsjcHPUxWbjsDXV0tKAXzShSTHXh+ZQ1Qs1s6hj0
EQZzaEaM40mLVGjbnz5/uRccmdZ3ni2nuAMtFf7nDhuuKjWE4fkJf+jFuIFO6kDubJOFsOLsrZZH
4HhoLQhWeVfYejY4jMKtZsijAiHVfEjVlYNstxHVyFO3RqrCE6rstRoRFD9n3bY2bTAQ8CRMyMjs
mtFxw0P12+0ixeSV2bCz7boRDazjxJsTMxnIN+lFQXBQmn5OJndfkCUYwT6DNBre/UOandKNOp1H
dLGIKhlNr8NWKRBlf45mlR32ZuXGDc2//x20oBKn82yObrzf8uWp665OJg94tvkdmQIOk5uMmpsW
0Waw9Oz8yHdH9lBygoi1Qw5ePcZs+DZ0HLQD4QyCxvRlLlah/NqSeONib2Ge9HsKucV416ZUPDEQ
azScNSOc5NAB3hIXtKmeLIRSWzfGApBmnrCxgIYBl3x67RXKlPL3LaWK0qJsZl8ASHZa9vIHwCYp
5eMJaSVAKDgF+pbLpwQTg9XbZyUW3kieD1eJwT5kz/Blt8XuYe1v7RPZGw0ww8EUmEyy3j6nqP+/
RmHUxq1XwFIX9wLyq+hfEFMI6QHlw/+SsYuUbWSYDsFdd7V7VQjMX1w2h8Zx1tmgAB0no96AHqva
fWmfjqFkLML+k3BluUqC2AOreignOMmaO6jfq7i05em2cPxUNk7iMhRMcVVwk9fPzY47FPzCctoD
YBafqFs/GJATvi9VdnhPeWeaNwTwcPCEkiqUVotyp6gTw+6NFw64nYRSOsXdk/mSZbyF0yLz9W15
fli3OFPr5acg1GAjzIuKCs6fkpt3tSYHCDlQgFH5OqiFaW5qRfLMhm9W/5AyXFk/nUnE+p+Fh7Fd
bOF27TwNQ6tvjLvKUDMIBLCoo6D0kLQgPKC5Y4UYx4+KLBwmrWNsSZ6MbWMQ/eqxpJ1C9++RiEyC
o5wINFoVB7ItSSm3L1j8SNMuo4U+9Bq/atKkGbhRY+9ShZIfeRXgPbCPhfpLEzm+gqNuA7wX6TKq
Hiz8bGeGjEu7fEc/M1oqUh85QgJHuNgpfqPICZE6yaIs8Ko98jrZHcnxbl6mIRWPx1izLiI2YnMF
V2TCSz5tNty/QCG9HbttdF4OUWxc2Qr46aXI/4MJp7BUWHVlgo7WIcJenaAOGe2HtZwf7h2u2nMh
uUdX61IPbheoMRxuFp0ODgvkRDzxV6MePf+ByXIOCepj9PiqHcSRohQmAs9RXUeR5DJTd4LqrcIo
DCS5z1Str8+ryBLneBE8XxZgMA7Iv0iFD34rJ6/7Rz/tmf2YOpG/BnAQIrbXIQJjH1zcU7rPoBeK
fOfHtvkdK50A2V6Wsijvgu/tiLmcqSdNGVcp0E3rzb5Pf/WcdV56zfETtCICMaD055VimvOSjdh/
rc3WRtg43wa7jO9cC3TzJVRG3KYwuC9HijwgORn2N8Gz0R3mFYoseGIkZoaCjqNGAG6aqAhYap74
kOOJbywWeUMjzKUxK8KH4U3s1WZM+CaMGfbzOpdJkPRs8Gkedw4uqp96Qt0ANK1/OwmHM81Dk8Be
XayJWsPerd2YeBHQUBrYsGf8qIVk/P31R3prrjMmp77pfWQ2PO+JPNpY1ND2JucntuAYyT1yhz2f
JyxW4o4Hhv5qDfMz00R86LQgd4n4eFokfa78an7AVWuI4bbbkPzP6TL5TNmuDrGQ6F5O4efuXxEI
6PqlO+e2yTYkCmPOtR+qzwpgZ06mevz5mxfLQ4/KLNS8XkitU0Ltibf3hWvx5iicTjLYFzK/cyTT
H2vNpkgiFl7LUo6IEboXyODarXsWoLJnGe8tHbucI7Z60wiSBWpfTodSvHy9I4GLIn/GkcC05Zqw
yjhmd2rmO8ar9rDXrrYxzfB/vZZg075KgUetSefoypPXChNxmfKQLQWVP9QtCk6Kw4I1GGN5/3nO
vdDYrx5m9G4IR9zXK2v0j4MxgkDtGP0DBL9GJ/nAvTQgROymrJHCyn93vtMw85uL9k1HL+fQct1y
EW9nM1gWkNUVNgxcvsUSiO7maC7mlrhDDYSUZuCYHsk5S0GszIJDdYwV3BSF/bFeU7ANMI1/P4JJ
9ZxRXDA4I4yM/5mPES/Cp6iOvR1QBY2FMLinLw/FaLdmUNhASstTfPY+VUy9qyMD8vCufO/5KRLK
lY0pMWegmjOrCwvQxcZK/7JKnw5LIARb2Y9Sz7k/lz7XHjCbakPtCyjfRPiCoqhG0vUWTCEBVXMB
F4yMmAJWYBkwLu49GKZBpi6LFIWYHr/HjLd7Ql6IWxTGtCQ/dmlLDXe8QYV2f25aqDDzIm/h6/da
O8GQgQGk9RjpKJXRqAN1/MBdJRvJ4G5YR0elE9+cx8U/6CmYjc7X7ZbjUJFYXQPXq1zXy0MkO6Nr
uX9+Sp/GvSFH62whkjd50iCSFpotwD/DdDq7JmVJJMG7RoFiGQqpBItdUfd75biAj3SZJksNKCTz
1oj2pRhpF07ohbTPWuT/TlzcrYc2a7t1pnqEHtAdYk7ZKDAnfzUkwRKL/xUU3GBPaMIevjPdnzyn
oG0XrSEZ8QsBIIPVWKj9WH63RWs8LxbOsG9Nodmmd4kBx8q7qCTyidoVV6aJVEeab5ctD2Xo9c3k
tsNyfP5MP02C52t4HNwf7d5X3Bh1iCN2KOdyl2CT1TDuIPchNYVck93QAMNkfr/do3k1n/+HD0eO
pixvUQssW9mI3dsYI48e5OvutSJZcTumF3REknfvA54430uFThv9pGZwmGJCs5kUFrOXJNuI2d6n
b62JglqaCAwWOcHaAQPT53rUvCKDXnzflNu844kgzUbeVEDwPw0lA0RSZ6Q6Y3UyonKiw91b6IvQ
RbwVQHev/jGLUCrD7jMCn1m815biVdcrHT3iWpNMpa3fHR02D1LggaulHxj71pyyL+/owEwnnNKf
/1J+UUyVNb3OMchh0Mvlw9uGRmPyKF2A5J4HQY7EhfsJrW2Xyb7q4aYEZbpusG2jUm72mHCowlcn
eZaxilOhmkbq8n6i/kCVWBiXHWncO8ioyyoH4J/KGEWnyHpDJ6fQIdQyrW0MtR+XRF9MEEFOJFA0
KEoHGp4aBbu0jFVMJbSmozZhwEFPABmv6XAeHWL0RMujeW/7OhV3yOIqtAfaASScCucOgl1SkGaD
iRw1KI4q2r937Bl10JdRN0lWNSuapS8jaMfIMP5/9xDL59h/B5z9fu8+wbJZduRZVbjL6I8i7MDb
kvvJfjeqJL7GGpDvXi+5L516r9fpPcVRYY7VnxwnvmK4uVF2vDLTt4R6JMqZ8nhZicnwOZm6EO6E
oimGXmppuhvYgM9U7A3EUdJq8tnVwx+00W8Btfb/Emehsc0tPNhdDA/H8cMlJ5ur3OqTj3q0WYPl
PEFSf3rzfEXSZEYPgFLRdRd4rfmRW8cGBPVNzALFD/nw2JLNulewVn8GMhUtp9tzJyWsNB/UMhG3
NJV59W2x5YmcaIFvuyU0M15enOHOOwzi0YzOyGMv6VhVB9hwKIze+skNBRos0lnsfyg8e7t+mYko
DDUUstWmpH8KR8rHbiXXlLM6Q+AAw8yVqNh8hf8I+XQDYPjjRfoz/MUkK6bRk8W/33W132G9rCM4
TZjm9/NbuSI0SNohOD23fmsIyLg460wv0anMLZDF7zX9OwxRGidmhhXcN092cnet1OsCgYtan7y5
U07KyRnWzsEDJgXinku+3fzFT4xw2dGL37X3lB7YgMAyHU823DLhS/2pJg542keAVH3zED2m4wXB
kIwD5YcKd3Yy6fxppoVvYcSHqfF8gSCvYyzT1ogI6QgOoboDuWpWPBvsGF1qTR+mQ9nyy20FKm73
LJWiGgZV5C+QjXoWG5Qa+xu/vHJ07Au0/1F4GROx/YviaxXoy6OFJ+tS1o3vdp5vzNBR9K0ABNWE
j3bUQcMwpDW4FuqD+LDcQScumfLZvgmPnYCAXbbwn37cWeOHq35mW3eQKvqiXEue94AXYVyU+54c
zaq0rRxTaU778CdlIrjGrD0o70uypqWWWUxQUso6b0JKwhWKhhupSBCAa9SHCYWwuoVqfV8zJCEz
fiJAHQWTu+Lk4f33wszi2FKIdqahcKoXySH0pjOgDeY/DM4a3SZtdCess/umaAogcZcUWJP8eqo2
+tKHKg/Ggwi3jkCM6kXqaWaYyplRDkUpINpVN6gNoD5hzv2iu0xsTq/zY/73IMJbIVMYPdHtcc2Y
OGBgI4g/Ol+Cl9zj93ig74VyIzuxnhRtvb3jQKrCjbo77TqYfpOrNe8StcODj6Ni16tUvHDXk9ts
CwN2g8rIh8W3coisBVqk9ml4+x5w1cFh0jBIc10T5JEW9hLPJ4F5cN5TBithmdkJCRjlwn1F8e5A
Hv3DdD0jzrJ7lTFHrN8KMak8SVxNZ9C/1c6ZsQmFwLW+/rojE6wjoXLV+qosH2aC0xp8tTuN3W/y
YTAC/n9yvk/U9/A2gDoCILkVwjy3YmwvD/9o0f63rAqU6Q815elRpe8f1s9Qr0HVm4MebD0dLiet
Bc/9b0JGR3JSzN5b7STrgMOKMckB05C+F6vokbHumxXe2raPiEfI0LaN4MoyUWgyodBM1DeTM4XK
+lpLpHCf3d/m3ifp910uBhAbSNF9JeUmsSgcjK1YV15z9Kp2jwneGVXb2vKrRlXcz8hXDuaI1NAQ
Svq1E7y6Lcp9w015DN38HOXV6SdvRRnsEqW+mX3WPZjW82vCgRaRsnYtkV6I6L1YeJ4jze9QkYxV
hSHYrhvlwOFY/FmbxYE3Cx5dPdqBIh7tNWvHcs3If4kc0XiJwcx4ZORYP3vgk2mSMmQF5njfgkuA
l2NhsDmc5dj2h/Ma2KDrHNbZen/Dkbpfr1oHgVUTWc2Hentau2Gdk2tdkZ6OR5ZHRV/jklWHTKPj
3iO3/hUWZ2d2kRaKWEI0c/0ztg5ZM1GASwwCSMbuXr2Zux2DQYSk70lG+5MOcXBnG7Qvg6Q472zG
+GJ0AB9IHtekwt16W9Q/KiljJYgsyussfCbVjkyNfEpPPks5mgxMDvxFeMtQE/bmPZyxGlW+IB63
FKF1+22xbYVI8teVjvbxL+h9Szwe59b7v7GKww3sy2Bs/lFIqWpYTsW+yOQ+yfXQbvNsjbbqxlmS
OYOHLcC+Exn6mlQK3ZSLCM08G0EXIjutqKMv34e9mvWXOJtr/l7Nd8JCnv4Layoq2wBFf6REaEZs
LFYo1fsyZLnAn/tn5G1osNIQco646QwIRAg8gc/jQeq7TWmLU21nH3TYPTDexycCsXEWzQRJB9Xm
5cIcf/af8OuVcrbMqLfe6SIX/1sKBLXpqUVdXqWL/xkn2z+ZAxB39xeWBx2/XIzqwnDzgh27/g9I
bA0IhqYnHEci3aa8LF73UPeGMjeyZxA1iDD4h5Q4mDUiw8T0hLpdbgiLY6HY2Ve+Agi9UKu4Kz+p
sR7BIFe2UdJKBzWU6YrReAd+9m0OO2tfejCF2zct5wX9+NekyzPRsNIWJqagfPKSBO3VstU+T9lF
6goT7c9abEbDd1AwUza0VaPu3OtX27udB829UvNAGz3GNrbvE6hb3536ue9xgWhSEauvUozo/bPg
+8jGAV1YvCSqCfWPtrIj1vKhhIDTd9zi0JMfIBq9X4G8UAHc6VJCSZ59lrgM0+JfZZ91YsJ/grTc
K7HnxKTlNMdhuD8Sy71t9erEp5yDi7V3phMtbkUlqv8Qlspbx07FzCP1LZZJm7CM1pQTCouWhnoG
26vQPwjxGh2DHb/BXf3VgffdHPqpTNMnFn5r6A+no+VtCWYBL5lUPg+fwh9SX2M9S/+G/uOVQsfV
vX96ZgyzvhyVcxrbuXZvTXs2kimw4Fj7Ialbcr5hH6oiGblrH63WnqgcKcee7eOZQrvn1AORrGGF
lVtW9OVx
`protect end_protected
