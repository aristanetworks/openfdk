--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
j7JRCQ4WVdJB2ofaZ3l4WsNCrne+AEt2Rlaz2YwgRDpaOGqFv/W7SyTU0oou5/Ma0o1E1c6NWYLs
70QuhDpMsmxofiUoSjzmfxS5NYY/M3/ON65aWTHYSMw8TFlrQaoNOmve+si1NYRPpB+mFbAc37Wb
l1Dty6fjNruKvV5KDB7TozRAp8PMC43LdniIoExDK2LjxdcBDdT7HSDtqE+CTBB7PZ+ma2QlhfaQ
jXBbs8MI8XtzFGee82DM5KVtJ55q91GY56XLQ5joLBk/yCkqY2+DmqJmj9BVupie9jAZ0CvnbwzO
i7Kf5VmicPZF6LZJrBybYgc367owHIPjx0IWkA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="svbMuK0uTivzb/15OLwtAoFY3I886A+m1h7ECjGVzSk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
iaheEMN/fFyNauu3vWYFaCBJgffH5cpWiSzkPjAQuPmSRWN13FK04KS2AtYN9+WR6mAl4tt8yz3j
drix8uXQ3okvE1nVgFIv76ot9bXtCYgNVc7xJ0NkjyZIs1Y6UJjrTCvXHHgP9ibNCb3i6uYvVeG1
F45Gx4ei5mg8k+X8/9++IVPuNt+rF0gbCW2WCClrrrIbfGy8ARVWohOq0FUcieUl0yq7/Vs2Fy2g
CEBcf9x5jfdLM68TmiHexkcCq7rXKZmIdGl5fgDdAoqcDN4bvChTfYkmhRPHnajZLHpyAcoQSku9
x0rlQFiTa8POPml6gKyN8d3N3km8hG3vuIIqRA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="ekbV589ycTQFzpWv1dtq03xm79p9BhWQUBV8e+otS4U="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6032)
`protect data_block
CsAuDvjSGfqxN1MwtDK/ywm8DcaMatvD9dXPIkSWqbAmbwBytYS+Ofr95Ae2xtGwyUYCFcdVsxIL
KA25LRaAeAa5YZCS1TTKSf4dNZIcYj33Ku2/KAJsyb06HDw+wjK2KYJKugmPBPKnkRiu6714UeOI
9m9EQOAanGxpMThOaQfp++pSewkExTcalT8IZi3c66JHcPFg/P4Q5/bBhkZmfoRgXJRRzYCB5oqG
qCZITaJALPIm+AYn7uk6waZKpNr6X+AnwvhfiiEXMYM0UYZbRD3SuO1nU3nlqet4CnWMA+1Rnu3/
XfvEOG98/6uz/bPkGOpNI4VXUB/e9XwjsClE3LPP94yJpwiwiLZ614I91DmvguJ4YB6kNR21JvCE
V5C4Gob8E1WwRwg8qe0IyRPialuxzBfo65rrtjAHbnWhny9GSt/+UcRLozMrtuZYbBUmfg1omzlP
8Em0qFEEtdA8U9GleD365xvaJjzxyZHTlfebcWoLt3fdI1QQEpRX0KQfyBQosKDeCUmWHBzHevKM
o9l/xtRjWsMl/S9Em0DfvBQWR7B0Kn0u1OlXTGEpXjiSB7LTzvMgAjnCH8EL/J3FWRKM4g7nhjfe
8d2c9g9uTZVf9QAaUjMYGJKxSRldOIXsmoTjtYuM7fNPAHwqzsGuGn36uKTQmOUK7RWlw3R4ld2Q
ANsZ9V3Pq7Lo/JQ3A5ww9I8NP/pIEJCQlm5SOgboPgxEiPxMN6nNIOsv6iNBkilwR2E/IrGVq2TK
awar7JgRIC0QmFlTrk8T1B80I7bU40IpQe/lY9amv/gvHTVtHs/x6EDzsNQ6pTj37CFeCg8Kn4ap
T2kN1FO4vMwKrk+o69xH8yY6WwwMDZi1n/QDkk62OEkNWtXluSs6HHy9KwkG5PMS01Wh+frHITDk
0Gs9EMmGJblHGQrQ1JSfS6m7/7ZTcOFAV4YWIFoJBTCMoMzd0LjBW6opBwkDe6Q1+H+1JsMqvVis
NsFaLVekHENy1XPnrIOK9f7f9veg/UPGLcgDzvVKH3C+N0AKqfXvEaCSkTqJyc8C3BmrevU/8OzH
feoLYvkIvBiSK76Jew6SSixwsz1a9AkmOGAku7441FDAtJsTJ7mreIQUIOMJ1qQGV4swTSlQNcLS
fBTlc0UH4j6OwDvurG9ZEZ3a/xQs+3ccJ0nf3/ZWKXL2g0BrJsv2oDxlMv1+QIPRnSnDgH3TE3Xk
KxOZCK01TGMq+fllCxNy7S+RREnf2Tuza3EHVjjGMNLy55OAom3uZCfm+iPK5xtmFlyu197ZDjN7
nAK9jyqIY98KVyhA4ZLOTD6Kvs7a64Nfa+/tU5h5CjV4CsVEjXbVdGLx25farQYNpg1eHIOwjI6y
lbntqSyL1HEy3QBkeJ01MoP5LSZUD8cACGqp2YIrBIz/Y/SB9+NfXOHRfqns2uXfSxuWPLc5Fkvg
iFkt6dMybymY0FeRIDnE9EJWi4z1/wN0VThL75asOSUUilJ7oG0NoHr4GyCV+tyhSqxddbJgYCG4
kLHJySakcQx26PBHV9hbafUmHVu1QMgb9ivdcahtVEX1wEsJfIPaTTg1JTwrd+mb0A5v/4T+sn/W
H5hqAPZoz4S/UeHbEzf8/OyTvmA1JIKuIaorAb1RHVEYW/A34gz/ahXvxxK73fxz7z2ARlvyXR3Q
3QO+gELr4BtExRG2kH/tZq4kmXitKvXxYv21bmoi8O8qarFXqzvWOd0L4cpe2J5acg+yA7RZVX+S
e4PPjpveIst4PLeL/TN2/Yr6/8yafTATf1e6GLYnwsOjC4sjrvFXRkdTq/a2jXzjVyPmLvE6UmIt
kV5J8lsBd60srNMklnL/cfGRMfRQ5Qv4FoLAIOJu5KbpOcvxSqG/V5s3hitO9/BErFyFd+K9lpiZ
EP7ZPks/wlATz1qPC28tgw6LRRD7VlLkzCVjnDtZR/bpSUwbhsok/8afwe/PI8W7udEsljOd2L4E
mQNHiM5r+dmkOiKHc4MqJ9uEbHs3nGaImc6+zHZlenzTxTr/DBmZLH3bGRLilJRgH2VACjNdwRLd
zYKHPSQyNWQmU//l7D/LJwYtgFzCG5ZNDBcHqMGqMojg8mFmtHPMe4nbOkusZwI0/6ScLk8twhId
WHxAD9eMHGNcIGcccxqY+PXoKggA1QcpZ1tuOYXBTa7ZCz0pgwuQDAQ4rlWfStM/4uuEnVKJaGXu
H8Lfbmsiyf6RrLdAfxgSK5flSZsSxep2XdcA49hUoEA7urTirECMdjNwrVMFVlklP/HeVKusg/UO
/6aYarIcdDTALg5WIAFsdxXUw51u5NB87rt4Vbielffy9An/EjyiCM7DRPm7/vqjrjhs42quHI9P
SqJNiIVxHhMIM+eiFntuRru8wbDjf/FeK1lRhigZUDLvDfkqaJEdCql5nXNQS465tqvg8VZ/8LqK
LVnGYWFm1Eey+py4oW80AWCf5DP4lZTOAQYn5YUkp0zFTIfUbestTVRzrS2iaIEJwxJMLby2mRnx
uKtEqmzGZvj94U4gOBXLtpwLL1J4opRpYYiT+pDn2URH8O9NPBFPBHTRGUkmBxA5Qsk8Onskjq1l
xnlI1zhCqKf4R8TwAF1WGdOmm1Wq2+jwANSEnayh9/v1wOpgv54MmBlfymXwNVgCmVvNm/1NIwDO
N/Mo7q3QX5oHTcbjzfbZuXsneNqCinyBOOuAlu8efAFtBz8O9drvO3OZlE4/f1DstNcKeeOsGvCf
LK5Y28KxlhDKN/IZY0NPpIQDGp8gnPlG45/YKTfAmzuQ+dghLRX+HFGVdHCEsTriEhlXtXJKRT+i
DARMZu6AQQSH+Z7btngVKd7q2RljiVp5vARGhLIsjvfQitiqh3qyHxoqVd4avB3hihwK2eugeu0w
CqjAChblfaBwv8oPzsyXo7AnhQU9azTXip1LZVOVEru6WG6JT2M9ndfSN8yoewAifaqlnaWUhjCK
AaeJ9QTAN+nSAFfhWijYhT9mO2LFGZvR5QjOAVrWkPnwZYC/5qRUi0maxP4W922uNCn+PuSa4XaC
3+za46yTxUtCyGbAQMx2oskbOCS2WxoITJu4hLat0W2X18uNePKIirz6X5hQTlgh6D909aRTfN1t
ValgWpgDHhSEyn8drt1QdD/JK1ZyWuMchJx3utKSOHHv6xdEr9tPvTkBuXRe1c1jgIcKa20EwSky
OLJK84E2NFwRy+Sn1Uf491yvC/xVhTuSYV4+frlRxp9Hi0mtibE3+Ls8wAGneRWsOg32Vo3TrBUw
deKXTqmtqMw54iymaHEuN7OyyDcyI/8H7rkhiy2u9bSw1LAwzCuIET/CDFxpKNZdZJrpL26suBFE
VMs1fxV+PWpXPDtoJgkJ6tVYlfXWUs3/uMDCooq3lRjKtKfcv8A3mpceQTe9P/w2npG+y6TRFnm9
4d/GH8BWRAwnvcUfq6hVlYFEl0m02+Ey05aPPr9fTAUBXl9nkBrpk4QOCLVAPUAXZCT9PLothqdt
hR7nmIMZSSZN0AUix+mHLtw09Cfm7I3zjXNAd60zjcrXKr98n7e2jAYHZqu9nlSdjy3vLLTNLX90
h04kLSGMzxQF6dC5993AALvEAY0KCCKlck8BHdSUCgqDzV6KI2QXtmtH8O8Y3cG8ssWqWaMXveWV
CF21VwkxCUl4yWYUcE239xcMpE3hSPJ4a5VTEI9WvSxF88Pj7WpwQsPOkoB5NZaRtWj5f5zCv72Q
nq/VaycgJsJIsuRzRVsC0aD9UGcxTa9fdOCSWa2+fiKRRYOl8WX+y+qlR+QfhmILgGWABA+icvt6
NR1qLQPKoo0Bo/4PA8gIOFh+wmBbzMM1B013BBoa2ExMcelVH9+ZHpl5aJYmYnfQABYZ0yuagBg3
bdP+RNtRFlb/Z3exoJxFCirZLmEWbQdSpyP2yWD7sjRzNcaDqjQESG4B9nNzoXxfsYRVgI9455m4
tX0LDrYlEWGI9wsTXe8gDH/2TOzFbUwVWNL/ghHySRJ1WxVSIZd74hu4U/6ZidECAXgaG7jhUzKi
ki9LNIbb2/5BIvX9OQDiAFtoS3miVeh69r0W3klputqECcHWhDREcvEEIY5QWDZfHj/KasAQKZos
/HpvgBfJZxB18zseKKuz6xNsjfSUgLaIqk2iZ7cI0w7b5ob2wSJ+/fJY0VnqLi/bV+XtP+qdHZMU
HWzwAnadj6WQAPL70B6M8tcPY07sPben1hTxIFLxYC3q1dGQBYLh/uxzmqWuzU/vTMuVpmkoGbkJ
58/zTP/r5BIHAosSVllwnMGGK10PGL5OyCd3LfzvslTyJJa+rgkWiaQ/ew3E5EmS+H8srWBd+YyF
xa0FO/TGaQl+m3Wqn0aV4f8S9ZqPGSIEVgaR8IZzTsPQ456/m3SVJMT4QZzA6nhwcqkpzIZEHjcq
ItNSzsHwa3b2cx8lMYQCaJ+NYZd2XrucNCMdpZcfv/nvYe5qrXpW6upV0DMJ+WI9Z33tdW+uE5gZ
AdNOtc7XTVxnSpYl27ymyMccu6hhao5PGgK8Ks38dRz+gLTO1bLQAkwMUsv3m/0GzXscOhJgZ/8l
FL3KD2XpvWBial0vwsOzSYwgxV/um1YJYizhX1hicmXz6ddN2iSaiPkXWyaNT0p6+EYAmcE8F7GN
kSMpLzsBOVzK1PT6eNFHQAU4ExTz3hcB156Y03KxHO/O/tSOzg2k1MLLTMdXNsgtCBu/YwxfxvXp
hdIalFsh9+7on38RzRPi2HXhcK6NDlYnuZDfrJdhzmhmjpUucxbUTFLX4ko6mjv0TTsMZhr09FdR
aVQ4cyGtz/akUGHa/LoHFHo8zMFOwNV5rLGDOttgpQ9Sx2MgaB9t9gUkyhqwJz/4ls+wisThHelO
EOu683w1tTShUiapOowxbFIrhAj2OM5AYiwqaqXmnQ+h5fgBcst63xFF6Q93NvkNJIcP+pjzdTpF
QsTEzEIUBf6qYQ824HVVXd+byXGrPjlwxjNmigjKmD0aRPNRpPdFbCvoaKr2EjIM/+sQQPDvFdfX
Td1uHgp1OFOlMNg0/8Vos0owNPmqPu49BWw/weZj0K2hLKfMsRnLraqoCTIWdY1ykAi+xKNJ796K
zuETUWn41myN2ULCREYGt8i0wNkctDA+rT868N2tK97AF92VzUJTxkuOXOg51c20SZz9qav7pGDl
zvjSVk7D8v6i6S/OUyqo/KvBzxudsyySwn3NqTLJENjF7v30tLZpTswan7LZ/awj1yGFURoIi+b2
kcPfVyNi0M0jdJsCiiXTHdqjpF3jrmfvcKcYpYJOJzhjUvQ3Yfld8oyjvs5gbm6q5FZlv22I9pfb
2Rc5RWLl+/ApMS4xgwvSILC7IZfMyEQ7jjwntIQBph9sUboIvOC+uMwgoYRnSCR8X6MN+XqX2vxw
ksYFd0zZjUypwm2D2pYx0NgG4djg+B/JJAQ12JZjOyjkdgYVi/tZpMFroCbVUCXzChviCmzIRMSW
lfD+htnUKR/zkvYrFidupM58W1Zsb8BboMeQQ+39SimTo2eskhh50k7z9rV+0EzdkGUOcwwB7GE9
H8H/BTARh/FipCabWmfFbg/uf3T9h6DsbBHw8gLW37A8kS19jom5H4CNRAzyT7t+TPtv3wKE8s6N
8G1xg9+qaKUI7lg67Gv3opL1SYGWfR4tyOUozsGz0xll2IfFv1KxtYZWUutSydA4WdUKAG/u+tfl
9bAWeQ5ptYvmInzQMW0TWh9Bu1Cdi7rbBY9u3wrHrLSGTvdyjQCAQbHtiVMAQY+HvfwKvbdmL5p7
ewvv3nF5RI4LGdh/9XWhTS5J0b+FrWJ5o1VBdn3rBHAcy00/hj2Kt9TNU5hO9Uo7Ti90kT8BcC8V
fkq4g1a4febgsgAtmUW+DVVAQ37CbeiTZxB98Xml0K2uExJu4D+T0TBI1eiHPj0El6iCka0mCVvy
K/tWUNU1xLj++v4Fn6rhUpU7SCtQm0pobXzmzGRWmme8whxK0ihy7MV3huciqPejq8jbp3JEu9cO
IAU3vOsCrlFVCCic8uolBiL1HDp8du+Z0KndclneBRqvYunCOUzYnIGfxVNAf4y5LGH6N5wCv86N
idwlUEz+XcWTWd+BkgS8yspjOMw+UCo4/m81YC2Ev5eJkqx1IaIooBRctnwxNslEWg/vltuwBQii
TAuDcTXjiYY+ozhgOESc/8LorKADEnOCg+GlSqoi03Tn2O0y4yi3Y8wQTAgAlNuxgSDVM+wzPB3p
/HPPuDPNIidXdU2EbKkvCVFgD/FPCfJh18zO3mhHcD6lW6y/PXlpuFBwGndA46OSYyIJZZCeO3O3
+3Lvipze504thyGv4uL4OtKszjMrjf+uAlzYQWa6UjgeLULRO3Zmrqm4CR3AoGTQGPWJiI9DhcGW
XiG8Q2Bk4Qhi+Cl7D+1r89oF3vGNZXNuKJ5zWaUSDsz5ii7e2wwi5DiIKN0gPRD6onrB0PDhtbgM
vIzI+QevbLXy5/+iEMhv79fPddoUT/GyElvZlfC/NVmiN+z5gxNJGQPXzcygpBgEHUpS5m//0RJk
AlRluvzFwj1d72YBEnDjn3jcCx2QYy+DuCESKcDELAvNXNdP0B5ibwqQkqeb9S5P1VzSNKA5OR4H
lxi7LAcwZt/MXswKX57ldq4UjJx+91ES2XzRDDync4v/zKpoebhHnQETH52/wn5XY6DHzWZkdj1d
keCu+ujXIrU7zt0frGqLvDM+iohcjL1D6THxvZLnqOH8riDWJPhSN60LuLIld1Q7MphT9vSWDP/g
LQNogpqnypwCpyRXSDhPIqFO5pcJKlOx8zcXOL9moxiKOlKB9SdExIM/1l7fGrJRBfjzaGwiLaVi
hvLy0LcCbsRs1bhcGHZ4DQf5lAggtyp1GBqDTVgW/CpGd6+WQSlZtCXR8zrYCCYv4qlaGNLvQlKL
lKejHdEP20vGd08RMN1/vfkdRXNeOeRvhuIPaIu6wtz58E81vHZ2g2KYdHaGY3qUWcY/mzRkoL3D
ecUEvhVyEDPIXEtwmK/Tj0Q1WwxzK8SEkne29KGnIGM31hdWXFErRBogy3YQZL6fR52vo3lOPxaQ
6LJkwjaO643SfnUBqwzWawwRDQPwymOCNmaaJD0EUgGZ9vfGguFZSYGcN+YwwD1I6FQG6ULetlM0
H6CgI+QZ0Nj8vHntMmG5jpFyQJ8/gTLBHpMaqE+UY60YMGFIuSYmFRTvv761q8bO7ozZ2dY1X1Rh
9E7TbH/S8ZRCJt4GwUaWcbLkSrOfkN6MJgtH+4JT/fDmXLL9anv6K7o7chkwy9azI6oG5YmlkZnT
ycLyAMVlw2sX9GryQwRs8M8tecCcjl4U+Q0FYmRLE3K053KO026FcJBNotfUKcy90wHx/sLHLBz2
m1X4uDtAt0ZGImkdICd6STNDXyCOHlt4IUeJedh+vyafPj/izx60LW9p5GtUliJtoh4iOStPe44c
t8s/MztR09y0LMwpdsjkEjTNlRAxBOBc6xYiNwb9aZ/5k5VDqOU6svjqgTkTrYJZjqt6Vk5/kwUa
2MewLdO4ytu0OdjB0YtTbCf3q4eSjzBBwpYTsBfUP9qsXX6yTNnRzzxDHHFad+/J/bgnPkPN/OTg
StSgJp4jbFAbZ3UYzWJCZQVRb2IhlSlMcE26DHvEbxaaFAHyW/UmaIszSPgkNFFqDuLJJbm+J46e
C9poMGkdOVm3v0ikodO/eshZXy4t+wnf+IoBeRueC2Vq8hfdnqiRqPbUCIReP/CyYCBRIKkMk70Q
YCvF8YoMOBZBHFWrmeGkriKAnXUwdtV5aKJ8dAue025qMTu2S7SE/7YtV5bkWzfiI6LejygIF9x9
55jXpAK5X7C7S8wSrJ7REdvtFjMb9rC0xztpU6T3cTQKmoRamYUnCzAdQSgviutiRl9ic+57kdRi
IndgEf1RwGt32t2qAkqFPoiCctfzyGkoZzam7RqXoJ6XSKLarGjoHIjPHM+pGtLhWfiNLxakuv2i
MklAwQrxW3JeJ6E6o72X2xdqa2n3D/aNLOWAz/sN95KOXWeIVk8PUT24c+xBy+U=
`protect end_protected
