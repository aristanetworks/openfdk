--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
P3xbefaF2wgTgO5r59QdFGTNdbNOPHoDpBzMG6EKqdFv9yStqsBwkjwWlGk2CFlNgH6k029/0Zys
os/HMeTi4yxvHebh1wKc94QeKzuaA0TqBZLHJYsudOvhCtaTPej1R4m3GqcBGjUafdJFUnExOXaf
WAqUhPJiZct730egPrrwo3Yq/0BDCa3HLcLiYVWwFsK/S3cKREmlRVi+ApUaTUUHx3H+mzqn4Q5T
hNtkr192PyQBxLedsXDO+6imFjvyMwcRf9W0979cy3IM26xZErwMISldCxGjGHJxlo6V5EzsGdRq
Y088Nyv2NpDUww9JZcgUyl2EQjojicEJq8rl3Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="tMaizQmWqWBa2zuF+xnsdOg4SiThFIVnr+MhNQ/0gCY="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
WZeocFF+0ZZxqepe/sNVPW98+bZy/4eQL8jGde3240/svGwnS8eIBRnWanFXzs6QA5RLosjL/2sg
yu4pf6CEgJgbghiXz8ZEQGvbAr7GwAf0vt8mtlRbkeqzWdJ5SJE5Fbou77sHPHSDM8RJzeLzzx1G
mbZq2oLi9eajzhuYw/BCSPdDGG7oc+PP83OHE8yAmliK1l+gwzMdTTh+diZOELWb14QK1YoNg2aI
9p0Zb0Tq5rGYcinW2Ps93bbYRxDkZGBnbXZJuW/V0XeUB1EiyTVOwD4sDE3HcUs5jKn8Hq01BlkK
ZLEpBAa0A4t21BqBG3jaKP2N42mFSuwE+pAWZA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="r4iDAruszBa6/yTRq8Dl1Jhj3Q0fCohHVBUUNItEXg8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 41888)
`protect data_block
MJWl3e0cRbUB83KN2B2IRdeX9GF2YbLBrt8XfSe7GmzJNgn6SnDsu11nFXmvF7XBf5uclWjXC/dY
y9Ock9Dfyv3aM71n/1dRdhFCjYszlajtPYvBR0hkTjQ4BvkEFmQ8fo+7GqwW1wi8AZ6p5uvx+Wr1
scaizl791fd4dq5+Bzpi/wkjItzzxEwo0OYwtnmSjJiwLydDAHZ1l7F02U+MyXqEW/9VmOXs783W
olFEvhH9ZwyDQf3gbw4DBMU65yVulHcQNVyxY289byERvCoywg2BCgmL62hxtDqacpYtL/xA+t4K
660moI6I5J0RvdONGLMDcpUURo9VJyhN2dFcvtG8KyY/JNjHSV3Z2tfYr0i2y1ceSE3WJyhp/dWO
GkXm730xlxxocswcV6PO2PUfFaiwzn/G1aYur/k7JpNLTgmlLvC5QMTIZGvRuHa8A5nFhmb//G8g
3ZOEUSruoo1jxR/AHcdI+rV3Bf7GqgPg72YoQNhqEhqi3t7BsUPe7mawuSfqjPZv52WWBfg7jwU9
xnDiBQ84c+pJRuwmDJKJLW1ZeUq6sckGKyVnx/DbZFawkZVqvJCCMT7mG8/etpXHk2Wcwu0jHYB8
agijR9PPE/lF30UBcbZD7Ub2NnEC5/Ipt7s63yYo/us+drZAyJycVc2E81k+DbzuB6MKg+cxzgvf
yGzoDus7GYUjO2Dt685Vy0gmCP8rwE0kw9uNz9n2F8nSLuMlG4/TuhPjdIo1JWoGfOAFwU+vMo82
6HGxmqXIpzpVc2kmmdF9/98ANBe8nW9sqI6VLpy+EmR16xOKkCNkxEIn+/mh/zBJRcLHo09DVgVv
j+U0xUZFSKu/PcO/8vTUqLOE3C1j76Hx10wrfFqp0y8gL5whOl8fqrXWG1mBYueCvNrH/x/aR+PD
dZQAMqh6RP+KuhQ7NBCGgR8HSEHm1E+gT9cebK2k5tahL/KC0oDDj7QFsqXMNskxyaSUI0ZKB4HE
MVMjSNcthGPQjskc5yR2niCPXL9gXq5n+fbvPeRhPIwuhJMsZVAGT03rd/ODO0dWrfOYphuIi4xD
GR2R2ZsKtWkqN8MoDoDwezgT2FlG+PQzU7xBmdhdgUZFxsNmTQoKsMICR+kXRem9li1L5nCfYpzA
9SRjNAzJ90NgG1C1NzFuK9fO8WftLIQNXJYL70RC6H8dXhJVrfQZSXpRuPuK2FeP3AdzjAsoRQVu
Dv1VbZwK6xxoOEMCQ8zrJ1OX8fz8gwde0vDEcY2WIgMu928ICc3qnSOLEJgs6SvkzZGlv9IHzaE6
YbTGiCKXDErAQeydQmFyr5oJtaltrwfxS6aM/dFGzhUCitOqZ84bll2pw0K7ZC/zuuvx3FTFSdup
ZZ3JiHV4yvK05defKzyKucnmvSEMBkG9ZKIZd/VOdXSSSnMHSzdYgmzv9iTLZyPiqAE//SIbMD1I
D/iy//7rS4h/e3hP2YQHFTa9XFhRgVZgH9BTTQuGW5x9Gepdy2uLWiUah04vkxJ6r9Cs6FFKIWRJ
rcQm70Sf0P68te8K50BUiBq29RS604GLSq81iFj9V1IDE3KHkEj8V8+fxhnJI38bhJeDjrhkSgL6
mRBK6Qz8FTl7UZWCOc3aiU2Zu42Lh5UbXEDw2oc9ra5wi2Ohy93djsbUtzuluRkKK0UrIZ+Kk+Kw
5Zxyapq5y0cmZhAlZuxHxqAP9C25tO2Of66VGNKe5sYqtQwwjrJxG9NWeAc5Yd59xBgCxwSxSYxX
rtnQRN4tez1ljX97UxGo7WwtnkjXyZP5ZiuSWGpaAxKJskcTcEqHv0LF8M8oKCU6BfYZSeP5qLVt
0OMVnQ9Rh+G3V7ShOTx+w22L740GYvWPuBNjL5bbk/AcqZDi6XUEPcRf4M3Mw7gvAkY50O1c40GU
93Kv+v+i0DIOlHovqhI3vuS4HjsxW3lfm/y1BvTS86MkpZEp0JPw6Np/n5gfgiKE8OZDmBYMmLoF
dWzmEbs9ZUPdUPCWD+jGkL4idy+tdefaG6oD8PxypKkmOhurheCgyo+xc2DyLKaQZNp2jcXpLX/c
gj7TWIWSfyYP58YuLjlA6nvCpoXRBLBKaEU7DjfT5itV7i7B+18vCC7STAPAsXxHzzGPTzbLAqMx
2YA6G/fOlTyIGeyjsS6m9PWt4603+slgpuDAQthIpAt7unsMpXumL8xYNTdTo67ubREnDc+bPLKx
tPFZHmdTb2KE0cs8kfP6VuVCLR0QR3QXfRmiLr4D/8ixJ3TWK1yF0MmbOX3k5AbncKx6q+USK6gu
Fa7lbY5JBYdFkh9TEa0H4C4AK5sxS9ML6RS9+e0yo7xikCL1QTvR2cXQfNmUgPeQ3tiCEDY50yrp
aaftUUC2cPB9aaQfuZxyYkcUMpBeIRBwwxkLaNEGWTyJUttoMJ4AH9mMkp8B9VPBJCtTMxnGCqCr
u8FXoyLOJessWyWfmJtQ6Off9t7MD9QLI4Zh+jeKm/k48m6YR3HydKZ85KK00aQr6xXWX04FICNT
aMh7glMffl227AuQbjRKp3iXh02p9TS17P1n9Uvq+eG1ZvY51Xp2Ds24UbjiHgSRZmc/Dw/rkDJk
3GL9H0XzI12o5YOQyAXj/OFgAFbbcEY6VAQEx9FO4OL3Ua1/2leaKnw4jJ2CIE9yE5FQALiUbazj
cb5hN+Q+sS4EXoR0G25LzA9q25JM7MA3v5UIoxUH7uvMnWvWznzIVOa4/srGId7Uqsxhg7xoQUI5
4aLgQiHPIfaL9Fa8FJQR+cTb9mTTJAEUDSvWpbIrE7wBDI4Bwi58RDxaCZYHEEz1DzWS+hApL24u
G93hZBKwXyuIIQocOGi1Fzhe/0EwGFFokGHOpGK9zvfH5+N9FErAXUp0VMJK6zBCUJVtreeV4JTA
Si+tD5IOCmTKvUBp2EH6nuNiucRDgCOjGRPWmlSJ38O2QVUjqMHBgBJ5VI35XlTQFBILATcOHyyf
GIYV8xHYLBm1F05A7kZSa95fCP8pAx1Tvv7Yu+E3HxL6iN57CVOoZDW/KKPp93132fQA9UNYnO08
fwO5Gvekts8aL+eG7LKN/KGw8oE/fj+XGs5Oc42AideyhOMKJq1E2oLncO/ttO/WVw2Kr3ZIQ6OB
cM+TXQUchtTvls5RNa5PYYzH4W3d2S+/qci0ufppSfqPiQG6fW5brBEj4vi55GByfQSoIEr3DlEv
pevDGuD+TmCtpUv9wWAOwVZ+PlmE6EMEtu1/TCzWwY0DQa5axZtdLq+BLdj893VPmkeyqDJxnmGL
sKOAtq46DE3IIItsZvg/j+efkNsUVuoJ1ntpe/3emmEyZG9sAgS93T8pq/kFlu0ZS9RXW0yFip+y
MfQqBt7KMwirRETwvcgdGWieupQHjJzq3l61CGORRdl+anTZjElXlEQsvADabLKx0ODpe++m5M6R
MksxHajIB931yGLt06HVIYJImSMusQoi2LYy6QobMm/fShHTPhe7IcwICm+hHTOj9xhfeVG/lg4j
YwXVyxIfxjGn3Wd6ljuvRfWpL6XpRUS8UNwwIPMjHdikwGwpYczDcXf5apRrwUB4/9gJAzIl4tXg
Yb65JYFTa6uxnzx9IwBZFrvOTE64O47wXzaqqwwpzea62/Pe3HptacuGkPvur8ohXM83h4M4QCCD
uwZZuloVjqTUI511ZmDiay5GJVj0j0G9Gd/l/LLiLX8cTd7S+6Eno6R7CEXI+s/AbHxQIeq/cU0G
7ZxBAVg5h6sxlXoMD9vokVWaSAB1+iJYHaung8/N5Q7s7EgL7/pAmuC+cm9d0X7rI6EvfV6IcN+L
0q5HdKI1JAl0+7Uq8Yq21yO9BrwpypH2zlwbPSoALUwBoFBRMPRRT8YtImUxsYL+ehjRze1IXun1
xwp036SAe8SMB84lNA6TxfgB6ilxNoLGa77hyI7+BeZoB5KKDzLK/n4tCIaxwSDzafGKqDN5WHsx
g0rz+QfwGrEw6MhYxrnQjWNqBod1EsL0v2TLnM6fjaSU1D12XLjAMzUyKHCPeYyRjhNUeyKNGDjO
DT1GInPDsf86JowvzkMLtZ6pWvA1dUQf3yEVAlIOpja1Yzq8VTh+X1M3we8Op2SfTet4egmCyRXL
Tb0ofpeKUXP2oLAt8IJklecTGg768Cbl7hMuycmhAqO2hFr+sn0uhj6+CPEvVsXptR4bl493W9W8
NREv4P34tRwRiHMPpFJXuRqWvsWCFUPpR4eu70fKrHJOABAfgXIyQYOH3GLTgHLRmpoaZX6EpY5f
8Edgc35jYAsXpiy/+nUEgrCTtDfDCHX/cgYirlfh64aTVRnKop1sKGUKQx9bqJwFzsX9Mx2vkJ0G
kUEx4emkhhOd2X4oaFIxB/2Wgxdh8ljhlqG1Q1+mC35WaCe1okQOLnPWq19+j5SeO+TeWFUbKQIP
p3Ufy4tL5mUZDU0Q80MHdDDiW9vlvwRuQWKovDFvMg8ICThx46mwbyDDTulZsQQGd2fmJrLu/if9
/9aGMUJmK3DIE8hyxXNk6iujWCXEEN4hVz70diTNlewh5RqGR5+p31eIgtAqAAjUc5GA9oAMMHAr
YboIrasUmgAPV+pQjJUPDOoXmd2MPIbb4imXOYMg4QgHciLiA0Gl6/TwcyMi14xosiq4DNf1Gznz
CpFOs/Lm4Kma6R1hdZUB5lYpX0tFdh8ERaGuCvZtlntm52uJUkV/QoIZtp6gcmFdGDhxSG3yHDQ8
JVlznKI7gG0w01nbKFFOsy3BWaHBovoJQGsAS3dDXuvUUL+kM6Vs83g3coD826R7nuPxCVITFd/8
/eBn2/s/60q/4GjtfK3o4FDcbz9ZKczijKeOcFO2pXKUyUf3Ldn6YjamZU+PFbl49ADjeC5KMLnQ
TxbIwjl/uH5gaT54fSa2XIBUmtOdilHlM1IgDMR7GODr/sdagjvjhKi6jm0KYrXgAep6XRNoSh+f
x3yvFuyTmyH4DJKcl/2qLdUfHS08SHST2aVKWGxVvG3njiKRjuMGVnYq4cPo1XHaxr2oICTsNA82
GfG6JVLMTGOKJl8PUZCUEt6RRJ07k3abO6j6kP6xbjMURdPcKKzaVDjr+qc3rWPh+Zeom+qyVqg7
Ufpv9NegTjPbm3TB1chGYuDKJYIOdBV/lWIu/DEsbTryE0SavJ8FtEgiyFjm5/4obtKZR0qL5q3r
0uU43tiHWU2PDl/Vp067mKfKX9v68vh8PiiFuhEfV68PkJYWKVT8X0wlJhKei8oTKe9npyN3Bmon
AwWVAqgX8YseMrD1lZEOaM7P7eWjy4s90kylpXMUyVxHWONgqpKM3EWFm+IXYdqfnT2UGlHqb4cQ
jMwNQb3VfQVfQLU1TWRC+quoBHRJutNBpLVVFIpcDkvlc59Vlv5cEn/33YHK9IGII7eikgQV2DKp
O0j/exIz9P1UxWYlT4shbosKiLgQzz4csSauBH4aVFK7d3sCy3n2hKmwrs6Mj9/zal7eBRnINtku
XmGeA0M2bYyAg7j8ghxf1ezzsfao92854XbfmYrKInfVxabVEcuDggl59qBKoE/oPQ6GLmqtrIG4
75XUj9NvoTkEi2cIllBHOoBrfAsks0l6qf5+ZEFUmTaFVoydJeOz2nmV3BF72/zMJTjScVii8iXz
eKlSTq97cceEYOo2azPewWDscxSW/7TSJlDJ+c0qjHM6AAayOBIDjTSV9OroF5C7WoNq/nkW7bM8
5qYlikPPfpatKQu4jnqSSsnpoabKuv6qkLmH96Y/cDjkfLkET2IEvBW9zqUcgPkagYdgaqHzzWd6
WCu4fiT5+ThNo4rKU3wEa7KHaOFBtcxJEylhZUTFimWVb3rWn7uciTuQnTDdCR+lrMM4DMu8Z1tM
eDJcQfPrH7ek/NDq9wYZ0sxHgt6kd3v+NL/eRTnrzhfjIdrkYrDcpvHqwnaiu6MT/QkfHLYawjPL
LgJYXkZ+T1Q+Gd9DTXfylD3T0ffT8gCM3k7KeupaegUBl+X3tQqr63L7CTaQGodiwW0yQ7NaHLJu
hC0tLgVGdrPx2wiGBqP+gq8u8eLMTIe52rt+uHfzyxisZyJbyOjWj6njrruGdVUUuZ/HUoye40CY
W0TAm5sSL4Sd++h41POJ7IHuk1XJPDOQUio6LmCTsLWNL/WGpJjpLL9IERG0AfbCJQWnSpuZxFkN
/SP/LUpiUQ9X4CD4VlNeKsQYsWNj8cIjSAcZVJNjx7Nta4rFrZpPhcrN12qPlpnMgMxeJeNruUze
4Q1SoZMnd+mtpw/le3pfXkciIP6eo4mmWR2/ZKCj1bz4UFy9sSi00eV5bMJrDpw1A5uKrhfIVOm3
z1KhGgDluib+gT01TY4+eQiAs4CUAFwl9Da+bvZ0Hb6mnT4ROgS/olPv0Hg2SUeOGMUvEexBBWWU
zNbNQaPcBbCrQB0ZM8+Ec2tZEsfpLQq5L1rGUsIwWF0krcrHM5q3PwmfbuWAmdQZ7WOpnjgssv6j
1fk2ivxGIGJ98fBHJdcIOtQteKk9aT9NkFGb5n2Y/MjL1L8Rh27V6aE35UUG9VX5YmFWP8oO0xcp
xWwrh2A2+WoNScBLmZi40h+xmQ8EDdRM77YWXaafQZ9bKxgRpUbqbovK8/Yj0mSCryIzSPd84T00
LwbgSWHYcVudfIFm87SATfF9BJqG9NAuZpuNN6FCAHQD1R75FgPepaWnUGtmmrQgqrCenp71sEWg
h0ZrDiBaB5QC+dWYuqy4oqujDM2fTNeP61Hud2KR7DCvXczCpDMA/EwFWmwGuDEg/rvyXqWRh1S+
IBzNnUt1sWv7QPELzNiYvMi0Yl+Vo7UBdn7snEnhhY/iQ2phn7cN7oxPP0D/BS/uYEBnrzMJqvat
u+96MQsHEMQjGXuKitCTr0bTCouNh0Egmneg+55xf/Vgxei0ja65gLWHgqQOUz5OUwkHe5IQeosS
4j4y8648RYA2cXqsxbTc1lX3ZGMTIyW2nkN4eVILrC7PGiEp72t6v1X5O/Y0zYjffjce3wT7yGyx
RzocGCv8ulBy7e9uaen5WLtV/LQfha562RZ7uLW4XXOkthjHiVDJb70jUTuomEK8zAGUa74N7LWC
w6vkr/QF76lOf7WE4oMV6V2/phXdWxMbvsldUWOEZvtLeWUusRN1y2boED0aMp/fYGWWE1sxQX3h
P7+1LnWd6uqLny3mz08Of8sg8ubg1mVp4iQfCoflG0OSrvR3gF8nyAjW61f2lxlv+hTRh6SAv2NG
LGljCFp5JHA2g9tHlMob89mEKwoMPEaK3OB8jSjuq9DoPbJUSObz+QF90Y+nzAF424NIgcw0avzn
705dXoR87nycpVtmcg5kMykPJqXGJ5FUv6HwFX0MIRLUdBi8E6kwvtKeNf8fxsXbot/j1licReEL
PdcwDGeMIyxEgSJG6payRYzNr41g/2gS47+kpG8YVgOobZQoej43KTw7yhihfWg7uDQo0Eeo8BUr
Pobvc4pArvIZEBUX9+Opg0PFR6yEwK53rJvypi4Bmp2z82Tmi4KY4MAMsFWyf6/grnMOge/7E6ft
MxzEW18ocFzU9l6wVW+GjRbTeandJ8CI09YnBl/NdniqbrbeBkD7lnS0stU+Z59yVUfNX1kE+S6B
YNBATeeStu1uzegZnMXTzLK4FUy4tTsNdXH5nJ/ddmLs4oil7q3WmJ/H0Wv/RFeLW3CW7uh2QsG1
95AofOPYfvM1T8bC6p6ROHXGhoxRJNDI9Xc/BKqyiarRx2fYRuSV47ogOg8b7uH+9M0spYclB0m1
NAZs5znL76FBaZxhSr/A8b7mOv9RbsY9yJ6ZwvgeEDFlEVFIOTocOmlTtxqWzj3czcdhwbKPOrPM
cRaunmE4BqjBkHT/SFzg+kIFNzuB0+lNq5m3xmpu4oXR0r0uLM7JHzankzWJKbcW+fyBB82uzTdM
X05JnFkiOwt9Q66LUbH04RsmPacKTaomM4J0zsp4ZzsI/UVuqRqWFpSjNtQ4AiNgUmSkEWNHpaI7
qhDLLx8O17PnJpCONCABcvuTqOa+jJ6dJiob/sNmNwgFxXfDoL6LvZ4LjJjU9SIkcNhEIP38KvYQ
LnkXgcwUnyXTFPHmpXxkmjHlpAHRcMPjezf/iOwSbYVxAtTaMJBZu/1zrcvaKotQoDf8VRh9aRvG
wWSvK7p11RlMF5KR+MsBeaWGoAGQsr+EZZ12T95Q7BhuylEtTY7aR5FOIVqAp4pX/CuTsiYpy5b6
JvaPI4knr9oVw00t5HD8CbF7hi/8n3v9Yq8XlfE3pbnq5VVjf4Foh8Js9pCwsxHUaMVTHe5nBwtc
ftXsYZQgl3hUd7rkE0F4d0CPuYQHG66RNHi126S1IQDDWRGhrKLcn+sakYikv84/AQSE6HT+UOp2
UOXpvTf+OS6rLqrS84AwWBSspcaRA3fTAcSiOQgmMcIW+29H4ews6A1tTcrRY3VPiuLCCRf/E/aq
9Q/8mwrHNCi2fuK9rvwowo2eXbMTy7jZPkAtGuACrKFuDxsleaBT/jboZKwlYiOZhEfdoZM4uvEV
3mJONAcUuk9tgDFuzseZpZ+u45VQbvXMZUrrNmTr5s+u3NyEFR+MkEfXC2O1NXM461ECMoijXByq
fq1UDMdXMh/upgsz12WR++bAc6JptyXP+bFGeaTeE9NnT1JD94uxJ8hNcMciR7cF/DpeoTtVHyRS
ujUmD2Di8brd6FQ6HzG2whCxBrzn2y4k8LI137k6qFHVUpCRNfzDnamGI94QUMEzz6SBlB+7Ac8f
6n62LD9TZDoFEz9MvRQj8l9vKOtt4WOkWrDZcc5dKWCiRT5Wuvqj3b7mCwSwLuOzkslEZa8DRECO
UbfLZTAU1t0S9qB2F0C9gLRQajT5GsRo2PGelfu2lK4ynjaSnTeSoGFtxdnn5bKBlpRrrNVoghda
XArrFSosiAj0fZEeax0Bp+12H//YKl7BXyptnprZmAjf08reQG/g6dDAFqZwf78/t3BGdCzQjpgo
u285MuX5AQwuRFxNPTHRojpwh/fjFSPN8g58ale4cmuLMlfSVkB5JbEetwMfGGW1joZAhR0k05dv
889l4ylxj5nQ3PR2isaaAhahrBvZZaALsAcD8hc/DFHNuHMa60tevURsHfeIl1TR5W8m/uQ5t5bq
/IHhDLyJsOBX3ELlZUujhHxHIqno/lNTJEy7YzTN+RWJksm/3RTYd46On93bP05vk1wcPug+LNDX
1/A/8PwZQlRVyneL5FJ4CT2X59wFc/l5djKaVCIyU1g2dz1rV9a+oGrdppHWiaHR291bSPJR9y28
Elrjz6icwzaUJXW9ZRcHNvqGzPzlXtni22afDh5t/wpM88BgP+Ug8YLym4u5M6LD4N9aakXJ+M3G
l2+/o3eBBK+fD8nrt1Owl9D/z7s8KJNlLCD8x8Jf1Tnl3gSQqsHOC/daEAPta0pvsY6VxHlSc6bO
/lKNondBj7yl+RRbhjAOzlMnrRHhjtGTMraMXbkCWb4eQF1MgyB2g7RL8xgtf+2yxlzpbgf7Wvt1
lfIfdPx97Sq/GHQ6N308MlVQOH2XCdFctkLvo32PzId3ybmNynfxjTFzUZnTtxEEMyckJLaRNOKp
EqZxWh2QTxQIgvvJooRkFGy5kwhomJJ+qRwPqMzERu348/nixfXSzvF9rmsxG24ae2e4WJqq9sos
4Vjemdn8M5HxKUATjYeDoRkjPOkP+h/CDRye6Zr6KpDVxFi1hH8iHpmIwYZmc6HQ/BGXws+rhdTM
GQsI8nxQVCUdJEN68ptwSdVtH7rXrW63Po0ViYNI58D9Wi2sFaZV6kNwtDZynyjOMjNHst29AkK6
rSCSNm18ZAa5GQgtVS8+i/TEvkvZBfELe1aZVkn601xPek8MYrz6tVOGysL7e3avTRKdUw5IgAbV
JRRd4ZbylmrmAik5iIodiSkUMgQpLdxI3ZLBnOFxt0w3mfOFsDYPtXmDNPOhRfkxDc84vNsq94KX
8mdwPlm8JX1TQwXjBnj+js7tveSDTeyhP6U5q8XCKmy+wcOu9bQToEuulNV12SXg+etE/9caTzyd
hEVtMURzbjE/eQ8F92X0FjOz41sMjRyO1f0xl+jLQBL50N20ku3yX5GrmVsZ+4KFD4FXMwYHOGRp
pw01aHUW9D00E8Nh0MnkDpDmPkq+UlZ8hCCS5gHyBNKlr0GfwwCO8PuLGb24pS8MYbxffdRqWF27
clGeyOl4w56f+olz8BBUC3sHHFN1g9Mvcraqhd4PlpQ8I2oSAF3FWZbMGxcyb0A97WtF0/hAJFrj
6Tw2R+8tC5ilbabW+LHqPwmLbDS2cfNbz/BOQIliJHCBgsZf3WhgiDHgeDn1NYUEtk+SzA04ya4m
ZCgOyM/5JyVt8VWyml4zz2t/wE7CzScwii/YmMS2TxfOC3X9wt3amYN4OqyEHEM8vBgGdYKyEL8M
GHPXZ+o9SUoLiLzdEGSB6rRfAQMfO1HvVaDSMZ4TqPS7I5Nbxdy962WN+7yHD8DnUWeyPjnGY+Lo
q0ZtUrBrD4MwkLMdCjUIWjfymmeSvU2VPyXzsCrofYknJceB1LYi3PQjkUocdZKDTAJ+60Trt3M1
12C8qHXAEXNrrt227YuP+noYKerHeEj+P5exb5XAtVNdN55LWO5VWpAvW52T0efiestCoDMqHqKx
WrhRsKEwSPYWsOBb8wFsoLXyibWDm3PGyoqagEOw+Kz2ZvX84ocz6QjGKJKX6j9x+Xzs34ESErzI
U9FDxy45DZWGtJynvlnTCGgYCfTIz4odIJ1oCILH3vQQKKrfrkbc7/+u5tz+beNUI7hWgAZh5vJ0
A+X0z9CuXMwW5z9pMJfeg7Fxf8xTHF0JtPpGcKGRFgcFamvhZFXZY94of8N7nmGKiO7cZwExqwJd
qgKjfCuYAdGLAz3VLa6t9BhWFUj/oI57qvOSPcu/qm43KV49DyNOGi6+Fm3LgQ6dJ+UWN9q7r8fz
Q3w5MP6iYHZt181hTdXpDfttc4Axgk/mmHNVi+3b87Mbfsj5pjMfFPtZjyWcxt2H42xGzItURpVt
jxZD29CdJtsjS6BlVIQP9Fo3bCAaSaskqRLQy9ROTN2KOC8dBmXURLlSRINF7JE3nokL1nMeAs1g
R0Bumh1jKs40+9ecYUlCqG/p0oB9mnKep9ICgHp+57nXCNGWdsDnCnop0nhFqYotNlnN0nnuzixS
cDqhAdCDG9o3xBNItfgqSflL/YlKzeTpn1IuJFw3RPTwYs96dSj0HeeYd6Il/g27X5gkIOwcO9ut
h4dk6yXWbyBhRmr0z0Ah2QK/07Uqrw+YoZEckrxitJjWjYHJQypapkNFwQCsBRtG6uZWhBOY0L49
hXZN4e7IZFtO0+iAn1emY1FA3663mvk49i5cEdaoYlTRhlxhcy2upebnm3pBQfgTKmA7HXrIPHXk
uUi+ahLR9kJVmgZvtxsub9rZMeW2CNosCakiOsahF6Su8C2okSxagtsht+BVOLOIxgfJl7XRfkVp
2eaqtlMeJZGHy1M01v35AO/FvzAHwVFLfkxp+JH4OqmmuR53Ccbn5QJL/UjoGq+couaRcMUzzM8e
G4+xcUSpWTgjKqDgPSD5p8ilUIy7MwqoO/x7rh8UlB9cKLZK0N0Szkj2dgM8YSMXOG1SPUgUG2Wm
iUdL+JVK74N6LL8P1C4hw4cTMB1aWoNtKExcjns8RZJtRILF1TQMJTIoTVvdzczXGmfzcDNwYM2c
BUBSUifqmHHPff2vRB6F9mCvMYGf56OiHGKLueeSxqttt7QflJoj7Mfc8Zps2/3KbapmFOw69T5z
KFCoIvYjPQbjNCheYf4RUNyhfx0t2fAZtvRjHbP6y87rkYSJj3cau0VXO1iPH9IXMltauvdT4bTS
AKF4TT6hxyo/IzcnsZoZBrYRDUDgdDWj2Wxjb0a6eLIsYeeE+kcGcjxZhzpX75tYH3SZGySEcJo2
TxHxU8748PLi2r4N81v+ZaPYmMo5P2tp3sW8jQnzZTnV93+6JmKoVMb1Br9pJk3p5kup6C+6adX6
UVmuSomo792COdwAsMhBysu9/BL0E1HNHrtQrXl/zVIIHmJJMTPMoRa85U0RE8kkmNWaOK+rcKrc
2T6r/eMtgFaLfMXRd2oCJWqOyvWSPH/bAWZ4EnYYuTaCh93pLBZ4Tt+VR8aNs15ZkAQNKRtSOd3R
Y345nqPeWYe9kXfvtYnGCT7T3vTrKaIFacOjAbo/80J1ZpNxMtXsFT1s7j3hAWbBCynpWXkFgKTu
yztGy/aZHIvZcR/MDNjTFfukMWEvDvisAnSmlJTpBvI9kfXDL/ak+CQtNDhZPI8Q2VZjejIRgrTa
4pNOE9Lt51bSkou296GGrgLTG0lcKzYCeaCFAfFjGrhlMIxGt89Y3ew60WDz1JUS5Nv6b9Rlr3u+
d7wiA7NL68VkKdS38z+geQrF9YCdrNyreUNckxY83YeocAmt+97a3LnqHsJ18xakAIMUDEQWrL1t
/xPxRd5u0cl00B3Ydjaj3MdFJSl/x2ceN7TUMVYTimfi+B59B68eSktTh1br+N7h4GCTmbeuqhq1
rM1BWzZq2RA4Bwy1THp4JI71Z4tCli/FOs1Rgeu5MPR7mzsyHAAopAe6GUyAAdEkfxaWot4LiuJx
Frazqe+5tPk54Yt732YyZuLEF4mYAb0q3IoRINyMFlaegT6mYqe3U71xuqp7utMdz1eJ8UkLSeEK
L8k7c2a1QaIkxr6KFA2FJEj7FLygQ5sXY5leujSJ5LkdOE/wptGVDz2Ht7d+qphmcOL3cWPXNuK3
9FXhW1BGfB9Q6mTBVxqeNdxHtxDqtYh9asQpCP7MvslT0QfMCI1W+Lrf1IJdWB5villLdA6PuPjC
IMn/J767rgLeohhDYmZRVYfmb7F9nHUrPJnFPAOnHk9nhkA2zkZYY/r4iv6EG1u7R05he13y4PKE
Khmmi2T26RlR+n0eRkzmWvu2B2LcXkXadb0jScm+76oJpq25lTv2TgF5w2ayCzF0szLID0o9jZOn
8jzjg0bpRrUBI5IRjxUDYtZjWGqZrb3uSE58Pk5B5+fpJFPC9zGmGZZ3Llo+n5Iym4xtKFFhPAra
2JF5+3d7V7SmPRzqIdTUBlWLY2qkBH4f+2VnWJiRCzC7SSPnTaINhgNSDrqd6Zw2MGTKR2Gl5uVe
zD8HiT3bAaencZ4PeEeoyuqBqLbIWBQUWNINIqz35JcFzAN/+Qss+RzigOaMmfpa6YvDGArap4JY
6bpd8P85nOcWy/PJtOhh5+xC7yzAe7kfmfQ1tO4adu+xJnHVe6E0Gn6yo3XL3hRo8Bn7e+s/r4xl
AfX5nUhupl31de7Mirj8IlXEDbl47fnhUI4n/MD95xu/a9f5evxhYZHvLY5ZjlOkrOgtR3aMw7YU
ADdmsp2xK9Xb70TwGll4jVlUbaGFiAQU7cxW2W8iasi8jApXBQqDa8BbpQTBZODxAtZgRSUGZQQc
3Pl3g0crQ/kqoPDCYFXvOCDDVOoJPSYViwyJtI5lBr00M9Bnm1wTtwx+3qoBoHr5/2SjTOZ20hR2
s03xqimaJfj34FFe/bDGc0kIICBtDFKaP5j3aeuf8XxC1+z2bVXeCL1b6mseU5VE1KA2aDcFfIOL
/km4egbB/APVFkTCNJplwu1K1P3Rs3lAwbRpiAAB2vi3UZg2bnRGojBevn6aYlWs0r51RRf3QXaQ
Om9+lPVs37iOnvnrfpfn+VZn4VAvlOreqvs6iY5dGG/vzcyPS40qYsPxesXdVUz/WhfjdujsNpLq
mVBJxGZEbFBnj7vq+jdOkBKemQo9h3kUwfqYVexUaMP0sUQ9cs3fRmJwmXnfQnh7CyiTrb1G7wst
mYgz4Ps4esIarV2jaPzr/jiysYK+38Vj4BIGMRQhM2t05E4LcrAROAVVuqWRqA6Ou+fUbh7XFdCk
bvRy7KqGWZ1otdrbxcdhuV0F3txX0YLW6PYzPmM2MJVC5NjHbNnVQyMkygs9LlZihsm+TN5IaRnZ
p4VBuSW/Jy5NLD5dISWA0asQqVhSf7l8EDdlNFj49bCllibOdEzTrVR7zDVYbuvbINOaAFWxC/Kc
9xQQmqNMEkyJ1xlQVAQ05rqIt4qEVZZx5aIm8Evz2P0eJFkQqmDsVMq5vQMPFF1y2PlF36j6fwh4
HvaJ8ECcUWWzm2iPbvxvLPbPK5/3ZdOiUfeM6NzVWOtp6xqI0QZL8C5gEisfClhtyKQzlRaqsgyj
Sakc12doSPqey+fucMU/ImM/P9VWpNNkGI6UH62apOuTLgpb/q+F1kwxZbnkUOrYw42hvIOYmdEz
Jk5b07M0GepD5sVj/5P3i3/1OmLqrxpZ8rFqpUnfXN+wrfTj+VqepHNJDtcy/wWKcd+rkDFf5UhY
CtMkbRonRV85BRx+ILh7HMQ8rMNLN8+OINVJjrS05MAxhsjv08rqfgeQ4j5TYTdTkIFhkXTk8QDC
XBd8fObtW9MORKexheV+odTkHOCaagRcGADvKyEr12CqalNcqrruNoZcLLoICRoOYsxC/XW+GZjL
0EZKDiyG9jkcv1/QyV89LT13B6fE1c25DgMYdcwtoJHS2nm31Y2uPh7tWmPcRz0KyincTG+Af+OU
RpLgU9XMe4s8Pcz62sS8uVKQ3VzSnjCzw1Eg7zXQhVcP0187cjthVMD5yZ6GU41blDiQitLTF5gK
Vkv04Aas3N8h6yo6oITwjb/WVXWhdOfCpH8UXq6Yp/a77x2PByYHxQqQq+sPRenZox6pVkcHUgBv
GRknKEVvHQlR2Ne/15HFXoAF40otv97D2RNn8BUZE3Jl243Ev5chGP56u2Bxl5mmN8OabWzMxtKO
hWSv10ZoUSm0NO5gma23Q5vl40Lbk2XMcxZxQk/vBCf5BswDZAdUWoPlqOtBSIQO0l3wJYUjHcxB
6JKrUmsOM1thgVRNl5a4YTAG+YrXouIMHSBmM1tVrf575Ybm6Ghr/nrbTQB+j531iS8eQcqoU8eH
BfefgHL2/dV9TKoBKbCUjTIE6gMpkG9C8YGkd5gnJizqYT0DoiUczDKcElAdChFmMA3CehItU136
EUOuHJSWcPlkzwVQp+WRZCsrK+5e3P6J3aaDUET1rAe6bKszK3yTrV7FHntUBYd+vCrVZr2WlwiB
YWHLxn2jFk8Rg0uF4xvhaMK9gJCduQcTWfKZXFEO4Lfmc51W48JDtWV0Dtnl3U188f4/ukw8drjG
UDvEfVF4dkCU6Sf1Y7qcm/+pK6gRmUx1s7q4eIbRLV/FD97cnpinbuDe3Pt90o9bQnj1VlCjVDGd
O3Ctt8ZiM6oyB3t9H0RZr2O6l2F7fhx/wf+UxCPi58xaFcSD88catvOYOfIBGhwS4uLT4/QuQ+zk
3nJq71o1k5WxGW542U9Cbr4u+6bVpcIc5RBCXY8wk0REuhNE9Xjz7vOw/gwCs7f0mjcjhVHPtjA6
A41ASXFNk3GU5FxxCO1KrpRse33YsyMaRON39u5a2MJf3ILm7fyn2l8pqWso1zBOaGlejO8/q8rM
NzsAQz6uYwSSwEOA+8gaNA1n9aH0qtLrYdbcQXHECD19zAAhoJP4vPJJWJdnQXyx5PUOm70elVUH
ibTLTa48nh/tdOvMt60jlQq9gGvcZ0oT9nk5aUrDudwkA96twkWGEx1b8ZH4YHq6K0nWyGv1uNbO
mNdo9onU7cvyotCaTC0dCSwf7l7c829K0CzONm42SvRVL0+rvkzQ7Il1/J2XeIxJvJaCeVHLFYFc
UcsnedxLodBdEtFsj3Iy855+iy0x5N+wdNu5uTgYuuO1BETNSxSHr0+WV8ETP3fkqGks9ag+kekH
b2OVEWYL2HHykObl/Tmn4tNeKpOfG75sI++DWW/Q2TbpdsIesc7jdWMXuU4lUpEtHPMJPL/wibYs
KHh3kmCbSka6dhQ9wZCU3zagohMHUdIcU7re75bMYfNjQCMNEBMZzNH/v742sk8y9JNmALKyMBgA
x9K92tsHVliPWTGhIzhIWbXzDfDINZDtMKlpb5zZ9IQ4hDiBWAhF4M/wa+9IIcDpT+aepeFnn1JB
2zsORlXKImt1vUh6SnWK+uRFoUXh2nNN29MoMvPhf0CgZUOL8YL1M10BvRO0Wom3X/LSc7wKJ2mo
UoFdrUCXqp8lasM6OmhgnV4C/eADCnz1HbezcYrEw7rFhcZCjiA3+0k/7SyspBvIrydtny5uoYgg
3zYtNyTD30KoEPxKgQH86UFSbGrfgTLPdtn9mmbapAc61QzByS8YJw8bpjDHpUdQNjknjpQaOrx5
oW+nn7hTF3Z+SW7lun6ZzYCHpUEZu3hg/PfN2DXB5lrPBBojpaFW6cTGZQ98/GmmY55zy3z5BEW2
qqwL08kQVs56GnKP+PJDeJsBKQ6GLwpyQ9F3ZErGrv3SPbzEwJvEwRrTwna8HXOMGYfWjMFi3mfp
ae/OdWNtkqv9222DR0CYfRUajm1IZry8ekg2HLZ5KkLDts5IAvL8E/6mH9MfSny1Fn7oJx+CsAYB
zuxkNtkHpsEHofuKCORgxmrdGQiWWx1dyor64ZnZ/tqHTctCg2acaiw3CxO+6vTaYC+5j2Eh7wxY
6thomZQgOmmjZg26iCsoNdzmBzAzZlmiD29LGEXgT28Bnp9xzclDCAnANayv1Ai2sbEj6gd9WVKo
U1hwK42pDhnfZ53lyI05aCWthExNf/5PXzoyaXhePA9psTGd9W+B7UBe612GuWM5OyrTo158PW0N
KKgKmdx0tvnGR2ry4a/WEmFy1ZDi7R0K1ab5f0UaAr1lrO8ZFYrmvWe8nnCxgpZpt3+Rn2ZkfvYr
mYNT9RPC3AVWeeom6zpb6MPZDpGPDTZZyhDWgTKtuMDG+hh/KEfweMBhD37D0dOv4o9F8VWTJ7lQ
NmhqiGq26GaRasXM0q7NVRNR4z1wVgwuXPB4EYGCyyf5/kmRtgxpRoqmXOhNCV9vJOq43LL1VgE3
FBx50WPBu8A7B4ycBHttbWvuPs+fR1bJHf4eo4i+HOKPbmLywEV3I2eZgPB2fvrKRGg6f8FQCzBR
bvyvAZt/R5MgPnJuluLVpKP8s6njOHnJG8YGOp8ngG4vO9nAkLmXeYohtFSEbpznG2TGMJjwwUzl
YQDaujsdGuCEvMchy6nlkqdelItJ8ynUxjbk5fp+d8+DAyk/6xdNfuSgqFPup07Hr3L9Dq2jn6sx
AR4iUZ85cawESk0Zl8jMkhdx2acbL9N95fnCr+T9D6fArTFpcmggzuyhCzuUkL4R75bnOFnGUAbr
XTdDOZJmhlVScepIi5WG4S4m/fZUENfsEirZijHPAwDS66j3qj2B/BDKmmwKkPZNzy8wWmx9accZ
uZXX1soci6VJznaJ4ZB4gfEg2s/I3wzXxQskltT7wKuaLF8ipZSchP8uRB45rY6Y9EmrY/PokkFo
FIFcFCS8zRTNbFRXpAjn6GjKvDF3SaqLCboQenS2AukU1o9f5dcCwucv10i9tj2J+7CCJPHQQVV7
Pi0aT0HkFyolAID/+1qxQdaza+MKFuJ5ptpqvOgnqhKDSU+QHmy9ozxiRtYfSeHfXPbGuH73BIgL
1DB4AvBjnrT/ToX5izPQdHhOrtXfdLcrW9DLEfNcXbwgFBxsn1OH3p7i9qearXs25mZ1QkE9+fNH
SL7IpwR5Rx4+M4SzkaZYzCSuNc2g/dxPz9iJaWRyu7OUrHcWDSBcTMAeM5utXJbR+PgMCP5sRhWZ
LR6536tj+2YyxWPoZp74NUaEyTAEA7rRKxAf1VXWRtIzdBNK7B2UTO3QKYinZGo4XoQ5Gh+SsmpI
bu2vE/r2nRSpDzcyr5sjsRZDX3FcC/U62KLHOQTgOa8Gst6CtulD6eCYCHdafoYU/xhtrQqulnut
5voC0Ua5MyOa1vTx6q643VF6FLKdbzTsiTy+YrTxNt4lS1vUN5pTHa3Tjqo1CGe3EcR5QDhXG/Aj
yUT8wE/Psmsnbh9FOvfjXmfCQiK19OxK4GCJx5DfMmvD7CcPlaigBM6UHa4i55/+cABMJ7DsYZMe
K0CBI6X+XLvDK4gjXyAbIS0LidGZNoI60b4ZEPk2X9S4VnatjkSCee6nVgNVEt2+glg/c0vujOYT
m38U6AAE49426h14G9KHzykfFfO/En7kBLXBi3FEN9+iSPJ1LfZvVPDPWD9vL6xe+MF/u2TRc/IF
z51SD5AXWLIKdKVyIBLx4wjEE6ChhD/n/VzVd4FrhHCm2Gg6eEVOd1fLH6FKFu9ji3j4X72Y0Vd8
t0RMsgdShkvDBtdelXWIDY4Dna6McQii+CsscOj2r6/FzxzuNtlqsKFkpnx3lMGHtc9JVj1zQVSN
04MtMfKIUxzLpcyLt/iJNnUAFm2mo32P0l9eQ8z6BOG87FFnzajCxhl1ioa814oCelziKJNqsHIZ
m4dy5wdxof7CrbfzJJ7qSg8tEd26YsVuoJX+Bnr1fbMvPgllA0Vm90UFNkeZlJjjVF+pN4xFdDkN
A4MxYd81OE/kDSIk6ZFugMJkFWFYongkKE1JwluLZHNywmo6lLsYVhJVtk/yitlLm7MIuAlNdZ7r
+rVG8mYdtTgEvbws0bCNOLuqgtGAPEIH49qt11/bwH4UJU0J5qH2tjz+CwWx2ZzXYXCeA7z+D10n
3JhRXjfzDnPgsJhi6rvb1Ua9qFRhVRm26giRTMzq/gL0A2W1FlOtXVbtvPA/np+lMfulb927HrzZ
0jqPab1wH13MVrhMN8mEvxwziE/pVzBBMydlmtakQH6B9NnuRCE2tgfaM4NHz/VHX4HqXeuXRZpz
166SSr226T98XyyuWQVznCkmxxvdUEtQ6DUNiR41nusor1mjIBCstSNK9putJptYP/aVCDY3rtXZ
agghTseqImpr2Eo3r5bVG90SsPLJWDt6RlDuS8oyC/3/3WiKCkzgmnDtkfI4fgagdbnDokoVq40A
iDdisgLCLsQsKWEaiTg1teduKDoM5Gn5ZBrz+z2DJEYVFmrXtbg9oKSmir09jH24qQZdjLz0tzhU
rbo0sydPYNfj5ZxTy1Slts7QOQAl/FFKaPl1C0fm0ojWdKUdfjD2oaBtICAEFJAWbrRWqzAolSI4
/reuK0bvCVBV2wc2UZ+liVUeTqwRRpg8br2aqZPaSxX8gPa2DEsWw+p0wDaurFnGiLWg1SnF1kO8
nOlNGsESrh9uJbGH1Vqkhbt8wLwizfGcIx8zDHBUfFKXlsIw4/zcXqEEWHxkAwa5T8sbSYf6Pc48
9KbLKA43asmP+95/GPXcFekS2/OQW2eFnoR0MG9RMw2rnvS3vkYBus5oi3QCSlOplfO0FD4jW62H
xzxVn3MuPMXF3GX5ZqBINP66AhRUMxP0oplcNBqt1+hm1cKazsmMi+5SbH66yLyfyBiAIVoWoyhF
Urkk4z770vLSDjbbBrjYisoNySaclSK6b1/pQM5fdPl3i6/HGQsdnU0Hc3Q3Tuc9xKsa4jSgFUvM
RXFpBQ3ML4KLpVVQg4nqIyPPcfoSeIrqxG8Blw1tzuu6+4aTP69V1JaSa1jPmak09LVrt/V4a8qb
ET9meHWVyYNPe/KZcW6rEzXw4vnDyTH5rBdWYjpyAvPWgEqDWl45q44wNHGLQ7DRaD877uTBnuVl
9/b1FSpW2+VRzwKsuqk5KO8ZPn8JkhfheOZWohxEXsx0f8SUjO4mCGFC+uqi//s0N7+HWoFma0CS
KX/qdeWjfev/cteu345opEomE4pth/TlEfDYdAOCS9NYN5bvLNsD0A12t3ZZDs9Of0QdD4USrnNt
I3P7NzJhXCUQNEFvyD0gfFhBj6dc92BpmTVKtjYQ7OOariBCQ9+B49fDaVQAO7mwymkNrRAyJ+qT
GpkN/Bwzwf9cYkjw1SbWd2UcmLR+YgVHw67l9nT0KLr2qXcUFGVBDnERhoY4ciEBwJ/duqnQq5Eu
zbDCLN4VwmtrVjWzQlCNvApwFUfPG71wNLpiRi8KhygBKU30wvy4KLwx8SPaw5E1IKL8mmZGkZr+
WLYcrMJPmznfsLOFhKN+6inYdAendxEKa3daAcNR4WUcv47C7p+hd3ss0HVhWEUHmrKhAfAysHwc
vduZhXSFTS09v0hi3cLYfY2/LKEugllT179/MtSLfn3AtZfG7DSQXdSbTfkYFq+ZgID5rbhEZimZ
fECeY4Kb8dKfSaE3eGSU0F8DxxZg7pbF982phlUjOYXbq4Atwix6GUxRFUcwQTCPhSomX7gkYuhG
w2rY2PXhBOHAOQTq+xP+qPAbDtcOpLQSIy+s1h93TsYM6/BLLY0lOv1ihsAwWmp8n3lHVPqsebSh
+BX1gG440pewy9Pn6PfgBjsKyAtmZsryYp/vs/C1yydnREiDaWpiT8wH0xpbqKlYQVjHoG0K81dA
huOY9seb2NGta0CPR5hjrcey3lsd4Cd1LEyv1/25UpNWQfAyk+8b2lo6OlHBUSinjCTndTdpQU+s
CU28ieFGrVHxg2CAztRRhkuMotFvqgixRQhf4VAK20zSFoU4/3o1BUdsHEH6pswMlKpKqDXORskz
ejDGJ72P8TI6t/kRierBJB1NLCuC4DBz5bhvSJ/TrOoh+b3gj9jQqkB4aAGv4UaVisZo10ANcXzr
A7K968/Mx4Dq4iEfoTu8P28uYiVn7O+j2lj83z4VGbh2q3BNBGainzlt2KfdafuOts4UKth/hZCJ
FI3Cqpeem/AEsJhButnV+UK+l1UovIrFriZdkL8zyg3dfUanccuqGRWRUbnysnOA4bxmJPnPNnM6
U67JuenT4Vc5QEJ4/GJdzKOYVYNJ+5Pe9N7Cpsx7PRNm/M/sT/yTihcsU6wcDgGBtpmnrgm4CvLB
uFpLfAPGMGDHdmxFPPSzC4UNWYq0btFdwls0Hx6SrDlyJv6vsklMloBNYKhn3fsBejkINQJGvjcf
r/CilBHKShW6prWQkJJZF+teK118d0Ogod7WAlJoOk9cOCO4BUiGIT5CRveMCNu1BkE1OAggOHF7
RpbY/H7zwxC9avw0AREQEiSWG4ycOABjT3ZOLKX+NUNzPEjuCuiWGwuvvSK10uhqJ32cvZykDFZt
mlw7eBEPRgJnwdKUV83cc6uM+Ql7Hacg4YxPNTsiDaUvVZ35m9pCKLYWnxFj2TZ64AfbstMuXW4v
8pAH0dqokPzU8QFSzpHFfxIGhzWiwIwz4lAYFhdMQIrq/FE/iKT2w52rHyBvpS7KimZ39DBZBA2d
mcZzB+T4bEk5RcCRNw04rSyTV3UZ9GjHidVOax4rnocdc7KoZECkp2nhCWRhtT/Zopbs6PAnXcWk
C0s0znLabsQacUuxJgcKWcmjxnddaTR9lKofAv1lu1W5WXZ1ujAWoQYO/ff8+hXrThP1aEBiiexK
iKBW/5+OsL0sZxWonh1KNF6wu2bP5DmWbtj9ysxlbRbpPBmaSxPso09qHVRb6yzXBSk83oXLC6Vu
XiwpYaJWBrUq9wjQR9DTPiH2glwopFeNLmzuI9i6GsF8qXpCvODTWqKqm/ROhrdAgfC1WFX4Oo+F
ODEf7f+wKQqgEgKGtrMIAHtqS30Jxepz4pJ8Jf7qqCbYr+++UYXbVvSD0UWSLN3YeZGj1PGmk2ng
SUUjacnUJXCePG+bFDptrnmb4WUEe0aoT25oG2J9fgz6ExIOb6qijRIYiLY1dcA9Skw2eaAkCppl
b7ofJW1xa45um1DhAf/pFbV4ttzlLm1bG3OS7HbwKh+tR5dYMZkPN+2QrzBPoAmntiVMS7Pbs39a
q1DkFNPE46zMkjjRIzbOY5XHGL4KQdW81oymhY56Uttmls4zoKAUT289NYWtiV0SD1kH3+KtW0k6
oxpdOfHz3ZYSlwSfk35GL2SUquJp65uhi3aX959Q1QzHI32l61rgoKVRS7xdkUVz0Zy6D2NbMyDB
Oomsojlf6XhBUrFkL++AaLkY+ah6qh9ZKRUWaFXYMgUXsEqHDQOU6F0ktvHzeRdjyHUx+yFClKbK
IbWk7lcTi3NNihOjR4dGMkvSCcjWiOACITQSOKzLERhS5ZweikNyMa2TIUsrTGd9gVOVQyCi9nZM
MGeuHtNABhQ01FrIM0pzwXlCc7xsfCSSaoV37ho6ziyEW2Q7tCIyvhcsPkjHxtcltzcdijhFoOhe
9oDLs5MTL4dbhu7dqp64Mz97m3RhT2Yt0eUYkmrtf4cbnbzhCadOvYMpJUvf0GPVFokWCaLGZgMs
N8Pqczx92eomLaIa/XMf5i8eXrzNn+NSY0OLYnRCmjToFSTBsyajVX5ptHbT4No5Gl04ZN/F1QNZ
d5s56kFKDvf+XvBmt1a09Nywx+28WGW7jzYMXUKONJ+nTzvvM2GBij5u3Nv1/TY5nUGZiimy0Hif
UOyyGrXcIB+zqiE1uekNFtYY0098F05U1H3F/5K+Tz0aNKrnhOpxuXWtt6qGbU10iykeYGIq3Iao
jeq3kTkuvq1OH1jm6oIb0lkg06Co6y4b1WuPuMCJdiyVPXfyiPn3WpPmvB41XJUwKpccnOCD0QiM
kn6J9DZga1Rvdje5R6LWofm7WW+FvGSWVtIizlvf4f47Crwqr+KyZ1cOgYlTwWBwh7IQVpeag1Ts
aQylnJ1zAi+KwIwQYg95k8N63uVZ84AE6TU4gbU/poyrHmVzP6hTTnt9Gd0340+6cXgfqPJ4sxib
GCEOAXq9BXZ+Ewikh7UDdXOMOyqeifD4e1mVSKN7KNsSeWvFwC6Gd7VTf5RTl6JEyLnjxvGVa9yV
NHPPPotSapeMrv28GSRxX6DruEFHxhWY2Qud6MfxqSAy5Jn3tnfJ/u0Yt4Q7UW9j5CH9cPZD9kfi
9yzkkVh1wt+grRAo08uwNBwHi7PLys4AW0MOmwoPX5rDvVZ3/8NMYop9T/BSSthPumaxAAs3vBGz
jERwj77qmah6T4g5tCfIg8X/MM7JzaHo5YAMbio40oxMIGbwpJ0SjT9lOCjKVGhKoZMvcYiRpZTz
FNgCXCpuEYJlv1iZskC7/4JF40Qfp58eCWkDWHj2tOi/lZQCwz3hKBwzuMCEsBUJii76eJ4yMIzJ
Fbm4bPaxz1mqfH9dnuvc7TkycMDd4FkcK+5ayQ+/9gldME5dugdWCQ/l7VaW0jHdshBEwc3qkdB0
xrnq9ggRXM8ZEvSeZuDM61RUWb7jMf7kXypkvgZr7DDD2cnKbkAgFDmxxl8rVoyaMZ+hOtcqLDto
B07jHuw7KfH69tfh2f3GHe9L/nOzyi0Ko0vpLhDM0mdi0jZC+CpIi66kxhQEH/MRJYVhS8X4zCYA
VXGSuUiFxRw2c4k9teF5hcDiKV6QJrVQ5KxTIxTKqTV2GRmscvaUTBIoXvVr+/pHBw6W7rmDQQ4Y
Cnrh++DSrGXyDhHEYq9NuyOmrAS+agEeQLgzqoQM9l8WzscpGIzJMjQUR+Ux42hVtU4K3igxkYDU
LlUEanRW5hyXE6ZD4TKj4yIBIWLQAq8YCPLbSo49aiAVELCo1AK3hrRg3YerOSvm25J4L7BdIlfS
Wf9FvCf/r5ajIhze8bNCSrlK4ilwZ+m79WnXDhlf7hKGePTgqrk0auk+e1l6bpvIn1YAX4DaXsDa
+hGtfYzoi9x14lkHR+NIuMtzA70GvecWwGuXZCKKo9WSxiQi0JjRAv7J4fSpS3SJqAg8UJ7G6XJC
QvibY2kx5tbIFp/eXs1XcEEGjWxe4iU0U36yXZZLrPSmEhcXAMAAMSZfsI3VRmzy06lUhaHP4OXd
5LZqu4DRxdOpvk7BPJ1G2vbcO72Dg+BK3+U1Jh01wpQoB+AXoADd79MgUlrZ2gVTY/a13LLEG/X0
48F9373IYwgmFqsRIPxdGqrOTN3IDp0LYSgE2NkedMjhM5eKK8kZjOkosrDVgOYknahyXBdwf9qz
KEL3KK3n3+0ksi4iQAvcyEL9AYwre9f/1/jEodjNwCrzcOUIJ2xgZ2VkEMHwKoNjLs2fEpFC/3K4
se+n4lDoD+LV0qysmVMKTyk+7xo+oFucRgfJfeSP6lzi+MJncrZpjy/h0EpWCtleHFQ0MCogFIUZ
ZlhT1d/PNeqcRzG+19cXVn0Le2JMxEfny7EtubFV3J2RQtiHOMHbOEInDzSJZ+fHwEgVX6vzn8xm
eHbZHBdpRFFGyPjPSM/hR+2fTkl1hz09dIQgTlV+PB3Lk0ThpqEFwHjKQjIJz4uTze9i7NCmMgdh
x724/Mi27J1D5oU1gfDs3spC0BPkVmImsq/4G5dTX2wZ1e3uIc3SvdvZMcHgIgKTE5P+3fieEZik
3bP3BgNUtyqta2MX/jp2mapkbZnjrzpBR/tQGvEf5e62SK7weZWbKbrIrmT3zEuhoz0tC2eb/NY0
N94DcGDOpcwf2A7fivRtpDA3B5uM3YF8HPrY4Sgfkzl9DFJgT7oFG8r+KcbpfHcdB8Gm7L/gT1/Y
thJbcDROPTYnT1kNGjfv15MGSmGdIvsCmt11Hi3Ks858g9+/65QHrB5xAugdGqClmGsynuV7xobf
kj+GV2q8MpVx1VNCTUutzOzeLypR3cAYquQKW6rNcKSArJReCnZCKJRwIlf6L8x1OuJ2JeGB3NTt
Y/5fF1eyiewBPHDtycmK1Ci5GHF0lyKRDcZcy3iKdT8yi5cnBZJo1UoHqmW4Zi13Pibge0/ee418
u4JYtl0SLqjIPgqmo/xHUirGmXPUj1K2T+hyBlK+N/y/81ZDgit/o2aE77XqxL5/OkcexxjZs+/s
P/AhyQLJa2+1/RXf97XguSZY+Voc7B1DM4j1TMdYHR95qL79FBZv0dYzYgExdxPyxpJU9tAhGhDT
LnqvWASQTKJ+iHK+VIaBTlb7G9L92y6K53lt5n0F+F1Qk9g9lWfH4J+zNJeH1tmujJ/cOwSbh2yV
6K8QNElkHRPwpq/xh7sQUyv7Ig8ButHtk56QMDyhCJS5lcNAbmUWSfSoszXWV0ef8ckMQZMTlpFw
OW6dg8UeXZuZcVChCxHRM7Q8sAofmQhWjYvC8KScfSVkNLJCF8YRPaSddQad7ER093F5VqJF5vwA
w7Axn9/KpaPkeiEFQe4gmyR4YOO1c1uFTovlFASVVwFCn8w4W7GHg3P+wU60OWEQG6LhfNmeU7XL
+h+Wk+mSyYBkw/ls8skS51dT8267HgcBeNKZ4H9iBrZCRFSq7XkEL/VVlW1K2SSGtRZxl0qOy2Km
zuCLhhg4+gjAWfr3tnncGQ1rdwPUTIHO59AxIM+0BXp5gI5ARIMvTeUx0u6Law78lRXVu3TVsiZg
Ktg3s9Th2laM+BYDWU+vumC2q0cvAnPAZY9KPvkJAoWt0hDpIYLiMcKmq+I1KofH6OZwXNKY5yNh
HM7S/FZxYTjFw+DvehtnkN+C36HB9KaELIyRoktD/Chu2QHZdNpOrvflMbAuECy6oBKRZNGzgEZx
A7kQan7ST89plDR1T8UYewuMUbYiqSyKkYsI6RgE32W7Q+FYvq+NNpE0Pd/L+5JKNXSGEkR/+B29
U88L83DgySoTBRrClS9M48cAJZjK+WJVHyn9lwXOTiMzr9CcBVSaWcuQHxBanRDSPHq3Wula/MnZ
MreQ8k9USVgiSUNqCwN1EMLHbHmGGP1y0OgupKZ9UfkL7q7QPIwqsGsPbNKORg6iOuCO64H8wOFN
Inse42zif/tkowRxWvJwQXXCvTllvFZOX5RVPsQo5iV3lnuoFrZOc12PKkW2ER8e5S9dHbWhh9OT
teEM3PpnQKASd6OhnbcF9buYyLp43ruPC38JygHHz4jMN+jwqOIsm5DE5Q1bPsI1FTWaOd2L2srK
OrojedKp+zId3Cy1uwl+HVxaN+E04tYtKAh1YuLd7FVJuU2sNMQC2jcYCJAELCLyj02DIWN5PyDd
t9OORGboFA5XjXGCUrKYBIN/wZ/qbroStY7srBXezSeUsmBhyBMxyBtibtme0E/yn0s95aFB7VCS
qGvX/xbgmZutVVZiQyZKA4UgtedDIB3qqlRYUKSdv5xvm0ohwxhMBWtYRxu7zqU4TulzN6SqC05f
vuvRFg7eR12e/LX1FHtqFesqvugrHiMb/Sk39EbA5g3cLgK6/tvgS8pBSPH5JTRi7NWk0uAWHs21
dy3n62rjLQgvNEJ6AyV2IHq7x/oP6OTvLxVPKpAXxgegPiJgf6UgMrL6JJ5WiIuoWIMICjMyXA1v
g5z26w/Nz3q+3qvvrZlT7S0JKcubbvJZK3ts++OoSh4ux9wSlZ2esgXlv3dM5Rs2N9RPACd7M3Eq
k5BhiUFHoRSMzehFh5jZuRXrg9Ychl279R2S4j9AJod/jarJwUDKDdEZiKN7TQQyUC0UM6CMe9FT
mGjzSYtmmGcgK7bthQ6nTrLK+VE3ocNyByjRA+jBKozU6DTN26bs9emTk2C2EQB0qHRQ9G/qXI+I
Cwzv+doPiYmcT8781pHu0JqZQTNc+ejD5Etm7xa5Db8NF390fzDDJA3XstN4Rfvh5H/4WDPp4+eo
j9MYHPWblM6+Ymp9IZTmM4UYee3nu68DKqNnQJT2F0qoGJp4W1sAOXoRWQNEmrx7KlPXU/XOqkJY
4RLwc4rfVL/4g22UsPgEukFMJHqqnE2MABwBmB1Jn04GBIKB/gDHlwpdkfSBrSGSvFGx2tC/X2Xo
jIKlhXolt7sZgywF8mHzFZ6e1j2/Wzq6Ex2X5Iw2ghBmZdU3sHw7E1eeTNMNRQCykRHUPIHiW91H
TXFMn7O2Rl+GFjEP7QQRNdT4HQc7yfzMMIPw40+JSebxUtWS6YVHdXdXiIyDN3sqhmgTk+P3IIoY
rc7zNWSJEZeSpVeZwWae30bIUiwVTerFiNbDgKTQfYqyOYA8o8GHsL6P2a8s9Zb0NEAsuUZr4HqT
Ihxx/Nbn5TPpvNUkeTJ9WbTuSmK7Sj26i+0jSVtwTgd5Rm0alO6plUjD0u0Ymt29l7kZ7gXyKhOd
jdlQkdgYwEZg11n+jB+vW2kzFCDkku0R67U1TfY6p3CkB4uhAzaiv12iNjXVOTp29kWv6i0qy9yn
2+9MZ8Gxp+n7XGUSs24ozgct5avLfoexkNhMMG4DRKVW2L39D8/ZYsG+xecyDLvprSWZJ0FFezTE
sN7p733ylLBrM0AIzbWkduR6kRsqAHhJfmGZwtlraPpTZkTKLGXnQbHXZ/jvvOMxrLa1c3QL0D1f
UT7tC+5tXVmli+BuuiYkkPQo0cLF46VOrqOEqHV8FkYeLFPSfgOKSkDxNAqOCYAHof9VXyJbMiAU
BcUazAMW1/oBfl6Sdaiu091kWftSIZVDV4AmIjadT0blZdEqRu7KEx0AIh1mwxR3RjkuvrUHfIoA
2Gu7+n5XcGS03NLmmQPSlhlorYldg2Iy9LtUPK6FicStin6gQJwVAUfdvgmYp0yA+pruRARUIWV5
57QNfOGB5i0xtWlNLE/4P7gbhuXNcuNt/CYTlQ2PtEwZ0+IH8GcFKhnYlP4M8y9WdeKFBy0W9LpY
WadIcErlfN4bPbN3dZjbf7/KTGjuXwieY3Dv/rJDW17CZjS2uFGh3LBMHthKFv4EsLRchzhoVCHd
nLw55Ccc689ONHOutym549HjvZEmXjtDvJkAwvYLDCyuoLxvKTHjStp5xyJzIG8DuZ5pltGZstjS
xi28WLEdUBJXCSqBk0Ufg3s/gmBojO+BGng4zjLBEc7qF/QSFcALDf6162p+NJWB/ioxxcRoyd0/
vrR6dwjBHeYNfkmVBHhoL0dyO/W6YvESZjDJWGry00KIJm6ivVYlMZZwDdja0mvIHXcqOphr5hfE
FFYvNPRYLnVEv//otPiCj1l/cmpxEceBSlEDS8FFeALprkL+s7p1Y1lEUUeSxFmgTBTP7KnBitQ5
jvFVEZwDR1uPQO/2SJ1J0CXmlkkrEKp0/1m9pdtHPbFWrB8FkiL12uEU8C5NQTHbEer4qkOSvJnD
dAoINmb+oOonVggstuEcNZ4G62DVER8hiWGwD/xbiGAz9CZng3GC5uM+0APeyLh5vpogmLTX0BLq
3XXw3mmB7Q9VrPwi3ot/VC8EAdfvzJG2kILZ7NAee3uTYl43dc1FnQGCx9VLFBhsIX3YLGbI50Wu
nTCAtRFfaPUwJn6ato2338BdkiYtTXunntt6/jwg1YUU/1HpUjnjofe0K2WjsfR8gV3RMBaAeUeD
YCN4UE/SHl0NSmMHuShZjo/Qj/66nvnAOrHOV1JrRrNtcP/e+M2B9d2UaLy7DE727PC20zGL9ozN
uei21l+nAT69uQTs0TYKljPYVsFkbNcFA+Ae3bWtTcvOx88kS8QoKYQgxE1TLFmhiRusXabdKOZx
fx90zfOjYVG2JBdMVBL7e60ayGswjqO4XD8M5mGzF9vzxDZNLwPFx3+uPoFMRgrDWBSB/zYRpyw0
OQfxm1mtpi330tsAIKafeiyQxvjQi4/TjEMASaR7g/po1KneDQact93d944A8eG3g2Er7tmMPz7T
iLeIl/7It9m2+ACosnNyEs56Xoz2OWrrc4+PqAzqFMshpgerdVPKAU2dJzggdR5kSxtJiC1+wiyR
8U9E2P32PbUfo55UlplFI8Ryi5lw0VMlVUQ6mJqDrj2TgpmjQ985HfSO02JTxZRqb7iMbxhmaPeX
ikXEUcJEp+JXQ2cdYMIXy2QKMwSaGBWwpxuqcYjQVVKM1Lt/FiB+MuUHWU7uXZOWG88fJ9Sjc9rt
gd2dGNdQvCSLMJ6RKDW6ctjaPRb/0mRjWYXsSmZ1FcBfA1JzZaItnFmLvqhULG7rHrzNLO3T+VAu
rvfzV+Bw6KY/UDiBm8kvFmQBmBZqsqM2z43LqfvXiFAL5fUcH3uCDncvG/0Nba8orZ4wlymL90fr
oFfd2ybUwGSjFNfnR15TiNW2JOD+TZx9v19j9riW3GMfut5P/0CwJAr9Y1eLdyopv50WPI+A3naN
vAPJVWh0TX8DUkr+UxjZwp6SuJPJS5I0ffCyt4Yyj7L1rlcOzrx7whSnykqCwdugHc2bnjkPaU/r
tkiIenPot571dPJW+pA+dx78Pmfg6FszfYiGX4Ki/yeKp/6xksddIJAyOlKWzZD4+pPrzy42GMsU
d/k9Tgw5L6kWU7SXoNf66cdAivhI+/h+XAbdta+xkuvVJ/CVo45H/uiVOzb75t/eHSkxdJTKqKrA
WuFx3xX3LL9r3LtRH0TB7r8b30c2su/bEpj3OdAt1gg1VnmsZPUi6Mx0a2kGiftoQyJ6k0+89sD6
P9pXwNm9TgZ2tr+VGyQ3SQxE6ivOU+Zcc3vrU1aKi78AytWYFgwVvHxB2H9UW+OU+8OoBcsC5lsK
1tjeRt6umGUYxJ4AQHbvHgWEOTDKi08Zb/TYHq1Ab6fQHpSqvWK5T+C10/w+Wui3EiMXL9fz1Tmx
qAGP7TD84XmEzPFpbSlMYgHSTI8rhon3cc2eJKUuunG4vJ4SBzTU8FiT10jqv/Iy80WgougzTu1H
ZlKlUPVqgV0BEElFbdT71L+v3CNcPppfvgN0iV33PnkIARiHfEpl1nuZV0kVpBWJrJ8FImUX+vZ1
qN3AbG60TMhxPLeFV71ycBoWB7SgZFEsP/EJHFd8VrBNY3ZvIS2zwEiPjXPC11EFDUeJ8rfhpFFg
xpvlqCX2ttSufyAuQbBVFDUCGr8m4ItxRM0h/RijYOE+K7eIjsK/VCvi4RlZ6ISBSWjslyEFnVtx
4Y8AgWB+ONnf4q3VZb9noGnIUEt78aeLg2Ga8mbNtjklNfwyRFTA6D6GtMt399B97TMGQY5GoasE
KO1xguN68buGdnW5nqfoEmn6k9InAj+NlbT4+bedgVXQoUy5EIMZB3j40TPLaCxfydW/mbpbds+6
EryonWUBJNnVnhmupOIcb77mCr7/yXC4lKO1DUpNZeTJFRu52HwP1sV6ZOiK5WxaxxMOHsxAycR6
nzFfRSPtCME/7EX38WnQr9YZL3zMrKmAT+b843c7SWqfm5+Gj/GEVz6/lQGO4tZe9JX70lMYULw+
aknPBGxw24qnf00qnujWJ27AMlCtFYjv7lkCojsVbeLL2+mrw4nUYDmeT7W2ziqz8RA4EcWrWSUg
65MERaKHVqAKVf/oahhY9TF9YM3RYJytYSsbSYi5DLTM5VWlb5OBS+TglMs9rOOjg9h0rGysbQS0
W5TD9rlXvYMZFzd4jiEndwPiuRB7TQst4E28RxYmfZ5We/Xodve2M996l6unZnqB1kz3LT1ZX48f
ZDT/yJIeAsISnyw5vT3SVfQVrpXl5UNU7xms5WAyLM0rQ1+N1zHiQu8XRJMawuwkhxuMPRcZUs8U
yclMfPK/HVgr6nyM57vOIjFoWPl7mGvVTpI6vRpWj8IqYLWmD7ehGzQi13lxau34CdeA19cY1nYG
WiSdkvTL9bSTCfI/VOwWH0QSXGDGUllWF6RZIhdV4sM4xMR7Weh9j6FXGFM9A152AtdCpC+M66Qf
0/roALE/yDIXfINkas4KAc1XRHTwXusFgH1lnL0OxB6YoCkQftEi1pK8BKZsDsAMnRBUzzcRnQJi
b7rHiAx3a+S0IiaMCHjUX9VzYB4eJTdvuCw7/fcka5PtSrH4XwWW/3+HTj+30GC6tPKj+mxuhE6O
mEZ/HN5W6/cPFhy98Xnf+3rnwENPLbSvwlc6HTK3VpKpI+I5KwghSkUwjjgsAo5vv5+qBD0qxxL6
XG0duTqBG8ZrbjL7w30IzUfJrzM05uk8s6nipmcwqqY/oJ6H4EAiNzsRe9YY49VTaLi26WwvmIgy
6fy/IVdd+r6sh+p3dW2WdOQlf7JSOAGUOIZUG+L93rXYkcR8f0V+fg0g7qVv/bnrBSeGMCep+nqA
jrk3wSsLzrOavyPZ9eYcsgEktNnTrCAMDalv0z8ZyNc2dkqjVNLDRx6BCDWYaPOZ4haHPv2V4trG
qsf+m6R/wn8Y24gjgZxfkvXW9Me6wE2O+aZQ7xGo37Z1J8nXXn7fsuy0Nb0h/igojbBTyqTG2PjZ
51BOU5qVU5D9c6HeHk/6r1QjgibfvZElL+n+mztCeVVgoHDwnENTt6C56UVrxufBnsQtDqbfyeLJ
4OpUjmlxlCTeaMOqCj5ZFbEKyiHos+w61Ai0Lv0CQqOf/IUZlC0FfjTbg7pls7CvU/uGE5G57Ieg
dMcIo9XVOx8c4iPFcc/dRld3Es8NL0sS0UH6FIKY6II10poEfgvn8qOmXgtDtmEOWdTKJxghQHSy
IS8cQ6rR6c5WPDiRNohsPIDst2pMVuI1pemJjj7u2I72tqmQfmCO8XqqeqKrphF1TQPVBiAwmock
9k5qgHzqPoJ+oIBploSCXfNMyZcFMYVSw5xjTvZEvphvphvgWoOzLdOF+nge7KJ/7w75tEuDEnaW
OkrGp/+N0ZP5EwGe8jFj9KTWztMBOP+ix1wd6eVV697AdIjqbvPw7aznimHQEYwNm12Le9gmg7jd
9RsPZ0IbtrEB2Rp1btbPZg5nwhQNx5yzCqWddNvwaHHD3HfLrvmSyl/y/2TS7jUv6V2psRnLllUl
6C9RC26XLr3wdjPKy8pQu3u1YXnPzEMQQcGrFircgmBI8LTpa5Vo9Hn99YcwGVZo9Am+TLFwMQft
5/44LWKlzyAiFVN67PEItRVT7asN+7O6QmlT0V9N8MbGjYyxIQguyPP4g5t14n50nIgoCroefluK
biVL3DPMknCuyJ4Tq5rlJx8tR7QJ/Q0frvGPUfNR5BGt5BPqCGb7Z8WOPtpxpfCz7XYrXxruU0ru
KVqD9slwhWm8N7ngC0JkpMURlr/FHV77Z6VHcoE8H1YzqTNIe1Q3FdMmEBFcXxsBLFDtnKCF5FGk
RezQ0Gncl0r8iSvDkUT0eovF0CYZFedd5yT0IOjPvgQLVSXcD2sKQsWkOn1+3AcwmnbdNkJOtL9T
fu2y1C+LQX1N9MHy353xFO60vi8qYNxqbh3//ZMilVtKpr/Ez99AdXJrU9aYPoa1t8nJqBUr8GaZ
dEkvPSXLMpATK/vBYtPLo7xGbfBvLesdzjT255tG7iZcdSFjXoona9qpEq01UcuidYJMVQFhMfI2
GA91BpJTNrtWkfA7yvzyJGw/NxG7ouu+SBsJeiQLRbUPQU+kwEv1cqZjIfOoRkabn44u5tlhYzRB
jYthsYv1+0sqYIa3+97libs4YBsOkP0bJNxnaQlavRw/Bl+ZgA/HsZPzM3LJ7KzJjKtb6zzzB03S
jPQmjsA+yw5150HlLO5HqZtLNomSnQJRqBu1RsT1ugL/ZAu1Uh5gbQQumCGkOXy9kHUr1H8bzw0o
T3owueYolrOwecFMsqsDWwzyxhVbNSxUJcD4SwJOc5YdkLgefGmn6BzP6YtWZ6kWZTjaGm3ItlKy
FUoY1nuvSQ2k0OoLs0EFac6XlTEvhCwOdYb1koTlgScXd/ObYobOv2Fkhd/RmqLm7t9EfX1+xjKX
u1EJj5R8ZQvQXh0hHjmvxSj/S1fexCtrjGOQFr2wcpX74vpb8Dytxw4XNBqa3UD7VKuf6SvkCNPo
+jVcGQEHhRuU/nod4mH79YWXCMp1ai7yhCfJSMPxDD1HI3wv5PFAVrrHaVoRyovtaiaQqEe450Ra
8HcVQgzf7Us3T7fvQ0WegWl/8CCIwQ+fJqy8kzxKJXVkVIcw9QuPl5oBdnTzBiwJrYXRC1z+Rbio
ZCT6UpU5LDH2amQMjDx8fGVgNkFnRDo2eP1yvO2AkX2wjcDEcLPnYYwolnycHnEkDzO3jh4JJwpt
YNiXbPzcIyQ+RDs9yVtRWsAKhq6K0mJ2k6lGlT7Tle2w4XHr4M85LjyhiaUhK2J65AjXU/K1xUij
hgfRDDYbGerX6WA8Vd7/p3dZUL7HWOrNVxQUFj4VU6uxizVJHxeBsqw1KfPl0C09kEvniXy9RvjE
qENRIaOnR/QrjSm5OKEXja0I+WixK3wmxbNIMN/e3g+dgI8nEuGiDS/SimvEKQKXkH1eiY6xYc1T
UX+tDgRZX7Lrvx5eKaNIryVnRvdoBz+ee0TIV2lGLdOJuDEwKgBeRcsL3d7g3S4JBoIDBsOD+wW6
JpR3g3GdmtMbn4sojjDI8vNV6PO7aKjQucx+U0n13e/lZ5a+YvVWiZhF8MYX6+vahDosDTY6Dgxe
L0BJ6WCc50Kz5fIHVGXP9NycXX64VhZzdKXPZlX95LuXfQ5/zSLUyHRKijomXWPK9H3dRKwxXNQu
mFxIgO4BvEMU5D7uo8KbcG0Us4cy6TshRLnkCKjanwWcEPtXbp2OG4dbab05NkmS0YmIBaUyrXFs
qMRF4H0fbnc5+tQEyW2+FaR5/xEbfWN51WIici9AAsULJSu583EfMZry3fgEmHBHeg1h24gDbg4y
hdjLfJUTbvw03Hv3IdHDgcxMWaAavTHjye8A7McMO4+XzhTyTHo9R/LhD+puoT0HnxlWz5jid8sG
kos+Fm7jeLqlSKmZTSkE+YFOJQ2t5RGQk58FW9x0n/NWWtNYhEarjsqUEyyXD8pysC/iQZ6LVuoe
iBJXbVvTYaAd9nHcPdBjyh6YDThbe774bk0KX/x83L6wJ4VRWmy48Ft/vWxv0l7oDAGLGhCVh/h9
+uNi0TjmgaQ7pWlZo7GYAGBFDprri2HEf637DWxnprGNgQRqbFTNCWxOnkwQ4xTAFnaspStQ1yQ5
T76ERARe5rFWuu/yDdi8AVz52bOGCk8hz3oSxBhQMoe85F1CFJLUuKkfR0oivshfkl5GqaiKlUL8
R053xEl4XdjdoimcoPvEKiVN4slw6C3arvGbAx8ejmVJB+Cc42S41+wt0Y3M4uGs7HCRuyW1o6Zl
xaqnrMOsTIk9OZKR55AzUe2J3NcRHlkyWXgRvtKaCEvv9Z+klamdtohPERm0I9Z0NubP9w1+MLJI
mjhF7vF1LtCUwyWzPyPWVkaynJ8AI8RaxKZEgomZuFeqxvMLA9MTVDIgrk3wTZAFuUbnV2SnK4Mu
L9KLqJC8AvNCHGzVzJNSj5TvSqqX15NjjhKxP9dXGjLVukwUorL1AeyVEYvMZTVnE3tL0b3CL2dk
6c4bEg3VVeU7xv08qCqm5vuThqezE6a3WUzg2Td9b55rr+iHegICHppoVzK/9fkSVUgZz8Cr3uXw
3blRJUA4TkOImD6GIdAV+uPZ84YAM1YFXPtv86knl1mceDsxlExqODpxW9j9RJLbzNGE+eoZmUxr
JCj/F+e+bmFn1xp9ovXqAFajdde7ibAoCJhbwAqf9pQYoyr/kX9W+Hoank+nAYPNB1wNNZ7TlEa2
ZESqU/8PPExwHPpqcCGyPDm4mAridwuYJE8xuJ5CXQ1P9EbxEOcIG+IE/1kD9+u3hrjWq7HNhr2t
9g6jtSmCgSmc2Da0ucaz5DbeANuPPRgr+aa9Q1/XDgG0JRTLvCdNQhF1OYrNDqI1GDqNm6P8DmUK
Ivo/8e2icrq+ctM34MCYAyvXx1ru6jQmWDj10mbGpZfaYCyki6hzvilURrmVLlI3rdjhvfRIm9dO
jp0zVHSENdyLz0nfXvf03e+hbleDdk3kFPm14iK2zAfvqF8YXQKhCVN+GlPumo00QM8gZ548KdIj
A5BX5WhqY4YFffn1w23CEC5RkDrpb+zZwXAaR9W+7eN5kyBVg2fC8rLAcYkclVY9yYOjwmjiDZ2F
rxUDExJ+1dk+UHZPDJLy/kYOp6aV1bMjaWEgXxPyAZd/vZ+jw7rdjeW/a6gm1BodzqkcBpEOUu/v
NyBtZlydJlCzqzQNIAcZoIcanJCC+5Oy1pTW+lmGeI9Kt4N7t4mblis72f3XlQGCBGi6XzE3LZ1R
VN1EJSaQtsuHB94pnklSOwoGj3RQyKcQRgZqJqkySr3fk1fxj92HLo70m1lnN7C+qL9YNGPz8FNb
6cGH2AIhW0UJeoiAnxDVIxwtqQ8qPlel2slc1XEXp6C+Dbm/ZKs+WJbrpR1yQzIlPwaTbY/w8a3u
453QIXxgJmpOfAqOVDdCUUfXFRILSI+oaria2Uj0RJjBfN5Xv6EIeyXXT3iuwOHmS3uMM3WQECcT
DRV6zoE1ZvM9ByTS2kwBm95LkFWwfmnYcC/vsO3HsVDTG4AwOMg6IFUa1AuhFyh6VELtMkKcTXTq
Olb6MnnJFp2lliSM4Hak790EnVQi/dH/lwq8U2FMeqNtX147w2ZRfw+wlHAlbhRE/eCg88CYQjW6
KE/ds8rC/VO8i5eAoz5LY41iEfCGlfgrQfcpOVlGB3FzXqfKnKwHgAXASsvyJfD4l6PfULfheDo+
D/gJJSNdyFykTPlv27qJo2C5yehOqG+YgGJTLnSZKVTbRz/v219iBS0ijVmr/Yy9+bwKc4rcvL3Y
CEUOZdUbDFXqOt+nzCMWcANIY1F9BvGl9DD+lZFdkEObHPjWdMTd/N4IRPEDOn7ANIPrbmWWgJr3
toD/f3aTw7ByiA2WgleWdvZdGvR+VIMXbU++y1Dffex/wxJtX4s5+YPUZq9D17nvh9XCwKP+KmYw
jfwrxZkEOMfdVMe6U4Z+jJ2f0g9c6YYC4/k10Rjgs1uGJjswWkSuordICj0nLdy6FeFR5hCpMnq1
v1LiJbc7g2vk1G5FxFVCwd5JthsTOtL397Un1b/mA7XPOM7pUuxCy6mfN05jFkyvS+mIfZaex6ye
/w0WVStTg2L8nFv0eiphq8d5VXC6+46EklwkM/3+wBMM43hTYqjRYOas4daMbnU/WVY3pBtVW/4v
ALeIB4U85wzyq7AWQ0mOQdWRHFdRxo04L9VoWz1osrx/oHn+uWw/o8l9icpnXMtxAYwNPWT62f3G
qyMnp/1DtvWKuenqSo9niHPhc/UxEkSz0cIi56edJCbEHuTKYxrgCC3Ac80LsrOvPrQWQRoqXoZG
Rww8sO1tYl/+jaR0uoYr9p/o1ypOsElrxc2qrD2hlc+MrRNKvlxBq0o1hdoLLkSUdC3kDbnRHRXd
9oe0UWH6c0D991hGSKJZepQvs32mSlcBb/5QSEjR9BwKgvtsKdoVHAkAPx4RFALFiTRbJMoaxAkA
4khqbiXxw/9bAZq/xYRv6cruP4aQyS2QgCMq642GxPLeB+ii/ymHgRmeETzSD6GhbBIA4XHY54dQ
ICfq77V3Iam1GuHVXdd7P6QT5MYBUw3zSySir7K/8kvyOuepzHaD3YZWObXYzKd9nSCmTdjYJoVi
glgpUxgRJ9IGCX0+7uITY63eB4yPDl8fuNkBLiFm5WpDoEkkD1FibGivwX/f0SmvSIcvwduyWJ/y
CQAtHEkoleBfwP18MedxeDymHF3vE3WJ++Oo65d3eZS6OyNOBvRtKBlejxBmIqD/RiY8Ws7t6YmS
V5cnnEep9/b0J+04maiZQFlzWp6lFjsSU85otegt0BPMFPztrAUie1k0pQrv30fFnNeMTXPMpLg0
2BBV8KNxe6sjMaIlef+GgWFCM91C4oVymukf+hyxUBBah69G39NS3pzSctEcu5LRQA2fuUPQ54mg
70nyR8a2XOPt57rT0Nvw0Gr42+GY8yrdCveSfKfn5azRBd/t638xHwqdo9myksPiIhEWZH0lWd5X
v9vOfesmXhSyvA78+Dw9GSHnCmUq8WFyf3xaPWatO9V5BaeKwvwX+a++eNz8UFoIAUmJC9oAaiC9
0TSs0sf8wOHHj/BtWBXLDQx3IEtkAJk7sZRJaEm1geNbg0lObtm3PTljo89nLbPdf1q7VUhfk77q
qfTUrTnEp1lcl+tJ20CXgUpRpDEGP40Us75ui7qrCzy1h/HhVac334bvXM0q5spCXXJnLub1y04Y
lOg7tf1jmh/D9tZ/YmPrJmJywZ8rqlVY+HyoIhycuy2BExSXspC4yM+KAOAZW3RlGXHM4FvCD66y
rO+O8YkigA5/1FUGUYNYh2GKYl6+bTh0rF+Le32U+hmtfYPUZ5OBSTQxFIvmPPsTRWgApbjfpjAJ
JWjnK9zp2u7WB6prYjOGiH9SUnZ69obRrZxoKsWGwUGpkdeybi1oWK+XD59M+WfmZWVWf8+XtO/P
RW8rnWaWCfIJyEohIaU0X+9ViH294Uf49/D0XTXlZnFhF87anwoomU3fgctBEA4/1ibeCiW41+U/
LMDRbSUZKoJ/581jxUxKKfS7jcfwi/eAVjtG3ZSIq5v6dOOXVe83dp2bKbqVzPRHl6k39KB0mSR2
bpcMwcZ2oboekftxgsAvXJcrYgufhlCBS0vs9W/5R8w4YPbYf3yqF21cCi9c2IoR4+XpROHBoy4k
R9LAgw3JrZuaCrdUhfMfmtuKnOtiQKNMOEhYi8ijhaAyCMWcw5f+x4TP1mBR/PRjHi6Q+r+tzdqL
iaaGdwflV+yARHLUJUbRDqquB9oIqSZH3oPKdU8WfEvEoQYg6dEjz3TPImYQOv8h+N1a7I5M4sLi
uT/66oSun4v1dNY47RkKBljfsYfWJICDrtW1lDgGSQnr4I0aRIxTkCxyWp5dkrRVkm0KrJteSoZE
70RYM9uceIFkSTlPua7iOFTOnyssqwljAIPsWY9HEOejVd8qs4VZsB8yGPIVetcEURQ3iB2j5sRy
4an8q0zmvoYrr/gN/RzyJ0I1f+zKTbgfMnRMcM7/OfgeZfyJ8/1Bv9z63p7SqGUk3A8KWmooGGsw
NOZJ5tYEoCWgoneln54WWEtDp4vwqskoQSuAxQv4oDyQqYjiQRaz0Too7YVX+EnE7v5+swYxd3x+
k13SrvoSGEr2ZxpVzjsdTinjDe+ZIaNuRb0s7SNcFo6N8nReUtwkHufdGk9tQtb05vsMRwIYtHuw
n6IccBk/tzg4f/bwNxd/L6PC6Vm+sW5tI+2xKe6jpeSedSTeXRsQxMq0rYX0iIQNCdygh25sDOn9
blqBzx4Z/tn/f8JlvAF/snMzfZFWb8E/86baJxtMB8P5WVe3CHz1QvbnOPEg7YO4bei7Limaq9Ql
IpNHp6inMDSgMs6m9/18RaLX93jQrJWBGnO30JvRPc3niy2OtQqiqQBKwwwLiBJ4Mnbuq9CiGcRq
byO/5H0a26GH4g1WqmFYcPbTWPqDyW5YXnWOleIReaoGKJZUf6U8QOD+UiADIe7w2b7oz5PAFCNM
Mm5yyKWJRO09JCQ7CTqa5hDp3jRfahPQXbUUbW3O4LyLMAvE+jNlE2dTgnsvLQR1kxzDE6gJ3UbK
nVRyq8SNo5MAySBt4GK+NHis3oZjsmfj2Z2aCimvbfIvt46AbAUKn7oXMPre/r6gE5L3QaiESve/
w3E1y07PrNY/PNqhSl0tfoEA1vAOnV17OxfaXQ941dzC4NJFb3p81Z2TiUsyZLdqL60PWOSQUwqd
OoA34vFb2zCPfbewrDPGA08XIL6u1A8YrD4aBSWQNIkfdNk4tEJgw9lcdojjc/YNj+4k3emLBUB5
+QTLBotMInkSHVrt5kkohXhwrPQpEJbk8BvBenaOYYHhqvtzS457xg6cuX34OYNdMGX+CEHanen8
lRHXzAXiW2Xpe8vJJvKdzPMf+Msw0+TUmnpr9a9vMvvL9oZteItkeT81API088zoWn1vH4BE7wRp
Onby0x1HUshRJNzFE/3RyM8VwiG86vIDd0XnQr6arMIX2vP1TDDPTP0csmJljSxnVHk8wgCWgt0C
5jgfvhVrZlRhmtsMl0NFwRRolUp6RXMu99N1/w+k6Iy1CtRMYZm24F4geU+ElaeRd1DgwaPc9nDp
6PjBZrOSINkYKgd1xZDb19E5vo25NvcVSqraJmcX9ykf2+/JwFvS/XAtVwKLOaWIPhvvoAqq0jt3
OPTZby1JygWlQTwqPYi/EgItGWqtXkdzsvSsjrATM4AU+uziyeXWN9yX1bltRnYxLcKr/GBl0HE9
S9yqriIYsT2M8H4CcaVVSdacZlP1yiLn1HQa/vTHGyyc2YePwX9cD0oeeFSA+YQF8EyvzSOkaNQG
X/7bT5RxREAiwxRhh+6/rIM5ATlTxpI8uXeNU2L+r8BEI+mwX1W8PalQiguHTIUMO91+uGgLxHqU
uf9OVoXB+DOsxQjQE9kODEr7GP4wQ/zdIPZ/hlQ0czHWozuv+O1I9bnjxx9VJoTE4AQOstW0UTdh
s6rbwIf8an4OKqOeUBjSW3/WEe59lq6gIhEaMywNL9pfKwGPD+vEdgLdQDL4XKCR0P425wx/9lGI
t50wEkZba1N6TxdmbyzT1q9m9RCvjg62LZ2OaExWKfJdP3PGEBD/ObP0d3dpVc0L3TlR1OfMjDqp
UXQ+GRocYH2G9Q5YmC18UvVVSRsZyQyMEwpTIi++i9rONUApazRsfPuUDgXsYjHcUSM6WrhHs3JM
MPaCuzF8tBbJClzphsH8bD/0rSvId1f/b2WzXGRXq89la5ZUO1h6MGFS2+c2VsiYYHbkipaF5OhG
ACUwhixA8BDCYkS/x5mvXPrrnUMOhKHsIDlRPjQOTadGsj4XWVTOy3ROUQ72KpyyFN9UP9Vle8uj
ZoqK8MYfCxLrg9Wl/pLkjs+cEenyDNU6/TCGN6+vAQXAoD7t2IsS9iVMdB0/F96fGMR4t4TJcNtx
xs/aF7bk+CGM672PRcHOusCteRbmxwfvG1BMvilGts0gge5cffsKBrHjpsJ/B448/d8H0+ulJxX+
5J/pdhzOdHs0V7xY9zhMcMY0nACuyo91ZACawwt1ACg8/OzFHodnDwk2FTkTBe3HdC03+k++ic+l
IQH0DLpYcML2l9cR58syP+0wNJtMnOzFRSu3lbdAikC2o2AEqxSaBlBntKfDrVC7mtMWVOVPD8Zd
UnSQM2+RnhB3BW6d0XxqmWeDB3FOzj4pfMM3ogidskt5N3JY92/jG6loTpUmy+ldw20neQzFxnF1
z/knJZAJKYsA4RUXE8sVjyYovktBAkshyc6t12KDbZrVTo6xCtFxPqC3/wa7ctmy4HE7pD1/ldb2
FmuJx3gxECdN2YMoF8MYwL6kcpmoTBRHBCBlQLBJo1ffQNQja2gG+YvhcXfI1yp2yiQ72c3Z7rVP
PjXY2AWyq1G6iwz5KDcuhzcSaNr3uTc+i4BiQmWCJ8xOPT5bLUiInewtPpJY6HhU/WTt1WV5eUAX
5aKlwFwMyfCQwj5kVICUG5jFlXC7vyj3ZazCVN58drgifp6qh6dte/vBNlD02TtNz1Km1EvfZAwT
NSaRgH07hVahe093WMj4tQhuk5lK6PNzOJxXklOd2qmdApzZU5cgQPjD78cTKspcxWSPYTV7d0Pq
+AwUGo2cp18o510zipkMMHzP9nlQRWdXe9DxzU4NdPuibyAbcXnsWLsc6mErJS16lkstXVqjyRYK
aW29yvBkBvPb4IeHLgnNb+T06gw83Cywoi4zbIH+PiNaGAWHRG4+RzYAIGcvR6Yj/vboUJ1EUlcd
MUMHJKpy17LsPbSYwpysz8RrNC9TSJKXav+10P22vMl0PpX8lvLgJ/+m9hp/Fp8Shlb9EAC88ALk
U6D4QA2/ZlBKfXZ25ooO4To9Y8or2z7gqUHR9lpBd0Y05Rvu3pDtUZYy2CgsMxP86w/5xIPDRZ8F
OlhFdKQwNi1dubCJeUvlAz9mOPZd5NcTA58tB0KhLh0FHjEf34eAJQAWduFoRt3MgDdFCANogGn4
raFNR9lp0Q7toGO5fFlF4yFRgMXvJOHyOdIJsJfi6D2RXNLqfpLU/ywU+FMOYvcsnkS5tW3ryOgO
4eRCwVkVUmvNG/PMoJH2W5Cs+r/47z+onSd+MvUgOe7Riv9j8MufRMiau7rVfWyWxdE8IBGdFwxV
Z3wHJJ/k9QFpwOk/m4NvdKGMyO2XNLPGC4oQqRwdYXb6k6XTYKChewephXHi18QRtWFczGRUbEtJ
aRQCyrVG43q8mUyUUEpxkq9I+Opt0+EeFo9rWzEAWoLFF3YolNlUw/Z2EHaOyet6M3MhoVFUQKQL
ZVIjFWMObyYSHlqFIA5kZ2w1eO9678Mr/ICPVXzzJlTO0hDKuz+XubTl3cIkXGvCS5X/+juZmHyJ
CVdOMoZ13LCycSbvJAemBqDjPbuHDMSvx18hV+qitgrzbk1aEbDvAmdidiw8ggVredT65zzBZUwo
szc6cs/qzvrjVRIVyZ80qIaL7sRF2OSfHhVwjv0scyuyzGhstn+SK5r311O+FIBT4QONbWTzyIPo
WXurCwVIsMlN3J+ySktc2TvQMk7805/6QqDArjEa34V0rtIjFklrFj/qzKNZXYH6PNn9D+L7FSM0
npIKAkRbH9ZyvkefW8Y5SeRzFK52pcuk2Oo6jno9gv3Ooj5c46xclSvfIxJ8D03Fu0StjiPxEMjp
sRJyJj/93WKUpec64rp50MSAM+RROPA4nPDmyMaVebcELoczlh6Wfr8iD3kMSagaxfGpgNxFKISM
uH8zVuTmnj+9FeTPrUz7VU9J6iAkK17y3BzQFoVWufXd1VFSXXcMIQVGI4xZ6XKlQsGZuuo5ushK
tD39/18uxjHDoBoXJTnkGe34obvFODAbnVYGaEsFnJy65vLTyTdPShkO1cWlWJmLFYLpZmyP088R
JJPY+tlV6I8Mb1zPOTuAdykeVQsy9FbxhsHOLg9oXyAHGNTtpnLZIfV+TgGSp8q3H4ekHGgrSF+X
o2hV/hmCKIFyTQc+AZTq18L9eOU31hUb/AJlQlSeA/uAmJLnh/Gg2Ii636hgbrGTGD8dOIsnbQXm
4mrANOD/x0z/ICzQr/jmAmes/zDvEtzeSmDA1/BJrh9oBU1a5vBDiiVUioGPOyjFeVui/ZRrfwbw
Dj6pd9bFdmzxNsHBU4AU9NAl/68KqpZkr1B+qaxJgd6X03sReUgklvURgFX8sanL+C19NmLKdufp
IJzNZwDhUMW12oztV+MxPuEIBgtD3OWBPv6N9vfXSuJRU9SAoxtot86L+LOo82RBEiX1ECoA4Ve3
v0RkPANXCoyqXEsg9DNZTbXcHTbE+3Vo1ekqmYv0cG5IXH6gvTXvtn6gx7tY5hbS1R1QI2K2+BrK
woqYatsYPmrmCq434HIFZzgriyqOPk7VBGPQkChPWZMHSowUodFJL963vOFQeGBbAvT8r4e8Fw+v
6fuLmZNuFS8dwxf9PG0qHHuBCHXAUvD82GJ1F8RqSaJNf8WxjgY+qjjsBYN1sBziEKk71KzznUIX
uUs7ZZ0zgoyrGZi0zUtaLOnxXO/vuDxDvSWZriLt4dY3b4Zzi3keT3n+WZEsFOe3mE3EvS9QFzAx
E6Bqhy1YnruSNy7eorKptrYTRQd9vtJfLScRazuXJmx7sSQKzQ5fR3A2IU6QwCCcs0FcrUQ9timj
Xj4oJMAka1T6fqsA5tlZf6qEZOF3KBNawZVs37nnzPA2W7j8woayQoO4aZs0lkYdmytzRLwuqbSy
9bf9yLT0kb+uVnKUTV1srMC3B/k85CunD4CptcrwTClvnQHHAi+UbfjSmcu7pORbVYHGLkXf5axK
rwA6ClMiqwSF5/nE2AjGJ5SyuLH6wMMc6h0XzjyvSxfkxgeBYGHfxrsi6OzZ+SwFpNuaumABCJ+G
PPdGUPdh+E0AhPVV1hVgM2LGxoBNh0rAMghsLThoA+xxdgep/nr1Ks78nPepFBrOkuV+vOgLAiQf
EQ+DdLj1OfkbiC0SAQ+yd4UKkYVpplT0jxZIS0ThCWAuHKl9ShcbPPz6Mpfvh4t4FqULfvxtb2tu
53wgIbPAW4zHxTNgC3gEwgCbOe0zBTDuSdKDVw7ZNwNHMpqPpOHCZwIdt41tWmnu22zMTrEX9YKE
7oOv9vrSg8VSbkqPsn4gDTzB3SDgcCZLx18v8T1qoEJw1tY2MNO7GtiP2TmP5mg9tS9NNMMJAF0w
O6UCpw/VnNMofjaLzayjqYuWTJCmMuPe9U+FQPzuiyFk5e21SJGfR0AZPUMFOp5dLMaDc+bKn5Sl
NdFbd1dL06wnQuZQBqz2tqo4/k9K+6d1Xx6LnN+guefXpQunbWG50GeG9lSmtx+aOgXYxByujgxH
7CC+NjzHKONu19wsA6+jYQlkSk7rEaQDnd1NrDpMvY9AK0qn7T3ITKE/aAbcDfbOpAyhjXDbhITw
C31UM8R/1b3QVI5BFivR5sodiHK7JDDzZrCrTXUgiqQEdZVF1nAQ7sBhg1i85UaL2OM8moRfe7mE
8Tw+7wz+ql832+6MwRmmD6C8kq+U8WyZtVEhHIL8C6j2yR4JY/GQuJfo68y5f8/khdQ0TipC7r1l
YSB1EEuq0SwsaiVaY6xdKOr6sQpIh47bQOj7scmAfBU1FLk+o7sWmcsy5E/2170LznHTKY2BBRGx
vAUKnDQGvASoRSiRGb0r4Cx2JdrTs3+O3TA1RdD3FmLCWPiwaLR5JpAYUO5Zei1X8cFGmUmElauq
04E3+csGqFyFHNWSYkPlKX7XwFQVm+58x4w77miIHiMF42yqoSHsQBE4A1545xFKVjJsHhJOGl2D
rQeUEVlegrfxVDwgOxRz3Tub10+FZPDEWmUv7/eiF3Sht5DsVO+i3wxq4N4pGUCbZNbsZVYDrwLQ
OeoBhj0SdZiCbZ/JAwbfIDgTxEtOW6jIC7IPfKA8tXwEP+eW9Dsj33NKdOkhdzPFX8Dazf3UB47u
TJebe7TMzTNuD7VSwl0aZ3tsAoUuii5mUsMZI/A95CTKyAVXYZ8X/R61sYpETQeZkk3aT3NNf66k
3Fdm9tM6cLmbHVSGTEtiSIqPj7w68SO08GlyKiyTpMWEyrHlsXvVCp9DtU9as0W6biTDgUe9Ol1L
/IMiXbeFtH6tx1txumlBew+McRlO67bjMWWdcIbuPXmW1W0rezAcW/YgLJL4mX39QaZRczUagRBz
veflYDOUACDU3KZZom8Ql53eBSNRWB7Uu/ptnjzf5Rm0VnHsSKHeXiiWRr6OdQ9e60m8CCAFtjMc
qc/NuVNsnrIwC5CTNwXWjZCQtFNL8GJ/2z1ygB1EmGUvgTHjJe05V1l2QXPR8k697BxvhmQlQ0ES
tyXeLYuhlTtAm3/kEeIZ8iNDAK4SbUgTqc9f/ySgzA0/s4j8Do9ykIpYSdPmYYZtYVjdWm3Cg9u9
oC0IZxj3qWc2/L4YEQaFSQdVFH4TkIWjOum+4ysP1a7GEd0rT1/7c18LvdWOS3tIUDNe/j2Z5cRI
UNR4v6esmxKNbDBECybo/AyZ2sJqM+CGe//MIHqrbptUHBXqjosJI4lQTHWMRR0kddqP/XTHKnEx
0h4q4sRC+TqQvELIz9ufOpqVDEmiLjwe9hubtEqyDrUJk86KD27x3aAKYSCQ/NDTAfCtMuLYYkQ2
Zu5NzoVfkjSvWZ93ukQK6Cxs4wG21HI/sgJi5+9k5ndyqsivWJN/yOPHOlzhd6u8n3J9nK55MEBh
Xr2X9Bi817LTRm9cbPWxOzANMfEY7fOvKMC9bKqbykXqDj4NXDP9pwn5j5kNejBWTyWdSC3E5ZT7
zLB7+9m305kgXjq9bouBXhMv5Rq9AgyDe1rfy85gP82puTFVDWxKWa70t5dG7ktyI2HBdebtt6ip
byS+FoGM0d57HC8/+Nq8kbNdNRpfAQZ1Gowt9JMbpt+bT5xcnaxCZfNQxG6uFJH1qaYP46UKYDZ/
3cj5GOqtgNvAfKjwUkvwosZKnZ3UdyjybWGsooOqGcDvOm2G9E22xft34ijPHM9hrtgAAdOwRT0+
DDfilik0o2vLvA1YIXnOZMx2JJ1XCoUnxyNruOr+geIUoBaa36gAF7yUoOPlNmns9vWvT+wbtLpu
d4ejeEl5GR3MbWKoySMnf6lyqr9iNsAc8VsAKlp7LRNvyy16c/vYBkdAZHtOG5AcSCHcF3g9cv5I
YuuALzrtOfL35MXPDhS46BG2WHmJW1PcfrnWqtsWML26jsD+WgcXI3jnSZiVWc8TI/bbq4d3Tp7z
bmggW4M47awhU5gYIi0Th+y/HtynTRZv84EDN1MgM9vww9CJy/Qe+PlPVUR9EPcXL+Q5uTAztnYH
0BUT+K5OOX4mrXccJxah1g97fabY9PmioU7gs6ANxCqMr1w6Fe3zsSKxDBJF6+0bPz6ktEhvAwVu
ITY9EVFXdLmfuMU6NrBejR82aF5yzey7T5Y9iuHWNiQvAFMppT5ie/48YpFABzmcmdAiwedZfmsI
l5ZT4LGv7r+vABuIXrw/nKAK3QUqh95UbbMUSg3efrR468F9BhoL8GEnXZEsa6reDhEKiXSVkKVS
pUG/vlBJMOOVul/yny35MkZQwp03ggppJ9WCoae/qAzXz9XDwVx/8iqOcy6oq17BBAAUBEd4NvSi
sbtLW1PnXxvaKfrZERE2TyNYSaVoSfGUe4FcOuXX+qZXC+p8emWgd0Gg65L5XgjbQxHmmauj1cL0
6Pdmh+zMYdjANd1YW1dcGhOWgkNNPZ0fjHaq6+pbOlybwE5Eunbuwc74hH8wr82P23t5wEi6FfHT
uI0WBF8JRqut2p/sBDqtF8ld1Gayq/mG49tOXoE62RtfN5s/O9X+/CUqCcGJrVX2lgD49ZpxRUTG
dA0F3QNogCnW9LV2liAFIe4bLCFzZTYgzCVhFyAFriTLbRB82qDkr+A00iQTU5Up3IpXhUzY7qZ9
IY6/1E7jXcShYPHos3BO3cgq5vZOJ8cpgXitEcQGk61JfvHNB1CHyIvy5sXCJcyZPRRq80G+rwBi
v4sezEbFwFWRgKONRV9ytPqakpmgT3i6xpwWQ0H8GEWSFcF7dvX4RWcuPhz2sjB+TDNwd96ENOTf
+rX3UjL8zViiz2erlYHby3XjeU3f/yGWq8B2A6h2rgcfNEUsl0wGGQYHkW3+O5HZdnqbNAaQHkpc
fbja9ZUhD07DmZMxM4g6qjuMlWDgLpwuyQ41EE1r0YL8JRuPCzEdT5fVOAGQC12ll5vtc2dFOSx5
ZkNS8MisxjtkNrrWB5VvKpCqudyEYprb6/+1X5u9lF7uX7zASE0BZjOMp+dpAihEeuakfIZzBBzd
Kap2Elq+HyaF1f3KdCJiGi7OfkRY68BxbP1UrD4Lcvcrs42fM/iH269umkEX9XG0PkdIRSlDh0K1
89hh+tdmjobConX46v44EZNqH0OHPc/tIF+8HPWYC+Gqo3+zwta2mtuOBMo7Ybv/iB+Oyz6b/7AG
PE4QIhNbeJnaB/YXdogWZJUAaG7DfXzNxymuYsEdSu6jIj3PyxZ0H8p0N7DcQEAt2ZulztXXpIuV
dtrHqIpbJrNDtHzauyHoatnJHBDM6uZ6eVjJSGNzUCTDvBaAbfPcg4JkCDgHnjdSmiu6KVB7OqDF
wRtFiZfZ+QV825dqYUh3DGH8HnVXlyDM5KJihKsLt22/NQpSAOWqjeBu4qOuKeOMhwCPZOSo6cxK
tnG9Fpi/vX9kmcecmSDvwn9inlxhAvRc79rYmQCnZGrR+cP/MjtRiKgModvf4BH1+CgK2SIwUdMY
LzlYDyiSwIiSm8WNqOXwm/dnECK+FdUNg0DrF03ms0e84tF7KelCEYXAvMzgjcmPXoXaejEO8MPF
52HcWfULQOhCv3UVMOwfVhJ5YYZAEwo5xLcI8yiZQO8nYHzKLthQkZ1aNHGDSxWISPR3vYZmnkj4
fh4DpzU4jI/uuEheRK0NCyYlv6D1ZiHVm8cAJla5tF5DtaKHhGMLDPdXu95eUHB9DcfhAT/W2f7E
JgbhMueuh5mz/5Gv/dhFcABR93a592WHryfwRjzbbVgmDzZNccdeYamQB5GiyqCp2+f4Y4KkhRc5
q8sb1MocW82X3D7S4hFd35DdInV9TjWuSkXokiySa4ggCmne3fH+GGlLGSpIeFxTsXY5tZrPr4bS
mTTORHzXSz9P6hpRmFxGXN6Qd5uXJJcugCjzGXP5ob3ILrpTQk8zW5Iv2g16qAcE/S0q7lv0JOd+
Oo72yCrSTm4r2QNBiJVNuGA1TNCZPtE/QrUCjfE9+3iL5EHykX6GLsNWs/MQSbNg7P+KlkZMxmuO
JLQ5ZhD5F71m2mVjt31EngApzLYabz3hwStzkHHt64cRskQFDdkkgCsuB09F9YShHAiYjKlEOcdh
z+5mbplij2rW3C5xgcFX+AuFLJn+EhRqRnKz4Ej3pKaNNKEFGm76Yj2V5bbxrkETYgQ/KJKYxbWV
6T/znOYOvF4fGel2d9Ox1J3KEO589XnaRu3GbXJZIdvEbAEyuBAd7idLrL5IyV6h5AH2M93BWx62
LjOGfX098OeMMnksucEPnSUuqEVqZ4cDNDrL+jbPS+9fICZVPrOzSdSk70dAfGmZT5C6iJ071MMG
6+gTkYcQW/6FqqDqhnr/EbSFjt00R1/exHDlmvbag3+tIVLbDtY08/v+/fQFAfSA6STw2KPXJOls
zEutJojljRlkqOBLw5okitW1qrEuG0roZ87YMr+uFsDJDmNEQQL32d1pKSYrkulMTjpXZ02YovdG
7eCo5F/upTUry44AVK4XYjvKjRDKYRAVWbgrVu0Gc3xFtj0cKuMZg7SS++1CLxcvcFNKVsx2zSG6
7WwbPZhF52PJKJQzUGEYP03mw76tOh90I6/c0eXyG7WRIMX+wyDQ81Q67swkEhyG2oyBcIPWwxeX
mlRx32qfCWS03gPS/MyvvMwDR5IouVMPAm7yAvdKhMl2IQK8mi79utg+xAh4V3Xy6kIQw9Wa6Ewv
PRaszT09Z0oC8RuSkCDlpwBp8K52WR1O2poAhqAkjBAGstSFeEFL+oUg4MfubDVce+eKz0ZTAw6J
HabteYIhaw++dukv00uu9hPvRd/9Bbp66zCYfzt0TMi1GLc45ZoSopaK0WbipburICHWORDJDZFp
B7shV/UrLacJLiknhADJJhDBhocaRkhm6bwkIWlyQYLIpGY32DMhq3JZf6Uqfiv5iA/e4Rx/l4pg
oua2AOSr5WoST6ffqORR9vO2CUlBzigzlOPwPiqUF6o5NwYWKAneosfvCRcLRy1s27KeIMqY7Nlv
SlZZhZeTLRQ5n9ZXj6NxwBEJlmtwixRkxIKlIjfgajdCUo6KnhWLg88bTrH+gROVjZugv/Z1EyQ3
1Bpgx7mk/WOVzTEvfDqfeD9vvIOt5CGlKZe0PxyqdTDvymJWw7EzVLz14z8obzA/KUn2zyLgEd6j
I5ycY86c3dVTNvL2CcAPUwW3ej0NWQvVdu/+tcxhRfFbav+RHXO/eyW51kknSrnFTF+w/XSepcJg
wBm8DH1LVdSuIeL03FkqAXNW2dMxBPmt9ukNAYL27kKKWc/2NXVUb9uBe+oWlS39Yvdm1C+QsDIe
PFed1rKEfOEoWsGPdKGvwXGEWnA/k2vvrbnWc6JU4pWhvGJN9rwppxZ/grV823rGwmBTejwrVh2F
icFj0Ft+DCVjASk6FPNuWU2r69xyr3EZpDR4gr++GEIx1JZXj0iYRGnnuvLFHMNCTpelkC0I8KRg
8OKZFN96epxgjrEJxexyVoN9lslYzdj0AqUDPR47O9EZJtzNpnZdVzj0pSgv1sqxanTxWJLJEpl1
yarmxLXjYdOl+178qgmEl+sw6KUQd38GVfPBY/PCN/VYTT1VAtDLJmC6e/Bbwi1X/UmWsp7Xb2GH
s0JuUZB6EqrZN3fEIzMFIH9qHSAJfDZSUysGlRlp/VylUR1tNZZF8hoCEVFpK92IQfgoemwQDKFV
LAtS4NrBcR0tdYthT2SUQBdH6x7o0jFZAZbvwPw/GEDpzGIyXkiJ/thREMGjVhqQ4aTKvRAEGpkk
FMNFkvMlEECV26YfVJhLrfxvgSEwWAU5IilPeBt4nNkw5lzkryucG0iYy5fwE00ZpW+yQW4+JoUt
PUJ6LJ0eQ/aPwpciFs9u6FnHz0Xnf4SYVKdcm2VzpmiUFObDhwfKwiCaqu7KyAvrTkYrF0itP5uc
5Ta6EZ8kwOJB0smKqec8UCm3fP2nvMDAXlmYxQ7M7aspF12gqSDspccRlObX/3MdUCAxOgFG+HVE
zGz5uErUkYEZoPJyURr2YTgj12awKfvsQBhiyPr+AJKVJbAuZZt+7Lu5AWCjakiP2b00oWGf0UCM
ZAHGOPp2Q3aDm5go3f8QVFRS7ygX6lDgvtbWasXIBqEFMNzXjsmSk0CHNxvqzF+QB791d/+SNypG
bFKsxIsO0G6+rWrqBvqyDJtCCeQCDqxvXc1PUjfyraOMqJHRLrj7XM1OnM7BBMZD+MnYxrZC5xUf
TznfJsDTogQoBjWrmabtHkFDoMoQ4M5Afyecgt1ichR3xWifWeOymnhsQmqwM+b+GHD31SQ2htl6
tTIO7Gm4cvCfHdS6DgYhrow+41lxMvKppi20fkdqOn9INvRP6VwotgjDwr6Hw/W5gkbAmmjdkk0H
iAbhgEK5OfcDZbuumimvR60LIcJ+dwdBcDAoW3kmCrTBHusE5zQ2htoc/mNryNTatkwQDQzWZFh8
U5T3Qc3pR7PcP2DscIGrr9e+vsh5ri0nEElXLkXZKUVs0PCTEt3czR/JH4jpp1PBLztylCbfW1lA
4zvziWqIfkEsZ+sxloKyhTz5eSIgm2L5NFUTxjhrzZ5D5hl+BsuucGxFlM6bqZMFhiWxoiVeKUGD
FZmVrW4xSM1jD7eHyPcth1kixouchIsMq5xwmX6S29K03h/NjwwQXrJ/rnkB9pO/7kC8oztpnd+3
m+IoueQQeTpKjIqtIkiBUzjMqRePGaJeJSqbNasMkAOU4bs09I1Y2N+8y3OehesSluLytjQ6p1U0
bUep7f+LZIvCOdfK+lkAQW5bBRMWUDOSwnSVANrYiAd0R09F4/MnvpNFZbLwvgLoWYmJ/tQD4kYn
hOxpYM//lXxWDWgEPCQVBHKl0mZOiN23gHj6b1h/Rdb6mpx0LvWIg27GPfpU/QCECaDTPET9KMyX
dr5esf6sBjRifKoqfo0AzjFPiNXy9wrwSKk7ZbCh3VKKtjNoqXjw2sAO/yNBfT4qBxwCmEW2s2VV
AzgJXWUIMnY32dudwJSbjtBGPfmm+M3CEOvPbBrxtHkSa3wt9q2T84ZJlste8lI2wtmP1O7kYR95
nYRvy/ZMMGr2PQn7wzFP6HY+FYyU9bhg0ApYI1+mPi/8lDvgroGoHhgco9ul4EHWnVNYLcOw4LxY
o2yHPNl8O4gaxHrMbtYJtx77vpC0LUVHRX8nbgdJHPsDa4m15eVCkt090OekiWxnxNHd62LfAO4y
0dWJrkM4S9QwVPtctEmFXoDi3bKdLWxr2fKNXGYD6X3NIvHBLWqtaiwrEyYwgvPdXfYVOPuq3NAS
cXXxFg1xg3irrP+VcgrqTVXTTLmHeos6uZpLW2ZjaOgF7NKncDScYuYPXH93qFBc1yu/lzEs6BGA
hUYMViNRZWvsjOmCa8AZA9ieyHssxji13hwvMVZQAMmFZvSzfyIexZ/rVUUZFGL6SLE/+f5sBh56
n53rzFhYqKJjk/7bfxokaWMrJQ2vM1927y5ZM3+SKuyvRG/92t0c1IFMV3RFiT/2J5nf6MAeJRQk
LgD17sYaxPVoeHNAS8enKWJTYDfH+ZeD4RTeCX/VI52N8+6XNd5M1/ZoxsJ1iztpJAobWDsRCToV
hxU7chvK8EVhqg7eoR9DVQ4muISenyLN8UDNoVfG9bVmrSWxNrZhS1g1KLIT7+/0ZvdJMYfpoEwy
NoDffd/eSXNjcHlyEEaKHZtrJ+vtG0VOUwr/iSk+GITg5z17F+kEX7jjBNCnMMvI8XonWpqZJII/
+mv5tLY+AhAFisMwpY0pwqJy7/sKS/yfNPwC2j0MPArLTkndSzWZkhi6X8NW81pav8o071BnuwB7
r+vaS4Ty3j5SXoCLSRGT/sLD+RAKuZQeERqt+F7mGvzUcJWItMLnoNOFyK5FqL4RRj8QQGaxPlKc
DhaihE5RwTJkj3aaPR0/2Cw6qx6nCkwaWwavBpp/8obQlVZw8B53QUE8ZMUrFi8aXUTOJXJw4sHk
ONobwgivIosM6GCZVdi+QGnrm7BRjr2TCaIEgMo1jz1+JQoWvnZGUeXjB+yMmXI4bnsgZL8cSSsI
SE8+hx/xw4NFWFBH3kaFVsWETbR9TjK50OvyVpD/KV9PXZc3ctOVtjoW66X6rHm+LqYB+lBN19ck
vsAwLhxSahOKUS6lm/RvaqPDjRUVvVkkgsIlX+ucTR+LuZrY9TqTfsDHUAxS2Q35YEXgCnuunEcr
8bEqaWJ7/sxvlCYucoQJDMfe/qR+sW8w3q1YlUwlpvNdVWTQxz1Vrh8WbGKrRGXrGuhk3dBRbtBY
Rv5B6pYZd362MWLxSENw+5ZL1VocBw5hjbxQHhDhhXp9Pe0vjdnmxD0HTWapmJYYgW709dboGogu
JgNyYj8GVptt+9RIPTpnlcPRQjtmeMzrH0Tsk+Geu2LiiAEFZEfuTF6TCMwywogh5EKPn3xvB86B
tv+bNOm0msjGwoFMNoaSmprWCcy/kbIFNrw0qfN9Iu4bXQ2sVhrdbvHcezFZf44+HOcMqGB1t8Kj
9nNfqxLXLxtFMB0nw8IHc6iqq74JbvBqVBqWUYUGin25uG4vrtrz5sW8gYeIkZWwc8Zn7zZ/Q712
cjsgA9MEZrxDAhSKb3U/zIkFEjtOdKh54+HKgtS6ipcjKkjLM3qdbBkaW7eyYO/qXDOsCGSe2iAH
ubFubgq5HIm1ljYWH5XY/b+2cyBgPOGvmpT2hrDXcIX0rUWMsru+qXE+62vex/pdFV/f9gpcx7V5
F5mmQ5vWaKKulNVqDJ+uzYzKcqYv50oIT/cvwQoc3z6haPZUV28GLGgW3RPegvlPgt3Qxbnmaok+
SXQEbhYSUAY+wQatPJwyuYoqUYQEulBekz/Alhwmq90lLkcCVFgVxlPLxevso4QDFKVzZF09wBYq
rPmu09hy/NyyKb7iGPDjLxmW0ond+HBn6DKqfbwdVoQ+IQePSt4tBbpe9b+EEpo/pKkTicKpBI1A
GC7iI3Xofkpt/syaWF0+Dw9KXm6tthBKjfbafsdjjhKSsQn3bNmLdEH++tUy/h+a54hneuFxyl+t
0YuLcaAZN6k1tkR1fCSoeGvkXkV/v2lB5shtVZCbXQ2LZwjIZm1wO0RWTuJuiZUEQq73e8DcvAdP
RJ8QWy3rEQ9+/U21hEh8gHYGzbVvX9az+oq7kxvOEd8GMScqXjVPmIRJXqfIXk5fpG9a6CoFf1MP
4l1ta1SgIu2CKcj2U+64e4TIXJ1bV3RlNoiTfnT95FjTeL+4608lm3JYn2PlI1Vq7vk43MICUOg/
vT/h4OSDbIP6FaOe4XpajkxLBOHqhZ/+/S2S4laRZmvXbOpJiHbYdRDx+Y0vtu6Hgo/5R1Etu1IL
MktGLTcHcSJPsi+po8bBZ0Gh/m+vOtwsIa1i+9xmJ70rJ2l8NZxc6oncvQSQaIwcyziR4c138BKE
H7lb3rXE8E2/gnLy/AcBNR8io3snukMHgCc5YtJsbGcolkjGGXRr72JibezbUWUaP16l5L1iGsvy
HLF7guNYhT9bIPNdUqpJaQhKNEQ8IuvtAazFVrvQs+XyuyXrIbETe/hdX5QTHkL6aNiXbUwlaFyf
4sMufKD6DOVsgnNnx48XHI2ofHuHRGXt6xY62qvjSwBBCC/w2WW1+5bODaUx2Y422GOoXBYv9a2f
hhWSHysB+egnt8NxVYBzb7g0CI4/vp7vNCNeUBBeyS+4Pj07Hx51+CCkWloWz7eKSveWTKhDMAfl
q5fcvH8vlTV7cnIPJIbCu6HU3iOVJxnLzIitjW9TNc4z04w5DtxbBncX1+JNpwY4VFrpJXWQ3w3M
Q0WXcNLisOXvuiEYDRKdAYRaKBZTbr5Cd2UM9hTyPqK2CpWxHP+fx95FhlXYRjBTIbNZmAEn1xNz
FiMlgpAA7Xuci+VkzujDhh8RBfXI/k0mtLTOhlVmPiWPFI3hO+ie5+KDtCudhxMvRMXxzW0oYSMJ
SGdNTwNKrh8vnCvabpj2aKJsBFweqzAP4jNoOyiQ4wHMM5pAc3HYY5RNbcepl8sOFjrKyzMCOUAM
Z3loCoBf1UNpaCNuC5/lNAobItHE8BuR5VjgYGKda37CQy5c/QGew3QLIfVogARGhPl8Mi0pwl+W
Db3e8+3vOpb30aKB/aIR88D4utQv7YfpfOMOty8ryr8eEb8GEoLnHwI4aAXWSS/gS4OPBCDIqS2d
od+SVa3PikaQYfhv6dJuqSVkDt+Ge5tiSohLNkOESczg12m2nbPvO+MQWmhJ3muet56Of5FDfCMA
7ER2eJqCoBhFTdZe+LJhOpxx0Wqct05cjDMnZbkmPd0/beTTWf5BYlAvzzw/7HoSr80aOSZFodMo
4egl35WMHDFK9EeZi7iS8VA85pc+UVIxIPMyu/gzxj0oowERpqXF7LF3o0NkFdwTUEvoKqY5kKdf
TqaOupYhQsWKhRqyCMBHlOGvoQ1bsDWSD53k5LevfInTSOI5/ka4IqgRynh8AbnDQNAhAOOOo1ub
zUGI9i0av4r2Z2XKH7tVVtPyEZb/LQ7w1E6C7czl0WGY+4XGCgcKySgd1RloH9hz6UWDPwDv+eYd
9MtBqQp3jfusgtUApNxFwMOo/JF8l74UVtJNaM0Af3SCku2NxRtE3c557CWO8rb6/4OxFle6BtWO
bZlx886Qz/wF8Ayxq+9gun9/chr5qFZot4fwRJ6ktS4Bfcb7cJeLHMGHueMYPihr0+BihXsrgeI8
s1gzebdhBsZ7xuKuhloOJAv24UPCjEd65nMOQcLP9vnXPTZfK7HJVTonqkB7UAXRQa2FfH9oPI6b
Iz02EHY69t8jZHtj7fBbmrz6d6HVsRrAZl0GZHxLA0+un6uWJgVp7c5qE2uQK7BDY8p9hi5ZmMhk
gTpAC7uR2VjrYFefdXPF5CZPBJOg+8REa8WUTsox1jR5eayCDXiQ6vSU6GiqVCxfylZXXcfhroTP
p6NXhXVw6VsTdPJISladH2YriBQ6cjsi7DrN8EBUJFhcpJlhkFcgfzQeSUpoVOrzUcfKsaNtuj/G
BsLdPlwmWzC4IiNi6TICVteIGQ7BtFrxUl6ii9WTGHVevh1nZtX4UOWVAHmxwWzSuAjET+VWiOd/
wDRwfmazZKpkdZFHf2AXxDLdNvF3eiGDfJZFZ3l/w3CfNLmzzSEYx700tl68XOTlUPp5rhrNu+qv
u9lUordnHGSRLV2FN+pEAgiqEQIPjKnKu7X9GNlGyeCHMEUJOIJyANq3NUKcnWS8Q2GnAEIWm3xV
vOZhCJimd0kwqG9IBw4y4gxH9Hm9V3YRkDYAcaeJA3EeMGsBrhGpWKkc2dgYRg7INy39NLeb4X3r
cN0oslPnLJykGGydLxyLuSeXoRkccO+OOugLk2mGWcA9da2xf5WhkPS+/ZSp1rtPCj+HP7ngVPxM
hw5GF6FFsQHoU6J2cmnUxkMwBvIfO955uukMpLOzuo054FDzr00v6wPXkad0aNumNbWzJJiseAYx
0w+ZZEjqAzQFygGgAp/y4jhKLx1QpPb0ZFxrR7gb22oFKetk09v+gY4ix7t4ZD8xLt+jvinhNxhC
BCbvc8yh6pztqgqNPs4+A9UROhLg6HtMlBUb/ZzYS5IGeleWQfYQxeDWl4X3hzF2YIYk5rrTUraD
MEHDxfmJDC915+VZqoatla1EwPW0/U7OG0m58S5mITQ718EcDF3k6QUfwHTA3HpMorDwpg/Y7GJp
8M5XvUFSoArmSX1A0GrMbA5bQmfcUHvEP3EJIv8aKIqnzcNI3IQX3OSOn+9drqf5Fbbi/V0XjA6O
iiz04RgtB4d+CCpU5WGyruO/4cZ7tNyDtgwM7qE86U89boxIA7MT6aGPIOR0JWuL31GlR+F3G3mC
Fis5cirMe99hbe6/9slsDB1vXflQef/SDGeFxokspjUgqwAL6SEP7lGCepH2Kfp0AXPboDYz7pKn
7QLfP42soHQVCMsjivFRfZNZ0JU1tKNV6eenKhLGGL2XECsYSJMnXXSYXzbgYtnkNZp1VJqWANYZ
K1ffamYY/CU8R3qKzwI+rcRM498t6jXRhW5qpPC+OTuOIgYA1lS390IupNbDJ1UyjeRVllqM1Yom
CZqoZ8XSUIXSWFcHn2qOaoR7kWHpIt2Y4Q6dc1y3pwLz5kBhK1a10fWfv3lOIhwIN4WwScFRVUmu
cHjEAtYTJaCTICAUcNxbtQFAX0a1G52JW5FPxHVQjPrD7vfb5CmKWLCJiQqRyZOyYzR32HDzqXrR
Xl+PgGzDuUTF/VMs6IbcpBRU5xa3GKTObl/v8SIpZUvnAQ2//bSTv68rCXGPtPYiPsSgO+O7oAsR
fnX4jfXBtFvv35ou8NhJyGjvb3AHd8+jeZDaCgpPVyb3aGbOw4agcx1+hRCK+805l7WxEnmPzJAZ
gQbi07r2aDJlFwlqWdSuid2Hi7OE00b/fztURRQVq4C/KdJAuaBskFA35JOcW4SeEt/cSnnPCRjz
a0IbUy6ly/rESTLHcTJ69uLrUPXytT93DLZbwiMrf9qud/zjlPDDyG+yaL7hpSQG3038a/UjSaO7
MMFyI7jYHr4jrX74jDfMXslWuXGGRa5pNsMxY1Oj1NDV13dvaHrVbJoHMD7/ewYYTJ3rcat0zYrm
/C+PmT63jKP1smld68ZVG4guNs1ps/ojl4hiBKgBfpKoP4xn3Kii4PxRXDLy2dJw0vqf9DPKr9Bx
LUBgpDHqZKwU6hvlUXnZ66mxQtGZuhGxO0GI58yLXyT36kNaFnKfcNPdbRu+eve0/x3b3xEdbmvg
0QJRWvwQWHo1Vq3dpbnzEqGR8M1W1SZY0cON85uNQRs0ABpIftRG7ai7Fj2q9ZkTcOtDvETtgCbp
4+KuiSPl/ZmjgfOhw7yz39AMm90WFNmliGq9AjcDDKUE2c9+FI3b7IDhmNk/ngRT/HeHWLZZQfxV
dpdfJG34uCoX25S6QErqT09ogbkcSPN+zKobbdOiDteH3CxvzxUVzs2Xm1dc4/CJVxQTLbz1NtGB
ESM+Pg3a32FcT+5EiSsYn9Tl2grjpRNo6JNmVAeYd+KfFEVa/3PEV5PPDUB7bb8SeiY=
`protect end_protected
