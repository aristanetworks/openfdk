--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
BUUatewsQfbmhc63sWF4OJ60gFCMj6XVOwIjWzp4Pvou6ryn9TeamdshNqLwPbOh5d2O80ocqiRU
ePjWfZasrruGlZhgcBHF+72QLyP3B/BRt4X5blQQUs9c2pWFEkxigQJedypl556XVJip6ZRyuqU7
Nht4u6m/P0hKNYGMbZkl5oG2j8t+aK6xuTG7/PyjffvR1LTzppSuAJGUpAq1GD6McJgtNdZN9SQk
BWA6IWRRo/wPvfIzomgO5bakVqlki3oCv2y+SxHwkN0tr3QvcL/EwiK+Bvo845542EbDEHUfBvdl
yfQYoLBAqZLCFJCtROXsNPcu62ORJbLDcaHOBg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="LV7Dk+lq4obf/Zu+cxjYmGhqFqWlmKm8h7/MRMohIrE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
mpIyv0D+e3LxNn2jGMQ0utqCGAw+SBVCemHl5u+se37b4ui4CnoY5rMjCyPUehrMBSH/A/Xaf5V7
LAttdMQeagljjVB7p1UZaiyWMIa5RLuxXCbkJy4uOMVAEaMArqcVOKjvfxO1fyAVN1qOnDB/eCa7
l/kYTDNPFvetfb50fKntlih/HDh0z5V2K18glOC3qCLRKA4vTm+iiBZhaA1D2TXYsgGweXzUASOc
STPt5wsNcrJ3Xn2HUVc8VKRn7n8nXAVs0dcmDYNrTZf7nEQ8lrtGpQyIR4B08FsVDz4R64Az8lJL
fIm6mfCRHiQVk4BU++9+CqvwbcuNhq43/v7OvA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="giqtXolxAEJaLTpha0a65ruL9fFs1prqW0mqzgHLrfI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6624)
`protect data_block
P+bzE6Ky/Z0thWR82gOkdb8q5AuhZpyIFJqpdvB1XsQRQQpUPnMCCZRNUpa4if4BX407w5sSB0r7
B4WskeppKKLmskqfC+TUpd8d6tlyzlrwo9Pe8hiYTaIcm7p3cleLYp4uPdlQXumX7WHnED6FVRGS
XEy5rOhrkDTce4mQMrW2M2UAGdiVZkvn43OXsoIHMI5ZBHwJ23OEB0fHAS1m1sKY/JzFxBEebhx7
MU0LCbB53rOrl1CU6RPq2BdytMXKLSjbSD6ZnecRKwz43AeuXousqgVMw7KoIRj/wTmm9PxLPDZ1
vY1I3jFwLsF+kiqA0a48ucMRT0Gqoxgn6tpSe19mP71HxFJ/bDvMUdkFlrK37w+g+VREOOK6b/wp
knp/BC7GTz5YZ8/oPRem2bE5RsUehfurYD/XHe1BFwGsmy2bShutbqKOlHngERgVIeW0ky7JEZQA
dNUqXHXc89NhSiIzYVRRqoCLlnLeIrfn+ViRx7YnHgo0geEA7V5hDWsxDSXk0tw7UjrDUJ9rP76N
GCiChXsjf9F/0xXIOtnj2LnsaMUiad9dkmfIwexkWFeJJXlkLzB7tfx6otM8XZW1cYO+SX7pSnym
fj7c4jePHFKlowKSjYyoPFk0WwHplFLVv2zjGCPfRcXg2zsSGdRX9Zugwp09F9dlIJtcbjugPuzy
/No7oXHihFvAX1+nWLZXCawDTlF87sgt+2nbLjNZfu6BdFH+Je3hLpgw90pUk8EId6fHnEQq9lkT
UQZ7bpgPcjifmH6hIDp06cZz2UQO0OMVESJubPdA6Q0WDYBi9p9XXT+HX6XW7kbtCq0UojahbRvT
hQdDdBZUxlIdcPCuy+wbjTpM0XjCzeNwrabOe92BD+1buJXkpFN26yX3IPbKwGdLlPVxIEIYY/1u
lsP8gnQpuEtFuTr0FlYt4oy2bwIeqv6p7pn1l5ZKP+bic/HJl9I03R13/rbFWmyzCfJ0U6uKIfet
AcWPv1DdGw969GkzllMfoSBCRI1zrwmEz6JrWpPJlm9c9l/EWotNwcnwv6eTugBdI6tMbPrtRl46
De5iGDn7LZB8NbUGfBmMjx5lNlIg+I0zlMvTFPBvOQKo0GLcWdXRbD8EDdFd/eJ+WFZmSWvC08Am
0xc8V0EwbY4UMutYRMe4CUkL7RRq3+TPN3w9+uEwJL0nNFGPRAGPOKFStEWkdRslgf1UqD5LTPKE
jA5COHaDW4Yy7G0V/5/6fmQhu7fh8/l0JQ6pP4iY4F9K6JuKoBxMWtaciXDBtNpDlRuESc9MHPrN
VxznJm22RFZp387D5KOX/Kz+yTHn58zUUDo5RlkVes+fSNEXgwZ7NPy1LqhGGAPZQ+u0b1cS0TeB
0Oi43/xVAd2iyDbkgXLCAcHssEsHgE63B7cLrnWDXuM3eDuv+LwVq1OkbKxKWbAxn2odmF+bRc4d
t40N7TQU6kAzRIRBGx5UUK1xxwH5+ykLpKr81C/m10rJ/D5nVyfg81Zq5Y4X58yFzU/YUabZzRX8
uA91gnrD7teoymswmoayvXvLkY8lr2083FXbXEGAnOzvjAsKvpWCqRYsVESUVQdDRCElKUEpczx2
vodJLksE6VlBbXXpJsqp2NjIxS8wPznQS9MJrxmf514sMzwv4FLYj3ZspS4qeH6PvoNPJwALSq2w
BSlUPSKBvUF9ZHb4O6rGslK/WfXsAK5BLkMR+aFrhcs6WYo5ViAhGiAlILVnmNkfJeDphxgXyfGM
AYzS9Prl01bnLWRxTh4X+yD3bRO1BhbtdTAnxE0wI8jXpI6c5WByw2qnRkmol4Kerp35LJaQHFR/
0jGOj5pCl6QKmFUYFxtfQFI/VE8RyYt75EgzG5jxK5I/3nDlBdgXdW9Nkd8WAP53/upPzVdLofHT
qgiW6U/n0WackQVVYDkIAWniJu96nTPHqjslCw4wsEjU9KJHCttcobYRTkIFdTkAc19mwdsqgsz0
dWGhzGvo2hWEXhfnl5lD2tjoViH+FQutBh/NgzP8zcbhx1I0qnfMFyLejth7I5gqdOr48ZKX0fnX
KpSw14z12nWLfuCOE6plHJVOjC7HCk9OIKr22RtIkr0nQ6of9AGNphcaX4FGrSblIcD5Q0c/HCqs
ZD2tY/6qyaGWmdg21wcCEIMpp229kE7Y+8fnpakSBd24gYnyRsHlx1aKIUVLMU+/dMEY66/sIUH5
t/qxI1CpF2ZUYPR43Ss9c82IgPFvPhABPnCo4kaoNTUaP/527+t48gtA4cxVepOincSQsi2Kbg3r
ZndGp4raicSnw2llfAGFtkxqwKRf2yF2n7NvCLwwGcGodfBpOyY5zuDWfted7fBwbvSch29LdSpp
9ZVlzCdhQYpNQRCa9VghfU7rvaXEGDWTDCXIsIS/Sz5GsdGD9M9zftFSUrftCUa1etFf2hs331qd
NtD+yJVeQB3/reXVXbSSTYVTx3Cc/LjCJY7c0YrsJYdk7IL8NuaeO8skCtY3fCn9dXpLu620IHoG
BT9b4fobiGgx6YRN4Y2TvD+9SPNXmn4w6l4ALCZR1sqC7vHRRxXEJDbJQ8fGMqJ4269oMOClQ0yn
RlM88sFajp2WAp2gBBf7kg2vFbGbZW6RMG5haujrzL+sRBQtGt3KtbG0x2dRm8zan42NQ6w/XR1b
dAakNt3Ea2/MNCb7msKcqoITohyV1ce45LFGZX+1q2pGebzCpvn9ovoqBVX2X58z4PyH1t4mQXAR
ZEICgsJPSj1K/f59QNe52ZHQ77J/H44yC3MtYTZUUPjSNQ5tN7etIWxVOe60/DdZslGlexgCuPNK
OXuNes6oeFq9WLKxGxKaTSU291fYugjnHA9ZpV7VFe8sObHR+X3po1Lncz+09w+jCmjS4uqNmwbO
4ywXP5NfmSTzAqndawqLHIR3JHGrv4QCO7vVb6aaWmh+pzPyPuToeSnZOi/hLaYwDQHCjlQu7mDP
QHJQwRZw+1NpnGa/aeDAncvkJKtnRvLm1ORFaY+e+fDpkrtpDyxTvruGhBvsnPF10bO7jbphRKzs
bZycVzPGopMtptByOAvKquIa9mqjSO+LF+7EIpUUZehlocRZ7iTNbanW2wsD1QNkwl+rjxH1lCGa
+9eUbSNUn25mq0ypRBsE84ef6EaBmYGK2niZpbWNyfW3UF6IV1TCNhsoTDr7NuXYhVF544EtlRiR
ab9SqmvMwBKNu+3KDp/LqhG3c4dZvzNk5cbJOfWx/uPxHXbcXZFEuZ85HjGTFKq/n+l/spDsCU0m
Df5iJ4QZBrgAV1o8iswfJ37Wl+5LAzJh+6vi27keTl4W8Vqte9mq5puKWVOVwnY+Y4kh84stFEu5
2qCBcmxOEw20gT83kvW5AmPPtI1pID+z+zIRLiMKXk8+WSGmJYAMmrJ9APptGUZtRVicQLL9Nr+n
8+FCUBRFiYS1STmQ5rsdPjKExFJiBoLjCy+0+MLYMWH3uFQF/a4FALIgKr2gzZzdgkgXSjloscsR
pHsRjcp/ayLyG0HRGkG+rP66UtXpZyx0Gr/QYHDDocyQVuwp2XRL075DYAkrdTmSUwhUInrwgx70
wK3r8OQxnwpFkAOk4EMD2ABUFJjoe/5HcTxfqppfxNKq6IWlW6NsL0kDJELznnjWuHywnN/VDLxg
zoEwu2fthNAXQzPPfC8OdhS4T7STUFD6J877nj8Ap64Q0J/QJXgzCV0hFpoCPHHlDdJGshPUX0Cs
9QoO+q9eulkHGBPkBFsgznYqI9sStsXBKLjsAeJZCjmrTIAaR29Ev1+1wXA/4I9jvJERL6lf/Jk7
4KcLcbaJ3tz2EB/xvuGW+8Tyb4uYeCR2MiIBNYhcIO3CW+AuUvpyCTh5P60VHoE8//rYfB2WOGL7
qyRaNb3v57fQZV3zDDMPVuHCa4kuwty36w76JMGW+FF+cGZ4wEQQT1Ne036MifysQxVS80PyY/zT
WkrZ5Z8a2UadVWmRVHCtjsc3m3lt7aqNlr4FOFmI3YdfxQ+DIGHLXg4uR4essLXwRa5AWyangzk4
UuQ+jfzgKiqSlkWugYsgKWr/5wOO+d2VFdzip2VvU2f3NMYkmGZrgKaFaCjsmrTlr2nhmEoqEZrE
glEArtW51zI+nV86NjRWhhaBGuZMyJEmKxX16s7NJ7jspXj6Ok0M2H5I8TfL9qbNo0dmZmcmx2Rq
hfNmA7UaDexNPx4auDW9A6Dpxl5tC1zQA3nCQBX/bImahng5HkqkRKLH6Iw/M8xiQoAMnZ6AX9gs
YVB61tKhq4axzqv4ZsO4ABEQF05mtIzNaGcj94cWYFxmRY8lVPkA7B1ScJoRnfQUdoQ1G6GK5HD/
wbJNfay/8y5e4TAAZUfckU+wW5QixWOrtZpnZfr5KlJMOu17GQbsuZZzFXoLAkgeUCjex4EwNL5R
6WD19uOaBw1H0MMKY+aW10eHzpZKTJZC9s/Fiiar7ObdVJcDw1sl92YgjB70ap4N2XFq3VRHDiFG
4gD91F3Q85Q61xgYVFCvMIJEiayJJ9/hiqJX2Nw0DSMTgeNd8caUKuCKf4YYSf9K99JiuEn+9bQ9
IrcUa9/YVpXP5qTyNJMti1V/SEnirlPkPpg3YNVCPxr/9oZg9Vg9xxzAn1wH4oIa4EDUpMGI0JKs
BvYp76kiRz1EXZH3wHkH8iQE6IXXj6mzpq5Xpx8T6EUSmhtgeuICwzRHIe4XObmVwtaHYRbIv+q3
/CYwwIEJz0i3bznoamDATPi2SpJILhPGbIQoITlVHa2DKAiY9jKjGEax8KWKmFuoY83xjNKzr6Kc
+qz0iIoiaykpm7GU2mWOm3xEpOVw2k8i1pjpU18z5zpN+UstwL5a4BcxHhw9jZAqzf9cZjw/gNat
isQVG3fWSRptbEma6vKCLr5G3uuq8PAr/DTGBpynPe6f4QNyGOdBECLSwi5haN5++TWel8CpDDXT
dsX+MzCE2nYDUmGrjz/W9jMbE/4n12mw2NY2d7gi9BfjhtSW9qaIw0drdyhCD16a7Tdjd21Uludn
oEBea1yiaBXCLdQUIJhHmla86I/OBZAV9NYuqBLtHMx0soka7+5kuf+ZvNyTQLAJl37ZgnfFJWzr
ouvuY+0sojAXX+0jqHgMfFeobF769AH1QYsJByv9WSCgHuR/QZhQQSnI+xSdLN4nKzlUg4xC8dTk
tlbNL9Kh5W9yl+RBM7w/g20e/euMiJRHKlA/J1T5G/MMRVNofGMm4rZjCjdbC7xLeJaW3ohTnPPl
nv2pX/opHyl1oogyIYf/dZkz2yDpTul8JNbd3beV0/qQbcjFMmCKY1Un9D0okFZkfOEolF2TAynt
wKbnFq41H/KY250FZQGVWH2aM+Zb28oENyNhefTh+qCsFEfwA+8VQ7313jzYt56rcYTEu/9lez6b
CpuiuXIUSyTRTiGXmJ13X4Qo/FMbWXuewVil8mEHQr40OzgOGMOBnj6YmfQSNZ5JQxBjjFaO8mqz
K8omZ2O2FU4/glOtwI2L/p+s7oxO56K1MQgj/kAPkkBSr4euNBa/6CJzx3sFfWJSN41BqQIuHWzL
oCZEw2uNTXv/6NOKVs+lh5n1XHs7/J2aWhDKzl2uLhVz+3Cna2zVtS3vDqRgxim7pGFLqZHssNnQ
PRmPk6vXl2P6JGCU+YNz39UO9jzA/Qepqqz2MY4VkHPUOOCp9iLWorLQlLtR314ER4jZ7EMx8OaT
CJWoCmSGACNKb6qbY6e7E+jtJ0CPlEdUAlsztfbObAMX8qt+u7Q4ojYvVJgCbXZcetBmIMdY39W/
Db3aTIZs1dGL4L03M2WBkJjoSS2UCHLUMDo1ibeKOGmcNuuV1w1rcjNXXSL3GhLrIw02yn1YI1Qj
365qRLAAUzndA5pi853gHjyyemjLNGUfFcvNYTIJxqLaM3mC3osGLuvhyx2RgN8hulWTgtpjyoL3
EoIDJ+t39pr4UUeCLtFjQhT73Z/ld+2Ko3cPBtY7R0bOn5EIBkUL7Jsr2rYzUoL2iEqtj7YJ0uiP
R5/86i5yYdWHpikzPx/FGg76bUW0eJ/7Np6kfWYjdgRN3EkByWUWC8N7MUhdZjQEmhR7DtLFqO77
p4pTzJDh3zwCOMi2hBUqppNp9Vmr1A/7WhQ7b6s7f2SOjzDdBnqVDS9A0W9sLzmzzAjhMFmrGiQH
xEm9LwF1GXEjo3+PxSYzhcDC9ahp/POgZRtwMvHscRDxr5bv+d/inv/6E9z38RkgagGwtAkX4ytR
I1o96suMJiYEUvS0JsIXChWQLv/wbG+XzNlcLyfxp/1xRjmHo3GuyCJ2Hu6wJkSCR0THuy1a21wk
0DuGJs/Sb9NCp+50k72v55C0xk6rc44X5aO9PD1Dj5hxOihWTltCm5U8w8lkGH+C9f0wBUsvnhSC
1LFKQGWXYFpFLHPMYz+ohjF1Wv+JWzD2lXcGs2gMVo2Nm8TcKBvlfnyLR8niZ7bkdurXpDy1gFs+
tk/HK0ZKugcAcX7InTpfNt9YsyUYRpJJG62MF6ekIwU6lsymOQmKM2vBBcM2NF6+6oZvZWXgBEkI
KqWIjyUu/3O97yWNLpFgMfaGmIrGcLm8ScmBFMfh50UHo6j2H+lj3dl3r98hI05a4NScML4c4xYK
iix9uXZGPw15vfAdkmkYJD+XeM6jZlQr4nj9VdJGznp71nJxWSDsugbIavLQ2dtqyZ/bAymPvpgB
ImBgd/hQmT43g3ASiLRCJraaEw23xD/7IYsXYSxe7A1bPuBhtFyKUX6q4e5em9HIQQwWy0ORxCDB
UeRsRjW7DKqAY3M2I/My/vpbMrvxt18KE+j2FMlBi0iX9FpoEawSsKp6S/5AlLeYArp0RqUJxIFl
d/evupSE5JU5WrKpi+dvooSmoIvpfUYHGpc03GO8cNbzgvTwuNzZgyd/ZkZcqz6Skmcl7agud6Io
NigpLtsQKnu//fLhpMEIte2OAT/7aJ5VJ9NeQK/mBzS4KgZ6nNkUlwkdMfvR+xvM+hDVzTVF/U/S
aGp5tAMUumRvpnc7RdxKBugxfWKwMNNPUMdEhuKw5TbriaclYp+EF2d+NUBUj11Uw+xxJLpz/IRy
mDBf+sw53GfzQQHKZwZuzEbxRQ+5d8oXLS7xuME27xeu6ADLmiLRzzgzSogRmT1mrCtadEIgL0Ra
NG3dWIhKps7gsiCOj9HJtafGFgGKJJsfsZo+o70Un7UlQescZP/jyDJaJzzw5+WKX0BCrFHWlruy
01qVo8ZcIJxq1okBU9KaflC6APPO/hbixy4t1k8Cz5J8xK/pPIr9AdftGTg7eC0b0C/wwXQQQwEN
h5ZRV0kslVytJAL638N/5+v4m63+rrZqvW0o/cgvb4taiOlflOnoLGl//wlJe+NlKiPRomgCN776
F35FdF5XJFcTBEHhQAHGms5N3A508Ici/wPTi30kWLWgb9NGvRqqTtqOzRvA79JxsvbFTDVJoQ0g
la4BWb8Efov6AkN3aBisb9CUVHD+Eg1DZMbERFYncUrEKhz5Qi6flTP/KWgGuUhZVEjja1PLfzV9
VXqph3WSPl/+jaa2XCyZmzKCdHQu4G+VmPlJzhu3PhioMTAKaLkTEuB3gj5ZmV+VxfKv6QaC0Qzx
w2mB0X6Ije3jBG25bkbrDxNN07rmA4NdhHd9YWri7GzBxIraAVYp3Lz6EPhmy4cDOmvyFZ6LBEPv
H0euoaknuHFh1T3JLRGCUsAPck5G2DNMY8O7bk4Jq2+yTt22k+qCryT7HwQ/uT5JbfgpL0kOL0Z0
94f0R39QigD9vxQevHFS1potXQV9oizD+J5tbZY+YNqI5ZRapV43FHeyqkvCRrYcquLolvyOizqI
L/Iv/CpIKp0Zk+oNm6Pw3c33KVsmZl0ZN1oOkq4BhOsiyy6T/Yfn7eRSfeTL88SuStRRBrFVhaNf
EI8UW6UKqv/S7SbANkX7Gx0OTGS0yscU9I6TXYIbLKDV6O1ots+tnEO9PgXRWyWcd90PWxj/EEMR
0yeQLQyFWkW5UJQI/N6ONkdiXvc/hk+CRELMGZ7O0urXZpLLUOlx6FLO5MiFJmkKWpeqlU6tF88r
YVCqWP5TEEWd+FTkbfdBox5BpspvyReUTH10LvP+l3VuMPlUSCAyeibAelaQ5zC6Psh5H1nHZ3SG
R+BkyoiFXnomgtTNr+otGA2jIec5mBzzjstTaR6X3Z/RUXsgM8JyBaNuVCub3Xts1mPXXr1YpC7r
YPoEiYypAIB1GsPgG5ifWzR2lb7FCMB3fuMx7LhTGzEKveOzbBNiqVKICGE/GL08FxPaGqJU7j2i
wT9dxwOtqFbjnXQ7R85UNrJ7i0IOKwuChhB+VQ1+KtCdOHAiaPwcTCl02vD2Sw1FvGT9n3M0Nmv9
NMFdezSkLyUG929s626hFlnRqiMdEaUOZja9fKqSDPM0pzIZF/zf7YKi10bwEQLMQ4omITuobqVK
DELbxi+3rBqeiXPdPIEvpaBeom3QUkxiyT52Nh2Zp9SmLR7lsxNblvDFjq1Qw2WW9pWMopXQjD4r
HiEKG9bgqAe9JRn9cbNW5C5xrpWuUjyPvQsS1LtI5zyBF3OvCwN7Z8GQttWBxihHPkpIJgwOefk+
hp8e4eSm4ARtCxqGDxLdHvTvO6ZhwulVFSmAQK1H0zKymxOUkTtacv9XYwC05bx2WtCESbwCAUGc
zcUcHLyV2Np48/J45lLPIESGtAJcegU5rDy5llTdRCBQI9sbMR8sg/nf/dlxTdDpBWkRjNX+ikB9
Ky6yPE3AqimqfSHx3RIanOXpJE1CSaN8gRroSF7gQTBJqWvIMgRetrBIkoq2ORdM4gLRJQSKEofc
NHEcZl4FtZHwcUD+
`protect end_protected
