--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   duplicate
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
DJOpRwcSc1pqt/j75WDZER4Q6cJ/1xwmRTQSU+9TrBSIVgWnhEw86HnwxOktMmkVRK86gI7EbaAZ
EamRgYDH8SbS5gUZ+x8C37haHoKe9XWDktF0qOtX3owzLsBQ0JMVTBNZPFVoOXgnCHbot97SDstv
S6eDQTeQxrzI43JdyIzMnVyiPSaz44AcHg4bowdmQ1QffPqBa6eKVYsl+T16zA8h/oUjf3bLctAm
ugMCeiDmF+2Cm4CKcv4sLT1/fPw33xjoSrpimAqpALO8OpHuSTi4iFnPgGoS7N0wV7yJ1F5k4rqK
eTJRuyVtS//5qDebdFNlFXBRYPxtrrmKrNGTWw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Pssdt6QwmFgfDRm7+MlSYb3Vpw6gPzO5JgY1vo/jDts="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
iIJ7vTfTG6Uhgwt2Hpvry7YVa3rqlHBG3DjQuHeqk9wQJxc1xpyIzA8lPUrSEwz0+mIPQ1bMwfoH
XjFC7wICiBu8qlwQY9E3CwdabKjjQtrSanv9WsJtZPI+MSvaBPjn3SxSKTOBpjvsEXTtm5jPRDqz
G1SyX8sogq7LjJQaycZ3TcXzwdATbYuge2wzMrC8Y52ld1Cmjk1z2EkQk5ZzRWrQpXDofe2V7qqI
x2PnwPpgxEGbYdbrmnKu5DVGMwZ/rLOkIafmYr+AtYA1eFCHIZCmRWm75pp4kDKVglOXsUZHGz6z
TD3knoRzjfUy4OnPyfx23hlEw6GwFpq7WLW23Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="iwCJRNwYYciNM7CTgBc0BHmjimUx8YSoL1ns1oO0CtI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22544)
`protect data_block
jkgiLkxcuGc/1XSYqjsVKTWWBkf3eD/0vp9lK6mYiXRkFozoTUSmKkbz/B05lbEmWWAnrIqO06Zr
CD69pVkLS+Tmd1f9om6WLyd3cypnmiVzjDY0wnKW1sxbsmINdCsuzVReks+CpA0L8E6U7FYpG8Vf
VWGj28e4v0456gtzpyvu9HkUc7JxN5i0GRD9Q0q1HL4YI+4vP9h73HM/vfjrSPNWa/ypjw72mQcM
K92FtgwtugQ4/m/00u6UqilKbaAI8bJh/kGhH0/oAdqHq5clHb+7L6ffWf3ln/siEtQ6O/uJebLM
JDr52YDvHUpWolWDLpDAJj8vm0dckJcwpvuhnapYVsjXjbDfL8Bij8nWMu4oZjdTM68PO0sCc2O0
/1CRac1QjiIwo5lY66twCApJp2eXZ/TU+ac8+r1jY0TkiO9NpyWFR18b1sPlIy2gcuu9V6tgweat
R/a6HkbVcnC5BRE3lWbX6jzCWaEm3HTQMBcMC81BEk6YGvTSq6YATWPEKOFb5XndSmpVqrh4LDYZ
V/JGNGcjH8GjPbN6vrqajfzSLpry80bcl5euI/cyGBl3oPucM40cVUPIepljTw7EScAcnSLjaxnY
HxJcWGdbLzuYeToDzGtY4xaXj+T6rZYc9rO8dIxkn+jnRPDX3670R9ih37CJWQtNXaBTB0CeFIPN
DXn/xE4rnPPNK+lrw2NlLfkSq63H95FvD2Vgc7Yur93ZRlmBQoZMBw/JhN7S9wt1F3XZ2x/9pIdH
6WwVycYYtq6KUfZIGZwD9XuN1MaUbqo0mb7uHlyQr7NvR8hvDETyPNUeinqDQ+3NaqCHR7h9j8Rr
mUuDVvQzMQmmlh7k4lOjvFsQtJHrmvf+Z1FwlXjQY8S2qAGSQW8KUnNTdwQhppD/TUo0mbVqLsu0
NrEYFEqHk/7ftRPuU05yKHj5uNCfuJpeuFCtXPvKp0rqHE3VoFa1ty2Gkp6x0NWTB6xGU0RxiW5n
vlV39skLXAoyYbggs1kx3NmPWKkStz4qEIy0swg+t4ElAtKyQ/2T73ENIP3UTzudnpG2/LzAMlE5
7ksY/vIL0UOyX1HdC2Ami4oZy4FON1s64qyQIlDf7HnVOPyzemApECMDvqTOdtAm1aZfztblete6
NUEeODa9Aij1Gf1/hlEcBaQDqbK8HNaNeMlFhPeWF02huHgJlbtclGuuRqTKztLLMmeMBQD2e0ru
AQQksy6G4BMm++rDojVDF/VCE8DFF3MDH/I7O9ep2SVj+xI/vhK/go7HIYJTUKom28Fft0NieHAe
4yBCUMWVJa6BSFSiICrHiDbDRqr0pp8uj5AkRhkLTqkDmeft3WE2mQxuBS/yhyOdRGyLscXvESxX
iOC/SiyLui0EYa/Bi25mr3GQg7A4v9TI2ZZvmEjdY51w+qZNC9lDns5oimwsVhsJ8ZVq1CsDFC7P
k/Qa4VKpa2zZCOQ0pKHXPpnVMbFwoyM4jU6Bc0WskiLJmkyoO1RbzDnw1wTLBkT6Wv+gTdvYNxwu
i0KPa6PZkI20eIuV4TdGL3dF8wqSDHEUFaS7f6V44mpXdIkUIlzXUYy/zSCgjK3vskEhxQ++mJ/7
+BRgE+okuk2Cy8CGF5ce1DQ1ZV/OeTqXgRJEV1ek8SDQFtpykcU94so7Hu3xdAbhaTnhNIluAFQN
FBGBPd0cJbN9bBMyPysrT7vTUgQqJpUBmKVjVWglELcfxoLruitbFyixcP+TexWPkvL+5OJ35cL1
164Gk5BqcZEKXAoCTwEggZr3OfPTzBKyKbk9n71VJ3VM4unYbD3yJFLFhdos0eYgXShM/vu41ke2
iHV/5SkThyAcfVBUwp/I2lRGJojOdUip6dcZmXcVXsUEnO33taLyyJf3R4nFNBcQg2jXh7tPP1KJ
CRUIdNeKIqhcuGE7xF967VBm2SKe1dCA0W4WXlH0/RTra2DxJpEqeTWZTdDWLJxIxoGi/lKw/U+7
1yVPkNNwXZXmUICikpAsENmG28JCy7q8yKS8VmgDt8ryDF7C6Lq/yQghdVE2ap34bUy9NMF3JeHK
7Kpu91HGvEstYs0v0Z18O3zdagWF9xc4zLRynpMqxRpQTk9K+OQpy+seL+3mS/PQ1xPK+9cDBAnW
Mjzu0MSeu2yoITzT8pgZlOJNvDa9NfOyODaeuihJs/CHFyOVodr9YJoYWkuW8W6+Wp3OtMdmLL7s
J6DJSA2q9aEBOvARENFtwLDxSHk9JiJleGocXcZkBDjmLZXdy8KqlR5i5syK1xM6tkBFXPFPUwyU
W0sbkXS5sUNudgc4mw6laoB7QNICb/OCQ3/xh3Wm61z8PSd5XzAMKLQ386zNQuZr2jgiDUk3lpOs
SDVL4zmsevMLV735h9hBfSIWwlBm6e8ru8RArUOkirL8rP6OKdFKL5h0A1Nr01r0i+IGfwJqQ2dr
50KXWaXpXwpvj2T5aj+FN8PvRXTRRxZ+PnLoiRWGYy7b0IWbQ0Z7oV2mtIbXX+PhIqVRnN78y6qk
4LIRmKnEg3l9d68afR0Bl/MifRKs8e3X3sulWdEYv3ABfoNmr9rOAJI26slKWrmxnxnmDEwvLYfg
uID9hTVea5LRCnxGIdmb3z1ALbvVFhM5ItsMJx2zDo1FlQGZq/I3veS26hdVpHzfU6qh2IarzZy3
CHCCZMR6cDR4NBjLOJyMVNqYX00gXoy6JpMxwIvmNIU8gWZqD/50PpNlsK6X38Bh21+MBGbJ8tGW
G2w1y0R16DFZHO+4EXgzkCP+FktaskqoXy7XqL2bmukH8Ly+Sj0q4QuFpgIv2MyMNSSb1hv6uYHW
SSgJ5i7MIDj67F1q4rvsbRJRqThjn1o+7j5eLXgMWS+Bv+eIY8TQ0QCDpA3L3mpYA9jzWrJghvf0
XG3b48Aj+hNcEnPvbcxrU3VB9d5N3Pru3ZO22MvKLDRGJWnPchNxmXDnK97qjSetPwyIQtEcPlrC
U8x+0lKRQZ5WoowM4zfEenurW/jojBOxAxNH/LFmTx9vIw/s75X72ARLmUAdq75/6Rn8yzHU7nXt
Zw7W/K+Oy0Wt7kJB626gumf0S9rYluBG1eDkofGXor0QFmH27oOBujSOUwnKDwsTEbNsfcmcNsLN
RPKjyjXTNW2bC5apYJdXUCdjbxvIFIpcuzNUrMMBQcdocYgmLV+jqqiKVmqIdKmHg5JgBq7MkfJA
gpLHSysVsoFRwPcGiyUPCDZgv7jyCV03lkcnS46Xn+eI7kOlPbjVkGYP7b2KpKVh6R8l05NtWRxs
TmL+bCSHrPSaM682ApVDzsIW2jP4k8xsGq1faKVIXM/KS/AQPBbXKFXlVmmLum6l4pn1QORYj92r
vet4amw6OdOjhLsjc5S//Iyx7pvxwDuKq/C2VJir5c0W+vjos56rXHQ4QAJBX/uF1hgFqmRtoHSE
fd6tHtLeCRsCggol/xEBp2KWV7U/bgV6252meisjwQMAPNMyrTlNTWaIjmQ/JLOgOeeQpj1JtoLo
Wp1VucCmGfsBXvgKrHMG/JOxCQcWpd7EVPTJj3jnOmFm2Hsr/N+9gWlooQPH+Ij4V1TjS++W8BBT
v9DefkSyn0oJJpNQU3UKwu4FrpMbVr7QM1uUNXDPAFEZa/iE22so38W9GPPEf/7fq9uDUWLwx89h
U7w8aERJ8MeLBVE1Qhav4PNVGCh/HTmlJ/vim0NisdAcBL306/hF9Z3Dg9A80NGr+xZw8VMmuOIQ
FG6TJ1q/io10ek7DVRZAX336Tf8YfX1HDuPYangwzznOsdDGRVVatDNriDOYNrQSBU0A5m6H7nan
v7TqcyIyWdVWgiMoLhSZyvqKohZk2XM5+Z6RAfxfyJMoMlIYcmTc1HhDclfkbJ6EQpaQqIXHy9cY
4vfsv+NBaW6wc4DXDCnHp9Pth07UVXdpEGqqI4g199/OS2+6PxfMvuQZtzpICKS9wxK3SE0w3ayz
6CoRhZRvRGeqI83NW02KYXbeVNOtLtvGz54laMAd//qWH/jN6T7woQ+h1D9y9LvEQnI0dVBSHjXX
I8MF8Prdn/EczTa9ddm+J3JwElKl+sYGgk1n0Vw/AhV0+F1YWTep56jQt2sv9ULie9s7bQesEmYu
gUZyUvoIMEpyK9lU2oMj+raAKJ9eofQw/tU1VBFvZeQ6At4FKNzVb7Snj2lUMYwlMXBb4PItXTyf
jj9xuRPIwRJCHy8+miK3mYF2+qpsdMC5nCPHdTFJcWpNvCACJHZMD6rwKlWzj0xt03x2NNAd/hcs
kGuRg3u6ig31t18VAImiNOPOU4Sy7LPM1IX7a3/13QbHeWUEd2cSf7ST1jbUF/EuSKGLbRhMiYrZ
RTnplN00YRNIwIYfGJl5pNSfzI+CITeVtlCZG1r2kp4cgauFP89JDkE5rOn4UDWtJ7Kx1dF85V9r
/RL4GS7fKXVbjFirA/tHUVWkUugl8kVzC0KVFPsq4MijRnBEBfUlBmSKBTXp9tyT2czaDpJAeCKf
oDGEptPc35UNO+sKE7UDpzwj8b+I7BPB3CTB0mzm5suySJ8UfSgf3OO0i8WbbUriWabxSOeeIbMw
i3CulQ3xcszqUWo/P5NJCeTy//aXGCEvy6H4qHjBPbQ78hc4ryVAgWjmFBqh9Lgo1bQWjqq/cUI7
0IrpljuJJcIXGSxV4HGnEVHL3/r5FX+18ctUwYThxP6q7oKdbrt7AZGL9AoQm3CHgeYlVL1tOc1i
wBjebXf6LwPlOB1YLKzVnKkCl+L6CR+M6IBnjYUZs80c7M9r0bt6EiP/o8jUK9tmFFCZV+BWR5io
/S4ooDhhV+LhDisVBCSwlHjNx4Tb57CTDWO3UIQ1zcRBEZYGj+yp5MWSHGUVaSJ6dIvWhwgic4Ex
LveEI/dMY6jagjzBzzsLHMDfDt4K5w7ud6kmJiskJkFFDhgexp7bzZFpIYtFge0IjGc3zP0K7sV/
jydgZPA6jSM1ImQqnrxchmk37BdKuEkgVarL1VSnfS8luiiCEkzx0kpou3JbktmMTXsJWV/MDOw3
Yxj8B2YWtoWOKl4jKDbfJYG62QmsJqC5ZKHRPbmsUuEaKngNNS4Uwa1/pxa09XLIb0B6oI4fwkBn
mE95pplgZGhKhynsmjb4Aa74qKDJWkUN6tCDFsw/oRQilwryFwAQ1pbkmlPfe0c7Y3PO8kYoNEyf
eCm5ds117PmjlGBT9MPWvqEvdiGskYKyKe+MdwxsKqaJr1r/DaAQr310pbaX1fP/JEHlqXz3IGLn
2DcdwomBiHiRZDnMviOgKfyhc22Knbvs1KYi9qtYYTyo2d6zeTb5Cd10i3cJRLZ0zTUaa+uSETvW
EuptCxgSzvC+imO7LhU7/rTqYxQeSXooKz9ruDD6MmXbwj7kApDIpAtACsTcj5jAfoC2ptDu0S0i
rERQuHOcxnhuM/0oNa4EKefeIZpUb00679vgoMFR0yPsapWa2GOdZGWIZEMclnnzDEOa0hse/i9G
7/kiCakChf4omSgVC0r3dbbbR5Os8kNX7m8KF6ymDRPiwjYmGlJqEsVrMWKSo4TYbFYxL8udnXuD
y65yKK1VgdK4G5TMTuugdYspDUoYnepIKlqebOIH8TGSi1pB1M5mToah0Euagnx4C63zr7bqxpSs
jZgmhYvtVmOm5Fwe+N0yDnXuwejsZTlHWwNLjDoj5j3gZBiOuS+prBMrATuMOMIDP3hiltVcfIUy
SjRcpzhbuajQnyP7ab4nAkWIP3GEQAvs/k9FQ0DxMivOWPUS2xN2n5n1BsCt3Kur61gkOXiOFD/P
I2c6HfJ0EuBDEhtxYGh0W3PNhCM3L/nHVHnppvK7c/mBV+Idbt2siu9oc6VnSKtbHAwHeAICyAbA
YcJz75fTgvyNS8wAqtL+pig4b6SuSea7askd5FEn7DdQkbq2u0tNKRRQeU/c1v8TXuEFxDf+lYA/
KxEMJ9wMt5hcQMkCXXK6SCDNRytAWbn5mQviL9VkhFsK3Y5GStzNe+WXckN8X/vWE2aLV5UZlfOa
UFhErwb/fh10tMXkmsvMyUkjMc9uZ4Eo/KyMc+LqnU0oqaOlZNqfOIYcvwff3Ei6dbqK2xvbZUWy
+lcu/6HnlXcIUx1umD2hslb4Z4psZ0WwBLr9aa019t2tApYiAR2EbqLaJhyBuCk1H4Hih9K6DaQX
8qcwQ3aU85YZ+9yHH9l2yPU2B7W8aipxYmcTTBv20Ma2vk7SI1Y5YdZnZrA/vjRR82lt4JBlVBmP
AkrCr01b+uxI+BtcovkHwDYsRhLThmvtGLnEdgOFIipQ5YXSm23qYijfi8lmPZlWhIa07KSEeTRa
b9CeKC3apBIjCgKvK+2UwdQ5s07jIzK1tufLUxO1X+LTjJlyLEpd/Qddq/npFJ+CqNSSnQkDfXWy
MNB1t8lM7/3vX+IbfBFL7xet97QJg39hyqNksRrPcenGrBX9GuQ1EJH1dvURqGEOSauTHPAR5hMJ
3aKKDdcnOviV8h57Y9cUGbmlMx/DlvOh9rKn4ipbzGGRyiy8LcaS83F3dDeC7FqiheqWyZlM66AV
q3fEPFmJr3vAsgaHhd8p8k319wzhQ214FRlBrzwEwpBz+mpsXC3uIlK31+QUq06TGhyUTlgYyEJ8
dG3q6SlyLt7ND39ZnUSt32cmJz8fxRIyXUfW9Cdn8kx75GJUwyT+ldj+GExT1WFErEw9HYV6ohBe
AJCq7UqoV7wLXjwEzAkFZ8VbVrLEq2ygeErTEoBM2f7NitTO4dd25Zofks9MDbAXve+Py4Zwuge7
p3NOfMyLW35Rji/g39mEYWW3+L2Up+JDCIDjUhLPdZDtXGOcuURhkTFtJ4QhATvQu1P+ukCGFwBN
OOZzjuHIHtgpRecZM8AkdemfOzdqNli9xIK+hdQMAauKILpTmAFa58X1AFm/e2+PWuuRCHyipZwk
MYGvvV5vFEictrWGlDPEaQ+im8se2f648BVE1UNTmyGQ3Kw5si+PmD4oWkVepfPBWAD2h3rGHKO9
IHi+sMHIro4Tn+BBhkZeW/mV7IdyxK5AFmlCnlqyyfQPHhsWBHbqAelPx3hsj3bUU5YxwY9ypKCp
rdKTDZEgqYbSg1LTSMoh1VQWVcIVKw4q6iO+E+u2+78IAhdwr0kIQSL9/KOc3U2w69Mj+6hFRy0+
E4ku3iH3wp82/h3HgXJHkOGtyJDjZKaVGSnnFO92kR/fqpaO85YWAUMKruHuOARP5c0L85gwqbf+
PJWv4C9PnDo+NIxqFJjsr1PZOF3PONMzyTGp02KkNy0BGtGpRrNFFqTn6bhv78RUCdjfimmXlGaB
vfYkRFWxEB3fh/Q1j2g+qCGDKy2JY/TWRSQFlCf8VvZhrd7rF45IQfuHRzK0hxEgtNHzuFaYKxCA
vX48VSRO1c27ZB8e3gjcFUpENsJTHy7PUY0oC5qEod4YpYF5Rkvnd/H/yAhRi3jaNMpamtrFv9sg
41NAplcrQfZX1GUpJO1L98g63zccED8eNKN1+bqY0oAOo23ihqq2DQym9GFaA1SxmFCROZhScGqQ
XUCvLpcjcwLz96Yp9x5N0LAEVnQFefY3HIaepjCxjNM+nkBMYMm4zqWZVNMJAubJdlZyC6quHFi/
IySPFEwR//21UCZG+BQ7ZmVsSEqgjOB/YNS9196uxJeZ8VwuwZ0rErblEtHiRZH1zB4M4VIVEJG6
bkDwO8Zc945/4k+JyvuPYVHhh557DDbr15hHLTArDNNB6ToSfIjUE82fTIH3cpDXeiRaoGtcu0vn
SWDQVgznbKVWCLo5STSKwnVwQd3ktQ+yFL/AjiJwlcFc8h6l2A0RG/GrIldg6NsRBILdgGaRGr2p
vewOkcpf/PE01CCB9YXleM4Moj4xnirymhjPuhxbdQuODd289iFVG///rddhr351UZEEgkkTG62A
lORpM/iPxCgH0YcyZmnUjaoZYteyyE4LkdCii/PZkBZFSkq6BtAw6QvxfsDiPpRQrX5OkPWZU8XY
V6Gty4g5a/flCUeiaEHtEf2eb+J2TbS/BFa2FOnzEO6FGZhrLvnJk4vRUvdv3N2TNbt0MjK4SAn4
Wczzf1fMLsFsWkVRkNj1HoW2nhwEEQ6omtXU/KwGOhrU7HehSBVWW52j46CiF4bLzYGQSqFECsO+
OvhJuynHlCZsVR3up9ZEbhefb/dj2NOQvSM82g02msOY0Kin4T8mXM2pXku9wN6CjVbeHhZoi3bM
PBEaICSNdZFA58LSstRGr1ynSEgagjeoaOQvv+ytCSd+obpHPFTFkBKlBAJ4i4nyc0rOKAgNSkrW
tjMOFtroF4Ibnv/ejvz3DiIDbzqqQb1GjCgeqBJ1hCq9bCIhgnnNLaQvxH3YfbXO33AsuLRf0Ktl
SsVNnu5tzlSaRruWbyCgLtkCH47TnkeeaWVnTvIctsq2HP+R//p9dWcJjw5s/jYL1gxEN9rLdJwz
viA9XiHVAJaL/aUQBnMALC4RhfLzUWUrL91OHKEgAUv8mCP47acbvPBuK5mM0SGn11azjUjFqMgm
ODmYh9cSEet9ZN02DZXWBQBkJ7adaBFAGlF9qdiKNKjELjHwEghrek2iw2nQkYL4WLvqxXkRJA5J
EF9Ajbm1Yk6V84RgQ175VEQpxBAepBMAVyVHgJ2EPut8/ICtjjjoY5sfqo9e+Tjl5h0j57nTmoRP
o2xy0AdAbqqwMIda2wMcYrxA1oID8zX10MiH/Pc/PPBfPCZW4/N2HIXDxGBqqtS8yhfUqjRdrl6y
dvmel8FhBiuUWMxHLdZS4DqbLZuX7EmVbDBrvQcT7LIbm8SiOUIZmS4a1Pw3jCfSDdcgIxFMGeNa
vqi8JsZkWOkKBWwMJ8DaNXg0kFiVc5G54fLKPcfbkTzcvz9cOqiGToTgkm9oEI6jyFG+yv/ZA/HZ
zt16V1WuxSS8pLFi8FeBX74lELTw0utfIC6C0GBseqrI76ynh0sQjfoaz2NZRZnRaS5WQDpO651h
Hn6lirzN4HW2R7Ghxu5zUiftmY1mNmmxJV9KWs2ylA8guwsPJi98wRf1ndeyyCrncPJ9EU8dzUYK
n3cd7UOsL95Wkp/X39uGAa04NWlqiiUz0QC/UB6XYkVzfn44bcPvyTL7oe4OnJ10MwtI3NaeTDVR
MSYA+rb307T4Tbzqfeqt0l0w7kNi0No5n04x50YRHbGEg72iXFsGuZ384c2/Y29o+iCa5rXwDV/P
UtQwbcYiPt5NVWAOuHHn3QoPaYhJLj3FF35/TAYSwFlg6RRiEAA7E7L0D79WWQgu4bnCsVHdw0ls
9K1fZXl1IXyjMPUCbfEFwWRPgotKEjXX7XPilMgQzzrEhY5QuHoOru9Ezkr7CzR1W5WW8GVmN2MC
rS+qQGG/sSeFvDkFYIdYIPHl5CDehW9KQkCVcyd7/j5Gk3qZpNTVCHlued9LdtT4JWhtq9tJe8QI
MHPoWeATH2ej/x8Fc0GVTX7Bt4pZYcuqN5bpDLgPmnBqklX+R5ElBwHQebtRtSdhxCe2nRPDp7er
vZ8ej3vUWlAqKNK2s5Net3L+YRtnrzTmOXbNpamYDZQcPDZqqxjoszR+Nx467s165ICZ57KOEZKs
nZDKpa/iCo0yoQuLPiB9hbjcIl35R99WJin4zD9U7t5/LdsI6+QdM0HqF2IUArPrgqTvi+kqcFQe
VS8Q7crhnYrQPgzNfhPgzsI24dcI42gcqZe0DVoh11rWMTq5xIIRPHhgnHMUaclvlZbFgZoKHyqe
RaqkYE8pT2WIMo80KUk9AmTz0IzhjVr9WsTKt1JKPOyjyqvB0SInNTwwgnG3mEvLA4ncXVuoLsPu
0YomZc7EMEQDwnrDhIyrywpSeroZ/tAbovxAqASYHRVIJBxE/BrJJG48seiWJzzo4ocBdfNvD4w2
5r/94Z6/eZ1tzR0v9tg5/Mpfk3guvf+yKpxRi8+VfcqeX3lxju2AWrqBvJzD2wX0uVNl8sPKTdkB
Qj7xHVCbZY/9HWI+pYWz+05mKe/5N5yTo62FWz7YqWxDlwd4k2XzBG/77xb1HHTEYawYdvUbxfIq
eZODvd1Bos98fD1A5A8kpDsfqgPvuJ6JcIghLgoNfBPjzaNsDSqVMytWl/5cd4STw5waUJK2Hi3r
Agcag9ZI/a+sxMlnov3/6i2rhNlhj8w0g8ZKx0igHRa4X8B40T7j+exfwBfY0XJ5zPOWs6NCsElt
ssQo0/AE74bWIWOPBrbS3Rsew/aO1o8PduBRLNPJeuaimEr92htLTkkqec+VPPfId57hxt+8Y2/l
hxs2uSEF9a/lQhr5bKYLD7umf1bk2CCmaL3cfA1CTZu+s7+4kBPe0R1DUPtPuHul3AeP4KUAx0ZO
52iloNHgR/43S69B42r9R5A4/nJ0vvC9zSSUylV3DinfaOmPgUVQEzirU0Us30e1QveLYzGnflAj
IZtv0ptZD4fb63yofMZIh5tBZOxTkaqK5c0hKAZtZbhMuTQCq7N/NKBCU7U9yFvZugPrP+b7Gys5
UXv6IREruu2N22JcpNWFgA/adL3ucqyY/oxxOTViWdUixG0DOFvDduJAML7WdJtuMdi2AE2JGvF8
fSoZaJxmOlLaPITHJlFWBKfEBk/1sTlN8VK5bRD5pjtMzm5HcFLV77p+MGn3VUVJ5R92TV6Xtxg7
lfNsm5pluHNvo98pG3RL1FfwAJCIkXypwDkGCQrMmWawZNd5INPlf7iVrwBP7cTctjWDU9C4tBKk
7nr3bS8n6K+ZNPMN0TolrEOWkY4GWZ3VpgC0d7YtQc3HQc5k3CGEP5Wx3mKocqSVBuAcWIew1n2Q
N6yzKzXcUAI/dC51YqwJlKqZhVEGZqlMCKSSTR0kJx7hahxCcSMPRIyAoI4qL8S4HuxK5Gc8jjrR
JcHIdLsVCdj+of5jULMJVUiu+3g06B5vs+rRBsIcO3s4NjY6AjrkGcajJme2bEDaY3nV0P6WbzKF
Hd9g5Ru/bvp3xkbg53wZ/oDISxmQdciV2s0zPjrIEBRfc9VwLD/rz9iQzFwMzExmepFNRwk0wQow
j19PW4yjjm7fl6+2K8x6l9/o+Tgzt+aaI9E7CmfuwJd4P9t3zm+SspDQkX6BLIPHzUCYzSB98gyr
LmRA01g1gfAbJmQ3bgZvYvzHgCzm9SbtLAv17EKv/aUlPG9wjQgaxWB8ht0FMnkubUGY42Z+NtDs
EJvz5tlBWXY2Ui6NEJVqGI5MF/NOW+07+IfZgMhvQ08PZnoF1sxGE4v99TrXFlzAM+glwCjd8mst
xBD96kmwHOr5MgHBjZShLLwxjpIPJANPl+lsApGZ+DmMEE0VyeaKWDYPa79f8bkg1NURqNyge3fl
FsMsWOgm0CdtMFC+4Q0O2s4xkbesmcF5TOXMRUDYKybo1yxfCzIWn0oNdKZCMirUpUfagZCedEoC
hOBGsMAOM87hiojSJb21+yZTSXwCdHQGoULU84QflJgd1Ghd/Zr5cXOE+q3T0lub7tuXtDkOkHZ4
xH1gvKWyqgK03oxS5ynoMeeM+DKZ9/PJEbhaRPLk223KAYs1LojHdESiV730INm980dvWj4hlC06
VnEYLvGFxGlwpgw7Bl+RrvXXdD+3i+u9kn9fYU5KrRCL4wPOXweXf/QXRE+lna+UzeQWi1pHeJQz
u6FQOpzfwu/8zux4ER3JIzQ/zl/1dYv1Yk+l4B3NtrtbkRrKB5mWiHH62K1+oTzHuo48mC3efOlz
qQDaCq9Gvvgvm4KkwEiJH71SrFZQsi/TOTHQTSJU+jCgaEWABE1bG6INpGCEwP+0OhDDV/++FCbG
6FCb7v1Tck0QfY7Bq9lf5GZ/3IcS3usBB9QUqcr6XAJVrwOVtDgCWgxud7hKLzOyz1xFVh/WC2qP
h+mzxP7qcFYdS6rbNQm7X5/5hqpi5JkfKrnIAMaEQ20vnY4SkE2y5Cc5Ops6U7fnsAptn4HvYjbI
6/2ZDnro+16GQCauDo3WU9USF1R0/wwDcSOq1t6BUdmdiCJ2UoMEAYYfrbzdtCQkX2dTC2K/PbzG
Hlnw2Oh2i+/2fy5tLeVtRja+4TToYCuOqeeZ9dosh+r3ZkGXG9gOshReoai8Y99mT8DHrWwZIUKI
r5zRQIg1QhtkC7LOJRT/EWM33jEJ8Ie5VAR7tcfhvkPgAF0zaozHYM8iId6Tp2K6ktZtwC7PSpng
FInPwacfV8DTHW5zSKfXilR6swdvzvg0pqtBP50QmKaSTrNFgCZLBMrlbl0Q9E0twLof9CMKHxv+
3XHiPKXiQYjrYoOoewHwj5Ytb6O4fXjT1xytd6mzw2j9tcZaAzvMCGgQMpSr2O29p/0eeLnzi4uJ
MQUCA2CT5evmlO6esEBga4efDCm6MVb+nrg+7x4GbAODfmbq6WWTK7HGWnUo6jVDPzDqzsu+rRZX
RHrwzuTTNbpBjAtExjKVyA7rgpFi09iXaA9i1htFlwTaT44nYcUmrcqIESxCd+69BmD9kDV+Znd2
26PlnqW4JSsT9V5UYn6spySVQWbM8Q8SqDdZiWf78PHOuEFX+HaztFJBcPuIddLmGpZcGgxgvuDb
zKe+RUZorm6qdF8rzHuvozeVjj8xJDKGWxmWwwfws7NM9nlXl91yovqFi9g+8cCBKva0936loTXz
aYvtANA+RoaObAVGMQzUTsxSbwjP4ZpvXxMSMy3ztTYU7EnMABAn71YKGcLG/7OQAdVKFeAFhGpb
YxC+usEWwQGl1A4Uwe/ynt8AtUXXGD2xJkP8FGyvRzRiiFFsNHb2Gb5LdUjkbTreOKGYotI0dThx
cQ4e66KTI+9piidCvBNwr3k6DKVM6JFsLpAxLzJwmG6CMn5Ge6vbmiHYZYSCFTlPusdAzMfh1OTY
vD1BESwsxdLCxKUXxfARabrS6ImL1P0LXokWctCH/rAgjnV98uAmjzE6a/wtuvwiS2AlxAvFTyr2
ZagSQPcayWIW2zlFit7zzscz0pMmGPItRA8YwyD/jpBd0eEu12q0o8s68mNcFWefFe2MEYjqAhK0
mfuVmVowD4plajCHGComZ1DrRa8Wto9BtJ7NQKNgpv/c66wI0QICTZjQCxg+OfERiX127QvTy5oZ
l4Z9tEaPe8gdXM/jc7TPzYm0DkaBt2sK5Fl2rK38W4MSRyOOJNjn0C6Lic9e+muO8oyB80e282b1
aogwuuWqkhqHAqtuq9AK0rrQdclAQb/I/JLKTa1IctnzNgMfHO4L1BMNTs/8GuEZhQbso5r9R50G
apGoUW0n7TzI0/gdBRQZ5//pYgimz04oKOKA+jEMVSD/1+R0wOHCUhYVK2D6PXQdWZ4MeRE0dCdw
3OVHff4c3GqqnADev7i7bL5LJSeMEX5B74R8VjShfVxaBfCACHUbbp4l/2ZnDNkT0+1J7d1B3/qr
941IOywyUSxMOkyhMQbGhXlAKIuXRkCKmTayJXatwYq/QszBRCHq7umVoX+9/IL+mivBIfFcJIgP
h8LSTvv7ooBb0EljjEeaNxkWOAzz0g8YEsbzzfTwf9RtaOvu+VdM/7gujFFeqbWBKMeWrURzytaD
KQiN3CsWy3uNE6lyu6v22cULEHelxCD2KtSuYBfgrm7fp6q9VYBrXyh7ykMEgyi6IfLbYRf/aL9R
OhZSYyX7ofv9x7nR4WPQUNMoETDDfpOnp8vdto4K6xOSZ2pXa8TvX2vaKyiR80glh3oaF98Say9S
JJf3lwzA/MeZiUKl4Wf7okZgfPrPgENz0Hk3iGhGnHUXatYfZUc8Nj+YuJlutYDfrOPt5CdF6lJg
W0E/D8CtGJBcteuCHM19xD+mbK/m/Xi5sPxAzXH0dEWXQsDXPDpn8bBWXsv3gXRtFK0n5BFxxJ0S
Qc2+bCTk4vaFgYxxs+l3scAvT/id5j/ZjFA8yc4JLpUSIFnAMko1xftaSzeoSqp3ZuXldQ+yOeWg
Yy9AHXgNAXoSgHrDwZ4TheLpJVO7xyvHER5LKFvLZ4lvoB/VCeUS6F1DW4A4+/gMch4ottILGnsE
FOvf5VtCh3Pq9ljuX1a21dGgC8aniXoPB7RHe2cYuLE5pfN8b4SQXGo3BA7vfTFnVa4Vx2dzTVif
zCdWfFh2DkfpLP99FDlmouN+/w5Dh7q4QPbBIIettj2gFCCQGQZ2M1V1kdyPwHpN35IVY2UvMoFB
U6YG4pvrPLOBhEDVIlo8VMVFbboSMaBh9cvdiBDWpCdMqi16YJg3SJNBf8l6VXOI9D+dWCr8yjbf
rHE7/aZrbwIHlRco9Tvmp3nYrNTjXCkgxFtkDEAhasGNdlaUyjsHiBHMBEZ5/UWE88aZZX2ctBKG
XQNoBo0bM3TTL3gxp4kMp5/C1+T7kpb6EPqxO3Mcd2k/9RQMQ9sUYjupB9JTuEpI8Slf1JqKjvdl
4I1Fh0FID10TgSmTb9uaXraKb9bXxoVaed2/f67nAq+N+v7NTT9vbGe/cEcGNngBDTt6yDf5uv8p
OCp9vvFicdWXD8qk9LB2h5R5eNA+aTj+n+p1Cb3MaJdFfJw0Y5KkCJCPF10MQcBVyD4OklMk61CH
WCfd7xYhTZBCK1b5NnT7yo+W3BGx27khlUc+r1fYW+AVPrCFLqX7icYsfRy/+4+mEeANbhqMm9g3
/ZWrjLsvXkhdpvEpZwJR0Ob7dPnsYODeP7b8Hx7GmtcipH04MbF0aGnNXCv8rfzcBXVbkwSEgkWp
N8/2nwxx0yxOcajHq+k9IQyF/xutHIXMwldeL9spqBAqAZcU98clJvW9y3guHgEVE0VVkaqFk6r+
KMK9ZYhwC6waATUWzdQ5L4fPFDvAAO4Pc5Lfk8uZfrQr0HS+XtK+E3A7VBsgqpNAhH5dFzNMyOOe
W65NHdEghV7UwFlU1UcAvgJlF4LwLELMwMPwQoBIntOB6YS9+SJ48C8j81tE8y8fBlpQ9yuCk/6x
MS02dcrmJa+Gpb8qZoOPb9gyaOGyP0acKlo2y20/cEKCg//bo9awzn+7CzZkWOBwJMDVMXnh7DLa
xtNtxHgkUyxp8S6QeYOYlvv0/uFdGn2kUk1Q+ghMTnwjqOlz7vfPEUsAFUrMV4YUSQnEFGNM6eUG
ISpO1fK56c+zPss/BVhr9wKJyu+6619uLdMW/m0iLMWpaAjk7LkJRbMBtz2dBtTbvUFSmNpVUiWj
kU02w/7oPHCuhdltc2djlBoWXogrgk+i12RmQpfn2ugaZI2tv2apvXmrwkPON7MJH4llwjrmZT65
GM9f98UR6Ms18uf7c/8zLQAYexiyHGFgLi38jkqIDL4O6LLF4DxJNtNtxHCrSC7+gbP9T5B8CHOV
Hh8qqWWZOtokuX0n9veOlh4R3CrZBh7LJeyJA4pZLedyTv3mLoH+nwzjJHvec/xo9krM5XI9t2VG
vlok804g2L0NdbSj36LY2t+1QE/cLax98OlH2tj7loRiZV3X+l5Fz9tLT2nYAgzMGCxa3J6fLG6Y
xXfb7vbdtwuZJHJ/ctc4qECs5I2OwhIDMQcuLwLU36ZMMxcYexb1ek/H7SfWBmvkoTtNSWlzApMu
rNdlBXtjO1GnRdUTJL01U2SKH5MMbfhL+01XXVkglGdhcmPJ2iVKPA63OtwzueEz+lM9WM1AKG7n
bGppY4QM3Z7IJKfjtBwtyZrOH287oiraMSB/yMKHS8hhYSsjdXhWtsG3OJ7dpChgVbKhfhGt1gO+
BIT3C/exex39IXUPFe+86B22xBGXO+K3swqEOzRoMBoe4MxSv1Yq+7rNG4Noazl57+wWymmUrJJF
n3jLCvyfEEfFjbTRvKsl9MeG/Cp2GwecBtIUHtrEhhXXeYkXbsCTpPhrGaZdYVvPLyIO2Iwci1Ha
nU4skh3MYy+2awzj8zNACsf9EfnLY7H0gPMVbpBF4qOH/J6UyAZhtlHZuk4NdKf9/l5jB/IE+TsQ
TQdqCnq8rpbHjjlCasgNZkA1wI29vqFXCmR2tHD9i6Gf3cJcSELFNYltli1OjbevvYo+VNeZYUXC
OCuMfFGSTFnqkTweAAtD/iW4XbJ1pCEcBf9AwEPm9XI4M4N3iGdCsrKjILTREmOd7u9hpiMt2Jy3
3ZDSaZNtmZndrNTY/UqSGfv+3U7l+lhZN/2u7GKBSxn9qg69Q/QwIbZkNR/nVpCo8P+mzwzath7h
1BawL5Fx1JAuokQnmwJ8OrdXx64VZ8EZiOOIuLJZ35O09oxOCK5EdzQVVIU3LKvuNMG4cUASIda6
xnJnUp9L1zExlm/OTw/0T0iwBsYF1/QCXHt2KHu1dqlR2TrdSbgmb7Udt7N8FQX5lwukrqMWuvQB
C6QclkTZxEjTIA2tHgsMrSGdWDvn48e+SdZvF3Lcissx93Mw8VFQf0RVuC/67HhFVrPlmuizJ78L
KKaWB8Yj4lH6iBods8qAMmeo1h7bINuREA/EoM2aTZYQEx8OFmSKYmxAQ8mHTRWWhRusTy7eaf9O
fzSW5Acf4e3TNGDYkbLhx/jkmW5uSWZx2FFanx8QaAJW4m49JjqzJFpKeeXnwSFUtR4j6pqVGtOc
bls2fw/1L03yUGQSFcN0HcwVYbwOisEIsL6UB9aX8rhXm3KKHHxQ6F8pOk1zlCgf3ctTvpiCUL8a
DX/9cjXPdaWlwq3sHI5OjJQfRjZ2btCDELg94sQF1V/SQFZm+Ncwc88hWcGxQzJrC50dvxdbJamu
QCYi/+kcKQG96vAVPjQLfPz1ER7a7OfA1BUD+f+USNGlNCA2u86WGFCcfvg42C7FTmUVly6Kvh8F
3BHBG7FUbMbJ7KZAreeU4pIpXGI6cDJ38EPsjVSbQFSwuOOsykoWivzPvxN5XcAjXJP0jChUiuJ0
ahGUsIyBJYIaek4Vd5HAE4B4iGgAEnvd7dxsyDrWlcerznZa2//FvlXVzr1fNejeQZxUm4xL8xOu
aH0Xfqwj7xHtwKQWurohx9dE1RbFTJAXfbABVuRH2o8jXpDe5RdHl2fdB25s8kvPYduqhc1lyzzs
yXQPd4Da1g/voEXKlir6T/XdboYd8x01u6YQK6e5mtdx0SNKt+xpxxEx/dhxPUfbbEukLD6N1oKX
knCedToj6IDSlXOGUwVL7jhvyGng1ftye68maZ1FT5UwHH0zUImMQJ9abWrf4Tig0UB2gOZUP1yM
YmJeeJufmKGeUHX6ad/jzljYblhhLnQWIZe+tQKhzw1A00k5YPWKQllwuuA1JUA1KpnmvkPp/fzY
qbjWlPPUOohsEWGV1JOaYniSzKVyIV6bt/0lqNzBXjg8O4nZaVUXp7KaKXQUQOhfN7SuEUhSwQ+s
YnYbNpFHW3iQkmtYqOfdNXKHhnPvv06L0gXixNW6+q9ABPSCva2iP3rPZ/+NEnYfoXOQD9Vuql6z
cTTuXbZ/IwY+QN2gu/e5ZexRgYf6Hkx9hmYdKyh1Gw2krbgL+s8Wmn4/Tb0peVshGHT0H3oqlt+E
QhcEqBCRvJlz0V/mlG1bkuENk3SHxbtBI2Kot/wH116hnBuS2cpE4drKibFzmT2ktfBlrytjjtqp
bfSdzfDkivQ+h9D/2dP+Ji+W3Cc/f5KLCXyf1NNaZMeLqcwkMEtiNkF3YeP+m4VAEoIuIf/ZEgwX
5BJOkiQvqYlF9cPvoT9uK6A7vvngOmX63A07LY91uSZisrRiopPVGVB3cKN7MX4wgmWS/tKWbWXe
XqbQCRv95ZFBSlHvDUYrxp0+f4IUqpPY6FGBHO7xJTgjre4Pmxi2PH6dblN7C37BWIcMu/3rGiAg
gwbVniZe61NxkROrM1TUMY/zMBFrXjUROMfnJu71LFkDtxTRWrX36NIyL3IYos2OArJXXNqtvWyk
O2kduckTKd8wnZbBB/1y3/YuJz6TmOvB2ohG5cu4P9bAUQrbOHWtvLDZcKX7NcsxIiwXKtfHIXBA
sJ8P3LHOajQF7uGj3WDn31AHIUDDuOO40OQC2UIKlBts0+aupUoYbJ90fMUHB6WUqm/y68ZUZfsg
NjJGFK70unnDw0JZDfBtVJzbG0FrWbCWH1aRwr/cRceUzFqMCgaXyeSKMWEGVovXYTy6fl8cW+z4
ZuY3n0IyTztZT8wo+lKyUWtbfRj/eXn6NnC0Ud4DSphPs4jpUj2Nyj21SrcGrtRLPJCAoqdU7F/K
N324G/aqOF2TVjMj1oEk1WtCfBjfdtBju2TfmBNHNNwTKmPVTXxl5YOEOYHs4mI6DRRUX6pjq5hF
V9hsUiwchig69NEKtoiOdhd9EPIaUzzGl1u2jAdXXn7VkGt8ChQ2KHMZpr0x6rpdPDwBzz4Bg839
SoA8VUZhtGJChWT4FeNy+weMOthKkBloGvOX+ZCqtum1JEFy85IZUtO6DcNnLH5VTMYAWjVwGjdf
pTu1W2VlaomuuuHRVC/+SwnjnfNzzuIj57YydWTqWBSRsPqdNkXEg3+lOZ1C/3n5mL9PwZcwYNUz
HaZaBSgvMawRP2EMTLNsJXLR8tfxO/N864WtSgeOWNWmP7j3pLzF9OQgXzOhpbP2/i1h3Qj1rE5K
eT5pqWbzd1na+t69UT6U34Tm9Pb+0a0Bo+tq1y1YsCNbyuCUIvV8ZnxkUGnMfldiVwiYBoHIthdZ
EW+RKHBUh9zme1gDfzarwnuD5sXINAcuOAI0W6kyTTAps4k4/O31dBVjzn1rHRUaa5R5s41oLjhU
q0rq28UIUshEq8yvejyBUMPYrxy3YzPk4XTbHzCWgms1OLRqROFu6vQ3pc8uWa24xRSgJ3g/HZTL
WqJnEFNHARgu236V/CQshR29Q05/NfmAZaTlYemRxKZzu3eyP6IxymHCbCw6uVfWCjACRSC/RGcR
TaPWwu42ntjO+Er0rNuMUudDcQM5tBylUpezg6mmQF7PRwaBbG6TDLt7+0G8EVMOmf8OB5eXlqD+
NWYEsl9MR5ROrjd+P4j2hlfICG7miZWJptHhVmZ8Q13MF2YpCbIBqHZ45PUDJyypJTayJt4nuhqt
voI5RfKgclagU8lQcmpozSmmTg3z6L3FklBruqTZAPRf4L56IN9rqQPfO8LVT/tIZ40YsCFDuR2J
iBxAYMgG/SEaNpA2WSflAWz9sen4pj9hMS4S1Y7YZehr5EUdr5jeYLQdr6rmb5jIpRP9JxAmX09j
AhbV9CIudwIaDb3lRFaJtU6eRbz47JwI54tL5RCH8BUtLipMrFlTK/QDVZ6x2sIcDaJXHdjTGED5
3UCDsBi5lY8NZvair5sOQP2pn3W6RiwZT+cZxtbciMr6nxvT/SzIBYTDat1KDQdCKX6A20OUBRWD
7v4HLjseGHfETVgbSdZSX19rIFtPRYl4GBybFUIv9KJ2r1ucz11mgYN68WMlils8hsa1K6XwH8A8
fSpVNGwbloa8qbzuaynt6RkkdsqiPHJTOpmqWGqiS3W/nxKTroLAc54T5T5RFHebwFC5KwtXtgCM
gtFdnVSZQhj8VdtgJJFjUddmw1BD0+zumR9daYhD8gzu/D7UrADnGfSchVA3BIAxs1KuKvFFy2k7
kasXafCQoSx3KvPqcs1M3Wyo17y8fbkkVo7sYf22aLtKli1TyyoBrXOuF9kFtCgksK82QpF81v0P
9Y1lLIKIoSDsHf5RzXOm2OxsFW7h2KLXXCkptwXkxy2+t5AeUi8lNz2drWgqkOTya6SdPDNgBMTM
zf3u45iBrqRvDaqIn62sVlrQmqG7P+wKZrlT24aQ2Xj1BomrKxwsJsY326PC0VTdu2T6Qdz0FYX4
XTdVg19/+AjOtTHDSIbXQv2jP3J4TSBg6n8gyDhu5KcejC4XBwg6vQuzlTlhN0YYNHBw//4ZXf/+
DYDNXno2wm3khJqBY5lWwvRy5NlMCj2D5+s8jrlKdictkL7FsJDCzYApmJYtbMZ5OjKcPmgnPQm3
K/EknzGRjFjOJInKaNssptDA3UmkndJykk4j60RS2a/jIlw9u7r5+wGSz9Jvu1Mypt7SWixJkBf0
8DrVUs5fbCCP3ZQeb6lJ6P7XN+p/ceOw12uscB3xeHofXA3BsCUT7D5X4PAFcqRCdDHnOe8wXwWN
D7HVorwTIhESWJ4NcP9+SfncqHq9F9y0XVhri58IM/9UEv9+4+9t+7BanttMtNqj9qsrbumWKbSd
scQrvXGSG5z5G7+cvyzC4dam8L8pOcQpF2RI6f/X3zvBV59Opclc5/0iIryZTV6TDngC65hOR7vo
bgg3UWv4x7etb8hyYSq9UUrud6AV+TNwwWo5gio9utSYx1ygxVC2b7RTFd13Ntfr9SAJ3Gk94oUQ
VAflvG1Zo1EAhOQVtSN1o+PP/dfTVUI7rcUHT3xchA+XFVJdEEUu7xHOKYazzadsfPtB9+CxNKBF
dFsp8v0F5UoHF+rDv2wMR8O4h7ExPRTTTwTgXYiGLPam5xXXBeCFoUkSHVEnlcEzcH1c1rag0aFq
rd5Ampgewom62t+TY+m4BT8UAKhbswjyydlMfA3EmR9x2Z1nt5IhLp8LGs4s7Hpl6+YmHm/YY22m
blwvIa8ydlsmvsKAvo7Bj8xK/H/OsxHQNmZa5LWSlVkofzktFngw1N6srBu6nWkdyXEv+VxS+mdz
Spz0jfjHwu2lrvxrVNJd4XWTEAzSfn6464DXf2VtIsGeknQhfHJZ34dan/Y4AVGFyBAvBlT8OqoC
1ParZuqy83UFHmoij7nsdueZiuVpOS9VPtmz6b5kNIhYH7aN6qwC4jeD+w3b8YfFZLIcAF78yFtP
sHu478bYpbozLr3PqXEL2f8HY8AqInoubzWDCcMQ8K7qMp7E5oIltvjccYrmgTsXXHIydXwS3qWv
F2Yqp/WXL00ed/p3kMlCDIJIbZHFnIziHGcnHVELBwjpG1NKgGgLAFThtK3oIkywUA2UwoIb2gK7
7WKyaCR6bY4j4PnF1O3tHIRlC9qvabv3fpmartTSgMzw7fiNb5Auo+fa2nmTSwORkEvVxw5mqUfy
FTjnObHI3ilox/siDh6eWrvPwiyMFZefE+x91LmyxPaDwjhBaRo2xo9DHCUlJ+CO7p9l97AcBbFa
q4oloVUuKXAeP5RSsT7yfWCuOxYlwLyckeVOFtUm7qy5STMsxR0PahaGrJ8tWa5klc/LtofoYufY
IEL9gS8AhMz1jUOKhvcx5ztE6cPcifuOWAQbs0Q7FSlyJM5nddbu70G3OrA43PTtYPsamju1QKbC
e0J90eNCib75b6zbmytARkV8Q10x4fa4LgWWaGDJ85OMo6nihcRLh86leyiB/lWlS9j0UyyLG4FL
f7XtphNU/HPcL4mQAIF+W1Bw8YS/CWSeuvKkWfPnRTXa1KjCWy2RCJYGwV4J6ItPcCIKGSQV0ALw
ufMn2Agjonh4dZuF9KpeaENoGkthhAdjQvAlhdaAHq7mZIL9LhYCpqtdunH73MB7nYQNEuDmtlAC
+diKaEXMb2TlhQaNnaVyjVHWomYvg+Xhk7jDtOCm/v5fsuf0SqKNq2GYz+ES9zRhapQEzi/yTzVW
dHeUWuSXCUlJypqyhjLeGT0UjJ/e7MobXfndOZBrj0NR3wejFvQJVA+cQAccq0XmUAqxg18x3ryk
geCDOT6LdB7KPn9MWVY7ewFom/v7+b9YvtHr3NM3V+TMZOF3o1ksCXxss4T7zBIJPxL6LrSXjC/U
o0svAgPtFRj7lg+KF4KqgxP64L3J4CKw8i5k4TMDNNP6fvp2AdVP76QrVIhFx5mkApVJKdbT+EeV
KIYh6KHyvsavkT+dwGR6XmntUyuU9kE5AFoJ0W1vOmmNIzjKFq8QAWTBM4/KwqWzb5f8hADtmC3F
xIWN5BNZ4uhorrmg7FcJFgp76x2bgXCezNhTjv4aVcMADhoZmHQxeqTWboNY306hPM8dYTGdgyd2
X+Hx0kGGwtr7GXskMkZ6sxR9CLEE5OA9z92QSmHhwRq+1lyLCQnZZ3WJfp8DicNXbEhcIPH6jf5v
UjoafEv7Pc0HrAlNtYakvU/+mt+bmgnCY2Oh9EybNbMKqVnk02Y5nZXwv9qm6TwpGmLeZOcFM49n
PLiEcWm8PKTW9V7tB3rjB3EaayHvInkQbwQDOcm5C1FL6LNPzO7/gDgb7e8aSIo5PpGws9OSs/w9
YDhQPpHEI3N6pV0uX6zC1d/pKqWkhNLDT/9W2FYxrkZQh2zCCMVTOorVVjFDenmae4rdpnbHwodD
1rES8q7Ij/6+gYXzpvDJUZCQJqjhDn78BSSSIG4oU02PC5I+oKR8QPDcslbX/U9Y+WRk+30VW1AM
FSXb2p4HVB/OPQM/3v+Be3an3XreH70bUCE20yxOqNW6PNyRe93wDwYFtWtflsHNHpYn/XOXPmjv
+oNiWi2H2csO37aTQKIMOzbSPKk7iCwWBVp5Nvdy6nxU82zd4DLDdDX7bxNb0zPDdTuuACHBz6zk
w8iFlrCjN3Pg2vvOO4DctisWuyDGTZojsNdPVfUwH7p8BrSBlvNCaF2k+3LUYwo04vq19F2w2UAD
PhZs+weg13e2y+GuxUTrhg8sLKhYhMeOXBxYyJG4nRGdT6btTZXQMSSVUdOz8FsIWIxpT17/d73T
RfhBDA2qqnkhzJnZs3V7V+lOIzfap4wR8CoSXOTD6BvIC4iAFWpvUFxgmDuVgeizU3/L8JyrnELB
u/561JZSzGT0GAthd6W50ujj0D/yknvQBqj99tvNCmrCkVgmRLYfY64prUj9NM0xTnZDUwt7etL1
Th1Z9xiUOTMptElP0Td8jdKRgnpCT+shcWeIUuMlqd6XTGU1xDwWCsyNx8DDjK17GfYxGqSNA+Kj
fo4TenXnaWg0f9RHjbu3jV0N0nuAvMUlpXosMTdtSuSu+c5t6OYG30EFu1DHpNOJU9Ch1wsj9Yty
oMXicZZ01MBBkPPeIOPs4WlJyoZzRDdv+wyukTG3AX5YXnubjrw7TnkhDIxxB2AJvEbHIaJaCIp6
aTdkutEw8NgZ4HZsJYtn7/8NYuMECKay3wRXtBs03n/7ALLE5Vi2wMJ/RYL4zOg0wkMn6FT5QwCX
O4qmBZAVf9ZXEEr7u3aetBUOv/Y44n4Ut+Cw0AzBFZfENidQRiAFw+uD58T6iMDKlKfvHYkClf4u
gPBqauw822WiY9/E1hNs4xFbYeC2Wr4rCJA4aMUJXstAy/uBeUrfvEBaknJiduUchaRIzYliNyzf
2FpTvhF1ecXcan+NEE/2rvoGnDaAxw7yhJcBa2oiQovma3Ipnieihh1gpOPHRCyI0WGC6j2CK1JR
TpGI0fArlo4expt90EDjzUKpLgr6cWR3RcbdkEx+UcFLA5LtqrXjIxg+UEeplKeASWTxlIRn/mua
YkAzBSZ7Ww+Svjv5xyW9CYIS44NUUP4oJkOIux1P+qQoA+8bxStDWdeYpVfuKZ91AeUFpgmqaKdl
o2f9SDura3iDyPw4ND6x5UL9AnXD6waFludsWHbVG5JYXFyVBjKZ4OShXM1JxVpFDhjVcCjZTUas
9iPw7mmG568fTfsUvmVliO2BCDOuTO59hbzbgkV+fmFWm5Vgdft06hqn6v2eh/ibEsReG7m0o0u3
+bGdIob0ljGOqyCMp/AGA6iO1QCzA34N5NO7yeDL3BMNQlf56rBvJeo0Y4ccobvfWiRmdjiwM2+y
mEwgGECDSJQtZ59zUPJajFUDmzOE01FIwHbCs3OPsTKJPKLRm6aot5462fgL8s5iVuv4WtKiLTrG
Iqvs9W+KpeVkqt/JGB0BltCJ1otrDGCUBeYTk2DUwAjhXOGP4r3mSH9S335yz/YZkjWn9iGOM11Y
koMaEN+82BjLAM22rRZ0jmDwrVXGDlFcRWH3pdhSoaGF302wXeb99Mlle5eAFnbt3sQS3O/29EZa
M2xTJsgAZ4l8a14ijteM4A6qIVFAW8vkk8ncam/AyDS85KwvMkYee3PrkcpgSl8vm3x9JN9TE4Hg
ABr0mf0zn1i+hhI2V2dbiH6JynculTlB0h2D30aNKbnJA3wULufOSyXWnKOdQxI/qMQI23JNyzvM
rewhyK7EO8fqaju6IxUNos89kzdVkwOwVjbDBorISswT9YJ+E2HdP9BD0KlW+wrVlpj279cHXW+d
NqgEfcPHB+Q5iABG4sp5XcQ5vEcYY9i2Lq0fZ+3RLR2X8/TOO+peAufWmmOaxjXH/WKOHRDOLk1r
9RnAcV/WgFCd9C+hbwMQxRzi+vT+DlNpuEv5jLoImSpJhTDnoUerUdF8mdIOIQ8QQeGk6Gv3WySV
g2EP95k3yIBMz0DkIid6ipcUU4InFRriGDQv9Yw6snz4qeentiEhNLftLJ09JAtZ5nPIGAxVuBMV
a3k12aEyHTupQ6GMerMj/Z37TCirxOAYIfIvi8KYfF2cvK1zvZYDTNO1xKnaC2e4yPUis3NRagOW
ctsmJHEVmwsDcPIJEYr34kfMArXHUpcy8EA4CmJxrtwgz1czW1yg+iHGAJKBSzpItOyyhMZlYvdX
r69LEWutnRaj0hA1f4PPgjUCOuigz3ypDv/kdC7CB/xmB1iwp7fSZ/8YYCuB4UkyxvIUtPkq/KLm
9zLn5FsEEpzMiR6RyM59T4spv1FVkAEKlS/WFq/224rNwrmQR49up5hpa0cL+o8uxoMaNBw7xuHU
cVvbW1TUBsMX5VD4gtz66g7swKHhvS5Pe93DlxSLQ2T+0sqUbhonOeX9vLCrvqFVVDZuBBEPRdkx
2sgQYTWPgBW/px7J+5ApPTOLU18kCISl6Di3H7o7NzJzgoQyx3DL0xXW8LlCrA9FHT3qUveul4lD
wzdkui34DoPpz+xzjd44R6DjnwqXetoulgPRZQS2TUUtm/0faiJ24CcfN2Z27ozDz0Tc/soq4sE3
8Q76nsXDzVOAq/Iue82a4x4H6tNOkzE2+OugqANcJ1G1fM7HkJx2e35MyNUNJQcdmlVkY3dBTVhC
kUm1BxSntAiRx3KdQa95ZE7EqTS6W1dsBZA+9pQtCWblr90Kp+LGV7qi5mFCFd7i4sVctLn6h5xy
cxSTe/Df8E5OTJxhSVgy9AsFsQhauLdCSyME1NseAHl7MIyJQCAvuuMPWi4yskYYq2LF0VSymi3m
nz6PlwwLHNp76fIgkK3cBekb+FL41ftc38tYDk0iETjPtDDDhQLa7hp0nd98wGZ56yL/UrTbcYXF
FCwwelaOnCRqyDKGmnuisgY7io39Eqg8r4NtU0VcoAI/S4gCiCK04C2u4p08RRyF2RyubosfKVtl
hlaK8UV8NxGWJgAft0UgB9Rd8Jd7c6BowkwwQWZIkqq7+ti1XA5w8YLTDX7u2Oko8QltCskCQFlo
uwCoCkRqru0VHq1QO3JT5faZ92M0l72hHFkFwWsojb5IvropV1rb3iNOtCXY0oM0HtHSAYxvmUST
BL3nbPwOIi7Tob4T/pQ7fGz07aO09dBLuRPfSitzb1OciO5S1EtoSX7aYX7GRGSVcJ2XmOzEAfN6
jfEWFCqdWkcR20MqjFcE1KGDDJnFasVo0ZGvKjb9lrJGb6mUWJVte922Bl9LA7xSDBqQw/lmR0AC
ggQ9muZUWSwNIZuvmkuiR1fvZ2pClwszcIawTUijK3Ry5YnxVMxd/JORJdkCARA5RdygHsn2JPWG
KnZNoV4WXqjbv5YOWjsWCL0d5HhC0n1Ayl5BKQN6QjhsSfuzfq4fNdfgmVAB3An5GqJif3qwquSj
esrR/vPYl1NApMa7jqrCX31MRvWPvlJ5Fyun1jJMAlVLHa2tgPMv/cFpzCoF/oFCdCMH4S4ZbUbm
JHGmDL9vHgi9xX9GSf2jqxeoG+PNbFXN4fOIq0g7IaG2fxkW3vDNHDkHRHCw/BHJ7+Hjracwt3Lz
l1knjCOro+37zxuaeQ4ixh1QJRq2Ro5t9gXddiPFuGsyRt2eApZJeIkXwe+zXr6i3ArGfJwXrLvY
bJsbyUMl0qtjBy1LfuIGj3oV9XCTN2fY5g/jjH0zSlFcYrsOqNJpnlIaZ2svmq7JUFzr96qCEDMp
KWpG/lOj3btPO/LECTlMzdS3bxm6+fPz2ytQSW1F1/5X9ixiR84nySjTRzjPWh75607EF2BeioLQ
o5PIedNCLyfhhJ+4ptCYOwLr992QEhRFiH8J2TRvKiYtH1Dlq7DB8t2/uvfb42uqG26Q8FoeXlmO
di0DPTk3A7DP0ShwpzQeNabenlJt/9ZPXxCl015uBhJApWPEu7M7mItDuqJy4lrKCtJ6NOnqEHeY
kSanLs3zGOYT9efjmk4LFAdd28PTMMCKAYNsDifg1LcHq7B0WetG6DVrTUjmhPJGwiqyZxUOMoVa
kGOfUSS9VKBA442avwQ0zVaZg9g2A1fEmpx5tScw2qRNNO1VDbhgNC7lRe9whoWS194K0zNNwIlU
BAfHcf9hG9swifKQK+4KGKBmv+U0tR0dbCkHyWxJfqZvSQhKPU7Wmcrea2BJ7VVLVdMrdPO8bn8H
h5yPko7uyapYeXsG9pWIjk5xdJmlgUViaFjY7cRpMGL+pchirepKBr6WWNZqXD7q1smEn2ODAwp5
1xT4n0jc1yJUOkDxNi3VXmJZsFi4qhUtgN3aW3dENp/WqVgAaX4h4X9CmoBisbjgOs3kvLN4X1QZ
3YmbLIblS7EsurrCIIAKw4JU0sc/4JnqmsmYrCDbhYJNhVUufN7qt4Bg96EkdLDut45256AFDGwm
ubLK73X5sKbDibULWedJqqgGit4vnwLPN3aCQe/G5Os69UaHWCR6ScPptlHWGQ4hz7ZlONa/eRiy
DTD6HK37YyLe4pRP6Iu8NWnKm2N8TfEvtLRM3tKdE2QwF9ZCchvADLx1bzicM3UsXl97GqsyAAIJ
txd04BTyw0BnFLFfUps5uOLJvCdi2+shbCNqeSDf/PEaMvBiE+QcyQLLDrYzbakVWpuFaJo1j6br
I70PEPNIRbI2ZqDd1KJwLErvIF3POXw2NaOKasMxZZKWk3vqVVzSgsl5l4HdsAR9CgOoxcoMeyJt
0l5VVS7Q7ptOLRYgE8TIz6wczpmZYP0VVRwCLt5ScvnRRab4luy+v0kHTkEHAZIWd0ftfQa5x832
AjvVUEOKjBuHa/c9OhGVJS4/3FbQpUAJD+uEmayyCImj8Dxx9orVf4lvS73qAsNHiKQzyamPPe9b
zCA7Mlzk8/KIVi+oPro7ytL8PonCapPk7uLKhSUCIsVHOo6e1qubuwxtZrq+f7zmfoZFS9FEc/Zk
jecNKHeI91cK4b9aqq1n0w2WyFVjJk79aOW6ObKKsdq8U9ZGolYWSUh1V9YlBVx94R/usKkpyN0Q
9PBwJolSSRKTrcYH86JUAAa2nAlNK9ntDQXWU5AkmMGHGs2HC7rATXv4i4t1Yur5pyieqAziHfhj
3NMHuGyIQyHg/AaMDNVCwbhGqvCxcYyyEQ3bvqBg25wwVP7Tmt5ndKaiB5TTlbmCPWgVvWn89CKb
pCERpoMhGv0okK8KsqdvxF6GU0FbjOZoWfm+vfRZ1Ga8q5YevtdlJ11IMto2QeFg0LtyvY2hZVwp
gzVIKNPTFWrjyPiQL2hhqCQwTzRhfo7pvlM3y3rDqOpywa+eFUmEQG2Q7TDN649XJ0Ety1V0jOEm
MSUQvO4M8HkmPaYYSuorvYlsDuDKfpUhHlFFsDgXPBI85p/TS907yogH2rDiU4uAUDq+deoKpDmQ
xLmqUx7ChKYUdPxV1yEKMrhWj9Ioh72Wi5uY8UFmmGyHH6P9y8a7ZP5j8gBFxCr9UBEKrbAPkZ1i
eCM5AS2f0VaX8gjCcAWq+Y89Ltp+aXsu7kJcHr0msf9GlzbltSwir5Q+45qmTFhI3s2o41uDTW6T
nid9dJVNrSsSrQ263SJvQ418CsPCu8KPbXN8GvJKqBqzjh8E+70Rm2ZTHzsfsQP/Et6JtfK/ucAK
Cb/p6dnVwBFQf7uTbdVp5QRLjYOWmWinWlSHK+Vv+dWwF3wY666lm3HAgahH7F/Fgrfv75UFb5kA
Lj2aHeVxDs34cuufOUWy5cet9ZBkZHvH0rRlaCfTFSyjt6EVurPJxQH8Xj5GLK4oCZDKl5jj4lcU
A/KDejUKlNrYDDCbcn4XsnbPtTpS4N0bmcY2xGhV3KpIWwiwRqlh8ZQ6ZCqMyNKOl0MkcsocGmmX
natXHMgcWGqQ5LPdgu2B3U3cGif/8UkKaZ8PlJGi4iYk9cAWCoc4dGU4jwOyivEuRdAsh2Nli+0e
66i2f/YDAFdgVDWNFV2HiHUJfWk+1WoDlab8yteS8Ixmk07YM89UAj3S9P2wSDpirCmeHx98cpgi
2gUdfcYdMoaPZattZp66ZT4szUq0vkTOg8XvpBiYyVCyjTkM1sWyJOuuaPFep3xqdXhaKamhXal2
rOux5y9Bxl0PbuztEdBKVr2XMsQm6z1zQFBhhr/AfqE6Y3+ebplhGapxmD1fYGRN7nLy/qq3AfEw
eeVTIHHHnSNatw1BVWQdkhn7jdKMaNXjLiQzr7KZFzYqSmLqtQlElbX2ycn+ROOCdG9CNGanILjH
TefInxjrh5xGyBA+IXsQor/ZgkLE4VxGKy6fM76on6K6CECJFI+7XJU0SRm+OwaYxedcU2+O4vN0
v2xNU+PRoRAoQWlXyytv2FsRd72BSlE+OZT57Dum0GywLZnXX9PD71lqU+nvGSXBBV35Diw/b7f1
l63EMGNar4GuvKbnFsWk5WePH+8gKKmZmt1GMIKen7xXuVEP/A0XF41QEHcj3fe2odMHr0C82MCO
P0xYyBWN6mtZVJkfZe9DihasxNIsWP1xR9QSON2xQaelHFuutt6nR4HZl7Qoz1IpbIK9v4rRFWjX
2ua7XEXmVMzXaV/60cmYIMPDjwqYuGuensWoQNo3uIukqg8qUadHOIH7tq5iNMXvQAICho1avb1d
f/xxX9Db+2FEISrgW28bWfVm2IYe5PnieVGydWxenow0EayWcFubHT/J8yRM0uI8eoP+cIj2soWm
0eVWKC+jr+0qIVQBQze3+dKnWyur2EQsPUo5zpdsQ388UpL002EygM6KviP6VgtRWcKkwrLWhCxi
8A4tRxSIHSPofTrzrL7WfOZouQKciSzGza4nmPJWcZIn3PBqHMGRhvX3Chz1tDtv8iIQGigu9lXT
icbry1OPfVlrvK+3j6QUCa6TCFsEssNNLzIgY75zI5iSVz2s6dmkIpBjbAES0pb4urVVAS+TgB9n
5zFuwJU7E/xqhqs0FLUPEooylrTX1H8r8MtIn7PGWXkGjAJ/+s23YIxUjOMMfVjFmf8sCzmvxrGN
zkTyUy7ZgMy0ykUhaXuJ1EgJG/HW65RBDKXpG7htTR8+r9i6ADQNZLACH8yELIYIqsx5Ci5b/sWI
LGhuMfte1OTgipTMwS+unL7z627JlivHW+2gsWlCONbRTItEMNxNA1ddWn4PhY1xqlEZV6uujGNc
kVFyIm4fRR1w7M6/iCyvnnaBX2nUl62CrkyfoUkMLnhp6mKcKYXG9eJ98GyWPm6AE4rX2evLHqRs
vghk/6oY5haBlgUuVVAd70M83hQY4bEC1V4s3FtjhBXNSSsR61dRvDLxTJuPUec0N7WwTfnyCLIb
ECiqjPL92mFTibl5iGgKxt+MnY5R9u2fybZUxL8Ij6Eem4PTy9obY1tgx5oYbojE9TdwwtUTsLxa
6zEAGA5Se6IizCp8qY/cUqi83g6w6CUkqOUX+aK9tf6Yqm90NDOmy4f8wKNSnt5Ub+EHUyz4Jxom
f4n3mDjcNt6ugzok+/DLeQtgQLTNMNLVlR4F+4Pr8msJIM3HFKgVI3WkpMtO+r9VRmio8dEUNBZT
7S/UAssrTv2uFxTF9L+C4rDvf51j4gpi5CFCp4jPdXJHjr0vrslgl6IEuj1GD4uGkaqjZ2MQ9zqs
kYr2tX8z2yScvYiSlPOZaqIqbR6v5WYeWty4dYrrLT1ToI1+UYok09rNUALO++vZqgVsObXKLGDy
J6PJNOq2ROHFplw7FkaJYkwFqM2i3IkMACPjhph/1qyqS+2f1G79255x28mQk3UMymU8zmwXGKDH
YbW96G8Sz9pJ+0BXJ8QHS0/Wc2zzTP8DnV95+/B1EebMrMy4Mxre5XOQmie43k2Ss1naOzMvYHuV
GxEeaURqZBAVgrog23zprdinYdN8ByqiwbZIm+c=
`protect end_protected
