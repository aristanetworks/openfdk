--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
nm15tvqTqCvLMQkd1vYECeykzvkaHkEz+TQ9k2U11YBiLDovVGkTIqtmMhG4RhMHN8qfzxYXnE3G
0OjhUy8/BSpKzlzz+3hvsHVL95P4PSnit2lkfr+uumzwas5vUfAk+rNbLlL6QdMdQVsuvBEq5ARd
XFDmUih+Wkjy8EeiXQIN68eN9wyWPEeOMNZreKcxx9nU0FduvvVEC3R0lJVXQe6Bu4XiQv2mJTvn
CVMS5xzSx2XR6Ab+zZFaUuz5BK2aENWle5Fcflix/OkrdsOTm+CvfoDVXl86fVH3AniRXyj/KLm6
H6peHljKUWdhITmlE/NQOTB1M/xwG8i/2tmbSg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="b/EAuj7qEi49HCBQ1McDjwYVUhEeCXUGEcsv53gtbpo="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
G1W1jVIIfjcvrmNpke9MIOOqmPJNd48vIP/cZqkSdNpC9olaqYKeUvv7vaKx8L87lbXAg3wjC2OP
WwilRVCemseo1/5hlNUILWcjveLNqsPNlCzXbSmQ7FoBcri/5qdTxT2w2wItRcAOPfB8pmkbvp2P
/arDgyFLE/xkMo0VJN3i8n+fv2V3dhyhOjzpsjeVckfKTeCHBnIEwKAQLojW5HrW5BUDM7aClOEY
sddXNhU8JALyAVuvmEM3SYmxC5iNgdqP9ApSCt5QTq/N2T+ZtI+7HYNQeJGN6TaG2FSUOOSlZ4Wg
RKx+wW30/gAGKY+OzT73SYv+oK1dhxwKe6VE5g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="cVmMDWxnDVmMZAjEAVou730J1+GeTKtkEf5FmlGbUMg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2640)
`protect data_block
Xs9hVpY2kKnu8OJI78KNTA3u24MSw/76zmCSDKu4hZWdwoTzRVo4K58aAICxFpUmrMtTHfmiV/wk
VVsi/xV9n09tv+y4GrgPqud1klaX97g3mpMgMQ2HWhIbV9WrJEMU86OeOGbOm0BYQf2jGAG+GOVC
ypbXTiIWIWqjLOFXM/y5wuDjONcr9UrlZviXhE9bdNkLN38Gj7wTruaO0haFmWPkivierUU2/bUH
KRIwM2Kb39MlE5POB4Yzit1cLpBdk1YDoanCicvxHw9NK9TSb+ej3rdvysJp8ZbTxpUrI1awNyU1
enY/Ofg1TSbZM9jCq0lWJnVYuD+j+sX/aX797h0iinqvJjWWCDOME6CT7NRucHJS/lTK5d3vzLrQ
nz0VuIRPZTTYguLppPZTWTgPGWzpLfWRlLQm/xccVdH3XZCBgqkSiUaGdU5FgW3rl7d16PYOTw+l
Sd9QTiY7L9pElxQZ8E3ToDFn5efVb3BEdmBA0zzJUGCoUUz9egiTWOYeHJfDaIiuA5lxpxpKZPf+
YmJng6RABuBWjuy7nmJWTxo53vtZPUf/Anv2WbeO5EhGkOgNh2/RClzVaJqQO+/ULddCpK6a6O4V
3DrD0t+3FJJLVPLdekCdvGRFys3yzZoQl/PsdGRNX660bBCG+m5jMczIc1geI+L2WSpsMptP5uy8
C3WhXtFtd9KQ0dRyO+p5SmAg2REa/y1LFPFayfMfLEiynwxGJ3Bge5m5x7MCcOXE2b3PrWAF0SkR
Z2n3jWVaPdR9aMGytoISU/8CFwP0PB8LOdGxnoQigBps1WkDSqTgAD5AaL7tztLYjqvBjWatJLxU
4vHUHOwvCOQAbQ8nYeteFML5K+wBQ1tCvQEJdJhvqrj2UZo5Kh0nEpVIqApUMzaQkrWObpamxMO7
9z2+IZQzsGWwEb1SVxtKFGfecCQaIB+6JrrHniT36K9m31rzz6Yu6P/DqscURLt0mq1RxUhWoaMj
YeuW71qRsSRAI2/vnutbkjBcBHphgsZqwFiCciNXqA/X049SAzXXud+XPHstCRBDKWKiwQUWfBID
Vbb4brcaByaqqyOBtbGuwM2tt2hcIUWdESBU3kEdSTatIxn9FLFikxRSDGOGYow2b7zegc5xw7Sx
3QHO5dHymXyUHTbgcH9Wj6/6nTR/VC523kEREVdfPQT2MQP/tXM1IGC66bce2AFtP6CqG9ZBpbWz
LNSsA/Xj7yrvT3Wo0/TcPxM7BGEPrx+13WnnIoKYrGcC2QHSdELLrBn32IJQ0FJYSgNan1+8xrof
TngEDLYoJGN5IMKHJ8t17y2hvzGT2Elv4UvQKXDOK0yvLlMRyPBJQQk7fMVBI3co6T0pOGPAzoWU
hcOfh1C+My/Y5+l4avZP/llkVdUzxh3CNd/jEIe6VmKRDZSi/MnX1ZNwT6UjXHxB3eLxig+d1dHI
6j1Xiu43Hqxvv8lxuM85J9uWDsSh2fIjBFOo/MpyorP+mXXiabuFKxWzDhXF2oiVyeOY4LLpUxkf
vXOb7t7foG3MUXCcQHv+A3lOicocbiGhRBWby80/YCalTzP31AzcdWEPFR+Ri15SBR4/7/gYRviA
al8GyCuaXbr639iKEQgA2M9ROM4t/ERYRCfifRk5IA//NxJ2Iqc82LywbDe3Hx/VsT/FK9HjjAVu
cdJ7LdT0Jw90sGyT2qVlbyoq76ZCDr1DbwnUc6SZGSiZvjogOgCWKsM2lf0y+vj6uYxhJgYNzvZ3
3lYGUd780f0lnhpPoSUQlbEP2heKAttyLnlLI60SPbIUbdkfE4btNZD0fVZnkEt1+Cdrq5CESaBk
4EN6FiC8/9zSe6OON8EluCnQpYZubKU/L8KeHIJwW27scNM3ZWI0BqF9OnalqyHtofrGv/xukRUv
UPzUy7pqlxHd+X2oc8IGPfUv8FWJwOms5mdhCY0E49e5mQeTOV1RE/Kc4QwykaP/4cG7XVdoM2i3
MevJSZnjz5fDscy38hxuB9zUK3Jf5eTmNahCS2p8gdC7FyFx8oLlgobBy/s6/GDGScA5+44+DrBK
DcekYI3JMKdN/uDm7w1RbuUkpL9kaEHdqtGG7ChPP7buL7PhdyzdgbcmLQ1tvEHG0imzbSNTRgVF
/DuOJeQkYeW5CvkoITbWrtMZavbq5RUNjB98IQNV7xMquotdHqfkB/adaHAw3+Zqdi1I97PoJUNX
yyMW1F+H+BjSrXNV94p5sMZQIcbgsDh0n+oeyGq3PmLdJfHcTNYT0eM5QOr+NTZPyox6lxY1mNu5
mWLYugh6LXYc0dalOOFg4MJO/1qQDqU1RoAGxhCMuLn9Y0S5Sl+WxK5vu1IujFIgPozM/+1GgMlK
8Jb97cW9L0jM067g9CDym6iML4CH+I4TNcMwbWhO9F0eUNqRbhP3qcfwDFpt/wPviFlSXxKDdNdE
V2yRvYFPJSWf25idTqgiw2zbmarwjzPIaGplpyJUEagf1zPqjDwF/ynopGuDRjuFqkeg2+H0s31Q
zFVOvR1G3ZPBXXyVlrqTwuZzk08JZvxL9TGm02dKkYBt3wyL3PC+cHOUHsf5cRBVJfnDsRZ8yBac
B8r64qfzqxHxcqaSIZMfMjVXwC78tBXMIE2tpiNseVLcD7sGjvgR/ftej5qsFw/RnSqHHokp9tf2
GftaD3393kvmHUAeSSKnOnbesUgmK91ILnpLqCpI6Gyt2NC71/OPNAy3/LqWMe5havhLQqbZUZDv
VHYcJeVWcxl+7+jHR0KeXKcFauhm/urNYm2txumu66m+h22iIGupI6G0Fho0RwSjX42UWF73wGlS
2qnFmnLLstcFuOZ/TZvTmXgdqNAOB8BktPF3ZAHXJad9nEQhQgDXtnHUyFIkBQPcmj4Jx2razFPv
Vkfk19F7EiFlfA8swAVfv2IByMlc7JasdtasWiHVhq6ShSiqnHKNS+PKZVuWj+Xk/zJB+7AKGYPn
K/ydw3fjgf53mxJo1B5+FEdq+A/yqu/ZmdZIyVX7vTsFtu8xLgr+Q+oHXI/98ORugM/S0U/ANtj+
o6HYLwOongzhRsNyzyeMIFTwz8oAi2xqXnp3k/zAER89TtmCdlUeWD/XX6e30ePNbhqfc5zgXHcS
1/yfbvnGRTLDceVJW7DZ73jjYL59orbNDAa85blMxPRRdG5EyIvEl6PgwKsgIkF64jUsCExxadqL
KQP81R2TyvAyea92LDuW+dJB3rPyGxIQ2ONlYKmKZa13mUu3rWpIFNNmknm7zo/wdPDFWJuvAawJ
pFFBe5R+yjD5KOaudPUWfE9rjFINaCo1IfzmIVA4ZkGrf7/DwKIjbDd9PihgrwTQ7EoMUSRR4hp9
7g4YZkIdlhLJSlaXFQUa9fyR90gPXTDseTyy1jfwoA3otO33zOctPjlPLeIQA0VoKbsqAg2Gp+Eo
yy6QaAFZSPmwmVoMCUhwwTrwA3GuqfnSK4vROIWG5vx77+TchQUhvJfnLIMz8/qk8n60OYrhfCaQ
qDaPwjoDPqmo+AnQbQT86d3n
`protect end_protected
