--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
IOI40GQU+omOiIAlddn3lBbBrNbXZ8yhyPFY7xwuP7B4KfNx+JfqLRQf45kwaqmt6sT42/T7NWNU
Y26+Qr/YS+/c1+GxjWOXxs7pqfjdvNuKdwfh1+jnZWCsaQFYNAu5S5ACt2FzZjgbGHs2I1uRDFdP
IX0n2greBgA6TVzdEoAcUaz+w4YyJAjVE6lA9Ky/Uv6ZNLx1BNv8XxsqCcGPK1k3p3ccUSvebCDu
u5p+YEVxfPBFWqdHcwluNReLr5NuDutL1PUFHtD53/3DdO9QWlODyI4M1OHhslJ8rBxceOXJBaxJ
MEKzh0Cvx9h3I81WgmL4Oxz6+Toua9/8iVO17Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="23Q6nRUb7ETwi+xfoDRgD+scNHePNFOtSmMADR/WViM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
YXOOR+iSZsyUkDaBxY9nZ8aNGlcTZ28sfKXTiOhR5HA3p6JXQk5J+2CIv7YIU6djUzOZfxPI05Z3
q/LT2Y3RT2Vk9uBtFt8gaAZ6181Rtic6sW6pfr/nLQz7gs+TIddMeKi+5ukdsC40KZZG+5cuKM6P
PJnQyJCWY6PLxMVEEoYKp6lhUyxYXxwPRvpLQwm+QLRMVEDXm2uVi4PLnXjeE1JMPylDMN/tDJEq
Dw4dVebCvpx8EsRVyKOVnyG/YIY/5n/mFzSNzgcy//ifx3E50di/eUhlvATZreFmpBKpDxxb9y/i
2Yl80n+6gcq8+nZ8ZvopcDoj+qFz9KLk0O/CXQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Qge+n4tU9eBcW4ev8gGTVEVTDT52KQC1z2GJ51DLr2w="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6032)
`protect data_block
c1X2sK1Zy8wvdsWFmUPz8hBoevQnjkoZ6ZWfBfv2/XfMUnIMtE2L7h3adPNWIREx5sKvy06bn4qE
8cYSXk3XisjHAschsE6xBtxUvlHFimzigkp9S3EROGSPb5SqtTiqXuZrDpUeVGy7KCOwqhiNCntK
dPrwUAvOInPXroqg8vZyyqOV/D4SwnRu3y+R9vVhJGkwD1GVSQRNppqaEkb0XunbPkt3bJtm+69P
HxiDKM+0aoJqMWF0nPUIL9PkNOA5G8AAyl3ad2cHDB1vBON888eb57+9a/ptHyAAHQTkWgEBnvNl
tStKII1Qn9XeYFloDwln0sIJ/JKbHKH4M0Zkss4bdzu9rlPbeFiivh37B5g/1Jdz9UazkZvWicWA
5rfdJ2yn/Z3Cl6Iv0jEOjYc7E6hfs7Gz42ueZpzVJhBrhvj9Juk/5PFssIVjFcjRZf8idcIwHKUH
+SMNkzQY2ZL5ZPIw5ml8MlYDCgUke6iIEOtA8Ps0JAwm9J1qCJOF0ihpaojBjx/hE1NCNEx4Bl1/
hU2LOBKL6cW32p40Dh+xkuoj9CoQHx4ivptDO7aucNB2fOtHsQOlB4BlJWHKs35bSbn6PY0y16iQ
JUrIcOqvMXhlNCXa3f2i5CntHRDCSxpkvgzDQPrmYuaIhaymwkADgtr+qjjkTX/mTZmc1Dg8n64H
KFANsZbylUIv5Iz3/Th4Dqe8EP/Vl7QAn3sYkC1SopJKDUFHrSt18RZ5RN0d6A5eYDauQz7Wfj8j
HmeoDvJH1HVrhqH/sTgM+wZn6Pei9iNvYec4PFCMVagOIjJdzF9JJyuIld+8qodRgUlcpkzdThLR
7F4I2R1Y0XxFJx0YEiGRzZU8XqB5juHBycEF8VkP3On/H2bcO13S/K9mdGgLZE8KmXKjQj1bNRc/
76/GOA06T7UNQUgdGfR97sTFOmoeuu3QBkpeTYsIr1/cDssGWuTpcAlf5KjuVTsWRs6WGYHMEYor
Mi/Ym6Soyqky6CEzNuPxv+xa1n+iF0NXC+0YXzFxCL7Wier4jpLPAZTolKE5NDR0uTx/CZwfND7j
na7wB6AEOQQcvmqK+Y/kemu9Z/INkQE2QYkanzJTjpkE8AmVJv9CbTwjEyOjNKMINXmZ4qwT29oT
1ngD2MeNVgztr/mMDEqEljbU9hZW1Ik6Mah5BpvXQulcwpVCCmnp/jPqBisaZdu/l1o1H4oOsiYt
i6fV+3x+CnHBZTVWRU3KRhyusPJ0SS7u3zG7N7Ylvi0FFJ68yRZw0aIW0uPpaBquIywXO+lcew9W
SRT1SzxNzge2UjJGDh6Jqndblc4oOdUc+iNe3LV9K0zrDGPLOUVHFTZ5AM8d9ccnX3U3QbsHWOXX
T4u49CaWCQw6BzfB7zotM/Lvb9pSxaJ0fLXSerf0aeLswvVo85A/cx/osU+n9fDx7T8U1FypJ8r5
kOuZDtF3b4Ylmr/it2HKIk38SXnWUuv23lyB7Ik2LkjWCQo55n5vlC7wFOWnyqH1xRVr/Y/4jEnY
R7Xi2o4mqKLNK8ZtTMBeKqPp6WifAlk/jFlTxsdaOf6/JNE9yTgjMG2XTFre4271H+Oj6V/sCouj
ENR6fbsxPkFITZ+1V5HoH0FmxCcH1s7w9KrHpYEZFiQnldmUbFyhpcq+sy3IDfc76zNanfXsYsOV
g1VFS8eXZcgcIg4YIbCe+k/uKaEplA60FxX3/RWgRplZzAiNVX1zQXBqrHlFtnDyOhJTfqqEdVce
0B8SBQo731tnz0t4FTLk93NQVwfujmyFKnNKxxtzYeuhKAb7QEcIO1UP9VQc6mWxA6bk4Z7DHd2w
4VrLN7p86ECpIzZIfeaa6N33WV1GsAaYhcokDv7DQNZNNHPgYA4UR2/eJcuc8OFdtrEG/kQdqJyC
XXnqaY2z77q94o6+alhPYW/tdruLqZIP8sETZOZDINVmB7bOCu5Gg7WFyx314k5OJ+5ARITB8bAk
RdtwEsDiKypdyvFA5Re+or+4p45xC5q7WZVdBwC6H2SvGwSkcXuCFErmK1aRIm9yzHJ2PGUF+3I2
Yi1S/ijjpNzpBrm+FRgoOC2h02IC0jDbs20esughFusdyzVjZ0W0J6o5+enwmIssY8Jp/dG2hF6W
zCTtuQ0p+GsCOVQ5j8xocBOI3J0IwWPyqkEO3PH9vPGJoUbsDXeJlMejQJrsniZHFK1ffVHz5Ec8
fh2U3fdyHmct3YZWD3/t8US8oH6Fyc/Zn70vXQ1gUtAGEjbsbMXIvItmLMnzuwJyAflDv8eFARkn
4YNdY5t+Gmm/lPFFH/4Bx8kvfbFmdGs+Ug3qlOs3bpY0R9oSF5zKmJqTOHk+9Qi9s6wkrg8jgfIB
kjNR1ZXxxXGTzm5bkdkbeeoyTPRO0ikG+zwBTgG+X3fFE4aiwlVNF1DNdyR8QZ7ygz4CMiH93EWp
486ctfjLX6fj+GKF6cu07mX88FaaNK651zAN8xBz6hc/w1N2C9kybqQ4kweCzO/1jwpLThdF+vjB
MURbZlB0ihi5ISZAgYksViWfHEHEc8yg1yl0SeP0q8UPl9yZxZZfrDVbxMAJMF0bHRcwBcbzLrxy
LSU+K7/NTzDdJtXUi4O1lDXtPesiYMNn8wKdrDVhdjBz5n4m+eAO9sLQ79EPypHSpKlGp1G5h6eU
ow5YpaWy+IzNecSKkkIiKrGjuTteaXHfPuQuTul8NjgO1S//L9LbJagxQhbeGpDnaAlQKC3No64g
OFeK+Qcg1orwToeZYs59RMqi+xHWoMk5WIg8aSguRJPlpwFYltnZw1KC0pldC5DD2iw4nObmz5fS
+Ovm/Q/WQs3QiG/pPFgBS9wu50ZbWn3kGPk7AMRVGa8crc0L0vPCGCg2i8ybmwKtmlv1in2ophx3
qpGYx0DePWPLUcjKSx3Czl4oHopxTo0f9Shh04jKknQX5s5oeBu2BUOdkmAKoYA5+xyT+lJA0BkL
riSyziYpg1Oq/zLZz/4v1nphK4ZIu2RLl8LxfAcdeWDuMl1E3hVD2HR4yT6d017JxC1xyiYX9YQw
oGlEKVBCFn6BJ4g2r/KT61GEquuXNgSe1CWapHc5nix29w3D+Z96yQkTA+GdvGbSM2CRxf0WqbnK
qXDyoAWYifD0kMtkG7KKVLzJYG/6JRGV9KqVGZN+uXuzzZ90b5xcBzmU5uOEmyqsWj7p5dRgldsa
1AnIRrUFtIZCsJEQnl5oEjo03sQjGAZa17u78x9pdD089ylRVAWQPzGy4cCb8T5KbFkt3W67K74d
lVEpY4d533jMGLe9gusr7iUlvURnr5jlWYJkm0rFXQZ0KN/C76hFT74c42VAEyGnsMCAXK5S89c5
hcTOgcumKT7I9qrczh23tHANYN3phiccyY04Jxg2NNNVU10pyYJqISSpmxNIIAUcggLe0soMAf8j
VnJtrv3IPS87VK13deHm3ln0PPqwJW0fRVt/C6z0Yc2fhlQM4UA+PCZ/0W99y3e2JVHQ2oZhklaH
M8oqjtR0+9sL/h7Ga0zAUx7YgPfxYI8EoUrLs9wTQzpQ4lyVSHrtAviqcKpC2F1CZBhjn/59fPoK
Znk5vjYc01P8s62u2x2L5Ncpk1Al6BipokpxaPp2WIkbcs2exZpPnU2kzRmyuoKSozBYd8wS8jiq
64U3eEGmcVA8f7mdvLCvlERABtcGsrBSOfuC1WJNjfUCp/bk3MQvlD0HGG/Q1rTI/F43kqZIkbM8
nJaquXaAZ9fKMWp9/G5yMRRC4v7va7ZqaILwBVeM9g8gUTVq5CQUq1uB0wOl/MSZtLB0VHWk5tUv
CX8owhi0RFTbXUBJZlUDyMiZhW1+8g2jfxEI46Lo8kxBWZeVJBdyTN7Kzx8Wg5/cLXMNGyrolO7O
ja+/eU3Np2SlGEuMqg5Q8AW6Yd/T8HOIAkasOSa0wBvSItRoe98dlJjNj6on8Cj1TuAeoU57Zn0/
SprmVdbusgZmSoQwQ7PujnmyM2e25hv0gs1fKQu10XFVyujO1HLpFthtfl1UvxgtpPVVggbjmL/U
tsBHTlyHlZOtTrjgO1bWYCn7G8kQGIdRklGyD1KIuJtH0WOjNZW5fsWXsx94ofn1nAYSLh6at2Eq
WhZ8b+hnFfJ0R+T7+OCwmPMCfQglk682Rz/I5Nqg1WF06o/F32JUWblOSWxAi6yIQwm7BOqpWrPM
xQzwWXt+dHw1ugce82a+JjL8TnurYwYU+U3iRnNQ1qaYlUvneOtE44Yp6LWF+nhZPefJ/bI2waBC
O4zcSiIA2UmrRJzCPXdsMFHiiNhGUDLspckIwV4fFcPnfcPtKSUn7PUm0kKYTqhYI3HQwk4N2r7A
6Sb3cZOBIHcVq70gdSekKK4ynOXDqPH91EDHBfnAiYlmJXq4SxH1wVdUhqDTg3r/AOqOtbzN62of
xI/2wxSsye74H93dmFgtJTa6I8pIy8Xcq1EwoHqgIAuRhSPtyJlgtqSxNjlE9a8Ru0vXYclQpVBm
N4jiBP0Zj41lO6jFKPqBRyvXRNTytkuIDE5OdRA6VQ6EaDiTwDuLdlJ43gDvK2FDqn8xSoOXI8j2
rJqF5stqvxDx8DzYAbymywJqVOAqHoS8JjUiTYuu8rmD8QLWK/b79N3n97kYe8eQ14UDNj9gv8PT
Pr97XjKEL+Mh2iSbP43b0tyRDHl/UsaOiiUvZ4WtGpZktAvmcXfSQQ5+EJwX1ipaNn2kAEmNyJ/m
Y4ePfgXruP7lfQMyKm2FnC6m1YWHL6JMfKlVH5HFLh/N1CCZfZUfQy1L6ETT+1lxoeisSOVPJ0ZK
SiwG0duw01zC5q/zw/NJ9kzfocpElqb7FzLGIIFs3sfGkyRc6NHKXGN8xJsEfvcwf3oydRMvWEje
2GRLs33SYlj3iJViGL/yS56xBZnW4sY8nxxzPiGDdmSLjORSrp2iBZyYPukzQ9LKeVl8uREPVU65
AtYo41yfz6+z6+YKNPu6AnnLx1zDJ9JBzkWSpolSJgghbkrMzLKEvXRp71fgdnFGCxuLsUOGFOzq
5jfTxCGv8n2KhLXHyz+HlHvFNVwsvxxAgKD41BpVcS9X7mLi/sUjkiDDoStb+tV25jIE1L28oV1V
WIfGTBU+H8rNu1YzmaUk8yQit9CuPvd/F16K5LCp/NfJw2+7SgSrcv5QNOARNX0qBbe/Dp/LCq1K
hECKFx+1UPKc0DDZK9yE31mE4EKYww/KWPumx0vipLoAieF3BLyxBq7TZLsetd5uAlq0I5LPEhIz
px2brSG8D/zhf/9wl6EefN0WImv2sQ4XANVrZ8i1Nxix3RT2fKGdDsi1rNAN9s4eYFlZLDLyTW/p
PiIdWxx5LdAJ37w029tNNi6rSlQt5IphdQOExonA8te5VLnEpm72TsLyZjvHKs5KfduxGkjT924z
mZGMKrw2+y1OMsabaluHMP1hVe9KDLi4Ygdw4YHokKzhgnXeAlkLoyFay/R6zZPygpwP7Cwl6H1N
7itg1mmC63LV+VA8MuV0DB+333wXnxdj40tcsLzK5s6Fhp+qt50GqkDU1gtzAL3cBrW8VLPz01wY
neQjUObFXkOMcwTH+EfgfjK42yATevYF/iYLyW0DlN5ghHMe+QAHsdooMbslt8Y9XG/pqGSp/hhY
s4Bbl3AfzZwWp41HhHvrUaq5G+8K+H3rtGiNkg3iZ5/uMDAW9TeE/NKuPOAjYFIr/5zLbqf1Nljx
+Xe4mlI2Aa5mEetani+APDRnk5gv0aGka2hExutByiWWiF4uO6yZxzmxxdoqOCo9sMcPj5pxRWEX
/cFBQvYobXDSuceau1Wf0zg165m0NykuXLccl/HERftxOw0OG7B/+aMv6UdQBCvZCLeAIrufvUfG
XGyLEpRQlGF+laieKCI8tynwCL+RHlfoGxVU7UgsBNpsn3zolm5jJ79xdb0S6Jr+CVfszRWOhX0D
lawsEWnw4/Zaz09u7hd2baNfIAMpvL0uh5adTLAGjhyEvzc7z10G8qYGZjd8Io9E0JzJFK/v2sxs
IhdYcf/dgfzOcn3f2guTKNssu2Qp/DNOleJ3ATa3fAUXlbr/K7xlsKLntDVvXyKtKNE8JlZElAPi
o1QzisCEeFVcgM0zvhnNK20HVyIIPpbJ9JfgwkFYb5MlZi/8KAp+Gc7c70nb4dvmt0qNGQ4ORjVT
xuVIL7ck4Gmqbf+xwnxn2XGKOeDQkiNcPX1cLoV+7Y/3Q8GiSgtx1za10rd7DCY7HNxxss51TK6m
IB952RNwg1G4wXOqv/h3WCEgZX+yF1j3feTtlnN66javST84z6QDDtGcrhi8xIqH+onMBvAYKMOD
ViW+C6Szk5gwvIzPTJHQcL+5o1XMrwrwoijh8Vb1EXb8EWZ8EbtAhJF6H3+A+IS8vE1uuEvEg/Bh
e1FGs1F6poE6DVUK4Yg/deXc+n3aZ7q8fmjeRk3VeUuc3OsdEH2Ko53YI9x9hnNWkMpDqI+GDhD9
JtDFdT+yJHlVNvgmvkc62YKR7dRInErCy6Z5lulUN8gjr++lSkeWC9hjcX1FCWHfo2asj9H398Td
PLV10wOvG4vov4EsVqA1OpbMtyZrdhYBgNtmhaz6rCKBu9YNboMJwhcerrib9IPuWh60IkufK1y2
lY520otYlMAGr/U+fZWEUXe3K6lFC2LD/sjAydp4oNwLDdf8Zd2Y2CSUj2Nj6UgQZh4fQ/XFt8zl
n4j92CWj2CnYBXNJWo+xi1aT7LwB2SuwcfxC+Fyo6QQW9LK0clJejBY9X6W3dHYPaZXOj3EUTujb
fIgOhT/aO4IIATL2oJhpBzSdjsD8o4JvJvpW1o1DotjAt86ZEAOdT0lQISoUvttzq1O1kJPGyo1A
g6QckWXUU3XPssGCwBrzbdLuMI8oEQpNqYBJBBPDeTD+nT7BdlnF2xtPbvB+dUgAmAXku+93ZQGu
3M3uJH74KR+feZaHU1tq9+qQIY0g3YfcD+ZaXB6l+F37/zQ6oEtHRFmdhlqJxLbxx8O1a+mM1/UH
SgQy/mxFi4imYkxTH1Ri4Vo7BGk/DtSKTHKnJtMZ5kkDBS6MFpoQuJd4ahfYB/guf6qVCyfgW4R3
tSev+DJGytYGoQZTHzkm5XXCl2398NHrk8idmb9mtVvqbZUsXeWLir25p+SnWAOCgypgQNpK8CuY
BAinZCAIoJQuTJlpQgGoCF2Q2xCdNu4QAArWMRws6ZYeV2a47DiJiwoEjbQEnuWCF0HO89cR7DIj
rG1px5MPO9kmWsz3B1a1JERd/7n6jxjR1UekiLYlq3z9st1KM5ZMdogxFoyzCTfl/6+fEANkwYCs
n9EC1MwhXP68OhFVZAV6+9lQp345UXYxvaevYo3kyno5YLTq6x+g1Igtl1Voj5pp8MNGqda+dsaU
I/xPmgcTL17wBwHMIvXdnl+ldqdI7U9w+oXDp0vzdPr3DjnRkTx0g1+SBG1i5kKDexgazrzaBCzu
PbeS3B/S/wsIocJYh0UgdOCCf+xGGu55s+MMcPRtI2zeSJgVZ8clehbqSHlLOwl7SKWxbupCKK5U
HKCsrb4rFvjtDvOxFXB2l/KkSZVXJjgmf0EhE3PVpH8ZEPEFpCPrYaHySAwRF/IlwZ0oCD6SgHe8
UEhn1oYzt7wBx4pbtcj8ITVtBWhrVKOtHL8ewMYyKTi64GYyoTgv6hmZQbMfXUH8n92I+h54Xgqj
nFGMWgQuH51S5QF3ORFMj+C6CCFe04D4VnzEOeOuaPTGRoUXwRDKQQP4OgA3c3bm5Z3tuzXnj5Tr
4iXiFYtA8VPvzNL14hfTKeFv/+pYTIxTZzJYkJ6zJH2HFOqYlRy9zV2HI11zjwbvFTkUZJ1JZtUD
vBD/DL2qX7sLGD3Yh2iqO/NAaZNFV0jcJ8y+4dgg89K+BhywvUZ/w21P7iplGtOH+i3kxTpKxIEk
C9n+fVEvg1+WWfVuy5//ahRVPtKWm+QPJZLG/pZZRruuchdr8i+J2NKqCqNGUaF3gKZq0LGo4Sqy
QREHOVEEsZNnDdn8tMVDwTvAsPAHUWD7Q12XIctp3znmIVQ0ea9Fii1Hsk46xFY=
`protect end_protected
