--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
KeFfADLEn9YddVhdi+GaByCvNV1YpYe6/Jm/rBgbHtMVNkP7dUc8v6sAMs26N2ymXx+37bOtTcBn
MlSsUfkuc0t7ReJ3NuLVoqa8qokOno73bcQmXU6r74rct/wHAvt+omIShReXwoh4B2pSkr+a1oQh
FAyTFmoahzEQF9ohX+9/H2zvljd6M5Nd/u+tHQ57SOL0nWrZrs8uNpPYIOLBP09oUZDgA3/AWRed
ZMOp1NTWRP9BweS0gui2GT9iVCRsNYKYJRx0HcGcpuhmPcmubEnYvSh9J1KOCrvPU36xf9SSkIKG
IdFqwmYt1emHbeeNkgeL9W9FPM34XDXBvosyDQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="k+AORB8sHhKzp3ujBxvY3HsxPfVtc9CdJhGypNd9G/M="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
bukSKaNf/9d3ZNdknxXPVrJTWAdI+t5YLejQrAyCASZA82nveT1yJg08xhd0i2aV+bqqtHCPA8Us
pwz5I8Nwuaoib1rs6hkhY0RSxSUcAlrb3WcpSGVWeY/1Z1DjS7vrFIATzzm9TMM6Hki/eCDxVd8A
69LoSZRUNJotmJY4ASIB9wevvE7p2cqxab11y2IiNRe+e2zwyW7Kf4odOFdo3n9lft9+TmRSNytI
A1IpF400x64alPNDSf/Li0K+VNoWDQskEewjcqaC+GzhYSCesFgb6e1tB9xQsq2n+FqFJIT9RUcF
BRZmwfxw9ij0S6dNkF4R5/g7lGY8E/mptCY+eQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="AbGb57O14DZSZxulp/yi6GoX9qrAl1bt0VHHOcY2sTs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2480)
`protect data_block
KoArePWAdaoZPT4n4w3qpjN0VfNQxoiZmPvkvnHy3RdW3qD/ku4PgpMbO9T36LWBYBd9jqqvhXjz
MhSlVCwVnvT+YSdrqU0hhf31s47Ygb/L56/l1F906qfzOdFXbmf/x1pDCG6WssBVDPnsNana6wxd
OXU6zCS2gAVMVzSg7sSyXHiYrMjLzJxXU4WT3RbTtOP6I78jdo7qiOH4ujUId06IGE6sKRw87gJb
+lAaq1ZBM7wwzS7vb0KxrQfbomFJPg3hK+jJjwjj4folqeDUoMnPsbQysiQAA3pjp7Mw8mTx+yCD
vjSqw1/0lyKHQxlzTCVTUg8dQBB/h+RQuNROMhBmD1EHu269J7FaH0UQ6ehSJGvwJBcI7G6AJbZZ
BSjX9GDPite5nNPDUjy3ntYl14bI+WUAbzPlzJwMSTDx8EsoUttzdW1Dcxoqx8RMKlp2XuOqsyE3
yUekbtsRlti+0ODtTIBTux64KzFLGJ5D9gn9rnSmKrJEYUxb11k9y3PgTlD6imYeEdpNBCaF+7r5
+JCaJ8O91xxgQnR9ndF/zXh038n8CKB1qQEWGGyOYKwO01CrHdsWOKUjSqQRy8IlaUP9mU8HyDzO
vv2v1ZDEj/9IA8POJTh9HfUaVLSBZYnxOh8BjaSLK+4M6mRMuSqmdu/SidQd/jHxjGuOf24Vzu4h
roNOxRtihvX8iQ5JH2DDJx44eZ/NbwErnoftDHGAxuf/gBJVycMFfAj7/4kgxl3MyhCswn6yDdY5
/bqYdfvS722mPgaT8+qXzd/RsYiHpSgbQ8p0T44amKNWhMnObynlYJRIEZAmpdQRQTdTYZBSzQb8
/aNDY2JmLmo1ZSZzjrWH/9xJ+g+Wzj979T51GgFAH1BFEVCaawenvlQbZc/+pfv2IXYdW6WqSavi
ogVCzJgZoxsNazM3muOcVEia8FfQ4redCMP7QXiyzQp77049KF/aJr20k6BKMToMsO+vXxSGBAfp
J3oaRWnuz/95nE9V8Wl9/lvWgAbsK7FxQS8k02EejT8A5zXNzksMk0cpeQmFiN6iyqZrami2lCLw
5kWgBGOv3S5F5IcJSCtt00jFnNcgsMIFqBYLDq+xOTQeOHfuu32MkD3/AluhM+8o5B6G72g/mKbH
G99t72Q2l6xawxgVPK6rFKSAI92x6j2xK/5W8gjct3RXoO7Izf4nVRv3LUt5sKM5DeU6nRoQAjb5
qQTcpkJoRxICSzAYJmeYXw7vAnaU9EijwLRgNV7gVMV96KpxDGjUADbie7cWlHnBJRKnj+Lykdly
T+tKf3ZT1nJsBH9YuT82Zl9zdNMgzySLUCsp3FCycDfpvl6CKe68qYzGgoip+VCGi1nazzkNCPIc
p+P4bg082BUA9HbgBd+5oot8XIjD7iloEAH+VrSACYFiAZHEFAH3rlwyRQj9wEc5qLiQiiF2JTEZ
5/Uojx0K0hItAMX1xmnhvu70UGfDFEsatL32ehvKX5apDZ1Ld5T2wJxQo1r+O9WqOkJsH+YscEjs
D2I4r+8cAxDY3woxhXtNl8CPvwpUBytt2HMnHj+7xtAx+9XErdBw2fE5OdECK+rtecfemmkOsxQ1
OiIiNQ588KX4Usv3eEX9sJFPEU5fdMkZGUHNIZGYMfX26XejAROoFkFzWgiAgp+Tr7gUpChuUk5t
VEpM+KS7Lc6BKM35QTyRFdVY2IEbQgeKn1w7HCF83sXYjD92+kaWZLWEQV+SDYif9AXioQwPjZLt
9gnW8URp/IoE4IdagDJjT+b8XLtN6rHBoRhkGRuJ5zbXTAQv4MTSrZ4QSQiRF4T0xQXYIQWe/qGx
8w58gNuZLSKvV5g4LGWDAEqLQH2itZFNnjlIhYEVs+7q53/Q6WdGzxYQkJP5Hx/9+yiDR1DNNtY2
GmttvJe4Rfh5xV50OKK+eqoyXcF0mdcuJRZqx8fsiVCVaNS/bHidlfAEeaazLFB14Iri/pgulkt9
qY0tno/BpWmaQkeU4/nH1rokx5e5cVaHXc/XW0dag2hp603LudSLAz6WptkxbN4dkfzulHOwcNK1
1fSb8ht1uqO66gKn0bzUmC9zdNhRWbY+WjiSbqo6R+6WR8x80+7ObeYVwoeetSmPP7AwRVhFbUD3
DXvhHIG/lFurk73nhn/pKaH66Z6qPAx9vptdrEznvBsWOaii3JRlmkTJ6hf/H0ANGAwaXg8KJ7eU
St3UbIHxrHwV0U4v+nTMifNyWh0DRx+STj47HculPDtQC0ZdqCGd1pZCSWGOEC93udXe/sVu8rYq
LwVChilheqxqT3Nyu8G0uv5MP9C7YRDhGX7lAm9Ej9p2FYH14gclOUGdbJY34QEte2YiRAkPTQrz
xjk/fvKNcNMorsrRyChnqMToCtnaATJb3bjcBNdDqBOpLb/eVXb0okXAdnnzxRdZgcExbX5UqfIG
NXx2/gBK4CV3Phkxl0ajCoRIof+ekgMIbuHICiF1eJAt3x+Z38i8g1gxKvX6t/VrWSJ8bZLoPloI
VbmKOiv3TH5uHU6/R7Da1AfOx0wsJx3Y5PDCSTeRik+nYmlloeugv2+Laq0jvE2FQjYWGkeZYkX4
/8J8ad/Jw88noqtBayGeKfJBho6e/UpFVj0FkJx5iXuhNhc2+qRkwpFI9fdX2F6AWjdkjdfEL4+h
79kJjRkkVo4pCpu0wRJ05pA/faCaPdgRhksLNH8ycRgi4/ZRrNBB3sVGGzmBqGdzXFu3yDReXC9U
RG9j53lTJGIIuamiiuiGSH49df6hVHikfUlt6VP/4XZrMq13ilSlqm12Lvx7Mufoju6Q1GSvM+33
bNB0BLP/zkCk2d+Uyh9mUhI1TeKMbr6PLELqNuolllKwx7FKSMrAm03cFQapA/8KZ5/1r5v8tLaU
ZHkZKA4mLXE4holSjMLVetAEnfOEzNOlnDOv30L8njKlPPPUJc9Aj1sho4weelJL8oDbOR3rm351
ioJAo5LN1ZDy9NDQ+2UmIuh4+eGrRLwdSzRDTwuSLUQQG8rb9LMI+ZRSHkX0+nUv3LbRIqTye+iG
l+SYfdyGapCWC9VaUFV/6ub7wK2TJ6DpAqi+dDuw8ei0gG1AQmXWO2gag+xsyGMTHDybq2LUrPmv
RL24eRioR7M5zZ43Ibe0JMVFvjsb3aubtfonlPENT/hHXWXfpnqOA2r6AtftvdzGRxdKnL2KwA8k
RiAO1uFQeK+pfEHS73VGeAwQNfwPLUJbgZp0c7w+sHXz760t4iIyja/NgbotY8y7b2DVReIjyP+K
Vd1yNSTOakSnycDkh9A2IRnl4sntm3F5sJ61NZ0=
`protect end_protected
