--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
cSLNGRxBdfbhmuaBnAEgG+lx9IIHJ0k1tqSAepMqzFNwKFQXBk9ScY23uyiZRg3BvbqfeRogPwzC
OMLEjqaFleuFzlVQM32qi4xTBw+ldSZrkG2lWTBAhSjrFbeP6RyTrHPaqvTGXwPAOsn8IzXRfcCj
U5TpQOU2v4bKS6LV0P0KjupuA2rIXy/tGXWoVoy5vuMzqxfs158zn4m5kkxYWRR4d3YAICIY1q8z
57Taa0ZYlXlt7HdV7Y126OQwHo8DUD8TYDRYH5h50//fIjruDYTjYG5vcdjHMyRuBynqmEd+Y7mh
wi+MgEUFlhDnBrBJFrfqVAo9OBf0h5asgH6k+A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="KyRfUl/xskry9SiRjLSdNMH72/1BpJGJsBcdETIxQ2I="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
cj9E6grBpSzAZMUzfRzgDCdx0qi46beIl480QRhCysab+LU82Gx9/LyJbY9sUKPF37mLNJKKq377
cAT+uYENb1/HEOAPz1nUd79LbHfdPHd0X+KM3Y0KyswZw86oSzicpKXKnayS6YI7pON0QTCsP+Ht
VTVipLvyQClr5CZOWCBNI1/8nFgp1Gc/AUkeO4rpSdx9UFlm5Kt0+bmRYMohYQb3ijCWcblxaIfc
Z7Kwc/T4ZNDvjY699uaYDPGK/tGbI+gsM4fHuZasiEvJEvBIdl+mVOf7cNW9vbElbOd999Fl9D0T
8SNejxrTU5MXVZA95eJ/z7+d/6rDv+5C1WNqRQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="+/s8R0rSz3AfCgQnlogZICevEyOhH1QFcrX+1JwwKWU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9200)
`protect data_block
x53oaT19KNIIqH3/7m7OtAwtCxrxlTCFHOd8bbWh2GsRGGsv0BmDdFUfKunZgAlj/Z2LNl7fGgak
lCGf36MB+lXXSsUKSuRzX7wSf+GlCXqgaOL7dXWYT/jht+qki5qcMDAmgFdOH879A6f4xhfpzKFk
gWdLsAZzP9x+zAkPpNsSsNGwOM/NoHj8p2MMGqiKhgOUGCT2HSa8rxOILHj3U7td9OwFPHF9tp+B
lkoWKiZBOMDUtszweDeVvgGIpTTtiviYl2nhvqNf5YXfehXmnRIadPbfq5Gu8MsZVI+ZcUl2rI5i
woLb1gC/iFa/8iERF+ZsCeBY239VnNzrQb1mF7WUbDMhWaRUvj8iU8jzjtjuwaQMrLYEL8vg7V8t
aOWFwZMiHntdt7rbt0y/2mqGhkGmTpz2gMb1W/MRYBNFGbG+lMTnad93k1Kn1swaowCPrV8dN9u4
ZZIDPQkJaECL+ctS59I2oyw5HoJAHWce+D1hbOKQzY9LfgJjZ3Tzjydb0PnJGXcpFobXRRfRQOxx
bbfRDzMbM0az6KUriota4XWOXgLuzgJ1AonDSk77sYKCpEW39v0VOPa5TbRnLbHktR750t6961qv
qzYSBRp3S8G1eqw/FAptTwFM3TOwLf/OP5KFduWSD9hl58Wo4vblzlp0Ml5UAHUZgXvZtuvHJACC
FkmX2c8yve2wD1fWM/C6InN8WQOcj9AwV+UylqIK0t1OQe6EHwUvr3xYbfKOYhhAlcEbwILgLr0v
GhZn6/vBP6t/PpmZn/OwxUnfyX18cG6knMFVzHOrlVL8wy7iy+c6VRkCCcca06N6O3hq4kkabyVo
tZHrvCtOWsslXugSwifdpqd74328JX/JW7iIRdgXu3QznW89Ws6xWD8TSEaNJ1ULj3G/3z7dgd1V
t7MwCGGzF43oKP0PmY8+R11H2+EElF8Znu2LmUXdozgN2k+ZtaXn8zRmSNu7c9hyQBR7TSwwiCoL
zSElM3Ndlk7VJ4FOyCa1DSIKbT+P9ZSsff5pqpf3KtmapcEpkl5b/ngcmGYu6V5it5mDmckO9XcC
LbvpQpJSqigY0L9BYm2Nof7xtdFYYiJtpl1KaOb1x8Dqo/aDrsCsVN27zuij+t8zgQSl3YT1zL/r
ui+4SDaFDKuvDEbwgzbC+FYPvOcgp/CoaY0h9H1w3Cj+14FIv/uM2RIEASybcMYVOe/CCMHDLWjO
Xiof0a8UgqrrtoxayD6P4CyekPipaCiy9upbo1FzgR69oOzFSCtCFoDTQ9MtncR/9GSPLp3XBhwg
6Y80ePcmA3DYrEuR0pmcqOXOTD9aKmRPqXrTxWxPjc4GWuj69e35DV0EGm/v4ZGStHKb88rib0UK
/B8KrzdU6mtgcgrYX8eE0rcv3yoNyiJCBedeZP2ZoyELGIuOGALM2D0+SuEUeE7bEeOpUgymR9dK
AhNyVg8APv7Drgz+qZt3SA9OjhUVJCeTSAFJXU5rCKftDNYx1lwoPQwVBqnBeeMG6mx/yxLTpnLL
Hx9LVeTyVEAxJKDMeyzckYSMZ2cf6AjpksJBsapDB9uJfAHMq1pL6hMOpJAXKXECaFsbkJ7sX5YR
SPN5UqbdRN+//e5R927OMvMDanQInXU23y0BV/M25i4Lmgf5sM4aqroH8imfJdcTEMn2ppg+8TND
fcLl/nx5wzG0Dacsi95KkZBpW3d6HIHFciU7tzI/D4CoI5nquSmQ7K/56U7XvXqpsNO+uOO6DwFl
j1JsAFFK20qnPQCoPONFR3twGk4G8bag4A0K+gSLpSAO/SE8U8ocWkNwCxgEuJBoVVIRMZLXf/bL
bNXuU5fd2H/OhzXJpTI3yacGrVkL6MR8DUZCEW3AYlsQqsr0En1ah6iE5iIuT8LDAFRVVBrV1FyR
gYd8JubZw2/0XEhwxrZkEoIYArdpllsEv3pdmufCPqHLsl88xWKtO2gv/dy6/NWz0myUYHhS+RP1
tyn1MOOLnMxlu4zAegOL19yp57z9wUU+zKrpeO4Ee6JBKyTP9Br/7xZPwwmtMpclTRg6lpGpPKqS
/WYoU6bajg4MYspU47wbPMby1UQYAcjHPgH3VdO0WNVdnYCiCFSwHhBehfO1PKJDxM3JTqF94ShR
6enqEo/ymF+QjA/pqnU2wx/dHOjFeKGo5W7DRS2pFEhuaAotbFD0fvSfcgq/vRB3//YO1OMxgAiD
/+MVx01zd573KQYvyBYqjmkXcErIPOyjqtFfcb9v9GjcRPeGtURDUitzAVC3fq47a1+NsOzI1Vl8
HBAwrfXOzWbPXFvctXxuFAfkYRayGy9STyHk0jSuyCCB5O/YC+qse9UR1nWBA/jlVQ3v4Y2brd8q
IAvzRDaB1oMRAWD56+1BOP1KFYFf6TieKFS9FtNnq6cPwnAcStbKHwXFHB/osX6wmOUh5G37G88C
qS95b3BMe1Qd4W/UDXlphvud/uCApy1/TVgwjO7ALJW98A/+22HDtkbjq/1Cz1TmdHnGxs7a3OPt
spZjArR6F/SFs1JDMpb5k6PqtockfbcHxMTp+k8CxKzZtLE+zZfHulwFDP+L/6MKYMOwhZj0NCjT
dj4qWF7x+0sJrbyXt8CEA1mm3bCYb1iGwG+JX3YdSj6T6w0xP4rWWvP8X6+NUPED2No4HuHqO/Bh
wocHJUZjA6pFOlcEwmyTYpwmIRYO+8H/voiXPruxhso8NbqZIsP9vHMujzGGqrv6rql1kcEOaa60
Cy5lvz8zIm0FckrMf/sbYKWknTRDqBKAFkKBmgRqmLoT5qnkhvB0dtIoH/3R9Q2TZRI60eYioEIJ
26i7EOX9CaQW49v7ZcelONfT30oN1UavrxFxKON67w4x+SWLhWm4aSEAZhhP57YY4k1ANuwqWag+
zhU6O96KaOCz6Kyo4T4UrpCMB3ajlwFjA80Jk5a8KXyBSG9wNp2yEQjalKE0coadbbLqNvE6gP2P
C2xTk3teSiP5CNVVEc5B/C2UR5t4RKpm1i57GfniQBj/sQ7pUXOcdoiIAhLXoS1xMvi2CW7fcT57
RADdvrWKUWZ/r4UO3ZCRL1WkcZB7W6c7jc/zx3Kw+xNyP1mS6VTZU9Bdo4AnM4OHl2R+ksRsNuBJ
zgsnzQ5o4kP+2+GlAx+w4Bc0hrascc9J12ypMsp5qS5+EYVm+yHiCeora5Tn9qOU2yAfhktFbp2k
7zW0me74KTwPmQSouO3KGWApcYomErqZ0aDtcWy8+Su1h67YCxgvrE0I8h6YpRkdmusK0pi1je1i
pEl+LOWMLulSyUUgRnjgT8wPtEIJbIw5gzNXbL7UDjfdcw9gBNik5TYiil7VJYD2s80wofd+yYbl
E37GM/WoBTnpJ5ddGKP8UX7XnsQ3DmSc6zSkStVnFST2b/EteEpxDkLfclGZZFh7DOJ4byqSlIgI
A0Tk+UYupZfGdCB5QDQahv0nKFyb+ZnxU+eG/iqEXkdNNmyXu/6ieX8poJdJ9y9bMSrcDPj+p4gJ
LqFRlFJnM4rom1j8VyZ+XyU/Ihi+fnQvLSJzFTKTizw79uQm6/7y9HeAGNfxTQnf69fS8OnpnhJy
CCTtUAyMcHbqRKskcK6aRsNbzjTvW2hHmmjM8LDnVKDy2xSKl3RmDXjOUMMhI2kDlOg06mJhIRoP
5whSrgcXYcGlZXgGvsvNx3/gE5T/8TzGCcH/6KeFOjIp+iMjBEnx4wF/7INrgMvojQTWpcEBKaH4
5g6RH8DDNkprmDIo2Bwgy+43oq5bNB4QjbxMGbjOhQkGVatgSP+ItMV/IIZI2US9GLfKr1TraaA5
nAeqz2ULBuXhPUq2AWGRw/ytI/tsc5LzunwMWivg9LJwznLmXnrqr87ll1NcmFy/HWUwM/nVTpZG
4XQozSlRyF69vThbV2OL39eb37EMA16CGHj1st+dWuhXxV0HfjCju/ylSOlGb2O1fn68G1E0EGqV
Eauri/jy7Vzo+oJY14mQvRFf0K+Fg2IUqmIJrd7QQPxK20fCUig3QBjFLzB0pq/Zy9XKLWir5Xsx
1NKqmJH2PF72/ou+02xxSSx5kZzzga2DaafWHfrCvFdETZPtbW6T50R9gedE/Tddb1cmkOI5xwba
IGur8qggVtknhX9lZ4+LF7cSh0uQKGAb9ezfrOBt0BLWQ9/0EKkIl6o5nnJMECdQrIStsWVMOr9m
S3TRai1DRfMgpWGXkOg+VNl2J+evgX4QYfEYYLyiHPuiapNVX7PSZsTWu4WM6q0g2R7Y+uErNW9H
0RXVQaZwrk2KOsXlmguJW0NjlTVO9Sp3TOs2HCfwkcIJ4M2ft1zDLyKcLMRaZqljy1TscvCW3u91
J2Nu4DsS4DgiOEzQgOFFNcB/hUumh8RzIlStRmQ6KhXcHi77ZrMMyFmroubFSA1D+pHlZTLpOUOi
SXsTR0dXGnJCSQE6G2i8w2byCDRLuwFkUD73te/IdmspjAJOAmEO89HRQ0uWnVKJy9ZE7hTRRN85
k3vk5dkRrffTDDDrPMk1mwmbr6HY3XhVHQ1a2f8f+hJHdop0mTaZs2tFYt3kuHFg3EvMoZWZDAr5
UeGs59mBTbuzedWQ9/uop756RxSnihRwDRxVRXilR44FKLRLuZcNAjTz4jMgl/89RfK6+k7axSL3
YFWH3rMb/GGZCS1QIQZt9Il5/++FwBK7eMXmnCw8oSU1ipur+UZ7KmfD9wsItsECGZ64Hu42mOyk
SI/dzwD29OjaimAS2Bp+40z3loLySjZKoOG2RrOPHQI4t1zrgLdpBek95LpUkhHQkY8fCcDkFFR/
9rCmqpSETD/3+Q6GpGcgllWq5Htkv/o/CKsXf3+bWT8CkfHf0MG0eut+j0OVWLZNn1rq8ZKoBBaa
cNUmJ1ilQXs7s8RLmzFg2lcfl3HFqa054POsqRjcIS8OsXkMPCxwE126N/amAE9gI7+xuc0OV4m4
Y5uM2/3dVACZJz02/G11XHsAEOrUxKcqIibnRy3dZkAlxW8ZZSc/Fzxha8DtTUVpc+gIS204890e
G9PVfrcOrErsuQwJ8/PfuxyNAffy7XjKAG74yq64y9KZ9si9tTFFmea4MPhnWgOREO5D6MCb4zAW
DAoc7m7BiGQKgp3CbyzkyDowIawjiXPgziYb730DE3j+e7zWldTKO4H41HTeBhBHJag2mMRL5hqr
/C9FLS9PWhCAQhuoSaYxKDfhR+bNWn5Q1Iag/MvaYUVs/spxkOuHsdN7Hv+7kidcxHyULVyVJpG6
9spOHkyKb6B/RCFZlGSNqTToRAjq7t1smRh6Cset3lCI5QXViGaIIExX2oxS4EBApr8W7jc2U85g
HadzcWdQGNQy5Nm8qRp+ZkBx0vB8ZCcwqQsvGtLXK7sfjGXS59B4C8513cvmMFfxn8BxdU8yDq9X
35qZPuvcvLpZNg5040uy++KKadvsfCmk00KG8v9l9f4MyF+/HPzN04aDfztL/MnLKdt88J9vnX6k
0iFLIzEOJmQKj0BDVSFM7s7Z6774J0prEH/3XuskrD94Nx+PnoT4D7+sH08bCTJbXCiCUUcC4e/Y
sp2HcdNjG9NoADifEOufPvJJJhUCDfcgf2WnEK08i+Wm61+wlFdWsuEpU09Frig694t1a719fV1T
YRS8zelzB84C4itn8mwSrjz2tXwAC4acB30+LIjZxG7x30nvi7R2T+OjLdYO++EYtk2iUhMlCErT
wXg1EmJkxSqEtYY3nSPfLrPT2LTPa4oxOr+WAen9f5A5lOkSiG+PtX8yR/j86qcyypSBntCHxfUb
P+tHRHz2fYIiA2BsGEOLJbbDaDeyGzzIrMgQ3L1acY9gswX8a062VDnuY4jF5ItlxluGH5E9Txs+
uxDIU+dw0rjU0c+jShjdIO1YSWY3JfowNgXNniLFIrsIk81JK3NtgDxP7Kk8n+7OErEIdYbL8hdZ
+ICCbcBpnQPXYL1Mpk4985Xu+ghoOpJkZRTy63+/cfj3B8k2XJl8H0+qZsnYssA1px1F11qAqrsd
lwsItsdh5bHoSLcEbQ9cCufuoXVHft90nQTiYX/xKua3BJGpzUoEnZ967hdkjHgbyDasqR1/ph33
Uib4jVYCTiWzy3m8Qdzcua6aZMtufTg2iEhvgFyqTX4Wr1NJeGJ+e+tmQL39i4Z01c11G7n5dnHI
yAc8Q9j/0Sl1eUhOlTwuHRu8dVUooCTNArLs/aL/J3bINNq7JXvYSEcvstYckvHL5Sh3bvMxgsI5
84mOrg+ERyKdREVafRpEt0/GPcvMij2oYA/bw2CxJHMGgXeydAVS0rZ+lVcacAxGpJx/LV9MM/4W
J4vITdski/ctjpx39udykPGcVNZxCwE1IziJzJp5pkEEFDJV5555G4UUW2ikhlp10liI2vVX3cLa
Xcn8vKqczh+Re00sD6ybUqXlKAnWKQoVnc+PEsLIC/PmYpPpX3g+QOTZSm+fuOnNjiGOIVTkQAo0
nzAKOKrnQolZz2JG/Do6WH4VPILZ1p+2kR2PSl+UVG/X3Q20SWID0asObMfaw9xR77k148d5WBeM
ZsITevr2xcuodqfDVRS8NgAQyHcOvSpt8gYR8LCr/5OqEyc8F6nh14vMKloYxYCDgAcLqf9/ys7D
7aDX9D2biJIFfEkg644jMtdoVvzSOoNFCqZncdbljH6PDwdlnOseAFOf6nYO/Kgh5/pCk8ByQeTC
OvB3aRnVjZn4VsCaRqC96X3o7APLDyF1DyzKXmbVqCZ+5e3X3LuSeIonzYlUK+H1vS/JkXdUfOi/
PgowUcIsKYFVKOzqGaq9BXORr8/ZAUy2Q2MFBZ9437kiV1i16v6eHRlmVvJ3PykrlW1y+Bx4gro5
gb0ORaIgL1JVV6QhJqvyzsj3VQaYiF9ERUzSnMOmNd1PUQ4hF0rF+EzyPzEeBu/LwPbwDdE/lyMs
kKOdt0quJLMoCFUTN1s6BDA0yisgwnkWoSJHwlPrJPG35wSom0uq2ouzKISPvmX70T2CrR4pbfit
/8adLiN4Vm1KmlutATs346SoLKWDCFUp45b+xE8vMJtRed+OrrQ31U3cfV77IrQQeDICKR/Pq2pv
//uxhMnSJeMaYnJeEjl6j4b0/EhDqCcOEixKPdWquLmcM2XiO7XvBo4u8C1wtYqE6qaiRK00L4Cy
oZcMfyXaltwdGEkTe19p1pjggYGQGg5JMPufUayzkKdB2vGNMUAf319a9Q1kBgdUwBL5jTd3s+SB
uJYlNyGPKkzoW8ylD2kKI5fskgz2s/zYnRVFAg67n2xofx6aApa7SfSxrDqyQuLNlbA31J3NIJKw
Q393u/l3xhkuOAglxxJFbF0Bl0i2J0eZ/V/ppCja/po+WORUb4w66sCaissYGLQcs68KKSCJbKSA
/eZKIutcpTujLPBxSbsUwnbJrcy3MoL5tLnhLtDWz8R0RQQH4q0OGSrlsLkK9vZk+ZyRsBN+etP4
1jufwlgHlYNrbGYHKMjHEJTlFDS4ul80AGTMlUKbXzmrxVXRv/gH61IXGf4vJcutWGaS6zfpLR7x
qVxP62ztE8ya1BrIv94PEvYo0h7+J3JXhZjzazG1NGHJTv6z1gsL4ksiEOAirdQKpIu23FeUpuZe
nd+LNfyJlwn0YdGnMSfyt95m2OWGFBpwFn67EyU8uXorEPhQQSfig0OrP5Q5tpe3FwDacFPjZl45
a6g4a2v8KxpZiA/HVxbdbpjIgEyHQ769FRYKpXw36WAP75ZiOfgcDHE/FdB3YZhv6Vmv6bB3LvLr
y1SrBUVGAApSCOQoG55JYV5ifYzTCzS6AprATUhVClYe0MhxwnFMk78TpbfKji8CA2cbM9Xxj6Tu
J6ybMwC2Eivl+jXo8v7pLSSuuyln5+ydSvsbhn44Ms9drEHFRJHGwzp7Odbb5z8imZReMQIQxHsF
5Xg6mBNs/MoFER4m2EyUuVPM6TioKpdw1nmJGw79lMfLlD9x7FZu5GDA3iWczB8rPOEJVncJrZJz
B+nImD1ebgc1PdHeOwtIyH0GGa4ISFmbuL0LjUAIIOJFYf1QuVrJpC4GcsQ8kh0rEFXr20p5zSan
DJzKtxbzaFgrxP9P5B50rnwqqw13ofXPISwrrensOSDx+PFqLdwQiKdEBm2BUUicv6aX6yMuznp/
4jwDLKaM6C1xieiWnTx6gqZB7RhObvVjbTXGSL9/BtcU2oqkwd3lB5uKDDWNoZ6Havzl7Ieywyah
pMoe6AAZJKvpOd8V+nSK1N1akltnHC1MxFVal2frDHbUiSo2vbrP21ysB2KaKzini/RR1cCEohfj
MAlnUKFeMsj8mitpOiBOiUi4rXb+ddjNr7kQVMC6eaOlqO0aJbCpgnm904hZf9JN/Hvyvsu6bu7+
bb5jy/xF6KHB+jVHjgCKnOkT5Blc8HL42rz91E8nhSJwpoQexSRWDniZAmWaGUlTopbl5NcqhBcs
r19lEVcY2f22BTf+sndWyMHxl6b2afOtqLoWBpxE1JtxTtNi2OrYm5GeLNAcSHWSqwHy+4N3O06f
fKuTi6x1ARBQYP0k1VPbgZZWFw+lgCLrwYwCPeZYVNPCXy1wtvyrmhBmznjBtw9CnsG5g//zjV2C
DFBJCUC3pbNog724edDIbhd19grC9ulsP+tqkX1WtK5ZoRR3xqtzW22+VnCBkwxZBX2aFcNyj9MR
EUnscXYvDBhAOlcKwfzXAoXqQMfSb5uaP4Gxnb7xR/WbY8RsRrMpoPAjqh9H9I0q3OMVY5izEIvp
Id0JvoTSQPrg/t+01cd8K6M0E+n+5oThRSh28nayP/48kPH8+vibAMJih3co/VStPUpEQlT3oTx/
mk4GBKV5Yc+lBlDG+xMXv6lIT7uoPCD87C6v7pGDxH5GQV+ofj3aCSPIjiXX3+fx8L7FFn1Bl9Vi
y8hzJzZjZeAFfMGR3W0UoTJvc8CKMeUIdrGw4anQmmQlfXdnEvCb1eqxtNW4WMwzm8hVzrT/G47g
PevKFw9Sc+/6EGw8wkiZ02yTweh+C/5Xlvao5v6+LGqYiLsoWwtKphTnwWyksj4yhCTUJIKzu8vY
rka//fYIr2vzRsMSbBiKZvKO5XfAVPEKQ3mQYSOhUttgZvQyAVkr1JhpJPlCIGLUWnjROz1MrS0c
OBcHpWwmhpq2B/ynRffDrN/kqfz/Z29vja1VDh4QOmLGOPZUtfxPnur6s+N4HzrjGeDaNO40XgtF
GZzYz19K9go0APZamnTeOda02HjpzZiHNsq8C3zFQ3c92rtG2/p2t3G990vuDZ0N1UQDqCA8dMnf
Sxpem9axnGyRkRJDyfwt4SUyri6ljOPT2g3RGrJJYpVawlYJIlUPSvaVqxfmCdQEg6P4Eb9etMET
8E0iB1+3FgJ3jK5yuXXz1XS43BXUGQ8pTa85cVoJco2fODQuDutGVWT8ELvcHj4YOlzSSyB77G+g
sfrpgI2L3D+sptx36uctqt7NfBvYL5dtYudC8HjjUQiazRshbPJfexrrdQLPNv9sTD6VYokWcMBH
4cWs85YAb8E/QwqFhmETKDMnL4fl681MmY/sSJtZcoerRTaB7R5rDSB+zpw0/J8oZwJp31xmCEK/
DX5XzsEU+PifUXE3CMJ6esuWBs7Ac0mkurHiA1Jl+SACPgO38g6jiVaV9QQ68p/fynlrLEJ7RTaO
MJ/zbjt0Ivq3sqd57ZBCwtpr7GHBsolRFC4ew7ybWRWVA9NWxekVyu2oILsVQM5bJD8ejelA80CB
o59wjf7rqyBvT1mI0v0PJ4Psh5jDDVqRzHhjc2ZUCxI23zViya1I0tROFGEhBFU1Q7m8eo/WXtM2
tLca3fa7g44ZavCedPz/93afNdclrkPJO4yScCj3/mFS4ayEK99iZQhdemLeaJfYJNE/QYoGz6vE
+KW73UB4TMhvkoyDifxHtMcqPbAQAeJb8WX0M0WBDw9cTc1Z6alEtFTlf7NLL5vt9oMBF34ss3Gj
isLnafMN54bGRZ0MGA8z85MFVc3eUQwYRQnjIQe+VDYneX2ll2Zr5cd54oaUtsADdjmyOL8VKSrh
d3r3yDj/sk8C3su4AB3oB4SRjbyfAXUG0Nlux0L01vfVe65kV2IHZgd1icoRefERfp2ATmYu1NhT
49+1CPzYZ+GJAHGhUr3FztBl3rkDSmaqgRsneaT8jwfZyMns4wUyE53hPj/7RbXimeK4b/W5XX9b
0e21dRCdb6rFT8zvjZCxNXGrrj0HYfTyHIIsflXYpISfkxLduraqDidmJDnpNRD+PNpDaU0Y0aYp
ebcwhzSmcTLzX+okfrbIBRShcnXL60Qg9DmUxEI10fLhWtLVyZu5ziUWhxaVYwVNtpa2pDvh9CGE
GfZuTM2tYNuwVIzmnBeiMIjjpL3Z7K1zhuJrniOfuoTILE5H1vSbbtz6LIZpSnWBJiXAvbWNK6Iz
8b/X5urIugXmibUekQvsI3pz+b//b3hNaCmCzN766S8wt3Ithee0Mq1hD9+HnyxML2opjWDEZxOH
lFi8NaGP3+IA5wqnhK+yD0zpMc3l9wNeXs0goYlTs1OSu37+OREBnZtPaqaIji/7Gn1JFqFYNFjd
Z0WoJ78fTvfE0pFJZfQMP41pl/nL3jYwbfyZLnukzwTpNEeDaFSCb5yLZD7ySAUzpdS74Z043M4m
PHoiZBE59EJ3wS7Nc/dTfqNUsShhTXtH4Ag7LgHupgmvPSGe4a1vnJNKOVso+p8ORyI/UvMpNyaY
53YLG2va+2xuH+x/2qrSV98EGYS+g3xqOB/SuzbcC21ZlI3FsgZZT4ElPkHXzbFnIq43r3vWct7k
cHuAyAv2gJdHnR+6HVUMrKiLbDqiAcpXr576d9ecsFh1hroGCges21KYsd/VZwxEOHko1xhoGO6f
FAltXLe9N4mbG/97ueBlmJfxCpfnwmOwuc0rq4PQH9+wy6XpXTVGSEMQyLAaKFIshTNh4cxiH4qk
19yQhHEP5QGNWMnDOQWEANJD52MVZQv8tMF+R0tKWHyYoJbRLKynRFvUJ2VnhffRxeovupSyMqNB
5w94hJbXvdX2DDcgddmvCo6GvrH62FAmhulBMXLx+68hMXrojM1vHVh0PW2gPVXlgFcurHR+9u7z
g/O9Q5A4WMB44vzKdhZyWBVovVZV7H5h4G9EGfTe02SFCPW9DpbcAOW8f40FJ3EfK/C50/46aDWy
/dzaToiqiMXrOIefpDiqmVCTMPgJVK/DWPBTPsDYwPO8EHYJK2Zv9cupq900veQX6ckGWekBhthf
K8VEJnhLpsgTvkjo0dFBcCQDPaAWqx6ci6tzMexpBQzaFmXM8GMCCn8P1Pmk1Dp0CKgLtwFA9VOZ
sO7Clumi1YonQbA/pN/JDUr4A8YS9hXyE4sZtaAF1jXULpykQf+Xvrcn031tjv7F79RG07o2K8/J
ZZ84/H+81lwIvb9nTPsEGsYnL/TFsPK4A77G9TboCLtPYm3UdI/7OEnqg39cBIl3IR0OYMuerFQc
tmsoV7FdBbWUaaRpX4r2AEaCGggBsdlaYwe1OU8bAw5it7KfnCTfAPbf9X2Nsjd6RO9u9UnJjDuT
2P4LixLuFzOxV2H720C24yMs+s7UwXI/r778JZk1Gl54c2uv+FT/D8iElkoqwP1+09iYrnnNDywT
7kjBY9XwnRp/R71mVd7XHO4g0eUkEXNi+JdIYP7LC/AkKpoWJQQ9zuLmGskSy++mJRgzonVf4vpw
/MKBrQLjgOSw7/3s0vbdUj3PvCAPjmJVI7mDfhMI3wGzPA+6LMsNVJ7Oh3SS1fqL/q5uRUejS+Ac
LwMN2j3XI/g9gusflkL1iXSj4BTosq5Z/sKr0URdtCggVZiKcz1EwExwkf1et9um2eJDMNT/2m9A
aEUoGfS6WgNfuXAb1gYmt3x0O/XiymQCxqhcPdt6udWR0gcJ9/mNx8LoCi1GyqYWIQzSiKaANILF
7ohjsEmbbwH5e4eZ0T1CMu3lcUD9JkUtr4y2p53MQamTnScO2usyNM0i0DUNy1FgpyyccIgz1bXo
u/HKND6qHj/+2a+UciObAw1KS+Puoif4jakG6AqlSgYVxMlapZP6ITXQolWm1NSfM948BwYmHCDl
Db6VMa4wM36vI5Pt3zV2OBGYbV3ZAqToJ+OH+psHL+5izNn5ErRZQEiR+3Vt2B9h1JdvCCor1T1J
+T0Kx1npE3fORlrVBVwxJUQ7zWDvoHy5VJMdyLrSj4rEbymzm+DykTtRTkXkMeg5ranmcTygk+/Z
rjPb2nWUamcQUQJNJ0nEO696IjddfZ0=
`protect end_protected
