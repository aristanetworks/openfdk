--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
TERDzJn99D4ldoGfIp6fWInlnZgyq2/+XWE1NOf+LxkJtCgj++o/SgJF2LXvT0By1zXBjCPmLNB6
hE0NzhQM4kBsl2hQkKFCh3Qv6YdrgMCxsBCr6dHH+YADjygiZwDOTUZyZfwsw874DnOv8fBkdeRp
aKwqBRl6ya9pW7bcHF8CbYibmes76rbAU5RO+gaP4dIuH8zhZS6SHQi4f6KDNhWu+8j27XYFLa6u
kpcJJRiyLWS/Sq0kIpYIrhPGqQ8+MHBWJ0thEPj2Zr2DAQ+uTcDmzNDqaKaLcXz9GUuKap0yYdde
TCpz2I/ban1l4tF3JAUkdmTliq41RTzTyUp3Cw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="v1da8zcZe495EdML8eCf9IgP0CsqR90FSrPc5K1T0sw="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
MIbyQaiDFZP7sWIYMvMuTjrQaa7XO6jrHWZc6/izhLttj9qL/EWVWynergcv9lwsqdwzJTGpM/Tv
KqKsI/sb56/3uTA2HB15tc65DyjivoSqBEkvopOcGDhcKm+KXccLemjNDlp2eanXQByz2J0dGCBv
88qzRCjYlbg+vhS3jA7wQPRqLERLoxdvMiTujMAEegRT+KA3GY5N19MyxCPM4Q4SNDS+SV9zmkC/
bbFHfEQgs31nv4sAUzhkaSBixvdBDeUs7PJ2SuO0o8QfHGp76uUo1qWCNqYBaKJd6tpZ0aEiRjgW
E8vB0FSfaPL84AXoQr+EtKXlK4eHLxB3sCMWUA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="NcpJ809iTuJae2i0v9LeYE7sQgOI4/nXFU/D+BggMCY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6640)
`protect data_block
NDDus26/bjg9tK/Kgf4kchugtlT4wfBbJ82d0qcbgad6JPPdevv9w9i2CK1Nv5NKcnjWvMJjcAyg
uNBOXiTWwtcfpr1OlZ0hfQUF8jxxjd+/OaTZVrrEQZHfQuMmdA0Iy2Hb2XJ4yqrbWlQaGqBRXppJ
Xh5oGbBkJuKF6GSRA8AdSiGO3Qpqge1oIf7IQlysEC1gGeQgx5w/uubS6pq/Jj/TJnKOfHyW+Ru+
TFI66o/QJ9sVdmooFWOiIbedEEMK5i92AUI6PivaV/V09LMtE/1uNoTNkEquJEiUz53nMneh8caO
5u/kkhQEd0axqjLn+Qds0uzVaBl/G9hWN1QQDCBLSwAcDFujT5T21mxiNDIcpkRCmuflQXmbleEr
kSLUL0pt8a9blgLg80x1tOWotc35/0QrkAjQ+M5MT05A7MJJTQnZp5VuR9jdiy2pm+ZhYwkTnOua
l64vW68WXKFP5r0OgcNIzAi4y3AoqpjWnEijrlvnHHvoNByVNYQg9i1xHc7DBRH9r/IP/8T+XU38
b3NDrCZEIaiC03tqUa9FyMK9EyeBLsn3f5ls0oE7uzsfxv3H196D/LwVwKUn+J7RMr7KuYLiPZvQ
5Jf07DiI8jGewdL22tSIoswA+vBhvfj8ha7aIcVziPrvd5eQbX8LvKBcdRYoQ9J0D29wMWF09WPE
kY1KtpkRlSSlpmzrxVCPWrIuNkGko712VYRszY9R+8gkbfv1nhk/amchI4ix/r4xzSaVm3dT7KiP
MzfUCTPugYbaNuluN6Qm4mcNEpmv4g3ZPLXEb3EB9FD6lwta3bVEuABxTcQEikf5zOfQ5MaPfmmr
Q2rju2dhQRAi7ATDORxxJVQtKL+zI7G7xWyQmQo4RlzudM8af/W2ogcbL6JsmSmKVX/ro32/Q+qv
eGM5Eoioed7d4ZExEKTKG7g+4OvyhE2dpwKxa747fmRpwO5EutbAVy3ukfy+MM84PycxxM7OTJ/W
6Th5vA64LuaS81rITfG4ADz2OWZ7QAE72ZVLGBLDZWbr876qICem89PY3nGS6LBFshji9vQEIP/S
kra9zRZdzAyGGpoQAmaJW4dRNR8bABpOCLaZbsET4jDTREirWVcQObxaIZC+/Ux3+2NM1ZaaoKM+
q68wV79gMkJckE/jbGzlg3L+AIIA4wMb1aypZWDc510r2D+TNv2saw2hfw2qnT2n5dl0D/bPiQFn
mqvP+kBrEl1mhAWXVMmPjMu3ksUJuVBeBolAvmm6Z8mx506QQkcFbYh2lSL66mETNrkufP9jcjBe
dQBenzKkn6EqHR/9/eQS14vbFHRhDYTZN8XnO9ngVX6dmTaZZbiX7UsSu+vXnCAAM0lgDikxlvCz
n89blGAvxeM32brr8R1ZgABzIWrUK1wj4n2S6p1ZaYtx+344lrquMdo7zq+eG3e+6cAsXKq90wFE
8PxQAo2jdk56rfYN3/PZMoD4RRF60BRFqwV4tN2qEyxGUHvfCZsMJiYcXYvQWcSrueIHb7LaqgQn
sFb2gC/ZDmEQhheRoEwJc/tnzTyn6Mpa33YbYvM6wBCBBQheJkLSUr6zdcW+jj0q7cgjA/GYVcwF
eS1nC/zXpdvQt6XOkqV4+d+QGd9MX2seGOjnTnILxJxvI+jnoDqzGxaAHe18rYmfO09IhF7TB89w
80eabAY/w3/Z6d+95q6MDbDnp41omD1DVT6SqomP6F64Vs9RXPCRTE5jISdXIIfZLE/2m5KAokQa
36kuip86n6vrFW77rQajf5oNTZjG68RLCrgzHJNLs4evEBPO7KlaBnk2o7wvQX14D5V3KIxr0Trp
1BN41T3h5kZnblsTxcnn57/32yHGSXnatXX5/M902vclrdn6DTJPgdyefHhgdQ/+x6+4HhWZqFzA
PReyivCczx08d0ooSaJQBoVrcs/L7vFWUpCl2v4YqEZCrZBXDIvhyR+UsXNzBle5I6DI87vJScrR
Jpcz4ZIKldD2SGGDyx/HbIuXEZtsdM9CI9EskxlaPr4g+LronI28L+yZ0be9fiyKTvH3ESJ7cUYZ
cCMOLppcD5CHR+97rRW6/jl8pQdUYLqyi/rINwQqgCIfSAklkgfLTGoUdYoXBPLhPd5EEBLgSfcp
Mi22ejl1aIg2ZxZoOIDR+UowTn81723tCMVItfFXoUwUx46qPzB9R1xatOm3WlXXS5rF8dGhygw8
O0CdflV0AYbJt/GOf+EQ4krdKaF3GP3q6PGlb97huXRJ0BOPBJ52yDyHj6ZFGnbkHWSALwyBA5kR
3lwI/u3K3lqIWcdFTlE1a0byyZy3+9/Fc69brTGuEnxJc8GNnO+J5HDrBN+8Bimxl1pb/D9AnacJ
kBmuGP5ygcOJFdKPL7Diriok+LGFazYsLZUo91tlH5rcOjbfBrS/J75csTeT5jdFxxdwmo+jc1GQ
CubgRqw/DTtz83gkN+YAhUCHZerwod7UILkHPtTAB6DtEnh1g09MZ37+CBIlyNNRIsWk3TGDNcoD
FkmMeYWmZqIPBsYiGp1RwecCwKHHHb7UxoD6MthPAnEecgXdn1S2ZqYnAeh2IlOifkHSrf75oE+X
OkgIV6WTy7pTG24Cre/PlIn+OI1KEGX0pDYTifKkdBoxqdyjnupHlLgW0s79Mmpi+T+mUqcouRh+
Vk0bBjuWofA2M8JZ4kRF3sh0rs73cvYq9F3KLWzCmidv2zRmryfKE5S9p0OSnD6hlwLGoAJSfHlZ
ifCXxx7bV9YrSNU1btZqvQk0UsbUFynoC4vQrEFATQ6T1qeisC0rX29hiK71AVjBjJr5IChRQ7Qj
MU+/AgXEJ+asI+LGCDcf6Ju5VEVAUhx1OupK+tEibWSyL38FzFTG0ye4jAq+FmGTcj3C1VCHd8/h
vuf5xiMbCr7G+9NRK0DyCCEJoI9eqiTi6YefCA7xugpBvNKNv/JC7MJb0evXFMtVi8W2Cin4y2fC
noM1w1m07s1UrXr5n5oQSxyKvOjatCxNFKjp6WeK+IzuW7DjM18ISgyeX0u7gyWK4oLnOkJrxr9L
5TgbBg7tpMGZOD44Bnenat8xb+Em17vWtxPDCfb5KwIsIxdQIb3BNUoY3ZCHZUwODeH3HYKwAvMM
6yKGiNNso5S6ka2/H5drMzYqVWYw2QPULUMSg4hxQvywzT8awZK6sMooaawlSiIcezL+lgLO4wyQ
NsZVsPIOCYAfiDcyic1yFSv9LVFWS7qWjRpuKDoooVH4D5eIbQdEU7BK9etVNqAyrEA35GnkobaM
NErwxN4Q5YNZ7Pr2m2kRCmEbjEB8/j9RzW477L1lY9GILILaYZhk41MxStd6pGPqC77cMGa6jhTl
AUwmyHx+CuztIuDv2RGqkEKcaqit6brP5PFhYcRKxUMqpI1/WsvMkM2KljMvCbVKqjFIW6u9QS9U
26pGXL/cGUSHTpLTAex5x+2vPPml5i2TOdZnqSUUGhj4/K4EJElxqcOcd9DR+QUZ9Omb3MHHgxnE
C46kGoDh5gbSzAqKxUhwrkjbXKU8A4Q2Ea2CGBFttzWoWqq69XJ8TvAu4sz4R7QX7ELTYBowAGMU
ohHUPFFAwN3R9Z1sb0wUy3u4yaydfOD8OnBL4YNVkQtf4/ZsnulfE9WOwNt0tA2XMp3IBHRHC4cF
ncDsxb2uCFKzPtVRgh5MOBSgEq/3BsxA9A6vTi0DRltlWz0Dz0RN2aBc/LV0Bb0aAxAX9sQ0j7r0
BmaUnlgpCOmQ3a/a/YXYNQfOth0bEfshuo7oTere2N4dXDK79EP69hEI5Si0EjDveXtUaggc6fD4
9hLpBC/ZyLKK4AnMISjUNVW6B3q+ZYSqUb2RIl++0Q7QfT8g8S/M6bScm4hbaE6rrTajGSGcMGje
xgGrQNHn4dGQTa4nGiwyTVS+KRp/XdqnzS5t1QXu8MHkkq1W7HuIy2tkEIAa/iv5MAdqSwRyyKoZ
Tzk4iMYGyYCPTSYgoHpcDLS8GpYeaRkUA4u/2BUHeLUIiXIvMJyQC5Ep+j6HtknL1F76JLqJaqDQ
oU5nJHOX3i8qkl0Qw/sJDi/anobAaymUoosJtNgjjfiXr1kKjmIabN/kxS0H/LmiiSdGPsIcpxJk
Os5OAy1bNoRgRaflytis45QZLegUcX3nIYlfGNnBoB/CLOaPATT8ZaghnI58pCXFPDq2BEn1a28v
3YKciVwOrI0wwJnnkpLWKLALoWOzjIyAKmXMsPYVrA9Xx6pfSyDwMxjsKRKEvjLZSNlLuJ07zLol
zLGAnEulhzbFY38CfBsrEDHR6H2h17a4z1Fq0orZ2QJJoKaC7jdpDugCqydWFpm9ZFAhafMcBsln
I4VOc0fi8mq/7xLtRW0yVsdR3bMzxW7n8n7tIEl5intX1Uu29j2bPWRtAARG3TRxg6KyJYyB3hJm
oDUeqWNmN/5zNvcsvjFNcXAmvgm0ArPjv019c9sAM+wBJtQTXEN4f2DUga0hY12AyeVrmLvy8Lr4
hjEMNHljIMmxE0ujjFbMwlph81lIKqqOH/4Efyn1EbcdDH8bg5gnXfBSiNP41evPBftG3OFYCCCQ
24xO9EGDMQdFFW9O1DB05Wlcj1RlLOWZle2SYnCfwvkZhzKRkibM/XlaE2Nh+Rag/HAd4olpt6sV
m8IvNCCWZT9+MmXmeeWY20kWccSz2Y9FUxuGcbfYlRGFOQ4+KAXJiEXrjnMvsCEOkoZBAQFSJL6O
czvXDA0+q5cEkS4JIyKcupX82Eo+3pbm9tbnJdqeNObUJv7NhVrEIZulxcjE/tFaqUe73QW6uBHl
jaleohcrIcAF4AFkrzu68pkrQ8138czWcIZ/I+GPXiafx9ONukOyRlsQRPt1ipKJ0oNmbsluTcnp
JSAbFGqEH4XyoEFrLqAcozEhc+pk8YdTQ48I//l/rpdHmyD5nuxzOPq+WvTI0vEbviHUmTDLMY2O
NEC8oPT24BGD92lMZ80ZvjaKlLujMULnkuLN+5+hKIRWSqXvKLmNUopyK0kdgTvGNU+P6Tdp6mKP
Mcv5o+2FjDspG7Wbrevqm5pep0PUl+56J5LQm4nWOEptpzj6vu1vexE+idaWjS7hZHD7E1QlTq09
SwjUwN0uAbXmji9prsBFGx745iW1XLDIEe8M4fs8TSlkoSBfn6Rz+2bE0hiXALBBOi0EuCvrrk8Y
AonrR2jOfTpMPTMQjvnWTWyYovbXY26EY3C33WpP26fLFsHfGjYvKmAJ0KKKWqj59361kTQivPj8
zp/MoOJXsmIsuvsjRb9ra49EffKpEXMKj/9GMS/msWCiWtbAxjs43IN880ZhulyIXkiDWnAVvRBe
FwhJJ5ZRnK3cO4s9g2JM9dFrYe/dz02//NEeDy2FRK6rELU5oMq6uF6GY7wBALLkbBbmQI35+y+5
UNe2A+44IETFLet/pyRpmiWR0gRS4TqX4PT6ltpyeECEZZ5PmwcysIwy4oszQOthA1ditOlUk7MJ
lvIEoBpWQ5Q2Fb51Rc3xHAaCioxG9guNwLokV3WH7cMrC9nmc2npgL3WvPWJd5wwtDukWNkIgRD8
ZOFq8SdJ8Ry8DzDr15+9jS3ZEcafAB8rNjlxLD5Wo9YoPChyUXpS4H458MtpY+whN1nsJ/YIdgOD
YueJM37uTyfXQ9qKKbm8i7gpa11Tv7UNDofcXSKSHppA0SUT1MrD2q3Bdq7p0Qf6/1SW905oueXs
0vMb2lgMiphJsLUHZRGEtb+DzirvSxXX/2HWZCYZ4vxQMn040V6KsRikyiPbWealyYhAuu9hZOIQ
udzYN+l6OhV5cbMD0UsuZPepy+MBfkVfnqn4aCcBjdm4anVN1K/4t1ERTf5zIDolyF2cKLsa3jJW
5n9DQmmaSnGJksU77s7hghOCVUiVtjlSScuWFHqgFcb65fEJp7m2CKt1GIdnC3ajC8vfX6FPHa97
Jz3r40fNGJ6aMactHlZQsjP4x8Jv21zcRp2h3lqNTGWBAe1yU417WTLabEU8FaTJFB/FMS/5UMY2
wM9yrB3cVeEvZQwORkNj7600Z1w7Jba62TuUHOEf7xOkdWhlyaGTasvTPc5b7PgjcucEihwZk7JQ
kcg4ksqUGKCPQTQ0izgHgxRFXwGJ7UmrokUcZdUEsf7FJX2B1Y/xAQNDtG8A2iyeN3PrVR6V6h49
S5TnRqXcU41LXTXD10f/vaxxH5prICGpKk8SAW06piFGHaw8cB9uWZ4kVZgVzzhy3z/BmhN07FIi
huRTZKxt6FmnlCzU/hRSqtPae60g9yPVjiYTBQhJqeuDQ5VSFhD8Qn2zb8feCw6DwA69D4Tbzcu8
V6J6MG0xY9Zl5hcWjD1iWYOVeKRN+JeKSYVMhsW8+MwmvIA3o8hhPnMDknw97flxuGXAp2Nte22g
ySSiZiFdmhT9dOFcLHzM27Zd62HUoOJ+sfo/X/VGRMbtxY5L75JXQItErgFDdWNT9REbXuUNUmQz
s8dftoCofnsXvyU88/ZBa0/MssU/sHj7+ki7pVzOjIc2IEuhY/c7VnTNxLG1Rbg+wdYJWKYE5qRs
Sc8UTK0oyMKt+ZNtXkUDoakg6BOnQ5G2QGo/77WPS8sJ+On8GrkKAP3s/4ne8z2loBztu3XzycOk
tgOU28vbhhFaNk5RAXphsG/pq56d7Xrjv9HVsJHlmxUTks0DOEeO2izko00UhEZ4jfXVbThYq+H+
N2po17I3Cp/1pQxMWKcCb2HvDGnwf2hek2JsHtXYz0P+ti1jyjibXLB6jgFnfPTI7mFkcBbq97mQ
M8R4+VogZaZJdGs4F56EezV53PhKmj6yaeIAJVvg+0Svj8zYQ700rYEHzEhyoE2FC3qARZQD6hGl
t9N/tOz67WBTPjl8SCanqJMWwZUFALaEMDMMtF03oYj2AHPUXrK2hFWPqgelKBSUICD9B/iD+7zo
NNWEojZ9F2n22YiK0/oCwF7aKiM2nb6IO2At9wWxUO1jvbHcAHOV25Q+Qo+7GeWkbwzwX0Mqx2Lu
mxyiujo+SpA4h2TyMaoU7SGmCujmv+H27p/QrC9Trme/WIaIPyA8qC0mz5nKMOwGITqoHMtZu2Ku
3HFRgtxCSTbxd9jid3ZaSh8KOyTEFcTm1Wm7xQb7Y1OarW3Cz+dVSm+bbdXoON5HBAs6bdHHEXho
AonVCu+qjqN5Q6vueFm2zPwJveOMKsQ/wH8R/07KE1KxR6IKMO7XrQkT7kTsr//LmLkTXwozhUf8
MI5Ja+2f8KGPOERDTtb7GiCXkxJ/y2VIvGAeQzFWxgf6j01DhOxiphDJh7vkjGNqHcs7lvzDNYCJ
12ZJmvsYpYUuCOS36m3R8bOdhP9sKxv36akBij4iAI8cf0pz1LUUvfvUfZl5eEQMb4rXHnRjy4Yd
Vy+F9m8ZFYFNlHs3Yrj4txFN0bYK3YfvAVVKTY7ZVyU0mW6nD6tXHSFOzZetlbV3lhctHNQfj8e9
Vj0LuGuW5kJ0aWozoWdz2h435/RtJELizCU5KyFeg7PkclIACZmu4TC7N7AKbq0p3fHQETGDJ6ES
BzeQSGZK7LS7k4ZxbbV6sHn4s9GjD90WkB1JzdoLx70I4G85Ame0gwrjKU50tGtHeA/Jy93sX/Cs
p/lkVuyMYUNE7fpOfYVuqvNDuc5XQh4wtQ5s27Gj47c1cxTL81V6eTUTl8HCMwHmCZyqOoYGXyEe
VPPVZ1WoXq6Xl55h1fymCmMmepqMol9VsFEI2UGFeE3ocDtxHUpgFoEG1rDoWEa5aTLsNr+wsTVV
YmD151i/GGcSgR6lEeLtPWH8pQV+d5J7p6+fTrIWi5CSrbe8u1UDyxq8FrZELByXGMvTd+W5bTPs
juq5YI/Kf82vyJCCTDVwyDxQTSNdMDwm+IumvG9w1UHLBAyPyE+cTJ0VuTp2yBcAv/ShFDF1dRHH
CwTzuaE9r9GC/D+lC7M+lQAIqdlKY+AKK0UxIJ7+L32+Ve9xXVRDe2603lK+JmGS3biuWMKuta5m
nFjw9vyroYywujl7/KYHui1GOhdZGLk7ofAzKt40Shxj87B+Q6hmsmOPn8nXeXUXAKScDS6whfzn
bu+96M202vMpMr6GGWMGPXSqeSjQLVLGl18pFY2yt7iVXikStv1NaN/uCM/UZVGGH7JNRkf4LnXp
osgYsvA5iaOCS7kOh4ruTII4dGNZNwcImXRSmpxGnbj1wmyPuYYuwcoin7BwlANuHSlFYH4cw0lp
rDqmQhGCYFlLBk9CvNK75W1kKQVAMzopqzDwnyn/mXRX/tSN2W0qDc+OBQPB2c0Tukqbm/fkCIhj
LW5iVlGTuIRQFZ18G0qTWQ13OoO+3NedjlKn2YYLvsGHgHmOBWb/up65WPcyvtNzcYXCyIsqxdK8
VIn30TeMbIF0D0Ay8CA2TsuzZ2J1jomOr3NBVvXTWXhDSacVDdXb4PrdnFDt9P1kt2VOG0MBE9Ja
N1oXxC8TWH9Ek9Whu/uHAJBNfSKpV4C7geQywi1M1mBSjuKcdi/OINIKlZrL2NJDDQFlsN81GZgs
30W2hFjuB3GxDdsVJO+HuBz4v3kgTrsycO5pAxePQIAJcR4XzG3osgpm6xWOL1y1EbSYSmPt2Dfq
e8Iff2/XgK5SMrSD6ABDRYk4d68ojgxinAwfScVsHxBg0cP1FfUxMvSgq7k0pMkLhv977GnsNPAF
yrDOy7FWtapzUYNDxxvsu37ShYiXJ5wnrBIBExitnVYXIcirHThO6KWSbIh8uBBKp4rJhAkwLYQ7
RIXXFfueMc57RWMlPZ2IoV95VSz77z3ZHccye7F7gYcdAZLuXjf4SDpv0+kGAkjx0nsaDzFCwgbR
rTHeM+A0/4QpKHtp5qjHgXKCsOgP7hgw/BScVA==
`protect end_protected
