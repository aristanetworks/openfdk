--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
e+0TowDitgMD5gyFOM4BqVHKpEA6OBKvFXVF7YlGLXQ11DpmeyPfrX40DXF5j8Ati+8OUpK4UNo/
QN4tKAAPLhuGBj6176NBSgs904McTyVtF8PFBWozFfrKHOlcc8QtY7S8L7oJWm36TCg1XVaYUj1c
rGwB/65lw8bM+regytG3RFjq4NqKPCRFcCF/p/QibewZ5Zj18GlUD0we7iu8VO085YOrYH1JM5nl
PXx4iPlZRcRiMPV62H8N96X4Z1+gFSKVDsioy3oOpQ07PXcp3ZNDlgWzBehh+vMe9Ek5WdxC5GLB
UsW0xHh6w0BSceZsF8RvB1rPPEtLTbHiQ6Q3RQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="7Ypo2rJS0iztnK2WHk4FmAlOrRK+azv29mlXJeeRh20="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
TVDYVeTNvlkpYI0HphLalQwHTBWaXi38AgCf126ozrVKRencMXXUbYoaIADg5zr5P6qbpAxRGyaa
GtZ1vOnSf1ABXnYO1ze4+cRwu0lpei/BoXZOEIfM0QZFhZ1Lgj6c75/fklpriYNkdy1fZkouG1fs
9vbNfGFJrHSOYcIN1rvBOQYYAOUnmyZ7POmtQDWVAgr9wTbNtBr4K5F6XM2G7UlAewcO7X0a5go8
klq6rmV2zTQ0y+FfOLsWnNs2D6NQOPu+GakIDxhMOfw1Brgvmqq6vSDggl7ZJkpRg6/EdFZoMIGj
v99deX2xztgtZa+iD7TpELnBRwXblsIhqvAf/w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="OF+sGecY1tRroim8Gvu44xcd64Tj1fgVw6OypcsL9AA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10384)
`protect data_block
N3gwXzrvehe4NmUb9D3HFbJtU9gXwMkbyCrFoDOP7skIjAklbv6Jj9+udErbVYwpfY5ZJOCXUliz
rpl2LlPY5ToPBqPwEp1HaJxXBcMs+ALcTQGV6nWMl+ZhtjjrESnfoLUk6Rr2tOkHMCIXdIwiI64b
Kq5Iwt2jGPDM6jUomPc36MQLU9YcGRoIHf09n+ysxcz3HyH9TZvBV7M5q+2lHD9Bglxv0gniBkGy
aqTbdrKSccdffbBwHRULvJq5sNuYMpl0GjGAk6h3OcQ2zOEAVFpNQ64QdMkvS929deN0CQtHZlzg
QbO44auJhoqJinm+paB8fLciEwKWgaua56Hpry3jIgAqQT5pf9XdMS/Aj5H+Ze7H/PpxGju4eEBU
IVU/2FvApKXHNWl60Jqy4nPaAsos+UPdJqsBExjE2rekX3OtfO8X5zUh2Z7SCFd89nmQ8vMDbjSv
/G9547UJAgiCjbkNZZVlyfnYBgqiLg5P2QoZMdyyVPhowMYqSCsN1Nki/hEyrN3cPfbywknkpe2+
1axhxJhBVdY2YO4JG/wCdvoaG53d6IJ0Zpzykt4Gu2P4RbYoUkNtjWtISbNUv6OKls0hXRjfPjrJ
061fJnQZ9jOEDoz36/GyeTTUMMMTV39EJzPJn4mlnavQ2HfI/p4uOSEwR8CTrmKmAKWkAdGkbgtf
by7MF6yhW3GH/tyqMbt75aFu1RQd14pWUKZ39DD6Qs8LyQrOT1gg/oXql1X/1WID0FIDWMNB32Un
7J/F8Dl20l/KJScgtCx2wSCkuJVijSM5sfyGx5q+uqJ9F5hADwsApTQS+HKLLRIV7QfbTwFCrO09
/WwfrJ6SEYLyN5pDG/+KbHV82FyihfPAIf5FnBTk+jGuyb77aOVAVtg/yWE2tSvgl37Blq73Z5bB
k/oYxHkhNQ6PnUkLQVWFTSbM0gx+EkYV8DNPOTNkehH64HW0WO9h3XMddQ80jsJOgQN7r9X6nIB5
DVuMjekFVxtTHw/8tylago+TcZCRRkXLpZGl45KPAEUSd3Io/1kr/DaKOVHlwYAbyuvwsFpIWUBx
CjeEwtgm05wN+40Pr6CohNUcthnpx0OqxDoaqrP0+xqLOECdDG48PMqrtejcTVmmbbqGh5BVLs7T
87h0pOxN1w41NaAfMrH3USM6CVfAn/EUXPRcgq1+eVgzstEoMW+xS4s4CxZGxJYQVFekaniMx64x
uw1ULBrZm7UOoTeH4ei/LGulzCsOSTdCj59e51VWU0OWq13eUIb2obGRiSCKmRMc+67B7Wk/nPWY
tnOygYTF7RCsNob1YiDNR/L9KCoR+ypDe20bETZe6wFghh+OiG2uf2TvUniYs6Y/Ef7TLAgGyKsj
RPRFDLXJ+HiV1WCUDZuqrXUri4GTluzfSF+vb9/8dSIjt1z6gR9tDfgkEbHU2uBwS2gEa1Dy4nZD
h1C5bSJIhpjnWlCQtXQvhNU/Q3xva8LhLepDmNnWknccqOjw+Iu5bqiFKuS5siB8qLF/gO97q3WX
nkptNLXXX59ApHzZmvuM3D+DQVdOkHfvp3gMRLAPmlDoGSK90SMrnWwI3gE2vkQZWVhSpwdqZHm1
gs6zKqWbFMVT08/EmurJq3JXNTVID3IvPC7cwf6/HhJh+Meg/OlZso+SDj23J3pInbzID75BVeWS
MtfyoHdRpRbUTUzpqHCshvDVogZbg6IB+ucLCFSF2mWFKHIUicIPtC6Tx13Bx+WQf6EPXiEags61
x+EohHskShO9AERkBN/zwswhFN1V9aAFiwWGJm0SlK/C34Fm5rYml6aRFXOkeyJVL+D6BvHcn1Ja
RNDZ8ZIzL3pOoHluz25FlJc+juO+Cgl4n452T9CVnnnZx9OWin5Q2Ct5kAFUwYlo0fu2I78vqtC5
KIvWFQByzV27T1nH2n+mgTk3G0PqF+CaibrOgbpC/KL+63UL2Qpr64WmggsaLxp6vm0Lu5gwn0IK
JUNcBxQG9BIm3indaXuLMRF4CAwN214dhNb2hANXoFQ0Wl0SR7ZwFQmcYgMhYI9G0dqJzVgVYrAX
xZTE6LE6jVP0G7K/BWkYyHtOiUKT6azZjzF0lIVKUXawAtXINm8kDI8cKU65ViTd5Zrr2ykbIghH
dAChV9FbFCig7MEFbygxDLvXxLvJb+McJQ44rjSWNDp6zeLdSqKDUrSmJtG4+omBkh0KxSPVF6wM
NQCbm4vZs0BmWF1FTckSJf1pLvqTQXP3QkNPl6+3j/BknFmk7t25QcUfSqSHckjZNJI3+1YcZdDl
F1of4X+PrSdmosL7kzxzi4xX0mR04NMkTx3apni3c2WGTmUEd7b70TT8hFxu+dOJrlCIS+xc3NiJ
sg9Xck40bmFBiywas8weScPba2t8j2E/jbbJcYgBvayfhBupFbh1WpzjhZ//do0WeaWUuyDZ5IYZ
OBCh/enDxNSUT4A9EMZL8KYxSEzUi+/Pht4bkdpvo7zE+r1V14ikdvBfSkcN3Dc83szpHCSEe0lv
yIAxVwlkwxUt7CeoIjQMEkMBsj73LCDO8UaMzPH5jFLUKKiSJINP4SElMyP1SciOTZia6dE2kfjC
SQtoLet3qqEv4IAWQJQEQnNgrE8zhIO4o2Ai2XViaZVv/LAbObLsoHtckm+XXFm9rNUJEhsH9rKB
vWxyLlyF0OAkngxjZRvg0f5MPSknlAOO+mqfxdLEU8cV8Quihum03aaepHVpxnItQeRZrLNBKTX6
ygT8Nh/LJ2/s1/RjAbxHlHNaodJawFVtfx2zkn9SCadq+89+2RuC6Ptgry5gvR2TOjbAc67rhrlQ
bTb2yGhvWQk2FKR1lz1W1/LdnmgLOQHiipBt33/NU7YdQrJy12GP9wfFjgtoSxz6wIyFvcfeeDyB
8exuhe0CgSqTrj4ofnsYYjzk3r9kvWVOpPSAVIShC1lY8gp1vbMZ+vHWhOZIhi02Z7HE5+u3e1Ww
8SKqQCDRpei0kGUfTvt7AN8tcXd1q2tplhWD7WmMNSeBf5ydDXXSZx5QZCLmEXptvWAIZbxKQ5WF
6VxtBEMWn2h66y+guQpFLM6b6gH75xqvx+wklfWhuHr3QZjaH6pGEMimz5UAL08IAmYyX892YAgD
zRz6vzr3Bw7VrmfpmegMAVtu53TjGwmVnNDHFrNkldlJFoISv6VF3Iqq0/KUJ5ekHCCKHKfCO48I
xA0VjuGYJcbIR2LQrF1kh6HGl4UKTjWHQHjp+wuA7U+6UZPQTpEeyE20hlhfdnEiB8CSV7qjsFu7
8olCsJLTzJsaPjOnN0Qz64husaO8akQhZ4SQYqZ4tZzcqGUok1Nvhcfw+vzYS33n0gOd7xvOZNRK
jUWCYHT26jSWRkP8yxTmj1scjF3JTAskuSf/zE9R4k15MSjBZjFphjXo3tGt8c7ra8teGMuxS0ZB
GJ1veMTZ9wXDVRNagDYY+/TMgWMmT6M5MGr8TJmxuvznmTPGtFzoZzGjaKLOvgIUwsLoQuX/1z4A
N72hwKZ5Zey24Qwk6QNjHrwV1uQAgZdsZa+PyO6rWmQWp3Xw1exeJ90joFJXJeMTqXhDOnIG+K29
rfMPrp5p+ivruOQ0NwbgHD5w1Do+ltsNjpEbTxc+LH3tTmExOBZjukndYK6y3XzJ4XK2f7cj8NCg
tALNT0yXhTH/CdexNgpkSnIVz5KkbvFPay1hescW1dgeezVN0Q+mTuj93hYfAfmtfzK/icYkvyYR
gq8lloyrZV16IFTbtOex5IOGPsVt7IJmwGvha+M9IHie7V5xDZtZW2nZQb8tQO2bkeGDgi6bBnE7
ugoLjmfsKkuDtHG7xTbEV5Uv7Xk5tlWOTUkmdb7W1pTodAQgH2Iw7CFlFpbEr7/qlX3kWwilu37H
VrwriTiAOXnaqkEsTmjQJSKghwMolBxgKUsRpDedvMTkxbVsOKR9hS3KD0Pkzp7ukqL9PF5L8FJW
0v6dSrTXlrQ4ieuy503cnARch65uvcNkbZTW5KAvgYOEjRvuxqXj/PcUZLpVpnsVr9PA1CPf/gXN
sbySSVvnJFmVXhYBobHqRaz9kieGc2ocDQRNgNH7/i/x92QCQmmyrRGgFZbQPF00EroFcEyHPwyL
K/Q23C+4H/og99BTmoe7Ggqh15kn6OzZOAGT58ag4fkPdAZuTO0JRgOXZiKK58mgVw7X0gC832eC
RhSBhZdv62vS87m8MtegWeziRbBfFuFsPeSqQNr/Ecqk6Wojo+AOvv5rAzyqOI5JwL3cjyPDSSqf
70jewSTIYOA0IdIIMHoQsXoBCC5awYFo89ypLnWCViIXjyGRC9ePs79ebArSw36x4+oj0hUVsdXG
mtdyuc8RD6D+TRr3HfsRtk4GnrQflU1OQBOvDb+CmnTphF2TjDUG0EMkV8txpFvIYkI1+BDe/HtA
XpVWSmNoPLk9vlgfThLH5pVCz6y64bAobJcslKUEePCWohR4QzOY17VFi826OwiPdEwYQI0z5rRr
XDcf0F2+thPY2LWLg/ZRkEXXhAnLEe0vkHFpm8MLInagn5wyehU8Bp7+t9A/KYuZKG3WrFtaipyJ
eiDqRAoguyaffVpyZsgGh84x3GnI62/rmrXsl1BtSI3QvzNxjy+OysSQFPzIwQab4NSfevfoEzXm
n6G90KgWhu8ppNRt2Y0eMb8VOUPBMb5ianPoSxf2qbcW7RiHPfKLm37bELSiCZ3gRBpvLSTaIfSZ
K2Q5kwtqFp760y45AxhQfn56WUgdu9c4OcQKrgzUQB0F8ejyjJ08w6pXmnMdsPR31NcppGi9ZtJX
7Y+ZU5ofztfRy9NHhDMEVZ3O0fooJIYBWCu1QNI1keCnV77GTs7qIWs0Q6GmtUBqLKDCdXdKzFQe
ZUq7e7zPBcie6DMdXt8yG2qm6Yd1+OeU/V3QIw82uDwhHL29rWSVYqNnNDekMjuYHL4raJsImQBY
Pqhaa9C2pCBvB1lBQkn49xASJ8DWtNexVv8MZXxUUUPV2U4Zdzy87u3UocGMUILijd49jrmbSUU3
HB1W1sxmRuCZ8RoZXYFqVT+y5fjPv/C63lSgiDYrsjkAeh8oBxiLsODiLH43nSsp7GlMVwnZ9nq2
spESTPNuikwMjVFR3Jhq9TZodicajo1Us2tWu9h80SfEwYTS8Se9OtgtJBsef6c5+qWzpvC8qeem
RKEn3iopnMhUF/Ff5e0QCsZxeq/JUPtb63tUP0LgIQA+zk5W8J4R9ujFlWPkkXrX/qjXjr/nc8OV
toR1U+oIBGRk8A7e9G0r9sSYOq+qenfvWOb8d0Be83Gl56+yzcqExWLWQ7vQ/zNuRIgM+UIWdr0f
A7xfWw15jMYxkqmz+DHo6rDE4iJ03gu2laJ8reEBZnZSuvwW6D5Bcv/Utd5Vkvr9ofoR73bW6ItJ
sCIjse3Vkk7Oneouzrtw/uIfX4PLEtrJBzJd4DVZGI3Di5C1qKLsUVqpe3OzQUKoK932Kh1nQNBm
ULIQdGjH4Eb0Rwnmp7KxqrPk3coRBb5P6/zCUhxmQzvntMQH5ZZtuTq0XSaG9bdMxUeRaNZgs8bD
abmmAw/OYFNnfgO4ciUezcdtaWOiAVbR3HMk1QVzxOai7cZVunoSqbQvuq5uf7FlMjKf4N0Ij7t6
mmnhBwrMHZRLOyklH2Hfg4Ket3ZR6marxW7+mW2TTr/Z0SHEh2yuxN2Ofb1calXkvaOr3qvmjhdj
S8n6KRN3p9Zy8pHZUHq6SaKQ1ghseQe4V3W6sD0Q5OEsuMtrQ1y9ijWyLdtE5rRiE6tjf342Rp83
umTIdgcuYuRzL79ahi/mG8jhTBLxLlsdeZkDPueQaeI+IVPWx5Iebo2PAMRAmBO6OAOTPnKH0wso
yyGgnBxhCTp+rS6fFZnNTASJ3Q99sT/xn/NNvjLt9IITklnTIydC2osy1jHSDR+1DSmjyGn2A/JB
c70t7l6Ux4fB+PuWRBwSSkD4sh4wTQTr3H3ThmSoFn5Z6qV2diwTU7Qs5Qc4g6CUo7Zg1lOlFGJS
oEV3IK1vBDttf4OIj9T9/ALuoBXF+gg/naaiZm5NZd63MzvoLt3EChYPA66xcZFMA/J5vhI3SEOx
znkBiPBepe/71jJLa+qovL8vEEFBeMRGHcUN3tLX/mDSMWjymShwlCnif2QaOUsbCBNTVZtlPIU6
niolxxINWsjfxYEKzmNlEn6NjYTduV5d7+DNs1T08IvOUB3rkxkzc5sngKmBOA8PEqJZqp4TS+Zd
va9cyefYCxJu6VfI5l+BbcTn/WI1zmOCAkoPDp0GbAqWmpFw0fLi0TAuo669N6KhsvHZ+dQmxcV3
EvVSFCgKucE3zRqW+UYePA01xTgESksi1rs5cCjNNkcQLPTIjTF8yulzVFQBAJuY/IDMS6XexTsc
n6gdl8g9ph8Sdp03m4dKzPb8J1SZ4KN4kgSsTVrk/LL9pdTYxJOxOG6AtRJ0CCCp7aP/ShOHAzYQ
71tdXuVHt4nAKGXqq5+2WsDJnsnD3Ss8CWyoV3lKOitPtckfqf57CSqUdHZ7mLvjCt6vqf0LXVRM
tG5VNv14MygBhSe5YFXkwmZ4An3Nc4jQx7aM84SQpBsT9Z2O+XIpD7+X0rGkjlZH34AiwmDxQ0f6
w50b+VljH5EJJa8Rmc+NJ5Adt0Ti0mXqQe1AYQBr9DsKOKs4tpsU01D2gL0IIRBV0wuii1vzwcjP
InCY+QjGVHKOedApV/OhhlW1PwseAASJxbrfCXtHXJiGEDtmFbglL7bLFzUhQJKM+OU0h2xae/UI
SagUm+PXqHz8aNLrdJYO3STf7htH0xDIN7VL2MOkZLqQzItRc70+17xAyp66nsL6Xrv9P3rArAnq
QSyHns4lBerIlklnDDy2xUKeKGE+FQI5fmQ7FgggLRC4JaCifFdrnha9fcBE3LOCvxrrBVLGK1wr
SlDPVk3uAG/NSw8abEevz8v84xRyNSNU0lfT3bUdnNQNSx6fGlzHi3ajGpYSks1Pbkxl0sOaBk6b
0m2yMKnks922KicKkjcE6nv3V4sSH4SsANQVYGZZEs14r0hXo+MMG8FG7+x7dBRWbc4kTmuczJZz
8H8d/uagQBbbD/AXm7+I1Bk/Qxr3y+Wcho6B2gLgW6ko3UWHcZCdjALFve9ZLpvRANQ9reEoV6+r
VyVjepDj2itaUVNYkHtQlVuxIN7gNrdOvrguIescv9C36+SmZ0EKXNL/LlUmDOXHX43J8EmJ83ib
LavXXaSPTnmJJotiz2Ov5qlgijtKQYG3xdEym8ZG3KPRCR640A8hKaovFYAzROo+mr0p5kQ8ZhGR
NVwzSJBAYrXpk/l2bJC+7/XH76tuRA5DuydzhoDFblZOIukGR5TpRK8xbg/TrVkXVAX5VYM9irrN
WY27NFhxKzcGxLAc+EcnD2sG6onBIL0g11X1jtgcDs78E+F0GK6jzigBAmRR+BZmobofhcPrO0Wl
TgOW20rMkVhNdyYN7qUekce6S5bZfzGsN8sOV0z1BxC66PjFPvsi4nl55P5/c/0a//SWLK4ShUNX
AteqMbGOGYAkgbvMq1xoSFV8N6oX/+I1lb9lUNGpZYiGn9POYnXbqkw+n/RH6Hi8/BK/PgSkpZ8T
rWQiWZV/edLprOlh8pr718LxtZrf6aqU/TpJrJ1rPdaVY2uMn3dBpJH5sbLpnjCdPIb7XPchW0pA
vebSLXAY5ZEjA3Zx2Vk0uc1GzAP+WSv1QTGpPhh7vl/Og0buPjXkPdQjAgoYs2hZzWNBBz0RBEWx
XigEjdhwNSjhhMGx4XvW6DwyvcFR4KosL/sI28OZdupRuPP1Jdys/bu2mR9Y48lLDkpRK58zXHPd
D91XqQHp3CriGX6AgiqnmrKqx715Yh7R3slXvSKCk4BappgKvYT/sLdKQQtElrpUWxTl92tX48ti
Er/e1t/CF/oXmBOj6s6qr2w0qv6OUBvOWq2PLobnL++H5Ov4M7eR7G/CxBZr48gPArHvpnBVwfx7
2X6hRmDHSgRbx2h9T2fAzQLcxGw+2/X3nZECISv6TDT109ukqbYsb3Htnt5COO8jS+qhvqSI29S6
lw+haBZPjngW32btxc8VVkqPADYVh2Y0UWFejonuwCjI1dfBHk3RemvT8H/aLimljJgs9EM4CHur
hputymnIE2svTdJMVmsWJfBd+1MiUuzZTxRpF7h+eyXgeiuREKKI7NyTyF0rrsG+7bM+63m86scw
boXKvwmQh7Raf5aT8XJ09Ao3GKQlsd5IjNcip9xk+Qi46nHHtnMhev55LbxHs1JZ7H6iVvAe7wnH
dc0jqdNzWq6HB77fjrBMmWBde6Edu7tu38niuZwSikJIR1KQru628mhl8lDKdLyk0eT8mzpPxGXu
6ndou+0x3Tq+wIn5rH0Gz2tKpR8ZS2QSjYGIyRyMhyjadLCSOm9zNUTgf4XbkzzjqZA6oVU9Rgr9
HU5ed0clSaVQTRgGX8xMszsWBFqDNvTrVv6V+ZyJReUU32/PY5o/bVpAXqE5R+hQfSbq+glLl4fy
IvX84b3lkwze4M/ycu45EOsTvPVcjdbeITHi2rgcy7HgIN4xVyTpEhuYtrxBF6CqLfNmIOe2wRdH
gX6v+BXrfTgJqJHsJt8iZJruzVBPpQATQt6t7pds8vgI6NR8ZcF8rqTDeUcItAKZZrhbdAhF0PIf
RoMoP5kNWQg4lHJ9rhntb0Z3Bpg9izRGNgKZGlYbcgrmbtItnVS9kw2psWRbKyk33knUac1mCUco
MtTLvRFlh8n/HYf5OMxRP6FMnUf1AVO1Zb3Mfe195lsN0RFBHxSnCHd67RGL7BXSr0JPPooOBSEf
OmUrl5zzgHq3mpjFSjQynsv/LL+IETRJvuIueG9W030UejqOvvRXd0SKJuIIL8W8ZCYtMMNXe9KZ
GgHprEuipe6+c6VYbh5hPWEIfuYNmVNUFvowSiYvdVT3MNs9GAyQ6ZnQm3+OHVExgbmWJPQJqIFR
JeF9dMzsHfCDco1lx28i8vc9iNjTsC59rVnDLLAnuaHLXkddyHKS69snHfZyTxyapn5q0+alo1Ui
W7/0v1ArbIZGp24F8v01Eg3mVs/WALnoCz0YLGxTxGSq2gIEB/+G0+IRdeAa5era+9RODdepmcTy
RoGrITikq/BmhJyO5q/3N4k/0LcdGdlAOdNxWbuGOAiu9KnW/BTyWqSLjhQ/2ISjgVAoRXVA+mtv
KgUI4eXfOGBjzpQ81DQ5ExSKU/srhgsJdbNMrkF1FMxMLKWMBuVTAQ4s28M3Elbro4XuHlJb4Tb3
LrjkjmiKD0WuIogKAoxUi9LK+jaxqC+3Goyp1eiizxnRPVVqKCt7c2B3AR0TUU6KzkvS2hCUEUQS
KH1PdGC3tbdOrKSNvKxxCo/9lGxmKHTLLsga7IrVi0vd7423erk9qM59TWMP8fr/hXb4D/fdIO2N
i5148YpgYd0wu4qFpFLCnbsZoGfr5na8DAxyLY0vaYyWo1p9NQ2NVVWt0Cq/Id6qVV8I1Cw+f70t
FpRxmWDkwRW4vYAeN2K5nbq7e9d5rOgs8lza7z1UidHwCzluSQXZiSK2heBdfyvpMbRv04UgC9Ji
hGUi5+jqbzXwY/VnFmmEw0wUb9Ey8ONWaUKwBzSkVtiZAcFYZoYccMTCTQBwrXmD526SnbKkvg+J
g0FJ+mNjZp1EJ6t2x5ZbyTgg/JV5KD9Qom/3OGLtU7TuCIlV72qfxqgHbjojNqfEQuaj8G9E635R
ZuLVldB9bMP87Gv7KzpZBpfiM8PyZOT5QClfjyMRAOC5cU5bgPq+Zt9faQYoO/dtkFLlsMLPdhfy
fVtmzJIDAmh1n4KwswANre4mRtKCcyofnaMnMn/FqbpOzfLv+wUe/qg19UUODrVrwRlTqLuMOQIp
opOejTldWh5gFZcMp70WKFihH0X8VDEPBi+iw/AjKaakEh3mgKmotxaq3THQ/aWaRn5wbg+IBnpr
uK/N+uMir90Hp9ntdwJrkQePcejMLms9efNYXufI+eyIlrh0aLETFDuqDZjNgdXmZ7cTpVWErlZ0
3vgcFo4UeEL2EWlH4neu4WuLxiPuTqnydhAPpXKih9uv+NjNIe4v/vuBWKc0QmY8nzot/G+14wuw
Apm3Skk7W8ZRLWKl548/dvSaPy7CF6v2GVYT4vXzhOAWEtSkVjzD6Faulk9gbXyS6xD1e0auQEtR
jWxjBpqbzTQ20QCeg25kNW++X6yremvR3mnNbTN4RDrwn7HYFiqzyfVyPNFlv8GyY5mLfr00kvGA
EtSe0ELesP5kn4vx1sXcXyJyBJ2xtr0uYRRtL8pSxO3qXu9HQn1eIsMNGNab4dMqoYhjYfnVprws
ZXaUQhywyUdgafT24jOX0uNFI1rqY/zu8KXxPBwu72ISfRlamx1tpPiGQW4X4Q8c25U3TCsLTRx9
KWZNtfh/knOThywdttZG2g3Uc7OHiS9rRqtSkvJBzLTpLqB8W28+A16jkJzOI28nL+iQxSyHEJv9
KjcVsbaUPTUAJ7kGLShUVMj3XwvtnIFN01IJrmwDuh4nlGPMkE/65X/O8YfG2CU/mgaqzmvt8i6m
Qhamd/lriT195vzxl+v0d6goVpUTHoZofFQDl+lwgHpLBwM5U/O0qV/K6Og1wRCVRUEWIw7XiSco
uU1NosmwpaiHJRftIAY/UGTJk/m54A1gdF3BmruvFjbt6ofNWjozOZlvvrer/JNt4y/2q7qznaPG
FK87Q9w1/YlZbuOPqt4HgUEm8W0LhOMnVk38qcij59F0dwGISxMf7IBFP2Vm989eaf6g4WlnB1z6
IFFylO+yp0ym+UCX6DJCQMcYCSSqc+x0G/I6HGXIMvCtuN7tDxd2TyM5Zjl41XXXEHeDVKbG1rKY
qYR9Dc7tlcBOcJ8cTcHJ/ISEQsfEczF4mK6ytYSTYs/3Gk6SIKcGwCqay37Cn3sQryIAny0x9Exh
W/YERSSqAt4J2lzMHEzQkzPSn1hLqD6TXcrND21KBd7ZIlsqaj53LZs1ZbjB4PVOKVPDfia0TqiJ
MoBO011jyPEj0v3n1kHcITj6F5+NycuqjkzSxevcUBPDapwuMJ0dsnnIF+6HqoL67RAJNFdWftSj
R1n0agfVZb0kLzYq0oRdosYYB2CAYDX8IVf+pf9Uzv3/IPR3G53P39b8DI66bjeZddymkXwiRZVG
dvl183O3v1GNjL06GAaTqSX2TMeeXr1Xs6q1F3l8X9Zb8xqO7jw8slCS7a9VxNx9wVTSfq5QBgOO
GAbwtFBcOs79D5cM6pdMuu05V920AVJHhb0LXUcPlQvgOx4/e4C0+lQAK6doRgr0bqYxgpw1g9BC
Kt94cpCaIiHk7zh0UOupKseUuAN7czIPwWzNU3EWCUW4cYzvpKxfx1JsNQfSEOdX0RQ18RRlc/oL
//ZUwfXipoeZysKN2vbyUjVxR/7QeqXzMC/tboezMQdBOuSs5n5Trounr/naeWqTNy7DIHa3dh6o
Flf2QIv8iGHcjV/9yuCKtbMoljjgJzOyzVygGGufrZuts81wCEi2BOXPv703TZVxfeSm9MeX1EMn
K33oxyQpzgZgHRPWKGnTlMY57U80CZdxPTLI8eFlCtjGxjfWJaO07+nxIzJJgpobXQYiN2fOCbMJ
fzsImP6185M+BuiXjT3BvsVqlWtTUtGJJ0Da6eBFs8rNSz/CZGGp1vBU4QsgxTRZH5pE2PawSoQw
wu5jtTrG8Do9PenMGHWP/MumXmkKGML2DCEYs2w3rqOo5nC3u0eBf8QiBxh8PrX1mRk4EOWI8Lvp
qvUzwU12wLCGW6wZ9eGnf9TZ0AA40jB4ULJ25Xd9rLTsp2k1cHDjrdC3sywK1nZwkN5XUZFdRCPA
xJjvVEadnccYK+pa5dMSCTbuZq9pkJM6mL5DBHd/D+PF/ZCwiB/RD+e4lxlzxs4dJQuJ1HVUDjhK
JgY6mHne/8UfqIE7ubHUOqNOuxH0c9t7Eh3+xrlI2CYJGm7GJBJuhd4GvCZB+Jlz2ebSCQuTExaj
N+W2yGNJqBIoMOWkYHiRZc4OboJyCWQLnMb6q8a9hLfGCE+0qrA4QpsiA1ZwCvp0Gp6YWDObIBN8
SUz+TOPw9+PHBKYN+DrBg+OA4g6uN5VVAAXD5J8yjY4awMYtyf34NXcuTfGtvN+B83/fPOHN5ncb
/HP61oIL2WjPp6v2wwy24bB15BhYectHrMFNUrokjuX/4fHqLEVREN+4yY4l6RRjsYaOP5OAH2B8
5xcWfmpY2Iwdlxczf0qCE9P6QHhOL5nxC9AFDlYRu12RRUoIGycceMT0laqM4Wux8OnyPvhz+mvv
m77LdWDweQWikke1iwAY9KLPAvHHfxsIE8YslNNMPcwKcjHTB28fpZemH3td6c1zEKnVKEs9llI0
NSh7XAQYh1eOMqlyZK/MZ7RJPUOaog5LuhvNRRDFhT1EgprfSUyTbFWsyWnCLl14wHJPkwr+bb9u
7+WbfL7pD+njQ+BG/3V3wR8iVljbELlvWv9sm1sV42ZTYPeqG4hf9aX4O9AEafg9fS6WoDksAG8z
KiwdMljHZoSght2pLdnILjwH/bw9MRw4/MbZf89wzkymGgDIOOyirvVpPGWXMW0SpC0zNDGMwv30
bXmS/IscsCkwTsJ777uaJxVDv/JHX7mOSiNZpfTgKuoRA7xc+07nf1vyZTY6xT5MjtKpiYkQpuwn
rHZcY3Dwc7BAnoKkP5BaYS+QhHOjgl40kIgQnvVGZIkCXkeynaSNCmUZAMsrYlmfrYTQagapB/cO
DQGHe8rxMTzTKYYk5glFcOSlQkKmVqCW5QSqdPFbYl087ZJIoXtjtPD0m66QezaP32QjEdhd/5HZ
5QNXqo66PbcRg1EHnPEdQ0jIyfhCPVlhMFRH0AVRvU/uu9F8IhIUKixSs6LjbIV/e3waJe/OKxMD
bwgjul5tKxiem61nMDai/bgR9oBPyoDD+rT3jEQhIPaEMx359RWYlcEzagV7TltDJQ+3mTCQKbf1
8/LJK83WBQxhfP66Epo/5wLQjK4k0LL1M/2mZ5KhKGSdPc6XM4dd3DAG7bUFBlynPEkQN5HY2rM/
C6yyet9CoV/qMaorLgiZ1x1tJoqednMN7uHkG+NzgP83tknX26WJ2dMX3qd5E9l3FfBLKCoVzpez
xyiz5pD5I8uz2flKQ+lOlBmjfJdY1xuYdaip3211R1rNWpBKVb58Jzb5I+ILjkG8bmPy1vvKaV52
RG/zhG+M3hcKjWxsFsLmfHYcgPQ2S1fUZ5FaSKhZcDRjhhphSvKwYCjJvauIHGxI0IzcxVxG9dZF
ixM7joNxEF7FkgVaAbSNaTdq1NUaXQcbeMdK1qaPFuRnO+REKoCGUn197A5rsf3nj+wci82TKsR5
yvn3kUTanV9hFI5TOu0Fgm3WyniT81W5cInRaIbmMX8RHoG0aXcYs4ONCAs1oMEcs67h+5CXSvlq
Izmi+c0gANri6k9dtEtvenPQvZrTS2/s2ab/H6QBft1Edjs1qQSA3Kuk8Et7p7MZOW8f6WgeXxQI
vp7cOoBwsPni6sjaEQ1PeIQ7yTLQfmQChAfrUjaM4Fn/wUkjaqg22y6FZ8VOH6TiTLO5O/WJePKx
xeKXL5m9d3GBCNyB3rf1aGJIMu7kNJmJ0ta2emnMqB5hSA/zp8y74bd4zy1ebJ2+vYnmUZkZtClX
9HUmpWZoNipOEPpIg22r3X3k3ct81tO+yR8Urp9eauoeQGwPAXezI6dipWAmytSsS/sIZxe7y4YI
J4uO0GjFGB/iYEYs8U/KfDw2MbFUuObvnjOe/AFUfQaJD+1i3V/Q5Burh5OzXiV9OTaWWOK4eAvf
pIabp1yLuW/uqQ==
`protect end_protected
