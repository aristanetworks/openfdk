--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
d+S1s8f9inRrM3bl8u256+DwB23L5ZloRnF4nzhhPIrARKLe2IuyxuqVwssmqL/QdjXW+eu1DuFn
h4u7xf1mm+ZpYW/DYuPhwcWnRvJ9hXZPcMXhBlTxn+OYsa6MiswA/voQYR5eANU8W7Sio/gSn3wN
eEupdtafs3nUbiJeyOZd3QY2se5BWJiH0FrayaPANjVmA2S6ajlQroqJnGa+0lIXIcOF1p/89Arz
3h7wPWQ1HJzzt90ujszFRsvGa3xMv7PIGtvdxC6IrVycKEE+opNQvyM6FHKr7a0zssyLah2WYVku
U9yyCL7rmF43LH/dX+dWnb8f4uZBsF5WaY6h6Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="hR8dFK1RUKOPUV88AXBru2lcBCeFOgZvty7Lll+c4QE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
jIztBXkWDdEDMZwWeOO6Bd7PvioozZiH0m2CdymPIQ0B65iWVzrh1ChaYVjkmUcmoxlQv6EuTExK
/DPT48EbIKoIW4A0aEFrBuwMk5Xc8YV6upHaMRUG2dlkc7HGsK2hJa1rYBJO96BRx0no9X1etu4F
k0SYj8r0nnHDtFKhB5+zSAzpwenm+tG+lVsVxjqwbfS643sLrvCdU9+3mlZC46uIoY0j5Ca628pr
UD88sm+QDf4KBddrJPpJ7e92lfKiswzaLsa3PgaYjolQcdCqTTJYbjIpNSBnD93aoIR5wEea4jE7
dq6qhlu9s21qLwo7OpuRAcKVJZpqcjDa4+aJ1A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="0Z35Ghr9wPu5+i6G0pr2tAR4gDe+MbLDx6rnUIkCRuI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8880)
`protect data_block
c6vxjFncpan8W3d9mG1fm9j5BvH3bQfjGg+zL7T9tOS7f7Z2WKK5be0icr68Qt+Q64PfPMDY2edB
mBSZC6KAPYCuY6iKC47982WSyOwXtc/R3Bx5g0J8picZ0P0+e1WM1UJnhkrgKvBNar8eA53/PSHM
WxY289DMdQiHsQrITmmkUYMMRs8AHv49bJeLkrSwHGymcI98HrrynmbXwmzAt1aepbqKnFeuTnNr
u55YQw72Ya+SZ3DnD6Rgoqrd1ZwEmejxI7Wm2lbf/RJj4rCWO9JpodLhSra1i/LbAGmuKrxE6chI
syvatnr0lNTQH232480vTsad5XpycQ64UPShv3xIgfsvbIsGRmdbw8yUtwXt7ClZ9qJAc//ABzG/
MARy4h20SJOc5A0Carwdp6FgWM6JlLIHFRZvX/fsK1vumCIoZq2RV8OOXmKwXx7W3SYV2Oqux8T2
rpiaxnY0+YE3fEPKTAZH+xMhdZSfBzi84POovy53Q8bodXW2PfpRnbaesDD3CleedBlu9m4hbSb3
8ti8aJFVEeCe9EIoQzdoj8dMfdEyQCjbNmfmEkwQcvbHG3ioDvNAXUzYeiZyh6yqLQORlEguZfxW
KVEcIvoX4MNpMl+wHaFLeEP+8qXQ8JCAKm4pICREMYgjZKHxTanooZz/dFIhhngO0xI49SePP9RP
rD3KV9zmq1K0O7REPh2fqk4OXtEU0nlUmvRQqycLM9Fc98wt1/Qld8f724orUWGHoTTiTl/26fw2
AsYgPIBAUHgQMBALjeK+2WYweGBcnjoZP9VmZGkIydt0KGRxQbbdQVpK4LH4MWAsDhe9q5rEslNe
V/4BFswiq9xbdTiDIHAssOekOOzkVKH3IkB2kSmkeJoQAhFoPmsS1XkK3qCQ3lJDDvutAv2MdN0a
3/asy2hhEw1wKjPlfiwFhomfB4SOeEBM55riSXY8bBGrwTK/gAKxRtilVevW0gTNdlh9UEfe0XDJ
CTGKd3/lG5YM/ewjJJUgmbmS03QbfyaKQF74XQWUTZhcYZZeFBHQzbXV8Y5UaNZs+Ihl19iV1tNc
yZIUWJcowx6wF+09qyAPmJauJXsDuY6jIBwPAyg/yB2RW08glLJ3ww5yKysUiMe4OyFXVS13bnAP
v4P8pg7QnpUGD3zQSL+h7K0QzRBBsQUtKiIo4Sigj+opKH3WhKonprZVQKlGejN7jpKuoqZyLf4X
68lMtS9U7TXnVxpjGgRqpP7HTYWc2T3CRPWDR393OaHyYCiTQevDezNrPpjX+LQgoK9Nu42P06MF
B5xLLneGkEUyCjispt8MpubNcgHz9THMyWQo7A4vKqjTebGyHRrDQFEviYNLKiwO7JqGLZidSkUt
lEfNIb/XB76+/yQtOQtPEnt4BEpOH9Jdemygvs4ze1rXXFVh6XsRzxNoO3TU5v60XVOs/PIcsCYI
5rgIy4NLCq5SRJ9uRVDOIMyRIGLTKIfNl748v9z+F2ndLHYVWXJvDJ9Is4aONFQs1jKehtL/JWyq
3toRMN2ORCyYpDfNbHmuKuPjcfHA7DGHQBjUMHxyDxlHBOL2W+VJ4cn/4h6S0qebuTnNLl6mY3/K
exywp9gDC8jHt0uXCNq7qfVuePx0RXXMIWWbax3ioKkvgZzX+X21y8bApIC6gvYNDTLDL1JopjSc
GErMUNjNJ8WTXSspLDEZgWkF2keWNU+8wkvo4dwVM5MxxQTN/704eFQo1X57jPFcbSW9dzNk0hsy
XZnuf0buWZaeusmiLZhzXekuEokMDuawsMx5J+chPJHiLFQcc7ROGpJ0m6G4W4ZjbxT0tpcF2Dfz
gkbO1HRjKb2OEAR470RdI0iG5abuNCrFu/DDuB1Yot/S/Weoqm9DxfZ2vqVIT/zuwqlYx9iykisn
0MY9eJUYzcagZ3tFmWo5ZWBpIebXco+yj5y0eNZdJ6jB6z4tqok92NKgPlMeX1SsqVZQKiAHq6CW
5hDpqIJv8k1JpehLluulLEYlXn6w06W2HxJgGhy9syJ/Zf1tbbmRJ8OFkgLq2eRQCdJrqvhg7bjG
1njokHDm5Eh0M3KrotvTsBiKapFrg1egI1Th8TLYxXHQKXxoyhlsud2VkyLT9ulg4Am1HRfZZsVA
J7jH6sGrQ6683SRVGfFNjBTzH0eKREF+yc586fPrTGLIzPGi/5INSE17i7Hbd3gX3u+GZ8752OnU
4ZeS/4Ac0nceuqKIwqTM2vemam39euCoKYJS6Bd3/InXyiEjMe9yX7WX76Rt8TUbyRe5g2gE+FC2
ozqtz/V+jfr6BgvwotzVYKxYoQJR0rYSh9h4sCVlMEcnKGq6xgQJsRNKFhQT6R/bwNUxFdwT2bK2
r58A3xKw6FWSSCZb7AzECqCmbTFa0cQSxvzkorjGbJjQsnkK5d3TXo1VREZIUJD1bGkJISZOy5cI
OhelZNDoTrPHeTqTgthWZWXkjQkOOpRa2piyDBSjxkPBrqZfg2YpwknVL2UusumV+K50st/RKx2f
SeeeGf8V5EqYwfeRIleQNAxKZCCRUNEi2HDJuyxkdV1XSfniiDTDGG19Ms8JNo2f2PTMxFhKKzbh
Nd2ypQN3VlMk0wZWf+pur+C18vPc1uBmq7nUg48g4sFYqO5CHbMwBGZADlzzWlCfY1lRO8CN6jwP
heZD18GWyt+ZDpB1qYb23UlneViuAIcAF5O4Jj+fDmClrnVVMWJk93x9JAXL6oWpd/9PQWzSsm6C
vb1WF/aq6+FeCkjGptS79g0qnmbA9jEHIlDQWdU5QIyLttgw1qEcWrwXLI+oINObbnqvF/BjtrgO
SWSRiU6X6d/G/p4/wvL6iiBvf9rsyw8/wvll2kC2jq9eiWqiU8f+I0Ej/5PeBWR5HL81AtQgMgVK
+BiClxa5Tr4r/Y3Yr+JO0PkY8Es49PIKsYth2a4d2iZ5zsTnDw5RUD6+uS0btEcqNx+jnOJF7PaD
nTDgIce/p4f394Vy40ob8parLcRV4CCykYwrbx7+QLwkKXb+Wv+PP0Omj1+Jp4IHf+wpN5NHAdOm
QBj/0xOoXFF45kBHN0UDYzCHSJI00J5hHyeA3KNObbZwdbxqA9wE2rgZGDpTFUf9zeaTkGlNsLt4
Q8EUT5C6KmgWhLDEFsvFN6IXu1Nuhn5eXwsgoAC7uZaHEUHYW0D9eKXilO6zubwMV/4G6jRHOI8H
G8foWlvMuAqEHE8yDTl3MJckAhN3DUDGzWe0BKSLLvBcK9Z3Q/OQWYl2i4qi75pF+2cOJ3VaRKB8
dER4jxuPHnwjrNOejfOXahZrUwW89fv6N8Y5/OkCb/4es8xZuBqMtLkXJYTtBnxr+ZW3V7oPyK/A
VL5AqFCWiO375zeRgJNzWgQ+5+SdBPqnJrmQr1AS3ne/HKCTwAYuVD3IqkR+Jl15PjtEJ5M8icmI
ccVL5nxjJ96eOPL69QUQcqZeyFg4vItUeodElBTIzSmzSsTBZwHIEiKRR5if72cd1wRxKZUHdwqj
GVcwbqcCMoFDyRQPwsfz1E9v2N3bOY+8qNrXB2J5aya1+8NZnR11b/fd8a0pii0/XP1tmitc2Bxs
NczgjgfhRncR4ZyT2/4uZmecvjwGIKeXNNJqF7ZjX4x+qpSOEben3Q2FwZ7/T4Vco3a1w9CWeK6I
XCryx/Sy9Ffku4CGEK+OkvHF1sl89sbhOkbM6AgCXEKFbsB22vMFA9N2ofM9SMVLeeUUYZXHeIsT
S2U9vahMbRx4smJ9ssy3mJW5x2Nt2MYlaZw/6Ytg4+Wu+ed9f1YYhGL/s1GQZ4rSWXGqaC85BucS
PEYWD/xsz/MD0sUGWKUaXzg8RwlCvtMOaMsmfYI7Ou6TSDdgOOEV9neDftmoV/aSdRvkrwBirJSy
kFMQRxYp2kD8S2aDV7UXOX23z7an9+LSPtxEMQ72rrRej5z0aCvFqyyWwETD8stvQ3L+WGc126Q9
lYx2KqWMhFQ/bQ7JS/Jp9APZymxTDEbRmhjh/0Xa8M838S7KqyZZAO2zGjHvA0QWbDxxAi1BGfxc
hauypL1uTAp0VUwe/QMhc/vjvv1epIcZF7s7O2ufuBdhGDD8mIOugq3bjElZvaTR4Ooms/jRBawB
MqWgfCwuBbf/Nwf5b89cFG0YFIzW0zyjWKujUQ3dbDac07/VRYOqxd5F7HYH4X/YN5vjqCQhs6dJ
nfD2qG0BudjgPKR5d4ut21pVw5+mfKtTgES+E8GIkQY/wilzCSHnKfuLNYAttBc9QOe7R9IaEY94
2Q+8xn87+fSRibV0neuzfpNiFOrxHbJNtrFWMlen0MXbD/9MSXityLY+KNuihfdf1k3iX1HbtMY2
Y3J22ph2U3k7UFN8U8wMWs9LNGdla4f8GegmAL11t/5etpPPHRNphA0OirOEEJ3KuAW6sIgfm3qN
K1JEqy7BKNdiA//egOuRCl4c1VGy7/GY00E9A41EenajC6K+02T7Y3/6KFsm6Y1XHCUn6/dG7DOF
ycxRZI6t7aIP0m8FNLfYPaEgBgNbDwQWlKJAwr9ZsX0VSVGNyKBxT/BS8fch+ir90xB1+smQRTef
b4CGaaklsWHNrc+MM+vRi2D2jHpBvlHWbPcC+E70/cbzoRE86/85z1uR3O9HNjF/uf9txVYnzRxc
AtdV9J1fMqhhpBKtH+em1iJvJFiLOvSaKlelp09SAZyEZUnLyJUvgj6FpyKs4gEeE0KaaXFGzKNX
teH//CTB7D+PkhaeHkZpuBwHjTJf23VyedHSIE5BRvkfvX78R0I7yKAdNQ4a/1H0gmpYkh6LCfQD
E6AYYZGZ/Z6se59cxUPL0LI+XSZMj/KgXBa1wFB06HYWm+dxgJzPafnRYjIijN27RAUqdnTb3jkn
mq3ApP4v3zzbA9mOET01cW6FUH6ueIGXIgl/E5T4AwuFkP1VvYsKOWelwKDBxVOtdbGQ13E8Cj/h
uC9p5do05GFRpBoX3Hp5z1ZQGJTN3ZjPSf5bCfQPxd9lNSq0+r+7PJB6w8eYvzWTI+Z430e3lZjq
JeDRi2+8fjUQFzu+qfKvp8FfLPYm1MAAd/DZsDWbGNfmblKQnJKwuex/KBGEkQ1ZFwrXrrOX4qoc
/snP+fpa1+v2sPH/qFG4U3n8y8bpCTHwTtAMw4Tisu440jvEVgERUZ1EVfJz3tvu6j8RhT+Zg70E
dLNLWV9/Nmtie5QUgsFjbJvXIqO3jSNtsws/I1qnUWbeNhmmbuypFKnMvCGiNTWg/6vntrYefDM6
nJ2WNZu6SkXvSEEgDrQ08aMkYfhvLmo4exBz50kIYVmLIIhpFBju6I9X2is4hE8rsXnv1bQbs/xl
JRN8n8YuRuq3pK2lFlrlsA1MivtK1A8m6H7qbrMohCSSZZpffRFCO28o79xufgJzPz9q21++Z8Gb
vBbtYNlgHsHlL/Y3lDQBbVNfApXecNw/ARMJl8M9p4EoNLwyqeLZVay+fpB1a4hErh13rKCGoeYy
KAzBr2Bo/D3q7TSXneK0VTwts4oNVF2yOS14zqHK18gaDtkJB06av0JJDXIL0FWkFnRweERCpgMn
eNbA3bGW8N0xOHeZxnhV3n75Zm+AyZDW/4U8meZuOeufm2IyEhqdQ1dqcehdDvGB7dpA+9cTXjX/
QtHl2SC8MbyjzruIEYNk7y8Z3+fA20Nh8hYJHe4ge8IA8cSi/QSvQqfdww83KxGmVbbiVAElvkrj
AzGN5a0D6NTOjUA6RQjQNxxoKOYwYdRFv4LNK3QF+LMOEbuYyKkmEshELGQ8SndRyCHLJkbrjaI7
u3JwqPyxRlfqj/tpnro1OGPJEapIw1NJBfw5mqiFf3whr75L4GmmQpbg7Mm6RMwV/BKHLYkkeqdn
0ju/YsTM8FrXlz9xV3umUxSN94flKRkM10oZ6zYTiFZbr0Nnr1a49NAz8Yn9qPkAoqjQsfdbQ4iZ
L2GjAmAVu1bKuXQYpqal9nutrWlZLuGSQx1CFumblhPxFB80TRES9HfmMU7DoPdM1ZdrWnVVfuOp
hhXFtJi+w9EfNUO8OQoPtJNSttNII95BIaozBEUUcu7GNPoVAWMMNoHHx6Ohtc0X6w3KOkV9wrCM
iQ4dGWJ4rtZacuXdNI8+LvjKNCB30rrTN6CTr+fnPuvUPIbw7HBpWiEynMGHiCQcBc1QnBCUz6Ao
y61CtrmsnlpO4RZCmbU7SqNelqv3fRcFMxz8unBKAUbLzTwjL0Bxo7wIh1EIzyrjNl7mb+3T2UuE
cxGp8pOkSlSb5BJ4qdpej9IEtezCV9MVV71r5BhXCyB6cjwqz/budkf8xnX5eeQZsTY4pJgomOuG
qXNa/3bZDewt8lh8jnSaFzzAvCC0xxDSSkzQAuJKXbwSNsCxxGjlnSTRaO3TX2zt3gerAv5sEqFY
WPbT0tqwAIwKipgGXC42E94xBoEB+5ers6RJCWMGtnamHV9Bu3t3LycUfOp0qdK6YZQv9TUqfRuh
qTD93DH2tWjJwu3QtQ4X2ej00Gfyxkli1lLKixV2lsNd761Na+YwxtCffSPgfwDKyXL2eQib1xdC
yjxeP1BE4rSbd7181m4U0yJ5lnBbX28eMZoW7TwDAV+mJxVqVmmfdOWSO2jcdAbqQS2Cbi98Y/nv
5v7Y8tICLj/oLyMWl8oXZPZMvY7qShWlAv2V/83rzdxX7R1fuPThnRZu8V+x2SIgJrqLbTKciY8i
7ifNu2QBs66h0ic8BRI2LnUbLCdqGtVgJwLmg9wNYg4D2e0nODtLAxBVp/BGriRtZ2/tIcDhHVf5
KKS1bIoGoZkzODf+Lf/whK4WCzJOfA7vZqWQ/8pGu8OBnTzeZQpeNWA3+UxwRU8vz7Ko4Q6nqO7E
jdyfz0uOe6PWkabl/aLE9mc3EpX6s6lqfGDdTerjwdEpLKyE2RzUrU7zHfgaxBweUG9EV7iGc8D5
hgrcynXR53iaWTd22A020WkPHuWtTGmJObE+uYU8tRZTU2KUIg2JxyC4V/3RuSIzDw6fmLh0Me1m
h5+XjjtaJiTxboBMsH7vHTKw8ZI9jFwK7hXHlt4q8yyB0hKoHncsnuNBbPWdchGN2vC+R5oY3+Th
zm2M0kC/H4F8I/XnSNgkQcM5YADlAJjA/rM56qwgJBEXWkWHJd89xipmfW79f2el5amuTpAQHn+G
LrClRizxvYBDxKrrXbv3YNfjH9fJAT/qidv/6W6uTltnPY3VjydJ2cF0hJZLIVsqDpXZFio5svBT
wJLg4i4jNAF9cvaSx2VmN+kAXKiJKqlFsEd9zEomHDdzvCTX2ocfIbf1WJs4m6HkF3rWfkN/Tpg8
2FBHx4Hsky1U6Wzh36xwjVz3Now3vLkQ5TkUnwlS6eJlJT8z5JY0q4QgLrMMZxJz1rV8/OuEPhvE
HI0qiu2BnVzPLb9skNV9J7vvCpsbe2zSu2NnVFD29H/dBuYcwQU/VUrJdERbgHtUfCPeNhWdKnlZ
XJRHi40ByxHi3McPRD8nxv6PIyacZKlfr0+9EdZ2yLuFaF09Mne1IQ6NIuH8VaonGgE3dPBx9OsS
ujoQlg/xtA2oDq68BMX1PwmGdkFUrvErGUE3JPlsYH9awWVSyKBOVOp6ni07zxbasgIZOaJRUw88
+E53LZlxWXL9w2RjP9YDDxN681EnG5r/TuYzzib2Ujz3KGzCA9ZQRPRpkdlY2PJE6b+pPxFOvwrt
ZXTsZnlWUwccqjk/QFMbMZpQOj3Bbm0bET1Knhr4kmwinejSbvOm6997qOdzwdpY/KvqJeX5+tt4
1mDIDTFL9dzIkkP6gVAAdnP9YKAo+oW8hS1NJaXppmLk+fnumhU6xykb/DFfI92nVt8jOz/LevTq
1SBPwhUUs8++JdFdL2LOS3Vy4aqQsRXP3uiGU8954I55epI1OfSfIflpIYvI9cZGB8H47DeOEK7o
Hsff4WUJfDL6Tm7YZJ6HatFFmOeTfd3YttI/L7riUv4Akwoj7HTZ2HROGbEPQzmpYt9VMAbMTej6
77QJ4k7ZEIIDpDAV/PgqUyUfRoA8LVwGgZszIpX4OCA8Kmve3+SiYVJ4cuQn5K6gnsMpz0tkwWhx
00DoF73PBeC8+5alk5eG5TT++p32gotKW5cytlguDyh6K3eI7yEhNQHIKPJvz+r9OCUgCF3AUyMd
du26+vQsu27kPnjr8l0ytOKbhVQmPaGf4JpaF4ji0rolLaCGhg7Ff/4r+6J/rb1MAl8IHXZu+/oY
rfr4ody6k4UfL26tW14eAq7uQTCR1+/fAbyOJ3iHljMrQJdT85aBxZ5WNqxtB2N89ImjYCfpGeFV
IVTHc34CV3U5j39nQDE3PMGLSfkH3ZyrKfrAvBx6p3qXvCFloDBb8ezurqafVgYMdTHHV+5PyKWs
NasIdulnYtitqrjgS0JJ0cejbgRXbLhMOdZUbFS6cgrZXG3Sq86wji5Jk5VTf5K1YofurVdrKtHB
HKjpNO+rxHlICj1rQsKcHNHAvU5GsJhehW+hbZgSgAtolj2WGtyhL3SxUNNM96PMWrPvUvAipPDg
Yx/kvqMzM1LGlksysu1zhJ18aYXHJdO2IGWrWa+yG06P42EGd9tUk8E9vHi17o0VYP4yhu+95ecE
vApKHQ1UIKA/PHNrvXOUkQMF9rSdHD2hY/pC2tIm7H4xlG5zmakDXciLQoTuCI4XMadNcmop6BSK
7fwI1zN+u3OYBl8DyNizWrNisBCUof9KpRCsCITq+a4SOpN04PUjaRCNT74MWjI8o1e/Jlc3nuAA
/gBUCTk+zWHb4KWgnSIkd0IULY3FAY7pbZwP2kMvz/viczep5epyceUn4MLy0ALxEB1+VwDOrwBA
mGYjytRqD0byINGb8ovGKOpf2Hv6gzfP+LoTuAXYpTRyRJbW3ugOGjMxbFK+Utsz6f7Z6rVq3v+J
FSOVP31SZvz539706CxR9ZUcmGNtWA7uZtSWxIzoBd3MnTXU/WmXSpfQZWiKjQE7PaMONN7zZhKF
3yGwi+nzJxv9PWThX46z/x5iE9gvxsJ81DLREiKD0FidFXO8T0czT7pxFMCsJ76sXhSF+g7wjWKj
G/os5Dini5nCcltCKrWrT5PJhyJN3AgIhKdtpRLOV7nLwo77sjgk2dTHP3b3RL+CX9avRPTl3Vsx
cmgOkJ0hA0e6I6+MNGuHDyjtCK32cz84JZOYe4hLzftCfn8BAIwJhZyzmN6ncPW3hO6zOJnK09jO
EI9qp80PdBKoKcfCtVxYgn+LL2g1WugPsCEFwQtmqq9zWAZNJLs8zA/0zHWaCGbOa0FF8jMYxQGS
VGBg7RyXeiNqgNO7A8V890KL7R0p/NHa6MEbjBu9stEegetf3RtRcXdNQOeeVBnP3iAcvPKN64Z9
sZj8KyJwZP9W39FvRO7JLIna7xtZrq9QWmxXJYUYaxHnNfGIvJPvcKP71OAqu9xPyMA94yLv1eO0
4csWvMG8vtpiFmZsC+UfSNvZ49Mz//N6PyfjvRUh3kmy1IoFDIu0sjnWdhcTTaFpdIGW0YsINHpr
N26rK+4ex6boZP5n6I/f2b2dB8qg/Ud7fqV35r3GH5PhYxN8/0dd5ijD8Zu+b+N9Ykce11SwyAm1
ju5HR93B3RdQqjz0EdlCU17bUgfGKnM2Z6gxTMAZT0AkMGaQt4o1x715F9OkpAmQjmzvJpSvvgVP
FYveA1oxa6BUExKTfhdikbl0cilNotkXNVHEB1fCJUuQ/by0TchvUOYi8HzyfcyiFfmnlSpmAu/w
49jYhcqic4kyNNS8X9/txP0V9A00sjxVnAEEEPvy2EIavk0p1ltUQ+/ba2fC/HivLZErD5Y7D4Gu
pYnTVKPkH27qHJ2bg1swFjEgMzoeM1LkwT/ggZ9BPBbPkwVbdxsBmxdk4Jfq5WhsgQRk+cGACWnJ
vRzT/Ti3JN0Q65FHVL8f2lNCZYQBHfzrOH/ggJfsFSTDHQDZyWsKv4GpbbVXvFF22sBrMjr6DzFG
oaktVLs2Q73gofeHAzjsqT541KpR2QW/DMYagAIPrD7fZOUBXKd97UE0PH5auFWD55FZbdpOC85X
re9jNuS1yB4PLLWfd7jCTO0YnVIhG2bcKib5kr3r4tH6mdx8n4FKNrOXaBm3BNL8mljn2YPZhFGz
YgIIQxKZydmHekFRdMNOPVZb/IBcLKADes3Ct0xeulArtk4/wlvCoSkVOAkuMVdAiZX9rf9UBJ0N
jAFyXgnt6xwdG02GBMB65mRSGloLaejYuZHJrPsoT3gCNksCVpcPhGWJ+CevzGpXgBi7jeOH7dpO
G2z4vBEfUQQcOPTlir/UGBmiG7+ybT5OYA63uF305rPNamhD4TeVG7U7Hw7op7U9z3oEkhZz9XR3
yyahcEEmgdp62BHPJacr1zPUXfUJ25u6OqYQ0x5qXDXG2n9XvKY0YJkh51/dcXi9Jz/R+s/WPBqL
gtY2zs+BEeU0uSW9xC8zjjZ9BIIZrWXVSKq4dhU/5+A3T4hE/qEhJH4QdXbijpQUXOMUpzf4jFkP
YcglRD2Z3FdmodPyfJqGGKu/L0EeJiF6LywRO/W8PDigwaxBgBxP5qq72+qHRD0fveFcgF1dW6NC
3J+STIWkbKJSzIRn/ZSlYYI6EH2HH9y2KJjpviiczS3liSFCUfkefyuA6rj9SiBZox1F4I3dLBci
pc2Hy9fi9W54KNHxTEq2FOwPnS41d9t58OP0u260zh8WaNybiffr1KnsgXwm8GAmp+AocZaohCDP
/eOtSOKeIZetzFzqEB//TqCW91gg6qSqwwWFVyt0RN/2zc25xj/FdT+pyZdF/JbU9w8D2x4T+B8p
jrBD6hkv4KEkpjNguPb27GhD76wxR3S/Mh3bHQbGcZ4EN1DA0t+kB2OTGXuJen1K3lVw4jMkFv2r
BJ7Nlvcv0jGoCPhl7K0kEg84WPUfjUZk1lKMDZcWMkKjRp3K0f98z4rli0HRNiJLDwyfqyprUsP7
Qm0TyrKli1lLxyZNlfnM4WD8PQdDiMB7p4kf1ySS9mAeqqaEaTY75ujZlej32CYuvuRI0lcG6F4h
47+nQ1SNSXUyikpgOQSGguF/l/lZhBDbq+erpvzCL1c8YVeJfIV9sw3ZEZhQlgbaiQ1V7xxheWuy
sG2RDzadcqFPiZd1a4k37id42YF/iWmwU5ovK+wa42ZIghbf5DqUu0BCWWyvH1BmaK+amFSUNWCf
56snvwxZGloHLXIPI5lIwhZdAXX4KmOs8Qtr6luswSXirzA+CgqnP0kvQDUOtD3BlMq6g759l3V9
664KiU2F+HoIA5J90lY5yTkdhfevLtp8c4iz1QDlKgqKP+ycKgS2rI1sogVNTmHkCfjHVxtRmeMf
YZz0/s86e3ikIr03P/1xy6tXhsM14qdNATyFiXMXdHwBsxGW05lJgzvfIhlWpgYrAoxRdUh7qppw
vvG2uKVqhB2yGSwG4xbR0ho1LsipZ8Lu/u0JLFwhEZ+IStQ1wI0MiWHxxof8EhyZU0b3HGrbB8Z0
e7npTmjJgLqfwF8NcXvyAf4wvgl4ul1Qu+DPdraNx+B7Xw1dRtFALV9uPy2RLHxdBYbJC+8I88AO
SlUBm8J7O0LUUV6+VpigFC+sHz7IkgXv1GOQy44CBOaI1nTAhJiYF39rB9RSbxmal1D4WaRFq2dA
f2qebgs95GULdnE4fkN6PxAmUz8S+hI3tlAW6QF4FbbX9vkNqPv0xgMrbvQNXFstR3mdWfznwus6
8VFbxJrXyKG87EcDvsdI1MnscJdv0Kql7ul01ZyK5Cz64k4J75mp+oWRgwekK3SWVyT2Utk39Qww
mphh4eQNj6ShaYnyF7T1qWJs9j8W86xG2S4/EwNjQ1MYFPVsV2WvAbcRkzW6
`protect end_protected
