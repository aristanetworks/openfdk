--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
HYMf52/f/uCefq0hUAs+KPzTtZuEaCVLB381MwOTeh6gXxPoqyhOuKGES8OhvGCbSdP/CQJtorP+
1fFCZDKPtKVGY/eq78F1OX3aEFVVgiyIQIN3h/dO0H5LEckSrNuIrSmuy0JPdGRhrF56RED2zxFe
/IX3tVvluWL7sASCvh+M+cOrDKXZDZPdlZccZoJZrLSntBTsczNF16p/nqORrPjAqyVnIRP2etbk
INiUjnmbhcKRwG3Sdh9nxurnKvMnV/HvixfmLPXEx28tAl7d0xwWfWgi+V9BYQm3cRTc8s/t8rCB
akCFgI9jDJHRERFT72bvZyJjGvpNf0UD0USMlg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="UJfYzbelfdL7NBj1J6H+NB2FFk7ggZWPJJV931e4JWk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
l9mcJlJRSeLdNNnMSgj0Nwzk74XvWvsRzWIjoeOAa65ZvWnOPu5lPlh0XZ3K/Zi+GGHh/06pYqYm
ec+OSQdntEYe15pAMRVCDBpFIyBL+RcMe+JB5ZemfRCg+TC/7u75ye1Ma+ODmqIUDYLi4Ue3KIA0
N/aYryAT6U0Iy/iImsY2Yz1lcB7XUAI7WjD9DZCvq8BurXZ5gNnNmC5+VdV0A8+rCrbkAYOn19BF
woFL2XuaUSJBKHnZ9iCAPKcboPryzt1yqvbiKSh/iei9mxjbnUxKaViwkgQqtZHq0PhrT+/uXj3g
afdKtMHOh+IJLswzncsCUNgBWzG142ZMPgPLTw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="01oFODi7GOrgn3wu/lzXwXF64AnK50E/eYz+OnFELiA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5472)
`protect data_block
1N5No+88K/xNvN8E2V1++kLcpn0TeqHW8aozcw7syh9mFsEmTZWfLuYbCv1WzulNmgZ2r2c7RcUB
gvJ2sT0VlfoJYveW48ex1+cU/6ScdUjm7Qa2pH+6ehukX+Lp9o4CM1wJG9s5UaU7hM6mvRP72SLy
TnjdaHaR+hSb0Ti2iWzRwF3LOZ0ppmRyM+rAQaQwl/KNBAYjrpuIVa+J4e/LvK5DU0qsyp/vD+6J
SckzZhF8m4EJLsVVa/UGOk3rvK9pnZSOWUmQOlAYGlgOt1Jf3rzuO5xralpDC7EimiASI13hTnNI
Flioceaoncx+QoM8H0T9aRfPwxi6n4fEPq7ikpj2BEHyzsfvI6nkdQPD3MHMwUK1NbKUcxGyLS2B
c2ZfDPM/oRDpteQ8chaTJCGPTTFAY7vcBRU0ok6wTNHIq0hISdAilWIwYUxhGe2nkw5YO/6Ytwnl
29csNTAVfe6oDmlEQpw30XSPcMnKKP/Y60UFmN90rXt9aUpjlefAXxdiViY0S5vcZKxYxEAetksg
hCa+e+razENxxCVOs8EnsaddZEELTm+KsSRTdmiOYcEY/vtYDuHDL/qWs6G1jWB+5xwybgj0TkKo
4Hibffvat+uDUevuM1Yyw3Gv1V0zBUuRR212EfNGPOBvE+QF0n05sWe8YWKbRjg5yNjZtqImjBZz
dUaIZKqaAXwskMONiFd5eVJ6rIugQ3vt9/8apcGhG8h2rBbi4MT4/AulGl3dXSqXGbCsLLcgg2Qt
KPmmtnr9PiDe1n9bRkyczBGvq/nxRldx5rl1P3dMAyzUGCKE2fEN4eCPt9x6jQINBoJC8Od1Eehu
+0hSE1TctIOGPL6fn5PhNVtydZLuwQMt5oEcN0WmxQrS8uwW967kWSKQ5dPVEo1xmpEPuNvSViH1
7Lqe3t4ihv2UaMnmSQkow9vx/n118R7DSA1MipqUHwLJZjX0NkaWNktdG43OqPcI26m2EauVby2G
DnAfccRs0kGCW1H3fLHlmO0lhCFeelHGO5YGuEqrD7AvoIqzaoM8QFEf4AvGwiSYx2Rv9ig0yqky
n0Jq8Sr7wH/nWJNzWdr/ijYA3Q8xj50lDM45MeCxeXS+MoakU4nIDnAQt6Y1G24c4ATE16CGT0Q8
7wKZtW8g96oyogqjYnaY1VFujdfW9U6M1LpiZcNyj51TmeBugnTSeb0RZ1L7DjGdr8UUQCtX0nw2
9PtNLuc2w5ZlIqpny5Vnd/6zHiiwPRmiKRjkzWb+SQvhqxJzVAf7BVFPZ/LMBU/hPGKzMdEfqPAv
Mfrg4SVSjO8syzbE5ImAvPiTzH2cMFDDraTQdZhM9xIcC/WmbbqqIRqfF93WOnTvtDn9YFyVx7Ss
NY5pZrJ5yeur5H1YuCfYPTNr7omBhi7eY8uNgEB2G51BH+JgEpyN37Ly7J33hByP8HRcHTV7udPt
zKWOqQOGDt8S891jGEQXRjEA5fDT5EcCCR27MyDkLMqKSHrW36oAys2fXzNdStA51UbXAyWPrfNA
z8QlfTmDwN9TlpBCgETLIGIOzKEIpR8MI3fpTztR4Pq2D0cfraJA/8iMaSGWZc9xcZ9B7v8W1SaF
D82aF4RHF5SrRrWeMhaJOQIRpYN97M5EUAZUbZKKgh6B4wrRE6I+sH3waBe3nXPDB66IGae5xdEU
rxLd0x9/yGaxrqmh1bp/uPWKy2Btrx1sQ4j55OFEZhIYLef4xgBatDHooI2mitPYQ6mRDSO9ZsRY
34wui/FXZUmCMm1kKyIIqTiSvp9hH68URYs+FIs1cZfYw5b0jTmRt5KzNLQvZndFT233ctP/C5/N
jDsd8aPy39Cjj79JB9aEQWdQ+ttTM0fNRVSqE4uFMpjZW0lBYfs7kLT9SfiW8I2ANoM6pCA3MEwo
ii1TDh477w+Zt4lYKj26SsOj+pRS8RZ1rzxKBddWtwj5G5Zy4zs1xUK3s+mMNuxO0ry9LMj6ZXz1
qFiB2naPbUk7O3uIhmNYilfKqiKu4ubCa0u5L1TPiPdJAEyZXLQ4gR1d4WcBUINWVghCK8NQNL/Q
Cs5EvrQ+TexS2m6eczck/qpzrJwFbDjOK0Dit7xA5yjGpd7vvuto6aP49DxCnhRgc3viG7lp3bs3
62t2zIiexo3MTZE/wF69H1G4WqmwHaL5Paf7nDRXe7d4SltM6z4iexz4icrMs+mlf98Q8wdaK9JH
uNP1DCThXpy8LcolpnZqOMyKj7EH3EanFRe8iBjlyOrjeOffdto9cRMWiAtxXBr+n3PhkkyByfGS
CA9WaJ+idsLbtOPDej/delxvK+yNb7VxFnUOTSmsXbhXfjJ4dK0y3abIDTp3aOheCH2OyCr/YlH5
VMrxUG3iqhBB4Oui2qly1sz8YULkauxWEPtjLdKNy1RvYRVQ3+kmivKv793ta+TPLwlqhXGJ1ywe
gyC7mPqqsKlZ4Ev6A4I1Y5lx2PvhjINi7k+4KLabpuE5fQNi9aoDPpAJK0J564dBffGuKGmFIsck
fQ6ccASjZSByOAPwvziOPas0OgVrN88AG/lpKVLaZEQmEncOGuuTstTxBm62CctHZD+0vAQfTcIQ
7oOFJM8sH14fVhvOG+PoZZV7RBUhNOI5YSPfVcUavN9MOs9yO2ikYAKEJjbtf08FoR3PWcXV7aV3
S0mvhmjzNCHwQoN00NHoL6WkG8KQ8H0xk3J7nZ99tb/8JDB6t6qwe8O10IL2ekhPaqZQshxp8EqL
KyORj1ckMU20ALki5eQckR7i+Q5bfCMQya7XfjFcbfK47gJiFDCdnN691nB37WT5GS8qL1TYCWwg
lnYsXNMwM35v+1qeX4VdgIZA10rjpLbJmctPBE+pQ9n3vi2uRHpqTDvDactRw02iYHpA3XGUNNFr
wPssGvFm2aqeoRhCSvM9afEOwK9NnxM9XRU6TII/A0qBJUgEAs9yo/Gb8sWoXezSrM8t0mrxY0oi
f72sD3DDkrhKfsfaaLgyqUARWOhXtKCldEh0lrbJDpW7Djqf3raCsGB+5Yd7JSgKbrYOEV0Qmoyu
QaPaLX+eQDvdlSH8G8viaEw8IutpBheG+X/swNCSncsGOIFPhai+QESRCw8s8ewvtPLZLJfx1U8e
gF0lEpQckOOcsCvWfiZjNyspYAczpV5W4eRuV6/fToPhQwuFKWK1letyrN4q7/9Gres1LXFZlagK
BxPP2V7Zc6YWTT+scb5Mj6B2emv32wu3g2jL9cJb1b1CG1DUjkgI337wSumm5CqH4wneu5vYaoVO
BakzWo3dTEh49SvlRIXG2oEyoAOOGEz+z6lZ+MSxbgMMNtngmekuO82jFeYfDA/2ZhscoyYGT9Xp
w20egs3pMZDnhAL3N5mSqd5JAem5WMxuJWQceTUe6VMG5BruJR9VdNPgZZMqWutmU4r1DhYL1cwE
+XKUNP9266gl4cwiULFjEbeAO4a04ZzmTUw0viXfi+SwkNDbtAetZ1Qgfl2VnN8YWy2qpCI3x6NK
J/PcOe/XKe79NTEEebEwzQhQS/erziZ85dokuwXs/2QTkrO0NkcbdP0wwKhDX45BZeLRidu/7KDd
RryFGRZwZ/2DXt6cgT0dhgroUD19IVA3BcT8k3L+J3ouZIeON9KSOrjyNacRIFbyp3p8uGi1o+/0
ir0w08cH/PoWuvVaJyepk/dBoSJeBfyFNK2p3cLEq5VgvDpo1g25UOg/O+3UJz3+qLqYI3vy60j1
OD1Y88Q7tpcoBXeR/lFLvtAzhyuOSzZForfoI4dviDB4OC+JdhAwEuFu/+OhwYSmrJcqqzTf8gJu
LnR+SkGqQcharLpJRYxrQvLyWD7a0E2mPMZDmchJF1yQXHNnZ3NQs9a1XG+LL7zvUTcywDbeo7Fj
EbEzfGWgWjQ9TaqtUMoJ0AS9MpVQwJGXLVQyhW15j1r9bySp9VNStVS3Uzhy//Nz4GJP5g0+7Poa
CpUHE0IcbayMV70KQMOOLcDgo+XYgzWrFHOPNY2oA/eahAsUQ5cVQN+2U8Tk33ew+cyrC3fbVdSv
5jPDe5wFEABj6qR15hgeSkqtmOlyHa/OTJ8zxGnTUK5n3VpfMGa7NVHms5vP2V/BjlaVnOYEp2RB
cR1cJEmtSXf8lYXrlmiawKoltJ/cP61KkC7r1DSVgUiYPhRiUCImb+uXBh3cTZa8xKnVSKywJnEx
2Jw/cSqBRTwCdYDXAnqI9smSbPXyD1noZTPiXwZhafHNKM4rQLmd4sXw/+4xn6xISk53IO5seS6V
Q+d9hVGtSEOY+qukhRFF6BpPQugH0v0TfZNIrf53aFGt/sVzFRIae4fuNY02kH+XB1IcdDZgL3WN
VMI57qCsJ4KSN3TBnSz1tLgZKREPYJN5vYDzNACAbzRdbcAneIIG8kBv1gFUDdT4hVJrj7QJPIzW
gdw5ZtRMn+jsLi3Mz5zxFJZ8wlXpdfja/moOHRHMV5AiI0ZazlKZbwoufWNbaIFiEUEK9X+Ao4fr
2qBnR0ZzEbYn59WD7bthxDaO2gjoI1NA8ZiUUpt3NX5eYQE7XttUU8zA9DAGYslg9aQ882EUelfF
CrjgKdimAfQkJwsbwsbuiah1OxZW7Qy7AypWAOr0FLnhmCm0EPzwTKRczEyIEMLsnQ5mXq7+kYuA
WEi50hBZKPVxLJyxNKqthmL6aAb69RWrQw7ZVeaOxGeOteCYkGjkKtkknOkOi+2vDMSuZk9Ju1pf
Rehf1Wnw/LljCJKpuPvLW68WAhrpzQWGMgfZcouth7WXOtmi0Qryy5svvSwquVxRu9DCSKrUaJAx
mEMShjGRPFbunQgr4ZPDcT//764zgiZZ0TncZvSwJ+vQV2xwYUnkbbeDP8B5p8KV5YzpXczK0Tkn
mHG9X4W5A5l+92RbbsMJ6XlLK4ZxYMsWxdy7/3FpfYqLPiPuepIe92RZzyt7jZ1gQ2aIW4HUrTRf
C4IVM+mXp/fEUk9/e1BMMPNWCPWMyNAUJ7Ru5Jrcx7F8+XAMbWiJK4pkkQowmID8GxHBKss/FEkf
atLa9XQTCwfrnuyy+d+CAW8t3fHWbicJQZgiYou1OWTWgDyW4GOuHhzaQMXntd+dE3DrwZoceaWR
WVCQ4OT7GmL0Nbv+qqffCuNu2AfgMoKDC56l2QyL3tQ1Ap3KtphdOhVCTzYoOFozctPfFbOZGCKn
5XXkybGe6aI/lbEbRBAysUsLuLBl49u0RtXbLBvZ54vQ+UsMJf7EdXGDJFoDNpN7QN0/hDdWWkpt
L95O4S8kQGdM3WCDu7mv1gSplLXbBmfKm8xdtSJ+cfeiM+5IG2r+oRPlWbeBDeak4NCriCX7B06f
3Nt3YtCzoHWnJVMqNLsw2F64fyY2oWvakv/6Kw8qNTTA3YiW8ypVv8VJ47/5FPyBHHAJuLv7lgxA
AlUIrWlFs1qODN1JOyV6iC4xoroqvtYUe1cVPnSHQDukrTYYWex4m9YtF98DWAKgVb8d0zLpeERN
rrdiFVlK8BJUOsE4S16snjPj7/13YOCh7JSgeh2RPviiaiIlZjzdPDEfY3mHZFpUXsQ5pFPgzovU
f2zWo1VvXSEpYTkOn7/U+iPIdra8lzlcnFyO6YFybQlpJgJJzTlxKqNmIepLAkjrH39KkPDNQCDV
8CDS6uTW/ShJZ5UGuKAXQ2wk43QOyUy/CC5lH7tM2I8v4cBaCGhMJ8EzOMgUVxSW5man3M+BJQ9J
WajDPnsRrZibGwK22Qhn8lE09Jn5EN4dpEASYEubw4G+4h6L/M6vsGOvVbRlW3mEwHh4tRNvcia2
xXrVxwyHmC5mjJL6tjhwwa9ZEqttjkb2yQdCBm26A7dy9bcFpC51ANXdVxx3QOvEpapANFTnlthG
o/HfP1S2Dra5WhnfjhK3SuG0Xl+x3+r/bBWscVaOZQyRWaxUFYvTO81rb0tjK1iQ+RtWwJ2uLLSC
HpPFIk6HCTV9jwyilcdldONryaH1+Yso9C2oNYOLs04XGJTJBXi9fNOBuZViodwDaBb35EBfarp7
Ul2IEmNqILFuflkfhOcJCcoutY8a6xOzD9pG3fUbibH6jHFzigDCqrHtHSp5dIjbGVKxyVF9MTR7
wEO4CQT99SqaiDOc1HJKScZqIq5Zp+MBz/Qe02FHsRolShewUssBNY5is2f9wV6sjng7+Acox6rc
5fR03Bvgge7kEQ7SGaldvMbxOpfEXte2bBs+VG9vOklW1bkvWx586cCmJj0/WWszrvIzpEnr9L7q
Ny/H0yFlbjFMrbCsE8W59JhEDB8PeRT92mxH+K2abicLW5wWV9Kp+lDiPkPLBVlbLp/nu8Di7Hzm
PcoGsaIBS0U/w1oVFGl9jdiQT32NHgE4VXauzeZqHdbcSwyX7JBEJ6hgBKWRRo3IIoqeQefX/VFg
VH1un2H3ZhvKadAOjhVEH5IB6TVjCGCh1/2AgDpvsrrquViDANZt3s3FfHnutQ5pz5T9YKt+9OeU
oUYZ40Pl27IumtvJ9zL93OMR2xvw2QTAqGhZX6eKBjUJkYioDyVbA00tmTpScoElhauZ7XlnEzqD
Y+yQ2UxPiI3xbrKAQ1N5gzKKPYLI0pJaunIylqMO9+ZNHSjcYmqDyZSGJOTNAmcL4kSiLM08RmOK
6JhEPLGZaERoL41apWesOG2NIXAcbF3smxNewXEH+UWrA5njsVvj4nFxuUZ/7pCUQIiz6nbVHu+L
SCfPt6MrcBrs/KrGn+ePu2N9kIj05lYjIm5BVVkL/+fYF7JzEJpnyuasYbd4tLLhyfUMtgaQ85Jy
8Atq8wp879URrBlA67Wex+QudUgpyrAKwzAeGC+FMTxl4QOnJShpERHeXXTVjIOYUpjzf//fMgUW
G4rzcUCtSTZTHX5fjloLV9lGA9tD6WSObSHcGQcpj08oxBHBZl6Vl1mmq/wMp4naOipAc9Xeyz/L
FNeuc8jJIWz7jUPYn7UnoTFX09CBieFqSavU6heyhCBj5RBQwpQjVnFzTHqjGAapwBCOaI/QzoYt
kfC/3+u5W6lPbG+UyTWKbdPWhPLYtOK8S70smKjqjfArKzuXDEXFBIn8j8PQTQi0a7oBOcXYdBlL
TQkoqeruNaAX2Van7ms7xIf4syAm4NKuHWtkW4jz8gh1ABtAmFxsEcVFxGTv9Qrtw6PPc0nNmRbp
lSQJPsPYmGDBM4hudrC6cbrsabzBGE4GjnbsfxkI7kCXvpIWCotZBNRpu5GE1BdUyj3NhhVI5SyJ
BdaE1ejf7Lx2jj+GxKhWryvhJym6Qcc5SVWGg5ado+8MdcFmtQuUoFFaN3T3gYfNtoSL4u6k81ZI
`protect end_protected
