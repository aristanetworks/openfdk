--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
iv3h9YnFO5+9zZ6Rksu89vWwfXZkBZeq6F7L3M8k/sV+5xBAVAD7Vo4wjGi4DCzmKshiBuAxYrJB
B13szknuHFHVI5zvMHpJnNZn121z8MK2zqeTuxlE586hMP0E7/IYbhZoy13lygqFhPqOf9OM4m1J
JoRQWfz3Q94dxi6+Kq89+Xy78IMM5NbwQ9r6LjlRXKmv/nqYoK5bIEykz4pXVHWjkfAldFK3p3Hn
NbiWardU+/FacVZT2SsqdWmkzc0Ncotr+nAWsNxZznhY/sROZSyNz4SyIplGRPhQs1oydAqP4mwU
XgTkfH/C1Xeum7S2xzFrvHcUMc8znl8xlMbw0w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="iIwxlqLQ8rgPsE7lUI1/Lz4pjyDsEEPHMtDT216ARd8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
N6FH58gEf7WJJjV31urDnbbJSylphyDBCD3DsV6W3YBtEorxSv6g7QBFkt61SDIlJMQGYfyu4peH
DgvqbycdV1fp+0P7HJMzHW0Qzw9SoRzn6ZCDlJCl+eA+S2dCU+pCbIH6xyRPa2uCC9TCPOKlPxPO
LR/Ee/lgcc9u4SPPf70wLPflAlHdw8CAxdoi3NXGXb43c9p4RvXYAOOBJkdQfqXdeiilOvNK2Hy5
LTPPhQNcpVij1iIGXcOEiWgcpspoOrmPNX9uRl1hJta+T8fb1sFbRwaWfykZfVy7iJIRXIfeukga
YNGLdfqy+iauZz3fknF9jqRqNSqZ0ORDJDqirg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="zf33bn9AMmayGqR3F5EtCzGi12szFYqEhsq5WnpYQyQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 29600)
`protect data_block
fGc74KmAoONiJYIeaM4zCoLXBksTF+6hcAOE3oKqJx7c7xvwOS1UqznnySTxMqxlzMGJQO/YdqhN
QHOk9M559JuXXk1q7EIKdM4bwoLax8WWG76vfkuf77dXX82I8+46JTHAnLDTInr2HeugQgM05Ci3
jMn6NZwYCVq5jdJLBry1qoGq7oZ48b+AzPixdENYwDQtuOzq2BZssl5I5DSoVo3XYqesme1tvH/D
O24LLK0q8iO7Mhsf4aNxTOwPyobaZ9yRxOOPXmfQQ6TDlHV9pXq4OD8MgSrss6jY0893CQywQr+6
Gaz1AB6i8Sf5nKqQ0KJ4ZqdHmfTFYW3WXgIQ2Pb6vGikY581Ufj2Sygds20cbpzI13q8ODRHfN/L
WbxAVD/n5lh0ojE0DFCfiaNIjitpKJbPjb69KM+Uk63x6xlBdnkl60C1nQk/DqT38T4WAZgrY+6W
FF8TnqWvhsDwuxmXGQ61ADyrr3tprTwspqmb3EMyNOfrsuFvYLmGM63kOIogu07FMK4C8qUZetgl
zfNOFuy7/+xtptzp3Zx6yZbSqR2kdD9SrWfAnG3yvSoXR3VU2+CGfSOjkqkSRGbbpwxqJ3JNqYw+
ig9ynWvtLOr6Dy7RwhNQmDaKNepE9qqpWO66gB9mHvXRTGfL8iJnFg26Uw8FepYaTeUkwITpORqb
e7LxUfrzLY0USQ+An7PzWy3x1+Aqx8rMWvDMik50wnI1ZG8KHDVFsVQbNHIgkfqoOiTcmYa+QrlA
iNW8NWQjTDGZxeKG5M/5U/Bxv2gIhQ2PdEvS+8FpMhF7VBq3PbyhNC139t08h7Zoq8bAsAT179pK
ounALVqgHqB36dGRFRmbj4/2yC9gsPSocNp8oaJCcM5VHIxqpQH/2+XYfVPkEDVIiiI29swAev8Q
EqpkYhcSvZ4k5gjx/gFGGy9TEUun2Ty56CJEHwNRS4OVYKy6ewLSn5Ymci+EUvr5vTu6b9v/wfY9
XV95C6yr+fot0WV+ICvPeSmOXp7/wU6LN+/wcU4TSL/QYDIaoHfNn/gYtpbwBZ1Hkz+YF5I5vyCb
4mhPa0Ot6aSeAKwU7OWOJwA/zWO9ERoLeRi+Af0GaDKV/fq7h3uUaxRRUh1AAAH/b1GaKOQEzDQq
OL2ko+tAFJ/N4/Cl8Ovo1Gnb25wBcZjYhFDIHxGY9IABYvK8ufiPbOnTvYkP3MEhdd6CeRdMQXOt
NFmd5eZjHqUBN9yZLS3hEv/NQULLVNuyroAxWcuMxmlQP49M23uRYMhitW6Fh7oT1CDsZXyW9RDv
zrOxc/kt3mbDhpD22EHYuK0m1yGuuu2BW3cUlewHsbx6VQIckpXC+fw6efD5Ydo43nnpuql/S73P
Jfp9RhZQu7uSZTOUjy8GGgbldTBU0vAS51EX0XcrDWLuizEGvNICJx1Pg7Ue1pkK4tDiH8HaBVds
KWVOhfTJB0p+9pUc0TyohTlnzJ6pJr+itXO6aCoptZ5r5uu54rOpdVE9Y+pr9F7FUan4BkkO+I0i
PoTmQIT6ec6l0TwSSm4th2myqk0VbeXl3x9S2hyOlYYwdWzUPt3cSJhl3d2e+rtnpTZ3LmPMfMI2
ocKd+sFbDwQN09jHVH3arlaPDk6kkM5lk0zUCVXr3UHHuM0XnpdwgJ7qAmkO4D+IschcBVqtS3gm
j6iJPIyvxNg3ktsB6JE6Ym47goE0ho8O1VKO/i+77z1QMdbHueqS0xjamRJoZatxxmWHahT6kPuV
1Re88JxAfQpBMGYudGRTkh6l0Ul3Ar5AmVSpIYlu6mDPRPMFnGTWiU3N861t+Zhp6D+z200drnqf
jqfjbaqesLnYt+vz6/B6aSDhVK2Vmi6BtIjwHDXxceKH7xEUm7MJRWuMEA213kjrnDkSwGYlcGQJ
p23FmLM6xzmJ7A1o0ECtLn3Z1NZbxpfXZ3dK1NDvXl6ZlJcOlTgosgpFz/IfzIdrDjtlCkTeltM+
dA9BucY0uCGqqlJqID4uwUk3GHrp2SioZPXMAp56sZRsGLIMH0OpgaHxWHUjSklNoMBLdpVeYGkL
LJNofud8YxAHO60a2b56aS1EZKEqadlvSx8bBPbUVMzXoWzOitGhGU2Rz/RTmt/VEesZCdkF5FLj
MA6mwUZT2w5WCMd1/MhHyrh0W3slX9b7PJxc2nn3ZnTmQoLF59TyenPy+R/XSHP8ikRe5qPM+8hE
JXhOZpX8CeEXLwVfoXLBtBwFB9lj4OQQvdt+9LcrAApIF5EPxQFLju1LYlWsPxuf90FQpvbID7I/
TxLj7dCK1m8a/FzPVQK9n1iVqYNPcfu5mwkfOM10WXm1kWkvRORYa8/RAQoVzz9tJwDuSRANkaRq
0TjRtDbOoz+heyPOl0JNPEtIV+MpNTp603aKGR+Pj9SKPziyTQV7e5PO7bFDbhWplYWEmafvpTxr
Nj/jjww9EwEAPwpJXPO6ZMDDbgLNkbS3sOC6c9fx5zTvjxX6bTBue+f+pSXtOJSAFPQGPNatJcKm
88nhmRO4Xxrc4IzVtsfxlv/q2upeK4vayH2QbvBh9+IczlytyBf7WPiKLhZbqYm8SUM/zvyL2xRI
dDA2YrNLZ2Z0KxVXoGd7UvmWp+rsstZMYeAECQKWdMldgJiLckZt2EZzYpRZ/Sh11F/geapb7sBP
FuD4an8bMeb1/tDSrxEgyjaBKd5Ts+FcG5qmb+3G98lc/IDlPA3O2UKZopIiNkLlLZqodWt3u5hG
d8CgZcijyKH5VnIjGIqD4M7OY6NoguWNh+L3uGwZ2AuQ3A/AqomieeqtxiVzHQ3S9B1vBov4tO5r
X8nrCBKBZUGg/PFW04T0wP8Lm5B1MVIq6blQO6kS/mnmJ6tJbjDyh4AXxNral4crUDHp3Jrma+Qc
yqtaGTnCpti2+FFQbGWtSNIoKhdTaFRfZ7J+Ghiv0mMgMgArYI1abPzm16uZdD1L8/AoGCeIJMqP
NBPcqEQ5YwyfqJ+Lb0mtkEcT7nFf+Jjo+Hozc2Vtl0vI5nCWf2s6WdfqebaH6EIL2uXp3LLMfJKc
J3MHfzzrR3XZa4V9aB+L2BUcYwntY1SSgcbTmOZlV+FRh1K54E44jnB/BPOfe+c5Q2n6Cx1rj2pG
+ZGgy05C0pPrPl7chJTu2JKwifUBAb6jk67cVvGRRkd5yHQ7H2v/SV+C/JU3zTBOTpZnno+biwMN
CyKbgZcFW0L6vef8Dsey8uWUmoGxh2aqQxV3H/p5dswVeZHixO2d/Ya+7K5yQ7FqASe9XdaJowOe
/7ufMz3ZvrdcCAaxBhYpX0+mGcKD/s7D3qLKEsOtgU0S9+D5hjMytCtVl2rvkmyt3GbraGnpmW8S
9R/4yQ//d1yZSboNcGBCnkTxm8L4IhfeIJ5utNnffbGOQcONcsxmv1Cbj8cxGsOrwM4TfpW1HtYM
3igqCKuftH5kYRfgBWC03FJ/ZYs7Ct7rLZKcTXy/wkjVwgEAnPHm2+OdBaX3tIGEUEWqY86h+GYM
fwWKp4Bez2RXuFPN/dey+XplYBIrI4PazX/uHlI+sZDZ6/TBhNInPRR+tE0gLBDzUqUSZDf+CGR3
eHOON0DTXGHh82kalvyCkajyTTFWr/Ujs+BVmLIP51DjXc8kdLfeGYj5gfEDuKEOMMMIcIiKBwgK
X+fR4LHo3zEJ7YCAGratJjwliMpv9Tp/lOkx5Cz1+SdQm51xiM3+PnF5o361ACXY4Vjvf8h9LkgP
dENcY6fTfsxM9n8e1Yan557MosA2LNrJvDort+nm5t9ynt/cUkOarD1D/Mox79Pf+jTJoPt/jPRw
8b/y5aiqVBo/6Q1I50Z7WLAM1UYkep2qobGzCly7nUaYvuRUGyIT/PRY4dlRKlnUxh/Xlk/DRTbj
wnF58YdoYi+S0DtCUHRZc+cjGZBaH916W6iYSnFe+Di55TDI+8963bL/FidOIyBaNGfS2YsX6sAv
Ryan3uGRG05qidqzf4rUJZehfQ8z2ieWf/9ELoio9+UE+rc4OdhzHzmOrBEu/lrfYc6uNb8bV8dP
aj9xfAD0PNjVn5H95ifNhP7gd/pj5S/KowSZn1cgjrZUE39A9s7ILsLhPMgHDu7RJucVgCbfN/Su
uYKCmGvLFBMMX4L42SL9N/N3CC9mrdrnDXz4fAfvzjqEuF/cDnNMIRCdMu10vgSpm7keCVWZVi6y
ZjHVqWJWey9jO4uJYNCQIk1MibORvWgc5UXZjI6jTG5xYXpTXQgrOnsoRFUK5S67lULIs8y9XgHl
o6Mr4+mmcc4q14hHWs2kCp4EeX/9qkcQUqBDwmDTUDwFKm74lZgHyBeeSbko16J1t77efJruL+2p
enWWsNrm2pmunOi+1oaq4KeA3T/1Gy6Ho5lsMZLFQNyAbOuMwrzoehYZRzS9sMOh2YspcOaEgKUI
JWfVZnlkiTu8qj9Hq1YUPnukPnfjs3RgsgwzJqT8Jn6MruNrlj/kH+3NQCL92CwoJMOmJfgDY6Ym
snvbl3OUAvto+a8kwc4TcCmYAVfTAeddrK9cdySb3zU7x7rZhngQAU+YBIaDHyFCPopOAgnbu5dv
IXACvFo4b/QtBuBWN3mZvCN+zfyR1kAuOH8x7GNMWrl1w8M/VqxHnSjZbEi1Q4tbLh7RpwVhaaBu
j/6kv/p+jHcJAegH2L6WYEoVhQyy22jZnyVQFwPZfLqh3tlViC85k9YehpAWB+bKKqBDn4cqicbS
dJMJXHK95dRwFWJGDjnsy7Guux2vBOKqmlJkF+Ut6GAuZsAuTjHbvHsSy7myrdRgczFy1R4SAbqJ
/yG++8RRRjxjnlzxvlD7IswSr6EwPiT/xvPIIvlAsxZnPcnANKhxpqD0tnWuugXlRrv5RIWabqHl
sNPodSZI3t38Keiw2F1wTM9ZGS/TkLgsIyrdr8vp9zxYdSZ22qE8vAvTgvSdwqktrgNf/rogJpFL
2s4mMDnNtmpM9GUoLEUcVxuoxqV/tt3vdagxly+FrpUi6NVPt5pn4ht3VOrD02UJViwkuUPXGN3Y
7HKofQGOC7AmOVXoYR74qzorXPB5PdWkdZdwV9n6vNwRNsemE68Yz29kIZSOVZS2eGWJv1BYzNPE
30XQNlHXUsUg1EW7yha3fJkd/68mqrADKMADDDTN7+UUqq5tGBpfS6TlH9U/7dthpaR44Ht8TjtL
0UU0No6fhoSD8u0aYKC/PIYNStgqK1Mk5/Gc2o2qlhfLNg1mxfXJNUKRKwGo1rtHkPdryEoFOTB/
iB9UgViAwyZFD2/UiRVcAG8eDkcnEbDSVhJhjjJkXYHng5v2h/uk/Gt7UaW4YrTEKBqnOKlmkNv+
M7zQketEgamwfzcyNx/LOxsNqCxs1t//rQxlw2uEv+V9ta5WHwxQ5q2MyPIChwfZooh09DNzr9by
G+zuFpCdmp4JtkTGK90PWxmc1nhQF6Z6Qtz++D5CLr2IHWTmOj2fIlNwpsLr1Zv3Lme9Tt8Qa3DZ
7HHsqmP0uKhmIK8/LEMVWZjyjmH20rMa+QDsF/lZx0nSAsL/GcflyR44fGgafPuUAuKaXYTccm50
FdvziT+K3F/TBEjWrAyAIRwgljQN3IOWhEd8Nvjr6Lr6eXKKyJs2mU5pZ2YjWxhXOT2kI4KyCdLv
cbDGb26GB2qTooqVk5e+NqMWKknyWHNcZO3hK0+/AqVq6KRjLlD+bja4tTu1z4GQ/zb0VUzKvzaj
7CdMRV0E1aFz+/rpsBKpZq2wg6R/V4Y1ArsQMK5ThOCxIKtIvaiV2BIspxtV2McQt8ZJ01B2yWZu
/XXd/npHx96p7ubatIzLMRwMqQ4UVVdcN2Rz7TXn1pyru6RXW3aI33gQl5pAnrumLpg7XEEnN8v5
Eatfip5e3wdmG8vI/JbKlTLM7kUglytdHlSYSclcWtUKLYVtOmxf/hhmY0wymsu8TCeqNdSX0At+
9kbRQftRlBlT55CXUyRNKxNmHn58mjvAIYxl2Vu2/JMdR93BeAfTwUDvU62ja0dZSyde5KCkJLy4
LNcj5utUac7SPWdnpQRWrjDpqJcbWZc+hjP3L5b7SVYX/Clv7yb2toZlUBaHGumFR+2ijnvzKg0r
P+cXgR8WVG+kUCWBsVVmbRoYHNwNOItw1oeR/lZ2V6H/JMlu7XBd6xb52hE2ZDaf5aFm3xvy9K7L
n3j/HsGegGNaxDPxQWOKRamP9/GHmsTcV6A2JBaByNicKvVuRvO0YbsXYvZbCCHlxD0aB9uwQaIj
thv119PTNKapuMnBV1PJtUlBq7It7DPzd4UQtYoVo7gZvVY1FDgcxCSq9KTMmhgFr+yE0DzDUqiK
5zmCbwY3cjUT5MQ2LaoNeLtyR9dg7wcs8TQCdwpyWcrHPC2kBqtqOzwa7/SjTTng0A6qiq3sBSKy
JRW5jNI+I9N6qwsnGaUiv+KnGu/JyK1FZvJ3C5jwgnltjRJYoCb1VGV2BkzO9JQvofGMfzVnmxs5
fMQdZrRigNNHt6FDgVmy8i/txBNSQ51tPlIkGGf0BMufwZux5jDtJV+qyhLEkbZjXcsUBMllwW5P
eoLbgo3LhZptAloFyRaiWYmBL89bHu2rtTjeDhgoxkOBA6QSEMxbukdy4fPx2lZDHeElodX7WAB3
e+hzF4Y9L+SI8xz9gqQXuumSs019Ad8s24Bq5khd3hYchKBSoR3ZyodUO0h7Eh/tnSKLRQaUptSg
kTviacVU0N9XfQm4LqQk8uD0DZOYf/xEuUvA8SEl1qiWWOzP+VCKaojI9RprRR/hjtSeq5STmWgS
xNKu2nlpqaMmoomOmW4PrDiYxDLo+Xq2Kvu2EvkJl/ahyfzfwN5RsOZmKk0rZZCyPUwT7pG0doT5
b2MKvbSIbAn+CaZoZZDqiBoCgGPEsh9j+lHbsNqNcpZHNyyHqm1CAwt/gmPRDoVXqfSX/aaEuIAQ
ukVyXKVzxxK7QFqy7mm2+7tyLhyCMjmNRaWCUd1Gg3nQuqR5idkNQ0kHyN/HtcHpgrKKgIg/5UL9
auLbcxywz2rz19VPZz1vzVb8xVYBNX955CSDI7j3RGZAHz1WGKE4RJS2ewkfZZGXqNHweSq81EQn
S8U/JarN3fNuvQMSEdYPDjVmQjgqjvsAKWqTk4oVenwbFLI3ti3fOwhmdoH6FEZdn5l6ttbRrvku
p6QwTNdMKe7Sc1vdeQWBed0Wu4ktILMHQSsZiMPdjGRazzZRAzuNqSX0K36S3PCuBHvRxpH+aHSe
on9nr4m1mTaEUpxSnnX0ZPxN6+pZewZO5v/ffXZDCSC+XGQS9ganU4bG9N8n5eMwCkW8GSfJPywP
SJN7gLXI1JrkNV0xmE+mSi5lR7tVvRGZdqEqNOUd2B6qY7sK6HeuCbEoa9NErRPW5T93X6dAVD+O
7PlgA+ftDzsk8WglY5J1YumoVdmmY7JxaKyFaV1yM2yusvcVOzVd9cV1PnwSJDomFto7jZsvt2XI
5pzyUyfkhiuZJnqOXtFrKOxnYl5FXJHFW+d9CIWx6cRN6PRUcLGotBTJJQt7Ap9pbxkspLTtBM3u
7HuwnyipGyF3kRClialMSOmyGKkc3agi9UfIp23SWkSzLoohkQU62zI2CyfQyz3+zQqxJIvPA6pQ
Zg9eZbvslNx/X+qgeLlwt7wQIjIN0s/xBcAG1bv7PNnmAQeV3pCtdIb5Fyth16DC9eiUd6G4nJp6
hBcmtxPu6pnjhG4fphEFR2mbrLq11zXvc7LuImcYlIV0LsxSoNttOT3N4sMHu+rBzn4gP7dPC7bP
044gpsXsr3fPjcEfVBOtDri3eLH1pXre2nFHBvfDWeE48xBeE7XA+W4qZVj1ZG1RNEUJ0043dPYU
t0CgyIzwgvpGA4TdG1XBd4iEZZe1dw4aR/FSH9zs5nk7NpQDfOs7D0TCxJQQzozsWGDbmM990qoL
WszflYOFd6yY8SSpeDgkIsBI2PeHwlgbXlfN8hmeFfRczUBfXDffoeQEveJ5JrwuXflxguZ7PDIL
3fdqW5gPUHR1mAsmoBU687NQgcfxjAmuhuYJmq7ab/pf81Q27dQs6htBAZNy25RJGpC2YVQgo2+t
Yea2DDHy7Fq3f6CLKtyaongaOMSI1r6Ymap9Lj+Bpf8AqKUkfcxnHZplJ14CNyYyL4fWvAHvsWk3
uu8Xi6OuVNNEc/o484O9ojydGIjcXGD8GmJGXX36pce1fJxMWfI9PVlrajvZH0RMn61Tq1Q6NUl6
oBxYYoeHablNX8N0Kf3gmtRlJpEG9mTEv/UcPno8AOvTMksCTMz9BjZ4Zk8Y5s2Al+AwLHE0pg9s
27ejqTImwnpGM9UI0C+I6+tYq+1sHJ/mVJ9WqKdTSFr5BkdoDAl9f28+jx44Q2jUp9QXVr4lLTEJ
Sg+L/AR4+2PK/DY5Qus+Btz/QNZvGLyxT9FaQgQTEbPg1yBTzHaJJB5HUXVQh49kSs76cD5wiEXm
sA6vJDpxyGHa31/wKZPreHZ3mea2ZSrdJJjvCyryVsN2gQokFlXjwMXjCMoFLlBbsM0wCGiyK7Zd
dJgABkNJGRzXOwGhAu7z1ti6mmKxpzkem576hkn107Rl7xxS9j1S10KtnWWP0B2Tx8tAK/m9CCN3
PJtyM8d/eu3A0Y1t0eQkRBzF/T0H7aWDenCnM1YtKIoU4cT0apr9IjV6988RLmEm/B+3emhDxqc9
QtkxLw9FTNgPZPyQFw7Zhp3dXya8Gx6vjnD9Ba2BBrVSovBPw9Uq38DfdOZ7YJu53OWSe4klmYnl
JBV2f8y7yy1RU2z/D/5HAjHb81oPGPrG/XMnNBGrFE8LVfHwRBpcjy3Xppi36K5twJBsfopxQzEq
SgZK8EKTapaRLD/R9nWLuQ3z6Cb0PiPj42BN/JVSNzhfFACcPlfgFE9mo8UEHTDb1ChJcegsPbBy
P4jvm+HGBGHfJTHJo7AFV3cLh1YG+v12R46oNKpUE8NaaLwpQGA+zh9xU4hJRrnntBTWfQfUw44A
5XDimv1qT8msluq3TJgVdRamEaNBm2Zg0DDNTwSSfbi/xbX/gaDH0D+bzGhvoKVVjXT+HiS4jo01
L9X8kf0GulAtjkgoujdw1dzX+/GoJ6162Q/cj21glr5C5Q5pIrOp1T9skxRreQobW7UWd8X/oXuL
3Uzrtn5i2F2CwZ5grzxXHZMRWZX0VGz50b5uMNEgsu8odCEX3NqCSJI7KRz2UN4UQhxQruTNCWl8
mQDHGb2zui0UIBLHrTuB8o1hjvbdbrRcA5XW4XA9TcN5M6kTQrrvtbWPXk0pIMAfeRvGyM5O2HVf
iaKvYVAZHNa3thdoSu6uWvHBzPgUYaqMw1wxsrHd4cqRJ2q/QUvPVIw+VLID0fhPjx2ZSN5HzhOQ
YGDIMZuyHeapGzDvEwXDtC+lFVrnCPqA+onBg/qeRMD2XSPqUrugoeLoBEpMBpM87gym77TQudLK
hm+DcS/WpR9+3qpAkXrPZerywnPofpw5Hc683XrYw8pKAo5oAnhPzo542mrMAhSNw93ICo+2AcmP
fRmR04G05c04Dwt8qOmUAMGYSn7SJh5Tnh0al2vV12KQg8UzKnOxsiiUNmzoxF0s7BL4R6dfeGJm
jcAShPXia649w5Al5f2190FKwkWaFVaAM6BDeQzjQhIw5x3GxMi8BAuJJ5EsVLnWwR41Eg+EEPVQ
TgDd3V0U0P8hcEmvduc6bss2KESgYoe4kptm1RPcCUOGYvRDHMs6jIIZ97GMhT4dj0Sh2ZVDceN6
XxgTj/8OiK/dNs3pbROQCONvxkjwb62hwBS+gUu8X19xhevn3gs0F6hY0ZNrz/RqCgpP67C2+MPE
/tEDyYIkXvihF6YWxuXlG1Nsio6eWfd8knneqo6T5HuC7UITC7DFfA8OLXReHNhORiMqqFeqrNbd
TmWRxEdQUD7kwKF/5Hv/uOSiagORiHbbyE/QYHGpvxfIes3RQisGCj8OhLG5ghgXU6iZKfpBk+cz
mcxc0vpz2Rrr5O51Hs4aixthF2/vKKMEemWBFkpokGeKSRbz5mCNgGUBsohCWEPymKO/G1E51S8h
qQFVYM651w5n4IVCudUbQPqR0DE5XhvSjxuAKn2FsXW3wQrRGW2HTu3EQT6eNCx9fIdWWd6wJTpC
fF5QUqnlIp5VoPxwxVu/fQDLdRirIVZjY3fLFDTMC3VqvPWGo2XXv8/HJ0lgzEB7U89Wn3tH2sA0
7I7iN+uUvQdE+kZgQ1r5h1GQTJ5UH+gajGHbp+NtsUU6RxfgJ2PARKzgGuQ0EQIlI1GeN2KYEw98
ZoxsIMiuy/PzTgLcVPx2HJYxqzilj7FKu1YclyqaNszG/ImcPvoRgd1p1lhQHIi46izfaMjvcnxj
dLsEiFnzJQ+RGvoXl+1kNaL35/GlY+6BgQS+nzZ1hqSCT38hHyNVgS7LSo05aNq0nKMQkzAkp+6i
EYBNtn0toRD61qmHoO0Vn4XbHQKLrbnEhf2BYLBccs5Mo/yfqDm3ZKDlIXpRXODuhgmC60fRHqoZ
7ae3A8JJ9oyt5TeSuEB9wcxhjPouTKLQoQB65Mt8bO59OJEzFkZsQqpW1LbtO1YLtStFmBVJIR9e
+y+PW6RWC2vS4WVmzHq/ihD/qi/ckR3i3tQssJYdBhGrGyxWDuZcu6999kurSAg/dS427OV3A85D
mG84UrnmpOs5lWFTIoEzWqDm95oBJGY2jAtTAfNv2c9s1Y6kEglLHkbVdaPONNKSDqZswbbI2yJ4
d+CVuxXuu/3WtZaXAEc8Y1HKZFQTIIweaFDgaOz8GwFHMj7h2ESGPeXt3rS/tjPb5y3bIuW5OvCM
LGW3sIotLGxFEntSSX5z1q6zof2YYJZ6MwQMuamzdo3Z0Hdcn9EaajvLOc6ikBqfdW6AceqjyfbH
Gq4fDSB6YykCJreGEg3JtK4dp/OrrJXfJqZP1rnRLsZFcris+B2OnnnUnoRL9janJFIjn/jUHd+q
bgndFUfycp9RXJsu4Df/ans6K2AhKrKPa0j0Xm0sga/oNmYByogRhCS1KV3t2HoErlqHRVFvcJ+Q
FuC4cVnDADdF9RpSwfnyNnEdVoOSf5fmADSOA2KpKF1GfAaBdb5Kvj7SxluhXXOW6L4sbwU978ff
zmMLAwdx2PbjFn/sRc/My/2+S6fT32My8Ps4yCoxpasiQmB8oQ4/UyIgyHGeYZXFKW2dxagNW488
eh39RrC5IOd3CbmrV/vt1D/1IhUx4c/RAm9OWyE3WGqiqvcpVN+pQcU/2SJCcQxTQ1uTDNgTX7L5
Y9CBVaQopTCY8EqzJslQKeCyFWopLta2aSgzRJ93Jit80BhNHw+CpmPaqWW0VqLVR5oukTxCLAjy
3zCIGTpjcS9eCpRNZLxuIdHpB7Hy8L6pSsL/wHF2ggjmGTrVC85KiGjfMZj5diOR8kcGcrqu64S2
WI5Lv6VvCp3HAZ5He1ByGQfY//mpTCBtpStUIvFJjrmUG7VbA+pQhwp5gb/GQ29KIg4qJGLArE9n
ri4Zxn5e0Lvhg0JHoU9MgGAPGpKGbXLvvBRNC++EnmT6Dx5l7R0F+lSMjy6H4seNqjKQCR0IHlx3
U7QK5NSQ8uIJFy8Ur1JZGyWjXpYbs8nVjDyipXGexv6qBPv8Hpk5jAMt3NwRpGHRO+ZWhl++R+Q8
awqejLZSQmtg94VbPjm6tmsUkSanHbGzfHj6yNJejtpD/Kl69Ky1kxwicrQ4kZjfz0ohYqfwjZG0
uVx0DL+BfX8XO0Jeapvn3VJO6YxMr3pAeUZ1Aj6v3SxHGzxXeG0KRC3nv5TmkOe/uJujaRy1zo1I
M5P9XUCM9xkoSEbb1pI+zflVz8zNrgC7VlnxlGOwYziO/2ovp8vCfjna1/kSv+KhfIZCNyLc7mrl
EqhjHabbakoG/b8/LWmQjwBWJS62F5ejcFWHKvZ6YLnCho/RdgWD49r75hVgk3MzZq9rDdvjX6MR
BLpORybKL+0Btz1D62DkxAkLI417P8oCaameN13SW0ElY2MjIWdNbBwXym6D9sLmtjDzXP3UCNKN
PJSB6xwwwnjS16iMEZTVUPs+XCrmiOvoRadbSZUfjp9JTiCpjyPd3RD4RzSTSlscFm7V0umc8Pmf
k4u/CYkK5e2VuO3s/HcGAQde8EPD/O/lLf2mjV2iXA460jIPh0oVQaeUYgYRXjc50VOvps2U1x+I
l3+QBd9zHVsphuKtcxy1XV6dm2dR5+MBlMUYNmljcyXZ9GWmQGxacFRbBFrVO9JlJKTuPkJmwMfc
WXMNk1u3F+nS5WlYfcLR0VgC71Z+6HnKKtLz/nSAZERMZjN/ZwxfsFbF/lWWAicNwFGxVd4BNrm2
t90Bd5mrCqA5zVTvnRGFEn/IRJO7gtI+kVa/muUEon7dwpiTcfbjslL89tSqSivCmiR6RV0n6p+A
ULU6soqrzOIYp4Qj+AhRIStaQEzNzQLS+zzV09oyRLUYObO3WOQC3+XM+herKKEr4lt+wAnqBxca
w+uNIqyRjtjMR9aOXyDfTSyfigE/iI8e93gioJ+Bda8m/D7Cab0uHj10QxaU2dqPjFz0+PAT3//R
ISgtaCnlzFbZTaC2r1mnx7/l2cwbartrxSkPsod62GABtJlZUwqKqhx0HaofWfe/IS/mWCOcioeD
E2yEwJ4viccBxYnJJZdpd/CvBivxFLXc0i6tGivIDl19tgLCSZEdPLk9ranR5n/XZqYHC85v7+DU
dw7hUILHJqfYX2Uemrncj7CyiacTPKIIn6NvOmHBrr8k7u3j6m8mkS8Bogg19fdt8F2oaNkoEuTi
o1+H/Gthd3nXRdhc+wvPE7qkvKSTwnkwPsPWOtcpWVkiR0ixhJWJe7HQfCu+FX5TeHZ2Ow8i/aYE
bM89chMctk6qh7ycXu5AJwmgizJEsvwVPbK0RfBnte8vlLUfI2NvTmhz7ZRqhvRn63xZxaw2sRDg
eUajNCo0b9foS4OlW/djlxNHmSw8ntGq0BpPyRadxMcKFSgT0iWC+eZ26tCiqxR2WfYTmT2OB3HG
m5uySp1S5exTPmGT3ER0pIVyf3852Zn0C+aYl8n8S4eoXK2xmKcEZa3qIQUSPUH8VkeaKzcei8ig
ZKMx8kFTPLvABfoVe764xpm6KWzgkCmfBl2kz5frIfZSG7UsAaC7vkDCeCwLB8nztZdqz57it6db
vDesuwkEkTvGLuc8y5VuKrzMMrx9R3XboY+d0HctGuoxjS2Nv4Fd1/cyivDREZ37XWzrvd+ugu0j
Wgf00GIXZuYiC0g6n86Pep7Ja0djJ8QPkQLyNFa2/+j4R96TWq2ytrSdX6FXRfUZZqCgVVWxKKfE
Qk/+tv3oznC+Uc7ogWh7LpoomlYT8hJoH5662ylL6mMjp1sdptOgPuPfdDI9JZmmGmSttrtHRmdv
cfyXvSKFx2dTTcpIYu9Ur49QFjedZQ844Vb6M7lM9ILpIPcS9ypdReJvutUHyMsi6F4jlaN0K0j4
VLgUe7dp9RN+NpJxlZwQjSA0yKBYidx5nsuEPqMbPWMP0EyHMV2RvJRRfdT2D6MZrV/uH58LqLya
vRP3txsBeMjYKyP+YrWTWG2rpJk4RQUCgaxl0W8rTodP2f3bZLgDyV2ipJQSNyuOK3BEdFtbNSNc
b9o3OJXNmHPpgvJ9d2waRIZqQ4Igqbx31ZB+60Qsnjp9YjQ5EjasTnDY/dqoOEX5ncYcJ2MCehtp
2iBlhdkhKC6OTJPfR3a9itZc5hFdhi7xxx367Gnx+VGDVTd/E3U4DaXjyPTGIQYne+W6SYhzqAwW
2bZCA29NOxYbZd8Ozgq7iOelrBkVe5+o1WrWUUUimVxzKWGmMYeB/EKi7rzSmN+iX6MsH+6CuKyg
f0hI8NxTjoZJBpUjAexKPt6pl/yOEydMmLnCEFUbGDYAs+VXSRVFaXboYhTk8C4RRXO46eqo+g0R
Ns7JD5pEYRM0dDWoWhx/mzwTrQdKirtBOkiQjZjDIY3RlNKWww9ae0b0Sny+epe/pJBHS+q0B0O0
b09QLo6yAZQwYQBGKmEuh8yK+o1g/0Njl+pJYEjapVzk9iJhVtMJpO0bbIXNmnLa3BrcHx8jdk58
FPkLnTmZLXUn9eTpUd06Wqybv8/l9CVe5lr8HfaZLo+PRDrGZ3NOUa40nwpUrCQAhGyCACNwHIcR
ehXcSy+j4gyv2/ZwCpGdKu5xDkTLxjxifUNrDgSya1HZhKtDF38s2GRznK5jh7cS19T6nPIgDn4G
aY1xsMMtzyZDlXUlPOdJ1T9SKZo3AUdoM3bnj/djtjS3lWg77iJ+jkklMzAs9AOoUXHn0cEpZXqp
h/2YkOzK10mkADJs7RAYMQqRf+8ixCWhf4iFS+gr5A77OYBB0modKo3KJkLvOu7ThpoYNUlOUSPd
U3jh4FO7FO2g3Jd61u5YzNg0H7qiJHsi3MqMPkBdMjR+qNybHcr35Y+200u1TfmIDmLZbX2SAC1k
Ue+ZiIDiAioNGehaz5SRE8qtCNNfbVfmHaLPqb247zlPYsHn9k5xZIySW/A4JWa39HHUbIobfim6
qhGKWISBlFgWcWi8QwBBrW4hbkpD7iNjjEKQNNwc7o1ys4Mqyl2j91rkOMW3kO4MIOpNs6rXg1UK
k7JeRswbQZhO/FkW/HMsIsSYDsuK3J7DH7HL8U0+50Bl8RrnXX8iZSHGJ5F4lq8EYVy3EqWV8HRM
z95bxI6BAPqAvNWBVmEvlBKJENBLm2qCHYgCmZuRScp37Hpbw/v8Fh7dszyNW1GvMOm+nlAAbb3d
PC3uBSzl1x1l+ZqOQR0cWdN2tP24o01WF00V2YLyY/zw8ZcctMeRFJKpz/85ymEG3zbVmKZ2QZ29
+SNbQ83AelVXCraejMoGnNoKHdyiPAj3+qP0oXSL0C9/fXF2brytjCUx4yfM0LeWljThkg+KAPUl
YC7cm3sl1zixxK78Ag4C1/uVmpLlbou3XuzlE1K7JrlO9jTQrMNHDm+YIqz0ZxthuR8FdzEDI0hT
0THS404Qw8/ubJoKNdknxeZgjhzQQfwHbMVx59zhaPJERjgyJqSEMKH8R9ROs4OQgMtOm0jFLkyl
fg196ICuWGlVFHVzw1sIzeo4i8K+zG6TYPoZV2Mrtz4FMZdoVAqo8eK3OFdzXziZoHMRZrftzZ6S
cgGJZ2/tZ/LDKmRVZTcijsX4qTPGaWFjeDgjrMSE2dFFP5cviEmZztNBZlS09LqTX5Duvhaq6g3d
TrXcaUd/17l1+spgLIbOMRBKW5PfWsDLySbNlmJOZYhAPDqcXd7a34/Kwsap5VZJCysU3l23I+fd
2kmt8vSm+DOOR2P8rKP/snPPU1pUXbfwA/nuoSW1+6r4Zzh8VFjFriVuZpac8tVikYUN90JwA1zo
wdy9dr48fDKcFtkC7283tcL+pBaIOM9/9YIdNoHY+BcCSlIjeTjGQs+Tz/GJS8JA4RuYOG6W5sgA
Zs3qPTtLYsvGwDvOEIiq6Ae7/KATDEbpB9+f69A8YhBvRLW1vM7ca4LgSIFvdiovxLSUy+OUtSdF
c0kxhssW+f6kMpp7J59uj8+yfzfk6ZshRa3Axjs4hRUrq/CRSveWwtSjIc9wgXKsidWeNBRHBzMI
hf/Ngu2fTs9bOgF2EatOGTIM0HO14Ztjk6VqqwTDbQgRsdwf1kfn/dvhLj1WVPlGQ28Au0MA89N4
3nzoPBLe/rQ+55VL1IOK+XLEMJEt0WtTGXi0Z0b7DGucyWJBcsoLcC8yJgZjGTw4DNFI8Tk8ror/
b41/lfh+ynA77mFOohnvPoN2TlJuBMP7Py/Uk8hZKLtaAFrW28jKnBjo6tlWseBh8fEUOxyltdXQ
2cwDjzhVf4o+d0sRb+3g7dbvaOUxUKjeyRoa9Qct2cAv0W2cWzEDoLo8tQF5wNRDJ4rApaXzPD0g
bJWmCxSqE6jYY5WRH8X2QNY8T+kI6Hb77dR/mOeqHKQuhrgpl+Oa0i1Y0Ys5uCAmb/j+mA7Oegqb
5KON4cO9kCYAJS42TZkEH+QtbpC9yNyD87PiTfsb9INr9z+0vPlnHNcNGOVWmiIbLAso6opNMNTF
MqvGDukzwELkFy1Kv6jCgx/D0NyyN7u3pJd8zb2BEl9wEg+1RwoERHB5p0H5bGNJsX2gH7yI6Z1L
KNERxMmOxqhRtMN+aDgiMZPU2sTuaevul+GHhl6i50HeFZez9ro6E3htZFmips0SPGusDZEMg1ZE
WfgHgPkp4hZ4NswKlpoAxz8uDQTbsbjUpV9MuhBj+9btZahVc6aPhJSBWBxb/8+kqQhiYnjIKJFq
tpsR47BTeq5CcxDZ/8SVhKGpIMDcbEMtlSdnYnInPV0gjOq66uYFM/BckodpEqC3LiK0wpHwTk8l
mGzDs1bKNuGlLguk/CXdD8DexmtqdtUAMwPZxSaw4M8Y9p2XduUAeGayoCemZ46DCYlsiSu9e8PB
sT2pwxpxLXx3ZrURoei+twT7SyWcVGBTFECarNa+JMknJXYLBKOv8BSqmYJuEI1Vn2/cSl5tFJYs
F3G7/fgxV8/hWqrmvsxQVBu9iOXm3q0qbALrm4FVt6BYK/WO35ZXkMhMiFC7i4YwN8IFRdMdt54+
Q152vda7EPcgJfgdivto4i0a7cqOC271P9qKeSSJweAfLXju2Hv2qVVW2FxfWU+LmNhHsh1FEHU0
JDtZQklfHWf3/9l3L9PWhNegzz7YiG20+hSTMNWrxcvdmKJVHMoCcufGZLw2MvRO7qDXjLDNIw18
/GnWexR9RQonMkTXPwEBdG21phqVLc/mLQ8f8seXy9qC7vQIuqQGxMnrPDSAVOTaLpU64ldIBE9L
7DyMNHL+MHvacez8KX/2NgWWGCFnB+Nhuz9vvcvyg7SyVFmaO4plOqfPY89luwsw/8iRQsazOVBB
GGyAWNb4+e9LsgPKP5RGbES7fya4U/T2QITJhSiIl9oGZjg52TqZEpy0eHzB9UkjL0uU8aR9DAWJ
ebXvxhLtgfxuSKknKj9xEtgspqm6OKRjMLyYWrhGvgcK9ShDwoBaImmXLfrjWF0Ha6HdZTmY7Ivq
TuvDTNhyJ7NUe8XhA+e45V+mdt9aQK5hsCxKVU+PMGXVpuAn5r4mQkTGTcG71XJcwJRZh2c0efSV
0CHXMa4M2iZAFG+q0+jWBGNCQAMzVNP87IXE/9R1v4fpFNNp0z1QYenjOMxA0lHY0JCX4Se095NH
onSYj/1hoHWYeAqL14lnF15vdnqL7XR3VMlkPR5n5r1bTe51eQ5mDjyHlpZiaAc2Ipn34pL7nZ1F
/2wMXv92nXJQDchAyEaHDzuAqROJw2MootamjP8Hdrz3NzH9vmr+fmVvZWbEcUBYe32ZP4TYzMJP
iGRuTCiBerOdWyiHuMDpLa5DIBqCpdyFn/g5XIVjDqv2vR8C0MJvF2MMkPuqqE6rTsQlB7FUwi4v
G5qo6u6GDyZfqYaIo+lTvqarfyJbyCFBg34FQoIMxvVpfJRhPAY02Ec8iE89QKqkceN7y5PH68id
2j4xfK3tHB5PqIYHJXWTrc/6AmvKik30TgMSZZ4KdOrnfOdgIL6ELlc1OQnze0Lv3+jtjOhjqmDx
FBIRC3IBsJBoi72bj8RD+xFjOaa7WVIaMyJjy3OzfdPkmAnsJmgPngOvVFggB4aYs9RTGA7TU2yu
wH7SqDi4Bp4lq9zoeyALasZoW/P6sW25pxroZ8o/YLAfbiipKqJD51+Y0qeAXliF5vu1on3ThIPV
NK4BlypMRrLV+FDHPjvab08KsCYto+B1M0RUEmBLyieamdKwjC8lAXeptJ/Xu79DlmDPGlO7gmSo
GOEH8bMX2tBCZfMffZLJR1JxNA6SGDhEiJLU1ifI5NZIRt+SXiAhjO6P841t6jcUWvTvGFUz9cmp
3dKKCyt7IHuTJR/qDEW5AEqQ+zskgGuMzTojGH1zrY9h7fg+lroAXy1daeK/GDy/Nz0jFr/OW/Vl
M6xRm+2Rd/InLvYtPa2loFS5SZ1d85dEpal2ZlniEoOSHFSoD78WixFljqw9I0n6BhJ2mHXsOW3h
Nf6zFF1jDFe2A5eKA9asnDNymTOYtyoo6aV25DptQjb0Fdw+KQBkFcXss06m8fJl69lO7M8SJBE8
R2xqCLLM9UjC9DdUnm1ys5oslk6QDsWzYFtOzHxlTIydqXt1FIdSMX1mRQSBX7Qh48TIFJwZQeqB
epVJrGH7vXQV854X0wN8n0te0W/+x6FvbXmcH9K6lCU1GhMxuMmsUHUe17HXAkEcxIepoai6EnFB
AgGOXlV3p484jA1M6nNs1vpPSDXHWmOiev1eiVKQd9Tlf44icn4cSWKETDfiC6vp++XOrp1Hym/t
WNHA79BVLRpYL1VsBEwzY1/Ohergyu6kKtrNAQjp/CBUb7QxeUwKqQQogzKj1q0lUIScJLBm+tRm
rLE55evhfYA1uBs2fBAtkkGdCMAUAFF9zFETe6OKGQNuOo7YvXgRvN5R/wpeyWOdbw6xWByRbF2l
kJSWTIspu0Lb32KSApy+ybg7JYCvgTxp3s7jMDbQTYKkHwX3xO/Fiqer2HiDlbwLNVs2cb9/gwmh
AOWyqJMxecXcCqt5Itk9oWGOlYYQ+9TeqNjeIY61CEldixD6OTYB/4o06+w9tFrTRKoUh6WxgW8A
fu0jmvaqBpSySTVlWroTlmRYiuTP9KFVv/VDsJRG/PFmlE0+M5MQeMQH1Whyrjo5en4osZgqVdsW
MsZcvpk8bKTuT4eBtwJ4UkwhelNXyWbNSX0fsSfHOOa2xyQfdP2ROGA5FOf8QT/jwHd/XwMNFt89
qhDEJkDw4uw7PvXBLEb1cCD6GAJv0UMMCCnapKVPquQG3YqCADp3ZmSNlRJWPOSFeJflTqmy3hiY
mdppAOsJYMs/+fxQlawWxfI7P9byzXlQhm3fALowD7wRG3VHJ+tISuankpytfY0bMcqSvaJkW4Jn
O5/I5filHvcwX9Nd5JFkNJESt5YPGD47bOLVys+iy3gNFcPeA46LfQ5v2IXk6RQmS33jR1fnt7Uy
Qxg8MI+EBOuOlzFjtmU6SJe6sNL6ziSTsKN9Nk3H9LoZidlNOl2V0fNC2Bu8AG/5sbXOq6BFlDTK
1LbsY/vfh6RL6bZUGsRbTD8uPd1mZdzLAPB9obRwE2G8mH77UqbdaiMLcnwhVkxwlkeRLAzufCTy
S2JGjNsOUrGd6uk7EKHoBhYfQjR4ZMUYfHslnVEs5RtOlU6oznUdAcrWhrxn3k08jMHjBmJ9b3I6
ZoTHuS1dxPLP6SThkEg2TehWMyXrDkhRg1lR6f3cvnjGBbITfZClSoOtuBhbqGfDfy6o9DWJSRRQ
cTpCdosuZUSA9PtbZ9w8qn/gVUMdMA35+BN3iohs9SMvH8pIahIrkl5xPDJH2zk0/IT5S63+MMRi
ifqp4Nb9JzjyDPLAoAdfZxYjBa6dPyVevCwlnAK3sWlJ8c2bnXF8ejhotwnGUrlzMgwdUYAKOlMH
MY8VX72XCeeRCQcUw/yyzYz+XFNQxe0TQpsKQ3a6YGe0P8a8sri9DiG9tCHMZinr0CAyknA5zugm
ITe5kx82LymIh92nVbtt8BzYPEg+aeKqgrU09pelB7oOyIwdL3o8NPaUOcwow7SW1SH5e28jd9rv
yORwBipJWgYgkvWhz4SnXaoLleDEa5QM51uWl7DuIx8Uu9irlb9uYpRj1vf/KN45GBX/p89C1AoW
I6fVlf2FGBGGqbeovmTSot9uyvqPIc8quiiCuaS3HY0H5V01AVmQwXjbaEuLPl1z26ZF8RxZRfVJ
TzjeZsGsZUC9zURhZzCpAoCQZ19Qvc77TSkkVZrQPL+v0Bq4xVsM1b3zzUfmhrgPV2rVqwjkpB/g
hz10RX9IRt6WDDuufipVpkadMfm5ctqbbaeL1FLfcJxw8CvqR1Pngll/4HFCtJvYm3cnZxBHbqlA
O9/qovaYT9/d5yWCAQaXyxwfFU+JchouaUyB9rhdIebXwEnpoHgeqUhqVnsvocc1VheO689nzjbl
Zny3c2DMx87/XLvKMZUIP8nQqXnMzAZVuJ0izxZsehSXJK6muUGp3exRxZQoA0Hvs7y8VM19YNOS
d9paDyw5LY4CCumkgTYTbyGdkCSCtCz2XUMhnyhGEv23fUvRu81kmJfDMGzjkmpL3PwsGsoWHhdv
R7mbuL8eb932f9RR30N6hAFIidIHHafrQS6cBKp+R+zXx7hw2shX7QP0Et64UsMKauRGClnBevj1
/LNkME8Cduj++uVqfYfkRjwMAXQPZstB9fpj3pUHXzRJxZjWyq4TolXaXCnweIcXalL6Chg8KLWK
wLdXMmMNqtSZBn63u+F2IxxhYkfFPBi3p4mhsQijZJt40jEaFljzgMm4ETmkTNB5dKhCorUQVJzp
RrW5/Xru7Ibimd/WJRXEafeJ878iVn7zINp3z1eA+NAfNaZpsffrZ+rCxbBSTHA7LchDiMF5/JYK
qGTe4FcqIYKQU0lhSqrQvWvYtYF4ni/NxyUZCYeSKcYBeGfvmC/elp/aPhu34KC3l0fKYgaJEoYx
2L805QyvzoRRzSfMEWOpqkrUKPcGnVyeS76KjrjeyRWJL332zFieMuz96tbodtbUzRUavd+sH6RL
+Rssub+aar6YtiT6gU+Pe2rWQr2tFsmeKJydYnsxa35tSbRnjEbeX3hj2h9mml49G+g1KCkyOYNv
ZZqM/PxClTgkk+kJFRtAlzwiMVgCQDrT/vPjZbmIZla+WtDc20+xC6XWq/+UyJ0eaLkKGDr9/BAQ
dpNysJP8KRl5KVTLewHNR5mRN8LWlP8qQxq+gwE+Vomzil5tKCfil35Ou9UVWzzze2VdkDs0eo9e
UM19qqgM0SSq6bpgemXhNcmp/hvooSFogwrTDKyUHnEf2xpzwyPS8aZFF7HkFNEUF79+flC9rtOa
6xwDmTM/8Bdys+rN0gw8/cWHsHiylE1VFfPca/5OnVYi4Fsa5V3fqrK1QqlpTDOwET9LqZDyh+b0
CfaoFdVuMxNgzRHzAAKK+k13a/eCOIYEYnb6MTk0d8xZeHPbOXJ4QH4L/UurLB3Do+l9QsEz+r9o
kU3P98EVPJAEjSSSpfQZ6YAziuy1g3DH+GD3FSE4rPyMXWkAqBpmIzc1mxiXKsN8m7jqoKG5TEQv
08op6aDs/sK8IMHCdlmi+NOEfEhb+Oy+CIMoMW46mhbi4UpbvEqWsL5l+EY8HqwjYbwm+7falrKG
ccQ1hhx8Ttw7xjzp/vL9P9wfXZdfV+BW/z9M+1ERNxmkjJs3FEEpN7YRXP8W4OBkPq0zADxGyT4i
gfJkd/sP64E8kXd6WrCJTIUTueWdLidF+5RDt8FhqoaHmY42AFE2fJHlhFf9mRh5S9D3bQepg20o
tjDHXUersfw5OovZYLYbtbbuvLvanYsTbLTg+Kf2KIRj8Ap8V88rR2wW0+Cqcxi7ICGkfBiJQNEQ
gtthB2i0Ppffw6sEEMuWPVNDLAMSNk5oEIuQOzSqWwIKT3PghsoM5tAYpjRRofEk2EvXIYVPIJTQ
FsKL9J+8HEQFN6JDmeBLKmha02QXaTwapqdEhSv+VybwLPXn5NdI0I7TeuPPoAUC2gU9A+Hgs8SC
ko1137EESlM4MiCQVH2KEQcBH6UF6+5iWaJVj5T3vXLxG5O2vDR/PrB5GjeVE9y/Z/jx4UDeNQeh
hkTc8fDFGoqryokBdo9F1RumIy+w/1HRF7Vcy3g633T7loLjQ7EZdiSLdPig0R8olCb/F0HAengH
ZQ5Oei5dB/aY1JZKl2ll3X+AFuxZ0FTdxCARcoZ0ntBPsy+HrqRanl5FSMMog0YnwNprEUb9XUhZ
eK5BocN3tM2WkLeKZrlafKoAFnDbH57si8MYjsjffG45MO9WhXYmuJsQCu2lUoagXbGC/8KbmvB/
LS/22Et/dWtfolU4mHrC3zjHawyw8yJb5re+ocafRxoitFFnYahFhXcmtHvSLYrsNpAD/2qJOLMd
E7nL+GXW8NpZWUA5ZQlKOAc9XC3+dcKdLuvA1tglRGLa7viLMHIBgiBHX3P8Fzr5/G449aOE7z9x
oo+2ZG0KHwf7kEk+frJU7vCaqnxo13Xuh1PE1dhSZ6FFnsW4TevNzki8a7XArCmuwL7a0yQmMysp
a1nUiNcA8LbrAq53u3INdQyd07snBC3QymGGdZyRtMO1n9+E2UpmDy9IGcDXSqL1TQnbY+9wkpgH
8wH8xpRQ43xnS0EfJTU07tp1IIKVaeiolMeiW7wUSILgFCx41jc28nqSrIJ9HLVcbzgmY9+l/xQl
mjARUGXjPglcwoRRQ/oSx1WfLl1SuOadmEueF2Av7lERE478MFyC0UtG9tIDcHmZmaRYm0cpe8Ia
DT+UeRdpNwxMNuMXMiuLbM6LslzxLLBePPVB+EHCSX83lmZ8bUWdRWoaPfccjOVfY5M3THocdPss
80B+CGbApLuQQBpd+4F3aDNSsTn2pVFSo3VtVarWE4ghS4Bnh00yAE9F03tXznXPItqSsIHQt6z/
rBTM32lIFN9toqqAxHpduS5bFrt16I+pxl5IVs+E1KABecFJIHr2Xo0XgjJJ+A4nhRwbpBegRSPP
NCijVMhlAMj1KHqnZSjYC9OzwtFDYYJYxfmEOZQxjD5zbddr/3JNyEYmKnG8jKttXapZXJJjV6b7
PHC9U3nWxh2VHU/aqM1U78a2SQtND24CC0NJpUxKWA1PsC76NqPySpNxHpIY4aDnvLRiiknJKDA6
CeVEk5pZ1faTQQcKppnpUYsFEbnlXTVDfTGP6Cse/6E1hQ5GfPowvk3HNXDOn46PQBuITrAalOXs
o8b9EBePdM1i3rYlDVkyDuw8a1QZyVe9xfoO9sM2r3dHo7/7mrpnppGrw65LYi8LedTsht7VK11k
M+pO6jdikuMiZLOx5EvJU6AGC4iLupMR1Yq4cz7txpB6jLYhDzIIt+QKXOOIIPQY4DAa6vWCOccD
CXtHjiK+gNBJfAbm/qK3ARy8x+PpYzkenWpgYTcvQcsAbAZWZ3kC5UvjToszri9yPnjMsNDyAD7h
RYdjsJaEI5v8Iz9R3IZKs50MCUAjqxZxaPsMIAI+EvMvXiK/6HFDBZejGE5vt2ZC9tm1zF/U2HIb
EBJ77yp3FITxy2+MvP3lSdHG1G+oaVhGSyw/ib8DO/mmUywB8Da98VILwbphBCdX8vmkJUvw0+PE
302IGS2CNQArsvb6Ww6IsJc/7BMyARHePEj++gy6yF1xbRpYZMdcwa2WmNzVIDUQVOKpwI5qyY+K
B9Vf0DokuRik2AxZ80U5g7xCRoOpkxDpGoW1X94gtWkt1T4LA+3YimGHfitcEtL5+8SosX3bw+S1
Fin7YEHtCtj1ysceZrLiPhPu83TMlIPjKngFrE+KsEnb5/dOasbXRkswpyoeybE3fc5MZ1QcsLRj
dWrU+w2fEc2qujKlRO47qjVPgJoR25BkEAl4gQkek6cQaBwzvkmSj5lkBmGiQY0QowVwLp55r6bz
QPWkqqR6vSGleyHuZ+ApLT36EmQF61aEamfDfq6gc1bDwreRHHod/xwzlLyRUZdTBEsePsJ+4QjZ
Ywr4U71dda1806s7XnR5hQwVD/8TD9dsZesRFDFrpSyQ4C1BcuBgX0RLHtZ4/PsFAxt8Io17ardX
W6IK2JTxcxorOKClb6CnXRc92xLOvZvWgtDho6pK07euegQPSEKugGp+r4+9lMCMhnJIvXQUh5Nz
UOwPNByvvNxAHSHgc0akNepjka7a+cMH7ZJas/7E3qAzPoqQUZXMjKTd36wSMsEuSDl2RUZG/CMo
NrSzR6v5NdoF2qSLvtBVmtZdKabUzQtkiS8pRRc7aY+BG+OZhmdgEDnNBPPtwJFMrg3sI/ACvjqa
Aeij9jzL+U29qJpNUU+fqwjnDkjrA9mCtiXGr2yvaP1/PsJCz4X4UJC72LtE1HbfWsOjsjhSnCpv
7vuvMnJSu1H8zRNTYffS6pu8E/LAOkDEmnNoXf6MuZLz9ymSHDHqp2PAaQhwTVT9yIy/7YmaHlie
y/30tbz/RHH+bNx8nFkZhPEa6seGbb/cmv/prV2g5TlCz4YtN5Oi1BGeL8i8ttUdYedhE1DS7cXj
uISHRGzOK4bP1qhWPEOFIYRlNikytZV5GsldUTF+EGeKonajIqbGKK7Epblf3uTzVH/7FeAn4B7a
nw5U4Ot3ug/KR3RgC7wlQ3ITKGBJiECiDdibGq3jTW7kd5uHYdTvfdYDe49wWNADLrAw2NiUVokk
sVWBZRAgrfQMhwLEacsdACa8u0dndBGReMH6ke38OT6iVflzS3RBhPOJmKCOga6nb4EqsTVgkzCl
I3QnBBo3Nw7MB8HHAdlzLPnogUfEXTZdgEbSksAKJXgrwswNE3mX6TGTcw+FBFa7a444xWyT4M7B
JysWyOS9C1/PtY71Sv6dMFt03Vnqx1FFcfPA7LSrTUa21+jy155HxgLV6DWPz+3z/USOF7wTEbZB
u4INU9UpPRwoyRf5BDKmZz5OPEtxk9FLJP+u2DQHfKpTsnse62E8hNhjvWvao711Fb+CnMLmT/lm
qpLSj39WeouaCJyxGTGAAppu6ffHu4XCjhPOZeQ2PgMlWWJilCIFLq4PtcCriXNuIhRH72kdxeCu
UlUEmFR6fFLTiURxktLdEeqMlPu4LhxiHhcecsVoOJ21W9OBzem1NkZb9sRe2thRs7QqFEb9SrTl
+61OjIQ5uMO0dia+u+TRHFpHR2scblGuskGS+1LndBZ6n6LhKR+Tp+CwnqGbOjBw0LWbCyuEDCUk
7PCmDGrMmc95+3BuHN6ewzPT9CHzyfvmltFZIsR8HXPpaxZ/unpsLF35MMZfNPbTCVuKybvFUueZ
4Fvkb7RaNaWZlVMva7mmIx0a/h0N3V2U7UiMpICPk10G27tvdh0KsxOEXczePjdPhIvgrcxtFzlx
PyLTTAkIMqMUhurlGWtTPu/JnDIQKIFInkmAJc6pnROLlPECU3Mwjy8SvFf6sNxvgBjUoTY2bjFF
ta2T7nDQPrWHWDGGV9r+4gkPfK5qy6hQpTa3sGjef3j/igas+hMunnnuWMF/ShBaS77GEZXS2Xw0
R9JX14wLdPHi5sf6W5cLrThi3Y/ShD3eiO4hNLCED8NE3H1BxJGKTR3TBfZ8hNUyawhZWEd5vCqJ
ofJr66MPYMNcolQDAu5j76SGlMP0CXoUARNMaBXSVSUQxGEqUc9lLUaHLjAzyGiRRjIH7CVZ0+/G
XnoCY0TUb9zI5ui0Xdy8wLesgC+kIk6QaQp+IcVTfEJHpqyurKLET6rS1GcCJSwcHN+nOI7GQSzE
WTU7YiQJ0KknzxblUagdnxTPPbdrVnTZocrqZA8YhxXaVaf115efHMGudeqiR7pJR6SFUvgjqSCe
/2kAc5K4eYL43GXvwHA1DMJrbFhMipklHEV7H/Sxvv2DRy9I92gFC3D7Kld4T2NKaivf4yUDlSZF
Qh+BmH5aCvR8ojxUEyf/8qx3lP2O1KQ/jEffFetna3OLYYD0E9LPLhP17vTPj9EI/BUL7vJFAx/p
NW3RccVf/gsiNHQZ7IgxxxIwd0WynSoa/JhtvCXxcnbqO3fBF6rWest4qeOKwXCdDuj/TzlwtNno
7WNJz5X4eyqjD0cL5iesxy+AQH0unLDbln41XkBxi8htzpPR/8/eMIjAAw5AQIWJOyVCwoh1YYI6
WRGAlPbSLMJG7NTw9Z9CP914/luIFRbfEuSNtuD/Mw/UIm9C3I2WFb3BCcqn4G5Fu780PZ01M+ZL
99q/AE6BfsNiaYr4khvrQfeLP67/NIUTMNMypH21fE//BPgE73hNNC6OJtl9Zu+oF0OBBdQFVo5e
K4LN9JlUjhehoVuJB8y6szqf1128vGp5t9H6MNh3UE2YPFOdVubmhS99Z9Hw19gAodXbqh/uin/R
UFIHaeJjpkCOctYpHWki7eLNgbE2rUTf/WjN12q4nbYpsaUqJnc91N8RGzTTl3EajFX1drxB8qfk
eN7vNhviIb/Z84zrs0dt+V8bZ3EoISknDNqsaHZfjp60o1N09x0r7mwFFQX4D8OM4WkKsoot8KX7
b3AIAbjrk5QZ/4taDO5vqiSjwFde8V0/+gn0Q0wA15zibBM47NslUsbGJMlqqvTBz3gj7/lNQmwZ
/dmrO/5PJMEYQ9VVdxmiL+ctGhGSg42aG4fI4hB6cjV0BdWcMIknoT9Tr7dg/sLLiF7RP7R9Hyk+
FnTsyQJQU9BxaGsIC1eR0xfnQKNSUSmCNUx7Osukl4kZY8fVRFeWgj+XcEczN7xicZUqfS70/A22
N6DsReR/8Eyy1iuD5Hvd17DEO1aCEWsv+xlsyLgJJwEzG2pfcAao9IjyPN4Emi0JDn08a7/aOeEb
BLwdyxm4WDVMoL+HmbrAvj8geymYOv8UWsya44dGLBNFxy/3mUdA1+dOWTS/lgD92qWKcDsTkHM1
uMUeZiiEvPoq46CZ39yPr9fkbF9ksIbJDfgyTFr4u8WFKyFiVClOPu2vS1brmebVgP5U1Rdq8Hmy
Gc4h4FHLKl85I/dho8IhLp0yocgF9LLNbQdUE32HnFqoYT6B2t6Aje+r4/VSIUSfjaiDRlMeJJRW
K1wFxZTYwzqaVtyoj2W0kMKUMiVjB+TTOWBqiP2NnGKb5QaNniET0Bpjeqe6FPSrSMMiuzsEs2eo
BrbPLqGJyENR109nUx2OIfgzUlDrD/QeQgRlEreMI8uicPKul6YDXDrYHSsy+IR2rB1zCe02WHZY
MVljOGfGC3jbBxF+2cKpSS5rfpXSLDm6UWbG0GdnPVgaY5dBHTvtCap2s+3uVvXh+uMAmNmVsGCV
Lh5pwjt4Jo1go+ecZDT/eDEJJPl3qvOnVi1LIWsVxiSY644rXOGdadyBW3A2B8/J9nY8vItgCf3l
lCBO4eZ9TlDtSAgBMdC59GHYlaBEo2JBvKhJ5E9nKUsr8/89I6uBZOOq1kexN6zuUh/CJf4vmGYx
upwoLVPjtSzN5rq7nMe7XZlMAf9sDR1v2Uz8crMzw/wCmxopcVQSbdHV1xKt8RADbogihommRsIF
pfRiS0Hg5NqM8pVN0ZD+gMV24WbVaIpYvvuHN6LnSvIdH3PBl0Xi0HLza8naAcChjT/Ec7T1+3ZT
klrlfvf3J38BdyBkTcipvKRqNk3NSQxzUiJQcDZ97IuKNYqoGxocOz7uwkGDBrWMsxtpdc4sqndz
DEonEh2vByZkvM0vkK8FM7K2MXYeMYd3yHhNN64zSts+V8d6LgeXanP33ya/JeCPT6YdW+4Ir3Bh
RXhaXP3iov5pHvd8zBq0/iRUI1Bydl9SYfjSr7HWoFJaBG/nyWnLcZk1w4B47mM4aCY/+J3Wbpl0
3/uT3eGlnvDcLkb/ktaQbK6eJTdlB0DsxSsMvbtSj/ZPNMOEZqKjsDRwpAU32CVCjrVKTtROv4bi
IX5Bm8M+Lm/fhuk4LrFLePZBbz2Q6LuxnvIAEQh44jT6yxLtVVQpASNBvaLUdYHDfcLvhSlgShMN
QT1jrHFv2c8I+d2ncazX0P8QZav9jPIK/656ARMEeGt/dw6Szb7z7ORCA1oF1Mv0SNTbxlKCBM/9
b2uZn+T5LFgaXf2I+BlokJ1uKxl27UhIcclodyRMWy0t9FfMfHM/KQQrSddTOLOf0Bs86doPtLdI
cvvNyWMdGRB/jve0xK8wyt+uCzYNpr50oi81ukPn/9RlEH+73iKBCStc9P/eZd/q+nG0Tb4LDN0y
yUpbKol+nFi3Dh+X6tWDuw3lAFxHsP7or1MckNjf4MQLCaY+3bFFQdwyTTl2AsqKmJ1vx0GTEykL
sbbQ4QiElqHfGDYIFWGOIgE0FOpqUIJRkm+CqtY7eoAcMlyet9hO+TzfLyCscT6PTDSUFlE5lLHZ
qlVOJLAYAKUTFBeHXD94t1a3/R5XeEy7rkAZmXujWQ24OiiKSHw/OUv5+E6ckedmSnsu7rZ0lhWn
cpEvfMXodPrL8fBcUOEs94ugbx9Q8TnFoKDtsl4xGIouZSfeT6zUFxY+wzzvGvKIU3RQ7JZ/cJqq
Iteh7xXGK9Km7ZGpTYuxPfJPC6y0TcPngeki9rsSInjlIzkaBiI1MjJL8G/+3diEsNYMo1J5HisK
fy6wJrhvoK9dOsQfkkKXSLw6ATvN6iyW0Qi4hPlY9ikmLRFOr8Tb/gYabxQ/J5K9puTjO+xWXECB
eMZuIo1UGieALbdTMmyaJXYzY4eJJB5EGR/+lkcquKuY/1mZhELdrzouI5+hf6X1Tyha4B4QJ004
Bsk+xuqp2I/GWb2a9Rf/pUNmoG3ztyReopALXqvQG+tPBOzf/rma56gsYxsUR4vQlkVhh+yqNQbk
CljIP5cT5By2Hpbp90AqWCGIyFk8tf1283yhYWcsyki+ud2g0EnEpX/AO2KcLjqKHRxCdabwSM4y
XDnq2R/L1F+EQ+kBHA2jWm2m+13z4n4GojgDGy8euulZU5D9tw9WCRDnWhWb7GcSZbQaZDB1Ws0C
5VskFGhIyI7aeKzFURIx/+CTXtO0Ytwlu9cJIqCc51kVQyprJay4D2zC0qIcDu1CqZkt1XNczDAB
yQUR9ciPJcnrKZCGibbFiVfh3gRkSdcsjdwzEjYzjIIG+Cg3pFuWgSkAKGqpA+lTNhMJ8iHufq5u
DLkUqQlgTtp2RrdybUaEGQE3gJSjtZU1nB/rw5oJZYdmJrEA8DPtj8C7RvotKB36wnZne+hqm67M
fNlQgUNR3DXLV8HQCGORgvi1UbA8K5ZFVM5lUIUKRvyQ8o3TUwcOR2xVqsF3Q/eFTEnAaXis6gy7
7rZtuIDI2YnTro82is4SP18skta2n3VLpoyEliGLW192XyjjWq8zvOw6gEx5H45UMGhzAUfXoilM
ixc/6vBJWPS2c13ZLxR+wPqF92MjQBhkq2mmcP5C5cMjMMLRWW+ZO1RkwODrnMMY4UyZEbxQ5TUv
+HoNd7gm390GcdOJLZfmxpEAnrNB+iWYtuqm4HPMC1jqaIoHxzjUnDZG33I4YpFUuUT5uqNPSiSx
ad4zM2Ynt48RDeRGJ3Req3HPLzbvUI5/5PpSxCWNr8ONDvCtEylIVnpAEf78xLfglYCSYr520512
i2ryuthZwQBWvXZ/CBcn1+RJ1z7w4w7+8imQeHoABAUJV+4cPPpZszyl5y6k62J/1ZbBq2R63cMG
E671dkGqISJbr7qrmY671MOA9roPPS97w9hxo6HEnU6BHiHBV2LVqglDHKS8QtLJgn0GGFsqP48M
FMAq4RPNoNh+NjVMAOmfPePt9xPVzO21ZGxVvYgp56mFKmIcEq7qPO0d9gIhsVDadk8K4kPHi7EN
9Rt0KaIOdW06eafHzTkP10pvG+3Hkz/twIatifI1slwyA5zCSJN19tbHkgfC2HA4ZmrWqa/fXqAI
2ectqF/nw5so4xmvhv9JfLdvZyrctvVm54mLcTeGCZfADcahD6zqvFgB5CXeNvpMSYMBxyB7LzzZ
x/1i6XuJz+R8qdVq4XCKmq5zuSg8Pj/pIuvt6t7ORWrD2O8rpjeCZK6MOrNDNmlPw8DKJ22+6Vxi
JFhLlaCgSWSwcij9GDanZwAVYO1UdelySCnJPoeB5OTRgaG0mYqQc+teiYhusGEgrkbB5mbXE3VS
mPfKmO9ZwKoejXWuUl06ZgGdjwiB4UlrSA67Z5D6KPt83Y8GXOm1pqVRn5eo+6aWy03HywZ7QAb/
avk9tgthm66ERv8znjNyHWT52LCfUoBGKVYZuO3EVORl2VU4XBs0267HKnCiVOtmOpe4W1wwEGmG
NfQ/D5xrdAwMoMB57dc32yVsfM0HDTq6uT7qGxEQc7fY7Ix6sozGmm3jo2XIkP1nUl9GwlnnNBx8
Zt933DPx5LYkrSkjDcsKS7FUz8GKCTYeJDsRcos47agVXHnqqR4L4YAinF1ChFFr2o604pEcL9uG
nuum6V+yZoossGepw7qVNGepfct9Csety0tsS2tmTb7Lv7X5cQ2BASyJJKD7fH0nYw6G5LXpFj3s
VGd/lECyjezoBn17TnWz9BsAZAmDmEdAYioh6S6/RfuLgoSoC9UxRKpGKcx2QYqOSb03GxbcYiJE
9paMgtNLT6WU0PG1Mo2aFN/6MXxQmkGBVrHaPcmzUeUGInGuKUy84MqUGADgD3gPmcJCvjJpmYtL
OXuIsnWlvcdmZuZKMcOcEVb7ES3gjXGT4OBQf12dUEBYaUYj6g52+c0ut2j3csRCdBnqdp9ObxHH
cZUzfeyPy7NYDFXTkzxDSt2EvgQqUVWiQBmgBSB8wTUw3GGi7OlBSWikRBtc6YShinZYA8pIP6/N
qWSxfenz6KtsseV1Qv2xeG/dbCbvf0rhdP549x+ectk5EzQ7ombg3HCSsaoTmih9OfIIHnN27zPv
EgBZ4nQAu7I2pAGwAzWMv++txubvrwfi25vqcGDxnfaj8wwAiwG43xN2r8pErm37GogQ67dA4Dut
4O8AA1Skx72dxP4Wmx66x+biEl6J5C5EXAcx13XwEp8FiRqWL6ZxzAEm9FIgx8Zs53YZMYmnt/FM
1d2BbdN/RO9/Tegs4+1hBA3AT3utYuuewgu2y3ka9SAv0yH65n9edqn7rcDvmniXoMZKrvdLmhoK
3PD4D2U3ujEsjo+KagNoC+Dgk0kRg26QSFv5x1D49/uFiHES6+rszFDVhMaeW4iFtatfCnHnkLjp
zcyFa9zHNlYwapoiHPOQ4y0jpuHpUFZ6X+SHmSg2gR72KUUT1dtRqutEGWI4DuHVoY1emE+tt85r
6EvZiygOMcczuHnYoadvYO5/eYRT6QqnJ4RhnqwR77vHYNUpI40sz+Seg4zqmNez2Xz3IWZcT5Un
UH+PwFZTrZN0XBKDJgZyky/tnym6OLTto4tdRSSJkeBVGXOY7G87ToXdlReB9PXyZg8TU1TRnu8y
zXKAglVv5WYIpS+dqcq57LktbV4tzslMWzmTyghDC+OLjsPVXINTWph8W7obikEyxYCwKaHDrt0F
EA6TEiTXFM6n65QvxJYI1SqyjOF30WLcjruiL/fFTvOz+1uOAEgZoerbYKM55H15bHeRDhjyqcmo
B0gGOtxwnhynTce5JiEjpl42759ymfQWNa094iDkco+JATKHl+4uqzefl9mOLrhFt0CWzVojmcYJ
mcV1PMZyGxgheQRjYyA+uePk4TTxKpR955KkNqgJad+8OuMcm+1ZQ2nA4ZqLOTNXWHw9HawT1DKQ
BlYbCFji8SCDjHxbLu4G+5UAHH3wrzDDwMjBtGSctjInK8Nx0XP1ThSin5KzS08p6Cr7eOyCaJqv
4rCqDG7etov2x9IqLRzneGql8nR/BjgXrase/jHOR46cNSKrw0tKS+Byuc4fFFvhdEuOgQDLqP2h
vau8BVEcjgaB5fER4UzUnbPBl4oqxj3FyaVQ91E2P7y86bAtO2DQ/ml8VyW2IN0mQMOUH5lOQOsP
erkLePjlgN3TEpb8TjuKOTe2LNVJ2M1zvDu4Cv/U3ZQAm9jpLye1XRrv8egvipaJzlR1HB67+Gum
W/igGNOgxEHySYHi7avlCw0pYQFNTSOuqZw3pqgcQ3XbOAAoZGCOe/tzWGtwniZP4M9EVvYE2bmP
qrwsWbGLZ8QOhvFKvmVgVJkKuF8n1jznm5D8aGWEjmhwSonDsenOQOOyFi49PP8ytWugWuCHmFof
AjGmIhRDk5bhzrUcqLHPvg8J0E+35VCv58BW+/SIY9abhhs8Zb4c9L5Adf6F34H8uOWb7fenOjiF
MIs2v/SLZgXB9SqvWuPcJCfZtUvLCc/976pjlC96WjkZyewVfDelk2XvAg+qz11mxRXG19FPGnZY
oiB/Xo8LbPghoIorp2u3YdFoASNmrHnisf3kU9tSfEyy3DHv+Qy//tQ5jyl+w/roA2b0lJZ+keKB
JSe1PJtP41Ni5HN5bKPOJ+/Q43MIEDvHTpgscJJv3Q3z6OoSN3luuZpQeTj5JBaK9w6TlTuIjCa3
uTRLNCPd2jeeeqLAg3HD2tMG/PUWLWq1o4sEvUS0sdOpdSsZnJu8Bs+fceWeAvW0eFGEtKlJ5CBG
gVfG+dz7S5K3IObUKI+34i+gcibrIxZUdG7XXBJwOH9f50PnJ8gC7PBxeJEOCL9wHGKlt3afpu0V
GiirrVlwOjtAzU5ePVfv4fjE1Gm230DBYO7Q4JW9MGcg0orglrA6h8ScdEA+zlljOWRxhdyoXuk/
diq2gxu6/mCqhoN43RKAfohXzxXLukS907Ar7uA+is73gHPzTF5Q+LYX/rbeyY0BcK4TqpCq7FBD
GKtCS6y9UN3tdwOIAJbablzSNnfCjeQGrfvORcEEz8SnAMnRiC8n4LyHwzFWaX53kMkc6174ZQ+e
N2RjKSGoGzGiFH/XxnpZHSycS4UAEzW9B/+oSQxxenVAVIK/S3iXWVecATQBTz2MCjmfqjQCV0Kh
YY9PU0kARcDJlLk2gFc3+IZER/+rjlVKny8dmmTIE7gcnnfOhAUvM+ApNB6QxtyIhswmXyfdEwZR
IFu1JVWHHe+aA+X1Gi2KCtj4AZjhMrgMiPMYBrvrmwX19JJgyKru0O/N2GJ6aPq1NNzTVJWwAawJ
rssQxy6uYLyBzaLziP+P/0kdXiL8y+ZvmOtOtcrBlK4G4xyveIK86lUatpd0HyNzppwRwFNgQ3fT
xKH8o9yGIkL9q50ZzDavh7CUX2UG9gGzn+39C0BwYeST++5NXKQU7iIAf1OC2Jl71Z3WBaH1VwzD
ugUFlXA6WK9gCJD3/TV3cJbjVS7MjdQ0ku7yjdFNd42W3Bh9xrdARSbwqyVROsQIEISPw1JUNP3l
DK/lISFK+8VPAY17f4LCfp+/3afS2bE1XGgO7eAah4f7ReCMoeWNRRRLof7I/LNvTrOR09NF77Ik
GHdJRZx2tqTaaqVnQvsHMVGN2JierrWvBrpc17F5eYC2RNGahUAu07w0TcVRIUSNUxOzATjiIgkJ
Kh64wpjJlzJgo0VI71eo9Nf9BGThR0iee2+gwHUzPu+FodB7hKE/fyhUNHkEKEmFpjXZFlBr032u
jhxLBJPX1Tj1DJMsQlP8zm14p6xOg0ztSOshuImavrS9Fk/lBrvvcZuARFrLMNUaecuI1+uzxP9S
LxFlK4Sa+FjK+0X7UJ34KwmtqlemKgONHROD5jVAI5D6F3TuV/9wqUL1yaE5tPKCSj9xLqzuDfKt
VmROP3xpptkMOgm+36Wmr0Cghx4mYiZ5qqtaJIX/J4yfy4miJMwfUFBqLuE8yqdCZ5ND82Kkzl2k
4CAi8loNdE0CPhgZ+TlRASTHw4ioqCirgI1S2XMAgvTvPrqj5ULivNfu8pdRLLVnuAM+gSq0ERHA
7Ck+djci3ecOvFOBk0cK29umqkDbbjiXDbYf212Dv7KO1cBIWP33Cks0399HwJEw/Ie/lOyUgIXU
oeQ4SYTJylHpYNloYBim419pDQz2T4nkRX3Cbf029+YnAN+F9s5cY4qELuWFfJPY43JCJfugCVC0
PEULnMj0Q7EO2Lg1WR33xFKtNZfJZBpVXAusnWj1PTOt5ojyfBw2FxwLfNFVSv9k1dTndvQsUWCy
B2KbOGBafc9PBDutvsho//35OgddZeuxZObwrqv646gRZ0nLzMOF9kNExg72pl7QjR5qLJ6kMvOH
bj5NcMbu9m93/4HUajMU9zsh0f5g/+qpe/75TNTI6L4EHId8LzO6rKA3Q453E1DK70IBbLXYxvUU
7wECZ99Ioa09epbSh7G4ZuWCIzOh5p7tgBh8N+ITwQWDT8VXwiDBmQSZKBN2yGDhaiKIZ+g/np3I
fQCD+QsHROfyoMBCDtIkFQ7KeOvn6qVyOJwy/xfwazLsegMb9kDvaN9EevFPuwwB3NtqL1fI9Jfk
/eUcMU0pm37vHtB/b7vfTqqmvnDEmtEFgG+dv/cnWHcbVtvL4JpaIMr7bcElnmoHUeHK2SiQj/gk
w4DhsirQNXQ24oIMtuZtxWdR3fIaHedBjjJOuvMJJiv1yf5g9tV01FmAPZMpWEkKKldNGI8p0eOs
8+/ngdyf0B0QcuCDkNe/ceoWBYSMyK/Vd8UHr5nZAoPTIkmbqdddXhvbO6C8pP+JnSRk1s0bzFqw
col/5lA3ejNcNlGC8CKah8v8VJQuaBpcYh2NU334/kv3kvLUrvjK+wqIpDVTN0+KispTD5EU3d6z
3qQaFhkvK6ZqBv47QKjSemYojz4pUjEgfQeLLryoheewRnDvy08hesUOr8MtXi+LsndZXFyF0Kwi
u0Pz+cGQwj+W45WMzYSbF/QivZzEx4uvbVU8gaSoyH4FQch+FX+HY9i6vixsBZ0bgwx3Pvn7K03K
SIQYcb6QecHA7CvNXPMma483klrx25+KDPlMUMhBTlNuWSCwiI28TNNQoKwDWZ5fSajBWByneaBo
p4LAGrkAu4lCy18PIRtAf6jX72z3QcuHGHjyv1FV/bIK1z3ONJGE3/27AlnvpeAF/xvn32D4RsPj
d5A1IoEoybyiS3X7g9bgT7VahQaCcHsc1A1WKZ6Uebzfq95YoroTLvJQ3ZfHM4rijxRYqdhsbJim
Vz5XGzeQcC9YDat3TXolQuTjeAxEWcC83zIabyBqrByATgHmWuJoIIiQ1rknJqDnNLyBjg9A0qZq
WtwIaLtclc3b3+IOTKrXnl6VZ5eQhqrebvQotGb5+CH89ROVtg3DfcM6TaXQHQBahi1BwMiO6qvh
6V6HzGTxuZB8knhR9W5f/fXc8VFywOfBUd+q19LaYYsgGGUY/fjZ+8djP1EY6lrgddtFeHUV/k96
jQkcFf7FDyEdF83RCC3BMFZprNy2WgciyuM+tUjpbKwTiIq8j0qderRLMKLzpaRZYVHVM9uoHlw7
LfIORNloiuQVd/Oxqk3hR0OIA59Zp5PPUmABRg/WE5bFbiahUfsEDS1G6Oax5vuuYxc0cJ0MmIzG
Cp9dh6YaXhmaNO+JipSE/xf5jwKny8qtmyJ0zqlGrgW9rgl4hm9ceBxMuGP3FnH52ZfecBFg3cfb
j+C8um5T+Twq+JwYjBCCh+yrDWBbjcPtQ4dbsalvZS4q7bxUkf7AeoQ1Eh4PXnBy/tXi3qgeTPDI
oP+JzMLZQeHYQ0NzA90LWF32g9w9y7Yl9dmfNhIk0eI4U2YyaP7glaSjM+G2FoI77TaYgMt91piH
TGVcTW0DBYl+y9jsHM/4WqPI5dn3N7wivmZ2h9jC3QqcFyjbdTaJ4Tz0papOfyyFm3bYE3ehpmIN
K5iU8m2wBWNQhv7AFv0ZRvYZgIrp8Y9wKIYMZl/LXHp+Ei+5V6r2dDMcXw0pzDmndvSQ4aG+7I2T
JvlVd66/q+MWx78lXCbMDHtV7SbVgzkxU8rK4r03JuqlhTqjDXur/FPRhhjCElWQA0droDpdSrHt
RhTCy5w7O7O33UFWc3Wc2zQsAAAudUgqeN8xB5y2/6cksTXnXcueysaHY2SJyRWdnTxpXTWCSjD2
oM0ydyvbzoYFbSueAxDYmO327Eknv6PWyzAEEo+oq0n4Hl4IrKt1nGPcZapk4FsTt4HfNRsWAPVa
ssG8JQYkmPKUkR0pCXNGXGCDPRNJ2KpjUGrvgkVLh9Gl+kDvrB6gnQ2XzIk5ZGL8AihP8uj/rlY6
Mq3jUjTZQIGEpqHs5glb7AGq9ON0nYYB5JgAv2IBB+SVygm+HnsEqg++IimdAbSoYj5wr44p8e4G
QP+iBW2fDy0RDPpPMB9T94AReZ1jXNuXAVg9xqLwtsRTj70upLIxQSPcFGGofy+bZs6YFjW6nkWv
YFAinQVDNhPkXr3bmp2imXcAjOEqICmKqT+OqxEOJW20/HQ8hA8OHvxCe8vKrR2hXLsXJQ+i9FDX
eL7MWz0Y4HtnyPFy0MBvCqALiGOV7PTwAKVLJ/RhsQR8o7lYD7sf9CmKXhu4L6tvKzZ7nm+HzTJI
c2OrPLghRrgxNb7TsYN1K31sykiCHXiEJqQc5psf+I1XDli4PIj1ko3Y3CzY1YDYlJ8zfnnS3ED2
g96wXKLq1EMzbD3GQiGoh4/0yPoaSrlqvt4Fb/FH/tRuFUdvVDD8C6FaP4NyUeNIS5dPfx9L/d56
/VsjzzVikpSd0MmfJ/hPtb/ME6+U8GOi0+jjleDaAKoX4nN8wBbtv9aUcy9+ThsCALPkN8mml9/h
6dtMdDlSKwhIK5nRbTBHPfHKMG9rS90LnpqesHGSglj8YfTDzo/GCQT2HGKzt9r/D9uyeKphQFp2
FEyxxXVBsxd2Q6p5tydC3qR3w0eTxg+I7tzGxCa8VNaafZRUFlQbtvz6AKzX0ck3AHxcuJf5oTbd
cBzT17npitY2jdYd3jRAbIn1I2g9Xdnl+LQiA03uz5Gq4SGghdDg5FSet0t4+UAgCDUSd5eeimV7
Xyv2aSsMykOBct9g6yxY3GipSCZBGD6i9zOAugP19LrE1jGwoZ1Zy7MDPU9VpRSxJSZh3uIbsmp1
xNeDlPoiNS8+E/KRQ2g49UbABlgFCzAAmnEU+CjF39f5LHlbyjF70CmucMcSWXHZap6QqMT8ZcZx
Qzh7+huWr7AfJRBfGqnVB1/tqHttTlPEyEFbuu+L64tN0/NEZ3ah2dGGOy8+qgmkgnPet+j7jOTb
x9fOXm7MQ326s3baskjb73NOG0eBMvYIWxjbk9/QS2zx13t4RWDqu1hTSgbJJ0a77vxp8K7Qqrm0
uwIJlbG0WRB7YpursQzwms0SQDVf2UqpANzzOjhxUDuM//eGCf+JVwVTe4zMhJhWzPxGoCohwupd
0dp4vPeuBV0bQ9nfH49lD9qChoZGoTdkKmTdDHRFwNBAci6fJEwsl1ptSkMQgD0llhE4BXG69/Tv
K4LXt5fr1edlGgxuoDJ4HZd1SpVAYp5Ipf8bnbFVTECa+zD6lpfngOZ7bRspRd1PWLTYWTPu7JLA
qEUX8j5Iss3jFWgGd2IBg+A5P/xVKqlpS9k1BB0h+567vDZecfbh9xchFUXCaVyce3kbyyf8KTFm
Cc+IPk5mPBXh3h03Ju9jGikdq1+IABklJCY+eC5CLA+IIb3OdrCovtrhidSBUSf6gDNNsNYOf+zl
0NOsGzratbyUOOt3hTZM9VYWE8fs7OWyy8vvJX1rXjPrzP0Xk7gq0hFH12euGcxCWQaw0Cv1EeU8
jhU1oCG6/IoEMToFePx8rccMc0Ftj6Xqato4yzU9aWKchBJe+NXUB+nijXYbC1p2Jk0hpTjRUWnv
Mvrri+r20tZ9nXmJ1r8wS8MpI+MB0j/fUf7gUBPbbfcvgLDoM7XiAtQ4GcxOIPRQXqy4ZDfIRhRT
DwxEZT0gfylizoqCTDiU35LXWTkXeMLWhSZgJOOLNyPgKghidTqq0IXsHCtuuN0SFu3tb+u71PHI
NMOZR++1LyXVNsDFiMKhKvR2BlS1kxqgaMZBo/9iRr10b+X3tb/gntw6bIKk6fICeKGdrYPj1tRi
SMgLPVILtsGWR/u7O5UjwLWTXRqSn50fTf2i8mrP3Yx/15UP4q9ZfWvWBc/z7bmoQuBQNmv62I3r
Q/TuRVrbpoPd9hJnS2W5romXDsc7yjZ6ITpss63OdZNKnI626Pqq7OuKWoPBI6vzPbVQmt9GqBiC
moZLt1oQv+3BGZBU1ESphrcpgbAyGHt5SMAvjrSFDC9/LYo/6xVJEh3T+JyTVG1n7qpTiLtdBsYo
DZagtcyiRRmYX/RrrlDsZEFGKgZWuWFF6On5ZF7f/OQb+anNr4qz3X0AGHOjheEMQXLdE/XfAD2J
d5vIW1LJ36r64ESAE4SAnxrkrQ2oLgW+jcE/6l/70zMJP0YdoV6jiDR6SVqt0OY6OaiFagP9tUp3
o3ItnmgzVk1nZnSyckAXbkHZw7Hksl0qYgL33VyM7g78V5P5SaqovT5TN/nVtOF5saxmLiDwa2Hn
65m+riLsgY8g20lKECOyEfJTSsoo1sD2RthLIrhQuvpaHTtugLqWVqpv0wRAn3RqnMDa3ojhzLsq
NQVYA/X6GA6Gso7tOHalTo19/5LliwB3REzduxPbef/Pvk8bwjpsT2KzbwHndTRPid+NbkG6OVFO
nuPTfaCtiVf9GbO2TXEOkZpO8habq9lfJsh0NOtCZW+Ah05VImJLe8b4IkYGyzeQzp57rdULjqwG
NxSBpRY59yUjtmqCHtbj/LpnqUQEuBMXC9PQiCYlI7ANULBxZbAq4GkHkgZrOu+SUYaJqlybWiDm
kghQuXZW7HXuQvsIxFt4zydc9vM6sBn8Fv/Gx5Se9wscRfGxyUL/UhM2SqNypcamjG6UqFQBD3WK
T9AGqdkGx1hAkzlZ58QwCywZn40J6AtYYsYqLMtwjZnkrbF2L2yaejGGhLMmYpC422OMDUvOqA5Z
69GD1Jko7VNCLn5uO1WQ9xAwLbpcLjIY0onyKTtvloca0b/dfP3D7Nl9sAbUY9tWAuUaiuwca2dB
uMKFsBf30SAvUNI5qMZ20XiyZqj67sEMOIoZ7IaM3OwV09hqwQmrkqvJNzVebSBFLB8I8L43J+Zt
P2+TgIjswgAnNcIuCuXx7zYZlFiB8uDbDi3QB61nYTfu+NyPKqFdojIHl2HvDnaM97WQSaPvjA+8
BV0psX8PtlGQczSol+VnJ1Jx002pxAdyIwccoy0/BXssIQE6hyy1wdAhVbZ0J5JNrEYXDkrh8J1A
DElwxwnFK1PfVo+mslLkGOXLsAZlo4tp29ayhuQIXVzjMliXgkqt7RpqdKisik0CxwAfUq9QfJj2
iowX+PVsg9AEOB81mPkOjqzJNp7MywNiQV+wR9HThe+zin9P5nKr7uLRiuQEANHt0EwME3oGULCI
jVLf36HfSB0Vuoo7tbYwmxlpLeeVK/USFM31cbSeyG+4Ewm2V5vVrarOUvljrjKTB9sZLu2RpkP6
b65/tYbkSNswvEou/S15jngLnKwKKLWdT1D7LQPjSbOPgHmLGPMJS7zPUu5OuwftDdFBNsBuOzTK
QqC3ULJx0mEG/q1jEFzYR2xKDDDH8sL3J7MHuAFbcwiepqFQtZK+USzBULH5cQz5Oj94HcIKlHFY
kJyed5HOdQhTLQz7qiCtS5xef3i5omObHByeWji8aQkoQbWgXOq7Cxb0+MEFroWmN2Qvz+dpX0cR
FSiAPx7KhQ25ng1g3FsmJVa32RgDIxSOmKJlmWm2Gjwn1lOb5goHhTZXvxl0wRGOPAGBE0kbu4Bn
01c2sjo3/JhGarlhvXHrLpTiq5dvjqSIbubLQtgLMTbjaySXb7v3cchj7cUYx0r5MBP7SExoTX8r
Iq+AzU4H1muPwVkgCT/DGaDE3DLyKOYOfMx5uSOu5CGPiV0KCSNutnB1lXUmA0eZtLwDA2IvxuPg
Jb+lnkXNkXYQZF/3z+waZtS1O+uljMbdlRO3o6merKmzwjjYZVzLxz1y4RTvb8m1CwzEbGgju00O
G8VYfAtuc/RtcdQiRJ/VCi0=
`protect end_protected
