--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Qkb772FZ4PigmIEp/tLKTup6UsFVx538NyTEtEJFd2xyYyjj98MOPhcqZWii9nSTaIhAVfPUxu+a
Sl/ZMqjLCHpiAFfZLD2kj1n+6pZaysWTfwue5DwPLaSqoAt7kI69KDq3zzxiyRTP0ficPIPQXDpj
5PdyK4wd9XsaJ2MoNwZUf+1uwM/HG5QWQfA50V6KnSdOwPnYC0jkKFHQJuwWNCYHIP4vLZAJsRPJ
mpGVNaB1nHT5cTVTqMGOtGh1M+EErQCbaZkGltuk3ODVR84xd1vCBeIVa4jUXN2XQwPXAs3NzbFD
izK2MLP6znBNjbDZODJBc3YlbUy4Cf32T5g2iA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="p/TLh5t2uDJCVfOhRHkkb1jTh0t5QRlZ1TcNzpN/oWU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
bquTET5KbmOIvHeoFyy+HVtbg6FbXct4eciASgSDW3IluBgc7I3UMHdgk/MtsCtez04h7juu9CmK
BUsBlQUvP5BtafC8bAvtPvQoQ0lgVlxyrPVLDmFO5gBNh3nBphTt9QvHMv2k4fDbM8XFpfQ1B6v2
dEnkr5v8UM4xZuedC82UIGHmwvj1kU/M/9gAK3c1vHohx4H+7qf5/PCtWBuU91Ocr/JKAjr8h8QI
B9D6VMUQUQzR97NBhLC/exZk/Y7u3dXCOgI0GzeVnqVOP2BxCLdxe7cfH34wqPIyI+8QIpzcP3/U
D8uPXq6vBGcMI8Mz6MBU3Ris5ot6x0YxuxbJ7g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="TabGXTtzWWjYanHSJZz2gaYTMPIq79A4656caZnN1Bs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2576)
`protect data_block
Y41ClKvfOf63tmLzWpp1DyaaQeNGerMPpRwDjbPnbl7oDbKfIuCgEFmQgiAqGxrhXgeIsCDbXYPA
5+XiUoN3UymQgF0/2coDXO9GXrTnzVle+kL+yd7uVlbDLauWyKjHuAi/JESjeFnmscX3wohi6G6g
sQ0bIv/SRj3914SPstgmkOwTbT91WoVjzwWAaaOzuLxcFGQHPZ5KnLSkSiIplIv/vnbgyARy9VPb
nlfKdgNFyCOKh7lu0g1Urwhar+Sc+J4UUIcLnBMug8C7I2YPXrmbo38tHJ+CvRM5v6Xsx93Y5bm8
tBtSt6GiMTr1Vfbz8TOyjREfB0K4yxaaF14sY/hn5dmcJ07jPRr3Jx5iQmBEAyTlEUj459Tethbi
3E0AhBy/bzsCxC1uywXiUi24yQ1Wy9en5Y6Awh0x2Vdtq7liwT0ThAQ3twPtGA/a5gzry2lUYRVf
RWgH9hQQSKH+25+tJfQBo3oiVnNWKap61Urkj4TW77hWt+4ssccUqgAhvfLTR7aYQa6Iyb+QOqwE
u3kqinDqJMDfj/52ubbRuzRuKCcQRYtsm8p12k0kBRQ/vOhqIH5BlcMUyTACLztsS/KHG4OsiGwn
Ma0SgKlCtU+7+H3sqPWgSa8TZa0AcfHOZwR8//VpXSFE0Ps+M/IYWcTSLT2vXH/ANmYp1tvHXSpD
Aqh6UfADBorxLwB9VcDf2aBSw8jzDv0fKjpfNoKpr2F4yn5CXjhvJcHosrl2wEzqJkDliQnqKRni
uGQNHu8BppBbFKB+mXnPmHnjh9RrEMCzw/26UmysHOGGTpCafBezFpXmLm1dsLck2K8xBwtvbKY5
DaemUM+EYSerrXjlS0fQSOeqG0lqiY+htvHkCqrbiSe9FocS+G3n6hCek4i58pfT67NLfx+PuLSN
MeZpwpK8PgIEmGWAXKcqxB9oIpenytsEexIMezXy/j08/VJFXXiKfsNFO63lUw5TEnOgqpXVjVYs
ZWTuy1//X8RIby7zILTRGoYqtqK6a2U6KPrKm4hRT3BANUcffyj/rOQk3yxkp9vf3lXVaoxOUdFZ
yaaoAmc8N4SYK3hEswTRbySYx9q/wbLJ2G2sNt1Ffmk5SG0q3ec38QSno3M0xWJHcxoI3Hl2T+9o
03UR7v36aDBCCEK5x/Knqt6kjat/rtTOVToerRDKHD9xfyQ5jEULcfTYFTQL3igkgVPcR0iUrAU7
E168IAtc0XWAFf2lKUWR3UCP/5oBH2G6z6DRMgAug/R/EylqQZWB/083yxk0atcIyi82JoN9mWQn
5x/IqERVHLnF73E6CDCPvpVJ3mc4lfFIxFuqgCskMW2WMS+DHLADWSvPTno5KhQco5WPsAlGBhXo
lhF6BcWb/0JJMcH3ObEcbGWANV3osU16rpSMK+PTRlRvXPnMWneSHLiUIsojJlmG4rMbZq09ndU6
WpLOniKbKv08sAJR9appJwRiknt7gO+t1J2cMLEwXNx6naKoSIYgLVQFs0LnQzpcjhhtrA3l3pVo
1upU7IIRNKv73J+LD2dzyJTm9Ua/g7C9Vdy2LIHupVInkgfZ/HcIwY7Kycf8zKAkEGz/Dq5u1EFg
CAn3lHj/Q1MRvjj/4vu334mvKL6IQ2AnABA+qxVS/XpNLVtZRk8bYDhxYCwXNmc2EA4iO7XkhDft
4swLaH2IVu0QxbL1PqKJgaOrZEGTXUJ/jjPcal80Jr5DI2Z71gjeB3ewRb7DsIswWE6ztBUiJkWz
W19sUfKOu86KtZ6xJ0lb9YQQROgDwvSyBl4ftsj/08XDvgUvDCOLUQjVmC4kQ50LgwGcMoINkB6X
WcIA2w7g/Cgmsou0UkFR26wlgA5dqiCK2PevvlQzwStknGW7XWLleFhMssri+UloFqgMexb+e4lH
vBQRw/o2rCxahHIPxUcQegMVjLT4M7qLBwy8YezFgMPtAoL9otrLpxBMjIn9Pn4Qf3XAHEzZSxCQ
2vCYZG35jkXi+NuXH/5AXNSM5oT5v7b+4CEf0pqdWTKIMzVsxc6xRZ1gOfF6gi8MLuG8OSIfZdXb
c0DpHKfVMckghd/fN/8D+9idez7dhCdGiSMHXTmdGmHhq5vBPIQGE349qQnscoqeF5/XYr4IyzDX
UyYzS9bRuS/ciKEUS90B0ipddmsofAT8Y5Lz05ASLw/723grATLkcbR5LJBEYsyQHFjnGWQOzJpW
J7q24JKjaA4fRjqHlK3Ljd822K0TbeFPWBdUgeM3ZufaOtSBdty/Jyv3TJ0B3N5zf7/5zHAWa2wm
S4cSkSIYGZRfjDbmCsVj6DgcStGuN/0Yrxv/xmUPh+wxpeES9Hq14x1aIFttrO4jVPBrDLlQBWc5
nNFAsD4iMXJSub9/QPCWuwpiyIQRvvZ32DOepi6VfSKilfWzp2zNKsuMx5b3K1loM9/pahZUkayb
zBsGWBiegsAu7ivENl2WVHBN1Lo/tuZ9XDA9VlUtj97Z8tcnapPjoG7ZOpGiJxaBh3A6c9fLnHgL
M2umJ3sOWiameB3T3zUoEZquBbjiv4xOYhoPVnwQQys8ZzwNA1n3lS6+G9vcMMs55+k6oILZf8oH
2aUH8ZuDGsF9sgkTK3OMhCc6hOq9IDTFiZ/wm6DenEJdYCaLOMj0uG5ZOkti6gM41Uk62h7R+L45
vh3Z3vLEJCCIkeCDbWPmmbFPJIECnnxCvEilS/c1+c8VVStDbS+qzWBVVcsj3yjwMg8uxFrGOPcW
6B8PWNFQC2hVfnGCLkdf1hoXmU5TH2VBC1TGkBHQ96lDBo8HfsEMyspi1w5CMU+apbDLoDy0iH2n
PGoXZtF78qC8UkLsS3msRdl1K22+02pbFCF8jIbPkp4zC8kGofLZv3BCpbKXmnvSUz+Vo43mwNhz
ivGEwbgKcQmJSHVwzAurlk7IoF6s6DwqTzShbNxfg5pmlI6DgWUfs2spBO0l8MuCUmewhaNJqW6r
raRY8jDwH4HHUllUiZkNTOpXj38bDZWHEux2kT0zFkIvTyqUokoWXPUQUB7qpxtdhc9sVB9Vzysa
gsqL8mo2If4yqvoevnD8fJLvVIosgJQpLP9IwPTqn7Bx/1bopkL1NcpPm4LYfQx70DWov3Jqi/H+
M4FmeiCEczAQP3qrYmPhy/ohanq63I9CwAWbkTNZZUFrwMXUSEGWCqbcWXieDTPdMU7xfywxNCCO
MiUNfxWzP9Fic+kwz3UvmG1l1R4tVQz0bAJm1T0Kk9GFt5Qbsh6DXIcOgEgt/YFs9B+A98Fdk+hL
uLHukDF9CHxiK5W7YylMsOBey+3h2PQt0NaEe/T6tJpLFoDHU5xwIgmIwAefMVIsPQWS73qFvvW1
CnjcgTLpqKsIoQb/ubrSYtswJWzouAYKN0f9BpyN8P5epi6TfCYlH9tBqb7gSyTWpHl2RINTaf5r
u9/EYjS6g3yeHvE=
`protect end_protected
