--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
NKfFd4pVf0v38MWE+cf82scL3dGc2lOEqw1kDpVaLN7XGQhJzT2Xlj26rBqz7Y69oqrhfgZv7XBA
s7Oq3RV5EXcNI2eC1jDDwPttWP+xmaIffqzJ4PeoMQRxzTJgJerZdHkTjfNLpYdyJe21cCFsoN+Q
4pA3pbFs4Vb3rg5j0P3K24gqwcmjkW4H57ClWS7TmoHorea19gAhZSmm6nro8F0cJo0cV1b35BF1
vxBG64dKlK8lzBmfMetZSVwb6IQDmziPADCRZ6BaLYrzxTxkPCylCFxygIbGwqbZnMzBIHob7GVt
FJuQ9+LgZXH3UiBtmaM5GL6jy8+KN/VG/EmGsA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="EoPko+ueljm+kdUrySBF3lSBKg5GVMQWaOlKZTwSqx0="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
DQdeZHjBrFQsZayARiM8OrfAbkAEiLBauIKVPuyoYElO0j/A46UzB0KBCj3EU3mBb5dtrKlmPF+S
AOK5xsRLntI4DXNnqKNRYjE36CzEX7ve4KlfZdj1XaNlhBeoWyouTuXExXvsUdLFRC01Cr7cuaFG
V5eRLgZfL4u3sAK8+4G8pRlldTbtuURxgBinZROt1otMRriTngKCxtFJPvR3ddAt+RzjFc9Vr9fU
eLf9ccfzMUIf8WR8koFN9XX39g5ih6BwyRNwui5YODUGa88DI0l37KEmxDsAtHqwDGtqY34doiKr
wqpbhl1G7BIz/f9eUK0dXX2XAALEit7l15w6Hg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="jf1tFcDms+lp/XGiKtGIsX4fOecWLbbKg7/TRB5Zlrw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2640)
`protect data_block
tgco4prokXZkNT6hTTLRYAKbRbUkT50mPJCgiFlNRFkmwmxHk/6md66HSLXsSr4xY+F7vuiHR5UE
fvou26YU9BKZ7ADPJV+C4duoDRKrT/ZASQ5aT4GlDpuYmJ+0ZAQLVdFg9i4FJSa5CgRLKNDwzxFH
XSNrdkWVCJOcIxyOkVud5eBI1Th03Sdr7Oq+n8eNGT3Qw5/POs3QlZoIYVkAI/+VJWJwflhjdTB6
dIWFEBXTNv3nm/5jZUT5gcSnF6kh4fn6+TwGcoe3wSnMQE1tICdEhk5ACbwdoQa+l19+dcxckqWw
RP3bi4sYQ9gsiLvjgN3npt97pnoJ2R5WqDmnLMGOePIhj36GpsvWaLUHAJMzKMF+JlTVq33YXWGD
9p8bfwtLVvRMUEiBZnMBo3aU2uX4nfHa6lD1+2qFnRsku2atwizoWKpEcZ1zOoXjk3iqATYhS65Z
gMELZNrBHFPvJXhXsKT+pyQ6TfswdeaNymfE7CR5k6g9e2s2LXjdGCBvFagov2SvIuBMFlZv4P7h
CaEgdtod7MS5ecOGg9VpTgCNsocFtfaDQhK0/Pcu/II0IY0ByniSAZaXAvsdXQcuALylUvk7vDTv
LDt+0sxmXJzYt8DPbhOL7msVnAkNrPoMPcMSXbebGsqynE+25uAljd1cUdQ4zn0M7cxRJN1omYT5
XRllV1wiWfCnyynV8C2GKzVkX0/f6+WPVnsp6vGU5Xft2B9a/6vHjq5cg55f++0It6rrE7QpO0L5
bwQtomswP1DAfVrkgETa4eQZ17nzv4EwHw0xxQT1MzLizNjuLJzLmJc2lS/L4E4RWIsAiTA1N2pk
ggfCapQxGMTXRSAIVc4VmTR3lOsdqlUKLugDLSn8xvwIahIO1Q/wZrv8vZvsXrpM3KbRV6nLrNOI
F6Vz32/wL6/4Tib3Wxidnsm1GkWx4ecK18Mg9uX1AVD2kyVVUVxxQUwT5eGAzGXH6a/an2lNbtFy
wKKNpJV2pxLsirBbN3sJ4+Vb2S+XkrJYIORGclRmmWJqyWHVnuAVnkqV5FKApkus/jOfrWlrmUNa
SKwJNMnE1oVq9OiPUaIhjJOJfAfi2F6dIzJLlHhNhPmkE68NariRPyrnCBh0zFND+jTrWdT+Hmqj
80hsnv7xoLlcNh63XQ6O5EYXd6II2rjkeApTdeZ1F5nH0glSnypgMz/FWK8kcU26WOa2xzltoPEU
q1FH3/zaBevQJxFIR89TMaNr4mmFEdLW3TXibPx5bOME6IRJl8NAZwdwgLBvCdhaCMWPXrH0MsxB
brJP36Ku2deWCPA5IfXyEJIv+aUuRnPu5QqrNll3ugJJ881Jk9xnyNf4ynGu2erbu//B4TPGY22u
O3m3SqMcNVktVklSaovpsph2lG5/QsKXM1zJEgGeP3DCdc+9XsshMlVc+Ie8bXACoSb/sP65Cat3
fIcjkeedph4rQpw6ez7jLDlNc24gRHxKjdxo7fhL3edvF6cJwJoLXZ0J8MHVCeP6H1EdxJVydzF4
QjkLY38KMC1GJ2acTo4wCb1fc71JnJkzk7ThvPBKriyYjS1ns3a/vf0hQwJSeC0oM+gyLl3fZgQ+
6WiCrVETJqeNFK5ZiyrIwJasqkMj2sE5Wz9uY3Oe12jCE+QTIOivd2pp+zbJgxzeB+ErRIpUT4GW
uIxt7m0GwO8+8ccWPViT1504u+9vJmWwnDNpIFyLDK/Fl3vi+5s/nCna4yHGuTEwyK3R6zDQsZrb
KVh0q4MVFEvHLAFOVU1fLX+KceIirYpibQv5qjbYFwe3ViUWiFWnn1iurSF9NgmzBakKijQrWlEw
s212jns/GOE2DH1VfU1/KWN6/CEU9fzHELb6gRsmsOa6PFRGoeNPXymx8y7iFb2LR3uI0zdhCGrq
J9dJkaq45NEeP2MuxTa+f0mgc/YIqWCdHcmLVQoOWcXlF2I6pkKZmOX/h0SjXJtMKgHb9Viprm6f
VDOUDCDRQa9wygkN3R4SJuEODAQD7jE/hG7CxiTb7ZPJHDPLxbWhV9s9tmlIDpwf030CO+GEi7V1
EdOXurhnTLFQufubVx4jhfuw1wgk3KBk8E8o+UZxzORsfxuACg0s5Om/44D3P2w5VvnBeGeHgNL9
7rH9455LVcMF3HdJiJL5pAZOzMPG+cEtJ0IKcWZvLq2zrRcc6KlHTlSJLtEmOyyTWVLSstpgcAla
xlCKaI2JnyNedklgwTu4iK/u3gbRK0NRZwtfI2kNLad7GrJkqdaq3kzS3H8Lk1+sX6QA0K9Satz7
MLXGfkhiBGFLJjSa9UaWNZd1EME7X9XButcQ96RemGzXoovokH/n8HlqF0P/3Kuj/SNmU53LBFgx
xWcLAPAGOyto2dIDc0BFzfxtW/q5Hpzux6NUAg2jVYRkLTRFIgT5VfjiXIGejtDVW11lYPNWg+is
jYzf8PFZsvF/zY1QmOW0gBCwy4rp/aBkpaBg3fB+5jQVqub6YM5MQpMwvOFZVFtO1xBUaz/XjU2Q
Po0KZxp0oLy6i0DOSLCIqDCTmUY6rQkCiER7GxnPJBJNmJCI0Km6TPUpp1Vx50+P5OtyGmhkDFyW
S17Dj9lXGCPti4ZiF7St093+tVCBaxw9JdimVF7MOxa8POODaDO78zLjnPjNBNt7uLYgu8qBqsxU
13Ilcc0EqloZDYGF71GbuUzpmPmza1Qn5Qie3Rzu5OlzKe0D77SNcFbJ+WNiPheHsqBu1j0wPN5O
sEZew2JJPwbky/HsCtQS3aNtADaxcwJwgohpxShTbQhtSNbRXj1ZZcWBGtJaUY4Ojr/WrltUjBrC
UM6D3lR3+evzsFWrFS2xU/R9vy6OZo1X9E9Uyjx1vzCo/WqO+y8BJ+svCvfn7UnifTg2K66oWtEX
UWrr0mC+2TrglC46wZkIRGMPblBBiZVdzuCiL0yvYQjX0IXA2GkoUtpHW0Kyp/DEX+vXAiSFD6Ag
wyi7nyUEP3VjGnSIwkq4544xji1CCLC4U9ff1mwIRPOLUfYcY/dVdTmlYQaFhopg9cpubLhhL/Kq
Ism/hTQdC/8WmyV44yDl5XNg/Cl0TS7So85HGs35dojX7lDPQbeV1gxcWKtTJ4YLT2yD8wKIJDDK
V97YZGn3ohHUnR9pPwrlC2+v/0jmyZopAsvIpU5DjEdfqRwDC6ovYxPmJVZG7eD+vBabvtvPCFWJ
eDxvRyT/JQs0JwBxuRC8MYgpnMELf1K85KcBNJ+bHk8gzdc/Qaoao52+fWgUTvkgmXl5hY2gixCK
JGTxVZ44ui5SAm89MsNHI60oSMiw+t0hVMkJRvxAF4arIjsijfP13F+Rcvhbsviqe3gqqPFCxoVa
GOycyWLAxDn348iU4xK00l6nD1/LShjo7skrwpznDmraL9Jx+HxKzC/xjsg2T4eIGDCUi3gOBjYF
RRo9gREtYcZxoQj/dFiwLPcuB/7Dn+SlM7MsAkciPiZnRcLlIdcujpD91uJwmHzjyeiKf/8mS896
koUdoRl5siIjhBEh2RS3ShU4
`protect end_protected
