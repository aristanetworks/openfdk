--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
iXW65v4O6JfPCFHQn0amNF7UlmAV34o9eD6KS+M70Yb4P9RQr3dHI3/GEpywJ6R6ss8Ty9MTyi/o
enSUXImu/b2BHsTIyj9Qqj5jCDTVp5E/DcCACYKDx+q3aNhnbfU5ohZu5AydIMzUnZF0gw2zmTJv
9ERyVnM/JDjCOSz3mQDMtd0/5IZQwp7KilRKlDUL0WGbhg3cv2Wf35EtnUngTlyfP3rt5bKHL0Kk
bYznkELe1vLmiImfWv9+cVvuo1jACj6dedSM9kRhFIdT0iZIwo+HMBfKzPTQwBMqg1oHMS+m1uDP
BsVc08t0CaOcKAZUmEKIrYfsmNTkYqOIpBtPLw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="UXxnJLi+6iz52Zik6U6m8zrCPoYd8ub7ShF0XwqGsT4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
dmZCQlmjmE07iux1RpNBT3W8v5fnyu4nA5jHcOc1BoCFj90knc5OXUiz9H9yT5VlOx7ikUPXAKxA
W2Frp1NwXiO7bKlcCIKTNcuewb8gzNXyhbZTrmUqv6p/XNpf051gziuweSQLN6cOkYS9HNm2D9m5
Lw+cIELLtC7BhybCuDo72zWPpm3Zua6GkMIM7xYna5NCQQ3S4jmzARWyRHS2CROkUx8sQN4BKC4n
BL9ye7mPX16EVUyDQRA5yH+NIWLqnkcUqAYyf6ayhWlzIofGosH4hLspqhoFaXr9R++i+hllebcR
LzonsYfUD+LcZ42HdE7yjqBeZzURNXV1xxraMg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="50gxVl7FHm8jtR/JF6rKi4e4KidXuXVlfv0waXKH5dw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2512)
`protect data_block
XDJ0YBVqWe4a2Ga+G3B66BK+0JN2J889n5idKcTogMyIxEyFT+/qo/DRMpHreaysdwkwo+4DPwtz
2eXUBUBxI5uy4JKtqOaEEDDyfPqUPY4le3DO2nBl3hO/g+L66BZPRgeNRk3YmYX7FfnOBRlSlzGm
dcU3zFTwl2fuET5MbrWdUSls3yXtpJcwc9CvrE1CWvbAkB2SEzD8a4OTx0bj9tpftQrHcFQ1lAIX
E8mEyjPuZPSCKsKgUCST8uDUL0mB8/i7LAEtPXgDl6M1W/p1A5Ly3evEgD7a1Urg+eWojjK4J1Mj
eKfdJV2lxezV7NyzBFgZsh7TIOYNhPUnTtuyPLWBG94WfGNpmMn9tM+Wm/QI5EUDFPxe0FPuG6gb
RYp1b3lSmmCXfv7FM6f8kYIzOA8ZzhlhUmXJDlrr0y3dbgkKdde3QveFBbkJs6pnXr+UzKvwVSri
YuJ+x/bmKsmcxIM+hGkTuedYTlQY2Mjn57HKRGGpwBpr0H79E4bLrkT0843lo/KDnTzn+nH4035i
fKL7sESd6SleVLtI3hnoICtdhfiUWhqnQscsTO3S6QwjQ0VOXUlk1eDMBMskBBXw5FeYtn90Kvi4
ZLBUsyMjbULxNDng1YeK39mgzP6EVwZzniqmYN+x0jklojSuh1KoU8hWOHm/qgq8XQn0zemU54tG
cJYQLH8vBWzPwr7PsxYop/RWs5pdE9u/cfuLBlBNiEsjQK7To+CCERiC8RJU+LlwIsX1Tk8L/Ytq
XW55hnqjxC4xKNJAgUMnIiYB0UUHpZ0sgqPlAfpAzabZrBwSIfxAyYVF7JevyvWPPuxKJevKSl6C
fD7omGHYJaK39UDYDIXc22pRicCzWTIMi5ZO02KLhtqrgpa2k2d+LPPbv0v6Wn8mVuTuFXXeMiBk
ErIKYEjJOfPzNKf9VHYdQWWkPxtr1/OIZ5exqi/DSkTV9NEyeFkaaXNR0f3p8kRpFvVk2ua74smT
NAG3ltQne3xwm2x54UzrPTCgurEWy0+0IIQlqWL6UAKwAS8l7SsnG+chITclqjyiQ3TZUxKX7Qyp
ZV6wX3mlmtsdLs42kTS4f5Tp6vqL2STfBv0LblssCWTH8bxGvCQzGVED/aX0LfQkIhlOUcbSnctV
/m9d1rgMlqrni8ynivrDgSc6AmNgbTx2N2MsnX8ez72try1CoIB7biDgVN0qlBmN9hHrbYXpIM8i
UtAxli4yHZSatNNbwTfr1+2MY4EC/sVA3f5eo/2+sKimGRvJ+pQtymea19N531UOO9ioYF4jyLso
7twefbFvwnA3QyfDK74WQvKrc7vO9LqjJooNsgR+Eh7piHbcTroZv0b1A3VjZcM141B3aXQmI+l/
XM7dUw1h1PmTXPaBa5X98p3YZihOTnLdynz9UInozDroS7586P7nd44HECfnV4vzQP43tT/aJXhe
kP6d2/BCrhS0rsBVI1gXhx5PY0hUvwqjhFgcUDZ7V1i10VdbIUTNR187LlUEj5Wp1NEewmCiOaJ6
w+UmLA7wapro6Scx3WAr4wZFCp8B6hrHZVswS1F48tcBL/Z+EU+maqENUKVMXs6CMt7CjqyGyPff
Dr0ptQRv0jGgF9F9E5KUTK4GyDlT5WpfcCUg4fjh1eO6MnvFOwoH5Ol/Gg2fPvLif1sv13Wsa1oN
LJb93AkZs0GOAgx/0w+9pOMOyrMD7jkq37prSGIYterSaRen/uIcPbUKOHLcYahOVNCSNQ5eemgH
Fhk9F4LbIEyB6h7PWfmRCbYdpgjkRjCkAArZVtrd+AZsGCHP272hW9g+0LlD/VEkFnrPDKCtk+Mt
sn72v411YKkRwmHH9Q2YFcLY8QBcTvosgWXQUk1m/PnQdcZ//d0E6MI2PnVPO7NAXNUxFAlaKWha
TpQz3HJTZ4w1nE+0XrkGpsOh4u0CyfIsdEkZu/jaZJTXL8v/4NR4kf+NbuO5ZbwVF46//xCxActz
dz1OdBXTj9DMNwmrqXKru5Fo7MvQzwX5pJDhypA7ZmpNFMyW70bW3m+L31uF8BXiQGXkUNSfQrrr
fEaW8GEOu4h27IUw2luBy8HMwVa3/TuLn3xMjaLsIkvQ57EIx9DJgde+RqY2DhhAPOEWLOiZ5DnQ
jkxL0rfA5URcudwNQ5T75UzROCvoZ0LVJlTty4Ojvo5Ijl8NsvEWcrrutAe+u5Q8I66XNBayShP0
ZbEv9simC4Q3/NAlBUlhXmu5rxI7aj0HT1Pv5UL9gQPOKDQXJXjqaJuswIq1+mbLhaQyQDSTB4A6
OlZag4Bh7+oco+88Viq4A7tZwj65FolXDl6GihfKY09aQxd7gFxbiYdUtYNaB2fgZ83AH+vfZKku
OJ+SDGtdShVl1NnUxcnvuSMdjCP9UOb1KQXfqc8Cfco43S7b/WL28QqyTl3nvQIvBsfN88/+eYml
erV3tIEPy9HQPcSbSGIfhJOvUdfWX/MqqIRLG7sgVOpsPUIRsy0tyCkUrPvXjA3IEo4uZFfn97OH
A+BHmhipz/jwfS+ao/o1U9eKN0EMDXFyHi9e46YORUgVVfDT/S89m1fNv4d/QcRHuVea77EuBP2X
HAlxwJHus111udsN8O01YV3Lxg78JMXvFHq7t4+04Spd/kzLdZXaFcv51G4xpCbl3HtQXp5pH+uW
WqZijEuFNH0W39sJK45Ech+RO7w9W13CWkFrxaTpA0SfUAkEZ2VgUBvySHgCqZeI74vgobcHdwnP
2dEQ1ro7rG8M6xfVdp8kH/cyky2u2LtcYeU1vhxCtGkvWj4fyKK65vaD1ba/cclK/nDnC8nYDiWR
1N4qJ/FJMPAs6o0I8BTOtoS4mHkY33eQtT7vbWx3WjRjVM5qvXYSWb8lMvmlCxYI7YTCGEZ+SFK2
jaKuMS7zn54fSpfv0JyGVDEmgqqS+s7125l433ZTms5awbE0kyWHcdLSBp6U2lsBdotTQbxUGLvD
JO9xlB1NfEgzgs2hwHApIbkdKzoxib4snqthZONqpST8yXFWMqbX+nTujSuK7k/3bhd9XhzeKI9k
5OcyNErQzxHrDgxhFKXh231oKI56+1xtcYmzTyeC29qKK9ZQuTY+zAROC6jNU3UOAg8RGENA4GCT
EO0/RLEh0lxICzBN2SvwvMLCmOegrchD6A6QiKnSPv4kjTjtA7DcBn2BUv0aVubO5ZCYCjkkBOZo
cQdjisd/xnlJSSxt7i9YYzT20ME9pZcf8Rf3kU3Q/kTUdKsTIPXiGy/7CDSPmCqZyrsj+n9b5omQ
eW7RDu9N7m3WT/D9xHqU0Hb0VJLvUYqTGihj6kOvYURL8Ia8Zryvru79BJ8GfdkuI7HxkxLHZS/S
tzjJcQ==
`protect end_protected
