--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
hycNucYAEgnfeHYx/KrUe+iSuTVXZItx8OZYMaLNm/ydO7qtr/ghuDFA/EY9Yqrcxze9LmV364xv
cbYhuP2caSOuRWBO5FMxA5KB3JuhqkMIcxF7mt8BtGe9j4Yj6Ttfx35BJP4iThs3gwJQ15Qn3MpL
xMlSe14emb1BCjXFkxkerh5ychfH5ZnL90uVx3WvCSwqGF9uSgNVAdXr8TmCbpjwSM5Bqd+Y1AVc
RZk49cF+ZNJXVpvQow7bbrDVctB6RwQhqY2kmsJj4Q3fEiOPNeQaI9U7PIOUBYdVu7+McwD3a+xz
gH3dJGP+r08m1q2QgSxBv55zEt9gf63nHXvbUA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="dd8xHtq8igKsQ2NvdxPRIiCiUjZUT0jAuIrUf/KFFJU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
scEmfEP1+bu+7P/uMoIz7u9GtkJ7erSV/6wAmMJu6Zk7wjxSwWCRYBxIwAhu3B97+LsCg1Be/sCa
Zu8+dBWecABNi2DGzVhRJd9sZmVaGSe0bBluW+G8GzKvp4un5ZnfMp71obNmfnRiMtrk+MZNzvvT
uyALAJQhtrb+HhmUSbS4fKEZwnkEYZEKZuIxwTVJlqM6xWugacP9zoR/4+Qj7vo9eevae+QONoy1
R4pQJW9Cks9Tx5utQM0LnfV5LFk4QrfFP183LpaDzQ7Ej4JK/iRTynwNjuSirdWzx+1fUL9fcNfd
r+J9OUh+382HEo1C6nVUNHaexnS889yRaCSE7g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="kRPtBvarhGxZ9HfMThe9uwoT2KnE45vNOShfRoPJMts="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15504)
`protect data_block
62wQjah7MISSsW3S4Zr2rs2t4875czohI0/z9WT0K41V03fxipGUU1j63s6ornRrPwWZma7Cr9c7
R1WIS+ES/ypPohumOAtzcW3VWYrf16brTU8dmejoNfumtFKAsXTqXlXkhAVhrVjPoUWq86MKlz7H
2WWiUa+BEz/Im1++zfxAHgphPQJy7M76PqhGS5SpQsVhoLIWi4OFz312IxO03Xi8laNaKJvsHGfH
gD0JslOAC6kt2n7PKolGR/QjmHREugJloREr1Zo0KP3BnD4HmNMtcPQ+t62Yjp167s34hJA0atj9
mwALWpjfR0UjjiGn1SAvpdOwkx+118OaGJ+wdzsDlMeiWHmVQwOrM1yx1IJgEXc8LUvvQLDCdP0C
rezFnh9Yn/c0fktkRsCYHnsqL24ZOyxXfHe9Jy/AB9DXmBMtP3LRPs/4v3z6mQtuJvjsGVpt39gM
Waunbaic9brOePDyGalUUicW5MnyuXYGoQ8AyOus5HYqXZ6KsDnp/gCG0oksvhbok+bMMK0PZtef
S08H1yEdLis2rPBaGSTPiJctYphwqplqQsetnHOze2gZjOOR1NsEFpsQZnU/aRB9ooSIw8j1TJaP
VLS6uSNvbp500zSxvcjhznBgQsb4md4mKW3ZdUQdUlLsGvpt5PYv71Lt18bYbFlgBiqGv7DYbmSX
yaQjwGxjFJo75gNTUUF2D254Dxuu7LQozD/OS5Fe0DH/Mm21KIKQefnJ6wgm6YywNJKj9Fhy5tjC
bOZJV4LHx1/6BJluL7LDYLhty/1cKEa6O4SzCwbg7fmuVuQ1kj1z+CWN91MNMxSq5Kwq63ID6FHx
vgDpzfHEi3OCLdAam4hkGRCKyfHtN2uj8caX34RCm2NhK4cvJCv+7Ad8hprr2NYpfG6uKLxfApLC
qgjK1UeYGnE6QTfLEfnU/ude2/joRKA+lSMkF7iXg9R1BFo3nEXI5YF3zVL3q8R1etndhNZQSsHE
xlLLBCGuLauq4QXAUFzucnFeDC7rocVjvbQz0RZRsZ4VArJGEmxBtpM108+IJidU0JgxqqnPJyZ0
6oa009NuVfTmwN1iaQ8cMyGNQhW8S7C/IrmWz/69xdJFAIemydy7KS4lsLSEXOW5JDL7nvjFA4FT
O46jXmsDzMk9BqCaS7eX/aNsMmFp/t06IXvC0yucaHBL/3mAMwQP3iTYUoZYq+w+27KhNaNMQsAR
+r8kuaBkolwb3o2FQaJ57RPsjVxzlJ39wZO8E/apoq/1HQZz0YMNgKKXPSeML8cQESFdtTygpBQV
XtZScXAbpbiiQeS4gxworOatgSfK1MWSaSrG3fdv01iUsgl0WkyanhUGFEDg0Sm0VA0yHJegfqUb
aqBOV8V7ZR6fJ3WGQ2BlZhllBV5P0ZaZWKS37fQSF8s8XvuhMFmMxzPKs5ahAlDcJQj+Blgal0Y5
KKWTs5FqrsgG8X63ayvMGGLVlgn0tzMk4tpZN1+QL568PZ2cusS8frem+ZCgwwAiElw6dUArfHbi
/YjEKx4Vf2Pv9feBjqfQBvdk9ws4nj7FiGqT2WF4P8gV0EkYAeGa2zjNC5VhC0wjgO3D5tnzGV1F
c/vqp01mWn1e/sEPhzJBxxPO2uVeOz3mu2Wr9XKttP3GDhG1gfE9QJFfYp0bobekzoCiBLtAZUCJ
KiWQrmacnTqM9oQaopeHjySVVt1L0SzP/vR3gsTqdjvYf6AHUP+KxrGK1QQBnJj0aaChP5z1NsLu
UzNJNH3L1d1oknEEJMM4lZ9BWZf1kLqVCXWYZswjQCNFWFisqNFuCKle2yDSu0RdMlcBgErYM4O/
y3mBZt1famPb/RvaS3yzK76UlCKssZRo4iOtF35MWc1yebynW4CDl5xU1vitGpeXcDMVY8qoed6F
gkd6xnupVP2kVZSQBaFD072XglSeXcQU4bvy0LKruRYp5LJTnGW6S2lcvRKNEJY7Rvtn6tWEGsnT
IAuFgnE+GGfg8g25cVediuU5E88KNUmqPcQyN0M/1mAS1Z0TtnMPLJc+cipvd7yrYXw9hos86kSv
PxRU9fMLQ7MHPhIx5v5KuKSwp51GXGuaq5gx2yWBGMg4PErMe9Xz++Xdo/efEQwdGIIh4Lp8HVh4
eheiS+ddZSTCrM1wSOL6lIfoh4ljvvmZvarhm1bClb0DC4/fupq3EZ5wcoVltTaTf6aMPvQ6J16J
4d2Ldu2W+xzEwsmQyqdF5PCyR+s7CPENHuC/RNC4RiYEzd+cqgp/TnvBQBIwJg6yI4BP6O5AjPwV
l12yuKcKXHcFW4ahzZ7c6Ew9hCB8Xar/ly8kO0pWCWOvJJ8fKR+YZp5h6UuZRdD+/siAj0Zs213W
MOoRCJTfGPsWN+kVg1NVCI88BIHrJ1x+UbeGCGMmiB7FNgMjU58YzxAk26kPKrSLbEXwwKE3fX+W
RoR/34fJbxm6nLlcJjNHhVi7500SETM1xMd4iR1OCanSXAS+uEfaSxnEuTm46HdBOY3I/fcxj3SO
a+yKdxIY2VkIMZJdHnFQK8jCMHnZP+X78A2jR/GXpGDkpiQhASx3sBFDaqqya49dTPVEEdIbvSs7
eIT7b3LQm+4Dg2tPBAPnyrUNWKRyKV8ok0LE8Q/61ZZ65fa6MVD9gv74ONyoYtUqBVQ1NpHpGvHT
qZHRYHn5TaxI5jPCcGeIkTs4jgY2wKSlHs/cRgcETJoBShq48VNhzTvjmDCoRTRxgAuxCB064mj5
/a+j+7pg8haUD+A8ZzY7pVcYsQKevRy/uee2lWRvf1NTWqxXRSoe4YfVfA7tu1VJl9IjF4Yv9Ocl
CH+CSaN1+q3BX0ZleGpPMHvaFfR4Bn2PkkxZSplTAgIes6AWsJq8khuoRuhFNDNIAmTlM20Yq1RL
bt3KzAxnVFb0EDFgyAMQIl4AcpdxctplXXeMkxmMBvksWrXHfmFCTtd4LFMt7k/aXwYDCzTYtvY/
Jopan3hn6jDPxYxLhFvpRgqPfvKfibLyEU/0rc11xApap5vLrIAb8B78Iokf5apYWkz+7JoTM3i/
ayPJbpACDOMMEFnSwzBdLqjhAMq17WmnS9vyu3UnNfS05uBTsyOUNuY/LWOH1ABVj295kaQX2Zoc
TZxDlfxtC8z+sO2vUwomryCZgu5VTtbg446NstbXQtEItdQYt048R8O7ryWWkUtIhyZQ7tL/G6RA
Joi9vRgt5jlZ3pco5+LR2KQ88PSfEJRnzzVvISzFTGu7J+1fky7jXtroKMm+MvuqA5tSs3sU1lyV
RWiXwC/OeAF/D+oDHBeqiArArmjNBH5maCeu1lSuVQTvC4e0FLeCMPaCG5TW+P4ZKwxzq5sPWwsc
cvBjgsnYlAPD/eT8NloWFOWr9FDiHVi0p+hOJguwNFi1jM3MeHDgNhlKcy5TxT/Y0FAuooOqR9y8
KvfyuCDUB/wtJzpZY1asBglZmdcxXSeU/gABcU9Dp5QsvLqx/F33CuFYB5Ifqy+MEgbPUplYztX/
0oe7RmVO2VKY5sf3y+7rfk4biQ5SWmZjA/UmkCsaRbs2EdYJVZnnfK7trzMwQTROKZyx3Ybu+7f/
gY4a9Kg7BaN5j8ebCptNdz5dO69RzslbrCzp9sgAKxENQ3ei5zJ3yxmRzop6VPsb5LoCa2JGAo5K
E+rQvMvy+vLmiy+KvgLRyNVx+7/szfzj4HMO1EakXCN1KfbvYEvygbX+7WSU5nNyIT8MSSU4VdDe
oC0l8l4hgsPZyB0GH6mvJM/unGhUPkmJyWyq1PsxJDP5XGDh+I9/5q6Zr1gAVxdMBRVcQLxEuq6m
BDHjaTE/8BtCtuTSWnCa8NmTEtBsWK4K2g045slklRrb3kIKMGNUQB07y1WQp0mi/YGDj9JKy+EL
gjQyGBb0ZKVRKTuE15ZfmwWWomo+7EAwsMmLIzDCU450EDUriHmuATn1mVMi3tpDxqtJr7L63ZrO
quGKO0cEZQCjuYoQhdmwfLMI28G5SNMzPuLLhXtz9qJBsmBcUuzuIL0f0IAG073PmFZXtobYe39s
l8H9EEv4QKvIUu0Mxtl/a8lDKw6ei2aNTaQplBfb9LxleHH19C1+g4Y4MefNivbpJMzoKdGpNyrA
tUshc6+VbbFD89aiYLEDjHj3kwXZE/kGNkp0Orxgrq9PSQl58lFL5vcGOIF51eiCEGhka0JfDYZZ
R+jJthpKr6rCT/nWXvKajZ1jHoDCP4fHPWVwfBY5ws1kC5RYBjbh8Diw/Ifwd6zmI30a02aypZJd
gyMocsRKyMRIkz8UT1U8Bhbf/F0b9VTgFBHzKHQLWJFGiKZaDDUignqNq+09cLQb222Gct271DcB
fGoAljcyu2xOJPIICr0Q0GErUoMeom+4UBKyVeYM1U5s0hrEKgURpyPJ3PFl6PDP/ZJS5koCos3h
EMaYMIqCfaAw+VmrKRLXgZa+mI/pjsQnYPe/0JW4cveFhe75vxTvwyh3hGzQe8597NQIlfIiDLT7
6Dg73mb2ERaLKlGkNC3bbfrVcSdR7BEBX3HPFFcx+yps/E47zjGHGJUVt6y7v9YOJSFYEXh3zH/I
YyXHk6SiTvHpWAuO6OiDdK6AGe9KL0eHH4OLeL/VJGE9l/rmx4ZYAiJOEduFM8cHqqnGna5rcdcL
NynLjP2GmNPiBWYq9jo3w2L7+nujK6cBliDxnOvWbatEBC/BhQ0mxJtd8quF1MTHq77ja7DG2ciE
das8ZyLKhO4oNtypSpc93zelLvEB6lYvIrT39hZPx7INdGY297V/1178PRqSmokzd2q1DKi/dAIX
KaZokQFmk20Pes+Ekc2e4XbGp4OBMXAVOtWfhWh5M4WMn5nHqQbNgxdqNSShDzktjDvwewHC8jdM
5j02KSZ4D3FLS6AaiJO3HmTA0udTKTDIshEvO6S/3mOJzAGW8G7APXW1rl15rewhCBPqJuw3HMFi
kzXI8qW75dK9nSuVx5aBw/NpFAwOjsBVweVOH3vazbYvcz+xvwuXJkgWbxpqJrkNBXqvLFMGTjFC
i4W0+EZdljq9ovxuj21P2wW/LcN6pjmbvRuLwk5urfrlx/P8TTBxylcepC12betTNj/G0laBlyZS
C3FMoT7+BSDnPAZD8sO2SA9suniDe/nq/wsRkMxewOtxm2e23La8PcrQ9v67O6eEh6hBoKXphiV3
T2jQhebu9hCz3PInLPJvKbeczoeZb52bDLG5SWwj3qZfW1lTrdVKz+F1QvYV73Padrsq1NO5S276
GqJ3aS6EylPvWI6SNVdPKRZK/KLcUuLSW2iwHVilvO+h4zNmeSVUIgET7jMyoY09aRgE9xwZ6KuX
Hx0BpC2B/2iwgbwuHmFpZm8b1PVi1DL/mxuPCdyhOFaKDPFmAokLbKURjOFN2DNW2xYzTRp5a3+Y
+U8ay0y15cGKeo/uKVINRK/eTmAONh6c0syngHrm0T9O1C9LUDr4qOFZCd3+vfdsF3HtQOn1AT3q
ZGp62QvYZi5+IhfQg6Fz3VufjuL2sQBcU7Jw0ArHiib6Fd28CNfZ60j75Iveza1Sz0j+mIREDedE
4TdcTWPUj1NtbyNBUUluJtvBbZz4BTtYNFv81RMrDiU3QV0mxheaLhrgLOv0SvUdjtXAyGrpvsgh
PLMDQMzPrA9E+aRZu2PSKctw0w8t56DNjjPQs+beQF+UNJ9hIc58npFk2s4Z9u+jhsJciujju16j
bRJ6tEpaaRUDV9ByMQ8iup/XfCILcaVZXufg74cLIbR2zyZ805zeNDf/y6rCooKUaAJt52pDQO/4
urDQiUqOGSkF/O0JVv8XR6xLPqosfI9qoShNsIpqLKCK5dig8ZsmpWY0uwG5OCaYjMt2cHWGP6BI
yQExhqK3CQBdf0OZ9AjvCU4C27CjrxuBmGvLy77t+MmfbLt/qFtYQ5yd0sckoFjSWeZ0yOynEOM0
RSxalHB/FRF2woT/fZP73bHi23PBeMPnyWxgwuCLCebpfnUD1iyXSM/H2GjjF9qbV99TuOVKNpxj
J55vWU7naM+Ety6kzn/76wr/vcelVDxVSFVuGFX9qRq57eb74o2Up6ZE2yeCSclPiE16Kruij6IO
F6Or3Vsn6kSRK7dQU/+Ku59X2eSEGfcoP1C0bLdkhJKYiiQBXoDoXH1syDQK009eIOS+yJS12oAY
+bex5Xzq+0pwz8fE0qEm34xEGBOYMpUAwp+mIjSaQ0CzetRM2valBo3i7EZsrOjsN98AC5zgerXE
A+aP8tTuP9E308QRcdoT75A/VJIFaQI/MIPOyd/FbVpv8TsPNcUZy+vSsr9r5OPphCU5Vw+j65hV
YlHQ8wWQYnO568dPi6AKNY/ns4e9n5iRCXoGjkBeN8eglQ0A42oEr3A6kcwjcEIdN93CqWviiy9f
lNGK5h4NDZUILC1mGc1lBcWkeCInLWOZQOwjKQusRrdqvjLg2ZMWe1t+cFBgGLNUmSV2ItSpisM1
BsPkePfWJeqPwakFAGezxFR/y6AWSw70ZlJpyf06IW4rkkGWBKG7NMz6zm8bdkU80cPoyStQMCxn
CVglyBBI7P1f2uAC/ZexEMaRwxE/Yv5m7OuGAgMTfBQJYArb4NuOm04wLICifg3u1/8CdevkoHuP
3m4Pl8HxXjhczEICYTC+GBaWEpLRgQvi7IuE+9N32KuHsuzsAnz6bKrtBPfT7NFKav1x8m4UGb52
AbqKWdjhYzYOfcYFaElHoKkGSMBxkHH44Rn0hHwl2fcg6bW1YwJ4EoyIOXIlGlr3nD6nRNh1cEIG
x+gIYKB+EENrWs1IqA9FGAVWaFI4c/a8CHtm/fzCboZcsUsv6uTYwXn7AwSYIM/+lgJf6wURGf/u
CxqLuZOhbu9WzFuuluqT7mxt+5Bttt1UvXLHxzIM1m0ICzxvh55NngGtE4ljNVIpKlurVonCXH3q
DNiI3zQlL2ygL0S+IY7wZFeauxs65K3Z+wH7XPQrZ3NXSiXmFsbaYuGQOCxSNC72WTFFrWLKzNO9
zTpaQ5ohuBq/fSqVqD8RMbAVxbQTGKJxT168srJDKudtsBE1zwJjPD7rPqQAixyyJTEWyrMssdhX
IYtXall09Pv5JNUy+auuo9bi7xkvTi1BIWdNeCnf6sqXAr81dY6XSE0wR9D9iRiNe8iLZWTcrPAo
5MKf4CbWGtsupF+8Xfj6ZQcpb+6OLsVYBXX6OFFNrycTOZrUnVutEsqTe/s1Wz0tdDhHTePHUG/c
+iq2ea2gbO2GKq0u6ph+Mwt53Yz23++bikCcvqHHN9mYvrXItj6bb+OlSvd1WIgPk+Pkpx28AAry
GabDm/sFIU1LqTjD0EDQOrtayqNnRG9CPaVoqkcyUQWiarBBMwUbJWqpY2EDDsJs74MpZHWaggny
ID5lf+7/W8NJRNMGObCh2eseuAxcm2Whq47zCkMUbL/zslJMcoceJVhAhkBiQxnsI4muNuw684UU
AQgBCHBiFeyYK3bDHDVJLlYKGaPBjOfsqNefV153ACjkrmcSmTUYUlFcvBFwINLlhFF6OgQ2U8WC
wv/1m8XeT07XENpx0KDBguVGrsV60iHUbnsj2vXVRbVWe/J7c/k8gI/fdCDon4Ef09TG/IIoRXro
4pdKOsR1MMCRGYPrb4nHw83n/wPVHtZUki2em9tHTVC8Q5IgrBfU0muIfAub6YwJwr+H5rlztyxw
yuxf9bG1Pq9mw4abUDHNanyItfA5Y6H6Npt9DwLpgMpzRgj0ThwbKUt+SXgZ+KL2wvmZsIHMZMuo
sOg1gqb5bsTJ1n9UMcWKww2Do/54+M8p+bCUkQ4kz04tADS5Vf89fOdTg7a5AMRUm60Uk6UOdwoH
YB50HSkjrqVb3W8EzSRn/0PGPx5u/rAEeyxmpZcZpDojydkboqYGRVefEmskCtc89fBCa5ew7JW5
6drXXxsGwm/qT7UboHjfbw1YGrpfZemkx3bbm0+aFd1yMBqZIz/RrKGK970F9G6YQf/ktQK3Rm/k
nT0dpbAxLZIVV4V+7nujqhR2+vf6w4NdpzUlyw6nwb5GpOIHc9mDKYqyAoQPs+FLsXrZA/tXT4nM
i6PFQxSp/qJXoYvBBQIBOKVoPu7qRC1Cm1nsw3FO9FZirF5+hwOz6alsAaigYaZ08Dh00kM7PoPE
wdpTDPzuHt6bM/3rpWXqgAEEibpfG4ujp0oJXO1fqRRwPTyIN4MPuiOxQgmrD6Co+vM5R8B1p3zs
KIXXRiLFS4ZEmyTqU+gbWDf+jpEqUOgqkdFbQZLNDRJLG520mNzOWPHGqYZv29t5BJebEUfaj5Ys
ynDgisd3XeGTXhAzltXw8kBpFu8dWsvpVnn2Pmr7Z7Lu6qVZaqpAmEUYj9SnsPNv08l6cciz77uV
+3udTPPO67CZQu9wLRQioA+x8zaFo3a3VnFlYB/TBAfORGarswTNHhsDG1ykoofRQYbQiS1c3PPU
Q7MNGnzuLZRGcpXv67sdSfu2vScBwd1eEttqVOip4WGpK9wxbilOZ5XZ0z69U7Iy45CKvsTJHGLV
m8P3/RmhoPeJJbiY6a11wvKLx/BGsB1OMs40qRbWwBrbeatk8ZQFAuvg1e26yopRfe4DDFO0YSw6
3mvjfZQMXpeMIGoEo696BrBmj2/T3FtGPCEaFqG919sfsCApekVw+4j7yaAdgK5JUQSGJvq2zA4/
fhibzN2xq9anV8QdQzMCKXr+wrrqmjK2vSNo4H5Y7JQWMeu9Qhe6hwf/S60zRrWZONeT6jH0YMG7
a+GuRGmS2Ig+0xbrDQAEDUlF88EDFIN/gpOXmoBAxNalP12s8tGkPqsQKWzJIEaqDrMK/9O1htih
Iro51xpFElYZGvRgZTsPnbLyb+4MyIFJYosDFv2kJWbUVPJa2fupIoAn1hb+rfVYyVuFVRJ5xL//
0cNFGBr4HoQ8Nk5a78kZ1tTlRSrR5WC1O56HaEAD210Ig23qRGqbnJdQqcMK/eVxwnpzAcgzSaKn
h5YoEAelWA8bMSdG5CnL9pXz02rxgcr8iPgAA/XxzCcTsBxesIQxHVV6ET1NwVzZ7SfFB1zZ8KCh
PgP/0dlmM1kXYKZFv/dfsup2Znn/NWQkwetZlmbtsTI5ivnWz0QybfKt/725jweGpyY/nfJCAKW1
fwIAt00f/dnBJ+wmK/OHbXlz7n2nftvC7kKgCn53Zs4URpL8Wb3EIXPItX9AcA2lSDki64T4bSaB
g74OQ0ibFKf//J608Mjd52ZcMJoniBpZUGwPTjxe/Gzg4GGr2dUnbMWzi2RC4cBNqIdVgNzwps9y
EQ0pxy+pKcY+bguhnM/Z9rbp0f9ssvlvxwfqvqkTnM9RjuIQwCLuhIcOBPkJ6Fy+oGSmGzpckepT
RgEc+GOixDlFtwWy3vxzW23v6DVFsh/r+RWJXc4BtTlgGCDEAyLk1V60ZX8c2FFV3vaFG26jQ7ec
i26D65bd0nXQ8Jsc/X5cD9bxiPmgklrbDL0DiYax8aNPDTBLsGeo4MToMQd0OKJbGpbELK4lfhEW
W+MPdIFeOJTnjAbQfFTAcjoHJyTy8VIf9bNCMIvS8S3cWQw2frUNvpVVrap8JzpE8iA3xVC60f+h
fHbamakuzP0mfLCwAVsuiFHwLG05Ixs90PHE+hJOsiFqNcqz1Cf/hIBs+QFMOi4qMQ6AI3mdD92c
TuCvQk/Ao33d4GpYUTo6GgtH74fCP8GrCrpg18uLn/7g9D0+L49PEe+5aG6jdXU2GLFMr1UXuCs2
wYtG0cdm9yikxBZon/30IhKjqlssA5F35x3BEfSuKAL3fnPsLQcKkE/Wzve7UEyfO1erpRmm5bFI
rYrevI1V7vnQbObaEpuVXkM3WGy7X2dUgKznsVGBVqYN8UgdbJqXaYdLBG3gENcohJqx/bVCxpYI
47QZ4NrjA1eSv72Wpqz4mMMCYnbAOjQs7ailsoOCucmMBCByk4EMijx6CWS/Zu187ys0MGVDQsQb
shpRy+HdCA0xTnzI/+QUhb/E4tm08nYyXYqfyhWak9tP8r4OH/ZSXh2hd2ahsiCTKEGk0kKjHkSo
apaIAWm1fmeTWU+Lfj9Knx0N5qxvOc0UskIyEiHLFJ9hBtPESxDTQtesXn8RlvFo0pWAnkI6JMgZ
D3NILeTsOZV2vbkKJ0IpdXGTpPNCtTT+1yZl96dp6hl8eOmia7cf6uD5lbb+ECaUWT/MQfbN4CI7
HVaPUIk+eWF0A1+0Qwn/zNBwxtaP0WM7wo2Gv7SwVXaxNLPBwIbl57xPlLnNdnofmXiLQ2jiIoSZ
lllmhIBiKbrwaYDlHJ0veWjjbP0N8BAsnJsILthZFgY5yqB23OmhY8hzoHSVtPbyfrshX9fwjfbI
2u5BSSfVBqQmO0NiUexcqSu5LQ3V3wsVdq+LdrYB90UORPt8CCM2D0bYeDwy/i89bHAFUaW0zOmO
G0GzPjdIi3WJsfFbd+X1XgWsWGFajZidaJ+KkWq2nkgLsXLhnFLC0Sk+UM4RX7rk1OzRp69Kbbf4
8Ye/wB9ddu6wdtb6IPAqtu2FmqHdGY++xxVqLRflorJUecxr4aulMvC1ZRg+LIv7NQsXxmylbR+y
FvKnJWFhkGynqKbbC5QDcT4tIdnfossRVBbO9aNUPj/xQHY3+cNsEMFCoFn+oPxauI6Pv/eJOpfT
8W0B6tawoeTOR43eT5Z360RIZjdjHI2tg81fYuemuWHI+Nq+l6iVorcMgtAfiYvbF9L1zg0zVKzA
SYXdwGYsgn4z89kWdk13fzWFCZkgRHpL8xbp9jfyjEGstCMGCoD7wsBUidQ6wcL9K3wC5yAboKSe
ZGT2wWpTWUOkzoAyhvSNB6JLJtBjvg6CGwnqWLtR9pGELrn5xM2WCI0dxbzGCr3qubRa5qdyqiiD
0pFa5ea+iDIv2DxHT1c+EZ1YVbCC1gfaXRYDOW3D6qiWoH33U/1w9Y3BpFiiYZjzH128x6hn0yzN
RjJWCMM8aLng31DPbrElvjPHKbgpq/UIiim6z8pL6uVyq5D0gubQFQWk22km9iMzoB6BDQ+UgiAt
B289l7TYuEgJE52+l7hp80yKEIhtXJZE+fYraSzBf52cL57d1LRUU1WsrkZdl4Xmnx17bsM1nk23
jjKAt3zgsWxRIPxf2WjGxkcApJ189vo61frdX7CDlPJxcLwGMV7JInB+VLMNwjf5JV7tsPiNBx6z
zmHaewCHFZy9aAMj0VLVA5TUoF+7D7hPkf7kDE+v4IOEV6iWdnuyyjwVwMVpEv19N5nGhXRa/MpD
GICLYTEB+mtMqUwSQeHCOixmXXMVUdYCJQPSTPqoxQyvgypuXFwaQnbb6KfzRwGn/a6vwbJK3FPE
Tzw9D6xfJGpHkMrwg190IBRFIyGRCMdRKIPMFrJAdm/UXWSXSEP9Qa+lc7JPSSqaTQ56f0ZUN8MP
21X/AtUbZpTkJQupCP/VmRyvse9RVucFdYTOUUxrh0xwdIgFxf7IGfk4huUHrwLp6wRxjdmESV7b
i1pQpwfwW8O3tPTruzuzEpsWGG7RevBe0cVHhYoSfmDqwVwbZ5KgyuNULlA9BdW9jlCPAqfb8eVP
+E6heWiC45KV1wfYFLMSNqe4jCqEmW7flvuurd5MitBJMlb36so/BGdc9lnNKvobMnHxQaAd0YEg
VsNx/po8y1HuI7X2T8lgYbjLvrqxKiSAMONhbNQSGm/3eKcwFPXEx+26izpEuk5hIrIurFUdRSP4
ieiDJCsQFcs8p4I/Y5smaIsU/HUHosDnpJ8PwXSZgiFcqDsH1dySqQ35f8/zh7YAXkXqe/OCCwg8
1LyO9ORiCaGPW4wO1XjtQXuWJtbOpcDDvjjnEV1u+/X36jbd13x39ID/5wGd8PFzxBoSbuuewqlk
w81XOtq5PVS21BFZicwrAPkSNwXoX6gyliBI9dhqixjrZTJjKBtJ9RWO1ig3Ld2jGoLdAqZWSqRh
ayQ3Q9FxjsSj3HzjRhDF9O8ByW9bkrQkvgxnZQAXXisAeQaQRHIVuGaBBzqlbqlzYmS9h3f1kDFk
uBEa5CUBnXdaazfmJkgnHPEiQN14MKg46hOVj05XuEGYq5+51+lgHWSYb6Ivs9Y486mE95laUo9n
GaLeoxp/VZNzg+qGSn7E0diSDrp2FUXM5qcDy/dQmiqf8NUTsLdYZRDWK+49p83ydVK4unKgbP24
TSXa5JQQLdDQBG6X/LNrzIZeoA9Q/bsNCWAsDaCCRT93wGtwyTE4aPeGv+qtLcDwqesy3VVCNlkR
TB+aLScDf+LXJDSUbz/amwuHqfiSZLs1oBSc13qVlb+4qoL6yqH8Y2HRWd0JwRE5GlawAYbzvIID
YHUBYguxbitoVJ8Yk0l3HGIiTfX0YJzxJmEY0q1XMpktw0hXIijYUNlHI1KFxmRcFYAMIwSGHJd2
uOkKmkkgXqd3BO0PRqFcUbmidQ3/QiWwU2d8sydohR+nfwlprsdeUGr3I52oiUdpLAfSTrj8ahES
CDDcj45slOkxbnuANwkGxn/RzOlz96TALNznAAP6+T8vSTLGuGZtpXHgN10SKiCUJIw1K9iB3VXK
TxyQHmk0FACIqxDzt0eqRBQBSfRGOw04doyTdElTMMXWPJ6CJfPjKjnEOobOiBuwqejjdoQ7pO11
3Nm+nqWf8pIn4TmygY61NYBgYfTO/ZRi0+DPO8kXmQnO9fhee9e2ALFbKyDXaDvGk+AD3rD5VhTN
zXPvaXQAGfIlPtgxR3plYZJ7fJFuK3hxLkIoYaGrhPW56HaP3k67TMTGuv/lhMos7XFu4k2y9e3I
RxXARYGWh8Dv23mblrECjn20Kb71hbCdQ0lykQCyRlUl4ZXYWBU4sXh00J7T6s7tfnZDQZNJhDxB
dCQ12e84BhQNeTmMlezgpLEd0dRuQgAetT549wdpcfy3zhQDKqe4GfXOMGsQiaFLvM44ywoGDTfh
2avG20WqmDmr0QAFLSFPoCZOo0YFl6WSmsruszhQK7hJXVka+EcQW+tOe3BZyEn01dO1N47OUSVX
bm4/hgr3cVK9B1k+DTPIN27whCYpEWCEjafyqjEAUxlRvvgIRxhBKUCxkLq3zKFLjj/JJiwHMpbS
+Tjb2pSOMsNHXxTCzTDL66OP2AV1ITdGgFjO26LAn9QhJ6qrSz70eDT9zep/wubHmni8dpbTeR45
uY47BaQxzXcsO62lTFkTh+GrkKGgxnq56pxLK5JcmHCzE+6GWHIiiNMT3vzRLBg5U3XviyPVT8zE
p9OBr1/4dR+3XB8gOBw/B3/hojd5Tu5MgdVoNnNq4El7i1IyfUgd5kRO1T+2ljZt770kIh8Q9eLo
zwWdq6nSwnniF4S55mi110EGjG4bLis0D/oPuAXFWsmeC9hXFdtwEL0dQ8XaQZ8GPQLtIXtXD0hY
69tNvrjRP0UZX6+BgDNDKa/2cK1QQTHyLT/PsTivh7oD1T9kxCNNb3/4OF9Fe44KAqbT1omkKsi7
T9zey6SeQAk9zGMu0qQ5yeuAPVChVaiDQkP7wRhql0BYV6CgDe01PZVm7ounKkzW7IYh8xaUSmK2
TilwBS2TfN3EDE5gwIerHCz4OaMeFMVhu1xUjEwXg9wAetKmgjHZ4novjOQU/dHgGCVCV9XvQegy
DiXQDLyugzLXib3Khu6douWWdUcGQyHRrPe1/8yrdqWe6BjjR0yP3KzmpAjg3dsTkgxl2kq2QZSj
3PKv+vkBzJ2fBbFnStkvZFsNdbk4tvSTUY+PaHXBmU7lYarmL2pj/s4HeAThPXZ/vtzJroz1IicF
GIM46DL8f6uXXUbsbuYWDs7SH7QLHiVP4KZwHsl/O3rFDBIi2BbfPxPybzTEEJYEX2pMHW9SXMl0
2uw1ow4JKve8UoSLYerdX4eNkp+pZ7mNV+O4EUTweNBvofc2Xqx1chCFAG2DD1S4RrWJW2qQxL6N
EAb7nwXy0otNwkCZO5pIxFPN//Ka9rttNqE9CtSyMWGYeHQBjUGLkhDWvNaoa4f2/pz4kKYCMAnU
8DcUs09HGB59rOqcIB345vzNZOB2ouyEkbyAIIYw8k7vp/LYv+XhQT40mo0kdy/gLT9iJJJthV3j
moO/MPeErp5Ckcb/CAFRMCSHmtTvtDijqPM0mZaqsrQZkEhyky6RahZLi1pxJ9iMZD1G7pYC3GL/
H0I7Di0TDx3bkOVaIFzLCR22GGmKsc1icZA8beXwZLzV9/KcOvJ/CbTjaWnIncqCTZjyjDCYN7BN
zI/2IxxPpJWBr07Haud19y+JrJio4BKXGYArLN7df5OezT/sQ/1kiz0pPRd9raY8WZJCaywdjoNU
tbipZa8zWCVKp9MZu05DxBQhdsk9iaNGGlcJXX4YwOV9zMWP9PRH/Oi3OnaKxZpi+ZhUCEZ0zVdK
x94Ghd8nPxehFwysiu90GWxnXpnu1UdCTI+SFSKBBVNIBIAK5byedTQcbIbM10iy/WzuAnpsSVeK
vhpu9b0TGYae3CvKgTcCO1yEFSrXkZcbkhOII5hI8EoVILoUFvhIs/baJ6+YQUNtSn2rQu+sog5Z
nwk+YFjAFw8R/bEV92v2mD8OiiElRYvZg0FbUeiuPlM7BEfrMdHuOJ8a6UR8FSsCHB3JYJoktEVr
iqsv6SuPJgFmWNLZ19lvPL97p6ynKYsNp5l3RLK6HglrIQrw5TdIcMK2QcvHZfU2HQ1hCTv356kB
LS+uo/1qFyWrJ32cuKMGAys3n/GHb6TR/Z3KjSVU+otd0kO6Cu9keZqf9FRwIXb74uZ5JHAaybue
qvSSNVzjTNoPx6y0q0EHexzTVKLhpWs0obvYdGhuNFvWraXkP7AYPYEYvns1R/m1v418oQ2cfFFc
BIJaOTEmMO8JFwpbi8HynrWRJ7ZAiUtiY/RocMAc41SNMvBDPwKwCscorw3mu+KZzlnxzJQcxEc/
M+TbntNhB8+Efx5yb/ByNJezaCQqdjGtxEGHNzoA68SCBjIO54hWPpUEtAoF73tZ5SUdgbHNgKsV
oc16P7Apwtbdx9dIunAE6k1kbHJ/q4VWx/z3/QgxWyXxX4ZBUMo0kQVJIum4RPIOid8QI8xXXAzY
5Ltt2jkMSAooq/BH1Z97nXFFudor3H4Kl6q6bsOs6gZQ0C8zn7wSYk0ruIr5C1LBpWAE3QiAidvG
Uj/SEOO8ExM7WhsvfAxvWkkGyILuCBBEKyAMPVYYHPRi/p9rcR2cc8e20+AmXU0tYCRMHR5YiLHy
k9W+Sws6Eav0/X2RsCZa5WhpFSkoAsk50t6lx4JcgoT6p9ycQmVd8NDTi1xtvPjYYzRHvJbF0Qlo
ZSqa/kfA0UrdfXrXY75p7nMHDQpBWn62IvlrGTF0t8Vh1jxeiBj4ueox18pzYhfZ7QCaGaOvFaDf
7PKEusrCDRMo+SUW7bp3qfuib1FjH1bjfPQDaB1uR9SYsIv8yO7kKbO/uDIc+g2fokhArdVIlfIn
RS/sKSbqala4hcKwir61F+LcabFs3xYqmsudXi8FB3Cf3wDK8IpQhmlRtAC6v4gjtAUEmgZHZFRf
zzEoyXr3lgIsCKlxJqI591UXoQnG0Sv9GjdlFheBcmeK6kz5oefrsc+s43ylKytWi5zlieVnt9Ah
ytMx3axbk1OMBdqEzG/v6QC3ivB8gTtG+WRLbJb1EtbXXQTKxjzvIo/7a6ZyE6JV6XpfZP1dWSed
HgBuaCEtEpb0m1d95CSgQBLxz950ame++hWqTEh2UVHeQOqYDmluJu0UnxDoam2hIxaJQtA8EWnA
tKzfH2tokXkYiGtRPqdlbm/oNzMb7KQpplFjOXPXuypciHoDULciI9YAYKUr5G8SN1cMRpTsRmDA
Do+MPTDyzrvEsxFeNJLni2XEUFQ6txRQxQr5eK8nzQBlHlpQxfelHI7ELxD7kbPK4nfcwGid4tzX
o8IO86UghMI/i0CfeWGOm6FmQiEEhew+SaGc2hF3xsPFO/kQ/VpFUOVVgONwQu7aK1eOGTOnE2Dr
0u8BicTxfviIRF6vahd9y6bEe4pBtRpkl8795PltQ5hUqkhIGbtwHGUq8GxCBUax8zwrdBAZaQXn
k1p+epjvStL0skY8kvCuaSutWuxn9aeGMqfpWYzAyXmEX6UQ9rUmp6hU5ZMv1uIZGyqVyyX2gP2a
7G9HoDW4/xrCx/lJoTvS9TUmmEA0EJMOunzwrbt9grIJbJI0M3Q9P4pQjbryb3MAO+PCfR3+18PT
m49arjblZP3ucQwyGgQmjCZ4jxJXBaXa4QahaNssDA7sQ7m5msuNArOLiVuC1xW+hyVrVGEh3bQT
TmqrtQAfk1TpeP1QqkT4ScGQ5IkGPRR6DcddG97YXS2038gmSXWLqylpTigHv7trik7/UZcVmPA9
+KWqgxRim2IqkRhiFS2UI1iZPSFMjuLeZWF75aKZorLwc1Ylxjgzi1R7nxwNq+Xc/kGMJzlN7YRF
Iw3mQG78CFWDyZygAwVVLiz4cYJpbUxq9/fqzZXJYhukw5cAZNbedm+WXGfbY9lOmvL4XyW1QUAa
lSKYZ6xIZjmneDZhJceMYggmT4y8Y8wIaQa9oTfovwE3p0mnvvFx0/uUDwoh8Q2ZJi7eihcSmul9
lyYUjsRAejZ+g7644mxaJ67vDGP+zGJcpyCEzTiFVDUnEjeWtoRiLmqdiLk70pp4Agc44XbrqxDl
koDDO2Y882U8i45yvjOO2KXqdR2T4BO7z4vti6hyaWTyf85zXqHO+xTMxLKlNu++NP6HSp+RuwHW
Z0j6oonJPbpeUluJq2gIiQsXGAjNHueUZXEkBbqe3gL3uZGtDM/feRd9Rv48cj2S6kNVkEwCljdQ
2mLE0JyEKBVagDmQnpDC3wBQfBNXeK2Nr2EBquOD16heRs7gJAjN9/FWEaZmdJKz/k3ft37+Rc5M
LPibKCaz+44nox520rSthszjlWtaEWrVHVq2KpTcrMgn8U4QCzpPro2qwy8POlL4sCiAhBWTJRPy
h44eEfnd3mPSe9wU36ETfNvMAjxriYSXVwMCgaZPCVcdLiDQgHtJZ9n2C2QNXTsIDraUlr6fruSW
AtbnPu8Vf9RAj2uezd86t44n7Ph9753phTSpvlbzU3TSl6KIQAz07dGlHKH62tYzQcr89NgZXkFR
4piOAewm5lnIrPsAV/pau0lixhyuMWk/52pNESlCW07BqSCVd8k9BT5OwxhFpSX9VyQW8kVBbIn+
pvKUur6bcMcliiSKXl1OLJ0hNLXQ8mv8bdU0gvaO2+dQ3VbwqHWvECZZwC7XZxMjTZ0ei1bvrfp7
iA/2r361CIR/NnQuiiUNRv5w2vXHR9MRLsr6c1fem3GJ1AYjisdASOYUqmkCobW9SkQ9AK7PDLgz
91Vn51ZH5mOKTfcM9OWLswNwstcaPmwY1zcSWwPOMJBTkete7NrefF+XBIbwJ8x3N8W5Nd1NT9Zg
fScXqJO4W/m/yrep+71XW+5BQlke8LdTKrcMqHnpgxS0CxZOjR9vg1HchUQQlf93rucSMiqrlwX8
2ykwpIUm7NcDubUh0HZoaCe4+IpaT+uulY+CfvO7JD/piXSvH8j5f/BYknP+YYHOiM9zMeZakjRx
/yuGU4dK1r4oJMktir9YPxvfQPNmYTzK3hJILRSwpepK8THur4gH0SIaAfB7/SKqA+O94C7QQO9e
fsIkEFqrAmfDCHMrjp0nIxBj+lEnR/5u5HW1R9tFv33wTAWhzaACZe4wdSO2G8h50ERxSl4gT7ND
hJB2DAi3g5/xZhDoYlqNCbkno09j225xS2PsovrqNI7BojOOqGJWLvh5LUwQCK4yu1G2LtNw/XE9
AIiq4srxhtxgVCt+E0ogW+aZn+MrRFx4qYgePic3jjSQKEE1g2xhlY2QJrC1TvaPjKTnIUCz6+U3
Z9WKYcbZyxupAOnV1wwdyC9OKE1ZnaT5zAd7YBi8BJ2xchNB9xb11l1aEq7aNy3YlKh84cucwric
Tq+YwsBjEB4ufHlu1LLf90JTRJDKlIfiVCw/zt0iBKpRf0C+C8uZWtC09+kUCYgYUi+PMNoWdXpt
DLuHGTFBChN6Ap1SGITaIS6jLPYZPJruAr/wyi0dleNadWbyzRoX513v8Hn5mYZhukDTAih/AkiU
jOnSzDiVJCnuQXz09YWbhWadWMafN36uzVNdUBGKiPLwGxE/3I6csgrSq9vd3GDgY7QvE6p8v7sG
+2BJ7pu36oEC6jPSz1e2cWCE+6xZiXfKV4llHdITvZFBGxkuyWecnwXkBGtMmojGLb2Ouk/Userl
H+L0TR8JEVOQFSL33s7WxS5wNMF6Q5InjOhmw6mEB9puBAZfTwAXWtZ8h2kZ5/fNYheEgMWNUw+D
WEN27bMxJly1CtHPkopC8mB049YEc71GLhDLYkYuPno0I0Vd9dv4WGke6gyh16oPPan2t6RY2VhF
4nP1USHcEvd0gRLIMRADzaaVsYtCd48Hg4IaSgjHdXnQTJFwd3yTCHcJZPyW+aAROeJIXkAgwbOV
Nrz+M6g1r7aFOnlroaznJTi4bgNHyWRK5MM4wRkOr0L1h1AwE7nxqkX+IAB/FVGqAsC6KH90EGmQ
dAs1j46HnhlJJMxrR7OtmFys4z/8EyDhoKixYogFqKyYWUu7uXGMetC0uEN1NZ6M8/jJ90xvqu7A
gPBSjoUgY6QiVQfk/HTcaLqAzck/nKcMTBYiU23anb6NpaHTW1vsZbAKhWgjdlUeTt2c8SP8fH56
6zl4NSDCEP07WaHYAWS88919vwmyZlgWUS0DzlF4Qwj1Yh8OvVFKKtzd4WrCyVCh+py3Ke0ndY5y
OeOx/M8C/xfTHsKRadzf63mXmTeQrSWxQb0Ow4T87xUSQ4Vb9sLmQikQt22Y6w4TpMMUdn+kqoaj
YGNOZ3ClUW32SjUfurtfpMku2v9qQmmVsmO8ygKmsOeQg6kKvf3gabJ0IsGwcApfWzEzkfxL/4Va
BmuF3tcMtys0ydQ3VxWy+jZvebfeuyazuSqdCxOD70TYDt1fVv8A8yw4oDmzvtzJ2lOpXtV+4hmP
T1+1J5uBbVql2rIdrwnBW1VdK38SC18RIAbBeOaTRoMpWayxzTpi+7YxcOWT2+nnkg1hs933Tvz7
BzJwRnbWzeh12L1cfqRZo6Osacxp0wydQueM0dVc/2WMS3O8nyghhOuSkIZW55i56tylq6s6QcTd
3yVPTDyhmocsMY9ny35YHHGqEVN0eNYOGBcq+0VFMhmhA1hi20wS4Xz0qnxkrNKzzwdg7qBGP1fA
bbE61nFH/JibFUuBktLwPegOyyhJrGQVF/q4C7n7lflcCyfHRmpuYdREQYUiGBlGKj70h3s4QKSN
6Zy2tcUByQcmaz+2FmJhEuYDz47M0pxo/POxP2N+DxOmuqQCij9z14ZNziw1HNAaqASxLIxPM2t7
+TiXe1ens+FOKZMF1/VS04jqlHYQLY4LYKvZWfj+Qa0L5YUlPNG6VxHI0P3q33oUral8wEHoTaGt
MIEaq69/aLvxLqs2hVh2fKUEeG+m1YZcKnr+RqyW7dMYKyZrJ3yr6xU+lLZIAgKWZEfQrPV9YW4S
P9TBfRELsTM3wA0kXtofFTJSynhxls5i9DHUr1No4Ph9uXJOwMqULrHcAKW1ogONfzoGDRiGdTKi
Q3sY2x3OPcuAGMOzwsDNUrhuRtm1zzSge+zyjBb3vTxLrzT8jwx91bhDOG8NkD0Sy26FByR9mCUu
7YCQTpKk0V0G/h+444F5DnYx4rNma1710xEn61axxnJLaZVFEte5HF4sdsDW04Qo0Lj6k7+lGQMa
LvNjve64ppUo1qMshfZXZRXECSnR39i1PzvCFk5gX47y1XC9Doro84RqOEHF0UOzg8NgLixIDuui
CBPE43zwjISRlX0OPhJdFNDkg+jjn23lBx7uPLPhON5amvCLikWr9J+Cpqsqv2heOyW4bd+40QoB
6T404ZiO0Oiqq0zIEqGybcq+ylKDrIM8cI7BKM4X2JY4+yIL6uW0591BZH7sDVWJWRWIZYp4vKS9
s2aAzknQwfK3884E2DxEIOSzilUAmtJ/Pxf/LhTAKfcQPLDl8KcWk22MNqQiiZ8uumFJtG8gROIf
7YisfN9TBl3XHM7isaLz56N4v5bOUCQPdnyrgziYL7VdaNQHzxuRSYWNBdg786nIeokgJwHCAHq3
nZzRuD15D0CHn9UJJL7JGeKwtEcjboyYiFv6y8e7DZUpn7N85u/a10Xt+tyDc2XPMC0G0fOsw8z8
tguRb4pyVfYF6HlmTqJm2E1FvKZB97Njukgjcy8+bzjvlKjlxkRLRa95lbNNxXNS9AU5Yfr5eWAk
JqbvGt8Tyk5bgwP7ffGQLloMOTUvlEJ6X0yoFYbBDLkzsg99PWx0RaLZA2Jg6b/RVoB5g8fUTvw6
wSzerEqpyEMmQaaf40+NwgP18waBmCDn5LoZV0w1Pp4y760X7FoHQQtFU0iqs/yNVvtX4SWlCAjd
Dyi/sxdMEYQnx0wmTSgL4ScCQLTfswFoUDerJ7Dty9kCTtMkRDQeY9WzlWBcTZ/sDOlkoy7dzk2q
zZNzf5VlYmBLi8ppIjF6pXaEUeHTPuLl/y/EDk2wIgfOjhlJmcweYSZwo7eHJD3jZXGd6zg+Oein
iynowS8XnYKPWBigTxL5EPlz6xSVOGW/DElYNxCRFkqG55ItBd2UtJMDuJe7XG4f1IltNfBfiAvi
`protect end_protected
