--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
RNO2CtPAK3+IJDITWbauUhv+o9c1rqhvqfVfiWPXFJ9h6tjGQ8wy5iFbXhWTkIOxuz/d7d6NMHU6
a00RKOYORyXAl9YHDDDcZvfllhXj1Lws2VCPjYDat+5J8FAqoaw8bY+MTFiEty5sc+jaLXaM/n+L
PZ1sNZes1HN+lnuhQnXTLojFg1BTHdi3m5AjArX9eExYjOx9aLrcNOsrdRNsvZ6GK9jwWmGgEw2R
Tl29QZCr7cC3VuelBQ3aL4Uzvl+fZP9ou7F3yFo15PtHDjSyfwkeR63El/dyHhDPYKz0Aruntr+T
D52p6XfHN07IqHfdYMLla9EbmdJ55zEvqUc46A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="23LSgEliz4jzkQk8Wd0Jn3rPkYVlN2SNW+ZCleW3yvU="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
YmiE1ZmqfToAhcB/UfEPXN+WzjyKCum++uJLdM6/imR033TpkeIwtUlmLe0rRzLyfDFo/3Kifs9q
ifIZKx6+WCyH+0JJTXGeFWU359Fk0TEvcpAU8tJPxHXWmb7wd0u5pTPlkYfeABG4nM2zo4UT2KCQ
IYDwnjbqi/o+7x+W6VEA9LUwd84uSvLpxks/0CG0XL+zyfxagFiePObFISnytGPaQc7woxBv0KAF
AMXmqPlXBwEPAM3059lsyKomTMVLh02P4fPa9cqHm4yZ94Q4Ley22LsAm5xqvJiIOXiWIBjdusZu
nB9tRqWw7TX33txJiYpw7eCpqI9Zlx57zsWCRw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="tFrGzRE2dGORr1NZ4GL8eZIp/2w+R8oBv8MIKdznmRo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15504)
`protect data_block
1vrWcj7dRYWUPN1gGxPr2dxl/HmGFuBPdQ6c933EjE5vuknn9wik1Z6yHkZFY0IwaRdYobHWq+ec
D2yhRbZa4wuVEEEGhwf+r1oAFyxADN7qNmi8FlVJRBjnUxGpaj2Im3JpI0IRiyhb+/4IZP3zzPdc
QBxO0Lg2ftgsPlx6SWcDN7GXDCANpLIQpOP2WRKyt/hWIs+eP72mMmLo7/YICB/Sk1yMjpg5kcRk
ci0PYijLYmHL6QcA1HUb6xvD9ByKabOUU/wsOIKyBFBfBn9NST/wxTR1KTcT/Ea84mH/AczDvnrx
nRainhwY7IUrJg6Tif3yuaqMDZCmRfAiUF9NxL31cPB5pQebkb9yi7SQXkURkCdNzzPFryX7+max
BgAJJu/lnKMnH95fH0MriDVt2EwYo0queHO63lz6PvU03xLA3aLjTQSW2xoVGwot1/XjRwcr1kvl
dCrbwnlpQoS8ZQ08King2617xQbEkjB6vnAyA+o2euoCrqzaLFFNUA0hOuVxJLU0EO5xn/mi8E3D
TSE+bMib9Rg7dezv8snuAknlLSeEJIhChzFdwQXDibefPVOGHLsLD54hMNfUZHuf73eUsxmd2OXl
wWoPjWefI/dgDAuLslk22awn1jLFXVL6zNQar7nvSGwGLlJ+iG4Vz2xkoe+MT6z1DCpQdS6fl1ar
9jmEh5Gj7PVRyuju8e1vvqTSbHpf5ROVOHMz+/ldSfJ6OmjbkLh41jbf8rGvSCZ1kmGIXRZ7rkN7
WTsO9YCIZGbybRB9mlJIzjIIYVTLcxtPiURpQbcRZsdz7ZcrvINeFoPB8Po9nB+cayEDXlooWMkt
AZEjiuMasBugMSvc9X2M5l4TD3TnwqDwEg7X+VwmnfvZvQg4cdq9EIYFzZnQetxLQsFIKKlXdrb2
mlfuB6xdOEgrcOdjoWiBwAk+VZTQJA/k0bjg17ra13DkN96nGIy62VIfILrhNQQjV1QJA3K/tuG0
k1yZXi5GgBo1dRgrWZ9syqrePrbZxx+VigTZQbzBCL9fauFHThR21qx8x17DVlI3Ba7K+XQoG/Vb
IgUQ7Jid7FVA47nTDA/sImBErIqWj6Z5oUudjTy6LvqjWbhFfJ1v6IOcJ29rFj9vSieUfhX5TEBF
RZkg/q53ZfGZV3iRx/tcJQIz1J09Uh5vYMriJ4YAoaypAv3FgOJQ5iVnV+IRv9ymDCBkLi2BcG1H
vLNK3DsR9nTAAC9K7Q84KF8VPg/isgTEFbPD6k1f6JMEJidCZNutaOxb3Xl9q921gZRP6sRMm4Iv
UTxyvgBKZKl4DO5dgPqmBzs27Eg+1sf8iUgJZvfTiqghuuRGjaZn1x9HvsXSSUweCjTUr0z/EY4A
TzdNIORi4o3M1/8V7BriS895QhOp1BSh75dI74W7qG9vJT45tcR1QyRZ74XdYdNRB/XgOWwrYGE7
WjsC/KMETfcrS7p9OJyu88IBVSueZj0vqzQ6xsX2LNRtl+hl8hdo2msjZ35PZ+9FleBjbjole4Oe
TqBwoBYkb49F59qKwrGE9C3p5YVZ/WK4n5RjT6Zpc+CnsSlYsEpBm13pfqNeukgKY5+GOzbE8EGQ
7Rpga/W3/AcukY/Ksxs/4+cvQ9+O+B6fenoke4f8URZAFAGg72nJIgFxsd4r2u83z8VAcWGgdPxS
M1xt9ukIGf6mWTM5nP2JdNxN/Wi1RSU2Iq9MUSEHyLQ6FwTf5KCeLuhZmg6wjNIZARubpa6Q/0xE
ndR3ZjzWog4IF/uqqj4X+e5udFKwBtIVRjLbhFhwdUbhwf6FAuUhOBwgy+TqvMafyWdqDYcksOu2
wlEJYmcLzOvFHxLB9AWna5LfXKGxerJXIfsMstV3VZpPK/2kZFH/ZsVt9gpwE1yO/rh3sD4HbO8H
n/t3PvzBlmdVHXLCfA4OWrb2X39PJFYre6nh1mwJepuHJTCDdYSAV2vss3D8tp9wSALhFJX93Hqv
RAExz3qB/0+BIcMzB2ZbMlGjHKvip+lLQ4y8S//Ep7Y8+baACf56KuL1lJhSSHbqH6HuWQgx+tZE
0HzdLExtcRVxddJ/BOBvoW3irLIW2++W2zzMsA+Oz5z5MetlWHnyk6bw/LF4/oYWLCPtfL7ocTM2
lu/QpPXW/0G/CQrsPZq9UsiaKTrm2Fn2m8yKj+a6qFFjejKxh/yQWvVsfif1XfomdYf7D/zzKDAl
y/MXP1jx2G2kLzXDi0Y2rNE/7RMKyMDvLEOVV4OVkWi5nLYD/iBEVqp7a4hiXBTV0r/vzH3sL0ch
KmtkL1FfY/FeZKQtZSqJRTn10qo9Jp3qVFlqnFjXm7bfkKT7y3nRMJxxtmZirf+LmNgh7uNbHR32
xpzXQiDwzqeGyQyy14X6u22reFRoVu67gv2lDAFjDqoomKEx8MPBUwi5T3qFeNZBwudIh/DM2cwA
n3ug6cNl4D3kjvm5XrNAcP+t32sCyFRRAuNcZXLbtJd/rBzsAEFXaqaP8/W/2LcFi/r9S+qqQP1/
24zS1FCbiNUnHh8IQp1jbnMQagq+6G4Su2NudLOk7Dy/AP6ZDfm+z06/J/34ZFzLHw2Z9Y7HA1yY
Ej3a+fp+dB51ezM9AYRSVl8xDvnE35k5E0E4SJxbLSJ4GR4uDCw6SU6pnyZnJNwfjkEclTyY+9Kd
HElTxRAn+b+B39y6nrM+Mhg3slSX0HLNJOyTnOJDCLXg82hMs/mlVXocAS8/wU+dykCuwXixEBJ0
qoQdehIe2sN1pIQjBjcrcZ88KiHUwE/K/N/XmA/um9x6A/LR/9F0fVZLtjDnFy2tsFvZ5KvF51SK
ND0JPQVxWrYoj4+MUzGwwujFN4WScE6uCpTrdEjlb3EB2dweKUpG9TqXR9sc3QkYDVEpp4A48xdN
Fq2UENZUB2tDR/VGDRkaa0yTokHyN+3Rr58VnG9dU7vNsxW816tUxnur4G+2+n9ejy5KtQMT5uit
StK7bXpSydDhfKz2NadJh3/+MwH++ediRIoLHIbCd64mb/1F/6oUGwTMKXftmTJrFeqQ/vhtVm6/
KvtujqvEoWwnBzhwT0ONElJ9zTjyka1twoJOjUHLeO8no4SMJI5wjSAp4vp5uhW2JD6nXzCzziCt
LHA1KQnUwv+iNygTIkv7rSzGJ6yC72tY3uKkLzDdqKdgNhDB3Y5qAdg+YXLfP98cLfaTn+z9hfK1
hXmmHq36Vg84IsIo6e+EYXTgTsZD7uRJdCaMRQSLuoz2Qihd4rfaycQUFan72IqaM6tmUzPBeD2G
kvtdV8/rPsaf1zclca/C87W+mUq+m54fPPcwQAWeFbnSaSl0G20Hc8u/H/xGLR8MuyfLdkZS6VsW
RBtvGMjnmaC8GoEq81SL84edawaK1rHFJ3D3r0S5Oc1Lxo0dNtRLK22ZYCX2ywCu/XXdsudqUNHI
QxPkC8mpsD09Iiibxu/zKxyyEx1w+GZ3rOvT+qnAwJprKjcMsfRQqHjTXscKGKXOx9933bvwv14k
Q32N2xSy1sODpDtg8tPwgg6ddU3dE4V2jnnH8qqvMjMAVbeSf5i5bIMCg6pX6TWPUH3LyEspHWBn
SYI6HdHnPRDNCEHPxp1rK7PuZ1fU5XqGefL7+j1MwcneqS0lcEUsUpqtVYEvTCwFEjFitsjsq2CM
8WMaPzlGHnaxQC0Qc0XYAUn0bWNXtH01NTn7CbA15tnPLXGFa/ow698JSohj95GtOSDyqa6uvXqe
ThvR49t98D9Ih6hC93MZoK6Cha6jReMj8rj+tVNu2KmCDCzbnAuZI6OdQ0ZqvCSBJ88PPU2WIZAT
DTpweoQmwQTvR1fZuAQGQPkU1NTkBHNWZQWdlr7mNzX510aNYB/AOFQ7IEbfUQ+zLzUvPSBHzqw5
0U+UGqM3XQ4chvm4fLbxOLFF7qX8+xGVhDImjb1iauzJ47+oLgp8QkfBIhjYxFFXoqtRU8Jb/5SH
d5uhR67MfKqvTYmOVc3vyXSiSjOgpQmCcKmLXdJ/PWn6TNGmdrqaGOCLwI/ToZPgxjOYEEL9cqrG
TRaozI//GvMPyVgNlUSeo5S2vodPEYAp74jJGDbCcnB+Ik/v4dAo1vup6ySoeOLmefAcgRL7GCpQ
5XAnt3ntobjjmhC/I0RT/ct7gR+/FKhIJ1hm4gwou++CkqgGfyxhOMqTIUwZxb1DCOW5i/N+x+/0
1eUbIKeScbuMoPKE+OLwCouY8WLRwnV/cU93FZUXAHx7Jx9GB69ShCfRrYYZlrIsP7hlGYpvRXGO
HLOGT7qdfbQqW9L+rSEAiAmYapZ5qZj3SU4W2n48YIo6jqZbc4VKLvMNdOPz8rzO+jofYk/3Jl67
8eJ85yBfMG5Nz76O79yFBIQ4vaUyDrOJ9CoSRAfMZSI7PUtE+TaPE1L718qfAbGpVWgi8VKgCYzY
W8uxgQ4rpnjCIr6X0lFK3bRzrPR8if05ffc7ZaU5zpF8ygMYnANiQQQZlx2AiAekBPKe9+7NyAer
3/imZ4RuoW9rpY/0VmDoFop2Aux1VRhKZrdObZSAyV3M7qjA4r5UIpLOl6qXWGmFQBB7Xc8zpyBt
Zgdsvfzxo+pXytrXIOJYm3jcNMx8B3MdWpTJ4qW4cfx8/PRR3Z3IAFxEJEniqbIi6vfZ5qk9JtsD
4AETzm2vr2yhUtSZuLaMoKvEmGH4zPfMv1lDOWfpyrTKdQJywrWJaHrZ+hHBHi2Gy6no+oZisEZF
23lYyLpvu0VSh5xQ1ACJTxcmcMg6MvXk0n4viz50T81DR7NxpTeJk6vzjvKXKNUphgEzeK7/Ka+7
MvPoI/Dwwgsfm6CdZ7uLngGB2HGYd5fGZHEH5vq6woWqy+hC3y6XA+p+fTHntzsJ7/+XTK02glrB
0B2n3bZPlNVBIOGp9s1xSv1EW1nJvDitNKPjGJX7J48ATlD+Rb1NU3xifsqdAgYLXwxvSAhuCU/b
UewzpoBCoZSpiPKUoGZxh9KmH1j+Qyfi2WZt6lv5S+E0ZQcisNo2KMVvlM/wgdHq69w9ng0FGvyc
9oFLT2RLcF3oLutkhtIm4JX39+6V1HGSkLCbdHDxqOPfBdk2vEGPxvZ+LgsZ3LJkvTqmht/UFSQZ
L3oEgPf8t7+Qlb0zxOSKNM+rRAA9WGIt+5Y5ik3ZUVCBZ8E3LRDQmDgwXAg53Rb0mc0DZRl3Wmdq
Q7FQbIzf6oT9Pdi3zPcTmYRU3V3YE/AetR8bI+Psp2OkZlU6gDWQh2Em/y3v0ZYzqG/7spjZQNEX
XNRxeGcRj3TNn7CIYJhZPRR1VsrUPi/07gfnPGg5BzNsCqidmhlF6ik/aJPLrF6jes9YXDlgY58p
R4sg56rCtvfHGhiwCtDF3mFwksEPWwWQ5Jg56xnk9LJzJ+bHtzQsDyTOcMNt/vcBDWNR5FWdcxSc
E9pfGwvJV/9n7duuH/9oW760BbBnGO9ouFJZwb8RwHFYDkVXX0uI+ufJE6OpmA4nJDMEB48rkDS+
6KKFSOi+79t4bCm6eFNW+S4999PUiPKQJEFyYTF5SWWTzofrXOGIdBEmLI3jYbPt/Y22uf6SLwuc
w1+SKhMCWv2yZNohYZ2z6yCv/wnTzva2GtaarZfKfodhD87Quo4OfCa4U1qK2TUmiln/K2qMR4rV
JsSDt5z+08JYmwUdwwU9KtRr4CRlzBej0i4oaHlo5/I1+hyOf0tk3Pws9xbSJSkk3bq+RqPp40XB
NZXCwnvGjjKKhediRIiq5arbw9hMBqA5Ug5b6IQhub2qYKSGgcYzVn/1+jgw0x9m+eMgTP91rtwE
Re+SpJLwH971nR9+2anKz0bSa/DYPAeKjpFHFB5VLxDJqvtvRD28pVHFFjppHMy+OWR84HHAYQB4
Efe/PXPHiNXI7+5K6VC6p38ytDZRYetP6FKbUzTRAa4dIVJKn+sND33S+SEOQqPCLzODdYKjHJTA
lRutrOvhV6YzDqkIanvXcdL2StIpkHzskHw1jETeaOcPlsprX22ogHGPgzshvD9fVVLkQANEmvmX
1meJArCSdFLaG47p40ho0dgAICGTGze92j1FGUpvn3LMPOMHxu01vRGhS/4qexWMBldirThendx9
TxSqdxVyYgJqbtkxi1UnNpkfLhNoiUnCzpk+55sTOSL2JiuDIsQA/kHOh2uqsTwYvum50cqOYlkx
HSmRSsXXG9zrYuAEA2OfnTzuLCMPuxH29S3P5DP+1YnfKNksMOf9LunygTsvZLvbxS1KWm1DxJst
MeCKjehw4c4st/+pS42EsVxvMYnVktpbIzfKzAsrZM6ZVFdrh6xSL9OPhk5dZcbxIIf/oUdihrEQ
WyN7JY8CLW3JTbeHZtNFSn68YX0pCfkuKtj5pLg4XFBV0TpS27Nl5zKQKhtxZeU3HSAptjr4WDv4
uLlcDZcs+7jpGRgOD9a1EaJYOe9cxI83iMTpzylR479xpiVR8ajseo1KXLQ8Ecugz61V1XAsJ1V3
0d92qznaTvLE3XJSw5lLXbRNvcO8mjtg/lnEdx2x8COPlXnH49HC3MznmLXS+nxJNbXSbK6p+KeK
eU6XlzUDimf/6+U5/dYDJPACtUPYik1rCF9IFNFp/F5cZvrfGJMJFhA5u2+rMcKqj0UZ96PFjifg
fWqd1c0WVYTW63tnUShz6KCjqRfCPl7CbdDKFOci5rPbHx4PMA/B3yvBNcwY4J6ogfWPUsxRzZiy
wnbiljsS37EYbnaJcmNMm4VYskucMIgnN54cVxgf10kihYA/bF818VGBEjC3I5VuW+lPEtOu9eNe
Ig++PwZh8COcpJs902pVjy5UMVYD/Tm1WJArb+PzoPO2QIfKp53Bvcp41jgka1CiV1pKdgX4+O7m
0KL4jV5F7qY2mtIscUQsVd9VpHDN57xmd1tV7UTNTXX8Eozz18Wyuk14/zmvMIqtD9UqC0MgUUdS
BequNBlMw4UdjzgviTAePBglQ1AP87Vhp8wjTcYodboN0bWXHgfA66/1PAvlxwVfokxMF33plhYP
sy0h0lWhBcEe6Zh2y8PpMO8s46NqtbhsebsEeI+S9yiX+fNlcN9MeES8vwtR9gvaTpfLzVDAUnDq
e8GkLNmhLA68iZsEuW+XVNyLU7fApONXLcNlP+rN4C8SChFJpz3SdtO3GNRkDjQHHG/8+TfqTKJU
G/zuy+kpfwciLemFta5XXJdpIHvulUTuzTv2BXKkiP6UfT0iFz0vIYtiAZ6m3ZurBT6jcH6Rl6uu
mXSub2U32GP7fJS9qAOfwChStV30jTSnDWgnQbwxcVUjKhcqiTl2bl7EGudkKcziS6nB9dT2hZ+W
TA8IEX85zO/EBdiLkgSsBPIjgq1AXOXM8SC7FHU3byVID2IvT4AIhhNG+uBkwPgdqYfFD7yaYmE/
e8bfFJxP8XxE54fQmTt1BdLMTGX2SKcRD4E3f5R4OFHCJ5FNQSpCDhhp/V4qJYbOPTsJWn/81SW9
znRBXmMZ6oeZP7JnCvmC2JRzcPcJcoPn6Pn24K4W/zYVIEmAlRYs6/8oxL6RHzwu2TuomYyPo7Vy
6HI5EEP4LxwRQA9T8l4JT64JTKWhDDLcFk0GtO8JbdAPjBd1ch+3tjnSbCcBiDAe1J+yWu388brW
C2G+gWuj2WvLp2amolY4NmDBqiH29HLquXGdcQozb9bDDOkJoYMSLfi6ZREF2Umpzj5kCtuLpIYR
k33iqiFsy1Zxxl5ktNLLt5SDQxpLtlSk0Cf7PywxbHY/oLB0MYOxVtyJesgn3AIPQchbNbQSBOCp
1e49BnmjWl6Ycbs8QXFj7sdDeECxySYtXh3M8h6R5FShlFssZ+24zZVnCNvTQAeDXBY1rJkQf852
qnr/L+d0C5oXafZ6or1YxYsFlzNpS539Napa3kCC3l8h/jXZbBG7lAZ6NRtSOnItxxasykaruC/t
JU9ZKLmoV9AS2lQP3j00sg2QiYhJEj8W4N64jg4JMXRBacOKkQXnWyfnRDIrKxCAKXKeHTfOGITd
pEnC9c/4rHdrKehNX/2OgKdE6UXCGFbhj9mIKsRKu4Z3e5IvtWvR1jN0OLNNHucczBJmfRx1kUUm
R34QVXd8VxPp/U/zEtUvqlbsBJCl+Xi6d1HoOiLvlPY0MDQ5d03GTnagH0oqU76ijZ+pSnRfaOle
wB7khoXfXW4Nagm6uoz9w75+kjv6DDUMysZN6Bcln/eCTeWOIlE8w8OqMbL6cUyvQAJr+rF0igrm
laXSaV+ove4fKYncYkdXkGUBtFyVw0v4pn0qUB8jSHIq8sQ6/R/Wz4qoXYeeGKowirY+XADPQgSD
CxmXIpiS65Q5eQDOBWFejvAgzOVm9yUl2NIU43PDIY49cHyJF+9neTFY6dXFyz/w6hHjNjlzmRtJ
jyYyDCnZLgRd8QqMEEoAegeoFtee9M5fRI07+Uk0umCL0r1ngQ3zebpTq8E3U1odIEQh01yU6xQ9
e1LzUNgesrLSayMbOk4pO3H1u9H2h+zJfydA/mgGeT1LGDkFqt9BB1Jp0mY97CGya1mLDVZX238b
Z+fz98MPCkOgxKacuOGSFpXo9NzH1KJ6HyF7wSJ85M9Jm6EGgyoohz4/3y31wb0t/jq9HHM4L4ms
99WNkTmpZN2U976ASOEv9EmNZGYFLzafQrm5fprBx68q4VhkgvSpqbi7+MSoZCamuN0iw7ylzu7O
Cbb/vJxIuEJ0L0EonikFt1WJKojRVPDUHvkVrQDXOqLKw1/hZFHZWko4MaaISVZiviYfJbzkZCVy
w6V8107iSordbxYmA1v6DMXNXpv+N2G/gue0d/A2p2Zp3Tjkm6aJgTVxWY3XQzgE3kBJSVHK0ovZ
HiG5Cyrwr2PxZA6nlUAmA6fFpWWZhpi6Y68Oa4lOhCx+fzkdgsk8dHZxOyRoqYo8XJt3A0Rorjzp
7ao3HObP2OP6Uc1yk9FVU1+lPe0ljIKiFt+AvJDQ805l/2HfSGZJcYz6zwS0X9vNaAQQDaCz7647
eH0ZXXoZwaqCOl9z5WzLRGGIpGzxrKm/zkZYHB+0VInRVu5U48QX1d5qDfh6TBTBS1O3aYQ69F6k
gVwl/Bk+aLcLoDZNuznuS7I2rBHpMmKF6rPAzKAVLPJq/GFkMLInQnam/pcw4pEa97Rn//yBXOHD
bkzNsHpbxHuG57+hyvbqIImX7CsdU4e8ibOzUsoCJpDKMvXF+nyZ83SvIU4Vk3TkpnLsKqlBfpl2
YgE8Y+cPDnRFhRBYfx/YV+8PVMvaL8rYOmjbrdO53hzCoWLsgcTgpnycbFzK7+a/01rH4VsPPbB8
2Xa5f/QLQSkOhA0vS7L1C0vIe0LOM8BH63Kwdff8NSHohIX1cayHGFdSpoWnZnDKyHbHIMtoAsRe
z37ppVvMguoTT9PYTTzX42oSeO5sAS1k09dvW7ogRvSk5LJISmVsbc1jyAIIAtFmoOfP1H9Wk5aW
mMCBJSj+8zA93tJDvWOsOnDLZY+9BLtLT6V95abXE9mfLuLN3x8fQujYGF3xTc7mj+tfG9N3xZXG
mzya65Oq2GP/uLqX4JQPSbtuq2r3oXptt/iWcDlF34w/PkoafQQw8mc8+lY8vqf8vYJ6Vm5g2mEF
IscWNu89UbhAzjwQySDvJTxTy2+JM2bnQa5U91FgTbk+hqxQ0PY9F3bTZHRIAjlE3pGFrADyLeBa
zALplHJs9yqZUmTN//XkNhwdR/1+lJoArDvsD4a2wTuzMUhj1+vLBslIwML0c8tnmjEFgr6Xmwoq
WMd0WA2mz4pmccymXaPYYgP0d7xhu1u6L4+sHicR3FcoHuxFB26ZcydfnRjNB0RxuNC9vTFwD/hO
4KrS8fYNhhXkf725myUck3cYp6a/2tT6tQV0ACjCRTMgsjL97Ai6bKyKTmsyA1rAq7bvjcMzT12T
j7qmfAH9lACsXZTiQv5yyNb3DgWb4DIa+1p9khaeGCT1qfjLiTxKaztNMzM9h85+xlJdI900c+ge
bCQb3/Mo9H8i1+VGI0Fpv+0oxmfJ4DnznOWTo3U1VjwnbHeaM3by6Lx7lLlS5hfCJxhCVC21hFkS
f/nfVQQZKhJpadb36WrtQDEoLteooXSDcfHJFjOzQKHZ7BQrRC3KToD6sshGRqpJ4V1t5U4bSQgw
b+mc/9BOJoCQgc4O/2LPhkNhLLjP2y62duiD/N3T2ayvpFXat3V/v9CtOFVuBRCZ4wXefi0adegh
0+wV3jp3NRWhiOfxnTSOTMXvlcqUA+ujIY/qPsttlL8GqIwp1XqNWnxKtfducW+8S5umpll5Fdy4
cEJLDAmJkPVoZ7ci/w4nLmgcCouu23GW9H1zfzvZ5mYIViTHmR0DqY9sptdHhFQHSzfsndV+Ucu0
Iea7vUudksj9EFiIxJZplWnSR2d3RTWNIhp6qWmdeYBES7QOKB3RLWxJK9ibuu0dS968R/TS51mh
skc1izSrKDZzxGyE2UtF+F+giqE79lAN/F3EA0bAAIurZVJhGbDtJWEh1YGx6hRLY32tXg3az/3J
EwzsRZ+NREZx50ya60hNJkem0EvppZR8eKoebHtGfqKAZubWDWkWg4HJFKUYY8PeQLjo2pgtkfHn
MRGDHdtFyMvZHFEVMsweWzenPzGR02/2QLCqiuGC5McMwdYsPgwNct2ksuI2X0JGHFWyTpBSa+BN
EakkoN4I5pszaObLPGokDHfjAxMlEuUngYECgUmAugPhipkI2B6kIMKwJWekezkJXoz5GTy8/t7j
kTsUL5GkbdiI+cRUjVaOT6Imld2ifS/1cJwqtdGkmwcrAwDcww0Ky5cf7MTPKBiFi/EiyTyGtCEf
HJ2ja12AlqXXqdN9ww4VDTmH9o+daZ5soHhoTyAqlrCkIB/gr1rxHaXkWCS1o6o+eLUbfrZxL0co
2CuMCZI0845iZ6aRDEEy4ylpql1aBk1Qv17HWsfDZ61dE8fxtvRLCzB1vXuJ/vIadNB3i5G3bXxw
4XpQcZbPaEye4ewJ2swSm8envS2E57pbrU2betU4fbeG7qQ3G/mcoMbBJJAgVKIs5UmCSozvTQ1E
94D33UQHxw07bsgiZcrNEvnq+nTjg9E71JKKDOJgER8bpWKh/6ppbiMKYEnpJXtRlqM4VN6TXzXe
e5GwsshKrXBSqYXP0iRVP1Wn9rcNJhSLgvmGGeNb+eaAEBuexsJSwLmj4ovBcNpUYU0v0ZSd119L
DvOQqh/w1TBiWZOu8bYGgUwV4L0VutPXJp40lR84ouEWfkYR4xH2Yc5QaMSu77LhhPJKfaSPh5vf
qx7mt15IRszQa3I8qWxFkPwussCwhGtxUfW/0rL5Rlgyw1ErLMmXofb78S2oP2XSIB4K7HeQCNi2
K0XaDp8hr8VVbPx0qdoT0EccHFaBS/bMRD6S2aHUBdE19nE4rBOxlk0eCAwXbY76deJBUDqD8qDe
zTguNwOrXR1fzHvoOSDK9T58H3ylswU9N0qhTJCZDvB49en9sXqY3dfCN4qxjJ/TT/uy50gW6RGG
7C/fakZqZXxNOvdj3vhethSbldADcAPCvnMwhOej5buDyAJ9yE0FeTbP1oidf7DjsKXMopSK2YYH
YxW9cO+OaUgldV4D5ZBpgzrGWnqh68HEIeRLJuLxtZgZbS1r/K0mJYqfpqkwwVt0bVoztojB4+Zf
ayV9voZXNAN9K1bZJeiGh2KCQpIHOrlM5/isEVJaTcai6V1rvbgF063CBckGCUs3pF6uzSI0BYYG
06bHoxxFdrbdJZd/FcSn570dNRGrUEYb+iwB3s9UPhRPtbqse/ZuM11LMicUpOtnOGEkK3PyuNmK
ZFiM+7AZhmitqBXUBRuXdrS0024Tji/DgO8+2XcYwqJgtAfpPexyLlc6C9LuhoxkVb7n/u63b5rZ
f0EOSvlz3yh8+D2mLgR0ApeTJlf3BNlNnwp7x9iXyaRbZ8tH3UBhhqwnnkShb0ZXmjxV15BpavBj
Supl7S/GnYXGEYrXIkISKg1qgpk+DzsXpMiwRODJR8EK29zpvfORuFmqMqKL+SD/00F7b0qaWcMe
Wtl3gjJgB5bZMVASH/t2K2DgDSfGfkzf+cEgn2XAonDlWSZfwiZSKnIZwuETrfCaEMIidL4zHy0T
YkF7ve/cDtAMzuwwkTczBxNYXGPaIlvI8rELx94xlHjsjYcjx0IOkYKfbKOsTAsxbQsKIZJpPSRb
uTUPRzrlvQp4bHEqtextT6qOPGtbBsUUO9661XLN1ooDe4KMj3JDfaxps1eBQLmzY/KGMk6pob4l
f6UHrvp08w6Ee+fazFMLuQ2jruWZ7fMbMUACGX0EE4aILi2eXt1lrEt6/CvK4n6GV0BfvITEjDet
XLwwmofAEuy31sbSOnP9xJvDbqdB3X5wpGseyQariUapi8TTOwS6ekqEaHSNx/K3kvUOjPTZKwBi
4zrKqPnUvD6F1HsArRrMwQIC8olJ6DrtihkBOHjRQFjt1kxjMhRT2CTKi+NHiN2WByTFsG30tN7J
g+ywyNpf7/FyeBnLT4erO+BtQIlMKjXBum3PeV3ugWPlbK78XYq6HwULcyJN1pmkNTYAd9FtNLgE
rEgly+PTgfSpmNKiL3UdyE4uMSfPlzfNgN3JNaVz0ovJsSv/axAC3Mx+3+ftDCGlL9cTT5JjstdX
3DiVe8QD/OTJvV7lq8YJWbm0bcf+Fy7yCK6tzyMPW4yCQFC8Nt0eNdfr+8U/8TcDdg9zUTnNxIOx
nNBFAdKEG8e7BJOW/V121vH7YGMWTZcZ4TKNlohtE9gAW7OOUZNdGbDXceSVHWllGHD0C9x7L4WU
3salG25sqgWI4k9aAksFg0LBE7kw0iBfLRVPCnr55845ZHkg24QfBqGqaX1eiPZzLWiBxQUIboaa
8XuMDLR0QAu5oNFERveB9/tQxV5wcHfEhU6USZk4NZAJR9mczJZ1M9cE0le25/JLbi5Tbht6mRaJ
3w45hWjHrftsA2Gk5H0/WQp8ZTZVRwINvQu4bWiYLPFNrdXouoRFuJ4Lf9RxjsN/WEggCa3cP680
Z0U4pJ74AsJ8PiLY2N0nGOa2G5j9yYu5iDnPxO+nxiSBBAJxf1vsIQNZ9fFgJg+lOrKLyOs7DBOH
zba2NWSnRijoiJz7fhECCIPMgB9Xqm6JV8RnkIe+PZuHvnhAPqwfKVT34gDeTnfpsodDu2hHsXtl
lHfHHWPzWdW+sf0v8AebPoxQm0k7VlVnMFqIxvglle2BYoSrXvzKvzTIhUMrVt1YBDzs5teAy+sw
VQFkEsPiD30h2taKoJIGlA4JXAsNi59vzMIfAIatZmq086GfxzO1As8OqtY6/7EG3Te9BxoRcDOl
Z7ZeRqf70WjdBdigntRYNLy7F7pPr2sPLUM44zSFMnEz81fnmAcPR0hXJTQ6qp5NRrbpibC8dwTU
AhTA94js5pYTimH+e7RnzaaYXNhuJQdJzILKbAcUPI8iLxOfnyA7HJEX3dBeMB/skIMeyMYPoZJV
7TpOiGVIYsFvRCQ6FLgC4teK/jpUCF4yFD2kA6Xhd5sZc2iVbuL7xnJs9v+GaIwirnFo9+TyonKs
zv1jBnmbP+8ZN3KUdzC8MPrJO0n3hTqnvk+38f/HfPh1Qy4RSeiOBQVKr9bNNi68L6Hhzi22/hk/
cShthQi7Hqc0qeA6TTDxBPc15kQxP5l2ZNmOMuIBtyRknoVGGz17IQE+roteLaVPQ86nyoDHPBNN
V35C0cqscs2+ILUrNefTBJ5gPJe+Y7wxBOmam6Kc6W8A1Mgjlo0anxOPdp7U0l6IDPwVed3PPlzs
v2RriyEYiGDAfw+iJGuKEvnfpD9gkis/lT6mKV1ibmV/UP/NPg/RDW8nariJJw3cANvOjSW7iJzf
lhgKxFyXgGPG6xVRc0obNj+goN4lesUYHTr8ETYyvfNpvOSNAvQ/Oi5/hliFYicFO+qMHT49b8vT
XxpP4X2Jt+3JhRKwDY0dbQYs9r8p0H4DU7zvOKGYT2Qbowuq2dvSK1tZ/+WZCcglS1fkqgy3Wqxl
nnxtrKIxfxYTR6SajRmwjkJvN3RT2psrBt/KGTVJkPO7SSzcjXHoNa1FMEOd10kbW19hHz5QHLyb
+yv+M8IyaW6QpYGeEO5K4gUsjECLEMF0HI6lLB1+yH3N8yRk3zn5YRgkNJLBTlednrr5iBxoALXj
iJU6GKPZIDMDrtBtZVTQqmfSwTIDSaAZCzWEMInb74y9H5TTI5KGHS1fg7C1qTVy8Vx+y732aMgK
0E3ZTUYe7YA6RclABrfXBV7PvUqXR8CujowKTMgmoxHFW/tj3S02dokUw9Hi57OqVC6hBhDvnXY1
pVHH2QFbKkCiML2U+tKqhiMa2t4HE0Muh32DY9MQlT3wjxHdkJUjnnsuZxMta36r1hbdYOnoww6Q
kQI0fGcXVtdJmm1cKuNDgTjWLImmJppwTAzyKUg4PHGlXsuEyTntn8DR8WcwqNbR3dVudEKLY7Bz
2p6f/OAZDkTt1zh+8mAkY6/Sq6osbqF4iJnhoCRkQIiaSs0KxifvykTEtHejGL5MHRouaoESM7KF
te4RSPXQOJNJWIcfvbSB60U59vUnFlXOmUyGKuzLM5+FOuWQPQ9zFE9dYxLnFdHD7zcqG20Gw2fk
DEMlj15lofzECzjWzgNN0KK5gsWWdh8zo8VLxYGsxC5pOcr/NyaIXaTmHAHr61MZraniEQxt2lmk
n6xYxIaXyuS8J/w6Go4M0sS7geu94xaftYItVZdD0XNG4bCRHPZxr8L9Ps+ZyWCSpq90R3SCf6H7
1OD0hf4w0L+quXsFece2RNnCOsLvGj9R9Z/81J7JyrYtLz5kFet0DYrCqbOIFk4frqaQmRhzDLV8
Rwl5f2eZP1aAfz6HNQtvvJuw3tA3tHHRhfm9R+MT55mjQyGZUyPv7jKC1peqjO2nMXwUA+tffdOW
/91Bs/nd24vrJKNiCoMCHhthDMzP576KmB/TgtdH0F4aWnQsoK5MojP3SAqz5yvveAHKIaWuW7rt
YBeA98PvfsfV4pNWwaVcwynK62iagEDdI3B5DRXlR71orCQB4oVWIojY4cQsNpCIDnEVvugsihAj
uFW9wNs6r4i37lWfaadDIjxfjwEybZQf2ewylzGXek/NjwfMRzuhAEfvhdrUFnpvQQY39IOnkNAh
AJ3kjUgXyXp/JtNGqM7YOHDDdj67K8eDkovHGsLjvBUiIe+yPMNZt3O2EpcyE1FJXOOoVGiEz851
scDHkob6uWh5OzXk6Sp5x6KLUwZ9kEZyrAn8vEvA6TOpo0UkFc2G3mV1sZKKscIg7sZI4B4aLcX1
vkFGwJ6NAqLdOsztC8XR742ZAB9dLBrt0hbRTnsGF7imfAIOAZYgY+BdjdocM3XNor2fQgF2fF8t
MjEQbA/BB6wW7m+ZhxNItUcMDLHRJKazNmWVINP1HIquShT+Xu+46rU692d6n+Z+4h4Nixsu7so7
TreUQ3HiW3bpEvJzf/s+13OwAia1AUuYkaSxpK47qWXmdJm4tRdGEvBEvmGStKIF4EHCXMZDXTM3
3tv6bApfYFTQ0E9PiFBurhlVSJnS2F4UTiWfcev8C3xaZzK3kN7/tAjsBBkGPxsIL6vCUYAaSarZ
QGuccwkXdeGZ/JTcrcCXqik7SULn+t/okN8ZK0/D5O1gk/rSGiUA4lQblanonULVVTpACmNgfGbu
VoOwfILUxbvNALi+zxMsf/8EsyrlAdN52TLhBioE9mMbql+OKMawmd1e+L9ORDRsoBXZ0wOltMjn
OqSDC0r9w3MiJ4sOWtXIOYY8PiU2ohJJQc0p2sB0tb8HAYuQdR0k6XAD5Azhw9+CzZ4t1SfSZBJR
m5J3Q9XO0EfJqqQLfIhlOMpHMSmRGhzCJW+PVi/RvpPpHdrCUZ9Ss0gdh6D7dKH5nZ/ttVOqwFbF
fhATTqLXvabGlYq3Vflm3QxIaYvKFvZEnO+uRV+KxpkPHg2yQjo1nGWsci21bpgcD8HIg61Uvztl
2TGlSdFv+LzAIlBKKDD9f0xxU534jF/Tb+yN/IW5Q82X2oe4ttno6vuvGCl7a+t19oLzUPLxMuZQ
sgfSGSmnZNQDSvAsMGl8/iBNSiCP4X8qfKh+imwthIrGbJO8TomqFmyitAofBNPQ8AXNUsG5yAhg
RBXEySggtAN85Qnvt+miO6mlNNSLI09ntTInhz0RGVPuIXACyYbL5whPjzvQYSSWCGU/2Tu0w2aJ
UH4XuGO0vZATC6J86/ZKiuPg69mMnIYj1uO1sdBtRgndueD0UaVN/P68xQwtoy9HShBttvtWu6rq
HpKfRRSzn6H1jFi0yekZ/6olqWC1r0xjI7p3kTpqbilrvgRu8FMBd/vMtfXFEQgMGW4Nqci0Ry2x
ADruIXg6orTT5J3FiSOSg0OHxfMzFB8atii1QtrgF9fXgugpj2AIYfuqy6lyE+Zo/O2OmnGaYkX8
40u5RfAF4OTekfEKrz73o9QaEz1fqZlLRdQTKQBRXO+hYZeiyczSX6E5ZyHTrdIY65cbu4bFkk59
izL+uI2tetAHlqNvEfjQk+OcoJ1eJ998nMhXGsHgEStwun2sxF+3SLe0XyxZAUEvju/Uw1r+t4/2
0yBWvr2bIgtKLwVg/PflmOq8dzP7IUULTy0kLkqB8T18xg1yk0p+nZu9wH8bzIqGUIGrH5IbVad3
knVDnypCUlxO+NsI1x08D+f+JEceDQSHm6l5cooKwK0S3/vO93QS5dyJRxQ/FOJqxsBKDHlMi8n3
OuY6l+6M5E+LgE2KC4MlihFf6QO1UhmOnbcALPoZBNK2rhurGPwpfYqgKRsHKdYNSXg/omXx62O+
VMTL/H+0RjwBKjz6eR1hYhee5Rg73EWttofFi08YtEEZ0dnQWW/du5q9cG98eiUcB+5KqJWLGhxR
U65SXj0r6ob3Qv24U1Fs2BMwBD6/iQpdRSxtfm95z+JrlSz0XjE6VpTfqvT1KLDapBvMD22/BCmi
/2MGG8PD6qbHX/iRzz0fonCwyxPpQg1txMBCNRtgpshXS2Il5CGCSfqGgB8NFS277rAq2meAgBMI
O/YcQjmofYZTuDZ5Rbbs3cDLVrbX9KoeIm0UuDxKpUH32aecdinmo0Zd3nKTQuDh/LoQgHFiLmJb
yRDpV1OBKAQd6ZmJEhXzPnjMBtfPh6rtTKmO9B+XksGqFBaeYPms66Z1Hb9UV1EPD/9XBnXrHGQB
qVojxYnn/1rc4hJFD8+iYB2JLTNLD5mxX+U1vrdulA2RDoRQvMpkMlEF09qXfiRdMmPDmpYLz6w9
l/8Xl+64By2XomHRSz5EazKJhxJwEFknDPGh16OqGlNcsEokbD11PAZWFbJGgvjNUOewGTmrNMrt
BYgye6gF/Nb9PYK6Yn6ngCZtn9yDrm7SwRXQv4gIRxPNlhJOPrn1oxWvlhYgOfkOYy4g6oiLNBuR
N68srBrQ+PfVfid+Yx+RvF2aPbNIZMmPkGD/+IZBRdBgmxTo7TkDOcxKK1f4ibVDELtag30sgc50
7E/bu9xRzYlcfTGgQTa49JH/Zu0rTnGnI4p+UNhzaXdH2w0emjKrFT/egwQ06lAH00lZs8wmmVB5
az4u+gFPI9cIdZ7NpM+UpmWHl4dE0xaSakxaDzVYOS4ZTTq5bLl8Nohsqb3tWwvYmDdstEzLVQAr
7X3c/ct/50+z2lkfdUF5nBikwoA85aubWGhhsv4qgJSWCc32l+llhN5EY84Z0S38o5H/FxErD4ou
KQh/JSkOinJJwMB05D2XeEcRbJ1GdXlUOqBrT0Oy3R+GN58Fo9O+4ABQaBTX5bTJ9dxOYXzo7Qm3
YCn+twB3RRqEpugOfbPNV368l4bWXK1OaN3NhOQjqPMitTE+WeLLMI96TCMbMsbUik+SS2IWlH+6
L/q9U7hF+FpJVWcYMgWtBhOfvwotR1Cw/0mz2DkkU2gxH6/4Fot/s2igRLEWATWMwLXMY3Yz7O1B
MSaiF6A1/c13Z39EeJDERufWAd8F1tBrsniYmQzcmS601QauE7juIw81emvH0s7+8amfm+h/3/ai
5tqqkPziIlIgBFB18Vfm3D8FUrEBdDSVan2P0/+6Gi7ivkCwZW4DcTX8HsDEBf5LPNCwepGgUU9l
8lAZPywfD3ePbnVZwuZk4JDBhynqmcV6UKNtQ7e5xbS3OaADrA4r8W9DdKlUohTxKITmOubsDcSy
C6UoGieHVnPIvWosqQJvS1keDlA0zBlrRXpmSN86M6uhdK80w3WSUvBFLtkvPK7qA+Q6M/nONgwA
S6HSk0n3c5mAf6yemRoc29UHuQPypujh26BgGhUK//MCv4bw1t8ycc/7/8M6F8SWVTNDSKA7ENdk
g9hJ13ZnuusORN+zB5xAS7/Eo5wPX2VQzN7L3zB8Qttmc3V4x62jqNTuVmybW0d/bbpMI/Ts0le3
SrXvQXSegOnnlmUABA94hEGFT6xjYDrdlE0li8R/6il/WQtDeb9BYIZanrln5RzBW7UUsG0RFTsC
KTG6p7oBu4fEPX8PNhUj64etYPLu/eiKmtJ99IFb41go3H5k84dPZJYkEL5q11Wu+O/gA7X104oc
tc3B7KsY3YyYTDho3stob4w/7CmmM3KNxQPLZBpMzKcw4Bfh9YmQAZ+rAcuuTfJzRh2afUGXCqGm
EO5WeFcoHBXPtjlwdGl36rYdVWnW8qScSG0Q6DzfYsLhlbl2y1bd0eqCH8HebrDiKnEJYBPgGHOT
PVgAH/TiuKjXcJovnQxSypsjHp8GL2mcRHxxEfJOfefP2YFcAFwYyacY/LPrIDmfpo39/Et4B9bv
VFfdM26dqvRi+vMuFt4pKyogmpQ69IYyQRZnlhpZP+EWrkqKeLSnvPEEZO4KLiiBEHwufWhdf/kY
0lPekVEYrWXDhjJ/ddaPN30tx5lfsxcoS3Hh3tgdc6X4O7lxKODXGsWqfI59/mElUuwwNl1aDsEQ
HQvYx7pq0e26wzZVZOccMcnkQnlIikpoCQOMnJKyo3sQR8qVSMf9Etzery6lrld6O/575DPa2KTi
W5Ol58L5MtITRUuHa2S9EJ6WWyV9beuXE46bSnOOXs2BqLZR5Q7Ed1ow+gwAh63UZ8B2fVZ7sTCG
pQ8w0tZFN7VSVpwr5DbAibJO/QgsJT0QcZbg8cPNGLOOb4Ug1djnWU4kg12D1pgRH7BX9vIA1X1m
8JoW07C102mLLbruYxrgYTz2bh4/3k7BgkhgZchTKSSAUy5wRZnH1FxCK9AUmNYED916d1e8dcd8
Sp0ntX2/q60YH5dn5O/HsBwk8bOtsIJpABL3KcsEdA5Yr8QSx1su1eu3BQRlIrgyDmePY9oaMw7x
iRxBkuBtqVPALJTlH7LXvWdHYgCisG2nm14dTsJwmWsIw3Vq1lzQFtwVcQoseomtDwDoEyw9rPGr
EIJg9GX6QBtKsXb/4bHP2aBHvi7TfX2zY09rW5WwkPVyg7IIrGQUby5JcbwrDOIyDDIjM/48YJBK
BB+Zp3v7L+3HUravza7YDtMZ7y0RSwQ1QiTufBQ6pKufG/2Ad5OQVFaVLOdU/KLvWNoB5tsS+OLZ
u55FcoIDYR479t/2XV4/G96F+oSomhnoNme0PLPg8kwwp0AJSBdBLKQC91FjUgQ6bwGTunMwtu24
tRUIlyZ0ozB1xjuvoDyTQSVjYyOoR2paYImQ8rA32FSmXbQduWBsGOw/dDmRI7/pqCE+hHXWQdn2
2mrm+dzfSigzaO89rTa9iH6zoDIggrRCv2zwrZnmBXJB4ONrHr5Y3F+NSAWgWlU5kofY7gujQP5I
EjbQVledQHhStD7ra9fUzLVHdNOu5cW2ndAEqQ8028B+DX+6xwz0H6rB4cwIhxXarothb87i9ruD
3nsozC8Q+s0CbVVKrxfA+0rsSbBstemDtjIFT0aPTV22SD/oVXRy7g1wxU+om+wWvW6M1N/oYzlD
lmAEwoZWxKfpLmPohJmeGSS+W09qexjmBanvBtnE/mOjDPmEN2XYbmuAu+8usBht184An73ccwTS
FAfVz1NQraYmXWPYe4pTH0hXdZjnskqdvGxKmr/Zw5ujCsOBXBXJGXJi5NpcnJtMXOk2uDBHCcQZ
ZTIvCI7ZoPCQzLIvThK7FOeMEWrclx/plkZxvUvgpLuc6PpyngwMQnQuF8HDks3vGz3M6G3rM15X
aUvdtizlkzGoXYWQZzJhFtGKLPvCekfVEOthnX1d/rT9rhvrvqaAhRyj1QsLM8R8ZC+Av85W2IwX
3teUekIc7UhfIwEqyUG3F13xoYWQ+dd7Ekt/M2unBD6usOKsw98lBAEsXKy1gsvl5eC6klDfc5dp
mnNGGOAyYAgN99ftoIx1wL5onOEXe0crSETu361eyYu8xtzCnEdm3mFzRqh4g/QeUrhEV4LF2cTs
Zo7ggx3uFSb+5X7qMKJzPHWCWDhJM9KhvwnHBom/GBj7dewvFJMtyGM4y70gRkgkqgrFdylEJlzT
dCd5vWc0xnE12N+OfuctxglF3mHh1BgtsRnDHgqXhwiQRoVIdm5CREIb4KVB59Q3m+EQ41FGOdjA
ycWmKtGSNGJHxioVU8MNuuREaNQVm/il0/aekT6XJQo8RMIw/wdN6Ho9NiWyExS5cgMBbiiUaxnG
L18UUIk1kzOH9LLjOIWBPoy+iBPTUEF0yj8fuNjbNkpxhLhz4mqF4ld02XGb7JaRafiQDKFGZ/Uo
`protect end_protected
