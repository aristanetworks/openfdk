--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
ZMURU7yNT2n/JBtja7/xnK2CmeHznyC8NWyEbaqrvMj2CuuwDEjZROEDUvBIp1VoUQWoRCWIRegg
WjJm053grUuS47uwyEHlNDv9SpIcOos7OUTaG/w/tPlruvBleWEU0sYZMbixS0heQWbJqHt1342C
18P2sZQ7wSNJwO9HR43AjSghxobn+7FFI15w1PJ8+Sz14uD5GjMUDQ7OnxpIYAkxqiCQtSaGHmhz
v/aQc2qBJRl4FTab+OMPoXPM3zX5N494HDGC/W3+0q6uXfKlOFX3FBTU9yAdo+b8aTiQdrFOoByN
KcGo4TWZp2l2qSz2kBwrLHANi1tKfK4P5BssbQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="rCVUgCAYD61fckEgglHi7/l4oimcQygr6afEDrpic0c="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
qQ4027cvZcYJyWKTDPdwFMua/PD+j0MiE1XfCO8QcyUrqcq8Q4x0biMckkvsZ8CIx3Sl7UASGehr
bfY5swgM4eaBq2+7e9WxvKQsE0y0VaN3VamMjOV8hzszEV6ZVKAJzWqi8Kqc8PF3Qgh1EAaRPOfX
b0WwnyUhA8RZcmyCSTgbBDmJxOu86jKSgDm/xnN/MhWYsjtpo0zLRQKvF51pl8cY/XbttOWgQueu
76qH8sLIKAJ0BBEs1QjsD/wFM2aaVhDIYZ6bGpl5x2wLsEcg9VXBqsydU+pn9f7coRjbGdD3mlFQ
PKIyZl2O8wrkv9xWFridj8mk7aAZuUChxpQYHQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="jjVaQa4vlX32uWlyu0swmIQY1/eZiZ8px/ourIrS6yI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21968)
`protect data_block
oHZyMz3UWZyt2vew72Nm18WblCiD861KNelOZsFxgnSaXzaA1CJeCXRlSDBcSsgV1Lvz2V2dY9jG
HCMxyzETsekVAcX/KP3mS5euGvyZQ1fbUxV142TFxbrmHES5wXC0yRPhQNLOkzXgrKQNQbQYVS+O
kdWNrErRwusuagVRSRxMR86l+VrycAaidr2ow+ZDmANtWhX4IBPJCpNg9lS/NDg83u/xHUFP3OXC
sB8NpN6T/MjSN3voXnoWecg2FgS4fd7JDS+1NMYIVkUUDGs3y0W7VMoAQGjec2dQSfrcghle5QKE
kLWoojlDAV7DinTmUFkX/Ac2RZA1du9v8nZKoxBoJPRuwxsNhsIaDVApBSjYs7AmGyxkj4yRCY7r
4YQtyTxVx5hzUGedDPvuEHiwVCoV17IdajjscflfR51+/xs04Hj8hY/UfcD0FJ71dhwSSuWE0hpR
ywYRPv3th28s1dVg7d/Ydb8RIrMD0PPmV9ssoMNB1RAwr83qjkeC9WSNffzjtv56K7uN5hG9WhAD
c6QHejEnMv3RpUHW0cZngY4jD2oSZ8N7LKDlzJhfi7YYnB0oAG10N2xcPe6S1eFAa4k0TZR8bHM3
/R1CowcdBy6a/ZTxnOmn4dVRZB432A2KnE1dwJ2WVF6B4hoy64MQA+NUKLkTOTOVynyNr5wCzIoN
zy7GBsuGmEceUIg0JRI6btfn2rtRCzwN2MvfB0NOr7Pr7nTblagSXMeZEX06xuSpUAPfwIxL1jx3
szUSqrpOmPe8MSjuf2VjunStYe8LjX12wSatRIf3u+dnsBn3Vbs+Shda1GB6pguqdL4Be4g+FP4H
Gdl6GfF8D1iKS8QqqDo7rTdsPilhHyAOMCKNIwMEHVvvnc3J84Fbv2obyg0ZuwLGaulri+iXmvvY
01n+J/SxQVY37UYHH6Q8SJJbaDRVIwAP0ilpm0RiwLBQpTZcDiuY9HJzI5jlAIthQ6JlD05a8nNw
/SiJrEJSM3ARDAcFX/UEojPA4hrnJsemasJscJeg5n0IkXkYaQUVx3DkHD6DDYQEFKXitpDbhTRt
snzj35Lw9hl1q9yQZnOTEiYFV2QPSwmGUXK5KOpq/DqLU5R/NTZ9EO3dKFSJtR/SH6CmESDlLxK1
Xd6uAIhXkUvOg8qqdAoX2hOTSMxDdvQNu6wj4ehfzINx7oLrL/GxoOLLreHZQz9hTFlF2bgzZ00e
oJHBHf6P8bWq1YnWxLWaQai1tYLnyX0kgpVFSvk8o9sGWNY9u3IbCYMb9pMZCsUshgDSpwewFWxZ
FpK7P6WCIowMgTL961oj0NVUyiuIuOA+fOzLpmNtvopokFCXyeyKwTZ8d2uK4bWfC0acamawQWyq
GoZOGTSF4esvFrbaNGryD6TS6yaFlNl8DFbtE/1jKjhlnWMV6AEZpkDOb8djFprxTyWQ2K1yMlVx
EME1MOmNUrtdW6vKePJHzV7uQrHadAbo3vLCpKfLip2W/FB7VNcojDEaP32e8WS9e8wIiAAc78Ve
nnPVW9gDr1GuBBGHvvvv0ua+zrCG7o0A5YfukYhvsx20l95Dkp2JG1v3cPkpN4hZpaVDnnQhgncy
q0hvskh9voO7EmCx85xV/hruEmrkTx6h7c0yLLA9TzBLZGcQRrub9ZWH90XNGqWDoyru+n467ejP
CoKvl3y3YQzrskakwAHZO6pgu9uraH9C1i0XWpWP45Brn9nny2pSIfQeDFvL3OW4CzgID6KubtL/
8Afx0FcvifPzqSGY3latOJk7d7cyXbzWh450gg6m04BGMsQ7JKmKrDPaEepmTEuOurn5SSYlRu4S
hhgjfwn/9tQYmHQ+d0C6wFcIlOsPY0Tqd16SHLYUUQKov2sx88BJs0U/X+Jl/YRWo3WYOGPa8JVj
CzjacdMb05Gk0HUEHd0sZp4lLNDW20DY9HBvPorRHa7n8IDxkzfYmtCPlgZKdR2DDL4vmchWKf0J
u3gA10dR80W6NJJT4t1jrQnvCm7S2lrktJjioWwzExeinxRibSWgJtxUO13A2qRHBQQYCRzZWNZW
72a4MKtqfvTwrPtSe7Uo88ayiq7VvTy+5hKYz/G3gD3uInyYyhEA05b4Skny0ygAb0WwGcG7uaV+
eSVIANsMqmkdclL2z8cIdXSt8GsLc3sAHetmPdF86G/SwEVqHD862QrrRbQfsXzDZ+jy37P1TDTE
0TRyTMev29hG2SolB9S+7jRRKlof4SVYE8ZNCTld4Mto/uM8vYAH1TU2KGje1iIj5O7IuV8q/Nnl
liQg71srN4pb9SzfV3PEPMn8fYNnRD0x5CRX63LxNuIZorhy/XBV2D13ZZs2FB3Tx3E3rMG328Wj
iAguy1WfKNPtPmB+msFFIBADIcclpociWKNfbaSPwmTfIOmRBhxv/ED7KAqV8va03PsTfkC2l0J6
oSteGposj6HEC6OCuQKu4hClnZq7ayPuolVY1eLzWfGouiRGkOmmgq5xXvUVgW33nvgBX//F5wEE
r/P5i2PRo0GFOyUrZhUgQKBGDmTtVbxpqELVRswT7Bo1gFQQZtZ3hdn4+vH1jttQ/Zb05svzKBZy
sPqweu4zkHB5B7RzZsbnYTK5C+4UzeV+6nFhzEl/kFsAyAJ4USMwJsKT6slSk1YXJVm6FhLhi7cl
YMuDpK9S4kns4HN7d+nNb36Hg7S9/Mz4VWtGrEcsZD2/fC5EMYovjjR5kjFAGCCF2ON4xP0iQavt
SdXjqUwmiD2RVf0H8SztrjynSQUkcwQm0VE5ELjtrGVyJZkO7zaevCLjfWJ0xYb43qhngNsmvKrk
FX+uzl53/jwE+E8xJJTUfta0Qevw/2a9CtJ6sajeJcF8VcM+rDUwXNf2PE1C5BbKMIaeaTQlcMro
cBMlOXATN5wohXowgWg0InLgb8zyvypHnx+fIBkdfGQb06mPOBLhFMotmo4xYtCJiFXlEAoZcPUE
xiqZg4XoD+RE3kHLub7zX/sCOxoog7UjP+mDg8lM8YifD23BT8/2EJyDsr99o6/RvxIzChjkI8PS
YbA2ltfyyRmUyKB1peUqIrOnLdFhMZU8DgNWu/F1PbOoghUTWF4p+eelAW2toFSMeb1vjBX8x7Nv
1iuDeXT1MW63fAGuwqjFJDWQZOEVBrr6dwV2XvERr7D8HuSpsWrPGiccFGIJdXMqt2g60PCe2mca
/IGQm5XA3EvNjk3UOgYimzL6QzTkVbkMk4XgJ8FpL1fFv9FrDgbaiRUI6DYzhrTOP+Q1JlxzeVIr
VcX78rnSRPF443DmsLVo5FZRDT74GTq6B/m3/gUqm1rOitnWPy7cAXr/+Wea23DVBS1CK1wMwE+m
TZbQ73koOC9o1x+SvJZp/jb/Rfp1d98njjFt3RV+g+3P8fP75IHtrQUn1CnOkBkRaBb0JK6QF3Ff
by0yHJkPN2c7PIQ43x30wnAy9LBGG78OmoFjU3Gy3SvxhLo/41v/MEgcxY8dBw65U9cadWsbrlJj
gmI7P1avSQCyevbcshtL9qO8B6yE4VIe02MZ7gvqujhjQojAqnO8rvJK+s9XLTHxmdpDFNLstPVA
5MujhE9NsXKUqtEuUHgcA2b+aKoCews6xVCz5NK9WfxplF4Y7nlO2QUUb8fG7TW9CZ45RuP8UpIF
c3Gc5nXLcxX6v6pDmSvYzbONBc8LTfia0Ldx2WAfJfm1/7XCfxF4j8l3snhOISVF2K70XSwZ3SIz
W6gIasGCSE51AYToWPBQGmRpz2thGPEVkr5dt0v92Z9piaYufVN2f3rsjxaAzJSkz162Su/35TrN
NmsUmvnAzID+4IESV41aVK6Lh1hCh0duhLfzRNhcu73wwm7xdy6d5Xtv+slOWWKKVuhk3OTcNlNO
VZA7sVDy+jXfztXeURSkHzUPZK5kT2NpwfsqYdMK+ThEmtG8Rnq61KxXPdzlR+yKiwJgc3C6CWZa
5KfwWiw3VJCS5GzbMr8bYnm0BwxjMY4BX+uPXHSjYrpb9gXYyfCbtg1MdimkJWQ8pXBK4WbdhBhh
TCCXbZg0D5Yzb+qU1/OAV3I6aum17FwM/2pIgtKqCWKeWKpgoQxxNtn67rJz+0CSORcLeg22f0J+
XiicDUV9TZLx4EJ6OcHk+k7Ct5fSlj/OpvZLrfsE3Qrx0r8NybfYOx05PNndAZPn6h4tQpe7+sMT
Qet1L72XIeA6mtOEnh/X1bfEeVDyoxnDxgTWtsQbDsD7+LoeTYcS1R1Gea1Dgk4vbpFtcpoFQu4h
s/6MgWSXfz8Qejv3Tp1CEAP6yEqPMecCDT762mkTsWh7+Ax3OhcWH5/cFaprxNGkyYyZI3GS4LAR
MB/J7aAhX8WT5qyg8sW9CswNWNJR4A+/IApo2w/O7l/S3DctC/d4SZQUHMoeNXvw24VcUKNwpLzv
blt6GiufIk/aLB/NHDErNMfjB0+fWbIdwfZ0e3vXho+kkYJ6ztkLtbv7+7cXsOaH3easv8QbTdHx
v0RXhLGSCvv+cKbIklPD9DRkQlj3eCQLoYf+iQRRvf4KnBH+FaoI6mMFh7G8tm6oYiqTGoxht28x
jVbG/bK0I8nAlf6OTFmccFjHkizI8ZeykPkrJz5gkyL9+bm7aJCl1tiILy1OuOrbkIS4bw9XvaJ7
eauHidff21RsyNfaLZ24OrheSzL6B+z85ZsxsqyxDeSWEcOunERQnNQ/3ZEZmyQom3sn+W6A2QnJ
UxnW27f7gxHnpR5fNxlLgsFK5S22tK52j+Z5EaTBMSOaDtHJ0o+b2yM+l5TT8hjADrOsHFhM8lic
ogN1Z+aRg8P8Vr1BeTv8IaR2x4xmS8d7IvcEKKeGYqpZHzjt51GUQ1UNYWJBFsGESffX4u/3ENkO
tcrAUqc7B/EmIBKH2IQZ0hMspLBkCUifuE5BidQAwqsaCL7wYdF00C/vAs4/nTPo6U8b3/lq0D5H
fA6Dk/QQPS2XJM/D1D6PoM/aqAVeGuheNZuTQ3Hh23qZgZWDVKwJsHXIfjdhL+Z18MgOG3uQhcWs
XV6dXLF0IJU/m4FYMxL/CyRxb6XG5qIvZWNZbW3obq9ysylLNBVgh7AuIMvkmT15ZWm7dhduY+PK
d5xgSMZW2sLpJSIeqd/Btj/10qy+B9KCPhyKyJ+rSgG7mRhBAOrN4Jtnu4LoxyhrSySLqrf4kRfS
8hp6Kwu14ayLc5lvJFsVVRvuC769Mf33Yl8cjBubkm5+G37vpiHV24WSmahjZVmhVNV/98gwVcH8
uiXaSei69j3fZTC5x+gEnGiNRdd7NXHEK3YN3/7DUGIjQAw8hQxbf7KKJKEqtuiZBRBRx+FRlf4A
dqNF5wiu5ER5VIwyPSXrPSs9qLCBEu28hZ5Y/FMAHr9VQJvnCxkWolsyZCgGVOYfu8pHzocQVnve
6WelmMWAGgL0aV184QdITtB1ZrMcJeH41iBJ4IoYBJZJnIjBCGOcFOZZOKrnTwqWtTgaXa4hzSNm
9J+eFSeXVLEWGRNQls/JlwD2jWVXkxjYEW3t7hkla/2HpBw5SshEL86iuBrPlB/eUIVWuuEt789f
m5o110+NsdsWXNtnrqBrdhDmeqKL8UZ9yG7bz9jHGeJi/hJnlQmgrBqgs8vSdqiL4L2epo1BH9sw
XJaFjQ5XTyM8GQ2toxjnohpU9l8I/y95UJO5pYX04QoYIvHpcqDfFAV/cRJQ4lgSJ7t33gI3Lu8N
HKKfmgt4MwVek9mistGN2esKMtSoXEYK7aQ2iYJU4I7KbCJn1va4M91VLwTEAP9CtFF0SUmxmAqc
5CP1YrUnj6YMMPVL3n4nhZWocPK+vpLFb5mmu/iWbZlZNbTsr5tKmzEbw1B9QC2vb261AjrxOFjp
FkAxwmLGKn38wPTOmwIocK5ngpdoUywlzpy1MwoYRTJtznHKJFFzf5rBo6dDZE26+dvRWgb+yTZM
a62DG5y9x+C3OeaiNiyIxhwU22Zc6sAWlDZJBgsFnRQ24zgiFeCHj2QOBzbKGKtqwUI20LzIcvMm
b27bUGoauxWR9zNPY6zA8Ym9FVV/G/rmlApo5sXAQHD2FQ0BKDjIBiCfaRWqQPsHrg+fSGWmQGvq
W2JGQsm7s8Y1iZt4H7EW7aVr975FuKVaFJQ21R4CGKjItSaMx0wn71GUKbwXvbrq61F9hZklzkHS
sO2uAdIAkaxd9LXszSNUlXjYEcwnoC4HUeBLpQI+2vkWTKdFB1zXr9KrS7WgGlp/6OylbSNdMj91
zbh2YST2aTMs3NdUUJt2tgfOIhqtTfTy8fhc9WNWm2UHmy/zPmE7SDrykRxEOYRd0rciJBfm+Uah
7VDqlKB0I7r/P95/uRv6KpDTk6EY2PUBCD4ve+xhyXX4oKtypl250LLrNiCd/KRWtV69VqSK+pWN
HHKRjMkh0kwIohuwlV4Ui1xiFc9tAbBd4p8k3mNuKNEcaof+bq1huzPF316DfrxSnc8loeCkS2Tx
FfsU9vdkRwYBrUefMPIR0fLJuH6pzh3coDgLiFwI0q0pww9mawF8YZcIdG6LA1XNoDrPHnFsGT1B
m0M7rHYAJfSxm7w+boN0dBV2C45BEBeycyG9Va3uJaZh3nhB6pVkLj1Z9i7K9qv9G7o687IW+pdH
d/N06nDA8mwIc+5hsFLZuKohT5BanlMRXv8Eh1GxXvsSdMq6wrVpKaGOSLTrty8WMnPwJ/CmW1dH
YURiEVzLNro09G9xBq4kH+1AGeqn/yecyP/X9/5CKganBQw6Ys3E7is9t4cyQJil/+Vdise9qLw5
7yrqp573tx99gUetn3a+Frk4PUO5u2/qRXZ30ebbleWsSRL8Kj02GOcMiBowqsvhclE+FiHr5f13
xwKfxTRu7i6x/M7GrPx15/ftyR4jz7AwKkG9uvNXzNdpivvLJ6qJ+yAeIcDV5+/j4pZRLfj+/zoF
pvcrsWZ6LQIXTo5jXCr86Wh1aG9YKPOOkOpeodQLZZMSJlccVIFhTXd3NR7kkIon7Q/Ko8VFkVph
RIs1zlUJXHqhaqU8XiE3Rlhy6se7gpihvgADvHD9DII3ua3axNb5L+mba9eB3C9N+mKWzazs0Ruo
f93ae1DiSgC9w/z+uLa/GNQrIVMc9vTNMlEFuG2ruRUwxhX03iFP9LOFXQj4xWIcNBcjLIVAVBtn
U7v54O0E2klQxT8U5RhVcTjc69fy6pPb324AHiYJFGEDWioZ312D1r3PiuaGoc6Vr5sO9BeTufE7
b9yx7clmd0KCt5Fu1ZYnCg10KcqkN7MsxCGbSmLQ4O/0Hn2lUdRa/xAsWjN9ES8wtZ8VarBapGzn
U2J8eUQXwsoEdwq3mBnLfg8ynA0Krt9fy3RsIhfRYTFwhKzh7YoiSkg89tvtrtmg35O7lEIh5ey2
Riz1/UPVTVmrQqaX9b4ki83Jh+5CFdQIE1l2nKHpFHriDMLS60QQh622P7li5XgMz18P4a3IjFR1
g30Ncq9RUeBVzi92WW0BuEeQuASCtBaHvR5gVSaBpTorpSfe6tqh7DUYD4PaPQhEtVLZ0VUw4fNd
2wqXKS3SWnQWlAqAFrxVVsJqatdiSdJpUDvePLbLBcWTiakr2kY5Y582ThntI7uydKLpcdxgTY2Y
HAWhP9NVWNCcP2fMrX2j1zlHjpoHnatA1DIUkthraFN4tzn2Kli9ZDuRjNMSkGWPUcWSU72dkfxm
VrAbx7GY/ye+fIcG6huKoBUuMlHU++1g4aKFBOOl/dqkzGEe0E9kkvqbayJoQkxZeBb84+/ALZri
UnEHaywdMBfJRVri6U7sfeLQd/2hdTHYzVmqgUAEnoVwF0qAgvn6ZjJsIUWp5ebGhFeIaLrrlBdW
52ZUUM4Et3IvTJNadu87hqVGiaCORszQ4u0LayqvZzh8qkeM2D+WWrNXLpSHw0Bc7YD5iNZtK+9I
nk5ffmOvRwQFbl6d+2IXy9DpK4jTwwThyYpYBsVWTO63fYlgFLKoY+qYABbbErSj0DmmtsapvyK6
R896JrlvMYFFqmlOgH89ZC+je8AQplqCnF3CcG3BL/uJbiD6nckXVQ86bQyT8byqInOI3T3WjOz1
8WFdrg8sjGPIdMf2Iz5IG+2k7+bZmR7+NS5GDwEG0KKkMFEEhyxlPF1/SXnyBkDp2WtOyktXVIqw
nTkIOiwPSPrTewh9iMN5Ft22qws0Dmx++ojXlKlqFdVXivv45vFYn7zmGQk60kWuEdTsv0G2ab5I
cZrNhVOIIm9ywJMYxdbXCBcEbNjIjE6/Bfz3+YQV2hifms83uUYjKK8CWsLzonAO0U60Yrgpkf8V
Z++zNJIRgEW+f5U3ZbbQCQ/C+cmqfYaZbAvYt9FQBYfHzpXI0JAb+rPsWmtyUEKiEFu+ZPYCEoUL
pPp7P9TJrI/lmHsK5giTCuWVo2PNJyMeGa1WpT9D3dqMRNfDrPhJTOb1KBHBuDS8rVvdkf/0ghdj
UOMCo1xATG9mgEibbI8okc69KV6SFg8ysA2nZWAbJYQovuieQ4yiF8hFuYwyY2g4afQLA4Z1EW/3
20obPWWW5mIj/y2vp6gC8Vr3UmR6HB6CmUJ0llwF9E+gWSIY2hUzt2sxZ/jHoXJQ1tr83Cb+gMQx
jS9oohlhQwKZjGacWpT+Lt5Y6MRw0ppqv3jilV0okyaTZSQZjt/ql4Rep2PQ8vJy1BW8ywNpgHUF
/Oe9XSFJ+2cacRE1P59xEEs2W/CaEvaU/9X5NmYO33B/QtIUqjiW/mXfzBRMKiA4EAORa08VAe+Y
JpzZT3YukP6zUgtYWZxikqFMAP8aCdPjN1NWfjDDkdAXoQoOqvYmH700owqtICBXSOquJDuybXWG
zx01Wp1Mrmwz+Wd0aE5OC7v7Ciflkb80OLSEt7Q3bxqhrfErQF8BcujvwwP9nzwEfXmUE5c3a7da
hBt08O5qGNta2CgzdP2MiWPjhh8CSOe3uPTnKIL1swFaAZkxasv/Tmyy0R1JTVzWx9yxilotESxj
lueq7C+jSxJUeV7bywhRXc4ZsBJXFhskACEbygQQGw+1Ggz1KaoPAb2REV3y0goh9gq9dIOaKaPm
26oOc8gfmaslxv3a/Fq02wIkrKZLw0sOcSVfFI6bHzj7yjqPSLWZymg/bDsZRmoW2Md0DUTuqMre
BgZ/dYexa9fW98jcTWZFneun4TOUC4zXT3RoFND9/VmKlCRZjWbUgD1sCzzoXzdyCudwbX7zel78
YpN31h8XTQzFju4Q9Tx9Wt/n6QP4WZ5bufEDskOm2rd+s1BridqbQDGUaslh0BCa1zELTPx8vYmI
zJbZHQphhphmQfXcmngw6qA664DmvA5yYVvkptnFdmWLBD7q/LfLfbbaOVDb3j6ENQXJEzBq8rJV
wh2j4hkIcBwcfXlWhjnafcvuuHolHwSREtqBYCcZB0rX1XYIqDOwXjmeAtgbuGAJDRNWGana3iJy
y2Q4og6Ufyk5/4DIDlezIGUdvgwUeH5UD0saiyoWSZv1Od4m3uBRMbxsraddMFaXfC4+viNkytoq
roP1y73O5q9HWjJHzFe20xiMT1dBP3CXpcAQ+05oliGSxyKtrCXS9ls0HODHEwoGZjOaUIdPemLE
siTtiW71z0Uen5+NAzQ/aUI71nqvXYrdmRWJOOqzKfkGuv17jf0zLkPSHlKbicgl9/h3LHmk8EyW
/13tuZmcoowEr8hBSfY7orcriBMo/S6Z96uxexWIa1L49nhpwMTiK9OymD2POKkINlx0BoJwh2BO
WgSJ+UBatE0U03qYcoD36yOBNJcyFtyzLmn71Ha5WoV4zkM2rMAHChmVGYE+YdTr2IYGN8zVxVNK
BoqCgizVPb9uCs7dwtuE00dyLlaDHv6TFiUfRj5mm9YjLFbMq1FGD4ExsZczQVHmOTEm01aIdeCE
gVu0BjhwGPDIB2BCrqUOjKvdiOuob2S6ZdUbs96q6EDKSvThmBryeeKibGOI2uH6NLpt27l34s19
xI/K9pvB6oSb7bwGA4HZ4GebBKlZ+C2uv8auakUncXz1ePX6gCpUrAgRcrhGngYR9yDmzYqcfoUl
e+t0mq0a/SoqLgaDgH7mrQfZWtMTLG4Agxlr9xX1jXkarKrLLZnOwxtwK1+HC5H2LSipADJpMrML
amGnY2rTd4GuY+8YHv2h/WZV7Jsrhb4ADDYQCPmVS4c7Cbu2E0BFIHy484JYwCx0+jdPcYqRZlkV
Iy5hSqXRpS3odse+LPN+fdiie9pX9HVfTVqVXwJojXZ4zjrwdh/7jbDJ+FMtjoACwJyTc75MfxJ4
bA3taNDR0IVuATxDwUxw33hNpKosOU9lu1q9ZwqD84moYvTQjF6oG7GJB3HByggbNQfSS7fKjm5y
TLsWpy68t2J5p/pstCpLykzn13izXBIQ+qMoFkSgMAMfdkG8WUm+2epHGJA3FwA49odjnFde+sVf
KeLdBKggO45/HEkqEdpapwktCwgOJPz7/ZbEmp7NCpoFShfSU7oVcWbh0Iep1YrNtZky6MYFQWXc
FIpisfReuvsjl35PJ2th3dvnCZsUfYUq5C3wxVEyYIfI3snnjrE27MEEb8QYnZAkvbRXVVS4P7Kq
qWVpSBrjcyLbLem6kPclJLs14yVObsdkxIS9NdYcUbitVKF/IFl9kcxKXlSBjPVskhZAjkEvk55G
qthnxnwzzJ/NUeGkF5MjESQVeH2M3DOkvbHU+IW8TUYrHYcOUc4pF/yyBCp+UKjxeHCOxKQNw6Iw
m5XSV7yu+5O6q4jsqaDYWWx6RW/Ft+hcHMv8Ji0rc0Bg840LZHsYUt1zVTGZRRd4qLagDu7PnAW8
So8HMmy/2t46BvGH1WRhNSl9IvtVb/IGNYxY50AmCB1lEpidKHuSUI3STEec9QeLSQl5yzSb0nsZ
Q0zJ9JPHd2pvurawiI6usdQitNycVNT6MKT7K0waPU2z7Bv7TjHk2lcBfeMbLd8Bhn0nZGuqd48e
zBvFF/lv5wBz9qZUjgDshRdl93j0MHvUpg24lSzG1cmq9r/+rW1juKQweyzc1Ho+O1hK2hzMzbs+
WKsOPTnzkacSdC97syL1uNzmYVB/V9XE54ZkMqLaMXXyCt0wuPn0aPU3HTH3Ya7S2MSG9fPe3iZ9
m46hhJ11jQOtWht9O1AcbySE8J1oJiDZfokcCmeJTpTVZc8dPvnam6I9R55Sn8X8QMU/VZUT7uM3
OdKfdYP4I4ixXTcRFR1d7+h0kg9/NB4PWF8cNVymF0kfeaZ/CYH/boTiUSsgU1cRhZ3q9Utj49FO
AFbzr5pCUxpX1NYHbz5WSRVS0tJFyzxqq6YNaSl04D91xy3Z2eQlU+ioUMFmqefz96Fs8c6aP8Ts
uPzNB4nr7PxQEjPQK78HI9I2Kk6jVvDnPoohAbKmsw21CO/6+d+hqQnQm/o6Sa45vlcQe93WQLez
ZqAjt+W0iWGYN5XIKWQyab+CMECG39vQCEn8oaIeCbDbdTP1JpJDwjy93S9pYRyPSo5tEOvUIlF8
CxZpQAj3dAuispnWEkduRa13zsFpBWPR/AIDEqi7zaDBKx1Ek2l9DxJviZrcC3/pLdtEYm+DIN1L
zUx3/cAdRXgO64IKRs0+Ko13/z9JVyfmtAjFzS6nUNxb/bRlxPXJg2znAsH9E0qJ3Zup5kuxV4T4
xzPrZWfBmVTXduqj3GrCFpcB/4txtDNH6f77ZkSDWbbueVy7NptxTg5MSDgqGyXDVnZY5aLIoeLJ
2x5tyaV3a9Hk+8sZpMZXIxM3gVCjAjtD/02sFaey0gC45dE9zHqmsOpUt/4QxP6wXZlw+puIlCKD
/M+vyjyx9y+lPqkAuUpO8Xj1e4HEUKvIqu8qdLOHGo/aw9+4/QCidzJzf3Gk6J5hLdP4pZq3YgPn
Vu2dULSDnSLw3Rzqa0s53oQJdX8R2NwoRYk0WplB61d/UZqGlkFsVoLLbFFe3NiLBKPoi8k79oa1
e2mkZhRTu7epyPKs2/+6dvM3gWsOxGsZwWsbia37eMrKe/EVaWeX9BhEZTzEQNjKg6D9QjDGiuho
N+y5xnPj/t2fFc+UyiVtC0EefGGrV+3y7diku5FtkSVb590PAWyZQ8EjCrzVab07mMhzKKWH/G3z
7xFJaU9KT5aXVi94PiLY0+Kv2YxSWsfoJWd8wrwUcbctEVNSKhg9zXgtZ7tFYIP+LwVT5oJNSmjE
N7hie4SMxS9Mj3U8PDo7a/J3AhKp245hDqOmJm3HzE29rMfM9GdHCkYv928x4gajJlhhS9+9WI8b
l6OCnVGhKeTXeQq3fnFC8MZbUnnSrBKw4NpSK69k6okL0HJVks9zwdkHkj//O2YF5/DTzkaFKsvM
8MBa1gVhRuwkqAxLbYUzDLXANZCUooCw+ePnJEfIutzfQE6jRKxlVj4CzTSyi3xODDsfygo801Na
uimWjJws6Z0e7S0ySWTbdSullzCkuZQLtOL6h8MxsvBlsgVMvRbIvpGkeN7fXMVl2NWt+qE917EQ
vMMAMm9v3RfOPtKXZ1fFXS914mX0o8HK1UWphksO/y5oOGE/Q7jk7mf1798SzoaOURcV3hodXMKo
P00NZFligNZbCZ2MtZa9Hb6Cs4xUdLR2O5Ct/tlIPLGuBULslArBto7Y8AIdiq7tzNbRHQ8NsfGL
WkvxwwZzuuZVg2levo7SEXBRIaNsMmmTqvCX5SFw55WT2Q/NGnMAYq+s4oys+QCXQqBr1JJxSasA
ULWFCKyiYoiil4thpZO7BCQvky3DmKPplHB0xYtoCYz++91SxcwEHiVy/YcceLD6Jr7jzkIbRaRY
Jv6Fx/YzLsSdc9B7jGVL50wHb3t+WFg4HWj8PjL1n9Q+hAhdNN6ycAzMx+NQfKteuzQwtDnFP1tW
+DbaOJ+zcciLHuswc1YBmerpXcm0wwUOxWXhHh/xLrZSnA7xYk0qY7BQbtEwbPVV0vZRARq+SzSE
0uea1Qclt6cwSud7mhYEkx5pYb8u5nfMzFEuoYnr7WyaREb54DGy0170bjPWvhrLgU+HbX4rY+c2
i+CM8Ghl2ChezumRK6u3QGgnMljd9x1Ag/Yhpg2dGWajswixdjoYxMfP+ROqUVbcf6SnRrKNFY1/
FJ3mh29DFtU55uAFuxUFbp8EW8rJkCKt4Iu6Se/HEVh22lT7JUjBilPHkCfNU7gH0gNGQwTkN2XS
wpvYiXppHSsx9nFq0JWF169WY54rbSn/s4PFLKWKbOa5Bq7wvlDnmY33bGkhGPV9nns8VrZU2/Fv
4uzKpJUx9P/8dioobL2GOWk6dG6doFjWqGRpevvYEG0NE80DoN1RCBq6eJ4xF+m1g7l6CyxPd/LL
vO4huQrfRgMdTt3CsH94KwgjJ2IwfBLgdrRiABteQyGil7RSnJeo36m2rwinlVNNN0jpVmMaRPPA
jyCnfOMagbbctm3CVIGqgKoN7CKSR2L6OdPa2He1yiK78xxK/loExePsJgUwBbNvH9gTfTB4Nmfv
kupCkogavKFQ5QlpwJjhjPU7RVkE20h1OPD+wxF0CqytzpH/CnGlPwFH6LLjXPlq/4aBZSVotf5a
AqlazfDtU08VJmzTKYzzWNVxnaTN27IGK39SuPk4vG5Ssf0qemEpdbW8ibI8Ca1GMzw374BzHbXC
vGFhaqSEcttCDIZqTFkyX0+mQPnUU71JbXuDDulGSZeBFP0Lb1A9bPLC9h5cuqnSJmP4Q0m+hx7t
WR9K0tCshu7SqAQ6HfbULSVOPKpmHiZ7nBHDeBuQrh6jyIvxjdB+z5Bd/6N/KEA/Yb1CxOIf2hc5
VOAMPbeGXpuxvzdBAfYHRtOYntyqNq8MY7Bn9YXlhvZn2qmGg/LiEQpRrDQn2UAFnl/lQfQjcLLO
lNdjSuNj3GstChqq1l4aoNm6IHfqLlmZ9OWbAcvhyECtyh7YLpu6jln1vKFGoalCokF+gqBnbTWM
jS40OCcykMGrYGw5gX9+1hcfBLazZ/b68KRJT2qWJC53xRtPYTEl+sYecapOSo+vNU9Yuk+H7+km
rtVQBB3swiyUTbF7rSJs7Ru1TmHCMTItp/W6CmzQ+C6pESPeRzKnmoE56fnFFYvyYTWONmg+7An1
59HpWiQKiVAEm+I3ESG4xfUSfyKTBZ6P8GK0cEypBUyBXjpqR6MFsb4W0iuejdAGW7waPTNBMv8s
tGNitNCRO/7/Z5Zn6xD3KpMn/Vq7zJlENlz2f/jHHIqR306EpzZlO074Z7fvprL2flQaoEqPnHS1
CI0lFzhASKlNoY+Wp8fP0EJqNEmg1qLfhNda19Gxy5dG6XsqiRPPa1XxUAiNDH9xS+7J/2kmvmYr
BK9QdR6C8w0MNLoko6leqDUzWSc2qnedYaN+eBdqhyn7v8JQwXhWnve/sZZj3m4v+bhxg/+3skU0
BxiHimlX3B0w6Vi7wOZCZMHDipS/fvsdBUvMWc9B8PO6H+s2mzm+ciI5545DeVOudOBFvurXc/p/
lkHAhnbmXXif/71HCbIkHdOjY507cRSvZaAU4G7h8tWD+EK2WvY0zDZ8JlJ4Du1VySL4EiiMt4JM
mJWI2Dc3PkpQqofKo7Kjr5vMsWy3Gwp4XNWasj+IQbWoHjNd4RWZzz+VgUKSZ1J92Oqd73bOIlpW
IdiU8WkG4r/6eXhzW9raXYf1pf69w1/RBx69/rXIMSB6Zrn05RnJDECvElO7rGR/m6G8Wd5mVLq4
7fp3/R4vR+p4Ecm3qy4bSetx/jPkybLjgace0Wn0eNrlswPZIB+louKGRpKDOeH3QSmbO8U+CNlO
paTMYgKapay8BPzhy5UX4zuPposm9AJjzyNzoiwz5ecxZiFrcFf4WkP8dXeOc7GUOm1Gm0S9uXfg
SAUkfWUNJHL+QTovELQqamCmn/UItwzA13QKZ/QlPw/A25lEtSx+YYERzNUKy/1ebp2Wvh6x6YWQ
e4D7c8Nid5aCl1Bfu/n4KiRZNreDdNr15avziDwK2aTZsg96EwOAlljPUM08nRKpan0dDc3o0Dqj
FP5SrBKCx0+cm29nRLxmWdjuZeqZPFcFH7OYMjitEnrt3eIOMD08qfUJ0kBaujfUmlxqYkpAKvWw
MMsiIeRq/sMlpNqJK8WzpWo0jGdO4QyWG7mW45tQMwOcYR+jTFwvirZ5eeW9GhXQOHH6n45IfyVb
n3aSE9izWV0xmb8ry3Ui6IXGfjhDh7yn+UpNllCWAAuXy+FONaArTMCqE2/Kh6GVCojJuTiCW3O9
lReM8kJd3Nql4uzb20B8pXwXo+yjxx02BwRNpXPdSVle7TtbwrDxdd1/uGDgBidDnRrys7R7IBXg
0k1k29LRyYA2/bf+G6FgU7S453TnFTGVo6djCuFxNQTzMr4YYyK+IugcajJVHtuoEvJM05rQeGqR
zvIrZ3firm0wO9A1N5eCNcMHyR0m9apqKfpkvRM5EOx1fBRLcSEKeNsxtLyk5e+TQJSTKrwTEvrR
EnzEA7w/Y/ivXRFyRhxwhZbG/m9/vmCe/UByfmychbyR8xsAANVJ67iLqUq64Cqucb/tZuXGnrSa
gyxKoMAfp6XF/IDM2OebSmVrxDEF5WOCpPNb1DQ7pwNwxPZmjp6FODwh6aU4H9H8MTqz7IMRrNgY
4fRzxH6s3wROwpjkNgZCgk0ZwMGffoxwZNUXSKbmiIA0urCepNPhBllIznvbZXtw2OXTy5Ux2ThR
xO562NVh/HYndky1dFZ0MM5m9ZYTQAHyopgFENHjl6Oe4+rQgMLn8ONV22II7AeoroBO4jQ6sBud
sY5y3O4+P2bPoaIqqicAn/48exSYXSebCdijoSmkLwlsZPe5ett1cMFClYMKR25H14SgB18ImU0F
SFGtXGUeJ9qIpHWqzbb0FX4JD0Ypq4HN6Hj3ewhHT4pfh85576rQpI+Olew08dfMxMp6y8a1CjDH
8hjihRN/uUOTzatnz/fLQJDDs5SIk6aROqVu5Czat2M5C2ypDGA2RMeI+bAubrW0EeXJYKJzSiQD
WjtI77p//+ie2vQcWkX2DgtV0H2s0R4GteKLClEMmYFXqRsWZXHZBsOctI8U6TAS28vStO3mL5hA
d/CpjaVlmZFncm5CB5RCQlAKUfrigznmOei08pRRuF95rbv4qBrPGVwlcXd9edBIrA2D59MgwuwN
DGexk/Gi4M9kbcnuwEU2jeqkyPsCiR6jch959XEn32TnaGL1TwqwvghH5K5uQU4rP0ZwYhvrN/MT
TRMF6a1S2PS6+vRtGv1T7VD2jJwbK3i1TQsiXDNLEDhrIIZd3urF/A4TSmFyb/JZJZl6H283LOdj
nHTcOBUsvRXsR6Rm/EchoH+U/w+3i8rpXqmKiOaZ/zuZVkewopw4pvjuGdJGpxATUQZwnHmaL30v
fOerRJ6zg4nr2NPpLHGs0tQa+4W+h02JXxkT4FxJur9TCqJavunZBsVEWMj27llG5IF74cEezIta
RBm79gM4pOL36UQusyaMohBIA1hrD3cfEZGCjM7iTj8HGpfRgxoxr701FwD2RUl5xgSnMSPEURi2
JqGyRCS6CnwGZPkuBlS4W1priMZEdUIRtvhTYk0cNfCwgcz6qRKT40Oh5b4mrc2ebtAWpiz/Wm+T
MoXUYOmG31dmJxX6UKBNUEv8mDPz1m33WxuVf2TW58KXByDkY5GMthnrVjY/+YcXvYMIHYFaF70n
xrcmnyGCQbNap6DZ8bUT5x0dbuncCCeSZVW3fY/rF0/YNGGTHn7B49EWdZ9FDO+QOWv5MrLZut11
i166sbZ+/FpSB89Y6LpyvecDDlfkESkO4nOjd9VDOxksJbippJ4p11AgkSfO1n+mpppY0ZO5Ngec
CZI6rdN+G+LjQoQF2r38zHk3POVqJPVgXQJeopEGWavO6aH5NwodSHGBzpeFGN7LTQ+b6cnn5+GE
yi99LXOVzfLLGrk1VUynAMwIwSAAqtktIXnfFxtH4o5Y31N6HwJZeRkgz1TzHopy3iBYaF1R39V4
bzgdStyjo21bZdLFFJqtTb9nJIhUELSbxfRsFuNLk/RkV9BTsLKDGWcRbPTFHW5flB1JvbL3prVJ
lU2ugW7fegSMMGk13jg1WIVWh/i98/9HrVBKXclHinkqQ5xP4HI7A2tyl/hmN9yV3T04GyYIIFop
PPumVC1+8FfblXt/MXHEK6zJpcs6qnWW8GMHixiSTRWxY2Avqzc/oR8pePqvso0jHx3gJunrpc7I
IP7JsSDF0RJdkw6YOlYaOHdrucDvFW9e0kZgJ4d7TuzQ1aTK7bMZvFRulV69yKuUtIem0zlxPnr1
mVlpWOY19L1OMG9EP6YdRxQciVog9YKzZGuMQs2R04cVo6qzi14LVVnb3/YU6ibHFvTJ6R51UUUa
ykTVrMDZ711xb81WugyaNsNMNgPgdKA2IKVq6DABUw89a3RhsFDnsBPAZQNMJ90TGYq49G/va1bS
hd62kZQ4wFFWciEMYDZQLOgdjzZ2pmq8JZf+Uf79ng6h3/aD7aGaRPjpO+FCVwj/npaxYWjSi0+w
1j3S0Q7LWWvLGXaXsOStpuIQmkmE1Fuw6WGA/VaDNT7+bL6ke751DP2YDoIaIMqFN39RMLLzjUg4
L+LuDjbR6GAvc2+YFLSbA6qu1w5T3b7xRxYRugXI8Gr2/pptNwzfuICKAtkh8ZJ72P7qVp5oqEL1
vuuqa9znBgYc8Wbg4vQdnbuhHuzyJAmoM9M3xrBQRuxScwRicYjfXHc0ou9QGJbv+zZjBfyx91GA
bnD9Yemkdjvc9K82aNYDVr5/3crVRyNlqdJ/gY5qe7Dz1zAGMgZL4ccE25Bl8/rs7oyAyIE5l1CC
6wDReUc62jtRdGwadr/eTV82DaJ28hPO1tGhP88wD6QK/JWehVcMENiWpoyFgtlyBFfOvvc/j3b2
W/TbJhjyGOtaYC8vH4sRj+DcMKqzG0F20eI5JgXT/wOAGXcOJWXIN5IV9fhZfzOqXz1zosXkA11o
iQPgB9e+J8SKTHuryoYVrIAJeKu4U7GOWCRKGKeYMmqZQCs7AACPo38vmQGu5RVsmIxGn8/ykYPS
Vbpn9UJwC+hBKCQDj9FPWhfYoTQygNvgyl2oZHQF6L7wVcEbh0Mu4JVgU+rMMfa5PbyrHgP9Cnf/
lpYCNjKT7I43OjPmGGC4QUIm2s3h4/+h8xhPkUeg5Vz99q+XJ8Ow7bUwaV2Ko1BZ0AhQz1arD/tQ
7T8KYqw63IeXXjCepKx3iCYfxWZ5D6sgmTvZtzfmcy2AohaEHzxN6d8cYFxXHTzJKYnGbU94eszR
MzbQqPZXaScH1XP9o5rELft5pEsL/aBAzOBeRELsV0FqQATp7Ea/hxmjqfcMEz0hHJupTNqbcyS8
Skd5LtCKTh6N6ECNc82sL+PWfV0AamZq5BEjvYqY52IvSq1f4NYsI1Q8+aPi0QdtI01i7edUwWcF
hxawj+fEca2dnBnDBwPBBk0uZzWc23oNyKUTdH73Q8fHg9FSOoYhSxdIya5c84ZFW4kOHgshWsaO
tTCym30M6N/Kq7V+L8XNCZ40Qc/tsHIrsEaXO1UkTF7umXiGQZJAZrdH4xbY4iPUwb9bWpeX3ixc
d9c7Ez+G9Rt9bHbXfUC3KkN+zHsALd9bStz95jxs1W/hJm6w8o9r7Q4aI8NYjewzg3AWpF/ZDe1Q
SK49tWeihtlkSAxRz7m8+VfXasP/r2kK+Nb/pF/mYmNVjU3XEAvpmtxQ5BtCZt9f9OW2DF4GbDN9
i1FZjq4sILlIgQKq+v3aG1FqANNdIdPfsl1nuVOIBzTapelOIMTfAYpk/UeigutJDo6OSBQI5tYF
X6SkVkPqIDq5VWvuqMlQb0vsKJnLIalEUQqiYVNHHAyEoKzMp887N+l0L6Rcp1hSUU/FLYHd8K9t
XJrXu9HXslXbAaJSkFK52FobYj4FBiFvgOu3H18MUcOZBxPFsbOGjN58Ih33L9jAoeVmtP/7CSWW
roRWTWbQ8Ce1N9xyO3Zb+TmLPzZot/7MeFuJS6HgGDl7RmT4KTE4AwR4OcTlTaWE9+yxc/qjx7YE
hUZVG0nXtQdbQnX3kgKznq3Fm5IvfMDa3FPnA9kqPDl2BJ/fo5LHQk24wBZ//q4itoDA79yxBDjA
MqguUVm8Zx0hAj2gKhPRN6sBAyAsSx71e1aXpL0NgZepPv011YZJrxX1u6OmEUnoyQtAKhryfBVw
VC3E2NIDcLcZMM9lXkTlFoG+qtenAhPK23WqNvPVyexFEmDS9PalVHflEEQhaszqqQzRgCYBI6WF
p80U5hR/K3v33MJkM/KUXON+/rfPtGkCvEhhtez4HoECyKzt9c+fhWXdgmY6z+Vp1sNRzZ9/ZwvF
ZAnLkIcjpXF5ivFAS7jslDxSapm5YHtgAMxtoCQOyvsjlIQEJ7+TDOWG5R9M+swyvMV4iaO5u630
culpYeTKxD+jJygYTCN1uGnCaStkLbGjjyul0iudp3xggR75nXQB6lf0UQCLjuvbI1Yi9KOyrAvQ
hEoJm254ftFqa+0TkXrh7ZvOXZCGwXiCcFZF9IMKHbk3n6AV6H/6B7alpmdt55gitBGDZBKXKfWy
wZDNkssjPiBpMuAeR4cbRUE4Wbvy2n/WMufuOIMudrFPhp7BH/yW9kvI2DouWWhHaaQTZS3rkpRx
NNdedoYFoPlGPKCkwnsF3vHgbGS8CupcYQC8HzK+tdfCEX7N14ktLx9m3ZUyUqfmKprTLBGLdCQc
RrFz71GltH8Jst8eP+NmKAKQGpcr/XzDfrkvfqb0OMaVy2PRyClVrB/owcmbtA0sT3ih7zy2eTJK
tmOceiBB0pog8zSToFvhnu0gwxpvY2r3shi69IVIeP4eMlUbUSBf3Y3/OYPFFr/yBiJ2RxBHlAim
f1PjwfdlWRq+t8uMIZXi2MHHxuUe7W0ZXAFla20ahPB1+CRvqTTt0dacWTN6VVCMTfTJOp8nc0zl
XbFs+34XcQIV3aWjvvxX+NllC3VL0syIB/zlE3etwBpHB3fW/VZ6zUOTz1CZ/fPGcuScne8SjoKD
PTVSJy99vcAcESEGBbyH9WoXSVXZ3Nyp6GNJa+Hs7ObVwkOM32Kzjx+H1ec8lo8fM7UA+CXKIt0K
GCH1fh0ceobU6LWnYNgbNHTdV9rtBzOZjvu6Ewd59a9/gaBGua9hT1PDfoUi0apl8HmMzjtj6ahu
BtjmispPorQMneqzo+jNGLjhbgJv+TggNPhbx6f5WtsRnDyLNkC4z/2qShgLHD5Z2kE8qiHM5gOC
uNyTvV43iK1x15BdqV5qb8E7v28p1yF06O7xngFsSjcTXtHiFVTtqBTXYckrgaG53k0rHKatWM2C
3dfQuuHJpdpd2Szjj6WxDo2w/5fP003mZg/yzZsq32O56liqPEHtW/FlwdlFK4g3SHy9kUwkbXBW
EpsbM7dkszdS+UWVdLdYivIAVo8Xz3JApy4lZB/0l6dD18pX+OGEKRHqdWYfuDu/9m5Zk7wxKESw
vtaRh8ndE6GatShlI5z6RmuWQ7LBBP/wTtu2lLzL/jfE175X/F/LgUWelEm1/TCXUTAbsi6Rc4Ji
TUeRLpvXJyz8XNxkuKyal03aB+pFrhzND/b25hDarDrvrlOvzg/HQwqlB6FohvJtxoefOpDHMLOH
kFKFNmpePKr72i1M/r+dWKcFjSCn6P1tWN+zeCFN0BrHyhM8F6OT+jeTuVp1aJB20WLDeWrDCY2A
YNis4HA86YYbn+g6AfPqzxPN4JmcBiTArsq/Uwc4U3qcWtswuPmNGnZR3KUXxVzeO2UCC/awSmQ+
JcN+Y1gPJSkqjkqS+43/cuHJORxgU8NYbpInNB0/LvJQQiHx3WBY0MYlEXY30BKPrjxP78LI5jPJ
OwJg8qjhyR17nD/xHa/F9tMPs2fvjfb8z9+9kOp/HU3tdL52zbzeCwIwwgvh7yF+4KX/HpBQ9VLI
PieQmbS4ZuaF5nDjQUrqxheMsm2GQQv08ZRsvvqcWV9lWIACRPL/bRAC8K4rF0gLrK1TnZ8fAp78
moQCBugkvf8j3wJHHuXIb8ZZqwtE4DARE+vPaTSqI/O/7ldNxXsVThnbJPiyKmSmHGb3csl6ZngL
Xto7skEoRL67M0uEQWbILmxt/NghBVnwnTLdc7RzxnmmiOS0lXTir1HLpxdmo3UmvGTiDxWjKJ/s
R5OB2iTiIMdUv8Pj3BUO1Uw5b1gHpa0Sz5adFmIZwsIYaNKVjc3KTXHoE9++sX82xi26VLtR4roT
sqW1CUyRW3LHQab4X83BjQQ1laTqGhQNg9Q24g+SWBj/DpRljwzONsg+FyjtamRiOGXN9gOuDaKS
ejAftEy6QklFZoI3E/hJYHyNTSBc8kMyIkHDHOH4fXmj+QMX8VWBBibDYUVp74vnPofFdEn+8jPZ
PnrhOg4M967tvmfDipe8NX13Ja9k2BnYaPQ0wg6KH7HBQr7YUgAJ2FAF0KFTfCh0vpS6JQ9F2XMc
KH6JqK2PJXnwneL/DhIRuKCGKt6mDEhSZC9ZgI99Nd2oE5J3Vbn4O4stEyJAq3i2GsiokmxvgIU2
fmY2KxOCENq9BNInBfhSeKZt1TSLocAeFWkV/lh6e4oqB9hXYt19J/cXre1s/P4pkd53FXKrr7uu
z00ZPfc6o05jixZwekduEcF4s5C9TBUMTkZH0DYdd+JhX4HJ9CIkuhZXl0Y1lQjz2JLg1Z7mg9T8
PT95vUNI3nklB/Yl/2VST087af3KqPlaQjWuRLRIq0jAvF17mKfVqqM7qg9cQPYySW0fVR8qXOvX
zjR6dN9diekx4dOJx5ijDtSaCuZD+K/j7YkHOiQnVUzc+JzzZlUrVuMLi+NrJ73dn8f+DcEgQimG
824I4Jps0nQa/j7ejLwOKMo3MtG61WjhywkFoFqFsCdN0X/0hCuyiRAw7XY3+rfUCjibVVS+xoM/
WXoFoc2GIG5lHAaP59d7RB9eIb8iupwIh2K6/ostE+8esbfrRYH6ID1yyKH2GCSxakdFcATnqayV
lw3UdLHQgDJ48HBbipZS4XPgpMv2igNPYT8grKIa5C7B5VeC2NBSLrqyD9EvenxK4QaS/ctgjqCI
a67z5SAYvkec0I7VgJl9C63z2vtssHrPmnzChWSnqbuNcr7N36DxpSoksrVw8kSRMX77RN+MT8ZE
faIkjM2VDn3eHZ4y6uIUPuqoj746myIA3YRcALwvrVJqMt3mJvSYs1JIWJoHYewH+KYS1giQ0z1B
6AeAcJlL/zrApesvdjONmwEi55Y700884DN576nA9xH8qYirfXwCZ5t9wowyIaJbE6xIfeKox+zp
zlKbXG2yUG3elUpAOtPvN3CXN5zhgNzc0MMVAFwWJ+nlb16UDOLhlOuNhthP84OAECXNvZ0wLr9R
9kgPhxzweXFc8od1YZRtGlwWHjIQML4VWrNW/gH7BApjqO6L0IL8WGfVyUnIbwGOniTcAYFvYShm
MqpF2xpy+Guo9jUbxlKRvUNnY0KeVXkVO18E5xfG3+stV5i0PmE9B8SVl9Ns8YqFlYYYU+VvL+fA
YaUO4XM3YgTv1zLyH6IZPzizfNPH8I8tOYprajuIV4MK4GmTT+48Q+0PpepRTFcHbdS6V1X0XhKF
MDhCcccgbJHnDcn4v/72jh4DUPoJQg+kOdiWkC6J0G9DBjYbwDmO8EWSlSr/N3z7044lrO5gNHBE
RVf9YVabr+WlqiNhoMdYgAaJE2RXUsBpXk0EYeyfeelX+IxuUJO3rToFxCALl8j5YONkY8WtOtHJ
rwGypnIGUrpjrMsjc3lfSrEfPZ3BHml0OFN1tn6oyC+V+foOUlAD33IvWY397gg2J4a3xLeQgqIQ
f1HzafpvXZSsWcaOclQoN7uG9oLVD5wvXbQBU9P8+PevdUuKqPPGWy3pu0JrBeaLw1EVykrInx6B
VYyH2u2fXT+HPwkjkQfXmzrxNtXDVUZc1Q/fgyUrb2hMUWFN12Hz0lKtTCwdiQvr36S0n0Cbu2P7
X+tnNlGBEYNL7q+mv6nad0OptPuyRcID8IuVI3XgEvhfAeHfLzQb989hvUlvVY/tazstZTUIJquS
W9UFHc+PtljoHTd0hk3ZtCI4rzjtzSI35vX/SjvmcFxQzHRQcwFvMhEJ5Belz3A6YN/ZewZhYHNz
fAMxESFUD9wonGhcPqAHSQkw2TChR54G4APi3HBM09qO0GdkgjaYfhtjrqBwJ5Kp8t6ttVS3Btr8
EyBpqoxM3dNsumD6gB2WQ986HCSeZcW/R9GOl36zffsPuM7dWGXIS9usqP7DpFwilAuzE7L4rxR9
DNH1f/SdmQCZI46V4jqOTebevBFEHbQujk8HX13IL+r17W4AFPty5SYSf/GRAFAI3kpRok8FfWjP
DQ5TRNbk1ihG1o0LWSHZcok0F6RJmLeolRBsgcSZgs3J0WKlczLCRfBTSwQ2FaYaZpid/WHhhsWR
67sWpwSX/kjW0A9WgIQE8i8tRWxNUwZr9rhIb/vBLJPE2LDVtK8nX6DJmoLzPmNHsUd6QVh4i5+5
VM9mgJ/xizD/1YRbRKSpPuVjH5Hbs9McoE2AkBmX4dNeFlXhHea5dqpTg1QfZq0gepEY4+frIcAC
s5AjxX5L6q0PRq1ndlnJ3NWD/OMqDkVjy8NRhoSFtXTHx+M2WcgMjP9+pAdiHq3BMAZim0y5QgTY
2yxaCQknBzZm6D1OvPo/5v2BlQTczROIvALlgbKtr2Uhs+jDfe+5lbHc2vpbfrqkQcbU6q94bUDt
P3QsFZ410lkh+A5B10iveDOOMZwCRdoMPLZnPVTKJkqlEr3IpMd5caO/Fs0xufZwXTDbN8jPWlcY
Ko1CrtzWUYhksbnk0RGX4ROTZpTaCqyAHcA+ilS7tsTFzODaQVtbeeF3MoIxSeIWFIPA4zkssQyn
gfG9X6/t1trdJmvwWFN9M50ivVY0DLInf2CNqdOu58vwW1CuR5XNEGFuGMF9lvAYX1OeopI0QwIi
caX9dAec+Lx1+Ed2wGDH7D23Y+LUGJUxpbWRY7VvOUX8yRnzziKE8LfxIIzpQ/KSXJu3+UG+M7D6
9D+CVBBOShQO1aVVqTfqdbNK1PKbwAsZBK/8uWcaHtz81h1ByGYTScPdjyssQjVLie/hCpFMgsa9
/mC1ExTl4fS0Z3RyREhMmLfT1e2RF2j152iwY6ARJ4/A6xAf3GPXTsUCzFYbnyFnToeRrGZgwNAF
MZJ/vSGHd1MLF9OYjagOVq2rWi3HndzegdlvtWZ72LOyDkUzy1q3AtRpQO1+81pJxhyBKRAbcaC3
OGxvUN47drKoKSHpQCUDswL68by75/yWC6Lm6NgtMk+Mww73omAQrAlJsYB+cyu1NgyI0D4uQZR7
VCmslzzVc4UpkFTWiSlBZeQh3PYpqMaeyfFCUpZjmaTFDvtFi8Xh6Sq76vjEsR1nNlm3RtYcZuNi
5HQCDX6j/5545AcI16E8ef22KMXlAUV4K3fX3a7reYkX+SMnFhLWm2IehZtG/MVSLQ86QkwaAjF8
qNqkMGwLh0TgCvNczRufbX2+dnljbBl2C6iWnA2YRkpYJzM7eSm7yfGgieVQVPX38WFDYmGzMgsT
zzBRa6RGBOe8jeE261hI7eZ0C4UoT68Il3QNM0JYZOZ+w0NWGpLHAs4xFc3SIhrWOrqi2PRX0Cjm
IIF6bWMS+p31z5Lq5shS3G+no0WrBYQkaybDFmAKH49cPdTMm/9VOTpQGM/3IrWDRraRfR2Plf9K
cM7RIi2uVMJD9ktKiPqL+FPcll4MIdecz6Bs0L/48M919hxkNTt2TJI4K+4ojqxvVi/dJDGdP0Aj
1DU+zzV3aAwqFn83MZkxx7JKzex/+WsCWIupez9f7SLhli/oC/s1tQxu9NWQHf/IsqtDkMH9QcgK
Si3ENLoXljXvGnnU+fXF5mNw1Mkt/htTcMo3kII3AwtuojEjwIfyG6AmkmL46I+7mIDERT9NFWIS
UWWMcwpsQyiMx66jXsal1UfGLIrDSZbLPtRAVsHouPEc0gTfFcO609FNpsM0lNlOtIB33L4OS9fb
BSr2iDTvxUNf0VV1Ho8bg5+7TP2kvT9KlQBS26/HfJjwMeOwNaIL9Y8zzbUZ1kcFgsMUr9lI0CdF
R+Z/JFnO3w6Lq6F6kjN80yCuQD5didbbRyQ71ab5xBkzBkgSsHkRbyh6DSO+sNJvTUI0+12HaBqJ
ITNVYnXzMUucP1CQDSqT/3HSi+VNGMVlKIvevxGDNy+RCLTi0wAuj1Qpoo/Ar3gnZeLvr4psEOCO
88/ZMKPKol7vzdSPNCb3WIUcxpNfGtd7q5WCUcWEZUbKul/zLcIdGplsvEVVo7sk2oQXObeYWpr8
cvpzoIfTo1MjsrWeaBhgG7NnQLcTuDFHFnq49fDtRgIdnHNOCHWyRH2jogVTAm8OYFjg8LwISxFx
v7XZgdPZICvRO+z4KuR986IPPm79kdAJmSnH1GoibrHJpnwEP0LzXRx1g1x5dWapQG2V+99Tqyyi
FY01dgp5tNoDW4/Emg5U3UMyoHKIhEJY+9vKPjWvSlJw2blry0o4LC2Iy3Qh4nNHRsEHYsGOm3/e
mh8Cqc+xLa+ScuTo+ThG4wz2NJe7WWrvzQS1X7lXaq3EWQIGuNVSOt+p65sh4eXHvrgTyZH8Q7+R
qbNxk5nPVjCe41j5PGsFK8Dup8kGjXRCZwYhAqCwKLM0rxtrd5z24fdRi0tnWwOhhcBx32wjkRZa
1e6Gt7PVKtdu0NvrdnPPspncgLi9IRakGE8AVejMfqnRuO6fZdQuJObpn9HuGp+URlllq+z9EuUr
RQTVHPcS37yIHfkAetcLgHx/HIni7ff63YUpgKzyJNVrY+vvUPzEqn153eGTxcMS1UgxSSfNUdpt
SZlGRltkbaKA9oE/EgX8O7wVILUrsH7OUDDFhOmjJbEeu8+jVqu2TtBxeVUZPwPU4U9c/XnqaQID
NrKIGgISJEDpBHPPpHd2j8J9e6bHc2TaZq5hxYnYkvyfyXm8C+y5VQt86BGlOtBPtZOCLF4WENwC
+WXIgnEZ/tW25IoMxZl59PK9DRMhMznFQhCVT6rKWfKdxgasLhGTmp3wb69Per0IoT3xSlw7etBB
CDLBEMN5WvFmgMw/t5aUwZROyS3/sYCTQl5mh0Ooe8qsxJm0LXc9ATBKzQkY/C0n2vibyRGdiN5b
FLmNGovshMZABq4EFiPdcnYaVLPhtZliDWkClFuXnisl7Ni9ekvTHPr7kESWY+TRSzu1kMfIns2N
nUsckwthvji1bULZ0/pWZz1LBW+4R93rCvVSRZtmObZlPIst+QbrxvUnND7p5PAfLVBeHyVh+Fwi
eOxUA1P+X/rBRL+KW1zv3ADGc5uOdbCrHePBxXlHlaRB3wbf+8NxnWDTEIZ3WwGk4lI1CozPVdk/
qFn/7Kt6h7ycfxKrje1m6QD1H6LmDp97fA/b5Oqe6pZQaxx/S9KqFG/xkSGaOPrY8UPotJ2O8hrr
xqNYXHC1N6d3BP74uwf4koenLY/QwVN1itj86fJly6AhtZ9r0fKFNd9e5tZXEazQ2q0wQUCqkG+v
7zjGwrslg3CS/txE/urQWZhhJYTvt0YnVElYypiTP3gLVw1hSKVZaA/OPG087UP62PzMK4pp6ie/
QDBy7tPGVfau7eoyBXDn+8lry1zXEakJowUvBQcPfcV1okXtbmyvu0nPKNgpmAjH+QPinkm5Djjn
BYN7LJTwoG+NmG7WvjdAGNSc6w71pF7u+KnWWqFZpv3L6XNcQ+d4EORy9pXRcFBv2xWMCm790uGm
UZ6pS5KST/g75/1jfLX+/P8Oj3ZGpD6h4RkcpaK+6KG8ZwrMZyW1Z+1kKT0AK6GWDQ6IOt/Pjjl2
y7eVI5PEuIIcNROhIQJsdp+7U8qChQWQ4isWid2vqBgv1hfB1DCKJbB7Al/p0Y9oOQGsHIuMh8mT
2eJyTfdPR1OYeRaksLK6mdjuUBmDMCleFrJpOe51AYZ1MrK2VWbrORgIgypoVMQph9hkXDqm4I4a
Seh0w/eNqQ5B3rGv6bPgo9D71csNhYFK3IU0gD3moBPNjbgOURutjAuqfZHO4gN/5GEy7mxHdl1B
AEC4S79lfkAfxMTJ+gaRLFXs6+rI4O9uSlGY0gkgoCcHMj4hEOuXNrfuAHdSBuDDnEfLeMQfEhpB
1iTQDGM8C//89RaFGgxKMhWly2qKqyQfUVUSMd7sg3CRtE7a87kT3KLvDpKZ9grp0cXuoPW1+AHC
sWkOh36lDWksewqjr9yU8jjcizGs711mH3WPkYmtOEc0ne6pQFQvQxXqxixUU9vQFjfM2EMFxUwl
cEYt0TxC+TaM2c+jQhA4GWHrsbvfiNW9mdjGHYZjhz+24knZinKDXGIR0HdXEzltsbhPUsaRDr0w
r1+r3mlE318M8QtnzJJmmGCRiNF+nza5o3VXgaBfEb+216yIm+K/BfaRKC3raHR2ZKYNdwa6YobW
Ntgl2q1LpHw9LXD0VpvsLPvsVnqoeEeVXhR8EM9iXVGSoXEAcOX+d9qR44ARK8U3E9H1rrdaqWqs
EpxYgYJYuMrkMBjxTC0ThQJl30JSnAyCgyp+fWggTOVWfE+ySBZvPhZ9r+JMlNPYyhWIvB2OtM4z
8vvVNXIhWeVqnQ7SuKVCVJ1OaX3AJvdGoRPHdUVk43U7Sw2snVklZMuWylo+rBa5lrfVp0r14hVB
RD6OHuIq6E55ph/e3PpUoczR1aKaz8DO99B8Sn2G52d/ryM9NxO10MnQ65ULvbYCa+Vvc79QYoyh
rKmNpoVDt7cQ6mBZLEkKSBpodW9DAibtXa0wj3iXurUf7Fal98hiDq+SzSRoNrcMZFnI0g2Rem/0
CcHHps0VLSwwgBZ64KBjJgmNS5Q25J60MLH59nanqnezu3iwEif7TaWITTEo7m/PMbLH/j3KSmfF
QcjA9fhCDHAn5zdksokjmiwJyY3GQKgtDjgMeqBggqJZUIQbOMkxcZaVkjAlxZmcRjLXmRu2OzWU
D20mOrO3cO/Su5ZHMxJTW8w/tzUl5i662qfNlxc9QyKKb3I0LQOauz950oeuse3rkF5DAK20Ek+q
Bsan3jUgvxfV2qzWA4vCuyseh9EfJAWF/gi2llCQPiNSKlosjCl0ArziFWDxNkYhT1XQJXBlFqLX
SCLPiWSqxMDESA4R1AkbEX7mqY4HgU8otth71uwuH4CQC1hIv5dwby/kFDKBmYCCN1r3ZoVdQnZK
VsBy1+7Oga76vLkfCEjE0uurTM5iYPqv+aR4y6RVQjWXQOy3ubeCnRtZ95Y+z21S95uQ9uqiJaIs
Z6Lw9xY6plCTDsTH+gWokNnIjxvafB8fr6HNJWpVHGXeZo4Gv/GTbuWPVNqxvzfiXTwIo76RNgfR
1T3qYwCg3wuZ3zGgxYTQqzaQFyXrtnAJWjGEsV2x7uEsAx3saA02WFiRzUOgdYgSibLRQEwwSsZm
8MblnIBRTbykqsVN2K84tQ/gpR5CMrw/tE1sZIh/fpqakIxrfbbbCUb9shu9AfxB3exFVszwxZYK
9uKyE13aVqsknxiE9fDXeFPsr8v9WEvERnSSExjkXrGoWyxEgqUkYbq3XeI8QUb0lgCbwxn9FG7M
fP8ttfSRH5UEdLy9YsOfSASy4eryjjAtjY/xYYsw2BN+ixTzjwgtJ+EAKEWbHA9A5PaHTQrP4pbF
VYrYYeVZF5H+Plr4Gdv4kkK0Nj6k4jui0RCNhPQigi+JwuGCnclXo2dEMcIrVZ1sAJ60ex3PpTXn
1dvSmApviKHSWpLfSJGdBac3ASy27Q1tMpHYk6aoYOY+dKnRMhAU4hR9DXWfN2JkazeqeiCTHqdO
eKqOSszd2dK8VkRDGfbzFn2hvaAJIqau+CDhL2pMIZO/udGzlhuJFW4VQMh9cdKSFyrtE6ey59yo
1qkZ0yBDIq/c4Jjl60Kb29eHO4rlPKZHG18oM7fYhE8ptbYsjgw3LyOzr9ohYal1SvjH6FqNCjzX
sLYFADyk8LdTy3uXN1q8gzjY0ybOSCdHsgglIVY5ssymIUfeE04jBJNky3MLMdAj0XDIj/LW0v4t
TO2M8hxQrwc2mL8tNgbt2J1NucjzoZ4ppjKQB128WSGRS5A/1OXg8zLp27sHkQGwKpOcjCHbHD5C
igqZZ6MMvQ6ZwkCQEdm4lZsRKD1JA+B/ktn/NaoMsxcR0los0sD2E6EUaVwOxAmexkeC5L9p82pr
PDRDqsL7yfeiJwPczE27hyQU+9vgBfuht2/Yv53bUE70qsOf4k/S3sie2wUfSAJtJzmQEphme3GD
NT3H1g89nUPmBkHRhEslSQlR1g7O/rc=
`protect end_protected
