--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Pb5f5BBkLTlG/YEoezhTkUCnapNzx98kq83m0cxMvPWC6QmfwIrewAdVMVCcgV/7hHyg85RAFLoC
C82EcnY3JqqjBXmyW489DGf0QR+d36amQiY66a/R+YgNcc1J8l4OnXnNBG+tjaeuamlh/KE+bKQu
jI0gzOTyGgV7Rbvdph9xlHCSQZ8+Q0QP9qAQ5PPDgwfSkRNhisFTYyaFE9yumwUPMHpVVKsgXG3G
KYYnB6aRwxNpcQRS3qxIYx5bTexSMscAbT5BELoe7zj9f56KRyqafBk4SDd+WqsyIZLgdwUfH6EB
5neh/K4tAmI1SIiQvnSZzp2iqVKcRdo+B7ebow==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="/Q7mPQdjtCN6HQFtcG/GCgyzuDBzAnY1koS3Ek/bHcg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
d5aNlA3bk+z+lNCGyLGIgVNxPGwHGVAm5hYXQ7/9lViV+5pZPdEI3bLT8aAyTkjItsUPw47DUhne
KbF63yuz/yGlOJGfdtqXK2irFMT1ws37U1k6boBaEB3xycBhXc7UJA8Ypjpw3c4umOeta1d5g0Qq
ns1z1gySCKYP1Aw0bTIO6//m5eB7/nrNKf3ErQxedtvomPjfbZuLyVSQJXWHFhjdBmByWyOn5T0X
R/H96if/LdI/UBo3p0AF3sHCbprG4m3thcMvolvKv5qVmzckmRlso7h9YVIISCpmnOlketzroWt7
aevT3C+79ho4jFaECJSDDIzOdLiiydrOnVg3UA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="x2mV/5nl8DFWqoqeWecwLlB8ZS4IRuj5RpvZQDHK1bE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2480)
`protect data_block
4U+K15W2cRkxTa745/5Pqn7j7MCq/v73TG69XJslfyL5YiZW1PVMUUUJK0TTw5748bSMIrdRSTZx
JGMpwWGWPozHHcNwZR7dKmA9Q1VALRwALRM/ovUM7uD0S0lw2N4nUGCKn4F8QU2Bavlcmy5HSd71
Ufj5P7gKoz41hI36Lkm+JeCheK/3Zn5HMVSy1deFO3lBn4oxHLjMs8LYcSR04uh8rYC84rCof4wb
rFD2xcKLecQP1iCpr3sTVjflcpe28NnPorKpawz2NilKoy1LNGWoQSYCXuCGQ9B69vdwUrdm99p1
jyN/dyCbbpej1MvF4KwKrucIo7giAFPmen5UBOfGRF/oBw87SCePqfec/TN1nVhycXzgFwndotXR
FqIdJ/UE03ESuMzdBr3PquXOdyEIGAZWmv4TX0hjHm+BoFC0R6U9+J+HNUtJp5Yg8qpDkH9EbB88
LwbvDoyP+Hq2rXLUCAE+rOqJgMqJ/fdnlqUythVmK2EuDnHxmyKor5b2+GhZQKio3fW3bKKhPi/z
zfrhEertmXt06OnO90siV3W0+EPAWyhSUMP+bTmmKIrW7lIxX4YbftIqjaqU4dbN+T3Udce/Z8Hp
QuPTygRnUGNOcmyjJ6UEEmw8XilXb/bD2i95MK00x83DdWTmtobp8ZD9fjiH5JsDuXYCtOiq0V/5
a2M5QgDespbNjpuUzn0wMroE17z4E4Efcwc70IIrQP4BvZIiRxpuhaWEb2Q7CZa0KdK6SMv+cW+S
B09gpH6wQ7HxuSoDa6y7726UecgYu/OtD+khZS1NLLiS6nYD345NV7AErncRlKbYWQ49ryNn/0/D
1GPfofYGAighWApcDtiW+xcqc7aBQGZwiKWHEPfoov+GErpSLTjF2/2aVTL+ZRb/R65/FkNZ65Du
Iv9rlGiOQPIWlrb1vQvk68D1M07uRHZi0d7iTOUUcAFlaRVXk8Qr4A6fpNLm8wphpG84EMlEiaXm
651UOhHplAUQMfK9i1XsIjf2lIrvtjwq5zmN+9OQz5eZmOOvBTWygGWJXJo8MYbGVLJMPv+3QwzQ
KctE0QU1vsfmQ+stoEJD54Ie/+50URyogDpRlAglXepQyqK0iwTGfcjuKt5hyIe2kC5T+gc699uo
6TUub1JPU2dght3JIypLugCwWcPWffFM6tlLATj++8HQDNbeIpyaC6M9oobTAn89Axmc6XCs1zZG
LBd5hwPiOS7Ie80sYu9xYZPLofaPvicSNzWU0pizJ1DHQFnUjPO6v3AIFiNyB4IvuxcMxEA7JQnM
sw/pthJ7vsnJd+/BMLtJf8Mh/GmWqrJocmggX1Se+UBsBBGU574hzVkSwchCK7pADaed50XzKyR/
HgU3LGI18Uzs9sTk7aNnPB4AJuNkbkxB7gVsXZeU8lkuPJ3WgZvspMlVu6fABhgcEqdM3/19BTVg
RwniNREYDlNrVRjlmEFkrkOMwHwaZuKrpHgzq2ZJtEmmv2BzM8iJ79Kl62Pbbrfi0Bg1Flqkq1Ie
bECk3fMb8jZ2ZsPKsHuWMqxOSB/Ho0W2GQBUFBDRcOw1uhqWKhjtZVbj2YoaTcem4evoaihu4NEf
6ToizSZQbD4+RJNB3cXae6eBrU9ZFoFeIK57d7rBwBgfKeQIcoLOmQI4G1D6yNBmAB47419AIvXv
0gz182ls8zG2YLR5u1UiGoVEE852jfG7nM6x8VGctjEYPUcJ2c0oYH3xgtGTAACQM3Pesmmb9c9L
YQ/f+k7h2Jv8vYeM7BK+aC0suhITQL+23rfG50vJ1LFnUovYkx2mIjpHtA7n1bPE8NM7Fhr7jspk
zx/hOIWB85atKAyGzsGbtzX/drv0VdN/AOaENaXcMCTOmz9OnuXp1vfWs/Ljub3Fs9np/8iXwmP5
RW3/NI6UMOe7c80/phMSo4SsbwbTrXu0dSOY7PkPxR1OkonxzWwH+Yi/VbcJTbtMQ5Y3Duzkov5V
lLC1r553lw2x299YJTzKQlSD69Ty8f0Or6ncKqV+tEmNzn55PCFAjLfWO8dDqOh0WdmcgqryQkQp
312PGz80Mi2F1NIF/asJlSQFXO6BFdfzCNinMrHmIv/IcaGOQYK2un1GtQpxLKSjFWJ6xl8zPqlO
iH5o/ctwaB1Nsqd6j5Dmpm9t+/jTXG7q26xAz51M1UXavi+ppi433D2/Y1TmKFKh6zHQ5wNBpRhe
aIha0nPX19GyNSl3bQ/ctS/NANfDfVHLcEbJ61TxULVKkS4rZ7kDz+SvaRDk0rES3K9YBvZCHRKF
fjWK31UQOv2cFoBV3X4Td2aunf15Y6I/GRDyMDXD9n/5oBiykUAzYgrRDvb0l0QU96nBHc/ueP8M
veRIdwfPOgT3shJrYicilE5AgS8Zv83eB30nWSxXjhU1snz2OG5e7hS++JfgTDTre3eWQyw3AVBb
+1gwHKnIsAQ26lghCrd/Mqv3x9732kNV/VUEo38iz/O2lvA9p2RqGzZYvthAVgaTVwFwSXQ/HInJ
KviK9ApOlERBqjZDX5oekzRangDZE0E+9i+C1I3/7giW8QklgsrLb/0fJQf+XdTM4xbqnk47+YNa
zH4rN/V2NNEKWkVuZsbXvzzwP3JT+qJLpN9d1y2AjkG4Lk/vKm7f0djCqQEtC/Z7o4HWr90OEd9p
vdYLs3JzCHdjQnp3NVuWc4Pk9Z9Et1K48NkHIWshrhFKQsuwIiheWL9ncqBhM8j61joW83QiOptA
FRjJ7Ffd4PGu98I6i4qu306An6VIK+HR/QvjVDelZAzqlohiGB2mZ3ImhzAt/wzCwD7+N9wNISoP
ixevIpnq8s5eoI5fwSwN+i2M4f4Rqopg7dndna+4nFYatoNW9HRJS88fsioTHuK/RVgcPeBfowFK
QwqpIpZpsO7PouixGdpHKSPXj9juavL+CdwwvsHtQSWbleIZeIkZocNwuaB4uaX5eOMagwel4ZQ2
CQ/WpUhom8uenpmWlnhVnCkHG6n5o4KlFGF7hUxBipUARg/Kd40heOBON5nHNWnD9NezSNMi275f
RfPOfrl03n5VbR4M2jeVzKxdrx5uBdq4U7EQyK9vdFRcxxgKCL3V2W8VVW3LwUEFaBa+giNPCnhV
o59i1kJw8encUE3D7LYlp7GBpwtB6qcl72eu9Hd1CB1cHx20MN/ayaMvCMzAEXndg67Vcyte0wNO
9S5kX+l0MOlXDgiQ/ly3C1K+1IWPuCIRkKPPKXSaDlmLdzvZlIAmCJPF7UUTbuPdmmfQdxcOtUAu
AesckJEyjfxyuiIMwfjIzXLkNewNE/EPL2QUnYo=
`protect end_protected
