--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
PniSpGWplZs6S7c6+sHdzOElBUY5JTVfrevmbtbuS10O3ri/Xk1l8nYkyInpjC4bSltzb1JLDSqu
OMzS1osWd69VyodklPZudloAX5yAw/HbeE3sMqY7oNyHbOxZwDHNST1e0YR982HE2P7TPKVZroSE
sy0QDBtZq6TcuKT0xFFbdCts5em4ENOPxCpVN2xZ9DIgxcHXQZIVGb2ZySASdSsf2jCuW8v7QKEK
M0eIHKsYX/eNFkhI30AuwI9MXDb0gCRA62zNo1kjZWX9pAf+IoQ5DsTcZncnnLm5eqqcEyqna7YP
Om9W1VmrUSHCpx651rYmFPI/jFay5fN0uPmEBQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="2v8yd1bUkGHj23OqQoRzSostlpQjHwMDdVwhmzI9HEg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
NdxHxAqJOt0HgFdhq6hvBWK3ht3ibbNLc/iiwZUCoqK972Ojin63+WgbX6hdJfaI+mL8XfkbhBcd
kD9sd9QF97eXSLA4pNMRA19B8RDUcVpSpsuLS6Vqmnd7jj55HzFnqxPEw24oRQRts4+W+7yPsYoM
CJebhHH3vzp38NJqKwuHA+ywVmrrVutaMBJQgAtO9W5adQ47wW0wds6D2+o0GamwotEGwiuSUbV2
7RU61ssJBpxHrqe8QW5Hc6Wnbn4DkDv0ej1mHgHxbHPc4xTzw2JbzaX8/zQHiXT3ItsVGUDz3yDE
ksS2AU3Av+Tcawv7lBUqOJYyA1L+k5WaqwYRDg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="fQRcIwaydyQ18aYQXtGkyuMNNuwAD7poCleYw8RuD30="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2208)
`protect data_block
lxEx6YkKIQ3P5SlB/a9b5jGiVU9uzyN0i5MgMBaw6SstI8Msr3itNelgifwQDvq+jdELlHV9mzng
5PVTWfkQUBL9miM4YyhblPBuE3q9IA9zUOSo/eO2nVjMCJRgRVWRotwdq68ComqOt4IVC89BCqcT
k+pTfnY6JWYZW+YnbHyN7BZPIV4Bfuk9DwIG0AKRdM0BOHL4GurzCRUG3RUWNIw+QuG4T1E0J/dl
dZzLj7jAmtrGdOUELQ/TqPR+BJhXOh2hsLzuhOkzeGc243Rttd6wvSR962J+mG/IP+czLmyVOt2E
y7dCbQV/ELeZWNbRblQ2dUurmP2IayZWf5uHx2tNuSrTKiUeOmUHnNPq9wgoAFTo5EcBMnuDYVjP
OD/8JrrSqOBMQEi1mO1RIIJWnw4NTh9gFUxVi3DzYIsP7bGTMyP1UoBwHNvbiYDRroN6CV8qIML5
8m2boSzSShbEhjnnZzyUdcJ2GgxRg5D1BbLmfO+DJRF+RQWaR/W0MPOQY02P/gC7dRL80jMCAHXQ
8fqAdjeh/Mt7mqpnnB90O+4Mqv0fNucFLBrhX4BPrqxpx0Dg93QSV/U3AEOPXVPVEiLVReL76af3
Sgh7/9A8t5bGNDlUh1r7/vvX/yMzdGBGeQwRl3hJvtotOgM3hbjEcHmcYgYCdkqaB0ny5cgHIxEc
yuC5AgevMNDvurc/D9LkgjccjuNfAyLAmved0QOXqLmp9BHmh+69kh5Y/9W/27bhuQIp/2HyF2jD
6JPlWjzEjeVu/faTMIy6jp+5mmIQdYaKN5OJsBgBDC2Ign8k5eg+izaMk2c1EMExmq5UvSxqz2G6
FzcLkND4hmbu8GzQm6KsEjc6IETo72zoNXgsng1CUcMuRcHvYmMZPCesAYC9QibbQ5xWpeUKs+nk
s57fXF75SP06lvF2vSoph4ODxmu2b0A1/h2dAskZABtf17iHbbGmyLmUd9eCxPWTiJkSDuXfjcAH
esJow2T7xjbUzM/anGXOOIYsEwEvSJ3sx1Mo0MRyirgARJHDpzDnZpzC71EFMAvRAYdi6h4w2rhY
+SQ/rGTt8IBdvKrDPTPcesQDuI7hpLuTCQWEnevk+kAm2LeS8mgLibE5uRGEDMZ6i8Tt41kkBmh6
zvnRARTQ+kvoSNXautRVKUWo12Q9q6zAL67RhQg9+KU8gfvxwkYukXYnHhjBDq4WOTM93q4JzQh8
1Bc9G/itB2yY1T0DyvpbZt1uQf/ESIHTyvajLbx2S9Q95v57GPB2bvICBtdYawIqGTt45MPrkSn9
NW5Cf/ZR/pZH4b5QuqBrVXZwBDoG18okP8d4AM9hHQpflak7pdjz+MpkM4z20vQmswgik6QcD19l
UF8GgKhtJpHaEkfSsvsrqzyz71q3jrlvnLJGQdaXvzkQXJlbi9shKCkYhLWH8nV65/zOmsJgsoUJ
et8XIcM13q5N6l8/IjhJ17CIu04mIKRJu4uqiq8ky5O37rT0nFDHL5GNT4JR0UKuhQZjddn8Wc43
V7HNhdsPZWeuNjJBkucO7pTe+TcqyWC4hSbKvWClFIIhNktavg2+JAdzUVc7v70WSXUiZhPeG/IL
pOIGf4yyn7Y3b6xH70TmQCy/A1aS69sW1K1nA4aHHsQH4VeLgNSofPxqmeZGpDyrRs2GM7abNA8G
kQ4gNP7aKSjNnJfSfqTk0VX8qv7XXodZ9ZWiVpkC4U5kUJjxEh94lHn3yhorBRv+yE326mcnzYIJ
uaCdbhdW7JRLRN7dGgbF6L1nENa60Vnx/Sf+wJbHze0OuNYN9IcmBu7PMbzLpXXuRdEBPN8NA0SQ
1xCwL/GIA+JzxItjmFKhChSTkCgMyScJ4fVdl600z3CrhQk5cvUD0GpHEW15pc8dgvBhKcJO/AQb
XxFkX+5dRACHBEbCZ6K/LcCVl0Y9qV8wDo0Szl4hiIGr7VYnGJi8rCwP3EMZC367DitSNGI0AKok
LQkxVrzZYMgaPt8p9c7o0sisze4IDO/o1ZYFYAy1I2rHEkUjxRBMwe0VsFufwwhVsf0afijuoxgy
99ESnVvsPNqtf8HjzlhbWLbM/PYCqNtAAz8BNWe9wb0jJ0dDYc0vSAE7gfQRUcHilWkGzWOauAll
p7KlGhxV/gbHVHWoeQpi7SljNeWwv8EwzCJMkx7ym06l9ADVAqvnaihU+FhezQz6bWXoKm3lxihA
t4xyBLu0L+qC7ng4sDV1EpT8wxLfOU8F3GHzcC1Ai1ffbOD7KGIpxOrcEgj+4oBI4SuDDiUehYXr
Du/ZrbbfITTIiF5tJMkMASOyOw1mzUMO2H5J4rKKxh50iD83fOWWprk+3+LmM+DerCBgdawWKyIl
qd7JcYxl9mv8EPnJYnfXbO1vjZceWj1aEKSS7AmQ4ZSIl0KHDE/hbCVTEekyQsHRXCOXTqYq6dkk
UKeWDCv5EOP7Nmq/ZE8GBoCsrPEgEvE3O9Cy9ZLLG7V0XixCRNFgFDW2mGk6Y5fEdd5lAML7xFDZ
5VN1HnzAYoATURNaJ1QwiYTNBr2+mQU0z+THexQ0coVI3AY183kDobx9aGCMYxoo6ozGPes5wbbU
mqKPN1GawvqbhHbM6paiWG1KId8egaz8gNqpp0Mc8ILiMgbqQrivDvNtI3oq4Ir6sOkb+9LhpNob
26g2aiXvQ7AZK+s2F4EUQ8ivb4Rj0pEkXbDvD41JtkhWl/mSrO3kA5KTi6LsRDedLkGsfPUfE2uC
Ef5+85503h62us1b/KEjEepIZ1FoQVLvNf/eiLUCjM1jMqdXUJpkkfwp/FA1ODHsCRuVXKOXTNgS
lnd1Xl7yt9lmKnECPZ2rCs9QUBeFkJ5y+rqyTz04E3fYqDotqE+e4W3+KWYEsNTuERo6LC+K78Cw
Qjur2+G+V0Ve030w1W/1qP4fg2jjfw4H4MKm/bvWAnOZSGsm0spKNmln
`protect end_protected
