--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Wik3ImSkKdHwPnKp7lK6eoKuzpod4or4VLuB/WQcpIVTOU5J8CkpHq3V53CdttsZEOQgdFf3lY9l
1Oszsqf88LVIdjKuE09pmsb7QDvHRGWGbd5leUOfw50i/N/mgwDHQsrlIbh3hWzCM/HF9ytpvWJF
FdQo9w+byWPbYJ4Ji+ZP79ixwD+dzQZRlYX54RmOYKVbphRjpmldePJcWT8AT52oytNfhaEU5zBx
Ab1+Dyt3c3wjaGtUpSXqdi5jlw9sDLhR+cpd9y1F6GLbS1u06UtF+cKN/KRQPPC/tqGFK7VYdXq7
7vP9wJupfYhSt4Cwik67YaCCE3nWzxtgXVga8Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="pVQxArrNbE5XtmeWYcKPUQsLqhvdohf4tVeKJc0ulTM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
ctrbZOq7hL8+CJf+9kvN0BXEdiLXP3fW7FMSJWfWbcOo3iuYWIjTcdy6SecyctYlZRQeve7L2C97
TyAjt3zeTeLvCjgQQGuvfv0qsYKrTat/rzuM6w1eLRrQXe+Fsen8P4akIlKoEyesrElRfrMvmDZh
VwWdERMTahKqUzkay2gD8+z3fUCZhWxDOY/DYAuCxBQFfRChZM7UVCWczW+vbWnBtSvvhQjVfdgT
oE71YAQU6HXMqjI3dKH3/eONJNNTp5dQfuPcAS+kZjZc1BMRyH0yeBZzVpwdVrhkQFB1AD0eHrUo
btSEsPsGKHXFJXZ1MqXlDlL/vOIgyaN40hhRmA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="2zZvLNfLPIt1x/UX68DDwJj82hDDOcoU9gKF/Ej4Uh0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5024)
`protect data_block
WbKMFoGE9on73Ljh7zBSeEZMgQW16U9YoU3rSb37orT+fxHeZ6GiNpojqL503bHzZqNP4wEazu8U
eaAWNMAJr4uOn84YqxucP2nJCe8hR7VHdWXoHDZ+Vc2gpHBQMC+dzM5H569JtcmSvZ3F+Bi0cSjG
y68vb3FqN/OUI68aVNk0TqLF5c1ruKSxTihfwkuOtg6Qhsg1BzhECPfxUqUw0bbLNGOtcqqr5L/+
HPQIkIMrXppFUZtMmgBz34zBQGIjNkCPAuB+WG1fj1p5X0n65SfJ7QSweB4COU4d24/Y88qr7Y7S
Fx6AT+qL0df5OxM/ZpEB6kz1gyhwUQlaqmgNcqj8U+/GTLNhN+agR4B1yiocfIZx7PHAIj+Ijf1t
Do7Q2dhoLiTY/Ik4RWz0WxSwtCxzJsro+46no9b6Htr9cgTcqDAhnlgekBkJCOJJhH//uuPzoDdS
DrKxKbvedTJyGeRbxSMzQZcnkpPLLvPrY1HZcY3SY+DJhiF1ECFGWQYX4w1HsJ+rfXH4xVVyw1Su
LUwkgcBPnLZuHE3lHwHA6OIJw9Ynn3HWFWr43tvIADNT5CjieUvsJ9e0uEdGT3UYSGNzaV8m0dzu
5FWh2Pykt7sEm2PVTjAty8e6fYSqXBV/oiSd+EcJJwLd/YfC/3eMIZgq8hoUxinsqQCxE+yXJluo
Gp5+m4YLHbu6Fbc81ZU5kAPgcfs4BiRldDZOJj+6GhgreWiKYnTnme30oYHRpxzuTiwNo1NqFeDM
E1iajjGTDfUfGind0ApWQcWgeQkcHGRkSrlwCdLa1Pvaw1RCWXfIGA15IksDoZ15tnctuzXAHXOJ
81L2eGXP7o/xgDeYOm1G/ubuyOOXOnqPh12FHJDyMfDnGr9flqp5sSuI/FKY2l5exyBo0lMPmBuv
0Rtn0ByOaQd70nHR/0Hr6AcFvHM/HX+Mpoll1RvkcrA/gqpQ7++3E/HP0/b8kkChVrQQm33f7ewo
R7WvX4d3dwUW4wsmxzJ0n/4sVq28dVB4LnUtKx9bqqqn6cdEzRnWQj2pzCY9SDI9k/DpQr54h30f
UktenDw9dB72Td/W4nYcnv84Ii7KbJ2CekDXw2kprfE8Rs4QwNAJipTCggBfh+/QQcaiLcId5dcz
ktIMDHv8EUBaJSQv/K2LicKYSJBrZOYlhZwSnJQjSnabDXziAgX7aFgEFWqd/so9FRYg9kkcV0B0
9QlRrpKAZ4/qKaru8WwTcReDOLJ78PK+kMZWci3fvxMCXxtAOodDodSQR8blCq1qyIWgdVzXTmVi
91NnLupspaneXr9gid5l5xLeid8WzyVh0efIgrEQVofxlxCuCZZ/W/frm5oJNqp0fN9iNI+ysiX/
LEMn0VQuZB8OF7iD/4So+3SMITXkCiatkGMW7OFmwWimnIkE+hCksDZC7zm8Xm5IIfITiuvGo/sN
7eiLx/HAooC5dqDx32LlewXF780WeghMR2jmjU/kmCTNxzXuCphoFKR3H1gXT/qXrrPmq0YaOFN5
P55s9SEp0IHD/xoFHal7Z9X7/e7fjzusaiCNcxNcNPGlefUKtW3c4+hpc+aUz6D9hvgyl8FV46dM
rP3G32urxx9UOYzesyNxFXJEeIEKdue/QJMN4Pu7MpwAi5687qTtjAdKtVaC87Y85W97EbD2VIEb
NC6bUye22VgeyhIE1NACAI+FefAVXywletkEIUkGZrd6Y7bO7MNJ7EF/Xgu7BqYY2Ta7hUvMmFox
ka2ywo9wISSGIfbilSfmIxAHy6P0GFiTszHIqSVsQKZHgo96lGMqmYrFGnPW8gxypeAM1WsQeUw2
1dG9Ux+F5bZs9auZxfz60tSpoLh28cUWPAhWHqD8usEPrb3AAe0eUUOvQONhnnMXH/IzlYFOn/O9
M8QJ1gD1t+MPUGVpNLRrFTuSCLwrrxIRS4PmBAUrLGxxdWETTAHVBNQ82IRfSoyNbUpF08gCS8Bm
KsIqW/Zb/lxd1PT62FSyOXKwmJ5W3UN7F9WZ3bshMP6fXRv8AHX97wcL5FgSLvxHsNSp0jYEnVdj
/AvpKeIZZF/cxWyzt5u4oJVGrCo7KjZkqSYJ7GD5Sf69KJcbEgq8hL5kiViKeq3yToKH4dIVh4em
yyiDms3nxhpOqiK5golMRDBf9tnmCkDGMJ/hYBTVlq3olsr1IkhvVTjZjj2B13iN5osrv3340trQ
7lIXrnrQg31JpAjZSsrkmJOOrWWZApdZFQ/aeFCUobfGbwATpOocHWF4dXoZCZX6vLZD+rIca74N
Jlg4QEFxd6na6UNVmHeUMuoYkzI83H8Mdl61NFJH8+916toUsIOopneW21sxm7bOwou4VAlBotFb
16ZDKDdbgQXbUljngrrI3D8JuxpbWtQcCvFPIMYu0r0UkoJfLG4SBJl/wghj8BCniljeZSJfBcJb
VS4Dx3NO0piPCQ0Y6VP7GRNkBODxPkszNLiacKc22i/qdHzyRbjgxUBDfsGYHLjF8/7tUVSHRRuo
lOzRur4rL4ilNJZWoLYpTChbMKOq0Qf6+d9GFQjAz3WCErnLjAb+JaHgnsySXlcf1SD0r67B2ML8
JwN3oRBe5lNC5RR4YRPkT6Z+hTantpr9BK+FvcKNnTeMjnaH72dju67Yzq54od01UrP7zHJsxH5/
joEyn+I8lInpdvo3d+B9D/ksZFnf+kTqe3IAJDNr77xEPEB1qfq4nR222pY+H3tkNuinJXx5Ad0Z
enmv22zktoKvpFMzg6+1538LuoZOiUnq4KuzQ5DeUrDCwxBQWLzkFoOtMDdAuJTnFolItYtQIokA
hVKkLtpbG5n6wsZFkRSQOD+hNGxEw7fXH7+7Rr3tBnHCK8i43sQQV8i188UtEro6NSN/8qjS9cYy
OLQLwOblgfBim0B9OIRKIH6VEog10u+9+DjhOGs18sLEm2VpO0OohNsiHjT2XxuIU1VcGGqgMLUF
PLunLR1r9EYZaViBlVkoC/ZDZm3OlG6ocxyN9xYcPt/QPNqG6i8mqomz+ca1F+SF2Fu8GB15YwjT
WeNuFuWTnCht9Afo9inmIujiWSlupx2+FBAw29nbeNk9K3WdJg8VbrBhxK+9k944wArIZ2dowfau
mYckSTGSFb/V70LYXX0FW+Z9foeevVyAoDo+ZnqOPGsYPIQML3cgmIshtwhJIi1s8B3yOBvMG7ce
cnN8WErneHr909JEGvPENUjt4zfk8tWkb8f6hf8l33NvTKULkRgoT50HTlXCf485vovF4cxd12El
aZj63nsUrfTS24W0o2SWL2ZecCtnLoNa7RwvjhWBKNRaH3Qx0tvm0n7wb4IJYZwkxF8kqpt2tD28
QIGpB4Q+HzxCH7e0uQsPXgMNbFZz0kPxbdpU6L35rZ2jh41+bYUiGJW/YvuHBdvqoeYjb4n/+Lz4
PyJQvtJuYMRA3tLZ1kbV+yezCkg2KhqCzZQXMXehy1Hrp0YYQ19Fnpn3o6Szp9fRPnJv4v53Tnnr
o4NSI5G6ZK/YiZGI4CWrX+pSwExQlm7X99PXR7nrUtABdUwZHCpjLpJDlm+nJ6UQdg7Xxa42bCAs
O7HAa0zy5T8Hen9bqoa6UAQkkaQjOorrg71un+1jYKlMk+qx7bzhjkJb1sfys7MfjXm2nVucsyYL
zdMgVSO3q+DRRf4fvaTUjVxhyGVJPqjTpPOUq2NeQDO6uNSYPLkdITRevkPSE//65juxNhdSF7M8
lh5oqwm8t9rvgSXB3PyMMWz8NEHkXd1YQM2n+jrHHGXQ76mzthG99qJCVdSaJ8X8mvtnDjkulY3M
oSCfWJYJM7K3mhEiR7h1JWuBYCqDA7HCk0BMQ4wlD7cGMIHriFP+NaNyqTTma3Z2YlrUhrzOx0wM
wB3weL9HquaQBZtSJoysLlzInTXSXSIKWI3IUWDWcJnjH20/LapBqur5zoqW3BMRe+8ka0QBUheB
Yn1d3iQOEr/oTPX32AdoPFj6pwRERnHzFZVCh+7UezB38xZyc2uRin+Mv+Is73gQGknGyCJJeZ7j
+HPkc6GvFKA65mwk7tLzLwNeM2Du9+0pPuRt8FfDhjZOxrcYg3AOFGmh2dl0+qiTz/lrLM7KGZNU
N5sxKD0T9iNs3KasXOqEAnyLnbH9TgEeuku2zm4yk5GzXp00HyiaixFdnfhfV7vt/axcQZ4J4STi
phjS3R8BrzdyUTJ8P9eWggcwxLtVWIzNl20pORPJRynMunzAKCV4qaOY3Ms3mFrS1UyCaxrxqq2Z
EpxOfCn0rESw8v1MwaDOilPdZEtFw9sx3j6hqtjukwOytir2Exwm/i75CIYcDfmzQBgUK4ODXBzc
e7kAog8s1IeRYM8UXKC3CyXresrFLlFC4h/mzsHUypdfjufRkeT5aDrWOqc+934lchCuDfvAN/NP
ELNUoBc6iUR0Q9sGPwqby1EL74yZ94HyZ8O+DtLrEFNJAnXXdw4SwXxS+GqhNqc+5VvSr1wNAxsm
9FNMIG3VkWphlzDG6kNvX8EA8YjuUvLKHv4cRK9FL6MrkaBZJtF/aszbnQ/TJBpBRxNbj7sxTrkX
HTwWvY9ocjAOXdFZggcVDYcCabNrWUNjWNdtEQRRH+sZrmGNcdx82j7g6n8X4op6GB4+QU14zIkW
n4wNmPHvtBoriXLJxRiwTnI2NrlSBO+3Ik1qJwLy1rUAEPiEmqbXnuX9rKeM6kvUgf8vNu4WnlLX
YiruXRgVKWENAsHCUqPjsVu8wWwSXRFNeD9lkU3PpgQySzjL+LdY7sz2Am5CRsHduu8BZF3oOYx3
SfO1j8UrYJzxsYKcC28CwMLzEQ1hw1sv0etb4XrvlvqInHyx1Dd/kmOfrKKBtvjuXkcItYHX3Qid
FZK7gM2Tl1EvkEhkXicp7JZ+xmupLaW8Y1fhzkum7zxVahH0bfMiUC0GGsAAt6+Pc9T3w05FjAq9
fmaUG483rdfjz79UuxuG5mn7/9X18gDUIo8hxD88pxXtnPzvNDWst7VSc3oqrIn7e7nOvcPIniBI
UCQTnjVkrJWeElqPb8l6jaHMaJTaUjW34G6Kp5ZPTTnQaypG7iFLaa5B2wWsaxUJNnGHU4aXjSfq
ImxNov+fnS4w8j0Vkih8BHpQ9y1PowgLN387jUjNPEy0LF42yoJL0mIcem14+5Zz75pRuTwGmkwb
ivrAE8LxebaNTrGZG++lzBzJ+2PkUgkRJDFwEKv+24nVn42T2axtt6UNjuyxx/vD7v3oT07DAX/6
GDD8SlBRH0JSRakVn7QCb1FGLuWl/WxgngM2c2rBS8ju8MPVoavVeAa5llZvCJHcu53lstdwpM2R
Pb7XHd0HjlFsCCjNqS0xY20fnrS+YEnHdkrsb5zy5LE4mI1KR4k9mAmfYmdihhbyHMeW09qgmQTm
J+pbWn1Jc/ghfP+3tRwKOPyWP26G1QnlegHyNRb7HDOYbFoDe425XhmrQXhs3MTzFtk3vv6IhkB5
lLOSio9SDp26zHPyY2abONvAVW4W6T9Vdbg57VlKZvE8i1Z/5kopbBRLKTA3Qgb9fQm0XbAfOeJG
pOnOvi4+SxHGTYyPI6SXCgXduMhqRj++YhZz3BdlCBVOHsGXpqn0bhGbxg1mK/iEXrEL+zIra0hR
N1YYUPDMSsH3IP8vQBK9zDDUTIJXN5MV9oIQ1oUwqPzjv0MQN9wiN/Hk1eyqFCu5caO+pfqv02vE
WPHVrOhxeN0RKHAkDW3fi62R0R6flrLQXLXilcFs6v4HkS/UL3JXOONiKhdpJY4VrTMaf2xb0nMF
9HJhtO7ri9WUmdHizJ4L9tevNUNwohDfDvI8JIrRPlb/e3952PAjuvXMSzH7aQ4hB2g8iAH9JbB1
03iNCUhsMYqKecnrLjt4k9MIWGFl8JYqFN1/31mTkCbFQ5kGf6fpBL1zibmv429c5YWMc5c9HyhQ
SJjis3vIHHQC21w4i2oFfYDZ65QVWBmH04lKh6OJKBKYlySNAQ+tJZX1Qqr2KeiiVJpfcBG+yJVQ
pgUT31xzZlbukIS10BJ7N5PthiY3tRlO+skm9seVCqB0yQ4hE5EKSjJEZaEQSvIGRE18zrvjKSrh
rdiGzVpFPqTQ3nEKWbk/Bn8nS+j/L4RCGDj+DxaZS21XQuTgDYp95E1hi6kmSWegGPk7z+jvtprQ
4NDz2OmSeEhQL/NtE3tzqcuLmTK51xhZiD8plA9nbYHODVRT1fLzxAO2RkCS7NyKouuwP2W+z+p2
NQ65NypKclk6SAwoOIBfIMIaQeuUD/ikkT7cDj3N44gwrTzGoYe3IYwPUm1WrYv8g7kw3UJ9Ket6
z2yS9854nb6XbyoHFSodKLUWhfYmMJb6ndmjNEwpHS2r752CwkQBpcNw1F4AouE5zpvkUgY/GAno
ulSocAnSq9e260Zets7aMN8km6eqgvpNvUWzPBpwgl8QGWrbhypOPyXFl3sDJjDn3yGms2xTTmPa
SxxKb7z1fmk9qKIBlKcwOT6nLWZeYhPoffKVta3cTJ5m22LR12Kya+K5xq9i9NB9NBAHCRkbnf58
+ot1+Zut0HBnPuPg5jPoHSRW71YV5BxGEmqEe/GdlYg+QssgMRUFzkN2BGu8o3Q6HjPdVV5taAEv
P8ey8D9wJIwRJ3MeRUEMbDedn+G1fXYX2vl7LalC3ins98EO5gMDKws17bhM/1qHhewYTWYBPv3f
sOW0YQ7WNHs=
`protect end_protected
