--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
lyE4Y1VraMepldXvOboDUBW0bqIZfmccpCcyys0UxnTGPSfv922pXBxo+P1W+pthnLH9e+CAt3o/
nY+TKz2SeLZEgaSizPbRjg6f02mCXE475+k1eJKoR5hpHSnbg+Jbh84BrvPcWeE+ZsBONae4fvzT
z1I5e/vjAwEPBxuuEM+DAOT6sB0DGiTXBZvySfCxU2cMLX4VAAsvk/1bWwDx3zOhGhTSH8Q4cNyQ
ul6xVM79LH3wXHgG5rSKinfN6v3CNxJ8DtyDcZkfeGdY1OxsLwhzxXUT8QY1Bss0tlRHNVRbjCib
VtrPL46ckuklzeIxiMmWEYCZohUAul12+B3i8Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="O0J65yEDybuib2iHXoWwwy5ARXixfx+Hd5S35tfAoLk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
HouCtMh8FZbUpB19Pa5qFeQ7VaEbW8jPe3Y7tvDD/m8vSu922r/IrW9pytK648PGCVyzA+gkt8hv
BJon4fPTwCqdDMovq+MBBXODrn/520AXH9iZ7a8nQPEc7SrDpIG38mZXkB9bDo35EQgN4pBgyhXC
Gkbc5He+WYf4EunP2pF1fii9yorYv5vO2fLjK2lX7dBAc4ZHyC4Dxt/WnVaCL9EO0+/xjOp4NAe0
Q5Ee7ZdBG8rLrAg9FnBGqjeAiwEgqP5rTIi6FVKefdt6EdEFJLL/9bhWWoi3GYNKFV8uPozmlbja
WITvk/tdpJuxghhpWzPzlZIofGR5gbIyCXrxPw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="+/PbmhbSluKCEeOlyFPT/lvB4kcNoJSN7+Ga8P5VsKI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3824)
`protect data_block
+ZOZk1QE06O8C9lZ3R1imZNfqbzwPb4BsjqtDRk06Rs/DwvlJSepZhB9bRFcOFsCfzDsostj5aWp
8fRhGRmrTo9rybqaMSs4pC23SbiJq8gWLAzuUoCzwhq2TER5S1AxqBiij5GepvHhtWQGwgG1Z/wT
9ZhwqfOt/ViJ1b5gtjR0kqs+QIkP8t8rAMILi9ltLi/Y35u9I/dlzFPxVAfLfh7hteSH0G84diPx
WllG1bGFshItRXp9+Jog29Bu+S4M2DJ/kH556pmO+vlE8HbV/69cEmoX4f5zySWywP22g52qKLP1
KrbUuabvDmvvipEC95lfJbFmS+cWzN8wC7/4iI/C1qOBknakVB1dMSiv0o5mtrN5Lr5XyyXTFEUg
lix9Ce+3YNK2RSXr+cQ+bc+ySk5sk7PC3vvVPQJAkhsU+L+oQaRvbidYnlDEiJDN7mjZtInWRAxG
Ne/XXxEaDL1CkmeXW86Kf3PGBEUrWdmv0+vL0FBxI7/HJyYzMzpCYFSKzuF2ppOboHui2VI7FYYO
lcoo0mwSQwOsFj+hWbhP3tIBmQQfRK1diCZvHx3mQfGu00ubOy9jYD6Xtm6KJGy31GFnCr6izc78
sTdbNEPCPJiScGmQp4xNtw8u8wrg+6BdZc/Zvqf/GKeJFq2dZTEZVKUrbjs8Gy9Y7lfR9ShtR8yw
AC9fjoQfFiC/ZfF5VN3NwniyPCVYVLsaEgigo/ruPcfOZuH5y1uHWuk7QtCcp4PF2wEISi2JVuO1
OJ35UrtmdzEg2mEplmOkUEGiCHvXkhIOpICOEZqOTCydRcY8p4Tf2EyAJNfc5B69qUFkqwaYm0be
L8WhOeblb2fpOxvmYflAymEWp7mpzGyGsP1O+8i86uWqLUDVNLmwPhbxZATdTUBndN2oIYWXjze0
ErbiEuDnibgGlvTDT7Yl8kqme92bwQ7Z6HJzMZiR6JUXDNtHmhKZFSGNarFsz50duYs4cX9EdJXn
NJUDqhuwhCd/99u2tXMwxCKYR0tAqdDYTzJxOL1pUbVPfFQP9uRkkpOfeS669sEPL+GMQuK+6u8P
IJ78l/K6qXIgIDm/dC7tzuHOJSB5GYJO3mC70WHsgz3iKFW6dIsXxVQ0GkjG3wUDw0rYuE8ka9Ij
h8WF5p9voA1cQna42qOn0MVm2T7WmcUKZHQvEIqGaUAZh5/a/cU4kObb1pIZBVn4meXGiwgjm1F9
5qesia5fbgCVqc9t8uourgPIdyUQr5Kjzzd4Zi211ESA+jZQkM7uHkil0BhmWQyfgM4Z79X9cTfh
NPkGW2qCKWEuZ6nWDqocBPOwgYyWaBw+v325fp9kate5YxGnZM//JMb3AZT2oBkCyzQvI1YPdHcl
9LHPZiuPOO3H6QAG2uX13iepxRE2DOkmzojeEFAiyXPmob4QAjhTdn4JnV2uD3zBfSPeC9F+fWWw
p7sxj1uK78fuCdVw2DnOGWQU1rbRwJlIYXnNrFu53YZCVg7WtsAbdt7PLJ6urWDPhfimA1lxlYOx
BJ3uSLcDTnGK6SvPbFKc+xD74AnbkEMGyzKu6Zm94CWjofy2tDGGU1Cvl0cnJVdeH+pe4ojGn8+R
NyCuOZh6igGtR9/cLKNMrd/0bYruF5gnXq0hz2ShUUzgpnZ2n6x3lnNJP857uU91Bq6UQlzb0M7P
4YJ7uvdICXsd6Hrdks4HZjTzvOCEw8AuTTGoODNVJNr9am3rlSKkmtNPPHb1kug2qK9MYosnphYL
iGjiCzACD1Szn0b5eozPnImlWj6rvJDqs3UIrPSpg/aD860jNjFopnlD2U3X4FDLPkgag4NpfM/W
tjvnQi0ZI4uIvR+BhMzBbNqMFmlkeibnPsGT/JsNxydcsNnRDW7D73rr/yJ2H/++J37Z8t0Z1sws
Btfvr5d3cuCYvCswRb9wHVyUOTcbHtpksODXRTyqgY+hdQxFCgcB44IHhpkW04FzLzZNIF4SZ0gP
9N3jtJ9oNLj2AaTDoWnpO2+KVXqP0UPPeFErQlqtw4huq71VGH7PlGwf4zNLqIxxPyjbOE+qKLM8
8z21B6+tuzwvdOiPCJOzzmgJTECaOHYVvlBDEkD9eP26U1mo4rJTcWJE43jzFRNax/xhGeWuK5h4
Psr/eZPzfQKgzWySFGZHTAVFL9egFI8NNAcsUGT/xuc+A3K7G9FcWvi/tGczIcEORjk11pGZNQWj
Bxi1zVrW2QTR90w7XoyzC06s1ePLBEqlGDLRPrTFflXlkmOrorAdNM4KBqVrQCjPcb1SRZFIha2N
em8UVI8ms4DSZ5OGfRIxNo60cmCnyB43fBa4d1jUOynjSEoy48xtHRSuoaPp2K2w2ZePg+Bp6exF
VoWHfeEU/6nTQTTsMg4mb7ZFXta0hSNYr7EX+/o3hlcFcM4BInAxszGxW9XYMS8KPo2ES1hx4cvT
A7TZwVIao7OrnTwVujzvhP/TFq/mTI3m+o5cHs1sGczXRpArWTO9WtewnIVCZW7wQzMK3jppEZPE
q+RVAKE++I0STMF/rUM5yJ9akZKvsFvMvxejbPnUdjEigTw3YMlgABWzinrzmPlzzFZTGHqhgkA/
esCZDDRvS6ynDagx8SQ/e0+sYsjUvEVcXOE3gYhV0wTt1BJC1aXfKj3Z5XzmWEdaxfgL0719nP8O
HZLbQfI/fbR5vSIPRanOb6VZjSDn7XUvG/iZCFoGD0Ic0RPCXkfSHhQIYpZ+fSM8AZTLkEy6ATpK
i7Rcb3d5nDZwy2/FFWcBfcZkI7O5FRDES6ZXnV4p5IHAKmGQkS7v0EgxfsklwGVfeF8Io9yr3CCX
GGHMEWDmWfRQlP5+NUT0a883vsFpEdEPPvOq1w4GajLqwYgEDqP27C2zJccvTNiYCnPsha9RPuFv
pf45hYmfAoHVP1TmFfkh2N5OIRF6ugxktWKZuG5rRVc8RoKkKREHLvtQt2UyXNGNBD12821rv8gf
nLxv6sAmr8bDR1ENsbS+wKA2EbXuRkfCXZ+Olu1fPvMOFD6QUlJNZXUDG3Dp5GN3SMVY/VNq4Iil
3HfimJz02N+L7IICWi60NS7FUftrac2/FEpzm1exrndAr9reXnFWAeeD+ubuMXyccToAMLXpgFMv
q9Iioa63TtQ4DqmB/BIMOGxo0FN2A0N2niKB6G0RvGRlMu7uqgehU57FxRTol8lAjiVk3jdafSqL
fNvdGaFz9Lh7tapihtP6ESl+7yyn9TTxtaLOqTv72LpnY+5oDb5VkoQwYIDbP7qIMD4zN94S2pZf
Ja03HUHBRIZK1ZeTpn9UlLn7MIWnIT88StB41GCQ/1CDX7w6oqxsBoQdfLeYsM5hSQk/wvgUp55y
p6ySy7/pej2op4OicM+tEIa9lmCD1NYUmMDc4b1rAatIiutIh6IrDnaWK91dUA2UzHCELzIWrKKr
l7AUCmG1ZEf6EqtA6Qkww8vDJ1QBT/90gUZlqVdQAs282RjpV0vF4gzb4qyrjYIbL0gBT0WKX62J
MWDfgQnYwyL8RarcQ5aLz1PjHjZc7zp+1bWi2ZWFBIjPm0KhBX1vjBzw2C9vp7QuETJN4WTyJ7bV
YBLBxm0ZsGutR+i2PFWpj0GBFCaaSN6Bngx4fGbeZu0XrPs4wTN2lAY8awnj8JsH3xO2Mz4SjIdE
S4xrE5x95KUCbftqT0u+XxVAoTIWDiWrOVMV0oiK6Gou/0Qrc6qg8VVf6BlFRgAP+EPvwXChgKMx
AzvcuCGI7bRPGNoGJSzU0tuHwE9PKaN1SVovSQAbZLUj0ycrF4vefTy+7E2l+HfaprGLpKpxpS1S
uT4Mnz49o0PKwVIvwBaTIJVEj8NRFj2bEpnNPeFJGW3hx/6k123gW6NiAcWEFRuOu+FC9lAK1C5S
G4++UiN2yS5BAezPQzKmobBCYbvn9BF7p3FO8Zhu++Tn2ckjcKLxRlpYwryD34puMyUgwpV7peI+
DsKtr+Y+Vu0Hk89YHTnZEawMBrff6+q115/ZpM4qgyk6Z61yCrILiM/lJmdm3IMYOgEzETn/nNv/
NQmEJhihpoAvdcUPrj9mJX4bFLy9aYj6dDXWbVnfmTkv6ZsWyx5/846Sw2jbf8IiG9AlpWdnXSvg
/dwZVsOHMn85fmjd1Vrom0O8R7ICPGheCC9wYb9vT+YyRhsS0/UijEKOnqHlKtauS7IfrFE7gKFG
hSsR6GWKbKcejDEEGcdfRME9psLW4NjzcIy41EZVCGDV/OCt9B9pb4lHDo9keqT482jOE/TAdQUh
l/nJUiETLbr6sGn3KxX6XhwHT/gdWuVhIfk0ACqJlQp7Z0/2SMwHWw6GK1Re5eov4KgpmmFEKKyN
a6cXekYaDkxzpybzTQkD8xfik/chbby7R39mKtL3HqO7ZfUxRjJ0rOzZndKA7ihCo44jwyBzMkSp
k1ocvAwr05Gb/AG9qS+GX306RvWefHw0dI1Z3NVfUNetoNKPnHhpRjeucj5xTEW0ogorntxAyT1J
JQP+5jDHe2Z6ANCqcGJZD5RtYu3m3ubYTtMWkB0HGfsN4uADBG7YVHDZ6m9UECxk9Xm0YPn+ae2V
rnigGYdpeZDwoTzSnCL8I1KodSXUO/5Boa1u8QMWzE3UdtZXaZxATFLQtozhKv9BqOxdRz1CdCLF
wSKkVvjqWvdS7JLfu9KGes/5yDk0E3SenLtQWlpxC8nzO03MnV3YxV378xed5swwHVpdwQ/236jb
pIUCgDivS+nKeRZBRb3ySlnVhwJFj01lmoJJWP3iUlqie/3YLVbxoXIUGeVq0zJn/j3O3APe1kDU
3gm/dpZmuZuBsFTYOGxEjHeLBd8ZBajpnDuqjeOBENZXUPiZwqhlC4m/7BxeGNzKLuTblz+gmRHv
KFdknjrvpBnYWFsuh9Z6ZrXjPdchnqLn5dHSMM/HAIF126AxYKyIxjV5thmNxwfgpmi6ZPQiI9iM
I2EXCtlQu6C6v0yKN1LiBsyrK6uJDRTGJh/ySKdbV2L/aFSebn8BJsaFkmnV2U4xzQ3TAWmVc00C
1rSvDdvytiDs/nHCfxcsR/1Y5fKL5vv0G+lqnAdRxl/0DSC7v96y8F/aigdyAo+fFlp/0WNInOrH
kEe4Ivk=
`protect end_protected
