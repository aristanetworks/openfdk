--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
EjFkgrkBoQXGFK6TZvN7JfgbdXk3+K8J47VGItpWEkZ6ICvC65Kqw50AVt6NdCjk377GL1jjZ2u7
QrJsKyLZpDrF3tEqqlUKvlFbh95VCJmb98Q/gXOyuGF7dUouAFLwYAK4Gp9ZRA0BU+MBUFow43YR
6EhUV1S6ckGZ3y+98XB7JQm1uGEizq9ABam0Ay4lRwDqMvGisawuZA9xT5gOi2OFedChTWNeJYM0
6JDU3tEcUdFrUAXOHrvANfkLVcxv71gKB50hkI64QhxQXVdb07gJiV3oyJpuknlX73g4pi9ahb0Y
dCYYJRrsWTL7fxkG8OzVU56Y39cYYXHaeHEClQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="r25xFbEcpKTypgktotz7TCAQP8KFsQVFZoMBNacA6RM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
SC42JqXPiZs1fHDbMV/45Xi8/+PtGyu5V/SpOZdWQsvdcQ9cSc0GkPLy2BJpJyAIzeQotJZXx+OL
/QienXNbCh9dnv8nXogvRcypmYAC5t0aZe/YRLpgUl6ChFoUO0US0DCpHRuybu7y1qzd2+CeJUt2
Ypn808wFULsY5F/XcsMYq4JITnYJMzi/iG1bERBAUFo7ThCpN9f3p2SmNDrIq9Zn3CGZxmqwuGWh
BHnAWpEcfR3K/N+0PeUOR6L14+ceDYt24kPT/fkYi1GC8xoR0wQRZkWDm27uXAiuR+sh9XaFvp8F
DbHXhzH8hq0I8JIrUQuGbYOIVef1PZb4n+69fQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="OB+Lx+AJ2B7VuRbw7QHPHOYF+sQ4GPH9fX9rqtnKmGg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`protect data_block
AxaOdaALiKSjMAKoheBBuAVNzzqhWKYavOnc5TfSZEX01SlWtRLFBVvUQsjZ/B3Wgaa26iM+SQ5F
2Uj+rs7n9jJFqNO06u8JQxhxCE/nDuSrLQiHOb8D8VBaPGBqSIz5oDYVRnXo77ZqOE+g06GTVnsR
IrHd4XMw5q7DmG7IEtCaDMrtv823sCR87oopuTMv0ey9uqI+hgQfYJ6vQ9x2uLafg1+4US+xdQ7R
jLGw6njUEueDtZRPTvsJjBw8X9iCkFbAQPu6cIua90dJUJdbcNz7RSwDXuo5mFa/5DU44NZCSuGZ
DG4J9DSaOfW20dXQP+Z2Qo7MulGYRIFYtkIsdCJBwRoJDY0bVtj6HgcYtdwh2XZ/xE+k24sCQ/jA
qSQenJlBtBHAbMFJF5VP/huhmeBepcZQGeuXmH/QHfNSf5WuA3G+JuvtbZWdEfi0AJlyGIwJildh
/mAIY6Mss5f8l341e+z9/i9BAM/iuQF09GL0h7T6filx015tg0xsP2rx6IYhZ5n7KeZvna8Crpw7
klCGAbBVVrEAIzg6zXKp9fZC554MzFonCYZGHP7RKoFfSmIwql3BTI1f3YHuzqjpgVHnVxTKwjMZ
0DmgJj72Wp/ZW85Lb4Og+SjrOXsOwI9u2Se6Nhay5kLtdcpFPROen2cqRmE0O3gDTPzZVelgSmzM
Wwbg6Plp/rxKCFMUw4bdJzP6ylVlYZ3h69v05NHse6U0SAFJ8mDx/L7WpSbSatlG8aqelMy8BXWl
k7dgXg3PHZqUWuuZ3higSjkhsYAeLmssrFJYxu8O0tj1aRP8Zlhyf+CS4F3m1fESOFcFUM+gaK2Z
3ywpw/SF7N9db/b5iOB2+I6szkXTZ7QGSRyA+D3jznqe2aQW+is0g5NuOql1K2nv2RGEBDLYlpuk
tT2EYTUfoG1YjieLJTYW2rSlSqP3rOoooaULTKKTEPq2d7o4ZMoToXBUi/WMC08ldAA6ZYE/KFwV
m+1iEbqsunY8F9HL1OF5jpCc1Cftj506gcOmWsdLYadXRSQ8C1QBCOv1bJwyJThJb58K7tlgmzCt
k+DgbiWctk20tRx7My/bMvmHh6g/vA+n4tITG5VHZx0ObcjwnEEaNSZFOExeVQdkSv3Jpx3s7ntz
qUQYa0ewWS0WxaHNTrLXBmC6moY/7OxMOOLYROBt1rko4h0kUQg2Ud9u8iFBQVw5QYKUxYBctPLM
7H5DbFEPYUo3VNDLxo6TaruQLqPC1yBU2qSwl/yHJCrD6NuAVoSCtNMYBgIxMX1K2mJAXaL0OTAz
bK5GvMH4pCJ64+WJp22cPtu/1mH23xU7sYHJT3Dp5XZJnI0Oji+lPAqtiPmMeBlWLsChvY+r2+Pk
mkFWODBsoiPnRlqr1kokg8D+vboMhtXHcoXXayLpSdG3EVRLuJdWKoKVQafoyJwMIKCn2h59j8im
22qHrNMgYAwLZTUMR+6b94SVlMWAw9XYJZySiULcrGivwJNoHo8gu2Oon3I66jtIouA+Mion0WNG
ntIpA5w5RvyhuEPCLm7o8mUxOrJB/78Xyvu+LgLNFUShjdChRf9kLKCblHDivnegP9B23K9C3je0
gpKvnMhZkAbr17p4kH4Lybvw7QQl0mLT5wUdK8IiMYI4jblcjrHJ03Chr7XNjtJ2k8o5dW/YCtHy
YNf4vmR9u6LwyDYfQ5pHMqRBF48Lu71VSpZ0L0zMp3ImjO2ZAwhlJKZsmdghzEM9ud9K0Uu5iZoQ
XN7LCpCs8ezG+tWCfP+l5RSGW98b/7mx77GvSjVGoyS3IPFw/EFEarg6FhdkKuok+/zLjS0EI+46
2Mu3J+Vg9GSXyGQne+0USXpkDs7E9FP1x61xG/JbPg9zcUtqxWkUyu7uBkb+ksntioiAYz9nB+p3
V+POlrJ3VAgvw0LeiGZKXHqBYs747CLm5sKp2zxO2ge6RhOQq/6nhhIBdc78Zy00pL0vD14cVq4i
B60Gf1JNv1PLK9ekH3toZe3arkeNFYkhcyWVisVX38XdZwV15nHbZMKg4LcC8HPYo8Sld6Km2DnE
fsNcQDHOggAr/dwjnAqqhZvW9UkaLRYfi5DzqR9jSpQxteZHGWikzdIxSgFktHjFzUOoc/OEPlCu
zrDyIcPSuhkPb7YpHNnTN+cS8sjgGoJzGm/ppUPyNr4STddGSmDpzoNRRr8uLw61YxnC49+qeBzp
SdGJ2EuA89J2B2uvBbuxIgsdSRLuNHHy38ZLK3IQyc16gfW8LNgqIfyRQcNDxSH/aWtIaKkg0v4C
sL+JwaT3r5wLT0eZb8ts5WyaXKPKOnS01nTM+/igQyy70dp3Ygw5d4Qw0x677z8clhWyRbU7bqWO
AyQLw40H7APYcum+n+Avi2wRXIx3+VWa9yXz4U13JsTriotzA6Z7cNfsJ7YCGFkma/oUvEBBd7+q
kpSJM4GeA+P6f9Kuuufy8YTwAle6X6ZnNQo28n8O8CZyCxv/Sdlr4FO5uPFAtSt+Ms5Z5CbEzkc3
RcNSTMwzWi6sZXbSdIGOwCO9tFhIn0lQYYVtj+yey5bki00cxDD2SUaFaoU6GH4/I/UTuCj76BUm
izdcG7jwBiFbWFBRbJZNnd0OE7KG2lcHD5s8qOJRTn8D/73WH3XyNePB/4EqRVhU1k0A8zeDPMuN
/aM9t50YqCexJQdIINql/rT/OWAMtRpZYY42lNfGJl7u/vcNu5CaarTEhdQHPkHMLgUdMrRRrZEb
4aK0EctubmaS1B7bU5rQg1O85fiwVM2LmS601HAP4XXm9sSam5Qyx+AkmncFaNMELi83yU2HHlBE
8P49SJNGYeUXRuqUPQ/s99/AZyQXZc+S91LLWTRytQZPBElUfiAXgTEoGSspny0lU9DlqPGb9SoY
Svs1BhZpVqgWfLLSNegBv15q9rLRPwVBS8c5BSgnDU60IZXHzuZ70Mf5lPPHD2SqkEHBJs/HGua2
OqM6xEMKNjTlyU8ya33ljPufL+1xGgZNROBed7O9ForGfjDbWvT5MCLd6xczn+5d8cI71guW1KO3
tSWRCX7N2SxsQ984rBNkYCXMaxvrw8kXzHRLoWVLPpXgWo1p5rc4yBr1mCLOpJ/v+1U+ZlTCKN6g
gIPFqu3VT3J/xYd4j8mMmNR2y8vYz1DfjPD1ta7Mi/GKf+qwVGm99+w3eNHgk53d8a8xJDWIvFej
mWadioJeHY01ZGqrL4gRSwOGnvL8acp9BBGtNyq9ku5L9K9wMknd21g/e6cfK/nulvalTbKLJFaV
DmbGUqSkmG0Uy6vdBN/lnwN0KDdMpR56dnCRBvNB87j2nQn27hewYWZ4HuKBApC8cQOoUAQUKmmo
FHLaFW+aT2Mrr1jwCZJoZHu2YNx5VIQs1HVcySwXDjz09kLmp5PaCoPI4Di7GUI+NvCiXhL2ZI+t
RcCrDGrIBgSlV/cDldyftvGGiY5In+kwRhxc4Dx36tPdrRa56cpHj4ltCPuQQ4qMIInv3sfzDSCh
4LreKQ7hl5H4CgTeHW+NRySN/C1V6pOOO0NwTtxI9W6YEzKghamvm8x5uvFYc4QX6qjHDF3fcgRg
hbJhB1O7+V3P5QzFVgIt5ETGC+GKcpeknLY2oAiFl+9RW8jjZ+g2HfkIkDPoIxnwEJYxwx+vcbs9
cxxfRjZ/YQLM57UKttDDnymtCgN6VePKNBO/kqW2+ue0uSqv1Tjgn7TN6UCaHZnV5CVlB5cHyNVz
OdFJ+VeoA0Fn1v9JpoabkzCwecZgwFEwIYt4mm03pldZBtikkpZEo/oMlBpVlVdjS/aaix22ZRv2
zYS5Jwx9rHguo8UWWVOClaiD9ks6JfVqFy0K5boJW6kojT+61L5y1Rjp7vKrR6qtQNbKpKe0ICsd
TGklCB15MO3p+mECQ9K91iDkpf1dIP4GqIvgXnkdHkzmT6o9Jqdb/g4uUMcFpK04KfeZ78B5EIJA
W3vKO/SRti3IAB996yCs0/HxuUMI989OElnEq7bTQIrL9Ap65pR0uj8EXoYyEI1GApsH4YKx5GPV
Qat8uRMI2EX3AWJksr7aNP7F1lNA4nk0W3ChFexwb/qwmEUobs/fjCD7o8R9aZHLiuPgurSl+gYs
x0t10xUfwDuQbN+BVpVLy/KHt/9HbJ3I3fk0gLKqG/PCQe2rGk4tCm7Idt9MCi/vn9QgLKLZU0Te
x1TB0cPiIHD0wWdHfapHyJt4/0OU79najAvTu7KV8JMZ
`protect end_protected
