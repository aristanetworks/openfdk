--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
LiAPjJRz607vXJZsgR1GrEBfR/hepFRlbbRwiqIlz/EgrW+Q2o5+0EJ6Hb1Ke/WyCchjxu+q3Ia9
2E1AA9Kf880EEqgCtBBazOux5b9ojK3wTXXWYZcCWUaAXXch7ZXlZlOcTr/OPfK+H7VmQKHbAxrU
1kna/bfvT2D6UgTwEblwrCE7wT73gpdnguxCXtWKV28Wo7PAXqQHhRs+9gFkSAXPWcYVJ7scDobw
F476PtT/iWiyjLPihhfqdmMmPcX9azjx/ETGydf0cs14vkBYPZiKN5aztRlVTGGLt20kgH0leVnp
uIpLAyIjXD9CuPK98Le5lRWJGYRtQ1JkVmC+Gg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="e8cSPPJbYumeibvaiZxdduaZ2OvOvMsBsQ6N+AZ1o6w="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
WDACHheyo7MfAyuVIN5bO/sy8I3dEoTXmekDjdxluKs1WzjH6prv1qKV/QMpVRcxjFZsjYmGsY2z
CidpCNXPkM8eXDXntb9P0SUAqAnA4xo3svY33tlaOTGZKibp32KbXHBBei9lTLvQ7b3eYSiW7Xj5
5VdPUHRNyUcB9UWNb6DCsz74cLv0OSRhTEufoyiJQ1MpF9MwhhyMZqhd1eCDpL4qkeSUZC/LjEq2
nWeRT59SnGKoMSbVw3fpHE1We4DXPSm77DKiXsATtyR8UWv0EGJTosGz4C4M8sXZxAMBlcKlegQY
lOFDHI9We1LwWmTzwIJTks65FmO/jVDNaGJs7w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="R/ZGn3bIzkqdHgjSwW1EYlSHr4gl1yLThXWAQjhBSCg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4208)
`protect data_block
IhpwQk0ougUbzyJ/eeFHVWbzR98LssXzzESZLoMW8YIA/cdGiyprIQA7v0cjNYX+JZh2WFnL6g3m
5zm2W4FcvyuzrLXdPiMMkMci4QnQkNwfbQS/ywdRq4Cs/mfHIqds7eO3Mfjx11BslESHaKwgprjX
fx0G9UWA1XqELd4i1xjwo71CKcaz2WauWbv0bsY7l2ruY1TmD5stFz6eQaPRIGeVuwE9sX+1YpcC
9biP+e57aTTfn41rDpKBQp86BgoXaNktBYkV/DYcQ4mXq/G94AyBfAPI+LH6GW6B5WuEJIqPP8an
ShCJ9a7twu1kPWQcA5MNvmwuDKE/fOC2cFcGwkmo87wJgsRX9a645KDqakzefZtxN1N9/zFb5UEe
3v9n3QV3Kk683g9YWU+U9gyKmPIQ8tf+zDWYEFX6raZsndKVvAhRjMFExU/fe/e3ExHquqmOUXW5
YMgR1H4KEMzf6i9vqnRFdrp9Ug9C8IVByd5/mE9NVQeg1JsW8zarbcVWAE3X0VjC+y30pcPdDXZH
6G3fkx85LJ/hmtAi5EKbaBVqNcwjYh3b/6T92NMJVrSB9qq0GyUclGVycz3rcaqFCKgYA6WJ/sYV
n9BzqYfq64svwo0zrO7VZv4T6gTR5fBxrUkgR+alkrb5jwY5PAV3G6+fkdR4+FEQ7FKcfWjBzsAp
mmEoKOS/o+GkducJ7MYM0GYq0iXVXa/ekN1qZJuuRtf837KNfOLdpGAlqcUID2uCv/lkZGMcfZeY
Ma8bBm8iwVEsayPyEyXTFWmGMlI4oCoKYob3WX/wc9tCFDp9iSjazrY3+IiIHrq8KNxJx5XF/X8l
gpXGMLY5E3MPhm7Y8ooV8haVvZk7KWrOVpHt2ajorIxvIHpTJlXF85+Pps+jM/aigCobRLvKaC2Y
73razgQiTYFNVoRIpSC0E3e1RvjxniUetO7fjLirYZ9O7wcGtBCAP37A01iDQCFTECS3d5UrOfsE
o5GQezFBp9qHRo6rIpygjEl4OXWQz71ongULMPCv3dRziTijo17obTk9Xv+wQQQ85Y9aQ8Ge5j0y
p2/t08pDGUHpEl+lOFoJBNJdY0rDV/r7XiQ2DuNu0hp2KvFveCFAkBrsxMlNpiB+i1qEaOSIZqa5
ARS1+eky/B6TmUNnlu4NKKrVxHFT/5TyW7uWAEKwVvjj8SV6sezMjNsDgYRltA+klyKjG0XkrxGx
Zw2UosgSP7Xy6+SgeB9ysWo3ZkWLqNHhfPYzUtsc2aT/4Ntku04h2cM7i8cWIWB9wlNZAID5GTNQ
iBWGYqEeuZeObmzljvp8G9Je/5JC+M3IPlSPlhlgyU4TLxMbRCgaHcvXd5721IQ1O7pUAPMA+B2L
IfJTsB5/qDTigCzajZh4yrA5L91/IuqVWFUYldxElQKTZ1aeJsuGo68IxT66MH7lzMJBb+2Nc5X2
fR7UACKuA22DPIdzBDFzjo59SRu2UGCAT4fMCmVikAjNDiHCe+Vx8yAwvUROunTV5HopMkuX/LZ+
xlowpYz4qZx2tQ7VHNoss37+BOSBZ/6iLDHs+yib9NMIVU0gW94Cr81by/Mu7WCLmI4IgYUXp1Fm
kTYBo2MeR8W3BGrTZsbsAvhMEOGtYJwvIUEfBrGyDTCfas1wl5OzDycy3euJwqMa3QC1c7Ay35RL
aFGLT7qVpfsegxyMaBQaoCtes1EfRIz9imZ9clJhJ4TMlKL2jqzcBhI9NMtG96ZHVSn7fT/zIVxl
KBpJy5KkxdWdvpxlhKJE4ECIx6F+MRsRnTX/QNKos7k2btsGBgeEvDrAeK9ZdUgKxYVuU8lySNEE
toazWVGD4CJIhRziaTV1dFy9b1CjZIZ1E5UpzBn2XTl668f63xJuTj8qhQlYPwWFJst79b6P5edO
8qBwv8piKJf9/nPcLanG6OctfzHcllPF1MBRaS7djEavf1bG0IiFvqcxw0a/AOzjP/jouy+jbFhu
zY1Mrvt/kLgZv9QLFh1rFrGZXzX5dk1dvLWKKY9w2Xud6GqNLhEZhriTpqvFdeCycKbBCpVaKvgU
Ixe9BXWP0tlrJX3vE9uhqJS+eILaO07ngWap0O/28v8D5YlgwS863a3Z87bC5VERIImXL7OaiOiK
zT4s9vKHy2jQnfaHcc1x04FYABL2/FvHV8s+3OuvxPo+K0D60a6Oq+tznvy+7fV+aFoRa2tiFRHn
ADCqHdfViUbAtK5s0DNPrbrg+YEn/M+JYUHUPRscNksz9eDUxTre8lx5hzCx2MtirLgZJtTo8jxC
xFznCaTsej2sQTCky0Adk+ztkdG/3L1mG2/p5zFdtfqwH2QYzxKbuKPgVWr9prtXUu73rNY3wTMq
7Aa9idqEIhTxWCDix7TYm4YaIetiQmI9HkiCmEv39kJYnYoSgY9hNymlF+e4V08y5ytN7lTAvQLk
ABQYAE4d0aTbQtVwlOXRUWABJY3PgrSGiAVpwHflgNwhahUyjzhoC/Tn0V1inIhTxv/1a9e5Xy4f
VI900UO23PsLqDfKL/aUx3K5nYWRtOTeCRH9H6UAGvHAfDuF3Zg3kPsXsKzd+gtJRPVr1dIsoL7O
OeGBO5ZPz9jjx/AX4JncHW4X3PPQLZXZifh6UKLu8i47gJW9NdwM5vHxhOJM/9sIhfTLrRCQylDi
Wt8Kx6zw/uo4GrTjGClLNWeOuI+5R3CxP5gdXPxkUsXsZG9NgzIK+EMSrkHxGClOxRUaeu6Q10Qv
GN76gbOJw9CDz7cxbvAUpFsyBJjNzoTeWAE8FiFwXvDsdaIRmeWj6s7tOtqwQnowxU6D4C6LYsVL
tSeL2c+SprIxLPIer2Ffy1zdlg2l8s+TjoueTE504gDk+/XcUSFjDarL7P1L6PMl+SywetWV9pdm
KKZm4+aqVh8vNwVNf1NK1FPpvIpjlNt+ESWJ0JTLvIjai0Pz2ObuuOZUvdGqb7JiNuEf2kWpaVad
2r1dVW374HqTwNcgQmWeDESWXj2tDRzf/jKbu9MVdqwUuCbxZyrobDUfP0NDez0BNiNA3SWaprpy
x5Fk6GV9alz5goBGfVn6Kvs1gxXGipdoS6+J/gLLx6M55k6vm+1h6alBqZG2hgDcPqGFtLKUSGlv
Qrz0djvGQfKZdlW7S5A+PPyjEPyUd4kPiclwO6uU3KTKhvfy3gELX2IZo3FmehlXr5EluqkM69Og
4+CM/0JvFwzDvvWkUQTq6ZN3XXrR2YaJCTGNm2OAMNiv183UnCiGiTZHGwX5OCKfL7VsPXFKp6Zk
hcXvmvxRSlOeIVC0YoAwwD+WoXqVTiIpbYtEZnhF0baNiXhnTdaV905dCil/fIKDzmM2t/9rvKQo
Th2BJrCPPkzCWvJ78eHx+rqau1VuBBFiuGmXvD3FLjegzVyk+vT9G6erPJ+UjKQ4CzcjBYsDdWUr
xefl9zPsxX71dlVC6SZfVImbEzE5H3GbDxFKsYzPEwxG58Rh94OhxL+YJfTTG784puRD7YEs28hB
g0ZWD4a7sbxLiaf3eaEASqtB9sHqoumgnwYQL2hg9kQWYum6cI9ZQyZWOGoTrb04dTY09KNgxE9k
1Ev5wBbo0Zz3o6eMe+VJlCofTuMFr6TUeIAYOI4qTHqPGntdZEIqfA9YrXghzvOmOk4cL10yvypV
zJgKsAbg4499KWE5tmNWRJGynmxoS5w39kkANuGYal3QEx31iJiA2sQQI7qL/KjJAUmtDu7insbI
RZxd/KwMSO3eQz5O3cfmC19Jdts1M4BxaiyJehlWSbyAiHPrHrFpFSRKORBkAuY6ctyC4EjisYhq
ceBjTx9N0nw5ByN3xOU06tTMqJqdkgj/hzJk3tU+gb8TQFWbriKDnlRM2jGfONVrlZo5UhAaTXeL
GWsFyXarWUXiRj7FyY/QtsWoCZ11J+GoZODIXdjghS4C9OJOpcV24UW587Y4gxxH4VPKfvrlhoMZ
QNv90RDirIzKvDNVeqI4xp8u58QNx/GEzsCKJIezYP04LtTAaowE2Hbs43Ude68J7ZrkK11LFgKS
Hg6N9YgZZ6sThlvX1gS3qzgF4jdb6eK9iLLYSmlrCj9WvqhP49MEF/hYwVaLuV4gAemsiKDhJOLP
CKna+wZYMaYhxD58wYoMgMKT9iIaAl8FcwQtcBrOKjVuwWdJgboUdOvoafm5yUrcN0JufEeV2PWD
ylFM0dylV/uD6r5IUabY+ZDcfwQULd2/j26HpXSyRb7L196uyfJLq7a6iSirhVbCdHgG+ZXCbqkG
Lpc5vQMQHMhMNZHpzLyI+ZzFzyUWFCjPiJJWm73+qBiAS5tEqLxicyYUpicyIVlRDCHmMB7CtEVH
F5D+JlpB7RNcFYc2wgr0OjOypWQJnsXSA68V4C5jQkiBqJCnik8WD0Op9vCQK2OQjdPowHAICk7f
eiw4Tgl+ZrucTaYbHqIOJRujX/cIhTXQNcvVCh4/Q6wGnr1CXvDFmVxmARm1TUrJF005ya+0CWGU
19QIJU8HCDOlI3RB5BM5BH2GJJVBgUsOTPjNZINH9MbcVtumiKJMmnYhZMZwpliC9hm5zfHrc9WY
12uKEac11VF1fGOcCvWqWW+BagH6snhpHCQyOzIT2eefz7GaCtaS6sA8B+IT8iSUuJqRPR6l2UR9
/WyWdMXg4DF9JY7uMUen0DGovd9n/JJDbyCSEN01hSptBsnO5Oc9oHpHWCbIfGGb7O9v2TcSD07Q
A224P/fEv/YgG7cXUAPf2ITYGJprADmvlbVLZtFweY2KkHBxLjL4C1JpgHT2a3zROCMDt48+ygOU
M8pUCyOaVOLv/uElTuvv14W7yqPUR9xmiSOGXwJe84VgyoLtSODvF7QegaB619XEZjCEMdgKdavO
BPedmSz6MeYB6onIQAZ2RhJslEwXu6GTThNUlAxojxpCF+V8UGcmzMSbCJ7KvgPuMXqJlzY5wbns
itGbqIlxEdkNyNnexa/qQhqSbcfVVhibduVp+vVA0njgANRsVhH/yzIE3ksutRvWxAIazMi+uEj6
GEiRVpUbMFHcUkx0nc3wbduvsmga7v2QQVemotyPmrn8EnGJYmb9APK1VsVh7kJnzMo6u0psncrQ
AFKWQEzqVEaqs6+RGHqDmB7e4exdmDu8qHuEgmz9729973UXx8jaDHwMu2X0mfx29AnkHU0YNqf/
0uOjLOxdZsCu4ywBZsraHOptSy0URL4Xmo/+SDDTkUEAaTWZC5kqAo/ir2z91clApYspqTmAytIr
D6qLEUwjMOkFC9Y+MY9vr1S8xHnNSS5gvpipQY/nC7M4XGl5oKrp7TUL17UtIj764NedOROyIQyD
KdAdp7EfmuoM01xILvk/DiAIMVk09LrZPPh2b9u0y33QuLzn7oqYeqvN0WUCgJCKWPgHAY6YBqIK
rr7K7tCVf5FiBLCdZ0I4T1SNYQ4En7ha7PDrCTRTy9qNo3nrMArW+k3Vy+bDUV3WJrEitkHef8rk
TQZG13ls2duLXRuxYOLPfH+42zMYN6FSBayNWbyl8Zsu1ZB4fVR9l1hT7VUvPOJ5P00pkkx7nDuD
bMsGQi/VvJ3w5cZLSr4/hyRUgxtuP2Q1HJFqBxRvDPzgp9ZqPI/qppW0S5tVzHA=
`protect end_protected
