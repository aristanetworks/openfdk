--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
GMMx/0jLB1TFB0qvQtCek2o0G9p6SfUFo4ySO6RCU95e/ZLb9dv2Pbi5ot/7H0m4XGvp/sP5Ptm5
Dx6xqn8vnMPgA7MFWRkBbYKzjKJRD320Stln7FpDbSwUIqm+RPV+janVMNHojn4zXKai51SyNb9n
cPM2EW1/LTTlncawZH9RYHuybsRNnvVUKTc6oMTMnk9gAYLxjS2zq+y+Wg3NdPMzAuk8N/SJBqER
m/wL/b1l7XLzj6InG9tooSP5c5c2DV6S/lDnc3aVx3QpnV655ipfeAJ6LT8x5zipTlKfN+zl0T9d
+A7ZGTPAhje4XyILCLGU028iR9542tYI1wBNzw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="XA8HiYE3Izb4dHrbCn/2YC1XTsXMN4qI2P2VO2ZCkHk="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
XT2HZl2AIyBKFHIwUCtLPG0mSoRz90BxrOgDb8Ceeymhm3XXjAN65sRg6UUliLh30ubMF3YzE4o0
xmFdBSY7zFCDfNgXdtWER4/idCIJqcaOhtrqX81yNj+CfpMr8tOyRzR7sMlMgXJDtr24WH9CUC8Z
mmbdsYLDQnola1i58o0LMHh3UxtDt+XoKxxXpWXU2uaUuHD5FSJlZSTvCok2Fwhqkt4/IdgsW+9w
7bRLTCJNASIiRT/S3PKS4tIW1eY7iwGd20TkZmiJcPZtxnf/OngrEfiagBUtRdmmMpdOO4EVyKq7
7tu6ILGuVagy3aMKXL4b+HpfVx9xLd/Dd1LdMw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="yBUrBWhXNXGGNHxgbVhiZdDMBTFJzAnBpcZQANBTUVQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4128)
`protect data_block
F+MUm02aTd7ucIYMpGrhs8NRvObbHmyYvELJn05ddvaHC8F3pXEtVnCftArYnqBKws5sR0PVCchL
Kd/z/AK5TOQTyAR+PUL40Sofey3P1SHaKxd29DYpCYB8bKEi5lABY5wLOiN15L9HBvCOvfGN1XY4
uZ0nU7TLdfz78UKSc4GFizPfqsVJHwH9Z5ZR4VQMlSta0h5MlHKryjjU0eIajaJHEBPCslaGi768
Lg3wVBKMK1GEExA1y5yHMD0RJOnrwKV+RDSElUZV4nZQAeewqv2JALgXqfh8un4c9WfZKsygsiuV
YQmY356kOsSVkizwC7RUQFC6HlB3L6zUp1fQcCdvKVrn8TzQ6RAPQyqEO6yvZO+O9NNzdiK/NUO2
+UBhzEGfV8h1jdcGNxv/wFEq1KdYLEmntv0twzMCNAF5Dr73nsMGsEcH1wefkhIn/eTyYT2v10O5
UHdrckxNos1wsswbE6cx0RGpEUQmFYbAAabyqol5HBTVGDs4BN2DdqFwh7CHRuxd0PVqw6ErIqf9
APWsyjUuNVq5wGysQc9f5OPylkDVG6gXz5aIpzCdZ4oOiuVdNLLe4HJ+bGFWVj3mtnWyTkARBZUm
jofUm3OKvPCLRFrSnEJ/V3LqtcVW3c0idR7tbJjKmXjiyX8joEYUJuusQZV7aIxRIFVoeyGROkTF
V3sbaYDPX/DSqyA49aUlWUgZrOTuxQ3r6hCQ9jLr8fdSd7vK8U74+IiWOJiSK45wtd2bUu7INpaJ
gyXwInFB6jhIYPz7Q0YBaycbD+PfuZyZdvTIkT9vemF9jyuc8bH/EpvKIURdvGvGIvNApJdEo/E6
HaP/R5Z0Kweu8tTxGitJVCy8xpoRcsPszMC9fASW9SZxopwj2+Dy1y+n6tEuAaQZ6L9uS5JPRo+L
SbvmJCpNEIHKVvu3IhepbFQjpJQrkviZBPjJNZCw/Us8NPKFimropArAd5pxrgOSsocsi9Tmysfp
890v+PkA72vEsQ0uoqnTzcQ6ZTGf24WFdmiL2lqLZn6D/H5GUiW72JADkybTS1Dofyw9dsSiSb2k
1UkTbyVK0VLWDxvpYc4F/J7xeG3IkVwP0AK4ny92kMN7MLF7ZmbH7GK3YkCf022iZLqGtwfYacc3
js4wf9+z5oigbJPj7n42H73z5bxed5LwZDZa017pZW8CPU2jWkn/nzT8qKoOX8VNjRXi22MG9/Ti
PlAL6MYt6P4FmltbZEC2fYEgq/kXf+VpbKNVzZ+5dTFrFBIKZRCAQ45zh5IP3U4sI7te6DwC24kw
MxTWTT6vbK7tvE3mclMN4A9zdlivJv2FwqV7YOQHm2flPDQlaNpx6gTVX/LWO5q90beA+qzr7u4H
KteWJIE/PznPWeV+0uc/P3CqucMhaWRnAKXFNzpRGkZPG6fSPN6ha8Spohm56XCkqN/20P2eonmp
KTcJRHwl5mksHnhiG7FEk/2jWPprgbRXiCc18MGLkD72XBR44tZplmDtK+RRG7XfCUzQf+xgNRtC
u9ijVhj/Ldw+w19wRbxh1KpIylQ31qwBck9JF6HmABBe1Eid7T8xMAIdecMj5mItyUaplQG1DPIQ
gxzbis19//F8OQwDo5A3E+0A8FmGZrZsonGvNqMsGnjUDKUR5Whq/1zNSSfQIr9Z6HXG1CqSi5hs
7uyxzUvQGcrM7Hz/VsckSlrLi56sEXDr1o4ZOchCOOGLHgCjFN6zoq5D3NjdwNsQsGZPRII+X2Um
yRfm3I7dyq9F22v7ZEC8yKjdAKgz2cnteH+OgruUcdeylXCyymLIPnTJez7WQPj8oTk74kQRoO+D
epmUExsQ8nZ39XsCvgqRAY9/LUTw5gSvjLQUXewGJYSzrx5P84DKi0/7p8bfXoghtilPvkihqQ+T
uDL3uUgHaFQRm1kGJbigT+fWWAuMKzeWjydTaNKe4ZDUUKySpKMPwYQ/T/WgbJMJJ3eIEwcQ4Dor
nEzYymJgVpbg7f3D33xo2u9sD2gAJntJXvyTGetDRPXebpQOQmjKaSBSRK+ffZL/0U4bRB9LQp5b
8qjRMXHsKzwZPJCZ5k5YkmF/c/nM+gWNNsYnziPjhF4xTTXsD6CklKfW6QtFd1PwiNz6tol0hc58
1asFQNPS02ix3KBMwhK/Yv0muPLHW15xFUiqsYmqI6T1GrXB0bjJoUYZCmMX0mLn/hM8OGlTHfAI
hbm7R4UJ3JG6p3LEOTUMzdTmcHPkXgdzvwWgQDhqYtXqSdYKyEpe/8i7e8iOcIHZH70dYkOiaHyU
tLkc4S4rovxkwoUqoN2vi6ZTvthCqcoL1Udv84NnyMbckWrw/ywosxjMXctVQ5KWXFBU3ei+U27j
A9z0oef2x2fr7wrFNFOAmcgAkSe7MTmEw/hbAxtPVLM+rhDYxoMIYxdYd+crIlCjC4pPA3PlhQVu
dWScU39F6xutqGYp68gEqFtWihzCv/nAmV/QsaVelXHf8syZB5QSrk6YjQZc/TzL6r46+N1ShxTx
XCVdyocFp+EfpVpVQn3qYbsvSAoUzqDqcZhxcp8tsDOzlLUmlEZRT2vhOB5JWvF1RFJFJZ0RUi45
79QRD/als0N9PjlA9gagM4mYyx76ax6bCUH0qMCRQy4Qv1xar9YGU2EJolY7MBz0b/3WehLu5d8N
YkP8JK+n8D2+HSdUNuW9QOfY2ASb/6wIZ7vvJjuQn/e7sB8dgaq0B3x2dqyjSplxblaEWYbY+wC0
oEqkUY4Ls94NmwMlcAfxTUT1F2bsVDFM2CxLg/4J+cGORUVmwJJP3EdmaMlVXUNfBIPZpbUW3ZM6
p7hYDacHBPqJjo/auBz2OkMlEjgpFFK+6E2OdcFGixFJoW3dg3FAmVXhmNUvG3oYJsKqA3t9+tM6
tdE9qfqWppe21fRz5j3wgkDDKw+czp0cB3buARvLdT6edQNQr8IaQ0lzeWCudKAgEXVVIWHff0du
H2Wkmi7JTX+zbw/jD+YdXyrSef7dLFFLrC/v4SI5S0JG/R75kI0F5PoH6kXVJbbcau+1k57H+1Wz
gYqL9tCJqT6qtZYN7mqw2uOJnB5t9oeniPa+8UVeOE1W8Z0Egc6s/uK4L2D06GfX4RcjOZlpqOzy
5scjQ89/klIuGS4TE4SUcgJoBltOBtp8tl/Laiw893yVFkOpeCYzbzW+7Ra3+RUuPzx9XRQie9bo
F83b1jD1y2resqZDQfYsM0KCWsh0iBGkoHStKjdm91Bke88M/88v3hjaJ1rflvOYQfhqPBBv+q45
2UX2YgJ/WmzSnkE0wIB847Gt0MDrW9G0ckG05vPPz4+9JX85is+WzioGOQ5EwVc7p2dIml2AgrTS
uaflWLnONeBw++Zb76VOdhReQFn7imtWJsHNGMk6+viSJjmHjAycmuB4JvRrOvb2Omw+/BDHo3xH
jjsCxVr7IxuIGczSmc1vkK2jdGK34vsa2Qy07EG3X3R3S5DiLe7CPkKP2gmmxH3tSIkk1lBO90s+
TW3uuBfFbPW1b1+ts/RFjJ8J5EtsmfC7oO/+7jwPuWz/bRXWFPlufo/07CpKpXs8aK3DvECILnzQ
saAV8m0BM1170ZsJQBTpxPTTEQhVWVukK8cX49gWshkebdF86QPe8k4R/y3ovAkPbcoCqy9hnvY0
Z2xBQoNtzCMcnvfHzXc5Y31s+hi0+TF8h3Q54YB2dExV7XumaW6vPPgi1WjQ7bScYxShzdhzTyNA
QxY3YVLdMw6tq00qEwJhz+JtimoqTyrkOme/ztnEsYE7RvzhOcIDm3UOczgZbrtCuIpMscJSkhld
B2iZUpuiS9Fm52hElTwL/2GoGYuXT/zpLg3owTO3/nkyhIDMc/2ZSUNP4IXj4kZuV4ZnbvKM3VqG
m5XLzzydw51TSH1hsJN2pHwUUr8ZAlu69G7cH2S3uSa8XpuYfE48H6ApdrYRlolcpyWNd607PTrt
JZWB8Aj/XyBAKU3TUPOM9SD0p7P6Wbb5pX4uuoGVHBniL1jzYoCalJKd08wgujyfDdHHcuvaEgp9
l6oCAlSwdjxyzxwZjI0r9rGOJ/F+y3nHKVfTxfqXfjtZ2pOKRDOY0tMxkQOhkmS80N3QyFSQfp+k
Ppo3QlTMfYGgHtQT8JX/pGhHn6gnxAVktcvCVdRpS9hvb4s8E5w1ebBb+F2IdwqBP2eFM+6X5APl
C506xOmjqhvWO3jFamcs1F8b5/+zr+9XsapMNDB+R6Fdg2fElDv5dy+MnaLQ7TpoNo1BUMGN+I+C
kJ4z2aocPo7BokMccGYHecJTnXV2gl3luqLoiJM1vnV0HmD7URTzMPaTXjhMqH064fyz3hqhLkML
WOwLOpZ3GzIQgLwjNJj4Hx2PerjUmhMvTXROXwTRDnCDhuuxUqsRNndDnSSXkygAUK4Q3F+rDm6/
2UE6VmRMrgHLqw52yZvOuTM+quGvdFm7BEbd4ngGJRnJ0Gv9iwhZIG3xI9Djol0rjlgBEN9oc0L/
tpqsQj9W7UzQdX9HPaf/WMtGY+kr/iq/lhlCEzDjxWgVL+go4OcRlPS+/QdzCCzZ2AxHUpxQ00Pn
zzSS1Jkhj+d2/lRnosA1/qRoqO5ubHqUMqQVz6ACFjQLyCcEPzPwAcfAmiitSijtB5RqvNX7DK77
bVK27IYZNevBuEMZEEOrckNibW1Q+LNjwd7JrgqGJeON02jAG+/ub0G9FaXVDr+vkZprGnFL3+e3
+vF/l08AitEdoj0KG66DyWDmfJQej0PDPIqBsi3Cf406SlavkKe+MfetmmUkxoZsg+OWql9b/02w
SJLKRAwhGamyvQ8y8u7oq/MnUgV8CqTjBHbvPB7wlxLJ9aS/o4oL8681Ho02gw1WtYHYFsgJoyst
dGKu76bhAIfnVrS1omu1tenAs/CCshFR+aRWSP06SI4PQRho9Y+sclNHHMpiLnzJU2lwuzYXhcwm
VYdZ5f2l1j77BXufUM16b6CD7+dT5riDJuGwycDAUjF2q+Uez1h8VymhEL4figa5pG966hCf0NYf
aSwV0p+kE8wUVyVtZaMQ4vor8dDZzC2CemoLmHAFW6xMtvapsoglIu171bi1bZzSuwKV1rmtUvuM
clbJ2phAeFNzyiFv03doT72SzC6Jo1akq4f0PRR3LQkE0jxKjGyTJ6edbyFpcaiIEEDsHBG6TjNj
NGdHI27GBou3Dr2xdnniCJmoRBjfpTNV0DEQyd3JNYbMdn1j8lOUfBkBR8q3FF5yrS0pP2GjtoKB
PUYuCTSlrve9VOeM1UGV4OlnPYQuNOXM3kWgWBSLLL/dD+FZMRAv5brICLAp+KkWUUq+U/BzW3vw
92H4zyegP7awSusmQh5391uZKhxzNGXATg6zmdCzKW61P+k0RBubaK5Y2nUTrzMoctuY5ubRZMAG
XyzgI0DB5z2+YX5m14bursvZQtqPsw6BqGMTb+MeN8jOQGz2EbMmPLEVCVJscGA6UzZ9BaGbIB1Y
e5om70x+PUzclblNw4FXB6r+Zqmn1aR6
`protect end_protected
