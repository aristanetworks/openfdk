--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Zd6vBqRL08cKSFW06v4M6GSZj1/tN1kvg58I358DsDag+JOzCf/KMiNmy7LVfGi+2g9B0Yh7L5xV
4BDgOyrUE4Ud7rdlqX7HdmgnDufJc+tKIk+lK1MHZyHjIzMqeq/PJzBqGlPAxvjvNQKvrEZ+SP1d
P5HSqfRqknZTI5zQAGbIgTifj875AgZ0G2vl4AB/Z5JZ118Ea5h6oYipgcYVSPez8w6LqxJ1+cAv
clnPp6KlmN46pTTV+g2qHMDSKc97r+X4NNvz0nl7+P7Gx4KJNQwyt5mEyTZatttzADdD45xNQk+/
lczDtaqNeTBDLFPiY8C7FvTstZiBTtMxc68HBw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="00KA+yj1d2QjnxjyUb/Ng3KD+qySe94V0DiCGZa25QM="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
PdPCQx4olA3cDod5I/2/O7lanpNu3tJpEqFPqJZyAq1T4nQnSO1aQSGSCX6JIXFHjNii8rm2Yaxg
W5QcmHUL1DnGmPoWTU/oERuGmzy4UANIWsvbPk6E9GP51n7MZw4AyRl4hE4ixy5BCEAJwLWvNGTl
dBPpUo3wmcgblVuE6hC7Lcakkdc2DZaKTryYTXNXAy0mUcEzMn8mE7SKQt4el1ZGH36+mRSkGATF
L2akWXh4Gh0GruMQHGBLNigbwIaDOC/r2XLmCGvnwbD8Mar9hRLS3YJQtE7gJGg/Cfz34I7NCxwa
zCPGIo03RnX0FxBSyPm+c29kSmP1GF+hi8Qhfw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="D3EptQ6zezAHGvLrgTwDZ4pMOJXWbqaUSQSvNK7WWfE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5616)
`protect data_block
/HBHCcKSlkP+pqsb+f8nfJSGmyJvnTXJt+rpbWboIcYqQKXye7H44P6+hdZ9eqbeQ3D1Cl3DEc2B
bamCEGLRcg9apsU1FoYCB2ZSNbx24TPvnEU4PROw70YELNy7xO1B2Vf+asP7PSVgofOUBmvOn8pI
h4oIIiiZxKLQ9YseqAlxAFmJc0yLlI5zMebNAO530UqFqIHWnjjJx3O+3iG9uAE6MITIK3cwjlnK
I+ICrT82XIE2hQrT7VGRW0kYGofSH80qqYTMOiS5gq1/By1+o+O68HYr2Ww3Sl2NwJVTIMzdDXH1
5XWyYtrWWkP4yDVM25+DA9gArp1cwxfKfKWjNDCI20aBhbATF5IPs5tEQI8kqDuN8neNggAejHnl
YNdTMNlPWc0/xEOh/OoFQByNtZrTz6Y/jkSnIe2jaVrbPmIkamvLxKj4C21DcHWw/vv4C/XLAKCq
+aTRQ+enpMkg4doNXiH/J7mx1LEOhozN+d5bIksXmwmfPXIXRIIpiV7vssyzkIWdcN5WwuZD57bd
5dhPUnwoAthRY87tCNlFpL4crM68/9HJWSLjRzok7kP5S1fckQwbtT6hHlGEAxFeTm46hkvlLImH
n1FLEGWP7PeWthVPMiE+wuk5eoTZBRTSXSYBnh5zhAkgfcLsGy+WV5rnmcuwoQqZZ3/yJLTklyRs
dIr3a0qAo8BZ5q3ilA9dbvWVS2Ic/RwT59WzUUZotsxyEQjjJcz9pF5ggyDYWZ4VrPkXl0MVJr0X
5i8u4c795nEuMmpIVlDy49vzdd+n+QsH3wBm8YA4iGoXiirmvTV0d9dDrHQo0NrE2QW8J6Lar0S2
lwzGzdCxIqPhPkRV5oWzXYu3Mh0xtBF0c2YLbM7MMe5rOpq8JtbRETnTmTAn0RsdodSSUEwSA+qh
NI1RhfXU1SR8LgjX3KXfEsGuwS46C+IT86aVTen8J9GvKWeAKwFi90cbdA2UmBrikpKqLnOeNV/f
z+7tbGW0xgt7aMEwAeHYjs5U8I6S3JjT3rXG4Qb+A1O7t0IsQTUQJh1pRg4FkLP1qn64FgmVghPy
di+dTU34ldVS4U9ndc8RBYC3wagLwis/+LBtuL6xTXDIQhZqYFEY80GoaUjQXrdFBVZnYoKAuqW7
03feX4lTaDUiXbIxGb8Z4RqFQHPCMke1iC0JCdlafg3cabRH0xp0OAGJQ3pn6+uBXZKr2D+QNAbV
Uole0WEX5A40ou7bqyTQyZnR0wedsv2kzV4+IwBoR5GFhcfVwBdJvFmIsQxKxjdN2GK+t7fZSKK1
GNLKI8Dvj9EAenpfcsHg5sQWXu6ZVEs0eLtS8awS5JUpcl6qecgxlIU0Wt9OLJg2GDjzISg5+Sz9
GSEooalPIox0tXR/iKoCwszpLb01YHfkNPmpVDIXfrVOB/PkV8wXRXh2yAfYnW/3rT+f77iHFxt4
MOnTjksBcErmUPJr1xrB1gAZAZGXd1wYe9AH3NsxE/XjILwGlLusWXz3yueglE3TO9u+rWwex3Jb
fuLseTVA+ijg4/dOps0qA2LrzBqhu5WWQHpJuyFtwdV7mYVXTrcSUDIe2v7NJMsaTgFgyfOF6Y9V
EA9+PGYzdXp8UwBHax17KV3qLEIvcf2APqz2QYCjE7V1cbdxzKeiRV51F67IxBhLh4fuFWMdN/mw
avM+U7VPv+s0LH4cZ0RoijRK5XkmKMm0jHAd7TTxxd9dc5h97oLPA1zO/kidc0tfj0X2plfcbLjM
cbl/58osY5+Ynv8w+V8BSFshyV/dNB9F9bfCuOYks5xUaCnhVXhqodGzPnRjbuoyu33zPLZ9PWwp
LtK/lg3QXM+qpayw+Iw8E9c60+reU4dOipiNXc786Jb7/zrq72rCo3hfyRGW+tPdlHxwudq1TSX+
3oMI/7jbOzpyHoT3yBgJaUpsiooiY3maK85JVZUWKfrl5mw6uSxFiV9r9h2lE3ZiobSz0YzHvFp/
oyknXZUgKZXnbphusR+HP1ufPjrLL4x0yOQkGUiiXVz6ohePQy9985PpSqD3ucXdxAveTQ0Qppmn
EsmcuFNv29k4b0pRiLG44KTxYK5jHGAPXfkDSN56FHXMOaxnjaTQDiy5x8gbVIOw4+yapt4QO9RX
AHO5cyo3XiJAOL8BgBv93LEEWRdi5pdKVV4ichX1Gqyb1rIXm6Uw9T3ZM6V4otlGGHVs4jgQOreT
w3rVH68tzVzCSih6NGbn5Eff43HmktZSFgTmIMY8aYM4VGMbfyAnQZzQRutq0wfHBG02rsAMU9QL
YVYNlO3/ClMNq3qf/z7xphmRbBFDE0PvXYtvHAU+is6gnOxzWumBbKQ0h0KdK4OLABTHBFt/1c5G
p41wDmgegIg2DFExLr+xP0I0Jd61/WD9L2vDlm7LCcNlKI4Zd9Ae1qNYhlX+Sss319kw88hqZAp7
hi8rJvZ6NXlWhgAL4zior0PFdGlpdRNVJlXXtjelGc9j2oluBax1E0W88AIQLu8di1DW3gUu3+na
XtZCmgQRuDR/e3jhvfvk95+2L+LNN8hEAhiHUZTfXudFfXA2PMcAcEm2doY5fWH6zmrmppy1taLt
pcl1RHO0ztF/Pg8Qo4FkzmBBX6p/HPcDfu4/Vv2mKkdHxAgF1iqCLaWyDgVoVL06cumBnG9R3ss1
deP0mn7mNOxJn0McyE7nn+zYD5OJ1RJEWnNGqOzPEhNqFe/i3VWBf7ItQ15KKlz6Siv0hmIOF/Gx
u+KD9SYIvfl32OhrR/T3h+qh570dpdEZkWRnZA6LUCrHuDKrkjZMpHSXbIBiTCtHozlJDlkFfpbj
JVyvahShgEm3xaWfMT5W3K+PRPmfkrbEcjPFs/lw1gyPkCq3sj4RCO2LVG23AICq+ZSYMWvIRB4+
s/s8BwwJEutkdGYdi4zTiZGxyfxY6tp1lrfFLXMQbyWTS9LugXK7xVEz0UGGIQh0xNtx/3HiTsEm
DnrOshd8tXYEd94JNePPKrWmn4sRDj9t9wSsRjfyb2ArAUuQQMtPpk6jKkdDkiQEYt3wWgHH8J2g
NyCvH6MVPFQ3Rh4grAVA1bZE1eBqGYOyz4todR10P8Z8nafCP2U8nvP0YN1VH7/Uko42qcpWd3ls
H1/EUW6IWYV9E/zgjTqWCWrQxcHfEbo5nMUYvC70PKsEIECuaLM8MrPgh6kdjFC6kq++QHTgtWD2
VaQWN0ogeEiHG9fOVxYKa24cGckLd1yXocv1U+Jb8XOGYqQTf1WwuZDOKOSjohPHUtE03SXQaDM9
SxC6CQypOjgj/1nLVG8a681IoNUXkYjyJmKbOkqNnReBZtR5/5JU9Y7wqpJUb3dGnZfr39aGNOve
nIYH8v32B2mU030URW6j9+eTK/HaEQK5efywrFdWq8fOXXJt2h8GU5B1VQhPYuEA7yTIyyYZYJGt
tA96Xq0G+4aGyHuL48Zr+71e5sDiwtZlGfdnSUqqpqCHeBnX0gkHCSrE3zsQeotRDdoN4v5kPpS3
36q/ly8qMlf4Xa6l3iMMvIrNSuiLSUTvVynja+ElV6nx94yyog+l71oObjUgSDqqpE6x1zub/V3W
kAgO1V107uofSgXbYymjLB7l5lCxLnze6RG3LI/90SkU2u2LM16FZfffGAMJaaKffEYFcXtdlIYl
+008sxPAuWhjiqfk4ehNGuPRjlUzPQQbn3TaP9Gi2cdtkc/38eOSRT2OxIJqQ1SZWe+opbqQaWPt
xr6zyuYJumTud4GiP5GwglAnBSow8hdZfbINFczU3hYTwOXoMvR7HSlz/rjbjYk36Re/BipYSQHx
K/PXPO+055T+RkJ4ZSBCTqH7gK97MlpuT+geKvgBUXi1t6DzynskpvpIOjDrju/wcw0YaD0MewOr
c8rIZnTW5JnVMqYFRWrrK118/8Rio9ilSq/AKb8G53qHXePnvvtoOcHKszUs35jLv3PQgOr8Mnbg
fFLVP8mk1hMw9wm1GJ3PiVr0BHbDl9+MViFhCC3hT9aoN7tVdRvj+q3y/hGKqnbc5lWN8OhSXmMQ
oTd6mh37aL25DUFSu1WSXJcEYhyepjzZzIinFsqk0xYMq1+78tSXasXfbHknCnbYw6U2mf3URVgX
zOE0WMc9YQBVmo8+CK8HvH4h1BOt61pTG51dnqtgdD1or+Dd3eEkmnz/dy10ffJpc5pMsGSXTwPB
2gA1s6mlROlNF30PFKPG5x1BA4JbAIzLt9OEiPsIO6a0uGp7byUGOb4n8U1NlGIa+r+EDFdpB46i
d4NC2stpNe97I58ZuCFhCJ65KVnQXo/9emjC8E073gbUSSEezzirQIn9E8fJoJj+Bk2smuAv2+g/
qh9IYtWLMu0eWRDgy0de+R3u6wqiKsgUlAc5aXwhMGx/izimbkQtrTXX7QI8EhOobw00m0FOU//T
rPU+HLa8Mhuh5shp6l/KALI8v8OIkzcqurzditORONJZXdsNQPDnBNaqR20kYt93yVzXUKHEy/C1
0XemCW4MSOsz/8NnU2xztrkYbCEgw+OCbrixf6w8Nga+skM0mgo8rzEgXiuJgOBvaovOumRFHRtl
vzJNgCZ3JJlg0t0X6O7RClJw6iNJC1CzKpl/5rtNhaPp7mKn6USP37cxjNtBhZTaWnMvGfRYRNye
VdxrGz0nRyYDQa5JpoI5fAC2T8aOn2u/YJPcHmlY1jq+U6pK7kNMhlHxrORm0jstbj/5OpNLUgZI
+SWdKdE/o4FRnXBvd4gRRmakQrm+gJRYxoASfowtZCxFFYWZ9c67gDF6rh0bjZ7nvyajDzmW3XQY
5PQGhgqY8vUN2LkP/PscuGslT9yc1xPysWoN3jKEfD+x7IBNrr2NwTo0RfK9wg7FZfljHJHKMNqD
0RzBzan1gGiFgYPP9d4Mhqr11pUfILaYIj1TJ3kqT4uammi4lWsTFTLAu+rOn3lrd/6COw5yooX/
ysQHqSXz6C7nes54omRn6kqFf9PbZEXdwsqBFfJMomT1xLN33xkRbcCx3hPCma/IUS7ysLSrAj+4
2JPVtcAMDKJboF5k8viAa9wi4MzRnFOa3oSswIETKwgelxdrRP1DVIhUDtUbbA8qY4KeB8/NHxQZ
fvfeT1xyN5gvQywfiLF5XMdCSeXN8+69uJm4uicva+HuhJE0JATqcSibntzS5Ep4r+Yr+9espxgz
6qK82Tr+gg8p7yUVMJPpUaEn8aXbRkz6g1TgTzdIPBtw2uF+udlyIIN+4+HRinhcUB5oSZU4LA9K
gFRzzlc+4yvq6547ycjpKFOAm1ets9OBfghuj+kpCfE0oNcMQKIFapCLafg4Tz/jdWro8m9fRma8
Rds3G40BCWyuEfml3fsFkkn10qaJx49hFEm6s2dXHFuDiMj+WaKze46pN0pJo/O5MSONEjul5QdU
LM0uXoY+ku8xrRjZE7gimXZIx6KOepyU/UtPx2WdvIdgu/ygnD69kYuGxknkD64WHYVGputeZUyf
P/S2FdY1S8UsC58UCX7NTNqi+RCYYFkspwAZa9C15Xn3OcL7l1dfKgrGwrnIjjlBYL3fI/frVxmT
qMdajSErCGA0TeFh0T3JeFqq9gAgZdbj9/hpdqZ1OlYF+SGsa/HIxo9Z0yCA6ERDBnZcR6LK4Rmz
JoPPPwEIlpi7inIV5vzkX9zUXgN8xjVO2AQryEow/3A3eETYnQh2Ay04IX7Wys54xnh/ZwkcPgue
AjODtuNd0+tiDhYPgOiuRJt2ummdYNFi8Q6arnBvhAL+Fanjs/kS4YZdwNb1WDRraoVhgDxASiH9
cAXBtV1jkh6bYzRP7DJ0mCUpcw/Xbt04yacM0U8xp0wJaL1xnEdgqD78+gl8U3eC4+QqTKKRD/4H
FAI2wugAUWKPC2aR6+SZGqWPIjaWBJJ+RsNcdrIJI6ewqOHDPvT2ApU/6Rpf5Ru1N35QlXwF/T2Q
vB8kxVQxdKeKZPIKPViO/idfJQ+CXVVltE2uyXg9nRwONWXpoIs2HuD/C/eaJ7c7zk5MifhM7D+B
LNbPF/nLPMw2DJLj0OWJ5Yh9uRSeBwgEvA/rd9BJsXrODiZKIONx+ure8/+ysNwwIXZ3UjbZoiCd
3TRYx8vXvP4+s1gpQuIejeFBGoDpTjPzfR0CbUuG5qwBxRvSEmWwvc5S1jdbaj+fXf/F1Bpub4aW
UudVQFqjTx1E9TT80K39ljg91744ly16Q7GVVe/i6ohLprKv4Q3pi6UMcM1GvoW/2ySZd+qn6y1X
4zlSNjOJFZH/rLO7n2wXDSsYt6OL6eQS+CNaRSYyw083ziBqj/rG9VVulAhw2fE/u6MW5utxCX7Z
adDVD6eO4nO38qhRkAiLLa3fWB+wnNsdmcRG6NdFp4tf1Z6HCKWBl/rM3nygUbpeOgJ0HZj8eEdu
X+SAqLg7nXOvkhHYGoPU8ApIFWTHV0skXVOVXf+hhN6Qi+v9ZT0EwquhroCe9/RSCyyObIUGF/eH
DN5h6Pmcu7/JzTEFFj3ayDrSBTa/rI/Yp9ljR9HTHOnBPo3AoYukcJto6MXrrtnveXVGWjMWtSR9
HQzQrMtXep70O/RrexzZS9H/FF7IDnMIyoa6ZvR11avxD8lGl29pfpZI80lPjVj58/10a+yGIJwv
aLhMPcyZGStM2RQs6yShLpfp6uDg2ReN3ZfWALrGbrJM7lwiuBx1K4evmvMwFLuDFwB4YdMb5Sss
1x0/S3Eedu0D7pX8OAcZuo1fYnDpL9q1TZjzagUbq9j5I/ofvpYLGbE/yomG8qOQozFrgIvTMS2I
NOs6F3doanBe4MqZB40xKPo9Tbp31QdaDl1wvRCdvmMoZRQFzcET0gmdn1TD/XinTCZ6d1rR/XD9
cGA6X9GOiufK8MsHetaDnIt+QcXh7xQ5W3RPX+m17lGN2dbGH0onSTijKYtrXpMqBMt4gbByyULU
roNgDJjge5w0g9lHEgZv+zNBkHREMHKq3XKyaI9KrKoYL37sQ/OTeGcIXgAJ6QfwLd556qStEw3/
LPw2abupK9N17rRbbilhKe8H365K7Gu5DMA/E49F+zKGtrBEykJRJFdcrIFrEze7bQOyYRsAWe/h
fHAzd7m/Vyqmt25FXWiik5cLB3+4fP3Yd7ZnO6TrtS7fOBR42Dk6yv3UFTw53EY17aMbh57ECb92
JDmwOI4NjuM8DKU6bV5WCsi2cHtADFCYdGGt82uo0wpct5+ALRpr79RIREjr/PL1nBGaUg8mU39h
LWqP7tvo6F71wGqWjmUtj+ABXktb2wSWjXGsyv+jzdhnjoGbIf85VwYghyWnKm58iRzgHGoQZf7j
JKXhy0QW5UoreRis7HklxcU1GJLlVYuLRW1KIPxcRiaeFsb7L/ZUgKzXVRXa+xKrQmsc3p2nhvAY
igTvDyAenqKhqAGHwc4j2cP9b8e6YyqhwMHtIXedcjZ2i5/sLaNMHC0+NUHQ+xZsvybrKKQ+pE16
jflQGZuT8BZNlAQfxnVHZ17ZZHX2WNridr4D4jn7
`protect end_protected
