--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
DSPSgprBUKPqF5UTUNuKwLuqHi7A5GMCeyYiS6nRsCFTrkvIsXa85O+jzIPQ3IKRrpCkiuIZu1WZ
p75vkp2R4TTO0dpYXDO51wek/v74PCDa3PoDCA1yl8bNVsP/iUB2sPecjyT+JhYltxQb+BM8crvs
NJBqltS233s0gm2kpNB1udnXpsmeF+mWjSGSLTRo43KPfMQfjCIsYQyKbWZMAsdaCZGOdYjwlzbt
22VswEgfqI1QFyKFtueHx60RsXZMUAkKo6egSoJVwjgf4P90b0UGtW5gqqeuyytEJQqlncbYZjB/
G3b0YSu1craMk2Y0nYPiBHXOxbpyFi4tfwxw3g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="DvFyUAahdOCtkBKz6g4xoXqkI3CttfQm7qQoQSuQOqg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
iVMgwp9RSs0fV4cdCwkBQLd+XbHK9cZS7zJwacTpaulpMqwuIfT+NJZ4CABQ5BKQPrBmvHSvLn7/
YSGdHUAFadHzIDI/HY9TQmpd0ELwCAzX2fLkO2hpAbSRBOIPqP0Ce+Okn3DySt+NoBBahpo4IvjQ
hVVFP4HizPf/M0M8GiarzaW+JAlhW0Kf8Y47KTQ11zBo+hUuY9Hy0y0fJh/9PTiS642QteEOR5tc
cokJ4RKM5KaLtnhqM2f6Tru0q8ublI0mnOVaSgE9Vwz9BrYFWXBJD9hjIz3m6qOpzX16wtw9kHIN
l5yBxZy+bveNeKdYhnlGf/SGRrCFvfhp7O353Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="iYhxywQTR7LnXV4eBNJjapyCiN62rG67Idd2uGkdA+Y="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3264)
`protect data_block
S+48r9iF00nhs2Vvd/IQwrEvqx4VwH0V0PUukH9Nby4o50zO/93fPyKc8sfgTIsIdMqIHhRd4TG8
AHsKJ9iubDce7/TPtk+AYgcw3jBad5cuVvSTO3LlykxYppfTb65Xo9PCJUKB3Awi+RKARwizZtnM
3gsqYmMzBg7ZXTvYyoHc1vacJ+To/zoG1Rv/RmqEG2FcSerhn5zEZeBTfwyDFw8Id0I7U9ELXKku
Ae9sMyzsxfLzd2X5PL+ZBckeio0/Iz2kx4n8xUn5XW8w8stH66e6aBbddX6PUi4w8J/KW0R59qrz
USkJ5w6BVITitDNWPuTbicKUSKQRyJnZDxfnrdcTXy8chEXbR/kWqM7DcVJkgij+NrHP5epvMwra
raQbHvq/PmkjvMep3wsq1xcPcQ6/EJVxPgVCA2XXAEFr67rdGi2b3Rn2L3sellaJrN+dcemSLFBo
XWQP6xhNYnlQE/noUlKXkJJBznXdMTw1pJvgunCChb0pDfunGrEwjIyT4nEgin3WzYBt48BljdOx
HMNA/wMuR9S6jWSf6NmMDUxrbXuZ6GDUv7KyzzSxvFjWrlMgNvOrTFuzr9/5oH/5vxbyX4Gd/Yrr
GLAB+KSi1nZQ08OtkyaD9cbQ8lvwifSfNk6sAoSAoYHkovP2gpPc+69/x+qV/C9WGr7MmmcMadM6
Uxpsn6LfqLYHc6Mt0wo0l3TYmrB080sYwI7lWelQYZZD0ff7BVdQZHF+aQXgG/Nf6n4JTEzrbDzB
jvMpsvmqLk65+A/oxtflziQSRD8to0jeEPI+hyzlbFuKpoeabAXIsKEnLaH9cPM7+Tv2Warl1R90
S7eQmVinPuNfp+P8O0eNepSfHbOQnm+zNCUSCEdm2j/SF0W8VPi7TMDkFIqQkpHQHeA1kIOqpcEa
01W4alVNhGD8kjjNSYR3IpOIFHwRcOPnEJdTPNF5ulIjOifCi231xAWqoN4zjCX4OQrKcWpMc+y4
S4gpL0QvvkdgWG4gL3Nk2s3aklipI+MVQLkPVDI/wkkTfhQHYhS/PLL5gkJvi+vvLAxaJwlHvkPX
tRYAdtLR43qTo5dPXyNbfzKVt9XazBbT6Wd06Loo9cW3Ot7CUUa2WbU26JL91BNWYEdZ68f8NcVk
Mbgp5KqbLwqDK+8EZ2PW8m7btxQA7WooX9ZYM+RlWE0ZBPN+mKW0wltv4fqrjXvx0WcaTBQGXPWJ
QR1yEXMmOR1B4D+0bmTJJ+CKUkUvPlhjMPHyJA+1s/94CGDoAaSPTcQntxkZ4f94tKzO1ae0hXn+
VRX83XaEQlf6oeN4cLGkDVJMlBVPRERqhKoQweJ383yOoJ3ZK0btb/wfYADZLf10+Is1rNntg3Ji
D4UmGscuLihV8TcAB44S/Nk8FIOjr5iRv5mjQOzlsr6AfvMHlxTknXDtsEAmkLWyIzJdOMsuB0sH
NKoDBBKiLKRLRPjO22hO2orM1C833j4h9T8isLIoFUb84dvBxbcJhZdgsiYPEaqeYFmyr1+QkT2l
1oI1Ltzn6W5cTmwXNOjdmSEcov9fqMJsMxQ0qQVSBHPTe7E8lJzTd0F0YlsxJkGDxocVHHqimlcx
/hEe6OdYa3jMzPWCScQleA/djR5B57u30WPvz20ksi54d0VBTRbrT/QlOpN6E2TcMiVmIoe/7JS8
nbJHF6ReJXN/Ac8A1paVVepz+J8uefE2FSaPk8ZDtkp0H92nW0Gjjn+ngIsVOr6RDN0EQyvzcEGS
+ap7U34NHaOdch1QjKYy5Oxr6qrX7/RAcdqIjvUiOvLAbdMItYuIb6oZb1my1DHoW3zbqONCvkji
Y4Lk7fsxDqCQuRfXNYOS72As4S12urcjCcMbCLS0D+zMaCpAzQg3OMDM+GXrQsVbfqKuUGg1FdKr
k1s/YJdAOCanGzCB0XiOtr8HCtKq4EPus6lHVt600cRZXFekoaZZ4fFWv0I3fZf+5fJVVPsn2dHw
/5eF8ZSP91vvbn81TB8BJDOQFZxtsCx6RZG6iEyOkEhRbAhDRo/cO004aJtUQDYdn8c0+Q5ze7/H
+9P9qMGeXaU645q+CV03ugy7HsG5gOfbmx56C5UCKGnlue10H2kxQR9fll7G0TwggscxXe/biM8s
4bcQK4dfn4hGaqki7I96/jXDVEe5ibcho8fMlWPJOoMCjLo03xkleTK28biykuohLMm0wzfdATR1
zxthBoLpdgYKNYNahGZNk927ZzFAL3nu2d0I87/F8j2za0TwMcFK83lGCrRL34mydZ97KpJOBNKl
vLaIVkBPTixuLxg+oRAgY1eTwCE4rZAbDHwuwuNhB7rYuUfs2PlwvyY1dSsQcHa68kluOJe8inpJ
zo9l14NE8LBMdf8ZwMjZqIluyB2QXbB72EsUPB2OvXhsVgQ6lfkQXyRTgfUUKofmxLJghYpMLKjO
1jFHCvpW6zyrgw68aJijMqDozdcNF3BC2CUZ4jGcx7h+5YArsviYWvvfK8kCn3j0JJBMl3M57Z8u
rtu9T4imb6EVbPtRbLoF+wgcNJvgFU3yVIrGPZhVea/lWOLZpLCn5I/aLA+95iDKckViwGMchP0T
PVI3MAblsRTkRmD7V77+pbKlxoUfdBrhCp9ESEtWrYcMNdw1Hvx++HQ9BdZtBnsWv5O9+NqGnA4s
eKpIGPPkk6+sOrcAPoCMuXx7JXCEgBisKBl4te7JfFneF28uxJN53cggDFCDdgQL5/ucMc/5QbpY
11dHNRxgDR+8VxrRqhhDzhmAk6xA1gPThC0VSeaCR97dkk4ETF1zrGRFwLAkmdavanv8aTHWltKc
Il2pFEzrzzKKP2dsNUKQKQyVovoeD+nY1VTHsAPR+r56U/xaOYK2DU5CWxtlNOOzEL1QoRNlpdAL
nlpbMn6dCzPOhR5b6ej19Arq4pAQ59e/RbgJGelgrnaREY1mB3+2i4RLx1JBECP59AxKriTF3+vX
K5OQPoNfcFkELyNocROyz9LhIsmbQ088zBQVxtRYGxxBclMGxduBnbReuUTlmi5zltYHL3L3iXC3
40yDKx02D5wNha9OHFtIYhrM/ywUqb0UjljsIgUHx7F2TeezUleFIj15HKFxIrxjoW9mc2tHjApA
20snAIRNvYbQjYSfbGqUSkikEToHBUMtsXedtHvTNiJPupXakbX1xRDTtQ33UHbm8/uX4zNtu4CC
Z/fbhVqVVCz6g722ZiAyfoTRJ6LLBc+3OJUqleFIXfIa+XhQbeB/HaioO5vhRXhs/AubXeCAmBfY
2Bx/g6SkmTT0Q3rPhFLfAYTuE5ahdE0EnU2p/3gMlxB2OHIZ61kpOsXZK3V4DAd9KYzqUmy9BYwT
M+JN68o9uGhQg/9vDnFMB+Ma4XfyG1cLDN2nj5n6SeM6xA+ObgQCI4GidZbXymRG4avXCtn/LHfX
WtkNIPQwpNls7qI8cQwL7THn5gWoByNVLHEIKN/QLbcn4M5U4ODHACWCeyYet1yE9djyjAV8Cov+
9zMrG0nwQ3WxMtvEk5TH0uiHRFydLRLTNi4yl6Ap+Ev1RmxV0OZtksHxsLzmYqmMjXBbgSrs+Vek
UqTirWhOGMaSH6jFDsZUem1jSXwlL5gRM3xxXCCRPOSgITOh7gyjCnvQCAH1soNMVidzSfBmExSV
dIof+QXyKXJ+ljh1OOPQNRxNjFzVY7YBz682DUPGoYnTsDW046zimS/xk+I7HGAAuy0XWXoqR/w2
6eaMAvbn22oEdN4ppX0kkgjZyGrd+If0oKYvBpTR8SdGWEZrY+DGX40r+1UKpHffBQjYHcflrkGw
4bqvbzmEDF5Ui362cZ68VQF6te484xfNBXmZiqKWa8/nwFtgudl7gJp7APiqeJPDBAlOZOHkZNLt
4CkUffUSe44vT5um1tWxW2TTzIu1hPhOjMNHOSEEo4xCIQ7sS08P5tLw9iFGChJxYmOFU5DdXhhN
3+Y1kEMRCuN2ldeBtnAokgrkqqSIx6VP8ERbrrXtYuTkosWcqBCBiRNIsT4JtqFT5Ydc4v6IUyyg
qoE4lFLPotm72oS9nqesyCtA9ABSEiZ4zW5BORXxyrxD3IyEcW3Occq05zoOzPjbLWrnPC5e+fiG
YT+VS8fCTwMtR7JrdkOEnsKujC8avHHRjG4eN8IlHSHo7FfKIxqtQWkbavSu+tovyCgxpGtE3kDQ
NrhErprp1MVAX2cw5KR4GrT625S1QupJNLyXAeYnkAAFKUAQA+ebsDvvvRDvH6TFOo0AaGG1BpIH
B6vBOSMvN2S9q4/OuSwHOhk8QDrz8bcGGFckSoqruXUUarIZPqU7EvVQQ6DPRf17eGhkmYHhKquM
Kn0Su2IN9LNhyj/Qyrp+
`protect end_protected
