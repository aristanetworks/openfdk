--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
mtGwnCaFTtDGZH5CbEuLLQoSrXCN4nyTOnxrKHTPvgptFQ605IIPTooizboQUtJll/I9e/Td0YUj
Q9a6piZm8/yZAsu9VheIB9Tmv+hQG+Y/ts7nSVRtk39OEGW1eVZ+T0V02XMlrw5/6nUPCnM8mv5L
si1j/EI52fHUpmdNUU8iwLzdcvV+UV0FDvoHBKR/LErFXrQeIgHB3mL7fZfSbVfExLGSRCMGtslc
Vjrg6mFD63nvIfmdj05OT0WM2lX5rTm3tqlmb6eHoGlM71cSGzu4uYu+lLMgvjZGkdOOXLN99Bo6
klgjD2OsyEIALoXieZulJLJt4BH40jmDxv1nWg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="UWMuXfDzRAKe6VImi/VX87XHCARa+HSiB5J/iG7ZmYY="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
GwUqlBaQ/znmPXFVmrkjmr3jsQCIpLyMYfiY5Kq19XTYGZYyQr+CyRYyc6su033oXpSGyiE9T/d4
pBLoQWn5HbTJc8cHGorgGdZOSuL64jwbetTk3qvDAnOLBERfgpIxSjXlS9jkvaJLWxdj6+RVWtXG
EGfQsZaPTVAnoYJp6hTBJxHN7r7UTa1E/2UMXGV6Ril4g5f9GhFgUfFc6/iCr9IEGZXqiGF8Jjti
FJF1WiXRDsNNxDc0LGeYHS8Y2vQx9+QcvvD3I8ODWNFQXH0ZIi2r8e2eSlO93NALM7QrOBQ7lzbp
wf6pYx6if7+mNYILTnAKIl8m6WTQOJaQi5vadQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="/iZwJ26unMCTHEXNVPghUhT0tcVc2U8qbgEFFpPsVsA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8688)
`protect data_block
IfqSyb9B09kR/EhvYhFLe7SJHDY1AT1+09XsMSd7vyYCBXmJzZgEq5ak6ficFnvEg+XXaN986dQP
srcCGJZcnhcpRzLa3YIYNlB9jJJ9TtVLCer0p6nbU8UmYTR6CZoCvtJ/FtsmuJgM54jReAOpYlOJ
iMH8pAlxSbG2Spr0AQrNH6FPoX62lXyPS9nbMlSKugaobqQkDx2A5xkhATJat0tO/0AYTWR1kYHk
n2zYQwcf9uGYPHd+Snjev/ta6sT9Y7XRQK+5q9wafntb5+7XIolB4Y6oJ9odP+XjKvjwofE/+CTr
eQFYov37zH7bQaTz/troHhu2NVb1lPYp1U7ox3xKX1CfTGd6Hy8YI5dvbpqLcqLNFYTdk1VJNvQo
UsRZLyvceNXRduojug29n1/NfwNaxbCaaooPt54CHS4A49Ptfj45U9rWkMeSMmqARoZyDLzqZFlo
eos7QlXnKo3vXbMLFJvZC2NONVhHbIgc9vjIOd/sc6DmKAHLG7NL/5z0lWf8Ovm/NhDKdKAFe/eU
KEnD8HIaeGeV5U+SMFyMx9hQGgHUsPcP4qPDets7hRE5FgR64ngx6iZ3/a23aqOLeKqukYRKf93Y
IB0CoULxJt79RnkI+tG+rmSolF4r0rIn6jMg8XMBmzxDoX6ebZeN1D4jVUZPu+Z+pbq9peG0a3fZ
pU2pHgXCUGimMyKfdFJjSiFhhMS23xH0p2Cwt+m2F/mvgjeOBRjPrTHbIkTzjVbmcsDs2AFeKCVF
1FiQHwuCTvkg5fOMT23ax4I0wwY2axkfIp0wtz/eY4EcjqGhQ264iP0F4r9eR3H5xHoeTMIbKCn0
uQzl5eEkDmPlLBPsh2mXCNR6BJsBe1o9OuZVH8RG4RrITyb8Yhq25PBoIRwiAw6PizGSngP8Sknx
5QLfshZuxkdhSplz+ZIOUEuYWy3RhXDx49cjeWjzZLC+PDPIuPG0vbKxGXmEPeMPWQrfEbzVFpTm
6AQ0cQKzEqgJkFEIimOiqjtWDMSrHYRk9FfHpScnJNzYItUzN5tKZSFkLfRLLtWjFnRj9X2Y31ib
xfT+vm9R8QqrHBW6nDIsWRHadkQHCoLUb4tgV3/ZSax91g5WctRXYn350yobGA5y/998RCJW8Zlh
buEJ97JZWSNphVzIGS3ulJUadTUj+tjbsUp6N5ij6lTAUTwXGCMKfvtshXns7QJZNNNX9BXJrCPj
XiMp6gUYEZ+w/lCk7sTe8t2nSEZsA7K4mw74GSougOyUPFeWSPeb923HjVwZsUWlSsHMLWT9++lY
OzR37xBXvSkXWqwYm4JSJyzv8Ea/tOk0pJk5rUHXi/CA3HIO4vCsgDSoFQEid6RA20NXPUe8dZ+8
/UupjtUjqCf3vuTzsxlv5vRANtljGI7IwjuAhd4OTZsPHzaAmdAH0WCdewAKUTBBGyblBzyMeyK7
zWwGUzAV1TwYK76CniOrdKv4VObAbFz5FOLX9I6yarRgKp2saU96X8NYr8bSvj6rLHAmg9Jtpobp
LKs/j+qZxMrdhOV2VJOWP2ACgJ6HXvmisVnDV6OxzfloEDodjSdn+TCMjhMCNOb4kpx3c4iIkbmF
BoK1YmWN6fpn5Z4VHEE1nmwC9Ehb14l0kcf/GDgkLvTi0xWofiN+QX5uoZfYaSLTKOHMqFYKqwNd
uD+s/a3IF5CLXprN/7UWDzoeHJzrLKW5ZWh+5Dgn3msaGNWdIQmO3Smgc7iyALtK3Cv4LFTGN5qZ
L7kr/p7/zWDDuD018p50prmgI1+pEs733664CLe+3P7RH5pdtvP0+Pe5T8KoWSrq/jynK8tq5DJU
DWN6FpXlUdHJFCnBSPR4C7/pXaLFlzBnlPmZiWt6mQ8voB2ftW3NMyhUbAFM8x7Ht+N0SEkD14C9
CZcSFk6U0vjmHKbk8DnHMCA1qCjeUMLI75AA3eikuyHW612nc9+hNfjaaUE2ten7g8ZR8W1QFVjW
B7geohbKu8H3pBnzCzyFOyh6ClMd+RzHsbXWBf/XYJZcWh44NS0s0Re5F+mZBsHBVYDEB36nvZRj
ajSg79JkeXdmKyXQajEpZ3GP+ZnvxUykxAKmv48NwJcFOQTU42aKv1Yw7QC3D9Qs79uWegoQzjQI
Sv/sKxBpME8+uWmMr8B+GJ1HhA/fB2wYBGR9iUUjlCX3XH3P3Vrc9RvpGI/bhj1yLRRbfI5YyV6Y
dMoBt4o7TuSN3f2TNrER/YV1/K6Q8cdzSmE+M7A2sKmq9vLj1q1tgflaehVoP3rDmM/fCAmB4NNp
8KoV1Utl1jyYS2nK4o/S3heuyx3KmPRO0RWQqoc7w5x78idjhzt/LDvEa5YIbgXJpZhrmlTJTvzk
mgF/ocRVJesM0qQEJWaTiq4BNH1WSiIPo7fDF1HNXD1+/wJIP4yNucOx8KvWs0TFVvxHxhwKyw+u
rPGlQdcY3QxyKUP/2jcM3ZrPB6bENPGU9DejUOEEZ/jonIbAjuHofz/cEOmxl8u2rkJUJ6dFT5lw
MQtZCN2f58m1TmH0WmFkOz1cLfoAnpW3Kc/gqsA70QKkjEA02Pa674Sk0GA2y/4L6yqj6hyb5S/z
p/+XAYL8LMhYnZFcV8srfFXiQ6+cHdP9Re22dut4zdChfXD+5cz4QZOa4GXLOsarY2+70YNwyyNt
ooexQWgCeRucBuasn/6FF2ZHX9O7PYgtaTTc1Qh885/P6GKu5oXdns1UtWG5XcsbPudbRCZ8BmNG
zghdZHS2UnKHbMdWeM53AnC8nI9pYIsbiGWEiRehIJbJU0i6Xo1dhcEW5APOPh+rbB6ZEfmcb6Te
vZsuICODp3+k9X3gFxcjuSlqlHTvBmDE2OQncobqrWoLIKpAMO7/ouy017y02weL0ExH5gc2Pf2R
kI8LjABMFTwXRqQIVq5khwlWuCRFKg2ycAD/2K+5My0IsChYxL/ZoKp/+8+cPkK5/dh2En49h9GX
J4pVhUY/Fw+R0gq8Mb1/BBjFe5bCeCkDFqdXBJXYJ0pGMjpy3imBtUmy+TbMB5zIdlFw+Fm4fhuf
bpj/0dgatP+dAT4YqHPPsiiONUnyr2gGKuAYEDSgfoX8GrFQsPvQyRfU08qC7Yb+v7ZY3caN4ghG
0zbihgvXqmRQNndZFqG4dpG12w2UYmWqra6907+kmL1dffsoJSqRXWAXTB7kdazm3Pf4cQBQwFn6
f3FVgyagSwJ4ittPyRwmi5CmPkBrXO0omYPkVHV1wdJfvRIV3jKbaLPFQqEBc582i/T0U5unsyoK
Et1zdIMVfUMnJeH9hOgieGHpfACq0g+7fgsQfZFcLaXNCFgPrYUEgzkRP70Xr9cJeILxDWG0xGo4
HGk+YU3Ku/Fw33NBg9yr3mQDKbZu3hZvih852o2i1MCRZwZ16z/jrYT/IhD08fEXE98iiQMtXY9s
Bwl82WC1yYGMYh0UARySOwre34aBiCJPTwA36FnLW0HDzL3mSFWj4sP94Vnh2FKYkjgTs7yEZc/a
EC3DC/ID+K8GQS3nJzpu+CFjWx21i5VrFXb3431qGAln7dUboUQodNNG8d1CzlFld+SGn+F5N2df
wRZ6irRjZJTeIGiMwNx/OtbGj7GMYepI6Vv2HJWNsTzqIBQAIfdYUJoiojLuC4Ql7K6I/GXOWCSW
M+hCcv0Lk/OSBn99ZGNv54JGUmFp2gz/bY1cl3KTt9NU7fnFMDei9jglbUO5g+ugmnJB+vXB78i7
eZT1rLUH+ZzL4VdZj+K3VCwvAl5o5zDoANGCOWqF2bGA+3zy8+FuZ/K5uh8MqI9rdAMw0MgRfBjG
UTz+1iUWJ/v0tU0WnacILBWaZxEY7a7dmf0OUJP+yL8DZq53QTptaEfLZQsh+qqFoLLYUbpXqfxO
fWvcs3BNPy4STjE2hKWvLEZZyrNBeBijkrdWvvnw0aWXOjgWMO+lEI373pQE/5CGCzqY7mQmf70V
7ZulLSbKE66vg3BX/q2QsvRsNIJMbQe3o2NDXolUArYnqVWtmhrkuQcujq/fGpXX7TkNJO0QrDOL
2/XLtVhVjJt/m2CapBRiFiu7LupxZKxi44gQ22pGDYI2p0hNKKWgriiSo/4YEHcgCIxKLrzU6Ycd
X6aUR4K97BchdhRf5lw4TLY/q+KhlR1IF3KHliQCsSEXHlXSIs+cxdF24jYvQzjRE078FZYIQLvu
QI1b2yEKRqMDCtkgJn0EVlNwY/zrYq1PsIcRmV9eBvpPs1EGOsZfA0IqDq5bv09AtTdq9xbmg2mj
EmmcF4LsLjmgKUviIv5IBqGz9R9HYt2KZPJrEnpCoKAvG5w0HduNohCpxr3n9Flt740B3zFP6A+w
BF/Cqfsd6CGvYrUKtyi2wFQv/3a71CGA7BoH1UapNWjevQREDwo65XAkRUGT2iZF63e8Xd9sDafv
r55sYAarwkPEXQC8UuhZ2pNPr6mxY2Ub7GrAwB8Wd1ohGyvguAYAKyX5dG0DLjNIArhnK2eSLt57
4ufD79FdPVriWxB2XVMeNFPHFtWeKvmW/CE7BW2+bAAmcLVf/1+WLqd8k7RmHmQUEaxDykd/Wem0
SaCgJryPq+x7wMw4v9uzTw2fxeCKXhFG0MxFuS/IGaOEWdIkFH06n7qL4BzCmopl/cO+y0GG6YZF
AhuRG5U637hxZdEwhx2cKHNmWleN85Gx97IazFt+sMNAfS86zw1LhISQnuBXscWKbNOnH2LO9rqL
liRmOwDheTcF5/6q3absOt1Mica8pv4q7UCuSgVVd387R0BhRselAsJ2FFjVdDKZYY3qxH/ZEcQ0
k37pgPhT4b0hq/j7xi6OJuLnnU4g0XEaxNqrL8Y0RL+tzitjz3Tg4ybbGQbqITND30jRSpqfZQxJ
QNtTQHTDgt1OCMYYD6wAHXGTlj3mys5NBSYSaAET7zXv91tezDjDBnV9WQRd5h0FGxW/oWTtfXRK
UThSjJD8S+aSk+tBhwjDmRMPAB7lA95xYzTi3MdAkbq5FZmhURFeEpOvUy32UHsQWp1vr2xv+DDD
PkucQvo/QZXDxQ5gN+y4ycSbrBHxBtuEVDRti3z6ebyNCz6SeSabA4SNkJ44ZyRSasQMaFv/T6JI
uMQTV5hL3HSrvWeEQ9ISr9R3wWaD9PYPc5FvjX2nGjrjo99/TQDgGpI+yh7S4ta53ICX6owltPnd
kX7QG1byKEh6fsI+R/1aTOYJrQoO4PA8p+IaP74twWf9X2aRLEoHTHTj6/NCSvFtfk7fJtH6DAco
UGnKfFFbJy+WQZ22Y4XR+ekcxiO+8JwjYWiCIjpT79Q66ta8k8dHQYgU34T1bR25hH/isxbgXq3m
8XWNPQJHWVSSTNuAOh6vbOOgiZH+cBOlNmpzsGNVSUkdS3EyzK4aXfU+W691lAYLAaFpBhNeU3Jw
Jpd+tb3rW2QvBF+wmMMLM5ljF37aR/UUSpSbtjlCT2yfNUrUI9kvJAs7iaSLPKLti2NA5uxzr8sD
qHs7xUeiH9QofwqgwZTldtb7FVqhc2Ikbw+wP8Vi9499LT1DGzTslkOdDUldci6uFhA6TAWM4Q84
Y/GZ7tPnJMVN88DYBARSx5ue8JZsj3MkBvnbi8qG6Ub6ZnYg7UqDZtlOWUhnRB8QYCkD0Z5vmGj8
CvCmndeUSOEvUp8x3SU69AkBZde3rSKZsJ2S7k2p9U8QZvkRceolEx13QiKPYQdNCLHO0FulVYsY
QI1ALpGYkMm4V4e9eOuKhIACEx3Tqqmgbd9u4HwV10qBDCB7Ujb44ESVmTo2seVZfKOoE4v8pthY
1yPB7V1Za2rhH/TRG0GDV34wAHrtDM/pmpH2n8gQSXz1gyYNmkvD01qALvoOjppcCkjyGrEXVAQD
BD19v3b557ig4/VxxAORtNDNcqhtVAsd2kJd7ljw52m1arYdMba+f3Dyudz6booWnp90v2G6e7Iu
OXKS9pIFRnnd/bIyWfgn6/GZh/gwxelRxjix5hCi12mJWXk37cJHS3GtwW7rqcdRBuXpjl9pfghr
HWN+wp7zARWFzzmjv+sKDXMGlMtLKbGQDmuJXZ/ubWZDBDNQLw6WcFvW3a6kXOVNTFBiFZgsZysb
keUFT9tM4LmSFlqHn4hGt8eBACO2QYnsfpZaDOnk8s6uAKjBqzeKuPWLENtPlzVfa0sNgqTVW4TR
3dMlkweDTY/EqV1mTMF/T5THyKj/m1IVJiAnRxfvAETRmEx+ohmtWVmO1rKeZAGSlQPOoLvaI7bT
Yvv2PKo0DFsGgmPgychRdDpfKAWdughiZ5n48+ZcJOpafGyNz6iy15H0uFBPbdiJ8o/dSl1Cm6qn
w4+gxN9sRxCT6ChzVVy+KL52wwEJBKunkNIzlHPJU4zHIa0c8E0aZnZPjvLtG2TwCOKNFzIVfQC2
W/SYYriPjDihIyvItHyoPa58urHzFTVjKJeTi/pYBFeH6uYVkPgQXIQUrJ0AbbqZlgdspvQUaJ49
GCEqvc80WJVvCXYXU5MZmK7t7/hVl1XKWnTSOIpJKk+/sr2w+UL531wxh/cWLJ5LCb/haFfHr31F
jZRwjJ4WkVOfoyp1WbweWJw1Yr9XdJv7jxUymAUWgl9rQnwMpU8SYwQ4QEW1ui+x8Bif/p3HMEx9
GX0cDaGIBsK/mOVnvXOLzAuqWpjjch8x8MnGnJoB7sz33RFx+PfHMavhcIrGMYonWPFG12d8nRn/
QEpPl+sgPJjEYdsgc+ATAW5sN1NXH1KoI5xk5e1RjmspbruwNJzuFjBWhrB1pHAeUMMjHoh3MhuV
A3AiK6ylSSd1BCpjYvYsaCRwSqV8QRHQDFDSHPw1IP45BvyT0jXZ6W4mjL6VBGssGPImVB4P5XA1
kFv+v+A5oH16sfyAA7caLqI2ZXQFpCT/6DKZh+6qWtHX9G15tXu9xdqw+RtIb+Q2dg+sUU656bm4
MzJHJKNLd7f8777SFCI2yFd0HKy8pDiQ4OIIhhSidVGjReR1zoFS8PTlqHRvsiWeBB8kHNSqU4IQ
MVvi2vDM2tHB1x8PKOpjFTZFf43XcF2kiK3R3bNRG0MfEnM+41fJRU9qx1rfNYbAcEGmjeT3q94x
+juImbOphTvMQ78/ssoozj14Q8tDwJ9n4VkziDQiCVaxEjiOyQa5hVrvXSEfKNl2SE01eQfobqCC
QWOah9G4y3cFMVWXsYt0c1+K1e/jLp/qrArdGe70Jzz7kXD8llL4+Hef2WUUYN+mZsONGgsg29yc
QIBAd8/Dorw4zG6tp44QVxBiKWFj5LUWIF2c2ITrJhs5Z+rLzu3PndlCuFoZodGQG87ARzn7bVyd
AbEv6hYIRJJZnUiKKmEGeejiq+IFsOyfRcnpyBaCFRNpPHgqcn4URoHgOQSiJzC+9rWFv1NlyNjD
93UYqkJqz/Ir3Mkdqt91GtgF14w3mrsEZKu/IIlBvXg+U3lfHCKR42Dx6ykt/U/dSnQSpisPNDax
SML3tButwiBr6dpkfYMsii6MCntvFw/W6mMf5NU285GOvDJP1xUf7JXPHcGUKSXcIkRy0zIWEQUo
d26H2ft5gO1ZIZ4X7JyYS+gjh2Neb4CqHTQDw6RI6QTwsjd5VSJysp3IXIMqRRIEFbY/zLMuQvVT
xataRi8MTU2727H5otXwj3IKHOQN++qfe5EViLWtYnyq8pB5RpxsvQBf/Ax5s9Qrh59vfUCuayzJ
HYGiSYb56PKW9pA+E5d4YwW7cmUjykBc00iQtubZDIQRWSfggOJ4q/wGDIh/Bpmp/00e3zyOUnp4
5ptvv/JBMIo9jPaiL5CVgjUvnwFe/3o8hoP+3K/NX5QAzFF1SCCxKn1HJJSKxjIc1ACBR+Wbu3+t
8q5pn0u9nSu/9FmQoBPTywYtNW7FXTW51c9fX5xdkM/Ug2+8QAtVBhQ1BWM2fCw8lgvJGEQUlaFf
MmGMGsnkgbKofceAFY1Q7VEs3+weA/hfApvkdJ94UxRC10erEbE3253NzXAB4lJmgQ4gDwfiqqk8
nndHYFpJxPBkYQF3d8RV8g7fyIngfBFe9BBnHpdtv8zlyOrsRZAKvMSSGvllNuS1NwyJ77jDSMb+
bwuzTEYnoJAyci4ca768r1zUS2uw9cmq9f/mi6e+7d2MDN/aFg34PVjP17YnKNG6kJGdJ/xnoRSs
fv+RKPUSqv51Zlhtzl4lhnERHKPGdCdTNZtmcA6Egnmz9w0MDKi/LPzaxRPUpntsnqV02uc2kjwm
mVt2NvdEnFaabIaAFpa2HwbUV116buxcZcYpZLBlITI5oOu+n2m+qpgoL0t+j1u0mIO/7R6uoPGn
JUk54FgnlkpiVsIBFBtljSJJZ7CuBzC1w1bQGw9bN2d7yQDQLoir4l95liUwvuxuHKcvmRXqHC/6
IJWOS/9nbX4IzigBHs4PuqLfGa/OKZOtLt/uFCDUbncNeYgZAccP4esv9fuS8OyzJSkQFv2Q9Gbf
t5yDVaZYbBbP2ZowAI+o2VcBF/qZHa+uW65FbGPGNK3OpNrtwcaT/+sbLhTmGp2lqhdEjzOWImx9
pU7nimAoXe79laDz4+Fu/wdIIKIbtV1pamuRy8q3wTJC/UZjqw9kL6+5Rz/+Qw/N9peA5u1S/JvZ
JhTv5AVlbsKhHKhfdZgZFlYU1cAfjN+mspKyLTh6RXgY4TsdHEdjb5k/Jh7UQonjYK04l4p59DY9
K3BIocE6FevkLiMEitWuSO8U2mFP1nxQYvNy4/4zGcSQSOu4cN3lm83VBRjp8zuTnRNIuuilAbR3
hqDARPMm5sAijydTlKk80id+FPMU40pkV9S0gZPljKAnOm/ybg+nSQihiW9cRobdWYlzPknVbFzN
0JuilM0JD9eYmkc+Oq0cTMDIn5Kt69ELheR5PRfdQopx8zZwvS534GBDpebsJNSg0UwJWcZBI0OC
VY7QmiiMRDNyCq1BiZVIm7dXEiI3A8/m0ktVQWohhjenytV22SR+NomVDQnRmN3fjMqsrxQ6+P8R
+wtxEHowBixkXF3x66ovyLIc+zuJ2dcBnIzj+JcXoPmZSMSHnn5Mtb6MIjdmS1DEWiM6ZbEpBrYg
gQeBTU4Oi95SBQ/2En1g4dhWB8nnGsw3SYSMSFybP+1z2wsPRL45u3Y6Gx5vx/O3rgO6QA3xRJVZ
NKkV04lQF2zCPtR6o7KC+NPusHPumezecvRdxpziNDfXPugNJeZZ95FKnFmkWv6mqi3cYOukcLhX
VT7Z1LNp81zG8d0bOTDJPW9JRG+0VAYSr/VoX4MjhXFjATJwPG/NRub1Pzc0UAELVkV1jY7ZbuBg
AXBG3GEVZyN7MYAqXLG3yziOLQAaVN0BJoBwBqezSvMfe3chXhQ7kNbt5qG8L1tUFvXbLCQsMFGT
L4f/yK2XipzLNF5UpBOhKP1d7dwu0aL+msnek/0mxcvGq+sx20y13Pm+wF7qxbG6Mgoe0DIg8IuE
lkOHsuVY+fMLLc8DSabVY6f4ppBMAIzbtjIKhmd9C1rvNsUN7vUHidaJwNmdCfARhB4NrO4JPAQs
GiHstMLZRdEn7P/ursCvKiQJBSDFGXTEnZcqtGq15tzYVyOwrlPxOcfVawdKbQGe1p0iZx4ZFL7T
FgYI+BrlQIIHHXHfKWVck61xp458/J8JJ/Dol5FZmkDCK6RbNzrvcpY0ICuRRhYpIgJ7pGWk95i+
jqkTITO2WTXjORXKBzEyF2sc6XxT9x6+ZIwI9ai7E9Vm8YzbtZAOcviNE8h4dmBAwsPUdtZXTg90
Eo/nOiN6ytFP4O1ncqsqCpve86IAGpt1fYRV//vgl47lA6/DZWFfXMsLGX5oEBncv/bjXgVmMPd6
uyK7qsa+CBLXrw+Zx8DvgNEuGuZcIqA09L+I+spM8kJAQ8oA4AX7dklWefnUUCpq0kro++TE1VMI
Y29Q6jMApbhbugrJW3UsUIxjH5aThndlwQB7cXLE5nGjSN8TarXHQAKRtmII6wyb9nAG5kDzu2Eh
LBJNEP9bghsqLMcPpI4WVv1uZSguRtbuL12T9IzMgXm9BwgLW3ZWKlfB0H8Kva2RaS/X00/TWSGS
Nc6OD9RYYfDMYgofv7pRtVT3xWCuPkRWZQC+fCzJVHw2lr9rTgg/Q9PyY9Pnc6YzQsa/5/0QByYG
EI5KPomzgxPc8bQKPC/yUPnE9Z6z40FpYGX1pXL4UV3woN8T1vjcs6tRFl9GSNtYNmvK7qCi7d9y
5FnrDdCdjEn2fJvi/jwsv5eNIBUhupbPUJZSBqGSy6HLU5XTyrp8uTI5GpD5LYMAlvfT7Koi7Po1
xEL3PdkyFLUVyWubIHVY4bEPHivBoiki/DLAQ7wLI+0/hPmAgpj9AE8gTYV6T2vfSwnjfJo/dnuE
BTDlM/Uv6JIJIyZKoD8J7212UQOZ9K/00rmBk+qkPdtsSqMWTXRGrwbSGCmRFIEuzuJH4TlcI7E1
4+DMr+0v/Wc6snXtUUz3yaynaUy9ZFNx8vxTxkHK+QLZYUXmGAX7cLyhcxTkGq5Rv0UHhqbW9gDg
oWcyQ+GvEHbmtaaI5gf0nXGrr+I0XRyxnEkzCGqa8eIm/AF9BbFVbmknKCeBSHtxYaqncBOaA+8c
erZR0BOjRA7LGew3zel7Odvj2wu7hD8Dq9l3rVZFWAP9I6IEWO2onpg/2ePd3FghB3iA6eJeJOcc
BA3yywM9qn5swMHDV2G6f0Ctao0DNB31mPjSUCCBGl4bHsSm5jH9xvEvW08ffX+PCwY/Mq0YY//9
uYz+i+z/Z75eASAQnTqVwRFFpXyQlc8MihuVxSa34UW7vxuMrpLEvQnE+YkGzT7WCYhpophGIe88
v5/+lsuoTk9Y+WTqLTbA+kBWjSmVgvzQlLrDweLJW0OT0j27ulzK3tgP1RFp+pKdlLDw7vHPD/cm
Uxw3d7gy+rNqYZVx/3zkuulZpaFpJ306TChouc0n5VFZtrAhufTpJF09X8agvlOr1OgpppAjiIWW
66Jn1tbNDNzvf0GI97yFHM8K15IVyuTaxr+ZLr6+Ctohj8neuFOaqRPGtZiV5eXAkHoYekEz611r
rfwmHxgi6YTBMLKldYozVcHKKUbqhbBITz00i9Q1aG968N+QVzHCzextYN9tP002nY/0nYCkb1BP
Mv7MAFvlhOkACg5nKttQ+vQbeOVTXDvKtam3mWVnhFoVJbu9k2ANL61SxUWB3V72xM4X4SYaFp1w
MLAlyqQBmk2+NoZs63ELKsibD0zJs4JREc92VjkfEkGAtxeEPWPwpKuFp3LXZ/5mZQvSKuk7d6ty
koBM7qGsdWxDKqiVRSZVhzq7OORDzRIguK2j6G3LCJVrg92UPA1GhzUS7sIGuI2aBK+AEA1Jdrfp
EKKrU8cpeObEfkTqL8NWF2ph5B/fg56eJzPhmIZCnELYITeCQqkp9DKg7tnbPnpR7Y6UGO8YXg6a
EdoN7FNYccaJPxH0H/6qr2wG+Fwyai33nxhQ7d5Y/7yi9FJXbTZtljWxHQw5BVYE6/bm9Bm+3H88
Q6sTbPGBqRiwAPyRssfq2szrxu50ofQCbxbxgLGgyZEUlEjULNe8dHV3J+C4+4+RG/JXMeONYGUS
0sb7ndIfMGd8R+AumC0ZgYRtCpJhxSrZ
`protect end_protected
