--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
g0Ja0IpdyxBqC3mY/zHi6frbPANuBquGuY4UxtjU1+GOXjFodxKUo/VWDB/ynFdLT3JpW/uwCjF4
x5TcLNgZ3pi9ex+mbrCshjnm+V7WIFDc5g/Af/dlP1onmvpgzVPUaMlbNbN4k8OBgBqGZC3a6Rhb
065em/O6A1BniZo3md4a+3xqfWtEC2BM8zj4pc//NVc+70QtCxykvL3cJfI1JDwd2bbMi8Jq3pru
qRJfi6g0cotoSasvvcyKw7CYFz/qUeMVqQbL5ZSPQdywUftG7cLR/NSO+C7tcR7cOIH/AP/fxvnG
jbtpV+kdZcD0npgVMCqRm5UQFKBvFL06sBLnBw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="bijXQn3eJZ3kmSgUEz5cfoDDkFu5Cmk8o6Q/xpf98Hc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
BACdrWlG6HKrB9fB4Rlzsus5UpSRQvUov1Lfr/J0ENiLTpuuBJCcqsr3T6NCTsmMeBru6hNdBt8s
Qrf33WRouxMz0S6RJ24tj1IuGXxTUv+pu+1AOyDmh64bwPRhDWBljjWyXzaI+PW4MAI1cydqXNmV
ZlWRSHF+vJKy9o7iXKl87wOH0q+sZeRZwNUOhc6iQzqGnRiL9lntfD/ZTnROM4tVVq5s9ytLu7+N
kqqZ6N/evoiHwi+ASfA2/OeW+xBgqLnDuCjkPkdyAuuPQtpB3YpHdBzJaeyKatpVYY2bzB3nlcC/
ziWeFiX70hlKLxQfL0KGita9qhf4J5Qc4VbuwA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="EA/DJlINcHOw5/FQM19mujrLO6Mlz4bmgTJZdfJA77w="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12336)
`protect data_block
2lfp5SUlqkNF3fcI1frKdH2SX4iWRs+6my3NwLFgMhMZz7j8ICqTFDlgRew/QLnUWs34HHI/SJO3
HQld5P2dUtEiuC4Z31bGK3ag6R/TlAj1a7iBlL6EsA7fNljh42PXm5Jq9tQ0kfjFGDYtRbRe2i5i
/gwRD7Z0j/pVmClp8R1EHn3MQb1kPTpowCBurQ6Ssg/6bxkAaA9ykBI8NQZDXyUNDoGieba42vya
/zGwSNFRZ3nmfnWF1foKfmnSJGLPFf39rs1N+j7i/0wBbZjygpxvJsGsXQDYa3dT+liAq35+E9Ll
/qXYfWicp1+hF+/JexrOs9gLCkyk1agNZdc3SQTJAZYdKoNavhq7FitenMUeCGyFrYyh3Xsr3XfB
OCA6u7xCgrg5ubO0L1UUcPx42c1DpXecdpXc+hq3tF8EjG6sO5lmcqcXPpbb+O5W2PRxrIc3OEDe
dAEaH4lj1J8DJO5Mqvp200RbA0QiTXxiVHL2cfUoRtXrIpbj38VDzwiD94JTtEJ3vxG/hACvjnm9
ztkNpfLSLj7PiEN2T/OSf5331e0DWcuiLDCeMHDpQAyJS7scXJObNUYrkMvB9Ac31M05KfScAdav
cxb/S0zfhJ1sfH9XYgjhJaPhZwJHvOBMqK+0rHECZTiMpCdZPoNY5ndTDSYPFcpNKaHvi/0KVW8I
59WJL7NgCq41VHTjl0hv1YstqF6lwevXSDg2zbW8MYQsHsMqlb1g9+1baJOsUGQwvKgatuVNs5kI
4s86zybO+2hWcI+na81w5OFfDk0yd8OodZdMSKLmBW/Z3C3Hezxab4V3QmMCLvN2ed9YOuAGZtfm
qQn6gHtpPVo3A+Drfi/NflcBzHFdoitKWHbPZmiRFr0uL0I4huErvHyIJe0+6fOyRehhEsXkgTh0
zy+vRVv2BdM/qvWGgf+EwAJTuvIR35c4Vm+q2Kir6zHqmExUN5yxa4/x07K2BBR7AeahSUF0Q7y4
o4CHpTu8K4L3WW+HmVSEFwjpJZrFsZkg6JrYNIyCKG0M7UN2Hi9MFXFFOlkJ7f5p1mMvnVeXwO4A
Qj1jR3kcpgpyEofpQIMncpvgqJwgjQW7Qjsx0cczZK5XDCVLEsJqbOBnIDdjQofeGhQJ1XhFdT4g
l8aZPdxyY7swjM/S9xKw5Ye135xUaupxVEym9ZG9zjDRNoBOExWA/n3adH7el3awJnREsjsY+2a8
gV6cbI6G9MsZ9+TBeN+Uln1zSOm3rL8FOqypZAap3TfFqePt1hVKMedSosGvUM686qfmF+5PWgzk
vBvHHnZ6zqoFJol1b903zSC4axwOTr5hIjDPdPZQlJSMQ2Xn+gadL+gon83sZM9ZJvk+Y9H2Wqsy
1eW9cumUxiG351glTpbWJKdhVn5ED3EkZ3emSyLxJG4QgNPPI4aaBn/7P3U8VRkf1+N8Ej+8DqUh
hHCJGB2uezWYFgT9p8OYyicPpwpbO91n1qZJH3FXIKCs8DkbyiE2RKBubZAvEeYOoVByDcG1aJGL
9+zEWo+qjUqJN7ruE3tELzy0X6maRms/SA4wBvCdPRkagZM/DdribPZlIr7q6HLNEusXYIFLddax
I3VZ8ekacWubCV+Ew8VE4cuJwGF9tpNK9c2BXsofAvGVeFeUUVezLgB+g8Vu8DzKq1nXdgR9iGoF
sHhZblf/ho1AH4RJhLwIXC2qDcyP0Q/FWiQx8BsGbmeQyxlEWSPWONOuPRXJxUo0W+HEIlvOFIzG
Oh/9AC+VEAwj6RcoRDYNZmapdgJG8bqAPBI/Fvd8Fg1JM/LW9fwsjpGgMEn6NdcWFaPJdlPDwDCn
xUQY85oHSpgDSQl0oIBK5Kbixir0vqJd8sDpnqmevRFL5xML/M+j9m7GnnI5xSFxy2d5KUA4fAM/
hS3WFr/KBZYI8sPvfExfhOC/H8tGxbSKfX9yWjpRPdJQqbm0SUn6qaHxGHMjNxQnVB47YR2tJRMw
rfwWDLb8tLu/DJGaMy4AOiE8p0gSFPR7AeVCY7xRLix+l1V8YYBOXyXApZ9YJE3QJyPtU3c8D3/c
NC8CgjeUWFxz7yhJCR4BuqLFpFElrCrzvTrMoPznJlTpQenWh56l0a/h8geAakxgIeitOO2oOcWj
FTdJvvstpqqpKsmd3eH+GHaWwG564IM4MxqvNwniQAPyP6GY2t687tR24N5N/Kd9Thp6WX3kxUF/
pyYM/RFsZxwV1oAGVpr45u7jRuaAesBalY6B+3YeZZtABSdw30HTT1808EzlVQcXo7L/p0QCOzoE
4MzPIFcy0Gqjldh76b4iGXwVGStMrFE0p4iO6HWzaadFEvrBNRuAfeB3cmU/UpDHmhxbFoK9xjAo
Wog+NPZ90Q8aH8iwvnNZnqgsHdJYjsUX+bvP0KVNvOTYoLWml53dVc5NHXNDgAHq8JG+hvWsa1N7
77cPJyTVVKRgGiyg/Pv8PWK9KCJkGEGS4/HHEuCLDNhqfvYiwuntJ7liuxsydjwQ+FL+Md6RMiXz
KlGiVY25lPETrw5KQxvMqXovzWU6v17xvIQ7AegtaO8pciL6bTLrwIEboN47+9j+gaj5cvZ+wnnl
/xFb6UN4IYEIoFza28+zB9uVWwmIg5bHaV+IEixNHbiiOGRE3/bxuK1sndNLKfiXZ41jL8XLebwB
FAgSJ6rZzF8rY9/vSXWvBUBNSjG2ZGWE40VvZ04Yn2q41BqzuOns+0/kRIXnLWHsuirGXFHQvCIS
oFPOn4/XBHfG5jwUvHY3P1M9OORFUxsij4ovqiNMzuNMm8xdWiq3GWkvDjLdnYV3D0EikerA29SM
q7FtgetjDWy52v8fD6nWJSL4oKyuB6fACjmf2ncNZxC8/zlfXAY9m8rVgJLGCvr5D0KZ3CC1LKwk
YxqZzCiw6M0Kw8yimHT5EeG0rL74SMEdz7xWDUkD1fYYKCZRWJDHAWBfPvrWarBXpMaHMfJvurKC
fHLF+1ndNZ7c0DXDpW+41bedMQWadz40hZEJpbLXq3xbuk8nBD+G7czM/767vMEZHxRycxR8PvLy
VFDshD4FocsM9omffzvIoEafDkTXLTrOHcwsTXDLRZ3Q2lBV1uHAjRXgoR25UxnrfdAh7X6jEpS8
Tu1D4otjcIKzhIdX9/9FDPPimQdc8wkz2m1RdQG0MRAqzal8nPMVp9GuxaDu37TyhvY3Yo3wvsMV
22vyN2dEwano+9Uq7q6CSfhxwv0Ft1THZvaCbBkeCQ1UeVLdXedhWwoG+vzcrcKjGALqpDhuqz8+
+FiEN69Jc429cNL06PN/OrTOPn4Rs6zu1b6KdPKW0xCtSb0KaVTahukyMAyorpo0c0zqjwOBZwVx
dqA5Klft+Nd10BW3lZvS4SmgqydeY4RWxraN3M737wV2sqF2174rAeyEtJhYYu7WeRO4GR2No6xy
2wmXTwOIC1CuHKlw790r6UsvemY1z+Y1RZC6eXEguY7b7ifVxUV1xIkIkJiHAbqiLPyizjtDTUMq
uMonFfa+OhDFyPXC3qnZl/ogx+1CHCkcYxVvzyl4FQ4fLqgx3xQ/Y+l1GT6Ufe2IrQKthhNclSnL
wb3ehVP1w4Yv0qB0qWuKlQ9hj2JKUlYHyEJoHtOhZKcCX7pzy5NL9RYKqHtKmcHGdZMWgJV8054F
/nFjaS/n1oHjRR7m5VNwS1tMA1OjR6vOn60iJCoQbcfKrppXfzFU8P+UiXTC/qOkgP1L31rJB2+D
UmglCF8LS1qiY70mSP0B/V+gXnzgi3hEhXzWj94ZI89UY+BJmusGc2YPmGH+IRbU9OIV8r3gfsos
UPIlRwOepEUGqI82+vuyPTaEahYePmWcZx8I/uwNTJJGGiRUppDDHnb7d7GOdjxitmlXXPnOoNss
1fSWd5cIquJWL9nzwZ/ZP7fc4Kwz3t2oI3kFin6IWR3gCLzlVqplW9uoqzxpPV/B27R+pG6x6lUe
zmxysqBTDvguOAUrvPC1zmCpmt88xMjwgycr70BG7jHM78UKyt8oJcUXIGsiE4XiJTxMLnYN3xJs
eGBPRR/NBRtNOdveFgDZUB2zI3+595QbbVyc2ghL7CKyytbP71GBfvQN4VGzxKiy7bnvhrl/gu8X
PvsCeF5+wShP25uRF+crkTokHFFJL7QFSsxwB+uKrgDBhYRZXKcs3nxI36eseX8F3MGgnSwZxtZ0
HKDFj17NtsHBgd//1Z5MWYiLyqworLxO3JaImBrOwbtoCV3VnC1km0Tt/SWdW+GF6Kku3hBlrYsL
1YZrHp/rhjfqMGhT6F6Usgp/a7gSRP5/8weVxRryfKA9KHVM5dmIBKFaiuhZXaIi3Bum+Q1ZGlzS
op+f9nh6lBmfZ4a0SD9/w0TJ0ZBVEgi5DMRHNW/c2tgsYaUgpI6RD5AwqC0VxhXrXR5U8+5MhMvq
z9sHgEzb17WUkBPGkk8kO3boIpok8FD/oMLKxcY+L+rz4KU1Y8GOVqTMtLo8KZHXCwKSdM1C0Ama
+ba7n8gVO9hmqqkKpsmvCGnPjM4sP6TZjWnlg85QWumwqOyxuPH+uvP2TG2ZqTpblOnhujr9EYtG
teFZbMML+RwU14B0XrFACP6EGcQx8Q4Pkybl4oqNGbnk77Q/NqqgMcD2yhCc+wS3yyZ6EfLbqmGX
P9qrfwx9RuLmwVqExBNdR90SGdPFWVL8rPi/vdmJEaQ7g7YymAkTcGOd0RPBgraLsuw6Nc7u5NpK
ffTWwMfkdEys8uIZR4eCLH7s2IyF9j8B8JoeqUYeaevvCUGWIBuMe7+mL38yGRgboo2nYP5XYRuI
iHMvt2kpKiT1y4U/XP9Vaj4PoFiCRSPgFn8xAs/rwqmVcWMJll4xILDhzk5MtK7hnLG7N6rTPxvw
2WUoqUC8/yh9lnkXBvL4nM0C5nXL3BlGm1Yb6bhnMhzSfqfmZTJkxDmVapuDp9PwUYQ5RQfXHb8T
q2C54E5Ek4Pe537t+KaSEDZrpLd0mq0/nPE1uWldEoTx+Rzd9jvfjwG7shawixQf1wZJBygILQvv
SDzf5Vnjpj9w3EupiWjdyNJN/7F05Tm/9Wam7F6zryUdi6ioTWsgQLdDMxpn6RyNyMZQIpEA5dDO
rZmhEJmt203NYVLugrTABHPvdphycy2dFv8ENRn1I6ZCMnIh2LIW+p2wPzVmjB2sMznM2+0PlmG8
3nnWyHRdIeBR38BV15JcZJQDOQf43Tf9LvUM63AjUzBajqc79UFzFMwB1iC22xXQkD7gDrGLL9al
YIuYTocF7zdsIqYS8yBYoyu7m/+gYo19q7bEOfJnuSuC38HfzrAd4WRPEtNBoM+oNbfKMZ1Z+KiA
wZWqIyW8cxkZj4WgP7XeqOHFQUm/zlmwv5CLHCkjKUUrCAiF5qu/a7/IXST63lb0PqT+8j1dPKai
UeRnplww2Q4atwnXPoPJKGQSvORGZyL1wBLBERDb8gl3+JbV3I5+fYUj2UbRaHf5SOr00WFgs3+F
bO6IbuUfjrU3lEjyJUDhggdWi90gkJUb3kx0yJAGsyl8SjaQZBn4Pk9q8SEuEKKCbZ0RqXixbWtv
J1kcKQPeYeyTluVFyW4kRyI0lAhLBQ5ad56LL8LqZjuP/Oa0vTEIZRdC+PQ7Kn8JErynDS5YWNIe
tmBFIhzSxfGIZPGtplt7w6nhiNNlNN2HUzyCeZFP8+EfJT9g/75yBs+bHgmRdWtqPuWWk6Ph5sTg
kUctVAyf83n7gmcDwoQCm3s3SBGnYOtKwfiaC60bw++IkD5PTIccEJGSIqamVxM/06daTms3MS9R
wEbyjNBzvU88TUM+z9MItHzbjxVOYgMjkvR4LAkwHQPPUXOVf1enOeiFvFM9SKv00NOr5+2yyuee
K436ChjA8rWnGn8xOkc8kGPgwcxdLiFCESVtVp8ujx3DMxyMHjUxKtCsGDrLCupGGcF6XxkUNovS
6TcZOqKBOnstHnS7EdcCejdJbXjgmIs8xadKdIIV+MKbTwjMfwboAphXodumHU+qTmLsoYaLgsoi
GBEgZPN1mFg5N3y4EhCgRD/dPsuRUH0oKWm341ymsLKvh1ddQhfgJAZTAqtXZlEpg/q15dDq2BCW
RuIMHVSPFl18WQgmPZ7uI8BTEBIN9MPddgt5Z2Y5RG1ucKHvVS1GFSVMeulAwgNiJo62BcSiMt1N
rrAQh0oWhenDFjHBO/MVxN6Tams9gPmWYj2mM3AKsicQheEkBMeXUlzq2828vpkWFMHGc6cnBPaF
/lSfXJYX9CIIT2lEl1yNv083DopuaQ5eunL56zBOKuD3CPyJJjnSdb4h4UcGh/wedatzeIOd1dZT
2U8KlBw0fnfrWsBSw6ADEZVObsezrYvvr0pJBV50VTNpWHU2ScHNflc9OgsLzzjGvrWAw24WUT/0
qdBH340VpddgS76AHjrHUB5wLuU/MgXVsq4xR8E2YMEgMQhiro0SzRqn4uSV4KfA5cvNGszSWobM
jnWFGihzJ+J5/adGOakMhUJB9LBqWm3atM8Qc8bNbtXNu2A4EdzWqvtokHwrJsZlAjnyn1wBYZZT
oE2s1X6up167xmyDdO6uZk/Eg4keghkBAbl8Ew2Gwne1judqBmZLEmLbD4jR4GS3zgj0StDRO8d+
8FBQSCWnnnkWgtTUC2tSUrY3BzBlF/qi5YylEoRVgNAiTRuxCTh4NG6K0v5qN6sgjRaQmR3KC5cv
P/glwHG+EgEZKPBYsoSfZ1CFDqvi7Mpqx/yypGBuQ4M/YKpp776qes76OFVOQLAPMIDb4DqbK8RL
8KxTH2MH9sh/D3jYpD12i87xc3A6qpU7cwsOp0HBBZJKcGS6D3NVA6UZpgJ5+W0+sLDSPSami1Af
XnuaPDVBeyme5s6MtlR5o3HAJ1LzvxIFa38XhrdXd2K35jbT4Xb2788TQ14th/adRhzHcGT74jbg
oC3YJ22Ya/2arPlsDQJloiFli2kFNd2pX/eGG/MUrbYE9uHRtXN51i8zTxPCPLUTisqCbXzYGjA1
M0z+IMmEehdT61jPJwt6ocGC5NAvtmuivsvuv0GyiNpt/JuUBjk2LEEaxIsmNLJaVd7TIxfBwSoe
qm2+NZQ8dIG63Y2TzlkoUajE0T5Q0NhVW1oRBYZCMfZTHtkQV7QTWJcnz/ZK6LYbcJ6ah3QLut0n
bQK3bSnMJ/pFw/1jU/S5NyG0wgA6S/hBvB+0ZO0HMg0k2LLedB6MAK/J0+URS4RJyJ/gODSru9eR
Z6ez9/DU1n1xh5ztfoHfQ4MlC4Ap54pTmvMV1KgpAqoRtThZrIl65fzF68VzNLjZh2hNxPUemusj
lLthitZSbWJzkPFSVU4956iQl55yP5PIYo1dipXlnAdOBYVBDbPwf/ZNy00c9IfR+02OkYyA0c+z
ZKk5EU4DxAZ3QnZoKsjdQz8zSmy0Ksgb7hMhV68rTw3jLEuahsxdGFhzS8tdbqcmfHhykbRVqUan
HBj7GdU+yPkSx6kJMPZR8RhEW8YZjgUq/Tr0W4cR2NvZEF3RhdYFZ/gxtBClDvSs5rlqTq0tEWwX
lwB6XpoAZBcSWfBJSz9aT1p2CZimf+ExSeL7uxbC0wntH8SchBTsBpc34B0uYkYql1hSqqZF7N5y
e0yMx1yDqkmsXJ665AMfKwiNsRMjG7KgseGQr0wR+mJxyZd/19Y8878rMvWEDBe5ghvMPrXHJJlC
mW3S5YZ8v0x8N685XLyiPWWkxqveWnNijrTf2yedij1cEyQ0ENWtdVmZsRTkRoR8ikVx9f87p+Tg
CGhnoTKaT83ckibDfO5LeQHz2N0ZTE+TdZIRIvND3VZFSYqbN66JW5LPoBUf0t5EQLBHbHmntRb8
lXODYDpTFPhwHfzvQoCJrmOsDfJEPwoip1Mq/NRZdAWl+x6uQVui7FRoJa9i2fV5EiNk1EATmhD5
YXQ97NRj0FXDtYB6SJ+BLKUCvUMNVEkDZTydCLrRdDezAz5h/vFY6MqZBBFiRKR2L9TIJEJS7/LN
MioK1L9dxp1ykiNXNRMr/F1cpCfdyOn4V0FWlv6KE/CJWMcgvyX+SVmKapA2LPS48PEPq22F8G+f
i+Ao2j71AvOQnMXU3K9sL+WgPlaHCO4DHU27YMYLBpr3EqWQdzZ2SWCGMNHfdSinOLyuBLrV+iEv
+Pqre7d6iIPoS1yLQjv/3TB7iA2/KWu79A3G/Yhjdf04uOI2KmMc/Wo75ZaPg0IIqYWIMpu2G2fs
pfDfrHAFXvzcvXxmz1wSfBxcwE5hydCcyfVVTZjFpnqoN7Ay+3EHbW3x/0UgsKZ5bta/1NE6UWNP
HWH11tKvqGtbk0qN5JDDcsXqf52SM7LfTODBtu9MJ/v4/g/sY9dQ1E/yNMN7Dy0u2Dzj5j9ZM0fe
RN04fhxNT528tr+iCeBR6txDeU/dHZlsgn81Z2PfcCgJXgB6BBGPVpBuT6JTl3cKhjbEWmwLjHE4
sXGTMYJEqUQ4o3NBtYUMlKy2INYGjnSNJCMdQWD7tbxAstlhIX8PL8fKLvVp12DURa4Ekx/NFeq2
T2vzApea3wiRJX6x8ZW2w4ar4mK0OmJgsiWoaRpptf1XFrwUMlta4bCewmRPLNV4ZXBVI+djf55u
C1hi3C1B9jKFMT8KnliOlWfx86VnIpBI1RjHKCDsYT2fUHi1aVjmbl9PzGjN7m5ZFyri9GRPpgf9
e6pnVKiz8w9kfb5nK5A1CkcxkV3fFLl3DGkapHwpf9U0XoOS139uK2BlDXb+oc7V13BbT9sNzYD5
XiOxpHkZIVIeZdqBmTm6rgo3cRVg/xjZgIzP8MK96ZMxLKU0wV2hZD4g0ZJfndOs2RjoRZHrgURK
IMJGCzLrikopzH689DHOrqW0hrpyqIBF0I0VZsM2r3bSQ7D5tHhMK++12JdaRczstsjOXfTe8KsD
iJD6CoNiWz1TXA+oVaSedtH125X1tZFyqb8kJ1YbGPGtWpOm8M1sKf+AvOGElt5/6ZnvmeCtsFLY
TeKx6lHhOPRvVxnfS/aFsHEFxL2ekFijmc7gOMmENPS57WQUDw69D0oy2qECcJu2+dIDkOpsQ0yc
v9gevwKpSZrO7SntP9GpO/g8t8e33FCOL3TvDYzWT+v1/izI7gmJzNVlS3vwhgVRm/GHU91C24Rf
kQTH7agJ6g31jB1Fh/URkkLBvP6brnCXU670F1uqROo0eH1+v4SqlZBjU5RouWRQMn7M3gdLnOHw
IN2JKSoX/BISrCAwHPQIzr5ZDYasxFTYH5MIrDIbAPJCaeyAHN5jp3tU1oDQgh74MI3GCKrUfaVa
QONH5RNORxt2sJ+waU+/53pjxhFEDE4ZyydnZJQdTDHHSFFChf1WucXn7dYOF02xxMvsCQmtSRR1
Dj2BvCLighl/mSSd7R1ctVHTC5gZ03rlncLZEL+fiBvVtsbzoQwplfsdWrBU4/YpnBOjXjUZ5arz
9SdGShLLTJgY/zH+2B+HGeoGVH2FQpXP1tabh+T0+uhy6jmBFa/lzZnCD/oHiIPmG5ejWE3GMfDr
LsZNSLaTRMkVhcYKw8rmb21NFsAu+/id1xZSJvv2l9/k/vyUmI55zF7pqoCgTD3z2SNBq9QJeD+d
QMuxm5fyl2zHB+SlESEfqbeDmHmStLe5PluDFFzAQlPrBjOPslrwQTdvLZtEOWAZEV6v7qaTw5RB
6q5i+X+b4ogtKROMALX8I03GZcn5VjXNP9vjk5JXaUNpYYIOAH5UlHepjHLJ4i9BeB7CputEr2RF
6/GsblMp9k/0yNNtvppq8UMUtXw/4zmSMsxa8F7leOpI7ZlRWdqTs8m7CBoaiGFEJpbHppKj5lMZ
Mofd1Ykr0EmZFOtfvSP3jMevLVe/peFUs1qarm13HR0enCMXxHHOiPOsYTFZwQirC4DAtEvYmQ7l
f7v/khcnTdaZFVAhgbR5gF2Uxw4SyeD+mfm03LG15Z1QSrE2ZVQ7ZPkOJXK7EZQvbVG0jxLfNCa7
xVN/dK77RIoJw8E01U+fmpMRFsrEwZCNSjIAVNik+e7/DER6Fh6jd/EcvDSq2gKxrKHtMkyNR2E+
/hP2E0830jfNROMrIfl3qY2yU7nJ0+cJJkPev0TenYHjVPs4MoMXXhjIHRvvgX0wuMNU1StPZ5oS
QkqVWvae6qKhSAVFrUlwoY0GI2EoeKXUJKnkHWwxkyAgtG90FSHrF9KnNA5OIu7nyObTNFpz2J6F
FHnZcg+Dzk/cP/Yd2N/NxJl+suvGk35mI20/lsdn5dAWfIspOYR62OVvua81TCJkKv4C5nlr7R4h
eN53mJ9+gnx7oGYo+Z6eHpDLv0C6kJZBabhkFHXq+2Iz36S8vshfTGDKa0U4M5EukTpBuJsJwjrO
eggMxk2JIfdE6Yy/btRCChCRO7z7snJLwFO2OPwz1UBUqC2tlPRPTwXtKNL/j3lb+VCjrREi7QYC
t66Qx7lx1RUp1FiDZe4cMS1dBQEEBsVq827CmBib08B6B/fQ36O9LexyERQnXOjirmf7VuXmhsWC
0mntCZvyWaDALFtapn/wGKdAhARtRA+Ob71EMrIqi2MjTuqRo6vCJlKQuAUEH3/az3Y4k7dEXYGy
pJirpau4BkBt+8dN7hiaAOEU78ZbLxikqGrCrJhN6e8DEoYdGDPioP2jEs+uW57b7QdMo7JUzvhP
8F7b4/spgz7GZLOmO3k2jzvE2j4r2JV7tcD7aP4h03jSGFIxUvCHjyVSP9I5M9KgYeoSjqP+wjI/
2khSZnJqXHF27ou+YmCvvPzO8TOgMBBQhNn4Y9Fxt2pcjySNvTE804GsjPsICUkefZBQEK3TaCj1
niFRseqRxC8uLoA+reZLSf8Af+PAoioXR96w2bfyx63xPVSB9BRTjKbNu8rFol8d4aTLxcR5Ehiv
C7nnP+lCiL0bcoXDHBwUcpZ5XOWlJPfXvwKnMkbMvWKdDed1pcdg3VWgRwFyicocIjg0saDxsytL
7dBSYUOq7HrhQRugKN13HWIJBzGqpZc7/pC6Rwv4eS0kKESVjDsZEFF3rTd7PUNu5v91fvGJcxwW
csXPwRIvFHz7qzWyaHxj/HF4AEMiQqit6s46jxlGQk6+3g6Xk2Czh5CbapyQgXeXWri9Hb76kpac
QOpE0wi1BDaBdsAR3e4q3RuhrD9NjytrnDba4mBCjcmgCtQB0Kon/CtfnZ+sC/uNRIoT9M38CLkL
I20owDY2/8NSASaaQO1R058a8LghskAjsBvfkaoFywUawos9KGyjr6K9+S4keHXuAPjN0BoIX4UE
xJV7fmR5WidwQqss++gyFZJFK3Yw+UxaaP0DQgG4biSpkQEqSLQTmM8rZr9nqc+rYXEYf22ZF7hz
NyYe1uHul2wQ2vFnZ+GPm6rirzD5t1cgo01SSK0r4U0TGMSaPk6g7D7k+vnOwfjDzkF39yNSaGEA
JHSifsvx3qcq/zhTdYZMO6jaMgT84O9iPTYqck3HM6Rk5xyKoZXV4sT3bgE2hyuagfNabIsx4XoX
dxqh5cnxVbuzsAquttryrXp+Hyj3x6l3w0W2ucMoiPmMhEebKxjLbj8BhxkMSannkkVSqGvpla+Y
XyhAcqKEMXv/MNU9aHQov9ZcN2KOR5b4B4S8Cvho3DB/en5rbEQJBvsB/PIjNGRLz1womdKMLj5A
j6cIwwgFLTdgYhUissYDmTiJ3sEJVmZP3QYHKetetZglckG3VxdnLwF6DNYvJl1del2vS55Om9WO
isZUG+CKDvp6kofasfzHz9MyzbRkkOfm+rcrlpZFFIALeeIuBO/76+vGpuxNIqq0DMHoeNm42XbH
CY8dtHrxhBq4m8u7gA3BYrIxMzdUAGpfu9c6w0BV1Y823ZOkLHQ8/tUxrKeqOzla7TdoSZF4Y863
W9DQCgiZsEc9XNCSPHKdY16kWsLYp6sJC2JAh1MdUNAi65JBC0gTG5Knm/0fiovrOdjWTqIou437
OjcYb3daG417oUxYoxwzMuXhPogO+knuW7YsIJTwB/W1HMWnsNuUyCjdM9rLRrGyc4Tw5xqTIOje
KiE7b29xIx51ZqyC3mPg3UYZljhTFBNlG6dfCgFtwRM9+WWeQZUwzockG7zzKlu3AuwX7dZxIN/n
JkUTnBUOu2+qONcg4hmR3bgSM8l/Fut7lJd8LcIdUMpEf8tTJx2kQTTT+D/j5PLnJN5hTfwrtwUK
Ze9ybSdFacvVdK/JkCKwNgqedl64A/UAxmuXAhhs/1MIJH7xeT9Wv27AHRFtVqOPqaR//6QWzcOK
juLadsHAI4hJfJo1ECYB+uMOGtcoG0U6pHvQ2dB3KZ27Ijs7DLS7/Xs4oMtQEj0lIWVFOeIfS6GN
ut9wPr0X4hZYjuraGTqXs6TalxTLboMkeH7CIPD/WYCYQmyW0OgZlZQdVequWOp6lVk2VrPLGK17
cYuFTnBYqO6YUsKHiFJcPBY0qKQJ7ptvnqNVF+Ud1ekHi+z0iTMN97wn8Fpin0sZC7tHn1qYWg8e
/fHwSZ8wqeLPz+iLFTJX/pm6zEkZgaLkGaHOvxXwoORQb6RRi/szLpJ1Yjd35hi7I3Y9kyhEWzjt
KLrfAYtMgG9v1/sJRrSwPU4Lehlqi3PR48CjxcaehLjhNUZ8YTHFLwz0P3I/fQhwRptHdMROYC1+
un7awXiUBCeiZgXr78ApTCaQ7C+dXHhf2Sx01irUjL5ub+jV4BqpPXoDe930PMp1It9C5ybKQrN7
DYq4Gof95mfOZJyprlDZkP07QUg45wgu4EigwZNr4DdS6uZIaEBWi0qYKN+xkAcQjQqtBSIZTa/h
UyQyaogZB3IoTMDITSeF9oI/h2QX8jCtt86Px8LdYfPH6iEAnwctfsWeNcHyxFIL50IQg1fIkRcx
1Qbb5Bpn2uaOyXkka44QTEGojbzyT8Y4Ug8M4/LlZ0aYFpW7JNXz9rNLB24282WFDpwqMYCVXKo3
qo53WInms+QEORuSkotgS2IOsdPKW83sGYv0hXm9JFcHwwezfhP5FNjHih+BWEqZa02JctQNe9rM
ljnmRMp4gkXgv45Q4t2sR4UN9BzCuhdLze/7tACzvBQkCsWBqS6mD1f3d5hci1aOj+LJLEPOUi3u
ioCLDvzNyQCXNFSOlq7eu36ZSJi2BVaGjhpPL2v1MdI4PZM1KnfE3df5BBkd/S3a2wVE0jga5G8E
w6nQqW1rJKI3Wr2rCsFKT4WuHk1VgJ6qZ1BlrwP91p0OZxNyNouP7/ug6P9J8Bq12qwUP4pMzank
enXLX9peJ5+AmWfAEDw8q+eI+vR6CNb5ZAopDPElYccegl2MgziqXB41eQsxObKq9/b0KsrDFuHX
+/AvczT1PrUXyp7NiyBNYZREv7iGNrBZk+BvSQXvkqVyKhtm/5Y89O+HBlSwi9gVmqhz7saRzuFR
FscCaRKKjW4aPphHl+BZ4Xy8YrIHXg5JpAeKG3Hgd2sNVhQF73jfEwRIN2zn/ruIJjwfMFfQYH9C
Mt/qPstIPyqTBdohWPdpEiz/vFxNMrjDrKamgjWnQsrA+D5/uuBFWChzPGb9iOgdcgprl5BKXu6g
Nytfg1mfw/70f6S01cZmlWA6nQrhTwcwoeEtpGDoygoyTtG1mGVQ329IDGca/US1KJGOb/+5XqWj
ChCPckdOsSaUTAVu+pK2bcjjqWUx1Nt3BOohw/b+lqGMRtArMlEku0ZivOaW5AD5emwnS6mB8KvD
M9f6hE1kkWvVoFGzYw+fEPR2d+wAet6g8G/9hIK68/eFNEb43GYle46ZkX27X8/uGancf3IvJ3oi
F9XrY4Ab0AC7WOjbI3Kz7Qjz1SGzY7X58s9Fn+ZzxY9qjNeIZcPbxsjgKD2QVVHDEJsvrET7RHx3
EKknrzjlIvwMm+8GgtWKY3Nj63goFefjEZVYWP0oJLSDm1uTnvMU+202+xrgmko1Vt8+Cq6/evKK
qP93xX9QNcdhLTY/kmcTZxxvtlS0+eZVg2xOUxIaQIwJl+hNHKjJmoG9VVvFzdI8heRmduSy43XM
CYxhT7LvbAkhc6Lc4Ynj3Od55ZL42fWkPm6d6poYhhzmrVhN97Wig9Dd0yFN8Y9njF2ItuYUrIQ6
gstdCA4SIGHynKMnN7MGLN6kPw8N/xcWa9dPPqdMUVtWyy6kUEPRjzsSGWLLsDZwivq66xHUn4eI
U1cvh1v9O+3FzvmttfScQSSdsZb47ioYLUIM96CQO1CLv8iuPQifKOgfyVPmhdCBp8RE3ok3PkjN
FByUdwyueAYvR2Ky+FdTRtc/9CUeUvxlspNVJ5m+bQWfCQEvooSKlEKH+eA4xgrFHcsx/4X1Y21U
/FSGddu72w9HjYgeWxVwVYkVuzTFLVY3UabkqYDNAuC5/zxcxQ8itvNdwvAbFFCAL6qwMcju7GeF
CE1F0Y9XLmKRTd2XZnqm+SuqYezgqAPBg2kgCNCxsji0iCFlFnVqAT2g7SvRCNTW3Gu3CWfVQ1B9
WS1VEhEfYTzToATwMIcdFrFzPswt6uQvJASbPtNkFSo6PmC2esI/Ig0RwbEX9EzeJpgzNtn6zEEb
GerKodShQ8ntJAXWbSjE+qGIDwaJswrsXKo2NAwbcEHxfBgjYE9ZTTDSSbl0TcGp/jj6KWZ8VNsA
erBQSQ6wOSNwkYdEWHQlHWdBnjvmouYQLPYOoC2P/+64Y72nxvaqR0M5pI2bV6uMI9iuIGC8SIFx
BdMk14kFkuyAtD1s0F8swDRvCxGBKbKNavQF4RYyAU2sLWkQNn4XxB1lfHMsP5g4B7BJam+EXjp5
bP6KAIq+s3pH2B9i1ay+9kGHYWEvOug9X19UwCu3fYhm6mrY+J0BbDUq4Fp/sddDqge2LRZhNI1n
kuyKYWo+FPLZwbdE8btskS6McpY1jKztKeOVZlYTrX+9UnKZE6dh8dWBw/ZlHzaPVtUEvr07Txr+
YN9WhF4j9Ix+hMT/dcYu5Hyo508ne4wr7udFgg50xsQdDfQnkpLmtcGNd1fom+WgwJzQv3MIOZL9
+Rv8hcsnjuRXocjsEHE2mVSPMbVW2l6Ki2m5fPViST8JLDJcsNq+qZxh0wKHA5g0ohkQy722QFYz
+eLxCFChAzWUicGdRQfEm5AAU5Ka4AW1wqgt6n6M8c+iQphyZfpwhc8sCRL278fkrtO10PTWUQ5d
U0UNbJGRX+lW7vrqqQ0vK7IZtRLQlvAo9yCccQVAVc86L2KCXxDcQmxCanO4NFI16ks9EN0lELfh
tXQRA0XkZDWHDHQTGf1kg7cDRDOX1quvU1pBjr2vWdgFAnwn5sr475iJ54GMfbGrvg9D25WnAitJ
AuCd01zTMbSRFCxBrprY0+E7OGqhf+/vnyhsK0w5UFgFmBHjlFN1RXf5m5vpz4y51xcwbGwFu13U
M/lVoBj4BN3OFTIPkXYpNznXzh4JiJgRgL2nCgEmUAcjP6Hk4V2VQ88gDJSXgiPExmoz3xjrXE1W
bCE4UqWro6EIW5ovoOLpFvxcJoagh+sUqWEaDBLIHUv6IEl+LvnnQInZZTyU+5FrcWN4i2pSZ2YU
zi3vNeruHn8UBy9hy82bxUoAgajHd12Vwv7xVAuRjUxVlrIqgQtxPOkpNiWTaYDIKYIJ1Ay7Sw5w
+p6SNxZbAuigUbj6chrWvVUQf6wP+M5EX+WnF1qF5WLgKya85CCD4lk9VQVTIiXs+EDmxQ5V3S5B
CMS4ZVrC6i0Qv3+OTi013HqigX2LXzdDb1Z+WJc6F7GHuiszhZWuIcK3vZmcmTDjRa0+NOvE29q2
nKIYsizZfEo14EK2zvYEa7ZxplZptM9McVz54m7QjNCYUQeNxUoa6D6UIhjAMyrzRc7fN/iHHkGl
DOJmlg/E/fVNicIvAVC/BdOl3o4Wj089L17qRcCDZLe++PmXp2xk+RUXwkMA4QRj7aPCG4BMWE0B
/ah2oqw5BzaDAOw8t1mNUkQgl4CsM30e70WRpY12t0FUCkjimSDs79sSsYb0ub83s+kpbewLzgOO
c0tJIOBmjgXOfn9yWnjOa/AIrlp2s60Eoqs1yqAeeoBQj7jpKfYn8qM707hl3i877442Wr9Pr6Pi
g+yfL/Q/D/mZhsyMRbU8CvF/2cgiDlBm9bNI7oaPCj4Rj8RkJf8aN4DBkTRwXdUiLhCcQbGsqtc7
TAPqt2vfwrJqUl5aXevWgxvWRZ5dIArYzA6Y91LawkG4QZkTV7FN7w4bd20Om3my6i/kcWJvidqe
sIANUymi0Ozx5uxqCPf0aVZknOxngrQ2Cq64KyTai3ZmeRs5L9UJQJpOhlufGz/aRq1OIJU2RPE/
7cGbDHPGMKpzs/4HHVOmk9NcyyhiaSKmTn2x4JMLDmES4eYcLODlv5LaaMLld6C5B6vq3INpBj3X
/MZEDqgDA+unpxtf4/RW+d8n/N2VShBEF25Obif43Bw8FfjZOmbCeTaBi+FZNcwpwSdANNLuLHf6
NH/VQVIExbqXkwO7ppPakXcxKvkyfRCb
`protect end_protected
