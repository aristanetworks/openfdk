--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
bVlizM9laS/4Lymp/i8kW2oNEXeFIANxaLJhRuvBdqKeBAu/BgHVJh75DPKufNL12oOERuwbZOdP
efnQBOf0loMRqqlHlOCxlTSVRpwPVQjDx7fVKB4ldtzK4rlAgO2DoCJzEoapF+dVKyvxDPJurJT/
mrNAkrlDp8wkCqcviIhyM3oFUnkwmH7To+u1et+4w37YawDR82VmTyoWwF/1hmuSgRrdDtbfokjZ
cOvxKIimtVa5tMLb/OwR1ZBvCLPEzAc9cPs63kwkazIYL8RBHGkB2Yrtw3miuXcnKvtKzcfGip38
fMmfK0EYvZlIutmujN8gsf8HtxYuoy4+Cp6YOA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="4DT3uOgN87313IGS3hz2ZtZZNpluiPiKi7r+VO5EDAE="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
BdgDXRpr8OtF8sQ00akap996O/sq1hP2qxGjJWMCcmpo+0QwKTLD3WS/66+4V6nz1/XH1K6Hxq3g
yK4EWnQ7BxigFBp7gz+9Cyke4R1GTiPG/hBCcDIwC6MHrXkxwcJMC2BpjsvNvQ+lQc8RHK3N7woV
KxOSHY/in2lKNFvHBc0JOgogwroBY9qEfc2G7/QOOjPdYJz5V/mGNTS8Y8gdg5mVFtj0ywnPNKwc
IYJSJyKc65uFo5pUpJIeuYNXYIz24Tvn644a2fVz5pKK07znLoTKLjej9X9+0nMrMlEjUR2+HhSc
SZAgjLdMlzpmqQey+iCS2VlUexDkxlacGmULqA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="0H8RIdx7TkUmlLjYLkcOhXqfIVbrU2ANuupbtyDa6eU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13888)
`protect data_block
qTPYfJxAy5ppUFlErVu/i4LTTeiZjxKZ9bsJW5SCH4/8/SvVJ+GgX405/ZMXgwXIVvwo6gJxyjIJ
UAlo188GoKJ35IvqGxuVSokTy5A5fqEC5FBZtrOZ7c+Cj5HENvgWWaV3lRqmFNd32TM3JUyz4TfN
M2Rg7G/DkspMyHlRaLC+JLda8YL8SW3CV3pgn+zPIPNs0C4F3PRTqLofsVUbYCPWcF54Wy3hZZf8
Gj9n6nTuu4JIIpmM0SFkfGLejQNypt0I0vXBf3Z4JBrIZAeWqm8bViWUz/tZy4ETN0J1hdA1MECs
2FWZlPeo9nuN4NEQs5Hkq9o0wDWPH5BFqjUzChIpOxjoiD4+xMzHPG8DefqPYN+I0CMdfZ16q/Pf
9dVyngapHXuI5r2SthmgraQY4wbd7QfgBEymWiYn9FW8cMxfSFfIjhFF4lrXVdwMzshtqj9zyLFU
4qLqo6laoHGAsbKmneX7JEQ9ruaBewlHvEWdPXFF/+tziigsdoYri8KGK777LUM/tnWjixf7c512
JrqC+0Nh7CVdB9dHimYJh4SiJ1hCVLUDNsWnSKAEgmi0jwrrNIOs8Gx8kZULwmMcZ0VM6ZSUDZ+Z
ctfANMmyQCdt/3V2HajD+qglHRBXgN1xrQd/W1lCgK+33UlYPrj8AjCMOS9Xzy5LYga6UD2Zk66y
AnqaIKfNroOVc/Mqq1qIYpBEAt/+V4n5fWielhkLaO2sOivp4xEVDdD7jhaEcwD5JME27XlDbHIA
H3VIzz+hSPigeKofaqLu6JNVVSHVJGD7wbq+sfGOeSzjrKh8aA1joE03s4UzxHOnVVXvNgJDXxZg
e6Ra5iiNVmmDyKP7W/1Ljb0qSNNCf8oPEis6QschBI12bxqspKILE3YizJAPbadQeIQbMinWREai
tweQUaLO5QSMhrpjCmEVFh3RdyLPjSRzdE+4Xwv1A2qBv0Bq3nrCnnKPOXOpmxTve8D4QUquV2Uy
deP7/jgkwztfF+k5VIpb0p+7ZxVg64oY3qlrhyYhPo9ZGtRGTnpm4fvdsBqN9+qQvJpV0GyJ09xk
Gat5THL1VoVzPWIdECtcPducJcXpzwtYdiUIiR5GJSEIiI7EbkVI/t0UAp9b3UZuztZFOTu7Wgph
rrQqjgkZb/YPFXSmBRJhSIX5/lH3Ep+4NgsWCw6sIyM18ePMd9cobYCiawpJwGMv+t/9GXPDwTka
xBYpZswb+r7wFVOL9uPf3I2qLyRWAROwW9TrgF5/B/zYyPxCVHvxQk0CSBLnl4VdwtEK3tvMauon
+Xo/X2/O9IGbFLGMBXzCkBeW0KanQJ4ialBUpvDrRSPfj22bkU0bNSUP9cqD1DIBfLfp02wayr2o
bzJCP7r4eVoIMcWXU9w34uoHA9fEmJ+Q3p7AcmzV87vRJac3zYE+k8kDJ243hVuKGsj33sG74nwT
tEt9ns6pVY7sczaTPpieLA7dHeijNESCmlZMWR4HEkNWM3yrhu2dyZII+cuFmg+9OtP1ycQ5O5bd
vtEvuaN8Hg5bWKD4iwkcLXaCz53bSxm5xLEN7TJOyG4PkaxuEBowLu9mB0yRnhDaJRxUOz22mlfm
RTEenQFYoNeYfB06V2hwTXFCkZ9g5Y5z5dg1wzoTK73eZnf/Cvf7OUNH1wC4I/oe569E6f2eHqxm
tXZZNgVoXKSdd8+3IPHHLkVDm9FT0dDAjLahCRZaDxOa1kj+C61QdN08Po+RqhMIjzlhrvGotBOz
lcBX9z0fSepy7Yt49TCPqyj6BZFphSiPRHAKAtvo10+2fjaVCL1EBPAvXUwi76irHGfcF4SqhwZO
ihlX8vAhfvZ3ydc0+N+7YRY7DqlUzzfg5J9jndsYcOYhYx5szobVvmtMtd76zSmS14RremXywng3
p+vVzO/u3IEWTyw1s4HMSMT1a7CWx2aao5g9fUEDppUuKpUf+OTHKPhQULYZGMwwDbvjo4SSNykQ
fkYV8cKWLLxW3OognOI2xgxEIpCRlASDvnydEIoyohkMzz0qiCskQJVtVNw5hLibszrk8BmCGXuL
A398mOU9lxfc6NKU6DaCqNAudHAxPnb9ppdpZWIdQWaf0yCEOqNK6r04Z76mQty7uCEskWL5mqSk
LfLiS8mGp0kSK6r+gNadMdbccDhaGe2hlffac9sP3v08Ycw4XFF+gHZ39ss+b9/sioKjdqYg9CwD
3hz2iDj9TnPSeVxxCkBohtsO3N5Y+HFaopUgfngl1YbhPv1bWdYTgtcw8eBnRI4q0wSSS+A1rDVf
TZr19fsJZW6qHKGgL4L1q2p9dEFxGfvORYwBuvI46mt196GROhs3jvXKf7LU+YMuSMTntR5y5mdK
XXG2WN5s2RvYapm+WMl4i/gcc3YsZ3bLXQdivrOTOMTeDNEsO2SfuboemqSWNj9tH8yD8lD26eR1
kiXwhjjDKxEpFEt6AqcqQ+Q8jeLtcOdTVcmw4uZtemmIzoX1RJXWkl3JJQQ5tPJbOjBMjJkTai9e
O1juIQVlpwnWRjmHd9Nmyptn/7bdvVZsNgnslTBJ9bKtpQ8UFdaGZUCo/agQVuZIy8xrZmBBs6F1
rhR2z5X1fq8dKXaR42xUYPRgROHCyBdAoWOl/vP3hh0JWLr2DPHHHGaxKWgxSxmFsEF6BB2eSM4J
V9iFTJxu6ZPNRDynn9Mh/1XTlAmcYMIsdfLbkDFuaUr4LRcjY8W3VeWWEXDH5FsxYyVLKlCs6zds
TubMmFYOvid7DU+6FWpyzmcFRGCiVjiki9c53dbtZMwj1e6K9sSXEtmgjFIBJSi0uPTyEyRHysDV
1Ffl/CtrlbfS/gusU4J2orefN8L6XQ0GsfSrlyX0/tAoiIxD3vkqVq7Gc0DOpojUFPJWHjocDSPZ
cpTHWnn/o8NAjrao+I+Vu7JjtizbzZeYswt2+eJ4FkArVxc/sHSHNr63bELUhjfI0L8xxrnlZdYe
K6Huvozp5fvudPD3OnBZ54pgh8mX/MpIt2c6x5+Daqx/JwfbWYCM05eOfmOjKR1NqeSlRkXnVwed
u64HT3XJucwF411z3bRsjvrRCG8LfVDp+m94694wlgcVH5TDYVxE2s0G0DS5Nx36qAscEWZM6JCL
F11GA6QOQ8FaXIS2WZfrnhwt6uzznFKD7jVf5mya+QbNluz8NfAhg73qqYgD3jyUqjyP5hIN+pft
IFj9EHS0+pOC7T+1E2CiOGwXT5PS7AoFHtoDPPebPjsIt1kRNuREX4nHqAJFFe7W3NHd/amU/38J
P2s67T/SWoOJr/i0pkNIVfOOzAO77bBQ+29xVtmhdkNoIkdX8yxAER4emMZA4PzkHft6ZfWjbjy1
d5lY+eHhw25BGAn3aNNMAxON1h2JOQO0DfFn0ZXqJKmrH9TMr7e5qfERQpP5O989tG/DEl+NWhsz
VMe0lTzXlhBIiywG/7D2a4WImjMUkdLOslpD4ECVbt49sQ9WVN5k18fzrFVq4Ez9lc66CxTENgBf
XMT+LEtY6/p7VB498Icc7LD3V8X/LgAIlcN6DYHDnIXj2VHSRAhz4GqjJd17N5rI7LYuPuj8eL5j
QEz72HUziRapkl/Axstr5JzKvlT8zYBPRmD60oLJq9cBIui755snviHUJkN2SLkv8tUXVwyhAQ7R
qZyJqVl4WevCm8ZZh2uKWb9iKLhibMk7so24ixfHoU/5RQ16Nj9KKi+mcLB3Dw+1t5iL8nJb/4xz
IRA7nlKwpmxfyUNZTLl/Fe3zpU2r5AX/SC1/pEB4NM0E3xgsqugI1LyCvzTqQN5MHjaW5bluVPE7
xg/iAbNhRz+8LOnKxGeg9ROycm4V5A2+pkNWdfQXTEb+PBBjjJBgokvLCATdXS4ZGPRqtilg9Lvo
52iIJzBVdJl49OrokLHgUxYRhvsA0s1Z7MVOuqnWhfZ5Y3iZ9/sE3ZFKNnLXREGPT+kKmIsrJyxM
OEgZQRcrf+7uZmy9x3PjJLh3qOBspzKotdpjDhyqMwYAQp6jkuELNoKLX9j9j31/zgQia/4Bc/ke
D8tP8eZZfvsoTf2iCREKyqU+I/9wuaaeLeOQdYcjlfmzpVlOuwBOPvoSGncQzbT4sI201dOa/Amx
q/xQQvyXwYeq7nJrb0chKOqWUlgW9W3sN/B0UwI49Ub62N1uREsrs7vCG+o/ttg28hYUKJ1MgkZe
z1VzlEmyPyB3kgKJY+j/XzfnAka/+zSz+eKq76+3S5LjMaHTmVdCxOPZ4UZZJqHLdExdDorTKAqH
FNWlpic5SlZmdWAuHAG/bPUQJv0bPGQoYFr5E7S/q5VdtXTS7Wi9u1FqWV59lbk9lLXTAj23mGXF
wUeXkjvHKgJ9qbpZYxcn3tT/gS24s2O0yoJfRH6lGRbQfYHeeDFD2L+kCuSBwGSwJ10YSKJOT4wX
Rdiu1KDMn8R/fmyA6VymKrTaZ7xmWYeU4ZxrTvash1mG5igNtD5JK+xdQGEoilzo+FaF3HkJq+Fg
1OTwAGvIsnXxMVTyHYAQs9cJv/YWWZObUr5RS55Cl1FvHfr1tGYmXd6RIw5lVDnrIBunUEXLA7UI
HdHEmtFCVuDuTIxyQ0UogngGMc7o5jT1US4oV3GYpddO9hrmD9O1qh4XetbTd/v7jgUyRhaAhPjp
0CY4rQhJeX2gmnL74h5ecwGVnCfEfQDWDuVYILEl1ZsbahMZQUFG1UNGpM1ZKxGbhkhJ8KZbsAGL
MW57eWklNBF0aztI40x6qhahgoGfyeamOGaNz04T0FtI8TbG0WaNQTajofOQi8XmcS4BI9f/4ahK
+AszemCXX7ja7LUaNeyW6VDvJN9R9yx4iq5o3DMQx8D/Kv8EGG3b6XDKVFbKBiI2/LXc+/tMBiFz
5SaFayg3+7IG+rTDfVZIVoMFgEYW2uMSDmOZ8Hqi92uxNjTcswLMqax4+icyFx/Oqar13fRbmFl3
dysawUzf9tAnlWOnzXwKLv9YZy6/SQE06P1xvguaAfR9Us/p2x56y8JpbgeYMPnvl1PyTmkFh6LH
bWTRBJZetpWoG60fj15XY0bkiLogJtuL+FXTWQLfwGuKoxHekh6XIrZmtp9WT7fstvQzyhR7Jj2e
mzHJRai4CJvPbbG4RgtwSbrEBj+b9dEXkL19guUXnqdOE2kHmw0FzYLEUN/H9+ms+C3J3N44feK9
28WY/3h+ljNzil+eNbin2Xd8E2YM0MCB7loYwg72OUjNRoRWX3uDdoIoEbypMaZJIqcAmg2Rz0TI
GuYG5zywHwO31F9fAFnPCJKQwGDv5mi7fyixAr/cGXQu9UlOkuHrPsRuHgJD6TdYXT7xU80ryqEO
tt8b7O+UcJuwB6nMCeEDWT5/muHGsGAlHVUC44Z+L4zZlGrsoAvz9yuFajsKZ7M6yEdJkrM6lp1P
hLIIdjAlrEn9JeNxFPX6H+D7UblGZJd/TZ2DGZJSBKpV0RVuM66GMBGio7KHlZYunyg+3UL7uBT/
YJOSpYfQlDrSMoxmxHjMRjoNEobDvZi059r0SWWcFI4IZysXIuaEWhFnbclWstqRJRdn33pVRbga
hYirCEbya/epVUkiyEzf0rvf2PkhwJduAfFa9fkuwa00duoPLLePf7gFcT49iL6obzmYt7kUfEbu
O+R/q6ncNjgOHH/8xWDfVpX/YStyRu9VcGNaMaHmC+g+HWYhDiqmTRTmfuLuv6NKjzmR8xT0+Pr6
/9mmnMiWyQ0KOauCZEIl478n3nu6+NRbXg+6aDWyMR25BJn7+6EI1hf4BQEmbGnToM5HCShNk+h/
rC0IsSIqT4/5+SQpsh0vC7DcpI016FubAi+mEhV/BStgiKp55+uLNbTmfnLMCwT9WSvNtXVSqYbl
P4NMkDYp0Krup9SEeX5f6CMzIe8Fz5Mlj2g9SJBMyS0qcmB3bfRcGw2PI1o1td3yQFbGoo5dlhzL
eL8sqJkG6xY3v30HlaQvUwH2Bz1PqS50EU9/aY31R14NQkbNlZI/zTx9c4TnTrJYFWSSRJ0PjPex
x4dHyGP1E1HP7kH8sHGZcyx35TBGsssVzQeXyVsUTrs0TSI/UMY8wgjaNVTpFTwuERwlxe1PW8W+
ZEcXGYmRvDJ587gG3U5wdDXoMDePaGn0VSpLWqYfl7xXH/JBtagvv/ldLTM1wRFnaL31gmgU3PyS
aucqopFKofGWAPVhn4hmW5Ec0FYfEi2BmA0bntXTjicK5Dcdimf3ExfUKmKuokkX60TozHtxQ7pB
Cqg1pVDza1Y7YKz0KJG9m9r+cIJmnQelI+DZ3IzE6COOl5eRWd99jpi/LAH7s9dBqu5Ph/5tLqfh
L8cZ5Y7PuwPtZjXhDvlKL6zGoxyhhFL/0drFOn01yBY/VBE1kpJixSwtOSh2MxdOeMqkqmADoJJb
S1LRvEiie/RjRNYSG7xjCyPjR5Zope7wvh36P4hr0WD2kRn5xqyZkNkX9Of5gufZcq9R9nVzuTKc
I2QJOQfqjU7Xo83OidvCyEQ3rGyC+TAS07x6viBdNWGd/nQU0wQW46De8BbL81GLOCRjsOpFoIBe
ua0traywDwXxiAp0LPqZfXKGLAVcv5AixHDdA8ILW+8+d3NTOzBAPviLVQFNne+mx/UGf3gbDCrr
t2Q2XXsLXsk+JQ9CG6DmF15m4I2jiMMEc+2bXUglZoBmGpd32osqp/w5JoZlsJkB1rlR0hXFmzIx
qN74/Qdi4m85Ytyt2Ih+HHNtwB3NqvFplw7FhLWE1la8QjonqPwRrSarYvu1W1J9rhvzI+4B7Xlq
rJGtOJUOFiUMDxZ0XzVS3FQ5lq5nTBx+SImdNGsM3kUBsOd64VBwjOXozrGu2NutrCkkl4J3R+Pt
Gq4jraSThUdXSiqFECF/+2/NiDU3NoS3ZlyLn1Yg49B41+hxpQxJWi0VFhw71Mfv1hZidUMV/Q9z
F/+yw0lIwTSj2wthwIAUGVVciPStBehAF+rpBgM3X49qSWO+PZO7mNAuy055TsStjxxEZTHquK5W
vbhS62tIarGtWy/Q2ztcxzSR0ndmsautn/9cWPs9WRMlOoy4I+sRxt4CIaxkp5lW0mCpFNuRb4vi
sSRvfclHFFTqJ34btopsw/BmGxfN+Dr2sVE5imGbZ9/Cb08Y9h2a763VRFKLS8oJtzT0Bx9wyjnW
pPLH91yMhDXl2fGMIBT2FjwT/R3y66V5pXQqDl2LVBu1lbq3VIIO4xKZr8GShdLuMGTtM38Aw2lX
zMLW4EB85YMF/pFkbExtdKxSYZSJ5+r/n+ukEeybSKcFqXHa6YwjUwSlmkIr3AQTyza7bID/DZXN
JHtE+VQB59KWm8ZEJ3YX7pw1mgcUQn99CzeKQPvi9Knv2oTlN+43eCapqDniJUPV9bIaf++A/6Gi
OSqAT1INsxyFkTCKzR3Q2UCySEOFCWz97Fzbh0PA6LQ8pHzyuO63JCgaknCixIxBrAaHKzY8k2X2
CJem+1BIunYEfsAS7VnWcGXHnfvJjz1Q8CHDJhm1NkBAcmxRyTa5xFxwHfYjB1uUPSevX5n0ShSN
5XcoK3CVARua9nNozUxunnwE2MtV6UTVkwpgxF73j7O18U+E8pT5oxIIG31RyL8+9sw+iI3lXWSV
Zc8Q20tuclMoGGdWxe/viG//jjEZfZdDDPflpOoEZER0ScUaOxGHyc8sI7KRQXTX1a+CAgsKbIXh
JdGxnZWZAj+KqKHndAdaMWP1YJOdJQIN6xv1d/OtjgfSVsrx21e4ylNITpz622RE1eOMvMlXXpaN
QmCzJ6/oox54b8gsLRdDfD/I2Srb42ABw+obg76voXVe9T5YAIe5EjKY/iyWYIMJE1K9sCLTcRLK
wr/0o1dDKBPkdRBYN3NqjeusFWuEE7fOT1DeZcrLX01P4H30ruSx+hy0xHYJrIQcKq3phfdhDF7x
eQ0Sfz6GK2PVKlPZvInP4TqUZ6TAf8KgReQ9EC7FVmshRt9afa5VfM/zRJOUYOIfHIKccVTKkY/1
YZ9rGHSm+3WTGqhkFY254ugqV0m45R9l8oYNxtIIB3MAdMG1+qaJp29CiHHR6zCPwBQOlhkfLAAo
9oiIuI/5UqS8KO/j/IMniKOjL8KzNAtkvtjLwq5yKBueMeFdGRkr7gnja3fQMsfLYbVPE441YQ2X
sJeAnMxvO/xvwKXI78nXYtOtqZ61KVu01x2qYXqXw0Pq8dZJw+eN4I5vcvArsHdp9E4HZfLDHFDs
skO7iVWRUwJtQYigWGPayaTP/Rub1FdOrYfHQdsOOAbPe0iT4bfTuOjeS7kzbw5qxNShaCJ+ad8c
TukNOnn7c+QAeok4a+8eyHsdN2xSXlFiEb8BOWE2S60atdRKWFwFMN5INpBvpKM8b5BRC5IgRb5Q
oI1m0090zy248exNEExhKO+9VgP1mUrmhK19FX6bRjddSbR98jQ8BT2VXQqfpLzThe59ZZ83MVZm
N61iJ+xv2ScbkqMStNrZbd9yUs9wvALhZd16w6iUtkHgegasq1mL0vypNAj265nQn/Rfxim1VeCV
D79jdZPSm3DRzemYG2imnT6AtgKpUOtll814t08LrGo98mydKP1ngG9jIuamDxyMr4bkgIBu/tFU
AXsck/A6mb6OOt5axnEhWoGZYS0JWfPSnKukIXv6lG2G9HFUxi86UrYTYr8zhJDchf6TpwpcLie2
yoAhzYVqi+uuHcbaD/aK6jw6PjCqH3r4ZlaTl7jXjzImqm6X9bb+nXuQprTXjEFHhgWuxYV5hS4G
pywMTey2L3RIemYN6e4UJoCSfEx7eL6+QvFwuCsstik2+OU6wxqzxi9A5innkBHhWy+OOES/vM5u
trw+hT0GfG+nFhpH5xy5jqGVxr4bBSaJjReaG3YbBMV+znuucWPBa7qd5vR+VCs78RBcreeF0mz8
WwNF1i6/bgGIeaZS3k+U34rSmXPIxsUxaCOi+0w9696y8FKeD/ShWX8BTPY1YFnXb825sqXEafsc
UvmpBsn+MTrsxpTo3cyaYsT7z7Yfg/XDeSmSvzhgz4slkLq5H7pFpjKe05Y41E9ibUF7Smjcu22Z
FPFM1RgQ/lSJD6dA/ckewg6JvQBmAeohGv+Zi9F2iIoGGTuUcvx7/zbqac68YtpvncczSd2hLZWJ
ta4YQAoZ52WTCVKnT8JzboMsIexYn7rGzytMWFCwmDJwRBIqb6mSuRBfBqlOgK7jPH1pIXreRob8
8ItvRGz8JOlXsAOVwSJ0wX916v4gSKif4n+fQkRwlPntt21nhp/W/E+jYbafZZuxvicWgF11+zJs
BsaAvdFZj75D31vhGN+r3htaOJzscPfsUq/kl65L6A/dx7ATlGZFaTI5y7hPb6Boy3tZW9woSPw3
lVMbzZ0khVdCLgvf8H65X/uJIFjzlHGjfdjwQi7F3kBuafks4PaqzHfS4ZdLGObtPR5jlES7ZCdt
q1+VGYBsCOQEa/AFOoTWPsvBSpjJoZSYXT2JCRIJpU2RMwJdDn/tYWBKXCwG1cmPIbuWUkurWfFm
hi4FTUshxhlNV3Cruwxcm6/JPYTEF2YwoNoXn3lbv6C4cKon7GvepsQ1upkUbcNXUtsJLWx4HVbY
ToeRS+tO1s0YjQ2DTbhK6vGcSyJD3F5H+CjdLLosCEvaQtppatuMBlWZgi/ili++8bP0zPhjveo4
u/0y8PSZTVzOzj8acQ/a6WXr+YHmrF27dZftAUQwX0DvwqbrL79BOZVn5f8vIPNFHZJ0GwODdsQR
/ZEL2WhlXpeNIeohwmZzrQLXgHG9icNfR4o1vfG/IMr+7pwROWYZON60EMGCDcth1OS6beOJgggB
H24ILyvAiRFyEL6sDdWvkR5j2HXFNhHRMA7521j5UPeqEmOOj3lg+jMZCINS8YEaueQg+tl1Zl4/
a3iajIbhrSHjRwC8/9w5g9mu4c79agbvb4tdtZKJkaGziNzAkxNA4Kx6o63KUk6zgRctkU64PdFl
YMtkxGIa6jrFG7U+xR1XI+dDcW+pkv3fhRPpG4yiRWHMbAKvBQi2Td1ZxiKyoODIQVdwAiBH7Ttu
4hKvKLNGj/Qbx2sjrO4RzC/q/341tRHa7j+ny+ZFjv/IL3RwNQu4FFKQQC7WZragdBUYQSLv5ZpN
V+wBPFukcPOCkSoWvIJnoHpTDwiNanohjJjxRFjvnPfn5rTAW88zl2hydTmzbJddsJ4kSoWtAQTm
u0vy5cdkBqC5kQIH/jpeKWzdV4y0X7lcrfLGUYAFARSerB9SM3vZS8utJmsKNTq0EV7Hbcr+00Ca
7qjHtLmE/EireAReytZsCr348QQ+yCzmLh/+cI06Eztz2H48vgEvxIkZg83rQdFkxr6pv4HOybxD
hqmDc6Y0B+X98jonbMvfaO9BLWR8duKbXj02yzCmjFqzNRtlC77YYp2i6qG7ZqBTSuxPZvaJWcB0
mk0twLvQhw2mVOSpTbp+3c844Md1tYD0bkK/DnTmQkPRoK8VRuc5XceE3fQHw3N9abMc8MqVE094
R3InEmKd+dFdxuiW6H49ctBzSEIaPQQygvIn8gmg0INx2u/x0oyp41P0ClOpxnp7Voc2zZr3tNde
hyynarKxtEuo7+f7EFupkx6duGbb1Pgwehss8j83nibsp6qZaA9tUwkQxRQwcRXbCJcMUwsDLxiw
28rhFEAEZfyRcQMjerTrGe/2UvlVoJ/hcSj5FfBprWKbgAJpF6y4Vo1AjSqlU4GQb0GvmH59mWfr
Gl9K0KabeW9EQ8I5ezzOZwfQtwKdtQk1zJvZsQ2j8WcFjSR9OtJk1P4mrCSBAJGvk0DeyP0X4LLY
ggDemIwNnCcF2cBRUREifKkpUtHeqmpvGHoWJPe2OLYJyodixOYlIgWzCd2r0tAlx4G+qrNnFn+h
T8qevxhDbt7BGrs819Bcj1OOBs0kMDn+ei0WGr3iY5+ywaibkAAP+7shoxClyYqYHX9SplXHdzfu
jzOamf+b1VGQWtSr378seJ6GABYahU29v5UUECBEEukERm7efzerEfPSRKLhCZ9u5H/aNjg9W4PR
+sITaINeayoPtDeNuLLB15S79y9XcBI5qm6zw6jTW3g/1c32IK1x0AIndaMne0n5WDsk+iYxszP+
u/AexeHWUibdv6mkoFw3wzf1O9SAuC5ZSWvJ3y0t91a00mXvtR9vaCTpnhA51pY//5pvg7OJfSNg
E/OLcmKKIgNc1eSGFsDtj/Lt9bWCaroqXt9KyBEByZNN65wvtlGl1OjrZh7FRbyym9h37AGU0RSu
d/2Ua6fiCSeIGtE57sqdhRSvLaTBY9U+IfkRSUQn4vWOHSwMC1vb2rGLng0yW+Z/NraiOKBJLv08
uMoJr8Dp8mWM+7ggiNgf5KBzvwciKSbRlbjFc+EMlXhZouEWDGdsAPIgX7CCi9bifpqyJNnKoGIX
OpXYvmKe6B7ufuG8wXyLje2ItmJ09a0z+z0xF1aYQNxzRfPrS8O3/HQqBLDvWiFYdSIlxDuv0dVG
zN/H3k6K8gUY30SSxBrovIh0W85FR/VRS7ZFH7HS+hu4718ml3D1WDuqagNP5xDQfIgbDUpHf398
HsVPQpdTCJaFW5z0m2+qG0yPDp4mpqHeXlsywlBfK8n53ZcdVaaJt1K4jqTEQcEsIWHCSVtRXJ0/
NdWSQbGKqtnetxWFiHj7F3hmfBQps2VtmbZH43O8J9gHfR2iCE+Ejw74KirFuMT980k6L4/PwaGD
4UpedvzJcMvFWEddRUFw6RF6mQGintOR+IaOKROY7y6HLXv1vXDRFiPYu8yW+ev+LgNDyD72RcpZ
vmZOywDLbObL4plUy3ZpvYBoZr2NbxMxtOQCmAlXkYiwZtI/INVEJsq3W5Qkm2QqYWOcpfvMELYa
ereXjf3dWE8kHSfnWrLQlHb+D7COzyVaUbpCphMx3iS88HC+PAAxaHz69pUC99n0tupfRbBiRICl
FVa+hP49fNVbp49d0dEhwBLHVvvsrkz9d3bM8xGhF0lvxiMRNLah0Efi09BO1GovCVkaCVK4vLow
rb42sur0fvTZxRE+KIgJDqYUKX6A0qBA4svl3cjKfVFk7upVdLfeuqEoDWATyMy8Ft7JMtULnT7b
qFi3/TubVY1FZ/WBRLHTmh8Mw9+tMWbpRigrexAJcPqhJMZ3hOCH7M7OxzFIeWRPVzFyx8r6pmph
5FCW++fk+MTksvbNrbW+4+bk/CTLH1FQk2BDjI8DjMaYNYPtOvKFGyzaDJEhgnXUwJeVl46OgrVy
Izv1U6/nvyk/JnHzAHTBzou71SigjXrm147Z215GasbBAFJ/8DnhqJzXat3r7S8Jsp7HQ8YT4ThK
phXTS5umvOY7Kol6fEYO3NaNk+owum3dSj28fdmpA44omAvXU76tsF8KLKnnbky8E/jaYiq3aqb0
tn6hjqyozVlG4MKKzovZ1lv4wtEFBwhK8nt9BdkMf2JqWYgGo9lNztQucmiSiszvUK8UVrheTviE
A5QoAwGtX83iDMDSa4hIsn9jYhMuMAN9xKhMdvlHXH1drRN3MkAVmk84GSzv0Skz0FItySsblj88
fBRQwjU94WNz2DAdjBvAx0vJxOc1avW9HGfKIUkO6CLQxA4bB45bPDPXAgk+IVJrdTlvUnq+e8I1
NX8nd3ZlF0yVA1/CqTEzltrA/C6BFo11rvTCfz9gQZGkFHkNd+9uTsPgDz3ESzrTVG0GBSMxYy7P
v6y9TcrA3alBSZBbN90Ar+RIlpAcAXutgbjNJGNO9vRnLGCSv2rwTDOrFb4M01iMNSAmxbaitYul
j8GZky/i0+03w+cQvz2MBh1/dqS8RDaHnw65KOLUlDwNZNmLqpMS1c/NTkfuirS4R1QDDVtb9Z9o
PFXkw1YjT2yBmtatwW2MnFPjc/dSyRzai7fY69D77us4ErPF4G28GoMQx/Eet4w07BVUQtuD4bDL
29id9cWLNhEYxg+xmrd+1qYh7qxt5H+cF/8QbVKNimVYD/RxmWN7H7SktqxAlRVVBboqqoSIesyK
851l9OnpnvBZ+e3K8O8iI774XuXd7SOK4EduKLSjeX3BaxHnEgXOix2JIYxPtbGcc6Y39tmpNyrK
LJnvsVFguS3SrzmLR69n39oGz7o6gceEotVXSbSl7sW1a9eDRPRqyWd1pQnSnca12tXPiLCkvJuC
xXQTmRmes2Xe8Cgwb17AMSFGFu0s70qC7sRr+4UPYVg7P9FFylFB5QdC6b99+nqmiZ9ZF0mdIaUK
NAPwhIfVUICiH1SwOr6Z3N/aL2sxm9OzVdJ+FiqhOElPAgC9/E9oTjrMka2JAf+n8bQDEd9zadWU
oIA2KFWYmnIOwvgC8e1QqX8iZ209LnqDegKX31dMuS28iQE6Ohda5fyVoTJyrqo246jMW+ERQ2S3
ZMZ8mjkSPIP4/1QW6ACp/bFOxPUtY7I7WKXQel7Lk8gFBfe+msyERmAVUbTUttnoRuBuBO3hwZzu
clbtB4itSi8SByI35qv8pF2e0GK/FNcK+jh52GbVMu9U1mg+1mfjgr/1VDzTHY5LqWqcCkqI9plz
xolBrc/wMG3ePkq5hFTdp5vZC+xxD0cBsGrXyVyzfhb9OwXhyuYUCAfE81Jc9Xp22HwkGoZ6o/LD
A/hSVfBaTy1qwaBsnx4j4snUGoov966mnRHV32DjYwHkAZkjA5e9HSLpj+VwSp23kl2HGn6ki47k
NuiV1C84TBpPWoCXGYQGoUxigmyNRgxuo+1bWJEda6i+VAi/A9LXb7ImqhN1X9e5l4ifet/dRmCE
uILpG67sHf+j62vndRyy3jNDwO9z0Xhb+zlK/2ie3Q1SgB5c2t9gA74H+rIZfngLzgD3sUfOgopA
09jmZ5cmsM8KXPZRwnFol8Ab+o6LgCsQ7XHHFallJXAcQXk70XlUnW1uTTIiCq5lmAP9V/SmKNXb
WEYZhskY31JJpkcIqnRahcv3sPBJAmjXiYqoKykbvOHqjeqUUuvh1row4Y+/0mfEFC8QoP86w1GK
b57HNmvdaoYIQLvyQngqK7C4Q2AEDJWQgDEZNchD2KWvSJhfxLing8M7WEPXm+UD8nL3h3otVxyn
g52+4e1nWtqsuq3zEs9zJhbZ5K6m2SlAui2+gQ09Ni7Ew+DNwF3QCaQotKJboJjBMiWKDL/pbQ6h
ydaeu0kGsmfKryHWNqvWr5Sds+kAHUK4g8IY50SZfswuGDvPVz33hfmq4K9onIIVhyIOWxVR7RhA
MDT3Pv4uI1LOVhe6PpG+6Mdpi/cg2HtMa5+ylz1AjV7Q1Lgu78rWlB7FOAhbIpPPDCa4JMrPJbg0
SzhpsuprAUwMeyBx5e11l9AtI5yBDrFfkiNY6gBaWgQ0pTJeEioTtW9w+jQsRvjw8K3UCgyWEGap
XaJmJHG6sORRmfTmzfww7+Xsrb+g+HllZW3VfMPLbZLWFbC9Teun9lwaRwYSwhDv7TLtaQtix+d4
4HeyeVEl1ZsuCKsKPJOJIe0uzPQC9SdRkwB9O0VxEYpct/3fbnffbp1QAG0sUHKzzAUZd3GuyjJq
93aHHW779ainL/MWbBuemYZj6MzGPa2Nlxwas5vNIdJSgX67IzicsX63k2FPquIhAc8dVQG7gTiw
1AYRdE0fgbqHvsErPCoD8mO0JuOKsSVV+OIyIw8iDznZg1UIj0WWuhzN0U4wJtQkawgTwL7qyHo1
qjb1eJ9fCn0j/yjtN99aGkj59HTziwg6qS1dw/uVALtFQYlfXSm2cU86wOvX4AgGtBP/5bRU4V8w
4YZimmgx/yX4aWPX+l/JYOPydzQClouFdUKzg5TA+2GQuG3SBJQLDcUI/CmNoh+84QSQWiRMM7TX
r977prj8ycMOqwagAP7jPqrjPqB17oGD8mA/EKJke2aF2oRj3Ic5Bv+EKDtPYvAO1JqkKceRnyrn
fOMiOsP6Pba8wJeCei/eF8yWHPw5spY8kCp26vwtIf+cvtMrd5r1STas0GjZ2NSzcMbL/y+zrzWz
muzmlCOyvcTD5z2ySNF2m2nnpGCfoywX6JOjxhigWcX7oBt2XwCHjqhuZ42j/6WowUe0Od7lgZhj
0sWsl1Fp44E+NvoK/iM8Oh5DIfePRw1ea7i+/8mHvt5uu38+5qahFoCoC4mHCKbD6t38zh43EEMv
IqwtHRMEbXByWq7LZ6Wau95H+sr2Uni9wyxZSH8QmJ3WtwFKQ8g0+i31jnFnuBIBhs688X+IKZRB
VPWJuO3NtLyJmNRyuf1kxeFgCZP1u/4rsssv4mjtTbsNpnxehm4Y9uEeiobsBnIkXKl/i/5frVnw
32VXYNTxT0qEghqe5yuahdGLa5PUuOBzoM5mkem+R9Ab1CfXMH83/Qel7Yk3+vJRcH7zueHe+5z9
IqhLsKMMkFE47jmwk0Ow7vnjGicWNf+psm0C+PeEU/zfL2kR9KDCcBGvjbLQqK7d92pRdbZZNUfR
wVEFoUe87u1WDRBEWG4OxHc7A1d5lLpcsKk4TDZjLI58b1NmP2JxtNtBRLYmt2g1S6UpcPLgCG3v
P7ZjRJQrF7ULV/AiDeFPIlVxXnD0Zewbm0Q6rUH7z9WjtTustzryxMlqaX4WzXMPxpmcCZ+3a+B4
pluIwiY1/KDSjsFQwwZ5bIlZmJUOqncCzV3LEeVAdUV4EknA93Spo9h+Gub2vNeiZUENPXn30Mu6
8nT6gOErMqKKiZXZicpBoqSyMSVwjs6Eg9LEGs5vh5fNEKpRP5JSPCnmVgQWg1cOwf0u7612c+Iv
88j2WLuDS43alkz2l85lcNlfX0GahUNEeGddNHpwjdBw8K4HbdINqIETnZBdTsuHq1PorJHmZr0J
jJYcshxzonTVHFDCpFc/4G3pUetcWNnD+O+qGjkqCr7xitpYjvyr2u7s8c5c2LuSOsNxHWCV9HHf
t909UNwnI8ARykqLXsmBcxifR/mCRrwLtGHtQsDPOjO35cSp/CDYQPvOtlHJsE7YDZ+ukd+/lXG5
Epz3Ll01Y9z237fXkLBR7BBjvVyZYVBUxPnqUq39RnnAxcAkQv7cMxDpHsF4PaZ834Cvf3Ie/XN8
ZebpauKWfyObcvrHQjgaNCQYkkF9xjguw6PCBWsm5C4x0DcrykT7LnLVck1Odr8D0LNHxwJciRec
YKbAicUf9Lp6tEwbSd4YG5NE19F83QDTUIuXNu8WCyMFS5U0JoGLvJt9oVyfn+ZHkWwnyTxY4sJm
TUB51xvimFCLs1spxglJlRXrGMHbttgX+6eXQRvuYbDdhpi736jjGhyKoNmERS/QHdruyE4RQkIG
+6YVQljwFU5QLI9HvicMZFx//Gt/QBwk5prEYKJlvVUNz0AMghc/hdo++xN8DbUiHQG8ck+v13bR
zzauz5orG9hfpUrMdS0qOPy1WmNdRrK+wasSqeDAIUySz6BA0mV2aIQvQg6GOlKO0uIUOq4eS+vx
GHp/zTnKHgJJGKQk16CgYe5WLp2Mi+2zgvCHXyDbJ68jb37VKndIcWGN4vIbgZ08BL9E3eRj4Bn2
l+DfFx0WaeiaNm3l0gnvdOTCfaTGg6flIjZPT8jeFa0KDSW0LmKCHCvADNQnIpu7zqrLcZxw6I7s
dR7p+SLHFNq9nP9q+RCJeDgB4xJrryAXnk5PI2o0mm/+kZvULlilBXfNlnFBm6LXkK3UqFQ/M2qQ
+ExlvpSRRcm2L+MVZj3x5yySuPNO+x23evGjGyLnkMNtCS5LqI6qv0D6BEZN70anvlHWcB4uzKM1
Pzp/TmkDp82nppYR4AWieN8ITWw4DxUz+dXHmkkIdumQyzwCO3kk0cE4lYGzP8Tswf++L+OC6XU0
08C1MI6fqEM8kMcqXrQ1s2LAFOvFuUKhnybnzFMXnObe3CLIOPz7QJZlm5a9LH1wPDZtx277UPXb
5sv6I9NbcZCGGfZi81APd4STsuvUn6I0Y5LfM2Kbtum64zkcK5iFcYO941TBM8M+HH1DcUHo/CXr
+AJ8dL5lel2wA9HZTbJaKsYj2ykzYp0EU6T0Mr0MtsNjJK6dSqH7FJP0yo9P4YXTJ+4Au+ZjFEkn
C5ghGj2s34WjtnrV2soFwteHkW4zzrnsGG87lW61+NQqIGPMiVT3oMRwlDzONR6n0qK0fugh6lvs
yW1GzNzonZx+5Ym2oyNjk0hpB8T13VzCHarHl7QmEPi70RbwsNaNp34yhLBhYCwEQyU1TZAHoSJe
Se8Fj8GL6I0/0J5Lp+Uq7iOSqTyZMowcOh9Dwsbw7cpXlr1sPl0kPm1k+tUaglVrfwjbDvx1U1b5
KicfLxhClLFvLBEWK84D0o8/kN2/h3qCgs6I9HNWXVlOX+u+MZig1TTGRdjpk72uy17u7e0ku2qs
IuyEvZKFa76F91sZW/VVzy++dB8wezludtbQiKe4vllfFgn2raxXvLVWATeKX0lPu2JCGNwk7X5C
2pz0a9FokfJCA0S0sgXaEgqA1zM38RIp5b12V9dF4F9QWwAD7VHhOOSLUyL9bCyLFZRqVWSCBgbq
VAqRxCwY9fxjjF9nXSYthvFLCh1eKSRvBMG+CWGZMhD5VHGkfrexyP4ySIICosbQlRiz8N654riO
lFXmYQ4tQLkkkoSxRBJ+PPE82FpRGZMEQTDLIsn1Z0kudwFTOCwAhy7e/7MlM5kudFy93YGKYNi+
+rcSHp+2+DJ0EZhMGeUN+92+PtNFHEYsyjIibMtidYvGsVWnD0nf5oBNjoQTq/Z69yPFzGNiFBzH
WsHGg/zles8QhNjqaydD05LeCVUUBRMIekzIPf+LTwU+YL6KCPatXmBxcGX7gt4fCcAyEbn1q1y9
dnMOvJp61bs+85lrBryUKkq+25pZH3TH9otthwqfXqU18uyhchwxDrCZJZ/IgA7gT/ewTuDm6VU0
4zCSKtQ2R2OtN61sjcPYdZKiZ9CAqq/DbrpijDQGEoJgRRpxkhU1B22RoEya0XxDF1vf8gX3gt4+
nknoCHvB8fAZ7IolIU5VKJa4HpMkfAQCZ9BINP5tAcztfFuBW7cN13D0/oJPH8ZC7p0otXZtsJij
pryQbK+i9g0pOSGCI23VCRVR3TBDIkb1lT3NFbvdBtqq4e8rO9r98GoGP6yExuAXU6QGSTY2d/RS
oGR/SVR64tBiyPoc5EeN2srWfy/ZPPcT0wEs3kTcw8r37S9xSkiPn8DJrnSciwa8DB4rFN4FzB8v
35W4/UFxyYcescWUthifjM+zjcLz/pfjZeTbCgPqMwSwZluxLbd9xVmBrqxDh61G6HEzFbzCQIym
2XgAWmxbQII0Hrp8eduJaVHaz0Iery6i3TIVor9i7axeCtpYSOx/7tYFL0WByESmfCiogzzXAlV4
uEyK4f1mabJInNU/dtRwJv4yRhS74/5NJ7xQht6buBzVbLRD4ah6xqrgwYyK+LLkxwE7O380IysC
avIHXt4qCDoHDwtyDO124wduon+IKWntrDCG2rWk1rX2RYBqrfgdxs7KWvxTn7vDMLqbtEnbVurT
KEutP6g9LOam8hy6/4Yws3j4mRiu/NwGsaHnw9p0OJw8vGlfPw==
`protect end_protected
