--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
Hya5Lrs1K+PEdiM7gi5CNuHeR775NsEuqW7rLgwcwx/b+HD7ukNueze20ggi5xYXQW+Zd7BkCdqQ
7NYqYbMdZHS6+g7rQQRAsXNVKjzV9TTLpDpTBUgkStfFCswhkQmtdKT51vRiMeOxWWc/vQJc140U
XHJ8OzVb3P43YNLRdO56Uh4cj3YA+Qlq5VLx4xwkFkj675YNWz/CCe4rUoBs4ljUKG9K1sdlZAfH
SKKH8UVilg8R2W+GMJOMxcC15U8RLazkdnIZ8AzOs2WXL4jJVUeGOVc1/M6RDzzByozbJq/4bq2H
pS9yO6VFN7AP/oHNo7hKMwhbxvw8UJTJ7lWPbw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="lwaybHBNl42pCW8RLmL/11ArHH/mZ7FIJ0ch/QQ1gZs="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
q9xb6ZI/MMi3W29XquJTw72Z4791VDniGv0Q9TevmFYE9t8ARmQFivAh8gEqRyZPZ1oq43Aop5Rq
B1wns9JL+N1JJBEt9S3d5B+prVSHqMAI3+l72Bfpk7NImBjObHg1PpPbldZEuGRsREYiLIUaTLr8
CYGFluZTT+5BGHHiJ+pvoUekWQoGeilbJL66MECDhGhmCFHYoMIJMOe269akI0adL9u1S1CDxgFx
MR1axTEmENuVJGcSnIBqpg1M2Laai16S1vb7/YD4vDLfb0CmF7RKG/NhShnc4ppgOolO2TNgNlRS
LcMeOaFwt0ticQ4xkphBT9ciulNwSAVTIFMaQA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="nDSrTDPc0rqmMS2rndCMYyOSl/qAsKlhwtWUTTq7fhI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3264)
`protect data_block
ABh0gcscSUssXToqE9Cr9jbPnXx42qXsawIYViDFqmcDp1dzPcsVMtcc5mnMVbmznUihqBfBZbrr
sLRIiyKQRFJ0giRqb6Qmpy7aJejKQR/9aEQB5m3EtiU8KZ2Hvp7U5jPvC/tLHnbtzF6jMHVypLrN
KwOD9pl67SopQlzEMYPSSPVKjmEhWa5R6PL3nD6qU1QKU1GsMYk05RF5UEhU7LQ5fULpdqCMpgb3
+aBxc75AdhOPHtRzbMsm5PoTtw9VYow1cwoqHks2++44hi4eEd1D8GBCwLMLYco2FnqyarDL001O
SNqcDM4aw2sqrZv1VpRsaZCPpVpA4ylQc/MQPUhPIKD35naq9nHGw8ayfQgSP5gAG9UYjkJ7Efan
YWRjhORZOQOjw+oPtNAOhFawEEWk/RjYWXEKMVgp0Qd/cUWxcFrj73im3hRDKYh0UI5Ih9yWUK8I
JbbHsjk3rNrWK03zIwg4xqOySFprvqXVB+gas6maSSrvcLa43xSzT02pa2M1jeJgETU82e0wZfU9
FkpMZ5erynPTOPfyGTVgH26sKhVIUGLhgqxDCg2GtGK7sNpT9uRhas9yBKa7bSveUg3i5iWD+sRr
Qv/pSLT9XAtaV4JVH3O1GAKBhKRK30BDjB9ac66ls4BceJRenYg6QYRggQ315isnbXmeyMW7eJ/a
Bn5y8ZVKoA8R4ijYRFeL9lzWsq+ZfoVesyFVMNBRjb/ytXTrBdl9fKCdGI3ELQu6vewvx4Y4g5Ed
W5pMWgB9Hhn5HZknafVAPkgHu2UDugQS3e00PJk8mZzkEUqNy5tanY2/dJcSCX5bivCRGrSKTHPb
HRHw90Q9uHo5hAnzsomi2wQHMfwQjODMxg91Xbiovbqs6FjiLEtHf+FtBt7cbAuimMXuAsi+K4kS
LbF21KLDAUZQJAm86rsntiFguAC6kZI05BiCJfQra1f9yF/ZJfgR8taQZ2Se0/hZE7UQETIXS5GD
eBi9NcMCQE03Jo2hAt1aJPm/QESShxH5apNHlqE0RJwYGeemGsdUb6pVqZ8n8XMeCKlxU3ihfJ98
2Q6UK7uBz45iGnec7TRWA25DMbGDkb0RyuV6tyOSBfCE31e+aQ8RpqlNP4C62Rj6qfYIQ92363pE
TjHMckVVsrXdRVvoUx/HXXc/24Z8XajfhImkrVKjzVfp5oeOaSN9BCOzB7PmnFmx2WtIMCxQBLU7
+XmP9qZRvD8rVWfDYpHRkkDbgG7rwPMVZj08a1PALHxIzx8375CAsgVFdCLCWY08qjW3sRHmNn4y
ufjU2QFOxcjROzMWKw7b4igKlSubmwM3TBSkyweXIFDbqUXdcZdpCXznfDjRIWWAwBjGWIFjxNen
x9rGgXihDYMIbytIoTnRBypUEKyG8fkOmkmXtL7pB1HnuBSGESGH6gOygjNZySPgRl817Qt2v5ms
vZBhFm6lEdG+RoBHZfsyeLd4eIEyZkY4YuhG/ApZmnQGhFtn/CkL9cKkwO5Jopm9k4SEuRltya6n
wd8ycfJNehhqhxPULGjG+plw6SjTe3ROeup6Wvn6WnaQFdFDuNkoUCqZlH21ww5jB3A413f5eUKf
6HQOdk3griCyZgapu4MB9XWA1P4QvWgsAyBXUWGwo5Z1RhYyiRvv5scMhGCcSEPni43V6s9dG96N
BTZdbazdM9H+05AcM9mWUV5+xaUkqbQWGxBx5EOeqDWEkySxbyJu0YtSkqg3tFI2uSdEGQMkhQOu
EvM5BD5clB0fCWl3pAdbHjjzdAay0p3eLy5lIwr5bhDvt05BGECvQ1gkOPoU7vegOGKv/SCJ3/Iz
xsLttGVyW/Rqn021pVRoW8dFnhxMdpR+oWIDgoaewaxNQZBLllvSAgjXJURUPbbNYVB8oMAOBYZU
YLlSvQ8r1jsD+OZk7OoKy365fbZO9xzQPv8d2HfzrvK4ugTw+g2bVyoUkNSW+Lg0noOrQu6yIoAg
e+GGxj94O4ufjthf6D2ReLBUFfKVKXAN3qj3+1wj4cCPYcPdwnEdtNHwYfrUCdPpkIP2O+8Wpisw
HQU5T1k8nN/AkpMRCBRuYZL8xwBEgP6/rAD7LNH1J1CcciZ+gFtLNJIzslQ+eYkKJw4iVLPTmXO6
GS4CQyutQPCCLl/uZ3KuYqdOnWiuPAB2oQDXungJySbfO3bvcVGpsyenbxRkuDRiBQdIiWurZD49
9XbZwCWKbpMHj2qTvL+iwLBhhSM9Co4YhCQ+IZ1+Z9LOTXM5fSp+v62Zly7WIHiJMmi+C0YzsrXa
B+cWsb2pKTVdIEThrkA7Eqq9CiStLNmdqo1v2A01/Nka5cCcfBgvV/UGNfi1aDLhsO/6ODhv0Uqz
W/T3NIXIX50MQZMm2tWxtpcK0e4ZgNzSyldLOJEYiVDklKTXoQcSfPQ4t0q2K1MTsh8oFcKvOVfs
HvHS6vC0OIhBWQmpB8N/oL18QJixr5IntzlJoX2lF5oVdiQVSoYK7c8gkMOiZmd/Dnakx43HdQwZ
STmdta3t4jdrDsFYtDPHIoxuLZ9vLDYMMJWvaEiWCMIezgtBAQn/8EHLJbIpnEVPf/bV7+xdt22h
H/c9TPW881wYpucvxtD+d0py6iKz1qWVCYKV9/S5brR1HROG4OV4n4vQMvLTZGqNIHSY2pLJXkHa
oXl/hgN8AXwD3mIuKJ3I0wC9FVsJPhJmuhTzaHr3fiIL21nnr2TkCTcQ1XAx97Oey2t/OFqInrv3
fd4SRKTqbGTXnKtpL6dDfCT9ifQyA4raABjebVsJQHbfn/t//l8LIqVJkqyeMj1JfN2c7igpeVlx
CZQOJ7OaKZvVMjJ+LQflJ3fULgIoMWiSDOHUK91/1r+iZhQiyxFc+8XMf689+FebPWebQFsj61Hs
4Po0YA5fPATMYskpheJt/M2dm5ykTHnZmGui2coRgADNavIlDcXh3gnmwc7gh4VTZfPffB40tU26
37z1ajvquctZAR65r1T3a7eJTqE8sJ53rr3CemK8rHR/qIJElcZ2C9vyJLoRUFhWWVNyJL3Ev9iC
yjqCMnqbqf09Te3zYATQ3//m0dGntH9xI2XwIkTg6b8Rlg/Df0DgG41N3dkUxq47OqmphxqIuQ27
69r/eZQPBBEpxNNyQ0SGxszfKoHbau6OFI3L5tLwJNu4Imy10ecjNu9MUvf0yQmoCX7wzM2pGP6o
szEFaS2V34CPSODNfF1XjX6G+QR/CmVgTUe/UQuYHn4KTK2dPEfdFgr4pT+3hfrqj9Gjfh7RNjzw
RDG3rRDN4J9kMeUCRgpMb+CVIm6xQBZQur3TBLBwemIvJmTiJkssenA8boUxVjK1zUOJPYChvzR1
PMbg7nvABREFpVpvo/adBgCZy/MRJj03HZi+lWhv10DMmXH6RZyUUrSqNklddrut6zkLUbaMhwGF
etYk706uqjvqYpIaPrTFuKT2lGFU2gBVzGyl6Ft9cumOBjvQvfDsGJQ5R+TwX29j4WfEmL9XXzsS
S/2y5EsvaaoFi6uPrxe28mx3eZ1KWoQfNbw6Hj4GTygkVkM2L581PPHdMtj2l2cZU9URX0953FCF
9WPHmtOdBbg0SH4TA6dqfsJBVpgQHQbAbrTJmPJwrTcxhxv25Saf7z+WmIXvs/wi8wVeI6pZMXXx
Ibd9aU2Vn5WbdCCYaHf3KB8xWS5b+MgJt6R2QM/z8+oDKziC5ntlT5jk9+gMV056mRUDUCwGp2Qb
hytbjkEBAX56JlGEUj+J06nXz/BnAnHuLUUu3U6TYMsl/mVkbHwMW2H/TvOHr3wS/Up0T56tJoCB
FcMSNbqiSlsh5rzH1A1OgH0MYdavs5U/YRrpXo9REH+Q0uBSCZClu56s4GOV3WxY5MaaM7pQcqWh
A1WC7wP/rWow0R5O7ISWtUgYsoOT9UOgxzfOOUj55vYCtxWkE9OEQV0J+A8W6+vvmbeaVIfJl/Ne
jiRTxL8OLTUwmIiasm3u/hQ7IjdzCFTMpyX6IctYrfnJFRs4OADIn3at9JAhU6ajvlJO2Qt1vrhv
ddlaO2cdtNh+SIt985jareX89EJTgxpHS8YVGuzTrEKN1xqEVsb4cznT2FLNuukF1aD5kzzJL/xQ
fXvX6dPBy2Dz5nb4QuOp/B+LDs4od8GP+m0XaUBj1m3mW4BDf9MpSSF+ScRTr5fwPhEFtQ8utHmU
KEj2aciPj6mvGtxmg++Wb017m+ojFQ/GFxisSb491xtAmj0kisRp57k3jVZ81IB1bO1dCQQfpU+Q
cBoQR5BIGIQ3/4TY83klHrjWyJ4F7qse1BXWoFNBy9LN/TGjjQaSOVZXEEa9fZGXDWH5TnCjCQd9
VIsON4hQUFio1tB2GQge
`protect end_protected
