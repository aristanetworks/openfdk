--------------------------------------------------------------------------------
-- Copyright (c) 2026 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
jqkSYvenx+hCbP5tvu0aqZJ6Dgk621/CkQoakxfnYwxPT8p+7Pde/7D8CISWWcA0+8CluCdqus2f
Cy1wUVK7sIYnDrsDosniFBikVn9Md6DdPPFpTSAVHkK5N0lPT5HxPsQT/j1ulE5TK4XxGj2Fq5NV
nmg/aSIiZ1IWkLdjttWdonzwqe1bbeirSOJoblq9tXUIuYN9yBPZzba9fvtVVpaO2EaUohvvziwq
fhG1hypdOVVgCnZgJugfkFyWMcQnqRtF7eL57oYxktnBqlMixAk6dJeJhzbB7AO+1EOs4Zh4PUXC
MxXqAuQw4xZxDswHxuEDMIWQrLPdWlFHdjMI6g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="/8nCq/dMm5LxkUWy3CPnpyNWkBbB/k1FCK2qT9IpAs8="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
IAdKBH5SRn9n2BJ/llHo2ARrUiwaJ1xQ6z9ybFcZYZe+Hvtor8J59vjR5cCZfIZmNkD6iUjMXlWs
olPiKNhJNFVeyNvUJfyo0lKnYKsRZ8nja1USkpXvSuFvn9SSj8NglacV9tXkkuYe7xp5E1wsl8YG
ofhJS1Pr1uFTdHrP5VeaphrEhFo/LfvttUW9+DcJ8EBENBbayGxEEF+EVKdDPNIFg/QpBtdsPe+g
cwRHnUfuiLm50o3AdOZEqx5fCdQHsVeUzXQmb/VIxvI/NCT3WQRO9sqxBBcZVLS531Dbt6cm8PsH
RXTCrvDl+9dvASZdPkClY0Bm539XiHRdCQwnvA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="ifC37cmty5ZRzG/eXpAsxW3jnFGs5j6m13mVOHTUWJU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5040)
`protect data_block
IWRDwdG/ZRz4+y+0qhLQ8yZBv68xyfz9f6vfdU2qAoCJDCc986opkBxnxQSijOhFbelnROrlA8J3
wv/3FXmiSFDeU1DW9jDVi9Mj0DqGW4Qf33dYj0GJSFH0Zep8RfmysgAs7flpeW1tFuVKgp88rIze
PzIWOF3VyJJhP9K2+VADrKjrdnWdD86DOktDHPpaeVjVasMj/gzoxBW8sr+TTXBL91iSCB21vmf7
6ZBfb+Gx8M/IYdWlMy2ZI4z2RsYdu2fCglMa+F9C1b5jNL/Z6DmDAsbv9qDr6TFg31KL9LC7Lhnv
ZB93R23FaQWYbAfV1emuHc8HS017jqHjhNyPT50d5+Ng2i+bB2AwaCpw87maijE77B69EEqnEDtB
3cTSjRkxHi1+rNyZl0Aqas0Ho5cy/AB8X/uAASZWd+mn8WqGv4MuwrPXzA3y/RDETd9OVeowSQR5
xRReOBi/zdhQnqR9K/kZXJRgFOw63O2k/hz+eF/wz9f/vUSz2fJn+EpS+avRfsL+x+MveN6+lqVa
Khe55iRtFnC9xrEaVB1hqrWPnGMI/J+ocPvZ57AXYuylk1nA/nfO3ejPPRgiAMJz8twSfU99HjWA
i7ikCCbOBSfhhddaEdrr3Lu5NWCFxeFQW5Ko7QSlM21/lMR+AtJDoGJ3A3lTDX7x+dfR5rB2EGXI
GHC9OoNGuzIDo9FOtdEsk9gN70M7/YnzdZfDF5dK9LiMRHd4cbufAclg8v0+WQJBn6/WBUTaQ1wY
7YiHsJlEtQoqr3Y9GDWuGAWCzZCfQxCNPDD8lDqtLoNqx36E2bfyfLvCNowX/ccZff0X10lhkv+6
BJyV/FujfgUTAjqifNQe3Gw6mDzTClNfGl1jadxrOOl5LJYUkDiAyH6QDw2XJNwShPT2BBAnUV+c
8jMrcXEzxkpxjssbPKkUlMpto4km97I1lyBw895Re92yp/xVk0YOMg2WkCUUh0dkZxzk6G2k6OeZ
KD1T1Y9YX6woEIPGhptsopPba1RCKPXXbW/z170axNwIUoUQjnJ3N175rbkiNoorjwwWCzMwVHS4
I9nO7VyYC2p6pKfInMtIKq4AfmuhqreesawdiS242U3g7geELyoDzx1aoaC189dcj5QhSFsnBr5P
HqfY5Vbt34FHOW6ohsnH3PGlhAS6Hx8W2pZ6kFBoqp+xXzFRW7yM6e1iYyZ2MmW6NDfOvvtJjphg
xW0oQq5pgvkeFHqoZ7C8BMbg/ekMmtrHlPVkun7haLefjf4YuDCI3r5AJSb5f9PYirOMs5bsTj2I
EgWfGTDz7ChYXGluK938Pf0vxRvd/Z2L92/tGv62IGgUVsMjDbof9i7gjHveD2Z6SmfBSwN5eWcy
uG7lW5YaUEbWVMiDhdA+5pOImfFIj05sTJUVHQz8DI+n8KwlkAbepgC/M0+NCSUpBCoI/6w3klKb
0OPtZjCh/dHtYbsB/TBlHEthTdLptoC6+7P5fPq4/QjWlGAd1QPePNpHPWi8JatO9ezXsPsMx3fH
vy2qR7Kp90e+HArOaqxbcvn7clac5emxxC/MY8pGOfNuM8xF2KaSVDEa2NiCOWw9l2pGAtmPlEOP
9f3CVn5n8oNMS2fwrKRmEybNBRYEiRS4ow1jeaVR80YH0uYBoN2Qtn/GvahXIDvoaotqhDB8rBKC
LNgoMaoZCd6vEA9hN8LWr/R17mYF5rbP9U+U86VeLvC+JL2aSl74LxRY7beiCBwD1QD02UjE/5S4
DiitdF5G4vKz53J5LSkLR3M7jlCsAAWAflTZT417zDMNgeLlXdmnV65n0aCudQVMEN4Wo72eBK/o
0KSSZvcWwh/Ps1soBsUgekbQZUsN1ReKS3aF1E71/WzDWOoyOHYPPKeepiiZwWazV70b7nmUpwQS
FwycAXWaLAm2imVZyT/kfaR3zum0+UUDyoj+6zBq6cBHa/+r2L/YONNBO6E95xcC2T7DHB8FPsuh
K3IT2RxKVe9LBYOKZ4bUc7Up89IaawOmfpdd0PSv9oS0PjmwnYIssuETojHCCs3FGMy87wgIdVOY
x3qQN+/EG/WP4NEjBsdnwMTkdm5Faz+swbplR8gA2ju23W67e1iVC1UGxj15INhCsKja0QyzDVZ+
YQvEfHsTmonqy2MM/SBM4pXppjn0FtnTtB49Cw1MOV38dIo27j0FvGjTpyN6dQw82wcA80aaGKr5
gbU6igPycdiruh6iuouT2dlx8PuGjalPRLT4XoiUJ0gCiBT2pZFxSMZXmqktl9N7W2oKjTAbGhWa
HnaQDoCkbPtdx14uoUGQQLY+7uQUQ6Q095rr7P06JQrbOeF7yH/+Y0meLe43S3n76inRhL70DtMu
9kUS9oPDfzozpHUBw72Ue5ayAt1ZggWa6qE6odOLlE5NcHpI6docWeeV+IZVtymgUXB3FcEGrio/
/dX/qZ0WF22sVaPZkXQobcnAvnAg9w3DdcyIZAv0FD5Wn8GWpgnZXvF9i+VHDWElGQ2itMsDRbNs
s8G5BuVFHWtKawCDp+l4nJmPR43tJRjlx2msXidTlF/un2us8p/rDFCw/aSGXICt3vpGa7NF1u/u
mQKBsaB1+goux+aCyWwwn+hfmWKipAeZEUL01/LqFr7am7axcqiGlEYNqM2lNtkbIc57d2NyIigO
OHzgvEZqpx/Oz8dI6l+Tg8VR2ZrTIkS99lSJKFNxyXya/ht+jgf0yNrGZkulVgA2EvnFd6MnrDT+
Pwh45MlO96iZhl7XDmYgY6DCwNSUm28AXv9GMNOOE00Eol9GRKvXHQFJr8R0al51bTMdQLJONPfe
lUwszAlQAXsL/ayrBmjenAenAuuvj9kalw7mej0LoRoyaSjHyefOAmFNmHp1FBk0vVgpEfmYvsJ8
BFvum7uu82ADWl86ANf284JhvIErHzCMPAQpfazMUn7eBlmPHVzIG6CmDEuDj4YMseaCi03z2G5N
vXrjLeCJAc0X5PwitWQFKS/yiqyX0hAE0N9YJ/c2F9q0z8JYVNqqZh2cvJLTSk54YG87N+/dPAyP
FvLEG02n5aboUPVsE/Qjbf3opMzc3oqHWk+BvdgoR6bTHWTNXkNX8HhUYPCKeACZepn6OTJHjDug
zhHpb9TH1MKmEaKRufPdVkJbePJRrTmobFFVrGlcTKA+xrsjhgdIRO7A7+E/uwlI2TIKPo1qB/O3
ZAajGqy136pqFspzHfkuBLBvs1qvKLw19agB6Br0ttKNl451QZ6CYJ0tPiADyuW7r+UE9HLYPtEO
GmTTvQelVu0cQHqM45GTLm7nlMg7+mkKbcLzGujUUpX+NBJoMlYvkVt+uIoh+NAF508mHYDJHl0H
XCa/E4umlIeD+KPEzdN/2ZBrU0PzjkyfJuQb9oM1ueoQKW0QhhbWK2GdJSuzy8psGHo5vnk0z0qN
VPfOMOCCJH04xx/rieWZG/lBmQHNG0r+AcpN9RALkA5KQxgpdN+k/oelqnhy8BA416io5UEUhory
FmbYJep/6sAO8701qHthAJaVSCrtT2beUDR9HX36Ee2weGcJmkMQM501D5cHyFPl/GppOUrOzeGh
Vg5KSrJE4OahNRw0Yhu2YQ9tAG8MbVJynaIZLiwXtCoc+DRX+rXthNdeE+qfGpeYQ9r1ZwTp69Zx
yx9AhvPltBpoGvlhF2EQ9B2dtK8RbxpYjQLbIHHFp8vly2PUtUISEnm9zY3DRfYj8Y9y1/ADV6nC
YvcRUBqWeVQnaXN/tWNW7nP0ZUc3XAG6wJwiqodEbDt/S2rNWXQKJQ2HdXm8t2Ra5mPVHzRRIIzd
Wiz1Sgaq1iEnh3U0L+iB4ma8/6xAFqyzuFQBZNwIxyGdf8VMl8K9Oxt//5N4kBYAu9kl77m1FZi4
aW9FYseUGrLxpKffGtPEPDfv4+hBVpXKQgoMxJZ5APwdqZePzrBCGTNqLx5ebR15OcLi4J8HA36b
zFofZaDn5oGzujyqaovrdGOp4yLA0bTtH6OPxbtXQmDTU02LG2Z6ZDtzPykZi7I4n/rwVp9TTEkX
LNQj7QS6wVaPlfcSTJsV+9yROwSR8XA5sVPpJH9KDjJA0Qr3NDls9vMea4QRjzbSqiqQtRQBD1sM
St0TUf/M/H15crEeM9Pe3Ml0OtFmS+FUKqPIOXznUe3C+9mtfjscGSsJuTZ9Ur2FwjT67Qorf7vt
UIgoOgZ66bVEkfT08htYydj6e4Qubr4lU7UXMzPb9QN053RHxfIf2BE4es7g+M+Kkp8FbOpf1hjx
VDVBKTrnCKYu43BGhzEMq3QJN7PEWErtldBUtsSE+BYuw8YcrO9ImA6TxWJHUl+zW/dfqcgW7EQQ
hlac2LqjBXhMyXGdC3qm3Oth8totNUmShrAHsURObqRdfIFGtFwun5MOrCpYuCz5ON6zDRm2fibM
RScx8JqBGWf233ajQosdrHXpKZWz0CBzU0A79rqck8fiR1N3a8ET2j90SoQQ7czUK0kmDDPdS/7t
7tsXEUx5I7aSUoGIdHNpR+WlMM5VN2XEklwyXOq42ecuGyjGObJY/Dmo9DvPVErDiO+Gmuoh5ty5
sIAHX35cf9KXBW/hkeQ36V41L+xY+xLdIkXpJHgJRVAe2FyQR9XVgLd9Ciz+ogfFpzgsldAnQ8Yx
w33dfd1q2NE9y9j08UvFm6QUe0h3yjnDwT+lsvoHt+NAVzzCx6a4yXkkROQ+jnjpSzNfDMf4TOiE
HiXn8hq+g5SAeFcOSlmJ/I6G9d++I/5EUIrUBSZXIkUUjprehdjhHPVB2v4xlGZOqJUKNYpvdSOR
x9vd0s77tr2wggvu02x3N5xH6Gc1FlqsnjOpfQCq7S47bP8WUf9O1ypkP9IY1kFlJGX21vxzYo7K
Ps567q9IUAvIY/Go3kpBg3wHztz3S2sHLiOapN/z4q78SjXB1C9zCPESWZ5xS6jbUzBYDahlyqhe
N/hSp5vxVboZ6ZlwNAfD27vguI5WDqHnLtTXHcB2PM5/rz26IxmyEvEx5qArDTbus2YmAd6jHUq8
FpWMOJenaUqMmWCaBFbCbAhnxoK5m6ztTj82S1C2DWEbE6uxs3f6uTu3GhAWH+24Lu3LMTBQa/3j
WbGvKo2XXF6GIxYeYP0Oj1PPq8NUJQaGufrq01XcQKn/BVTlIwuQ/13nudGSf8/Bnt0wIKw6nZPv
F5hb1c7oSs+8Y6knUgt4Y2ZIjGNoh/2t2XTF8jwOrQ2hxlIjmAkbbOrAtdbFvi6CcPEL0SIhJ2Rl
6QT5831f6klYFFOAZdAeQ/i/jFG+A/9wUHVe61m962iZvvUIobW4qPZS5lqn2F8U5cvQ3cR42voz
lI+kV+u1lLM2/XNYeG26I4eyqEB1O6CTn/Z+V/uH1VkoChTUe4vuQ3k4xPbfaogA9ppKj4K+F02X
73Xe7dA33+Nxx6M+eJJu021xqZqnBQq+/8dO3DKsOxymTQP4BmiRP5vjPPUD422tnnstL/5yazXu
RplmtQy21mMGFkKDrdxCYLW3oReKYrAWK4ryXN3QBzY1EPF5tC9i4WpcgbhL8H6CsFyWtdQbzbZ9
i/qWY1KR14Xl34JL+PiPljUE8QZiuJsLEXrDtKeaz0h8mT8zUCoeikC3lL3BoY+B0/8WfAujYwkv
RMbBAT3797oEcbZtJVPnyeLu548o9xBh7+IgOasYI0Wdw0Fziumjlyyiia0j/uzN0+DIi92Irm+/
TrpD6rTrwBb3Z9FTzJgaivJ84LvgmU1SHchXYDWPSV1s9awnqCfdiNr+b+vQTlaljn8XVkGiswCh
te6uARvGhy0VJpzrRAKvDAC9pSJPkT0VP4AZRxdF5QdGiK2QOARYzwHvw7sIFAmjD494eUllhGhX
gy5POIIKqUTDIZ39sWt0/TQuA0QAGBTRtgXWvVOBQa02uG8tLh21NUU5v+WNYLTW8l6Qi5V10c5I
AlP+BPsS9O8Rx+pwzax2d0v+MtXFCm7ju7mxZb9O7gtpFXN10ATUdmam1A0yuLk7rzvq+eTx6VBY
ZY9v+MhJhQTxEj8TehNcqP1Hayb6x0pmk7LH/dDeYdVXt46ru7D4p8fEsXG8njlJ0I/UdULhbg7q
OewoI417SqzBVdWO+dS5+beyyrDaU47jkQsIYJY+oyEqB7ifjoW5xkEMMGzyqZBYphiaGeYU8Re7
heP5+sES0mx+3vSWbMp0VFRI6rK6+1fXkN1kEIJcnPt+rXJl5p4qIiBhRkHf2Ivn4ZbUFK9Taxso
2/LiGgpu6hIeclmddHJKf51YLCNJM2qTkjvCntF21Wsu7Go7sX08UuKXjPbPmibuNV3EQkl4GS5M
iox1Vb/4cTwbxyuLKPb3nLPbtwDNhbj3c5gkS3Rt54/OMs0S895dGEYzudjG6CJ+8OdtXAzOGrGP
Ty7UWXIH1vibI2oIwZPu0/LQGvnMk8+TyDL5O1u7/P8/79ilyZsJybZpsQk3soNR7SvohLo1OdHq
VbCqk11yhhwUbFfB4JfKzRFrdAcJSUtScMlbZlgv9qKZhJqEZmJpGb8WHOoLi8cYXtJhdk7mOT6j
2jWY3R30UKj/g8qcY7b3uXrezbJEuk03FbFy7zRQg7F47A67kRko05Y4HWZCvvNwon4i/XTGFgu1
wL7+YBEtZb2pZbyqLBnP3knG6gTka/iC2dop8SLOduzv3pWsG/zKjfh5pRY/sgaXVz8SDf1futPG
U9lldl1hTLL76QSHqreTExMDN1zjtjvD
`protect end_protected
