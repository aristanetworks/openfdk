--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
NLygA02B7Z/3eHtYTQ6eUdCrOgczK3iu/ffXVu4hI1008Vpd9GxOi0+7Oc5iP1gpDTY2DVV/gul2
EnFD5e8h5KHphpd2N87IWTG5XEV13YjIC4dO0uTOcbyMY2vE2ewiWVorGp6+g5uarF8kWi+7xmUJ
D2GyWCLpfV5fFHmc1o9pmvtIs+lDYz8fPogL9t4iWy5sxO04pKeq2/4GY49o49o8CRkXbddjv2i1
ziEYB1AEU3ZKqvOSplls0Dg8CMADKUbTzaVeszaaiVJgVFZjrCfPDYrB4TwV9rjho2XbGXyf82km
19GX15XMMx0uYBTLjF8mjs1Lgiq5FT62uhjbkA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="1Wo9CrFokvTqo3JQzrpcdy6TKHHoCNUSIJ+rnx+KSqI="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
mQ8Orgravf8ZLdE746UNStSbY+J/Pqo5sLvRlQVJfS0hiVjWP127Je8/cEmhJb+ouK1MUEL+b016
S0lJ/nUgh9dh60UM1YwDhF6GeTZOlLUOdxW1GB0x76kuZTj/EFCcylnpx9uuMYpKCvNYGeDjAXcr
fYYXWNWtLA/mdl/9ifzc5wQ9UNThf+9v4vYTaAKtsR0a7AGgho/BBQ3QF4+A9IuzOS76Lyw5W5L3
9VYohuAeZuEJ2zZlhOqiStiEI183g24CqeyGQTE9skrPgzBAqHKDxuFEV1mQ7CKArAMXcnYpuYnK
vaauenkNKIDOJKujYKHggJ/SGb7iCBluCGdmpw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Q7c/0sXnT5X35X21huFU+41RJU/5YzSyL3U2OXtMTos="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22816)
`protect data_block
09KQB2aVWSm88nxLZJ/YHeT/EMZSrp2GOO8zvQrVEg9gVxwDZoVRxj2ororgIzITNlveATqn3gZd
dmI0FKg1kVsYyQiq/Np4VH5SiK8OhTqsao+hJzBjzGIgxeEDkrZWMIf+6PiyyuS3x1qFimkllLBR
86dBHjrb9sslBIAvOuXfWRVBMfQmMeqiFc9+zHthjJwmHGXl9oPnMJrruHn9/sATywaK8lQwWIKn
dLnVa5nJDqOycxD3Es9o/32lejan1/qtGakTJJEEuEJHoPb4P0DSb5UOercWoK9H04+GoArGxEFd
Bcu2CGdj/fyZmjLGcMMhLmfyfL/SuelCGwI1jtwuq7T5Dqvqn+TgFPGWOu4m42h/xJVYsyfNKXxR
I6KFBPBI3S85lyumz60p2CaXKletiF+KzPdtVpQmBuSg6ultnKpPR1QSle5wuyZmZp8bftU8vzXk
4yEJt2FE02I2DQ6JZyBJ2iGy4wv41YGxGSHxat4LraG5uTpt7jW6RN17sENB3ZQOFj6zuKxzWrRa
26C57EgRRce7jlv1LFe7+x3frPq2EmR0grKHxe1Jdktwujxg4aIpol3TAf3oc/HqfWW7Ks9nVTq0
0E2mUndyiQJ/GmBHHhNl/HUv1aU705jyaWM6D87I20CVeZvaSSzQUQzd3NJ1VkW/gIVHxMk0XXrr
JIaGwH4dXLBYFghpHfWP2gw1IluB/tYdATwyqwr9Wyh+CWNaqAJRHHVMYlBzx213nf+rPw/e0G20
JznUZwFxqBKaXjiISTAPnkqgsXtTUaQB9KuOGsCfmx0bxVpPv6/k0Cbwpa7f23q3af3bPvoyi2vY
/utWEbu1a0O1DhiemAYwqnXzaCu7PR1W5gpksb7B832UZUoiAfeVQC3iJ/dCT7lqrF7hAJ8kz2HW
tAvkiTvMrLxOnXRBBb+r+voUSh8/TUAdA6+flv8zqQHyRpHkhhMUL+GiWvq1KuMI0/Gb/n3ddBr9
6jrP5m5XJiK9rVI9FR3hrDOxceZr3dCfWy6SFqSWYxMne+S3TbPe+JZVEvUKKfwVjgj/zSMqLWke
a6fH7zgzV5oO8OuUAR7HmbFNrxCfyx167/eEHyzzVGocE/0PFt8rjMsbyHNPVWHkUx8PoFgc9SXq
ySFBhL0l1PB7BBfHzpTvIQMWhLGbK03aaaCSa66EvfyMwJbS5FDxR5rtpZURnvUtDnYfQllpHedH
FGiURZPU7TkPsCZgtBA7ADeX5wTWmtmAWDAXmT+16Vl+lDAeKxXiug7LdkTILClWc0LkcuCe0836
7LauR+ZuG3Kwm19n4WLnv1JeY9Qxn6cm5+d277uakhF42V/O9prxqUFid2s4esIvU1m5FwTxPcjM
8feEXeODN7rK7SMFPgxquPP/lvbtx7SlFcpy7GaGBDe0tWVW6SfMZs8HMEsFmN4TkN8ngwkNXAko
n7WBNWuY4tBQOpiWYTTO4TsofCWciayBP2hUgLa3vzhe9mFHArB/2qOpKpjKKmGQLH/OjZcFvmwR
fnoO/h9ulxEn1YMBJPOr/D2XaL5e4QuzpqtCcmjheD7Ydant2at5AE6YUL3RJ1ej4fiqSd6DjZdr
swIEa2p+pYtzSJzYXyl75nZeYGNstRbKrjTj3pDOyAo3cG7qyiC278CbqDslUer1WCgUe/531PiK
ff/p71TjcMkgYjD/qx0pHdnpNCwId7loqFDHe2/zS07cQ/4j2Bqi5WVR1Mr/ehfMu34JlLyuBr8S
P7H91NeSDhhlArqXCBOEWS1xQYdCRBllPZ6Y6sqNzD5xZ/QaSAOBXW1zs6RytpPcpGHQH1OENwUB
mGM2nDGCrIuZETzd5yaLIZ6xfRXklZHNWfG2K/Gn52+++iC/cgPS+9MCBzW01O0aqoJq2zZrI4ej
bTtfpsJmKdJ8mPJXk1KrgAg8hfXJepWPpaCsdaKiAUeDwXnu0ytt7+3m0iLKBH59TjqTOC7sLHKv
CVNYSCfsARuJoOvXwD1g2VF91ssxpDssCLXJtbu8/3N7W4yJc+QL30vP6Xu1VeO+bcbywUOtF3CL
VRTPmGo/gJwW6ZbhD7F8Q/crynzt5XlA/kBJ9XALWzuV32d7Ze6VTG1M4PIX232HmNPycJWnagCI
nxJ3YY9r5pDVkKh1xKz73aXoW6n5TDSriNYqOXeqUmglOEE/qQWNl39avFrrEkm6ZHfCqCcAFYrJ
Vn5qJbIxXUM9FLsc2H01FT0ubuPHvh0+r/NrskLFEhcbfiIhTOier9AkBLumc18dNOv9X0135o62
kBz6dMkBvC+Lte6YYi0BDWTwCj4AfpNthvJ7fT3254AhXe9UyBVUg7l3zC206cL8JEsVVLiShyij
3+KHVWfFVitbAKu3p6gEk+Zpo8dld4ymoQGZZyPZCnuCkFoFym4wsqMXyQ9HwwIXnae91RRO3AxF
pzxKSoonlNfpax4UeNMPB9rB3v43/uExn9kkWNHMiNapzGvjkHHVjPhmG90Iga/JMDHHf1dR1ICC
LChDRd9gWbCn5QscS1FCiK0gbdNJTlBbF/ZLj5m9Eos65YxDuuwtKdxWNiA5TQjx3TfvbBPT+25i
86ti1WcqFjvA4F1UQNhZfQWbBkAUraqn1W1tnTW1Z+5hD1hO3lGxs/Tw6qSjq/myADvlhi48/mdE
nUuAGfpi+dCP1KNtOcJpwyvX6D3+SMDkkQxtAct8bp+ATRG4doK3GaGQ5oaoGK/veHYIimIrBTFc
+Pl6mI6yf7t+x7et8K74Grk3ODzyxxoORZVkhgf57l/usmFZ7rJZSmGNCaqqa2ApWY8T8SMBKJ6R
mCyn7MUUMr7pyhhQgoAF93MYcT8TNhjOnisIO0fHV3tRv1KEn/1l/93AjcW5WsYWoS1d+2ml7gBj
0x6Ga68ZohmCdW9XI6A80u9wYEFYGj9w78pJ2U7CsvevaO2GF/M6CeHxQhz/e5kQIc0uRua5WoZ2
TtiyOIY6Eu1ub7gKtJKJwRA+mS0rdHT0FH+0zn9eCQDhuPhm/cBV6hgMI+/H29nqo40cAYWaCYja
OG39cA42cRdKcYv5izPFBfx/SigZC+nWwwfNElDw1rqXZqOuoPD+/adm+B14HUa5HhMcJ2YZVh6v
VgWeJ31rNBQTk7rfQVW1TPvEmudf6tYbC4A814vsTNd+cMnpmi8bLRhT+xL7jCcgrQaJ+55I4fSt
X3thYGPHucWG3oW9FKjebLAQE1gWcTgKCV2XJtTCaCmSyFR7ZyptSzA3JyKKzTJ9KdwHbgQj68at
/76Y1Ybv3nlWtmNi3jUJTr5oYEd6/Uy0jpB/BGkpaN0/pbUnua3AxmyOdgmwCScSCDTnd4rA+Zm+
jhhradrwBv1aevbozuQdR/4fp/imgsjhOeyMYGIEpLwMwkouLYhmzHTL68y3UOjaShO15nMY2srg
k4I1rOjjydoVLy/vJVQJ7tYZQIR2FEjYkHirtMUdVwbh+BRinXBU6p04jwP9LL39l6L+UDvHNrX2
FD5+mbE5y66aq72WuX0M9jGcxFLA2Gn+BdIrlIsKk3yuRfaGc29G4VbNV+Gny3f+WsuUbW+yJpfK
8/xXAIN3hdse+wku580VVsddw71w/iYepkxVCXhP96m7scVXntOj2S4IquDi+frNQ6pZCWAPmywj
EGeaMfH0Yu1VC2lln3RKwk4w3eZBAjzCTIKppj4pup+IrvgsCPtGHIgeLEB2zC1dWCNo/IbrxU8R
lsiW7+6mesqopzGHUvh/QGn/BbOYWJGy2Ng1klL+9DuTtc0tQLMBWKrMeOm+jpDfcrPwVSBEhXVW
oOe4CJUjyVQyq7rAnElNQz01GqDuRbgU2cARef0B8x5NtmqlkBz7/uuUrXdCz5MjpRIKNX+90vpY
43jyuvZ3waUEbw4/XD7JQe02LT8XaPNwf35R+YE7ouQrTbZ35iWNJyUhCcnvJlWe0LIw9zAhC+Q4
7WlBBz6ynEeW2WmkbkA8cNybnqLzs7xCOMRK3jvSS111Vxu9sCFClx1D7jxFPS8FHn51cyo5kRlx
MLo09R6viec/NbhWr/W5VYVgpdKh0D9jrMGWvaIPkflEy2HLZFXk62gH+/ztGrQJSjojNedi4GTF
4U8o+IoF72g0j1rD4X1VFrnyb7BXVl+Uuh78cXUiOOCBxn1EJ2D4TEEUMpO+84FYgbAUxfKgMk6a
tS9lvbiVHbDXPfcQAQ852jpWR3xgltjFTBtl3gHoddFW2OV34mAQMgnM0m78xHM7XP1G538QVGxG
xaQBIVRrolQvlannQ4Q3H8KnDQoNAQtVjwum9neNH7r2+XU8BfbD0Ndf4x3yKrX0zRWfiqZ+0/hy
HJ0cG3qUS/glKzS2iom0HVZMjmmW+N7O9G78vVM/aWdB8lCBzEQji/35i181a/PmC5Kpm1Nm0StZ
BRVzDjX4Tdk66KIfGI6wxP3VELpaE1j/nckdxk8IRrdYsN6wExc6C3WDBvQnP8Vbms4Oe9hVopr6
7/OdYAZElb1vvahHVG34KOduXjFSgHTUX3kUIO3w0FAOFIWI6N0YZ6cWDf0XgYXmxZyf67Mb8+6R
e061Hx2twr5uR/ZHtr5sBqB5cVEC6KmRmGADzkSVLdDEPnFyd0z91T1HfAcnhV0hc7keK1B0oR8Y
pN0FUya757yKTcc/0Gl8/MIW5JVjG+DGQYstaRnGrNs93Lhnn7CzEjFIATnkLcqM7FZiJSKVn6CL
Sd9WQEJ6L30o5gIfjKpMX8U1bO1c/xxyIP5cKwDAHLXiolB2wCRwPyvfHKgnBNL1uapWDZPBwoHU
hTnZeS3vHfzqXvBPmRjVurWTv/5d4kz9U6oJWEjjHaeM/47bUzCH4fkch0U92OPVPXH8Pp0oacHY
zbJBzcnK7m1x58VD3X6UfLfWkdqtv8Eemi6+vaJqUywHHT0YKPIkaXwtKJuc7RktqF+o9yOFUXW6
cgbTYDNZEjno7zEFKUHVT740eqvAtC2RDne709RYqrObnWxyHGF1/HYrpkzx5ib9DpCETbaxI3yG
e2ydZhnSt60MZjRvk2uVQxexZ2bN28ZirXM+CaD1EA01AZRA7xpKYF9a3msY6rp2CNgNLKM6m9EW
pM49gclDIWPiW3hmSv+nb3uAFxTfyXVn3CwayBTppqsBonwDZruLShoErRIoaQT37SyjgjXnzoQK
rb5IjLlVibZqL/4RsCf1Y2BVhEEV9EPCa4n+9WJ4nVJavrAMLUB5Z0+W8TOZUTLP3K6VwJsYfA6t
G1dB33BvmWv01XEWAIowHHY00cbZeatPZb6A33J2Wu8HG89edY8P1YovHrG5cTr4u6FOa7C55KWs
hxNuGtfHn7cvc9uc2Sci12kgw1cebmmUVlLjKLZaPxAJ3xzyaglj2mE+FcS2aaVyEtq7HcyE6N33
MSrB1aVIlONQPkHyO7xXQfgllFq8rF3GA/3JTkZ1DOEqD+n+F3rBXF4vv7BnoQTI4Okz54tloR8Q
Mf5p6yFBfr9RLoy88cMmWGtO4nc3cB4Kzxse/2qr0giJ6e9j7hqgRh7IlKKNmBy4Wb3GWQQHOrCh
p0270qBknNiiTmfV59sqwHDoTB1C/ywvKaUox5MIkYSfbqlgIufR7mgSz0wp/m+QmKy3lTVbjlPo
FX0mjk2PZ5MKHMKaRjF8Cf48Yc7XSbIGT3hXGQ5hO5sqnOIOG16Gt0df4475sbBOxJq/0bPOAFxo
tG6fw+9EbsInC0z+IT4PPPZeqtpW805c8PxLo4rF2jQCdSEbPUZ4dTELpktwOAwacxNKpBBzfsza
fe5n7iyZB5LkYIK/Q1aqaW63xRCsW8uiyixf3MULCIcSIxnV4L1tOwUFaOwm0o2MAK6bLrV4jQGv
IrIMioowPdn4Wtdh5Av1BFv76wZ0WwNEz1XSqKcWVY321HIL7lDGia35gaHTJ03Dh3lWOcbg8udu
PEo8sjC+U8Gri19PWn6+1WH/NuW/oPGTKeRcvD3LiPpHy4mXqtbGLsu9zuDInwJTQiMpoGeEirF0
B3CnJUc9lz1B1fwoUP14Wmssq6uw42ASwm9gh+sNEskHy9uY3VYRM9PZ9rLNgAJRlasfFYkZSjjx
us7Yx2ngOs4uSao5XKfYmO4Q4wKgjbfcCOwqY8FeK0ncUC8rc+l+Uokf2zRHMQrbtpWP0GW6ZUlL
+ytBFWRrWrN4Q0UgEsGxYJ7hU85XZ4XjYQ/0dk0R9oAXnCY4kVofyTiAouy9RbumUOKTLWRULr07
7mP/+7+42jSYcxEg4EdIzGthL91lgYoV7mRkih7O/Eg/1E2G6kxTAZgVEKK2I1TiIJn5EDcbxzv0
ap3Oet+/PorMmb4ImixIiF1UJUQ1XpitT3YM8qPCR+IwvgjBWezCDYgH+q3wlOz78gKtFyvuJK6y
sjA0PTUXVkmFkjXrIsTqTyuryuetjS+MWuk6aEIzWvvEp2UPMAS2ZcIgP5IzMcd8/fxLcirIFXeD
DDBYo2kBeT1zznEcT2qUE8H8GOE3Gw3nSOrwJicVEpo1tuMmh/DEDORjEVGJreDNsGE1AnC9m7cB
hkYmWjkuM1k4HVQh4ulIl6cJgvZJdzBrk97j6JwtBI7Y9y+PhDcNSC++xlO+sw0pXorEpLJ8SWv9
zNttSoAAJ9dS1rmyi+09Mn1vqL9TA9McnqgREcok/Mv114fC1K2Qb1cYhNmK/UInxhyG5pzTDKRJ
VtAZZ+PaVgAoCGHmfzfI0LOWfQjgkM/BrdOviKtZ5bmBuPl+ieCcsWzvjAsx1S1Zo6KJepGC+GEL
5CDNF+FovQRZ+oGb7BnrnL65AnqlYiyduISM2I0nOmPTjbz3gXK+smaI3DuXoPsp0nIfMz4dnl5G
+bH393RB4EejOoKy8pENDf97Jr674/tu0/U0A3VaK1xHGnL1w/IbvCN5aLbtxQlT8WkS3kZGK43n
GqJlcknyEpeqdS3ldY5HlCwNQFXTnDvIC3SRlMNFi+vly62Mj7m2jxm4nB37fd0G0kSdsyzS7oZX
3uBxKPOPLSE7MtBLZ/WVujypqtMZSL5FecHPhVAKRw3K9vx+f5l+GaXpDGDjwtUk3SoGw1bkwdEX
mpSH/xEE+oZyrLRRusIQibF9qce/unXzP1rh4taWI8em3yVL66A/I8vlVUQBi/lEieBR/RsoS4kA
10Y8dGXM49gOazshQdSbt/3mNENZztTY1rrNW0eoUw35FFCQtIefbfx4GTLS2hKU+iOl46VrGWKU
jHprIx1LcMd0KE6DdyQJxDhXITNpAU3vHukVyEoWsvWEHx4znpUxDw82j0Si3VW8R9SxAauZOkY+
49n+JHUKwLBPOrl1A3uNdp1Kr8fjwj2+6HMq3swVd98TYUUCJaOpjeBxA2aNYUIqa7Cyh4WGOr3/
pSeFqDdYs1t0PF9PR5UuuDSSVkcpApQIrOD9O7EbXq127e+dnHG5VIyYsorusdEkTge6Sy4JYSXM
a6qholytSm6Gx4Wruu6stx1yB2l008RAgkn9d+Auor3u+a+A3uMcYRXaUG4pLwDSesrt+XhpZERn
FeNyjeYoVbKwR5F8yLYKJXsLJ8yr2kDrP7QjYgS5sp89A/aUY2pXwRY8z3jUSCK6R/GYjmiMDVD/
JVA5Ui4OGl9mQcwrmLQBgtAOsoEFCeAWGzz+xKNVKhRxwJ4NHwlmPINC2fHj9eQXCXrdW5CIN0X1
8LBxmfyt4liwBYCqamhW7tdJDHkJte4uWtS6qmHulQRq1JVmP71xZxfwuY2qj/nQw2DPSDCEm8my
NKpu8aoMsJGASj7bqhe8ohSb02ZOaFfZqlPZY9EQZ6jwuiLglh9soekW+7rzOjk3feX0fUFkuiLm
fd2tCe4gBq93bMJ1pi2/+iSeKWf97oIcreQ+Tnq3zTajgoOz+sOrXFCc4BEZztb95nWp4/jh26O1
ZVOkBr4N+dXc1T6yr5jjqU6I6qnpTyfLNP3qbkgP8zURSWmmgwQTp8DeC6RyiviS9CUOmgAA751K
XQgPNRkasxeqpoQJHLNFwXzIdmoaxmESMktJETEk3Eeu1vCoF1JBJJrjFZBzg1df82JO2kDnduEo
goSEVfjH+VNT8gtdAUNO9hQGoDp7a5L4GghoFTfXP+lUZd9NOWw78tFqCjmQY/ICLhodsgxqMS7P
7OIbfWOuPGv0Rf6r3OA+WE34XuZ/Ec3ceIqUQ408KSqc0Aiia8fFHcjDClxBfuuvk++ZmPHcIVkC
FH8eetWTqqrdUZtaQQ5TXGyh3H5xD0Y2rH/gYiSdSO2v6BykFpnDQj9dX1XYxedALds3E3bthbEF
lY/JjqrgftaaCp0JT3l7ctwBczJuyCeuQhs82pVXhcl9aVfF30Pn32rYOyzn/UHK412iXKFzqw9Z
tLeuBJnD5OozkzxBz7emmXt9/urvl7EjuYGjv5uGaIHwQXpCp7lAu15rlasGR/ApyueiLLt6KtAD
NTMUohM/uCs7Cm2JaaH2I+7/g0dkKq/sVS2MS3/QrRxBMB11AsUpJVqIjQL8ejavNpVNgSFFDp6Z
9SJTOfp8RTGJIWtNAu3i3fMfGHYtahBlk7NIrBVAa5ndjsgqp2qpIjGTcOFifHHf1bJsnWaB7AEZ
EDBhEtYt1Asg9LdYLDPea/x7VyTKevfPistoE6Cso5sajNmr+jj/snwZXjRTRVzDWCxcOW1FCNi9
nwKm8ghIP5cAJd+sd9fp47TDZzE+QhEtGuLVD3QeDsN/gA0efX3jBMUpp76+Z+lR/3+n1zjOH2K7
qODG9S4ZRiTxmQEluD3aCPyJ230R5tWeO4UCtll70AZHxnfBPbsV0UjSsl/SVzFi+BBZ9myPro8Y
dRFwoA76gy6sWoh4u36G2iNSWOrwN4mh4ehTEDBGfa/6ebbah9AdKd+mPm1MYlTKPce5VZDC9hF4
2Ec95f2gwp9XG29pW+yosNmCZsNo5850jH+OyWE72voG5kbF6O03s4CieAn9nbfozBPEy+/ZpA2D
A1yUXTjdqn19xRZsxcfJa/Nfd3eXIns7REYB1hMVWFRHuf9c0eeMRoXMUD6g7x4s7MJby3lPqlcl
qhIHCLWYv80Dlh1gQ0ee+CRpA821tqIt4SPwfOmrYy5Xuxklmwb7zIcI8ZjG+zyxS7RwqOFhy/aj
J2//Jp1qI7yTPTnKEbt4yoYiA/5nBB8B1IIyLPFQ7NOv7oDKYJ88Q0ADgcMFHsguwNDBFAJYe02A
JNTwZOCR5xPR6iJ6OybjgxMEkCIPGCPDsrgF/vzlfU7/jzSyr6o6o3Xx9yP/tj+1Re3yq6+upQd4
l1p90urNs37pLKwi2DSFgSQgQctiIdf68f45i5EDK4qF19hnGexNUErmjxltgvA/J2QmLeyOjVjj
1gaQZSqgWHWRNgGt2ypVEQhrtac0FvJoPuOClgI+OS3mJ4bh8yDs14BnHDv4u+MQfpnnFz1eOm9r
Q2K2zgHKGGVCg4qGmcdKZgtkc7eLzhIZOl6FfISRa/VSYG/enbiw+YtT8+JjNnn0mjAoq8nwp1XO
cob8fU6rH9+kDNafsH0z17dWGUcKMtFXcWsRQ0q3+7BV5iJMqNwULQjriaEpafvEdFyTqHh21tbI
glyGB1CZ14V3rILLw2qag9c7TfrxKP0/luAm7Rr/WZFkn/RYLiVzdDJoWUmjZZih5qdR29pGywZv
X7Nrs0eOGe2MQhXYU6CAAeI4skmQq9nq/078LZdmm1a8Hm2LYGYI7LhpXEwio7kBB+BtuIlqTNzY
oiPQyCRxUj+o+xrYWydtPJ6d02oP/m69FoS9UFLaGPfhMbDclY9R0NoDiGzBZtcQHbohTZwM8Oos
sLTjcPwDgnJNISPHz3X4Rz7NVhxD5JhhMT0LqefkF2FSwnvBXKkw58T1EBqroGMiCusY4g/Nhvpc
AsOt7JCCK4HGeP4pogFMPIqlMrXM/CFVDTLAiHj/WG5DouezN07vsWK3TTFFvCnOXnexRNaEL2rA
FcOpS2GTDj1uXzT0F66muZMgGDLRAf/+/Myw5SAcMIDiXuZJJg6CQBXd+u4d68stdfQq6vh4YT/L
/hsz3hq1jwQ7P7v+1sPQIZxrnlI6i9V+gF04btUAzH9VI4KGd45xpVAWKt8/jlE8FWiYVwbtzeM9
NcCM2yLYVANEu/oc0W8MzxuC/FpxsRxwONlfd6G8zTlRzyvNHKZfA15ZbHPZgSzLvYYuJDbH1OXf
PksXHuydWvV1y2Ab2Ksc8C//zfoGNIQbz4AjvtxMVf13GgCZ4kHE9ooQ53zjHgiMnsvNgoj3MUOz
kLqs2mi8Vb3g+Zvnb2CFcV5T84wq8P5iNj6JnNiK3sw7uYPD7h0OARyepJO6CAIukWcQFr9oJf1A
9v7JxSxckIDPrPjpVoSVohVqaF3ghchtlaDovMl0hIu0QtFzP7yQ1HcO76aDHcLsdlI+hL4viTsA
SuSNJw5Tl0vYzemvlN07Uz3ZFNwyxIRfRN22YpevSJewV9G6cRoVGu8cBn05kmR7COOsjgFZ8kL7
9BSjoct04OCptiV3ReYCxZjhr53wF63vtLywlqvQ1P69tw2PKplRgm53XZeSMGqibKfjF513P5YU
8Jb0vgAHvPGxGMo5IKapv7Ay97aHymozr62rtwzmpBFiYB2pGK56OcUOrB93+YQnVYUGPK65eheh
6cEwh5ve0Wws/WdCl6oFG2KfdnjnGvkiFh/8Z0rrvxvt2+silnt/NS8NuuemsyD7CL3nvukWSI3m
PLauvIm6lDWyv5S+bVmU/W2NA6gpW+8ibdJDQoxf4zfM9fLhbyAwvYRCN7Ol6poM1U+myPTSY/m1
dVWQoB0oYNi0MhxJ2jYUEcG606dWqCxqa3oFUFcy5QsE4FjSjmpyDq1Ai9AIgu6UZQOpWT9iib92
UTC3EdnQlRXAQBHYXO6IE9puMVmkVRw7bkFZnGpGOJpzL3sIAjKzmVauBHQpUVZDrFNYf2fLUZ8D
389WK2GirH/VjGvQLjHkSLaEZfR8opmRhWbsgbwTUFaJtZOY1Hm3m8x5INVpTgdn9NOqiMUdwP0E
oV8sVIxsMPq+9RJ0UyjAuAUboGHz3819AuoiSFD5HEX27qacHTr8pSdLo76eDak7ASmuUxoSjeB8
uRNK5ORVAwYP1a8RQ3TBu/2U/J/s685mux6mrNGSBKO1Pbqctuph2Pbktn8Fwy/EK2Fk2L9KJN9K
X/DsqgM3RnRI1pzzFDZdTNQEmP1bG483myjDMBnIxaWBLEFic7qYo6s6lRc5wSGGt+QjYGWquSuT
1KldHyhwEYIBETHgoR6RKfgRw47ZTTaJTFDGO2NVgchnxHxp8OaeMWonDH7DUmyuheSHqnTiKG9g
lI++LSAl6/c7Bfj0vN3fwSyBv7ASXtTAGU+ekXG7IqndwhTnd6gl4mUeJCUeglUSG9cO6V/BbFVX
Xhj7x98S8BsZNcrOy6JPieJY20h+gYLdCsuDo7GQIxdSJXucrAbemCGdn2z4ElmmNGomS/aQPYH+
WFeq9dFF3xpSlB5zqM3+kSWtmj9LSwgL9vUJ2gAnqp/YmoQLvEhBS+1Me1SxVcbCU5DMaH/kzHHs
4fJtJpkelp8xIcpIchBX+/KI1u2EcZUh0mNL6jYLe5FEDXBm49QrCwIp/MOUWe2anVnZm2Q79wPB
ZQAAqp+Gmw2TdyaroHs7FYfGGBUqAv4H6uFFTDBF5O4zNkCLe4NZ5B+CuRHtd30dwCemt6SU9pw7
v4l7NqcWAlDNcr8kBEuWzgFiTNPeH8gP0DqEsRgiVlEBlNauaaNP2xmgam2xpwnYuXNoNSzPcv31
ilEZkSo15a4hct6jdgSrnSm3ruu7SiJpYar0LMPJ+TiD8PSvDLZt72bxgWrz+GfNsWIDYqXAGjqz
BG4QeimnivY4950/v1E7vmyKgIfa1h554uvC+w62T7DJmgxgrwpcu71l0rbfsYhbB4a70DqHUKEG
Cy/IXxeMLCZpHvKeTZdgs7QoxpWOjBG7CiNjHBINa9DXDmSI28deToah+rjBA208j+X7nT0LcdiT
t54jzVTtRTswDyUBIv5mMKFPw/k1fbsyTmhbroiv8WnryYaziyzBgA21aRbBGSmYUWspXrvy5SBQ
tRLuhdcTrTe3OhZ3u4RpIhtP0aRAGtaDXlb6xFPS6OM7pt6thWd4z9I6TSo4MygNzU5LMiGdp23E
gGTQmc/sFVhctF1trn5A+/nO1ODHoou+lPePPiPpTFsenpgwb4EeyRbEKUCUa54TZwmyerQZVmtK
O3AolbKR1JBpu3+X91W7GxNLgJoUY0HVZBtmy8oCp3SyicgZsYeaZZ/f1MGA8wcuMnEztkoDucpS
03Pxn9lCSuMkk+hq1MEISKmagGVTnRnYc8Q7ZUbtezEEXo2niLefUMbX+xdQQ7VngeBg+CWesW5o
3dsukqbpzkHGnLvh9uLNmz4mZALxDstwdoXFkj/h6Fy+SZoNEVanHO/48EUkAnbaCTNi9fsUzxdT
CJsVr1+pJJTQK84hJIhIFGyI2CcqTOUPShfZA+/hWGClcQwhXAcCAw/9ANYDbCs9ev7NUtOjvxiH
oLCvudRdJOwTJ5Xgh2XadRxrwG//WZPr7+vKz7oByx4u9hzwny/xk0lDsqHbCpxl2JAtmiLWmtcc
31DEKrAhuJZBWh3Ewd8reGPUChmoK62GBbn0ULf0mNAkVVFs9KTLXNJxukThhmWrSrEU59DfpUOY
YsS4hLX1LaTQ0minjBlgzU+fQr+Eh2Yi3yb5nAEw4L3OP0LEJYWQdAOfZjqH0aGwx5VTfotqq6l+
diCmgnHbjG66/3QqJSFLu4CuytNdSbIsh44fntMMX+64fhVgdByRSjxG7sCt+R2ximxtcJZkLELM
WT+iwBmmD8R4koQDcJ/iB8K1gcxKznpG1bwrX4X4mhxoSiyYqefGA+2qWjBX3NTwXj/ImCioidA8
19Op+SOUh1glTdjm7WqvctJXJBOrT3fKuulnzy7lGHkIM+yT5Tcq3rZsXBki3JlcYa6TC5nhTXzg
uCojsoP4IY0+Ihy/z+uI9IX+nA1/cqp+6ESXfQlV7z7UoYTbklrqv8zVGbpD7/VRUZo0j5+1FWS7
1t6vEal3KSptAsRKwc2vhZsCtEK2dRkmNgHh5GiIpBBfspAS7OItEsEmwN7bXFf98Mqd8SYyy3Ov
lQodOE0xoPRbeg1yUOJ3Zr0Lp3SAFs70dUUMIqwxrUD97Eb8L3olo+3HC/QhVBTy3t1yj1GpX+qJ
k0sA3x7vJEjgFvdTJ52kGTfVhilZ5TUjR3A+GxOKmdbb7qzl7bFmc+fK0PZcIaw3CwIEp+q/r0D2
Cusw1eDZAU4FZJA71TwezOXC5z0SO8r9bpmSDo1l4hJbrC9/GhHeqXWzqM3Ni3zX0t/yqc84ScCz
P0x4YlkWPiyFgFMn2kmmPuCGesgwtXcsu4ZpIxXWqaWQoarOWENkwFSZiCWrWLc0qetyPyrr8yaS
a4iWvBAuZ79XSt+TuzR+LF5Rl50Qq2ObQwXBDsfbCHLry+hoTC9qL7eZVwfHAby2q5uOt7TTWMzY
QYFyEDsEQnPqCXZqcDYRZ1Wog8h1M/jHY4APOItHFmBr/9I4opsslY89Qcz0GaiRVgRWWk35tDZU
Cmcb8zoZukNjcSjqOKkmq/JCyNDfOsFrQBDccMpxnD26Z7v1arADo3AglufPp33Al05YFjhubRaV
DDaV1pT6DHYnonuTlOwwiPoW476ncVE1lOxrIjF0KUvxFLV02RhBVd7bLK+9jMMa/Dbcf5p7PXAP
24eryFM8rcpiv9CY+NKTpdFTvejmy2LArzATI4TjXzgQRPuiS5G2lNuhMBqWhDNQbKrmKUh+vvHT
og1rnma7dFIa12QDwOVaL6l8UWpK3QC4XIjW31l5sK8TsXgvXkyrVGnga0Fymp+76t1dQhb1YFsl
kG2VpdiXYTUaUEQfFkZZn/hQlOgToWs0l8AeujnCTTx92TOXN00ahYGxWUqfe8oZY8JjSM0o+/zj
eGQnAl9FJvPSMaXtKMpU6HA8H0xQbRfQ+s4GK1Vu1kK5aUB2pAl3R9MbKYS2e7EOgpq5nZIVv8D1
FLvhKtjREBlelqpgapy7RbvxbmWA/5WR3K4wEWYNz/AvNfKnyR4MkXy9ku9oum1byyTA+0ZEmuqr
OXJ/GlITi5uoIpfeqGAQojavcctaTaCAUMS01OadRv3wIwqO1ia5jaEVF6JrCbi3GLzyDY8slTW0
aMiNDH93kvdB4sXV707SN/2OLE9iZTHpi5j3e10KZ3lXc3NQ1/5JKYt9cemcKoD0s13Tf9EWNxs3
4JZuX0iLwkcemKCjKPHpeDp0na96tKgsumz2gcmDOfjPUeKgxGW7m8uMXBDWIjwuUYJILdRKXnWs
4f1kCZIK2SCg+qkDPAh4woQEPoRIVBqTUBfE5U/txBRqVrHtwx/li6j+KqBZzMU99wqB5RwtkwKy
iEBhWWSMt3oVuU5Fp31IYRVtdE4otDLb16iCfSJ16vTqneMiUugsDvQDPGcCrlYNu0XaZWvNaIdd
u7UyAU8CJoUrDpD4orQ2KaIUKe51qGzIDyTGrRMr44GQo3MxrV17ulXLlODFyz0y51iZdyi7X0kY
8V+xqa8UuVx16qDLogT+mGm5SJZoodl3UauMbTmd8TEirTbFYoNHPhgtzJfxlMqlcpnyCLga8i2+
TF6VrHwC3LnK3WWtSRkttW1F4+y8KCRRnWiZdtOCMhqvUEknOP+BE2iad/2RwUduXWTzFM/EaDzP
7goKzC9tYrE85EWDN+DZxQrkDvEa2nEo7UmVHMFoKMI4o4ssDvyC9VFSuXlbYq9ErKT2y4ISPxWC
w8f+JUe0RyK/t1WJaUwXG3ub1jf8ZsY8sH0SaBqZ84toq+FiSC2koYMIghOuoQepdCvkzoBJ30GV
FunpHJXCx96lBEVEWLZqhIEPp+UeVN3xl6Syzq1hCuBwIACBNgyA7oDkLQ9YdvKnEG5D3U7epPQD
lRPHIQyve35YE3PJIB4S/m7VSnQSAWP6/682w9XJo7T2T9dPAT8qXhXvT2g62JlVy+1jmqB5/Q6v
k0Qh9uKn7d/C78zRIJOC2Cp0fyxPLUYuFr1liVwk8otBHoAtimJQKbJn/MWsQYXzIjrDtFKTyrOQ
Df0Itmzrkh77vSROvnQRvKrjf3hZALRiZug/JAEEUys0+w0qSF+K1M97GTObGt0sXDfojqufcWV4
paMTmDoHP2A8Qs6ydX0DWtr9Z1sYf9dBjPQLjxlPyqqdqZgsLsFImSWymxSmnnUViJGT2L+env1v
/hOspV2xiNKMfUSZA9LO3oZm4mKm/I5sm55xvpw3niHJOoiZwznE2vRSMe02OeYnRqyACNc2e6fo
SqHt0zgzPvrBAbNKP85VZVFDHaZ2t0FHxxTqKsa53Nle4/MHDHHgxuGQqwgSNSLDhLLJqXHwCii/
6xvuWJd35wmvCIAFOGMFHubXtorj6sV0+d5al8uZ89fmNxX7i2TKc6z/b8xssoVnvZZrn0tzfBlH
yGpmU0+0CfFfzH4HefdZpLcTeTzS/HzR6wFIqacgRNov3hoqgjiPVVzl4AXjpeD5GO5PWImiBlHU
mln8EAHOOq4iwbl83OHF+l6P/jNe8b0SidZsKc6QJMWBBH/S9iV4emCXAHXeNdfeqyKeGx/t9STD
YM/SMjBPbzuDxstTFt6Cm5psrrW/SbfyeDAlSfoNX7A9TH01pkrKpzh7MMevdIbWUmZ5xfuflHjr
BMS1PbFPKK0u6eGDmxNmYQDP0RuH9DHXlVycsDX2LOOvOPeskQiJtcNgLSBWl1CF8H8Jjdn1+XGl
8eAatN818EHpTmCCz1HPGhHSXEZxPzhFaROnSEVbHI12O8NroeyfDE+HQo24349avXHlgUKPvPGs
nWbkiNNR6YJylIxuwzWt5V5jOgONdlsWSFqXXWTa4ts/2Fg354s3hAQVSkVN9N0/Rq/321DBpx7+
yMXhK958lduqTFZjbDyelhZ/Ib3x25rbnQbHBr40ztsK6co8hmq3Nefnwbc46nfPSxtpqKw1I0P7
3LsoSKqRhqWxI6Tc2TsJJQ9CmFkD/JvHDvGP4rFZv1yWAUdvwSSF+NWbTSKGgB1fCBxgrWtsoTN+
5ctMI0heYawF/zqpUvWE/raKgcvW/NRyi8gUxButi9IgMWCUwdMO2HTA421GjxDbBKWQaDgI1YpF
aN6QJ7hIliMAD8hVgcIXVe1MNBGrF+hs1IZUyCeFQoyD7LUK9E5B4gJ8SqpwEhhbpH8dqVZy016p
eKFfDqnCCHo5aTFoTkeTOJ/HbI6Fsm4pwHWKGhxagn3UpnYu0IAy6jLlAwu0+5s2AS18p7NEkFwT
U7P+ayIVkvajvkxTh4QShZV+9X7P7qYNUqwsmqdLcy67KT5nZ+ObASBS5T68kNdDiMoFbe6FMikC
PW52O8POCumw1XLb6MBBm2a7kKVvselmuX0UP7c59J1tKMOzSabTIg+NtmfK/6r8f/HOTGN8akVn
hJDxZ8sXGz/rsCRgVomBZfmGRFvBmqVbCiMFfAWHBf4YdH8z5PjFK2O1RicurVUb+iLi/KLNWhXP
HmvIopvSXCAjtgmYH4LOe4efKI0lqLgb8Aiso0dyp7QEVzoM8H2IKfnTy7/H1ALex6aHElzY1TuX
eOn0JcOKHxVGo13Djz41//NPJJqqqnsRFD6PHF2SxRorOrgYbsNRcev5cdRv+ovgitftrlyoSUxk
Rfzjcds+Nz9W8u2JkmTQZ4AqsGlAstCc1Z9I39k1f766mg4jW6jHVvq6vx/KF1+ZupkkF3+Yg4lV
ulYFP4OMqDAgGBOeFwlUW6UaaMt1emHcSl0xwFCaAhfc8DczYP7XyzLaRUhDEzUBD1R3ChHG/zrf
4N2blQ0pGSmlOU/FY96YX8nVdLrREA94mfEX4BIt0+t2EH50SwIc2DBvNBDAtX5O/nk/7KITpPYl
LWb9kbJnjJtDAsy06wxH2d5fQo36AeMm0oRl5aiCi4jcwJKcVRccUZJdZ4mr1TbFQtizBFhFYUtP
O614x3s+IxRm0dfPAEKNStvnD5fea03YyXa0mevCXLSxK8UNyMpjZ5Qwh2HWZm1VoytQL/EHQRhW
riaLlhrqzjReBJS6XkDqMRkEpNTynhQr3jd+ilzpQf9CCk8eZU0LTWuJB+Y8xV3rjCThfn0SaFAU
OE//N6NSiB3cq0qScja+7atxzQA42CVVFLw4+OLjn+RsuJjjpzhQRYN0umas4SaiqLPPJ6K4EpaV
1hJBnLT8wtzDPWykwMFSoy1FmqCSzvetnfukVEkXugF/KxcQRwhKvmRX8EIpc5AK9YEVVDjTzeOC
0Qmo9RB+jVPPNLQbNvSPlYxOR5/NOQymPNegckjY32V+5xgK5yLHS0zFHL3ELnyA0IWOCkKi1vZB
wdTNmBa6JOrY9birrQJ0oMWn+VKn/9mV6YsfK/XxCJICwUuj/rkBx9zGMiJAWWdDhAIaIkzkme0y
b0dr/JZqyz5hZXz4hnjtB1PoY4eDTLLZZ1GYTOachVI+NlQ74df1ftsRKuUBw1oXz0D7ytejta9s
I6sZN0JvxnLySuPnwxSScn5UE6LqkhP2bkV89+IkjFNz96zqd8d1XWKz4gH6+7o+5SgbInJPJXEj
ZXFWwEzQyuGHe0taZ9f/VcN4RdELVfIG7RhqIHOrYF0lO2+DI1rCyzwoHCbxGT0TMgFt6kxroNUF
cLeKwo8zy2pUmLDuJk9oeKnjhLeG+t6iKOnuo4CaHsToLbRJWbFA8G9WkjQhDOuwBPCuZiycqFpI
WB0z5ao4pglKJEu0908bBFyv3q4gaWGSsca1vGKsQ1jYZAUsLKq7K+s5cHplfDvpPHbjtNMeX5IU
/6jVkCkhIdyQJ+1H3ETjhbQurihgJezURkNepNO4ONZuKumv/21YFcZN4ivXs+oxAE7FW3JRSWI/
jKy2zv94WRpoELYzMt/IuN4kDZ55b2PyqvZLf5HX9NSZwnUQMpXkPRmquMXCJN5OO3ygpaHt84Lp
LVno652mU7+uW6OsIfAaPKSPOswTJJjzPFUpp/Ft8nxUNSgRIk7YY7guEehyQKku2x4ffUdw5F5D
mMUNRGFMmCfmIea8fEz6vH7noxoCbrLvoaQ/R19Bz1c56y+faAyhUG5UAijzriCXA83o4v5AtmF6
j3RnlFM5c9uMplde2GuryAxtqvBKNR53YVhp0QNydqGNI1uXXAoBudCAqsZ3L5yP32kL1+fPvrB7
pkceD1GFJP5BMiXtumhZ472Wt58VQuQ7jZYb49xAV+NWj4PknvYLX18TIMfBArwa9qyP8fagxSqe
tfk/WEHcwd+zvu8hHkHft43glANpGg4fm9vNRni/YTkNYru8MsYIvLmqvCLMbqJFVzDofbpULULS
qHQfOQ5BP6xILOgNlzdXhhFr9vf49geii+cbdx1LVbSBHu+vPuYcKEpPCwK2bnd9uAf0oIIN9uji
sORkyShCQGXxBOdPrTsY2v78uudKtShrut09NnOhNwWRvwjtoIABUeauRLiFfBHjAc1U68jdg9lX
y6Zm2wyZS+RPgX9+rrx9qfs00pitkXHxMc3pYVVivJs5npvZ2BfgodddTy8aXyxTD23EDHTyP3fX
j5DzcChwZOOj4MJOLqYqcClsKkFC3DPSfTdcni+BJ36CZM6XMMur2O6gB+MH15K9x/KQU2CwGC4C
YMGaSVEhzBuP2HTJ4MNQLvXUoldssx/3+6x5XIIOEpL4+OSYr6xIPde7spBqtF2dojr0XkGZ0cFV
Dr5pXpKxbvhom4Cdn2kn+akJ0Y/C7ztoxxt+fJRkbqov+5KhWfCaTnzugET7NFD9S2TqCBlNhaQX
upIW8wSyVCB1AGnPqwf+Vq2fbU50YIvsCdXtd3XCKFpJwO6zYUsNILHUABKp+puJkgNyGkZRv65y
c6bI94CaQcXMdFsjiOsVsc/j/iFy32tGuN/PYTKc2u7SJw9GnoALAUfrXfpHbBAmNjBvJBBG2Cbr
S+LRVXMYqy3+0FFVtyR5jXm1rKjZYVrw+Uw8cFE8xVG+YcZtdGQ+L1JPGcKzsTfG4TbgbGrUxyXo
7V4Rx8SO7vjO42QZGGAzCAI972agRpaBVQa+GmHz6nYDvdWAov8JqXqPmlKeC4qs9kN9DA+Mvn+x
raucfJXGeg8BgJaxKQaav2o0YvLDG3aj6Z1RFpWjVx35+r5HBxOTQtB+S23/SpBYYDva837STtoV
xcAdRAYP+ZZXtq/w8lvSly94bHpZQMoy6ez2+cVKgvlZFQBCHYBahHESHdyCnPdVCwALLhf3CKW8
zNrKB/QdyCuGoqVX5FI3JBitLPBlMg6aomT96V7V9c7wV4iWuCHD8g7POJ+YG9zmWI9A0g6rWbWk
T1tf7xu48ywAwNmZ6l24xdisI238a+0b+PlZpnm0dghIJ5zX15ocqg/In1FdzydyX8nb9RpvufhK
3DI9zhzDjhrHFiZffFxJH+npSiICKh2UMntb0V82bZo96xdcWaPut8qRpx1A2mxfn4Wj8GxNhzqR
MXkTujyIba44T8mb1fcVwVmXY4VeVTv+li1Yq+KmLmUuZhADeOf76b27PIipCSU92dfGf4OVLIwu
Uo9sNeiwoLZHysHCd4lFrxryAF4nmH/P3kuD3n0CgPwl92mJtyIWGA6A9lhiJoG01zvFfNMLEP+2
tn2D771j79HjnIXzqGGGcpxXZp/Hy5U6IJP/TbjSfWlK1dtLi+KVQjTUg5w0TRyYAEoYlgAo3H+a
QFJFtunlyRt8ue/3rjHbpuqMlWqRRlNB7EAaDxwjQSJ1PXJxKrAb1sQjcQi6aD/rXpAWD1kNriAX
Jk1tcJ9q9ip51bZlOKo8DXzAYe/1NyJGJGvdsp5gTpmYd6cjDqtgH45Zllt203ECW+Y4V4ZTIsCX
YFmzdYGZDOhZr1PMoelb6LPWOEuRIDCwsTgBVH3oo+IwgnI4eJjoa89qe0Zy6VX7qfIYtJhS5uqC
TruUGWhKzwMyIIrwNllbtr50jQNgjxZO0BaiCj1l8Qu9XF+xjNc8a3Bmu/oQ7dCur2WSiVOsfggi
z08jxV7Dzpj5pyCWl3VvfvTj4/trt5wfXD+im3370oB9lDd7dcrpTyPO5IF9xQaYB5uHtTl9Bhbu
EfhH7Le08k4yPEE0hU8iA4QewEhPZ/fFwINLaPlSnkI15SZdmXYLOtPwdLUvKxuSrhG38C0o+vMN
xR00gZ841VyCJDkkLqksii8z3e+4lESRzAspYoA7YEzuEmN0AcUSYs0UTXVEW7S6ZESw24ZbV4TQ
p/UEWC4lRPLkNDWo3QyvDlc4uJ4sDWSnTrapN6zJwBL9E/LeGOzsz7lZZOeHSQ0YBVPNYlIwDN0B
WOduhAXpix64uZ0CM3EjFwu3qTW0B1RS9dpmQyGofG2DL0PZqMUTojfjrnRLWS4DiLPfEUbpal0c
BARgOuC1RC2irEQVbsqBmCAwDHguk+RkJ4WJEFaYWO9rXmYZZE8zu1q1mHtby4KLY00+icH6b8kh
vn8JAYVcMXiiBW6oShcPicup1lN6X4IUWvBxdlPWBmxKb4LWViK9RqIzRFUVahbWUONLQ5gzw2wi
/ja4qmMy+rNdhiZZWNk1gVYajYSC3jwhGgr4dyqrGydy8V9413Rn/yjf6wsoHe9SHCxMeAs2RYCs
eR8DRNSBkYUn/OavYtbbL00/ljj5C9ALw3qeZKCxFUy29amSX+7/FEhE3mOQ5ypAlT7LShSvm2ck
cz2LUqwzRpRFd6OgWCWFMd2FvitbB4xfGTmLMEOuDACpLm7R+C9Vf/XjPtvjZ7Cfk0G3hsiTM8vE
v2TXshGB0b//n1FU5fe4mkNpeHj+5aoM5gkg+dgqJa5nEeBbi9oE1C2aCssxKYQCfFM4Y3zZ7cRW
DLBbE55rHXGjDByPisT4bSbyzloEDT3H+S4CKnJ/Sd3iQfRavUtg5/k4kF5Q7Ym14rB/D+4E8PSU
uKAIZ4HXWn0OQOHSBAz4M9cEcMR0hRjT1FUOyISEW3llFpDPITZOo8BcbA1ZigjIwN1VP8dYi2o5
0wrnZda9ojJdHVLBQ0bFona/0c1Ri8d9mDyufw1pijApORRjogcRguhNwP/yD5IOZihH+eToplSX
E86c+GlX/njO4fMIdU5OTgDeYH9ItrWVZIK+EQQOv1h2TC8dSTeNqpo6LU22zrY0mkaXf6yIAZii
uWZs+aA5Dn1u4B7L4bwjszCMy831CpoiYJV9hbqy9xWqok+J0+9FB3xW9TLCE2uJ6MtPBkTs5LKC
Myki6rnFNolSl0Jt0XfDK5mRFQ/cXTUbhfEw+TbtxFcpn7tV0eedKpZ22TjlOIHmHcswX1NGbhU7
K90PKGYVMwnf3ABOC0RNkdKDFTRoSHodP6aFsC42uHmBEavs14c8yHBjzAmpY91JZ5pJMJAPTzgZ
Qjdpb2Ru5ShdE5IRm9ycCmaybbJR97q6MIigoT7pI0RsFxU6rHzX2VpmTqpHtxBll9kAjJVpVgbg
qFyAHKa9CgM2zxZfL24zl8HD2Ich4JYLZfOw9f7cuKzv4g9wnrML9CWciTSMYYbQX56avHcQ4JBd
y8NaAqmU+YwCcOtnHOmwquHQVuRUHbMq4lD8fGhCwYCLpyIfLJP7RPHskNN9jcntQ2eVikwScYLQ
lnsjJiRPZiRG7Ov+vGLTJLmHm9xtSx6wkqOjEAY+rgTf8BLxyhXC7wQULpcO8enh0zPCoW/u8e3t
MGcMnzeydCxwVyM0Psa3sfZkFp93ecxQ3WgtQ3LGUh/TEPyIzTSDm8iH2TSSIdDZDefQKj0GDRBX
Bdt2pk448Jcc2l3y5bbtO+ux71OjDGr+Vr8BjFwAzTLd3BlpNvmPDQmH1G+qiplmq7mImDhxUgFD
iSE5Sh8zsWcjOZh2XN6fC5GVvJ6uv6WtWHyfSFGpUWjJFi+AYYfh4/xJOQC9qRpXEjFZ1IQlhB12
E7Mxb4bRSKWghpAuaZajKRDbkKKaktVtQsv6rC0YkqDiFev+MLqnB1fK4PQeIYKFumdWXXRbVtcB
hmX8BnuRCm4yEhoxh9xMWbdFCwJ+FC/99fEHG5fRw+qliSFVDFPcOPzwpNTW5nygtUutKJLHfcFs
A0qbmchnro/JUvm1mqM/r9pY19fvZ4nfbjvIS/1D49QOPcutA1Y5svpse8gUrlVNqekHjk8bdSLI
DH9Jc5szVIh2i6fe3JEPBGUraaktZNfYioBXVN6a9tuadfJeqPnrpDmkqsFVbw8nSkPoYTYFXiBq
wrDKy4oEf5TdZhEq+aaSqd9n+LaUDIJJ6kSgoBivJnVtCI99LNliDYQizHdUG1W03hA5+Kz1M+GJ
nKGp3MGHIni/fv6i51I3votLtt5SUnloeZxOMW3xlSrdhtwon515NMtO0hGjl1CSp6KN/VO4VC3R
zmdmLlbmI0wc7x9ZzaHgOUpNvRtNmoVe8cL+t+mGemWs327TGIepBfg4vtnB+3edFTSuCS0Gcp0x
XW6gjwT286dL4EzatLODPd00feDdlDTp9PND+R8hK+YSqLEo4gvh9LtglhOkTJq5pRGSyvyBdyt+
7d4mxbhQDzHvDAqc4pNT0T5hjFSdXQbrBJvPBT057WnB6UzLOgWqT3Y5/nRHDlyDpezcVZyDnTCx
j4z1B9JkgxWv6r0JtCBCXj7oFghNGWUEzxs5Doc2sZ3DGnPeIiU+YSnHIXY4TFOd35WkZffXvmcU
j7zxzzA5EYO4KTjJMPvE/jgieVaKpvEVHQSOBbyNXyXEeXd7MyASw360Ji3XqdHrx3GtioEXoJgB
PQ69iuMRMC+nYpsJ5iz+oJmtSARmq3xbhCnzVGKVYTezxnsJMXK+N2vk166KCThlhRiGYq28spHe
QCQN0wO/p2gyvSOCGT55oxM1VQZykTjOyR4XPx5GrdvEZhXurHtyW7GnOVUDH/afOoa4vACB7LGy
Ghw0uZ7L2VZSnLOSt4lfvO7/rEQkA6n1PLsZSaUPq8pexCNB8qFZT++1YlAJDhFHGj4nvnzbdDBM
crPElKIU9KLTZqKiZNoYeUZ2GeTRDkwQJajGKrQTskXWrQWyP8ogArZVYST8xt8eywa0NCMvtV3I
Zigp67iZgFOJlgRyA/HyAIJ8SFur4x3GQBjHe4FjDJI2PdFLgYVFd2PqL+j8BrITVQGDhKJOoEY2
Ig4mQ1TgVoe+/nnw7wPaSsH8tV5XrA/x616BLgr12AjcPKFmoJiwCAEQ0NcSLsYsBBQdR+r9P3Ok
f8QKNtV00mO5FYj549oTsrwgrC7TRkrDejw8i96zR+uFdlagCErwakmv4oKu9XT5cgcfhBpGUbkB
xFljxci/jpOhI404alBwwtAAE2Dt5twD6mQumE1fIjLlKQNTfN5MdblC0clnOedVQT+I8BBSS9M3
WmZUiWUJG1oCOPBEM7CR2nwK7G57Q7UvCGY3mSCD/gU1y1Q/EPWOQp9XOY8hUiGOa2n+cSIEZ9h/
h3VIgIh4k9RjY1mTmM6usZNN9RuIvwy9fX7w3TNxe8PMaw/TEsO76/rJP228CympRAbiHhu0xD8l
9HFepnznuuQoSu/C3vYGoFNuWWkd0hcMAvPPMkcvcKisCrxf+rAe+OPld+yatA+EnzFyEZlTwB/5
fcD7KzrrqxYtuc9fP5dzvNhc+tEr2gF5N1XoPQaAc4Th3GnDX8BRm6T1IPK4ktvv9ds3AjUGBFTg
IhFGxep/TrNZHbjD2ZCLja5QJ8qd4JYtjZE1bRSv2WDYVs4Fh9XNenSNh6J2SqFPzRyd/8nCjtbM
ZA7IA4VK9KLlzYg6XZffx8rA6xXJSMUmpKpvOvBkm/t/zsZ0WEjnBqOqFPjZQVMgvp/ySxPNTOS0
/+oH/Ciyw+1H57MiN+cBBNBeltgR2EXZMU6gvuEt7OiIfnvKsp0hiN1nJPvFmSvcHUPjf27Fd0pW
R+iF9BrdxZQf/fy2tPMl9KVF2CEjLd3Mg42HfrqXcSyXSZaZmXewh7AjW5hPJE9AEw6OXQ5AEiGy
VJlUz0NR1ZgOwe9bnVuUkK8C/+016aIS96hrVx2tHuDjkfpFs5u/4rUgps7vCoeRjfEcOd2+O/tH
hQJnwG7Ltm3T2eh3XYx+aoJsXyEpXA8GbSxoYBs6YL64ZzTfBnReUnbHF+j2WyZkQQvDsgduCYFy
A6olTsCG1dKH50ZxGBRFjkP8ioe9T0E2MmLxJypsdjyZi+Qove4nooJ3/IWVouKR0UwBTe0zlJby
hL7G+F0iL4EqMhhL7182thVILJ6c+Qk1amFBt9zGHebWrKQuwA3SVM/vQIAr3/4NoMFU3fWOIWgz
RU9qNVuVW+jzNQ7z0IlB7UDuIeRwQBsvmBul+pUOZBlSkBW+zY0X0BqlhkpE7xuPrbFN2S4SS+cN
B9abIRgCPocnkSZ1vI1oSlodjuWgQhawF+pvbzSnvK7vNBYty+NoGKyujc3vFvcNGanezlF66AF+
e6knsi7YLU3AFlwqCoT8vPuO+iRQ3Mo1lChATAWlYXw/Yrme6TVtdMsyjBy136hEwp8Od89FBXng
kieqspR4Te701fwForFF/+AUuzPplnkAppbwl+oLmG0yaSGRhbRtOFvpgnkIFDrpDtzoVTBsqC4w
BGh5nR9Q9P7t05/3JqdY5k+cNqofVseOPROjj0vAMQOAlVe+Ns1/oZTfIgChv+EXm6OlEI6Ao4mH
o/iP3RdUe23VJbb5CpZbhJoxD6Rrtv2ujB71hXpT14Sj3ZXmWbDgPQYaYUY107hY+JWqi3qLdyqW
sYLPHeBw32fWbbE87Pv8duMGygQILLZM8rR5hnyGVBGY2WaLOfOELwSkK6ca0eOS58fVHeSOpTTw
++q0OOsXiMRQAj8gBe5O8qjPVBemqx6aWFVJMkr8+Jcw1uoE84Yy+vOy6dHB6N29QEmNumhrmRa6
0hU4uSiqDErq3fwGR+TRFVIuQI72S+TK3zNg9RhJBZwp4B/vBgJcYBn8/EdvMCsVWMEqKYeJYSPO
wVQFo5utxSWRZHVKMHftQVoM8715Y2/DoY/sMY2Q5MJf9ajfE6KQNFHjEMZ75pBRvRkacJphruew
QpB3ODZM4hbT4U0wHhQjoOWO3n7h7OXAcCj9LUvJ0KqZym2u8MbYVGAKcdF+X63ItfIz/QPqdFUC
3ZZFOJQAFFcsWroC+oDmf5fArr7qzJ/4JBR8fzjq9Tkb7ZcgEDecDdeLfYtB4hhopk7GKHqNO0dQ
bUs3m+mPqyob03FUgcZQg6BruCRH0slXKjdoPmC3Uq7Wrpb96C4AxFnhQIf1UOYJEzBE+Dxxhwhq
PY2VAnfB3xFCrVw/iNvzJNy9xo4HYN26XCoIll8RxSXtWq4V6peD7znHe7iB/TjrgegYqhBeyvH0
9zWRYeFiJanhaJZ80A6cO/OrCJ21krf/BBknqaBcKO6xDKSux/wRmM7vYTDgkUfSstlTKla91bVp
5JKS5Zs8u/Nd0UAZB1cssJkcXmJcQ/S4Kdn5zLaECPx2PMdUoEUJZ4TkZm4JMU7yRvgISIl08k+r
dJCDfmZ6RDacb23eIAvW8A3AhJrDlqE3U6l1mF+3BW1Fsl3Vq3CAzdpJEGG2yYEn3guFl6OYYXNr
SkkoBom6A7zBjAf/hdQNZ4Y360z4ai8aFGWj5zfYutKwzuQJqPLw2kOJlgwxK30mj7cFdjqK/SHA
xXLpACLrxSDxh7Y/uSTlmWcTO3hXTgmw07c3JewvD57v7/GwwSh0LtlN7udeyo3eu/zDBEL4mUE9
NgLuYmuKiP5N2cMCjdBdpjAwwU4cxGnaA+dYWqjTfuj3xU+OnEyAePtMIQiOndM0eudu+sDMG5n4
bbmvhE0HJCwweKY4N0KS6ugj6FRAogP4m2CeWlFl9H+xg2HxmgjbU6LmDbO2Np5D1fP2/q4Q0+pS
ecx49rgPl9TL+Pa7ttCUKlkLbUUT7TnKZVE/J4Orehv3NIW11Rpqjn9WSlevgR7Ly6rXaCXLcvwa
QpLZnaxmR5/HNdv+zJZyjnn1WXnBTcK06a5B3UOVhzzKEBBJA5axxUmRjOoPxCNkHmXhM5tFcXmF
o5UOHnu3SRZn6JXme7Y5t3E8cgfDaAT/dAAl0bKQuMLfnvx+hoVJZXTJYlyMQ1qWNkBSb99YmNSu
Cti4yON8M79EVmiHpK45QojnCMa9k6Ja5QF55XnKPK8mObymsUPKXz4fvXeZNcBl1mWSH6LcDI/f
Yh6DilLJbi+6IsimHbWl1XOicTgGreG47usCYmovK42WbBo9nNPVM/FAFyHbwXyI2/ipDyJag/WM
sGpy174cbj5Dn4U+Mug1UFcVG43GC+YeIvWvkAYpH+rEv9AFYIYpQal8r04VS4mmnhBlo9muqCaR
qGlfNllBP5QBjO/3ZA+u8CM94oOOdt1NTSy1qEChHS55OkdEFokQyMx5ex5690fG+0e8LaSwjhUy
FEwMEgk57yuGv4Gyzq+276VT/oqbSsGD7ewdvWoN7Y2pRqyZ3mhaF+EPlC8RWHBEfB0hvzszgXrJ
4P1JtFLawe+hdn4Qc2kpEYLZfrUoNU6zVmH4+c+fDW0FDw1kR/t1+cJtP4fkKfxcAx1AaMQEQdic
cV3izlmmXEmyk0rC4scZ8VQrIWbaY2CQ6G+q8g8YYDZgOPe5io89cUmlcEb+LHQlGjvSh43gwjmI
YFtumcv3R2gzk6Z9JiFaysaovSpYKy3PsnAi++u4P57F3nDG0XXA2AWyoaNWku0ajYYUQdUnoOvu
MEdP3kgP6OHjNWhpEvv3DxVfCYZ5WdT95RO6frmqynwBz92kbDH9re/HHrqUAQQcYjMMDWcai6iG
UXUW+268FnAxOP0DcyvQxTj+RidrguuTuTiQnCqx4EiwoqeMzOQLzFyYEKAtWtpHDNoQmwgfIc/v
fA/8Ds5PELncDsSpBvOvDkfHlJoHJtPMfQ85lE5mEp5oMrzYMZQ0SSGvYmXLCKBiAOrUfr4VAoub
MKZtFV/aIBlA7WjM6N64CGSttMptsdCpPnkBMR0kvEoDT7BAMCHN0ZxQTzKVhPtAM/7qr71cQPzV
dyfweLe2rB50B7KrYx5WIx7cwmKdHqYduXqAmLISTUsse9EBXCW8jvI/AKBas6ykMIvEOENnNAqx
DhpzbuIQefRU0ewtnfoDDrgIKxi9TpfoY0AEytqWbTEm0J0Lb2YZYajtz8GgU/PvUxcJnbqVA6HT
uRE2Di4tpOubeXwOPTx18U5ELn4PNAogYNLe+VFrMVxmt+TfZcoBdnqNo0HSact9Shlvt9rV6nu+
EdCok0HMjSuFJ5YMWnH2Pk9+yAv0bHWh7Ws43tP7zMUVqmhwj1eiKO6VpDucFuiQCXHqobB2KAy7
vfHZ24cQCq1O/5X01WV5fVPn5E45ggCH3VRLINujdMW58J60iQEPvPfOc4jYusonzxqhBWxQkUMm
jmUyjow9PeEc9Tz99WbKA53IuUi6MzaTkg68r1C/RkZHoHBSKv1kOTVT+1ZQIBOt49zXPTLSqUX1
kONkVrkYEwJT7dEMxI3UmTnnOC7zH7jiDPhXUCJvrEDSXOgeyla4s66fiMAZYTspfilSa1A8S42X
6UtzB6qNQT+ySfdiw41dkpT5OUwqzQlsZ6qPKybZPituVK2ywK5glWBaBrqaDt+JgMayXumMIM/y
dDUtqeNVCU+HQUh2LN6E+AsSgi6kkoAB3w9Un7aoO9cjwEoIT9ZBxTwzXxVy2fT8P3h39ew3lsGt
0KokYBVX8a1HiLX63/HAsDVg1vxLdPNPgRfiMC0bG5pwUyMKuprMlDD7hPCifJGwN19/ySOJC6a7
9ww4BXs2bEeEV0U6z2ul7l48PBjEiMG561+HUjKohLTDB9QIFqXUXu4lhUveQ8c1/diSMzj3bSs7
2jqfBkps8Jk4tNAG7P7fNmNOcdcytRat0IMnKaG7sfB+Ob5d2ueoh1Gv/XCfoPErY4MgYbzon4Ve
mpRara1582Nz8NjxQ0BXUxV7ONdaZLu6Y5BzaYj/FSHg0d8j7uq2roG/fKxF19ujnmzir2uAZDex
/nUCXRlamqS5I2RApQabwvoI/XeqK9iu22+/gMOXao89bJGOA+KdgK/3Ig/5mBfXfFkNCcNCN6W4
f5SBit7N78kXumZKam3ijvzBZDvROryuka9w6pSGGz8QkM+JP0DwAWe5qUAoKr3cDHDknnx+kamE
7oBgAu5lC4fStzgbFBbLig5TTAXx6cV25aA+0kSF1yCmeA5e11kzfagnJGPgVqTkZ+5TmlJWb702
zojRwkIOXjOkXkKYYl10J2bgzaHm2jozaxHb37RZFJBABpvfXOSuRCsxLVFzVisgBgB0T0b2zK5x
Q0fWrog6ZwE1tXGXTfEg7RMMKjOqL5qC8sO2fOqOsXkCoHXcJz41IWOxccixiJbANCf4dYlINlVX
KG6RFWW7E5Q9lMJGxHhm5odgTvMLiwiC5SyYloljmpv6/bBdBelPbLDiAAAy5Zjli0xCetgZ8nsR
lOG3Pt0v+SZv3tm5NGr69V5wfLgj69uppENqUSua1zhvfOkUB3n5SwEoYQyYGjLz/jzzyr+11C6g
s2cv8O7arOZ2+5S9PMIEFA1d4xemRyGHEwqcSM35ce4YqsIrO14bcjaiW1OpQuS9zO605hftYfxb
qd6Hag+S5YjXojHvcz0hP9776uSXh4wrjGwv+rkL4U1iIMxN38sTUYjiQmJmQX+o+3aL93zvSrDx
sL0W5nPxmbyyuAnAOyovfiJJbIKtWVNGsNz8cHlz7+SduNIxBWL4oS4Ah05ndgFwnRtnS9Re3fmM
tUDfA1wTn0ocOPomXcZjolgN5quvkq9VaVCePi3Pt6qSTWW25S4fFOAyuhLWipS59RWjwMhcogsC
Ew8a1dFycO3o3k35TfcE6O57N4NXV1T96nAEGC0RWcoavLApIEKyGsMThvVqiH3ha2taXZoSvsct
mmzg4f4pS4bVj9kHnfuG327gvCHCVUojV5dr/i9BXqqcttass3KzpYEtXgskv/wdUq1fryEWcFWp
uRjatvsiTZWBBYnQZYDCbiZK+ORIyBr8KkkZo5M9mci/4oh9BGfuLUlA1a7+ApfGn9rhOQeTfyXC
keYY6BVI2TryWKosjqGQuUvagC4XasabdwhLsyWgBnAs9RcB8N8lbbuBSbHz194SCU+ezyBVCeHM
zCeWOYtkBzY0uoDx6FfKcURvu9zYqT9mVhdt4fTLq1QOimQYRsbjsuCo6aQR2gyO0bKr9coaUvpt
x7x8hOZy0KbQtPqxYYGIhMzCgVtT/8Ag9jI1UXOFbN6xIYeG0XLib7uaH/eDsr0jmHoS1t3Z36dW
KcH0ek9IJRP7EOeTF+Ruwadnj8ni0bQbgEUMX0ljjh8NSI78doRhzEL/D23czjXOtdWLjP4Yb4L/
ZmeYe+ta65Mx6uogM9UfG6kgs3yN2SgMmDDDEtu/QGVR+/MmdswE5LqvJc2mgMbNRzC7VWwjXmnH
KiQQW+dk5FbCgYlxwj8pi/vrAtZ6ZxcowLfsDy7PnWlbHXQOoCHzjaKcuf4M/koj4EewzQy+h4ZU
B6sGWEpZkjgy2R99Zoin1igaPyQShhENnEWiRb1n0qut9zNum/p9/Sqw33k3pr8HMOY8o3NA4AIE
spgfLEqAZi2J2BVzSP5TpL49hZlylmPJ/sRK5L81z53AKJ15z+HCr5p86BsV9LhirgUmRA+D1og0
u6NonqmTZe5XqNqbhn+QA4rflzeKzT/A2qdCM85x95/o2a9yCZfDxq6z4l6pLq0/YbIRoiUg5mcj
mUOHQHU6WwOmFrEV+9aEfZBkIeIJ3wm/N3buJmal5xm2NZBcGzS0AhqtFWFQB0o4oaQqyvZXYS2B
3PTBK0aUl4amYiiV7I5MUeva1TdylbBQJbtNfnClPsQg8aKMMFZue78fEDGL9LOERyYkm3cAwMY3
tJ8S8i3DxI3OihRDWoXgKgpEjxS/ekAHuk3VE7rbJyQ2jkE/B6iHzuxpZMDIKRhGJ6JJXvbEJR05
WglPHORuM94Cu838kWDAdEbcm4PrOGDq9WWlqIiScax+4j9IQEUfT/lDPBeZaSeuGJQDbT6WBQZV
INpXW3KW7iEqXTFpCGidoXcXehooW/O38kBczvtDf8jC3M2gPmRqYj5xoRCnU29htGPxfJQMGAva
lDtRaUQt0bfPPCYUtlSvFjjREcQHge1CRo+jJjU52Elminolg1xZKIyAsMzLuQGzRayVBCo6dsiK
s3LjZi7GTIkjQYHJ9IvWyW+uh3TtGi8Sze19JKK1TZXC1r+fIzH1JnlDiv5JYhZZcwNpV0dgp1wH
LYnLBlqmLFj3D1GWRs6l7OGcisHtHwNL49cEX+uecSWH4j8meUxlNQRCykNQOuw1NiLEIWi0Lvk6
0Z9+N6pQGYcyEFKlZBX8Hg==
`protect end_protected
