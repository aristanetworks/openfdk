--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
CAqoKu9mf34DwEAm31jFybWI9y5XOetf39aGL0Hg0/gm74heB+FfoCiitihyrJxJhpfCUQYqtFZl
FgSOeLciX7U2y6mHErweiKqhhxoxuOA50MOVzlR4Ydp7SDyAP1/onBljkjlVh/xXK189c25Ag7ur
/4vXdMNjFJ0q5XJSpWSAH6IDyiTvkoeSak8xVE1pLHqx8ZtO0EQbgNmemJILwhRj66f/Zg8aXfiw
hmHddEir7loFPhXIOlxZTXQGWr9bCNwAD0tJNPXXV9H7XrEUOfPlNuVDQs0uOU3p+LzspgXqQM/y
2Kc31XFZ/ApagbVmIsf/phXmM47KAuDQIfOpCw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="heM/zWRGfWv/CPNJ8RSlN/ZMiY2QH5gi7AU+sU9s1zs="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
bc7gD7WzzEhItvbvMDcPVrXwMvJkHH54y96PRMmhQqVuNckpN4xhtMvPzxtWppo1gXQzaXVJzfLL
L99kE2RjapgZ7mb/ap7FBOkUlhfHcBF6i8KLe6SKVhRc9RhTk4Fm8Ev/pQJvQlx2mFMIRC1+3Wjo
D3EHQbLGNvdoR60GRxJx9HvvY1rDeIJDPRLjmA1wxoa8gdld+e2lI4+u4RnMgjZL5WuDoYVWlS2p
+/qH/Qa1OXwaafPiy5EypmqY217edX+FVKEuRsgcb9LCvAFQSgCP+LmVWTa+Ru1FOdR20Ag5gJ0z
/cf0RjdDVEF8djt25pNEaQdVKPdzPRNFasZhFw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="4OkF3j5GUYC8WohJjUcXduMrcSgr7ZmWA+6ncCdDAL4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9440)
`protect data_block
p7R1Fi6ixHktKcOEBvoNdspOyFY9rl1dhtTziEDoMnspcUMb3rJe/YK41nHp7eNBxND7z9TW0xEn
9uMwl5SCfRpK0xCnsP9J68dcyy5bt8RuGYiRa76Y0IBENfyJOU1oWLoT2TQF04H0RKwJ8eYPhnS6
G3T/+tUlmcOoDJB9z4DTmpPWVIZ9l9qfKh4GCbPC/pVQfsG4wVd4o8X8zjcOskRrZ6jPGOmPb7dR
oNfg5iVBlftMgeQGTaDCSG9z/OPSREfxGSWxQxnNN0ZagXHK9bGii1L8TmNuLhSisM2pSMamcRkd
OBa8veYndd4VYK2/re9PXOktXyI8jg3O/oL+4FS5a75DfgxcDvd0nuYwWsQRpv4LJXQfhjNqbcuG
XTmhTTASUWxqtvKQQMVorEhGzaJyI9OE4owEQwV//ZeT+UoBu89SdzxEMJohDhvKh1vg+m/LcH18
uIBPaiTy3iyK0dWPYck/WPe6x2HU+vDjgvQbmViH44LT6DGwCkygJ53cZRfq6NMNqgJYBRhJ+jR5
yvdt+HA1MHR+/tCxStpS3x82yVRQ4H4POwUVAh3v4YBF104Zm9MdoDbM9kX4ivUggoMsvMVJxvn6
3o8y4n9IkDzgoDBRXxYOgjgtDiwc7g3SoXPWzqC24t91HF0DxcFqtEt3k+FlfKPharv/JQAhkebC
InLFh9oZwPIuK9HjpC1n5XEi26S3H1bdCOqVP5ZN8AOPh+M52Pk6wDsH49EdYMVf9UjFgT9q4x8d
p0Lmzs8GJOtXEbZ398tVsfQfcYzlMfW2FmsMwD6P84QvzGry92wjm1JBQdIw7DQUFp8VONiOQSnN
QkS2FXPNX6A8s3iO0hJLK2PWozHTYdrqFraSaspwNMNr6/UFAeihKUJTKbvWbMNgo/fE3awFLdAn
TBGbdnGGcLe7WOJ13gOKyzgN3K3fGt36YDsjQV4Y6OxVzX6bSJliE2C6Zqh78jPH6+ojyXhhrnn7
d2Yw5mbn/tD6LVJ7L+KoyX++xcy1jsa8iN5WsccHsqjglENnvKt6PA26ZgxXIUVmO/2lAQqFdNu2
vtLF5015cXE8XAX5Tz4KqahyJKk86UThG/GZGIeyfp35qq/IN0hJ1XUrlPctRdIigvJtlI05bmnR
qdesLkR37LIGwwX1K3RIjPrEHzGRDW0h04VpbbSHa46OFetQi4sMdoBwJ/CJJK+YG4vyCBnuuIpr
1IPYOEjFjG9ablbUEeuYHqS92mylVjpy0U5eKMxmMNOqGi6meBsAnhFsFewjqBos5oLGx+WVmHGJ
ASj8CbTZP3YItXb4KjICTlOVv8VkT9ad1rm3BN1JbjnmmsDgjA/WLSKRiNbB84y3VMzfDea0jV/e
K8nfP0WEDVmgABNrIsO8XHAIg8EkfWondFzBWrAsBp/dKdmRMrWLsmsvIDG3WJz6I+u4X4WrR/IO
FwmZKIKeX2JeBPgWI2DCjsc0AQV4Pl94rlrAD2hqpgKtA/XlDX1DEHyiissoFB2Ib4t8jcppYBWv
k4eeymvwrLyeCF/OkoFxmoclv8VFtO3sverwsRnjG02dq/h0mcxNhoJJBc1atNBw15Y23v+imK29
QOOopYRMR9Vhaut3cM8a+/WL4ArQ1TCAvg3fe/cHuTMWlcQd6pctSuOSf6LLGz2NjPfx5G6eP9HL
hZTFA9IC8d3SZBHzkFlebAgPSx92BzW8QgNkmq3x/8JAVLut0ITmJKBBnq9tb3nxC4jcfxtiPTn5
16w5RCZh3oJ95neNlHRWc9Q3Vn1J5J322itJu6W+wcn/PSwJJL536nP8g/z5f4zU2Rh+bn1ZvMGI
F8V+LCqO9sGPdi3JMBceds6I35tIncIPh6w3Iao68nVpzsGcRrA5phpBgcIdWtyA2ZihKp6Donln
BOtsEw2n5ZuPM406OjMJBcfzstMhHGhHAZgoZBxw+PLuvJARBOFSXLu78oKov2J95evyclShUdGx
qWN+YyOtoKfgiCLSeJFDEaFWiZkM3/Lf3nLR9aFnp56ncSCt3QYIP7vZpDW02GGhWO2FK27WQaIz
sdJxxPMBaHnxvKd6JgP0QeFW2TEbDpQPLWfzt5FPJ9C+6sn44NkN9oIugSYO8ESM2ZgdpcgleucF
Efu1iDIK1Dji/wGwE4ltXkoC/gGV0ezIIb6hyMvFjZVIOXQP+9NIlSkGox/3kgb/Bpn8FkjCT/JC
AhNrk0lBRDXMCVmJWzoN3mFlWc32OQDIEk1DQSDQQcquUWrTT3zd4AKz1FZjsI6FAzEhwaqX5QsZ
g3ndGx7+Vjr9GKGSzWLtmhbQweMk6ltOq+Madnit1hnKqz1YEg5QcV6IwlwkkiSqDf1OCkO6z/x4
LGq7fglSgAi6l4NmWBKBFxQWfy/WI6vbDBoYjhJiF3CYXgcUCoL5DnonZ9UOfiqcbrbh+ijT+6oJ
J9lMN1XmtRxBciMH0npGa2Qma2kfWBk0AJBTflZHqwkGuw9pn3gPrAqFWInaP6XjBz44ClRGH49Q
0fs9p+qgrj69WwCptmxiMGGXy3fFVfC3XgUdi9LqQdN0OskagnjZHSzm8iTAB/POkJx3UUL2B1w5
cFLTXWz5R1I4cMwsnXUNOj1jE7pN49DY4PB0tu911oOUbe485r4/ea98ZkXw7xNGHt71LlGnySbT
Qcn7JxlD0mvHfxGeiZPDK2f6pANJb9YFo90Pehsdt2WOFYdrtw99yK+8Ay854uuE7EYrggD/fHWR
IWcsAzQmIcYoh2d+AqtVax3dBJvbfoO+15HX/jAP7lWA8vjSUTav4bF9+IKkJwdiDeniYF8Mq019
mSSqsHPFRSt0lr1njOlhAKmUmt8MPxArZQ6mpcGEtRGINxEYy+mBzLhTfo7mZg7r9NLh9XxRc5pN
xGp1N8Fc1HreRvu09C+Qu4LBYcOvTEvNaqqEWIQcU00dwstQ34BNH1MEP/+h95qI0trch99W9HX+
9b+LOA6zqoUEu19kTlwJR6Ky0mRuAi5cR98bNaB1XKIyWYkmz6NWrfv+/tRWbn9NZ20jjvF0OUKV
iykvxjq8f+wrhZqIMWTj7vrVibvVUUKdcrdv1KqlkKFOr4cW0Pz/fRj+O0q1jOHWerWNo+ilWMbC
XlxGJNpIEkSBs3MEJ9SzybvFxjb7EjuOArOEutBV4v6bpKGCcHUNjMGkk9uhJM9YncUJqgzi8cXE
kZ8Q8tFD+ueQe74DwcnZDnRWf6LHSRNVKOVU7/lY0QAsF7FkqQMbT/Soc+AmfANz7uFSEg1uIB1T
CNxjhGoAD579igRIEJe236vvQw6ziS3Tkb6YYaoPMlW0h75lYQKBB7cIoJd/ofo/XEDLorCjlfi6
uibHVz7NokzRA2NojlDGqxKASZBsqfJCg6OcPuN3zSo1X6VisY4ItxyEE6PKXXRewwvuMfCozm/d
VyRPnCrUL0kY8f8pqoHAkL/1mjWMt5mepFrECyClphPi+sBnv9ogorV9vG246nzExhfFfa9ByZxG
EfgTSth3uILXS9ziZAQNxMKtaTKoZFmRJb/YWaTI6xvtlcfuQNL8YvdX1mi0MVGSxjePg61nEJpQ
3+t4MzdL0en2JZ2dNwrga8SDf8CfTqkGBXMW3U6WGfHG3XZLHAqM4AJaCO2ULhIknVdUz9hofnTS
qSIVT2RyVLVrfJfSJxyooWzwEWYJJ/RoBM/uaSB5s8AqgoYuBkk+fRz3QwngEGoCbI/JlayQLil6
lKfdPgRvSxlZlr5XnwdqbdUoeheAuwUoQaFzvgyMfaFqKDsK51ZGtpFW4FiAsz+QQ6p45Y8XlDfQ
lxrYSNtDPLEfYkw1xxo65LDK1xs2oJfD6CSKtYcHH+9wQVTKErzO4kSegBAJ8FcBYlcuG3kPWMnK
/lmfZkumrXRGBTdZnentekE8xocXaDuYOFhFngGdaIzC2z3Ixv1F69dFtVHyTnZLxqChQo08xYBu
iwuf+4XHKlCN6+rQSm6qe39JC9z8AK9zucvrTWXOn78Ck5DhoXGfTfB6ATKdJuMWUodVot+ZUenM
UqwLZvcezRz9/1nW+lRLdSO8Vfo5AjjCglWqnVqH87A/pZrY97Cy5PsmuWIFNO3rEASy/h4Wntm2
WfEE3kzIZ5PqPFMgTK+kowv5yy0zLC/au5XLyZRZFG8yh+jxsSPRiR49ZKZDC9k2thRvRroAnHH5
VaTBOisFMmoqlP8R0p5WkLmi7S6yvNn0T7s+2yOih9SvGgJXkYWGZ2vUEcgbMAP2DjImlcIUerj2
yl1HKlU3+ikODCtJLZix4Thxng/NCJiJWNDw4R8YyATVub/mcc+wM2aiJW9CNGHp5W7wMRqkJ2IT
aSLKHO8M1HbN8vtYO3wIceKh7Bn9A6Aka8FI7RtiQsxxH8OcZ8iJJSd6zZXIYjzrBAjESt9MJBG9
e2rdjNkL7riFgvt9ZeRrSyeBFvaHOcbrXfGgNjjHk0r8EeKAPh/JHiXCx9i94NfFf+aKCriVQMtz
zp+tBmjYNfG7S37N8sEG6stqWSogrmjNr1Qmk6ggUrU6c7CZefyicrpWIE26SHq6YW67qOYR51Se
Ep7bVe5a91bkQIv4/ppE6nIXxhVSPAL5XgNmqZIudm9+MK2PEmahuc+TvPzJXr/BL8gnCrO9ywIk
tmtqSkWoLZcdiFBSm9LP0knqUmH/Fr/0+o8Jichcjw9tLRWrX3/5IHooSbC/s8MFPdvUHB6oCh6H
CRBfUlU65OMXjWX8brcXJ/uZ50A0llHFJfL3nbMlYsyjiW7It91Pb3MRqA7RsECifoeHeyMUHpHZ
RCOjvX91aCK/MuDFODpgTzgQE04twQtmCkmmvC2N2TYcF2CghOVLXfW9MZkFzPwtLqffgm33m/88
C1YrFMmfJQ9EpfV7vsLWSgmVqeMYo592psmEpMMmQa34M6Z9Eg7xA4z0MXPI7fd8JQ6NYCdDIyD1
Gv/WIFwdsiRY/V6CSgGhOyKUD2mge5xZkaBHESUe/e7pnhxPPN5h8Fw6F44kgOYGM11gIPaL4eDS
PlO8wQZMPJtVf6D12h8jPxy14M882eLaMr+w8pv6yDnjHeALdgnTYlu2D67zbCG05a+EriFdC4Qa
yNur80onrip9f6502fLz1fFkxNvK2QhzL6FKmms0sLBOzVKlV1tL1YYvXi/cjSmrrmgvmtz1qWU5
WHKKOaC1M9q283Mn3ZtiEe1ae+3hO5BLL5bjBUyjdCOd3vKIYaNBgZuaCpoBDc1tSRy2KTOVTRJc
/3Q8Gv45oRHGs6VZRhrWzIeAuMiEyZ22TTPhvOU9BPfWqTknuXVfn3UNs2NwmTuiU7Ld6puLgNBU
5+IwlT56tOMCGF9gIE3bh5/G4tRiNg9wTFvzRJ9puJEzaxi0OTnZ0AlmzwtbiKuxUqBx1VFx6CJS
1ElWwCzaW7SQ+ln7gDGZhpLLSpNUkjuRTDVqpiHLMdeVbXf/GPA3bh14TLINSVIT3KMjcGpUEHxq
hG756cGqb8Viua8xUZP45sWSIt2qGrYqXM6B3aWbueyDjXc0Q7OW1LAirAMgw3hanhiyPBXnOdHK
I8VQoh7UlfKMX7OB8592U/HM1cJYb5WYb6iMq+qsMY0wAo9zGCe21HKj8f0+j4v4gMi6CLKkWlwY
eekzjMjmleSCNYvNXSfqftMsJLNTewIMCtKiKChuB2WvAwZghtK8RkWUcV2QSOuHFC+PL6D9V95m
GKvPjGRDLHGp7UMAcsWQF0xrR4JVzhE9g469H7Fdp6580XmrMduq4YTzQj6Q4hPiaSGri/lVee4y
ylf1nMc11MaMxmJAeoix/CK+qFRIi7N0ndCTlyg8toeg4btaY5jYsjCN5zBhinNyFvi70AjiEqxH
4czVoKu5EjIH6OC5wYdF1VicO7S14UZJhngeVHDAW+YIVmcpDmYpLPtcmVcwDDeTNAwPU1DOndZj
txUjApZ7tfnCvpPm6zo+1eXP3fZNAmAM2qq9vZv+KEPv64ZkUxcaqMl8ZQW2XE8P2VjdTExMCWVz
O5Xo/ovSM8ruvwMpXXOylOEKaDN9DMjt852YJI3NMoqH7nAPJaaQu3j5e/9wt8ThRPsiEVXAlGPh
I2PB3Kay6BwCGLbr+kCI9izxDvF103p9+oMt1uxtSpPkimov2E0TcsTFkgLr5RbPr6mWf09NYcE6
ogEGY5Sr6oDbqu4fHK+enSvDxHlxApU6ZxI7/ywsDFNq+9uKWGrxMZ20MNL5kFHTPauuTglcc/3B
WlXA+phZ6jGRQrEfqgWPNgUM96BPZEh4mNxUKEZ4gAAU2kwinWdRLy2qR1eATzHbF0QrjfkMyCal
IPn2Zf9j7QmwlFgvBARhvKUxXSlTjErfqL2fdNzZLApZzBz2JrAqDBCI724jbS2kRNOBZO2UgkPD
DdyN0jlGCQW01QvpxnUxMX2N2O5Qvd3KMnj/dqTz4ZiCklwOndMcNy19IobNh6jx/bajnvuZ3dzH
D1obbSiJveMrfgfTTGf/tMnj5K88QLiUcsljmtLMr8fHPxe5zEHk4zPBBfM/uYFTSTQ0Qsd6hBqe
vhKaBdmkV81ranKYgJI/p9yopkeJioNr62x7gP7YDZ7fLA3/2xk26usvfrzQjm3Y3ZCL6+IfFA8x
cbt1hv/posPQdZrG8NLRRTyyPiuDF/dLDf/wIngncAVtrqiLZsIkO6IqJtE1i0kUrHizUiiDtdRd
X8FEDS6IerGJSGc2heRQ9dATq2OlxBCalmU3qkOAtlPac1dSBbe35vdwHcDNuk+J8YAqQRJnKKrW
P06v0juqj3Av1WIPi6EUQrvi4a6Ss3cZ0546lNLXbTo00Yz+8TBmbA5pJLoGVgWzzfv2cQx073E/
PJffh838/kMnsobCI/yOPExWchV/bxn6860UF+kzNisiJsY9mF+DfrZz+0TNfgzX6hKLfBT2h6es
vi8JF532ew1uVc+RWHaqklxoWMkdDBZzLZ5JC2ni7vb2AYP5Kc39XqJiY/CHHYUWP9uNDkEPMlbw
3uEOl1hlqiy9otCM8UFYH6H1EZPZhRXRVHj9JLdlUx0i8A6AP8EO4vMRGxmEYJwq+EnuacSCySSz
SklMgBRgXyqlCkfkPKcfv0paEygAA6y47aywtqhc7JzBER8jey1mLZfxZXcKNoWaUWyEeXNNeKoE
GXIEy+TyrrEuuB8T8a3f4ajsabljyOjvImhRtDrJfbyr1ykOBiDci1+vCF+bfB9DUzS82wA39Rpt
15mbUkWdCMKq1Or4VoE+iF4vI2W7uDSXmyQ33jA6GDLEt+ytISRv90GuCqSzw9B6pzFA/mc1jbWT
Go03vhKBjPv0rSlV1fjzo/g2fiXwBjtZuc9d+XJ0W6KCPsFr8fQWiIuDutMAc7fwqpOLz1HmOCX0
2x+H2DgD1SQ/oWuGtvNE/ltBz4Z9JhtlThw8PPXhHUVRH4TOpF2cVQxKO3MxmMiujHNGcQjbR+qw
sl+5Ja2ITJVZ4qpHCU4EMpdWu0dyduStpb/dBmPeGol26amQ2xirbqn2gEjqi+QY9h3Dv0Sxdr7r
39JscJmZU6S/AxtKNQRQk8aXiOvrkcgokXYR9ZVBYqM9hFtRB7IGBD+WvSzZYsJx+96Rci6dK115
xlPRSMEMgChJcsUCa3yeTax3Fku4qFnqMVZse3KytBINc7FMUlPGmeXnYcjRod/CIUqQSvB4/3LY
RxZJpaBXoXyPeQZ/tQBcH7g3OCDqKxOzMPp/brqQwFaLbpZYzM907lkl/DVGXzj6W7AQxraiEl1t
SLTronhyURRWeIjMVlD4AmWT2Tu2gohDpLzmOQCycCyng1vN45rF7+UPkmyf5yVVQkHjt3th0nXt
AHc3TBw7UevM28bt5ivSB5xVyPXZQtF3A9hzjgdJ1k+fx6LfQc/ut6h13GKPwhRatJIdmyOzVNkW
JnqoOBgChj2IxF1NwphZ0ZFjWdnxRu/RxmjUe6B4ZFOCuJkqoLA3AS7uxGm9rntQcpM3FatvCBdH
otrLsR/3Ld5j/utJNaTX0hpBjnNDRDpZW/0mIxcNY0pBy7R0Uf4DPryCXrij3nXi5k/JgSVCsdUy
JwKuuijKG2x2xmg8PY1CA+y81MnZ6wi/zSiDLLIxDAygY+mXsmWnMSwiB+2FXIaYlg+eNXepTZ86
omqjN9rTMzPlY6vC67Lk8HbwChyBY25MbGH+lKuzZd8Weh8IWhMmTO0xSjZ6sTurBCSzmEjTICL+
uGPSSHFXsZCjZjMwu2tu8jMtqIZKiLCSDBJbM85prj6oYR5mJKCbU7R79kXTEPCvW+SkZ4Df1RB4
hoYfeeXEtGnmNS59MzoyAXf4tK6JvpCfAkuQg7lS4hthbNCPqgiaiC5w9qlc3jJO1BDVtIL03Jnu
JHT35s6hGI6rErP/gHf/RLHynP4vQpBEl8FBiUuXn61aDl0xdGDet2DBk52rW3EMupSd2fKHmEzX
KCf1jnvB2A54wX2dCUttHOYpsQbe5OmCY9oXQghQfjbrrQG4QOpmNDbb0ap0B4fbfYBvCUyFgs6Q
X19ArJgZb3LX1ap93HLP1EyCpNITGrkseXBXweASxD8A4JMzpIoYyqKTdQM2pBAs5wdFC0kXvGPK
FTu/mgYFesGDcXNZ6CYjh5hWvqFFa2AuEbhCE5LDlSzGe31sCVIimVcdSUnVubgeQJLU6La3mMr7
ubISrZWewB4MmQeo9xCo+pK7y8k7GFH3ksDpGRy/wkuaZFQbiTrfWPIA/NHboYS/GWDRsi5+NBAP
On/dudRY1r2mZqbO0UtKmc3kQLXBZQzhBEUk70DgvzEfdXqZmuWpTaCAt/DCSq9tSe7L5hchxol7
PkHldb18zSMB4aQZvxHVJ02DMXKCt/7mU8K9Qyt9zuJvXEnG8aCbauc7K4x6AseDY4LbZCe7DnCp
C1XkZ22EDlPzacuxi5I7MJHT86+yxXxlmIpv8CbQGzyKCU2EqIwy4H7wb9PF7kmsPeTNSqUnsnJL
c+cc7hyE01vxdoF/6X646s0WPGSS8Jwp7YrJJw/d6AvjQdzz2LaNePren95/gDxoJXAT/iDCdr1K
Frs1wzlmLxjPWZIe0wlbX9aEVbYqjAKOWYq8x3/JSk9D3YdG/qn+TfPVMYJnpRM8VE5pM+DqYGHA
97x96PVob3i+6c5qClYvEl64SbvMNFp3v3CxTo5uSQVAa+8eik47tVA90Aih5O4j2uX6noRNLhKI
InTySKCCfUA0R0FVSrp1C9GJseTZy0F8h0h4LTcRMI2HDGUwEcntm9sCXZzd+5J7tiLNZ4y/sbUo
ULdm6PCYo50ijU03SLqdvCHuTn8qCfhFjwXSPmDhw7rozMGiG60/b11hYJOI3kl2aUQWL7KMWS39
o2FmOx1p4fmo8ukusEB+9Ue0U2TQJ72fuICDL4fAJveZyeXkof5VZcCoAjhQC3tg0tMFtJItpwud
GMb684ak3mY2V3cGZSXSroAoTsmBk+mniSwxhoF2HXMeShj4upDodZQpkbSPd4CdaS4kTOEfVayb
pzjm0ajPPKc59YpdmyafKm4HACqO8SHyYQui1qBQ0FghxW4ZN7x4fGD900GJLDdEx29q1zu/O/Sa
EopmhYXI+s8ve/R82UIIwMp9YUAgCPxvJVjV0bm3Wj353YFE2KY9IOed9vCTjv8DQulRus2M8she
oiVorpTnV7rnYjXT86hiWRxaZii8eGJe+nNAZbmT2Jt6hFMpLHUD+iX0FTC2D0nC/OBsVzCYeFsV
j+FEG+GW6y+Wm3jHNkL11h54l8OrWdr5WCC3HQtbsooFNOQoS9u/dHEe/k+s2l1xALBtuO3sIj5g
AjFpeX42VpwausAp2OE3fuEpAkcQesGfS3TN5cv7SiAd3JaOohqikP4wrjM3JpU8/YmIld93LSCl
qI9DEtp2EJXPWvaj41AVDTuZDML7HTHfiv+4OMnyjewoan04k91NxhI1f96u4Zw8auPMHlwXu35I
kj/maVjGg9LsXL3QsfwWvvyc1Y8cYLVtDZfGI4D6EbIj2v0IXYn9iN7JnhKzRmxjqxqYBEVJCd/t
Vx/NCX4SpBa0/is3hUV3Inm6DRbswbJUDI5+uuZMwjc9aqbkvMojd8gYdwOouCWT1WdmTHfAWKAP
XSCbGYSI3npq/Y1alJdtWje5BjFpw1cw7qzp8bLObM6rA8jXsKN9t/TW4MoVaTVQfN9/7uKXvNkU
pGVVPNi6KjIsXR9Tmjf/ROnwa1hjnh53C6uPgxwiqfQQr+D/+I3UovrTYPkO5gbdA/JnWkeY2v5V
BSOxMWj1lf0uIBGVv8R2HPODNj4Fc/U0oljB3BJ0+a1Z+j5emEsuT8/sDdBtGoHjJj6+RdPqQawa
Zvt82hRsPufzhqp68eHOQjLjeEw/w2TxVyXru21qd4UdZkjgHkZ/6F55/Y0PNCVV6wRwtgOhyKNd
wWKsFOJYj+r9C3QfAW2yTydD3AjQe3jEd4ffovn95YyPCPSFUZSnW4qkn/K7RcrOMq75N+NVOdeb
vXBRDu4JTSaMyNj2I/5dQse6vI1m7PsPC/AmAneBVZQ1VnnMInCnRwlNnfYETi48FeQcq4tS8zFm
MaHKy1+NVPY6+zVTEa6VYZ9uLKWK6iAjs4uuF38gcDhde/y5Tjgd/NgoXs9vbesvxcwCQPJADIIC
byN+dSJdwXVyytzXWo7oTB2Bt7ZHjxgWLPTo2NkW4F7bwUZiakbSNc4rH0aORZ70MZT8UTIpUvB2
0Ak9VXzUxZyTKQcsGT/aPGuP64zBStQF+HBJ/kgyDGWkmGHeFQHJ7Ty32wZQtyD2y6W22D7dOehB
1nzwfCngj3WrRjYeEed/ZXnOceaYk+nnvZ+8OtPUCgyr/xWp8iJNyvTGQBQHqUWAsqTbKimlEOhw
DyAp8fBmLb/L4dsx6fsYuF1dUlqMPXHUMSauyQ8kUzeiVdTMmYbl0GG0kaWKWcviMfQ3lmLhUCnV
hGpbPKOpDQ8y1XvzYQ3oj80G+3t7Cxs1pRWIhRTF2EgWjZ5mTfdVR7/Y2989GmbHa0LpUCAA3OeC
5XUfisi53Q0263UTNExyhnxSKGncp/8rsnzXosoLfM5kZdrU/ayliQDceCHH3tHchHobSP3c3Ql9
cShIDw+jLPyZKEsjYRtIazOZqlOJgwrSgRMbvbyzq2ButyrCdJlZ299IVOcYKLBXHh1Go5rO8BqN
mVeFQelk9W5cV2oE0/hhcRQeq7TLOcYI3K3oaVKEVyah4Gypo/RMoa2Yf/h39dYKtwbQEyRQQpex
lBeK+TH6AfsCiXntHwxDO7/mpCXqJHr1RPFeW3g3nIZ2SnLS9Nnic3yalDCjqG7mnUEiFGPARkHi
Aq/iT9CfhCxVIXg+IAYZCDUYOObdyy3tW9mdnKo/8SOLqpRMAsLw9VJyPLkeRT02EnSNRADtYlY1
+3t+5h6Fzo8wL1nZEKkJb5WQ0tlaKPQ6ArKYk415rwWCPfhB//tja+k7jsz3ai0jyLPkkZyoGY+G
fNfTVaZl7NspoSMkAnmU+xVlvjbkDqENgwVhTK9YNFin0ky5rz9GrxHkHZHyom54f7cZ+yWmL2Nr
KFprgF7gv2pBeu2K71LpSSRJvQ9GwEIO7JK5jpUgDGAoqZGJLgoBN3oeSmv2W5mGJ2QsAgIJDCYq
18svaCjVYIpvBE5mxDZF0zywlqqbhh95w95oN/ZOD6Y7RTjfULH2u3MU73rUAYsg6TCM8LHenUBx
5iBTImx/ETXIeJbVU17987Y67t0D5HSIJriHrD9aVovD6iy2hBTKxq8aqqGkgA85VIMPMP/chEYN
VI6e3GD7tUj50rtra7a1rYoOS4N8orxuwdv1GSFugYyxVPnxcSyhR6mLXhpMeslxydrHfXJYwlRe
LXjseMlRQkwCJUg03k1L+yMeM66tBBz8S8xdk4KDCNC++I9J1jeeqrMkQkRZyBLseDBMpOMpe63c
3JdfovyI+HDcMNICJ7o/HcnOkq5Y0MgREOpGwPhEXm6OD64p/dhTLwP6lRWVI4JPmoif00NHfrd4
2eKK98Cnm6zTtQubYK5G6YboUXpKKseBkD5XyN6RK135iN0MyAVEHaZdOg1kmYXfwkyjK6zk4DZi
oXSw4nh66jcIn7u4fFfyIh+mJnQ1k5R+EftmRXoDFMeLwMsySoSdqLd6a54IPZFCuDqirT0ynW6W
w+WCDqcXYHTTHCbW6YFP1dyPeB1hZOtl84YXlea64fCm6hya2fh43m8+jMyd/VEPu+rQ0qlJevx9
acVjkyPcy5IN37CyAc4SsxQpW4gKe/Wd6yzrTQBWIBCiMqmrHoxY8zINj+gDws1liIo5B1oXXZ+F
Nea6Ya4C8ieFFzf/GYAvr6tnv0J8jT65AROBbACTjSmZxWQPrgqeh8q7sLX0xcqnxzFWODm9YaqL
KFUzctZG2D1gZell9S5fACMxWMq/bJIpdAPM9JH2b12wmwawE9hJ7n68Wm92IR2ohsFs53CVX1g4
sounQpU7gqZjf+3LoqfPGXu+scAax9twKs1BPLBmXJqe89xpcwHRQo8DpoQYEuRpigqVGCg78A9S
TXCWbJw/7tIs7GWM6EVjQzhKflMtMmXZmTkT5VfdAZf0aS8=
`protect end_protected
