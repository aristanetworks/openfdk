--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
WDJY+k8SzTNUcEZ73X9a3CVjTI2HOpxBgUNgewP+/7je4hCyvG9JVQ4uXhHaFgxAkMJruVuBntN3
esUTcKXNc76j7pZnecdL+z+YJksQSZvQ4E81MB/W245LrJxDt7DMczU/XrNR07Y+WU+Gw8sIvr2p
BV/4sIjFtZATB/2Wtawv9X6W2Eqthu/IF8AQJ/TeNao42qS4plrhGUkjPhQ6ivo4SDgR/nMlTCWH
vAQyMSNWwx3Fthjfjey3PqGSYX19sxSX3Nyu8kXCnRVHgxJF8gB/25KpN/GiT37fhDpcMsNLSSpk
QUgWuP0/rK90QnJEacD5164ps2Zx/+fwmkYaVA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="V/1Lcg5d5/wU/c8MJxlg1dKiN/xE/QIpxT4drq28LIg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
mBYPdqm7T1kZ6FzL0HV4dXdKLlQJB37X8vsfzUVILjIZ6DwPUX6NXJkg7NinZJr0rNy7nWKMj2c6
UMLBstKyuZM0K0+AGWSF/eMRh3CgKMPOPqZ0XiqXEJjDxT8p44i0L2IsiiGnxos81iaxUdc5kWyr
JzlI6IQGVoyS3585LIBSNOScICAnfskqD202jsANmaNrbwRA7qGKMXgzigi+nKkzzCbQOoxaatRo
dQywsbkfkMn7GPvY6wB2sxtrBalF3vkYJYe0COEi2+u7pYFgsJNzN3JHx9u8cExh2Bq1wE/Evik7
cwFU+zIIsI/WzcYZTVJ3QT+cXLzMESRCkGK62g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Di7isR8aYISlS8ypYcgqGUdFsyNNwjlGF8S8OLE5mrE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15504)
`protect data_block
v79EMRgIWUX6bOp3kblGXWrNir11VS/y9PlmsfPoqyOgcgjq0i7lY7YbpiWybcsA6FDb38S7J9d7
99j6s+YzJNp2JNMX5yRIeA7zSbEZoxvAcPLLBoxg6KP2VBqPX1nisoAbKjP29het5adeGk4rdgOI
wOiQ373T0TQBcSv0iXSZkA+/CTGC9HV4k5tpR8YmlEU9bIteNXX8AIefLprebJO2fQ2H1THyJOXu
UUYJzwRnYzh8FAtSQg/E4+EY6MU0U4uvenAjAZtpB27ztEzPDqQOBPHDQg1NdPhY8c/F3WeLFUGd
oyP4CkAaZYYobfGD0OXh0ZtdwxnkZyj7++G9QEjT4NpS7s4QYSc2ede27mRCZAxCAdTv8KUaXeBi
1IQSMXwdwNrNtiqQ8Tq3+hL35OBksPlKTMKq9yXGB1Ga0TcQBZZi1UK7lJfPXcuwDRpseQPSuwQa
R2GlO5zSy2LUMajBq1Uy75Ddaq4TUMpM++neiSi7KnoreLyWyeaQQRL4HinKrm9GeNmKR7peOcC3
IMm7/Z6UL0DblWqhF/dfjaazYEeCO9U0cvh0waVdYQL0qMAYrjtXe3+RGWGZRYehS6YCTivvglZ+
5THi3sCMguRpCbvIeKyctijp+VAS4vsZSwtXTv7El0S5L6kaQZROyhu7zf7eWHD8deqmHOZwN/Ar
jS0y9oXzsJ2QTWRkZaLJaVNK4XKY+RWExP4MHTAq0riv1xIQzxppLm6UR4DZNc7vG+LYCikQcHmV
wHT5FMj5TFK20AZR+TUP8dfMCH1iM98U7ayrYYWpb2uuWVcaiunVmUrgdMizV0KB2cidmY8+idXj
YGDnVtXXYelotozxx19U9OA/hfxw9/+3KQzBlvKu/FrZpKHFtTPMTdMtaOUIzgvkWT88qk0TAyh1
OYAU8ZHKPHai+ZvcmygysSaBodgjtWaoag4w30opdsajStLxtPpl5GHniN00FP2gqKkz4HgoML1n
gJa7Q4gltBTcRDXKBRO0v9SwDTvuKaq2VNmsXP7w/eGMqqhE4VbFKhfl9J56nLXTjDtt2VjcT0ov
+otV1RNsm8oQW1MHWHVDUP9e5bXTNHsxf6hDtG2YPzETYXn4UEEVvp1DiVc7hus2XHPq0h29/5Sw
oHOz2bNVqc75UgteA5ocooT67Cw/Hbun4lcj/CaM6Nl/HPFkgE4S6VsGVG1gGfp9xjivEuHf08JF
kO9cG/ZP0Jg/07KuLkrQu8MHMekmNfdCO+CPzAORGnmwrtA/0YWOAUUOKokb4UNRh/9mynOVa4PZ
4r7a1ZcnbJCEhmtoxXwpwj4/StWLsxQvNd+0Dn6FTGvXWd1D7hKsa0kW0mww7bmc8/gExr6urA1l
xI0WsmfOYVtLO+3GwS9xy0160HxRA/gs6zBS/Ge9eDHeSgnUZE+73uxJ+gVi4wcpQ6aaGTBU4p0C
+bEobXtcRnCW1h6OcMen6CJA9zHq9TMirDfIv8RQ95wfjktmCZxPbNMQPmb+USKWTiJucptSbBNA
Yy3OkY85/kStAMpn5bA5J+tn6y2FuNRzsuB+uNVNmkPOMp834r0fEyWHqz03s9+MDw3i+J/VOV0X
k2CDrVy1xnRVXCGGW2PfTX369vYDwbRF2ZSI2aLaa3mlDY4+mrFMneAuR4jIKtN8/CLnal/cmJoK
zXQJZBlBY1F3UUcm309tM/vqouJ6etjki+nJxbnWWq6qKej2ZYqFqR+G3nV/PNS1AbP64ojBxMpt
8NzLnpw07xwlHrOlDuxKsT3nrmyRl3iLPvLz60siaOnp1YjibsV7G3qHLdQHsXjQRuBd/Rf0FTtm
ubx3+ZaSHH0n7zzsZCKEjv8rjxbDeKIMh6xNnn/hvts5JhOsuJxoIKoprdVkRNEeMwhO7SgktJZJ
h8M4O2s8MCix2uw9YNVNU7moeN4Lb2AEuWsxWIIHs2t+rOwWIZ5u58zrDrw5n2DIzgTSAh/KVN1H
qSfy9CwCDbDxJqH/U/f2loHK5/Qjji+scU9o4TlRPeEEhptg/rhPYsoYNPJQ8qNxAtGAgsgmwUfj
XGjFoGHUg6zAunToGzaTKFZCF84eSO1eG1DjpubTqmGOJJIWajAtTtKoXWi+/ACZH1XpBUFr79/D
ToPO1iU4ZMkTdM4trwhzauJRAOyY9kvEs0GbxWQGhnhjAOQfX8oLK3rgoFmbIFocmXIk+yhhV5bq
OgNMtwA6NJFT+1mFVohVu/z7Jj1pm5wO4cdcXdhFx5uySmsXIoPOKya/480g2os7EfwdAOFI9sN9
3pmeyyDgAl5OHyGXpNcQu/x6hupy7SDcdMTXn07cOegFKtCv7EMZc6taPZzgCn717ex9wHXSHWsc
CiCrc1/VRdPTIfWhboqkS/jjmLFjOVwNckQY7wZuydfzwIu7xdcPPV4/CYrhMuctU6UoKmidH4+Y
11Ps/BlWW0xgOPNAbPCQwBboFqAvYfhCD2tq6snNt1V4xOafQycTNc/sj+e8DG818qD5+wZVHfxf
awtke5QIkEYLXI+436DHYP/9uLToD59dMMjZNVHFFJZH7rKSPp8atJycSvmgfYoRKNkgrO84eoHu
hb9tej7HgK0btQdJz2UDKGaw3VhlKOie5b3xqn0yDL0/bjggRFzXeMqWpynQ9pSL7FtUdmgoCmhA
m/2T4aN31nSPB6BVfS/R28KtMH/BmsBq13c5Xiwqh0yun76Is53MJm8XxHioLrLM/O9v918ewg3L
0Skz/uOWkmrNJv0g8ckOx/sN+PERe0/+tQ1ZKvLJcEV7nrgDG1MCVr0qMyHynKjaKlKPWZCMVEMa
wNdG9co7fJKAKzEOtOr1Nn2a2OxxGongfYi75ricwMnv1at4Dyo0RhnyctHHB5rYODjyUskyJKhQ
VNo9vNReXfHH0kKUSQ1V56MZi5GBOcWySbwTC5OFsHCXjnxxqoDtnQYrxD7i5I+L06UwgBLWl2YA
7kKDfVIqJ9ZVZPB2JukLbSQRB9N5uIZDtqewSFMI4D/mFlCB/HTDPH6I11MUqENGA0PrTQeoOaN7
OQDt2LClje29if9J9N1tBFK3S3VGGXO8YY/QQM0pBKZXyjkVSQK0bVAqE2fltK67t5K20JYlbEjL
OUw5hc7t5aJXOISw2sSI9FqbdsckdIILEar6GC2jeS/lcRmjZmlhk8GL2V5s4jtKUvAfdu9dAYyb
+EgXgtXQSaa64tQNhLFGaj27yxlqHfKazAAgwfw9IcqXvKt2SVBL6r3SrqX4jXXPmLyUQKqgyWqc
qdBCoGBm17x5v77H2nKS9Na7gq2jVn8pWVCBbzQ7d0YDOYMiRWUSrIj5ik28ZySmJE3Uv0dvG/2I
H+y7OvAKzuNrTUHwpUZCvAg4PKBTKE2VkV4zjyYE36eZt7pYBG5FJRgjoVSjlN4D7//lWbTejng6
w4ZvLWif4c1EAc3bJosP45BZtHocTtFF1xvMYcJnXZeiwuhQgBJA2Ou1yWmcYaNgFpk1WMeV8Xv7
0nIU30Jq4JrXOHg0wPjnSRwmEHz+9tsNbVGnvVtdP3CQMScdByAyT2P/NAjS9SKIG1P6/Avc4GY/
rzZvnsn2bnDk3w+4QZSYuvSyO2/+Vdn8RWKlw7h4VAF3+MIDWcmvS9uD4u1q6eclQ2qPCfa2bz38
NKht+edxx+mV6ZCFm7LDgPP6yYT1cGJVFca4nMyV0/0io9y/QkBH8wij3jYGxc1ClpSTqqEuvmrx
msw5ln04OHhSGxd71Y35XuacsTwN0Vwul7Y0WNE/yFP8WgUQDlXTxtOND2eAIv/9QuNJzNi2eZoY
N1NbYSLORiVXAshqtf7/yUjc/hi7/pWYc4XPCozVkW2qQaMQlbt97MJBkEc5kYiuLAVfWnDLfqkH
BZ/LV/DfOIjrVbmNPNuz/0EoPntTbUm89lfYQk5Ifn7rXCypROQDQMs/f/jcXvcV0tEjLTPrl3Fu
noa/cHKYnt4W4tBk0T0rodkqzaa6vQJfmCvpXSLsB3Ik3g84p+MhSuJj5xhwe9RGWQmW8e2kmlIx
XByk/MTUYnnC87jxy1hjqRcj/eGoeph4X3Ua6SlEzVBiHjFjBDaRO1nsN9BAjgMl/jaGFvGKubXK
vkeoewaNh/y3wf/YuUTof3jq8StK/xlizfNhi/9f0SsXMJbNXnCYjyGJehTfNylc3FtXnAETN5PM
kf7aFgxjOgUJldmSHUUHKxJMauFe38Se1TxB4G2QjvmeF+FXN3yd2pxlfiGcviLHJ9pBUWwNnV0i
r78FWGiUMarBJYswoNuGgF7M+Raa3IL0H3YV/zyW/JLV9Q3Wbtr79rlFN18N0ZuZjZrzTE9Dlo6p
Qg9wZxJ5vo5VoRRZI7BEPBglUM+7r6OXyQ9rY2KOnpZhh7b27uFdWYHXxUR2OrOrwCUSl1PUMztX
691UhWFgbhjI0X0R72GMdvLa7I1IKrzh++iomiffGdoGVMntUkB1rc0Kp5kQh2j5TEUnv7UkETwC
3b87AOd8e0zryU/131L7am4daAEQGSjOyHwHIEf2J9iRYCYpAIolR1/7+ZSel/QyNx8FF0NGCLIo
IyCER86TU9mFIALMQm/cHDMb6z+5ZrXVJCoBHr45O4fNzwr5PchWAVeRwWHSiugLdVaQ12ob9a+s
qAdrY4SW38DASd9n/Zzwyiz7ArEjnGlVRvux8Z1sBpoFTxBKNrjtk4LElwVn1KA6BWs9dZ+PN8rX
gDFFUJl69Kn1ZbVYT+I59QQo3kWpbP52ZOfi4ZUFCzXqLjZdJPv4rGJ7XNEfGtrWq0vXTAyAOQct
wzBE4sEHHiptv8gmOBxcQBmd+suF7SMzESai4pmJnj8/WNtyNED3j8KV5tJk6PzMpjSyFbNC3HRJ
RTVAEgfMh0NGSpQKn3reE8tI3FVNaW14LK/VFZ+SR79NRmgpFrp/V46kBZ3BXQF8CCV7wgWpIOPV
6+8kSZ6OGjtuDTZPGavyamutE/WCaRTD1utEdLkNXsJPksGsUdyhJLVq740iQgz6Q0khhEdaKrwJ
6zPHlz7TNWUpS0JGzOymGPzqbDBf1P3JgGrs00C/8ZX1ziwFIForz1SXET6of1SHfjuVn45EJ+Wr
uJo0cEgIGGSF4QhMlMNESJyeg5GzN3t5gi72EqwGMy3Zu87SdInXdqoykzngFfPOIo0H0JOVeONd
6qFgyZC5vp4ZF/3Tr6K3yfo6vh/Tbk5eY1BdtInzd7JL7tnUdeWgvxFN0prdEzbewTnqNAsc8g3T
rECSMcGnB+hhx/Y4tVf9RDH+elvw0kPjxrZ2sPwmfhHkmFYNujljvRrfihYbgm8Yo75zr+U1F1L+
H7QSK3fd2aZTz6nc09JexOuTAL4S65FWCDccYU9q5Gxvz6H6mKh13IL9n0yVJjxsoiYQZTVqUSQu
M5dzvJ0r2QYQ2BMWuoTggrnzhv22T+RkcFpIN1jXtOzCCRQzyfxQRGW4n6F2A9Izq4B0oUjQNKvr
NkVq+SChWXlYFROGr8Vi+tcPzHSWH6nMpAKZXHbfv7NTQj+i8+R7vo41VeDE0GlfBgMwofR4st9L
pGVKg4NKHYXZ6fudChyJm3walP8w1sCfTgR5K4RYP/y2+PNTeH+LnY1w4ijumDsj5Oi3l0lqXduk
7PNqslX2ka3zCiXcnVw686krHvPSN12nxD3nFv9z0K5999rEMfJkMEuI0YNbjheW0TyRPaqmdAPz
iIQEy7KafJmnWHnyKvQvs5jFRFSx4xHvtenUA9jUfSJHzsfgO3HLcxPJSDik/W20sSHRisoLCK6u
nB+sskCCtLYB6JHKQFOwk1drNzA0w4psOZlgI8GSukD0pQwrcBOcbCrthOIehHG6CZDI2zs60FOb
YYW/tgxzW5fdbFCwWc8awLH2FpBVTlSy9AJ4L4Ui0nt77qYLJtzKW9D3PCdPP/raYZ1/wyc6/fHa
RbSVcJWZWNMjQVrEDwtX66u57Ma56eg21Yl3v4dV2fmKKuIfT5/AtwfuFOz7GfpJtY2p4K1ILxne
NTb9Lmesgje7OYM6c98ryflr0y1pK8GK6pxAyJfMQU7qAInVeyhH1bECiF+drODn3A7ngeTitu3w
QUSR5i8j0/HbjqToOvtbGteA0wgGbi1RfilGKLJT/PEjsjZtBDvQPRjNIfW+vIl6QvqiZFpfRmJ6
ulwrEnc+9C7lA1U82L7CPkNDje4U69di/d5NG56zWodG9CtBM8IFoA6YE+9AlMt9iBRhc5YhH4tS
pxStJUt+HzMms9OmxbsYIFySnP/yZZyrM9wMz2KAZJVk6nFUj6EVKyCTGcuNXthrES8a8uNCWzkk
TuoRZ5EvnLDiLtGNer9ULAOmh8905Rmy7EXbFnQkilrj6laLSyjhmgdXL+IijhNVMZx2rHI6TDoT
aqlx1pAHi1zcFkZkzQW4Rvw0i9UMJgWhqVQkRH7C14r++sREMxUz1fF1h5MEsmyxjqWibRXQFcfQ
d/TCr4JQFu6yfqxJubpBB4xA0Wh52vlkEJd4Xg4qYUbcHIm/R6HkPolQNerx6aswoOid5HpYHB2+
+MAeNeBpSVDtjJw2iUiHx/ViZ/0hDnCXo1hw5OKA6qJiXdPeZis1nNpjf9VfuGulDoX90Iw9JQPw
wUEJQKEwbjgHh2uz5SPPrjI2PizF65gtoAhUNdzYly7SCK/HGXTzbrd5UpZpli5Q9+4bZQ1gnJBM
woo562bWIWjL6Z4i67189zr+8gf35slX9d4UEt4KxDbr4AMcuQ0Jb/ed4BhXb8R9T+8l1bhHvm79
uHoQSf4955kk7VVUA79A7vlSLTa+dnMd4Ccufnfmh1Tq/YaM7mUMQ8i5GnGdtLUGFAAE3WWTEy3i
TTULwfAZSxTCFa+EoXr0kI7YnfnmR3Yo4WTsM38kS+5rGI1tN9zTVWEVZVx56AXaU+rZsq8RN3AQ
XW6iwh4GHergzefUDq16A6GCaN35Oh/yahMubMVwnHVKLb6+kiMxxqnE09qlb4mK5f1ATYkx5etM
Lx8JHLqY43VaGnILQamyK+v3yqzKhnqqwg+Bf9DwrohLEJFIqGCKuAeL88ISofc4WshCDjNElaFg
t7l1oa7mhN9enU/woKFcPTYgFh9yx4NpyzxdSnUpwnbZBC6w91Sqmjjs/UkS8bKxSsefFN5fIxd/
wKC4Qsy9Gfv15SGy8wYGMYbXZQhPAOqCaXonP8Io3Q2Qkek3Fk7hn4HdpF8LyqxnRvuyK/Gh/kHt
m/u7ywd9p0EPdo/Q9onTOME6FFmWo6FNpn4R+th0yMiatFce2g9zSBVp6WACltqlTZm5YAuHOD5h
3Il5TyfXFE5779HKawbeUdh/+PXK6Rppy7H3aXD1rJhHuu9sy4dAyRllQwf1IKLLFFfnONqN+FoO
ZgET+ye1/i4NAAyyC9sNobh+Mbmc53j2NSQMqHyy5/Y3dMhAAHbMuefACW0AbcrjuG9rDRNZ3ilD
w1+COXTxjUVbdpVh9V30PC1VaUh/2HDgXQ0TNYW/ie0Ctg+m9/ou37U8jZs/LOgHDwdxhEji5kHj
yD32ByvDJmrzKxkVqMboEah+bowQY/j6/s0s4KDGFlr8edNZ4gvbSf+d/BAuTU2yDbtZOkYKWrI5
e34Y0bO4QD2xx2ywfKa2PSYmYa4bs7lVw9Y6hvCFWwYaYg+sS77LWRGi/mtM2bLtyOWpEfOkJgIc
AkzbfUXZ06aaigsgHP7vtyhR6J3i255jslWCtG2L8ETp8HdTKgfNcr6QxttCtAF1/1HcZXjh5uc/
U0iYjHUnzrdy32nj/X7yVTybeRhIvbq+5uGXx0bVE2kQU+45dEUb4zVdNF83I10qxDc4fm+1p+5I
FP5yAQNspXm5wmi6pyoBhhK0+6iNvayyDtDJJiyPJbWB8wAunlP4uyWwAVy7f/rMnM6YRSlX4VMt
8aIdkzEbLwoW93eKgQodPImZGDTDJmAMLc+VfO9f+uwZb+5RThLtqg3bWHCXdn8NaBA7Bnl0W++7
fdkld61eOsIlUniB/cXqpiT4qboGyfsMpiZ/YRyW9VnFjB4D4ZZqQegv9hQGOoegiuBE1XaOKaiS
zyrXGrztPfyASbr1VO9DEu33852kVdQIAp7pii4SRlPaGC2txNqXygkNFaf4i2EjqexEGj9MpZBU
3BEbbD+tUIqxv4tWV+DfmUCBUm+QV/nDwlwqH5kBQlWUz9yTxDNYbrbAKxIOmn/Mn+yvzzsF1Dwu
t+0vIOmbCx+eofFFMjBxGO1QHLNpJlETjFkkOwTDDdtkadbIM/Wc9WnbyUBEnLj0Jvmv+grtHwvR
9laubwNgiR8rCr0HwySsvUgqQZFYxRZNUer6bRs4gkpS6UC2aq11Awo6+AxbuVjjfEFFr5cu9aPD
spHXSUWa33os4/fVBOizR02IPFBnZ9W+ioDDn0ayIdwDkCjOTnXV6Tig/jyfD6JFvDcNvIRLR1WY
HxT0+so7wr7xz1j8RBD16aSQZ61RWlngD6Y5y/ZIjzYLGpT2it4VEuLVtX6iR+rD3e3Ssc0LLH5u
chhmAGWSx/c0/00ZUOmz4kREEWK5/W3DtraWu3HbIPIiQe6ZCtZLQW8xZOV4s+KIU5Tf5OYQS7Nn
fjUNDvXNnbCCSqFsHjdicnb8jKr48fIhgoyZXFxjSFTqf3CStDFBqMqhbOgZ0VDfh9gjN75nvbit
8AyT587YCGKSKdi/FdCMbsmUy4CJikNBdJTRzLWQuoFXBL6bL/l6FFZNcw1ZAYMQkRzt6yd2U0Yl
3kLTEAiX+ppUV3Q7WJNJw3GjZQzkG7a47uG1oZuzKUpNqAtJWcN1TymB5KQdVSYm3QRe+k8syz7w
E3Xslxt3OPKFjCkvk90DTJz0xMGFVjjWpYyeQ10SKc2JT+13t1ARsV1/zIWji8LX+3WDNvxlgG+3
WMrtUFSBSC2PEuDjoF4wDu+k7YR/8f8wy0/TA1y/an7HanVpUybYUIX0jVXV6gmSTpBCwa4Tabj8
CXDqn1JosM+9EuQvRXbEUTRAmpMUpK7tjUOfxL+ix0+32JXEtc0Uc7FOjXBPl8x+22pyz4phKAce
hVyAQvlZSHDsaxnCsk1i3EYzA1LBD/c/x/Z4o27NIwqD5gadsHbIoaXpyrpLxz766qpZRKtJYgc4
Lih8kfBz9PV02QTQd9oCrHAMsdvl86qzElk/lqg/VgAlD59XL9RVM+w6zokrqq7WHRSiFXhO4FBi
WHZUyIJADcn50nov6y1WsK4gDaR/EWEXtPQ4PaUJKqDeoPjpt81JatbZotU8Xhgik0D9m4Bzjw2a
FSahfD4CTU48awZ+tr6i3XLmCGvUT+HIgC4Ulf3UHSedNhe260Y3F1REwRkLRV890V4ZXPGOXX+6
oc53rN5yUNk8QW4mOhWczWYIId3Y+S/RMyncD7MFyDxEypOkqYGXxYAVTC0piSshUVsaV0uF0f/X
bFVO7iiixsocqwaPEhZNuiUrfhA4+qmvvvGolkS7/MUIZE9UEZPa3XdBnnY8ahhE6UbkZnMgx2Ta
hbWIjOUK7q7rtq8XTbnR8HqRRr+KdvvFe6PRcZbGaQqhiRCjgbduDLHko9nTCGG0dGAW2VrzP7zO
lSnc0Xb4QJpGzr2Y7QNa1kT18ghLAiue6FXuati+lE8ptkhIOxsFD9FvWo5OLGeN8wNR5PYg5PZP
pERIf25n02ocvhE318XwIEbjzgo/RZc7Cz3cSyeyNZfoABnThuN32wny6Q327XRurjcY4/bj430L
X+c7cpsF/WbaB9CY21VCoonKwW/bp2W4GGFyhhhnhNrgWLPsboyEgNuIEK7sl1tLrdJ7C8hdsV/j
gubngqaMvEB6wz4LMIVOuW7D1VwIpLthkuh2thIe4PyZvGM6fRsaJ8ZwZrl3sDM08RwBkoYnaSJw
+Ja97D6B/GiKV53DopC04re+/70uItABBXiDZCRuHrCzzTgu1yvGqBfnH8Un4y3h717hJX5nkl0v
lwMRYfsJkUzJBoIJxEwk+OHDBPArfUY0KDtaM0DGmYTkPMPqdvjyk8Gzl5fo9889dPwzpjBVpEeq
J7MgLhodxK+aQNshbD6xTqS+g6KvGWJ2Jf4J6aIr06r2s5OpJagtH+5kkyvkZosXbmp7nUtzSFaB
m4x2FnM1Coe1FPzjDN+aOJ0NVYjXGt+WpJ9X2TLuyRrQOIaLeDpXAMz+/9cTOjEonxx9fnoYV7gz
QG43Ihy8CkAd8yFdl+cm15D/pMbpl4gA4z2Jv98rwFpBSigLU1WEQ8Y8zbKdahrCcyBO9sF87W0c
sY5/94OcMIJ0+y2Qm+lopNrrORoeq5sMZO4dZoBEmMezWcHPOP8Mr2fDvJHS8TDZEZ5I8/JX6THg
FRaZZB/3STC+MpZcYuXaiMIiQg/aFi5L6u3CV6VOZj5Ov3fhRkyCadoOXSM8RRM1xqbmGKietOm6
UJWc8u8kV2u5zUEWn/S9mt79ZTh4jtyAEos5iAp4DhTRasi92oSTTEROo/FbZApMwRAY4UdPSVA4
UCkBU5wtmKEIvmz1P6tD/MXPMnxgfutax/X5dnI8OIjcG6Ix18fH/IiEoNXj00cFsuDMXtQm8woY
YntQY8F6s7RFwnitmd408ww53ABiJfr56UAt1uxeiz16b2PnsJ1rGPUTz1lp8MJQlExH7onZIFKF
nMZeolpqO1QNRBCBeBWRSBhy9bANL97rJRMFFKmZybFYO6IokWsRZGhFAyhFVntXiPg34X3EXavu
cOubaSaD2ecxhVNtehmMhsISwG+6lQyAAKZzqZ6cg0baLjoN82cuLkyaMhTa3wYUcUVd/kxoUtlo
nFvPLQJeH5HCFtA5nAm3AqfVUzKTtaSbNbT3q3eMX9/fe78i2C5SygRK0LuEmsxilb3BQP+igV8o
1THy3OMBOt9AEDgVbO8dDDaciuk//Ksk8FhWnmeTC6OvQ7JSmk00KD3dfHLd4qESfMlAAW5I4VZL
9XjSL3mKtDNuTmkFWBw/p6eESj/YvW8EDW6DQ5p2ls5AzD8mTWusI/CQT6Du4CSKYIaloXVkqSc5
vJrd1ODlITqnV3HT61hlG++4Q7lMcBmcyXVrtOr+y3deTFdxbHPTtJ67/i2Ck6p1Lhb3Q2QzU5ue
Fc2CxR0LKI6NDX1OPtgD33b0WgWmX3Jt9AV3G2lB27CnXe7cR4eeCQ38JsK8u2lkps6S11CGOjGD
LDRmNGyrbaFFtv9rQuuy5gkcOB+y2jByhT+wimt/1wQ6TVCrk6aD0YUMsNx+j/VftIuvmTHNDtDi
8VAH+Yv862SU1k1cAhUacKlscgxfo80kleaTJySV5Wz16KT+chLBpY1nVz2TYwBffCZ+IMq61Dif
SZuDm+q7eFIClBRQjp3viTGTmDoe+Q89Au80CsE/ckylF4zjcZ/BxZCgFBV4VducgUzu7WU39JY4
OrMcoCSfDdMIaGf49Fp3pl1Fn+EilD0TSlWOuCy7NNfl958RcSF5HGwjMZaKk9SnStg9Hzzay1Xv
GQUWYG5EbCiYVj1uJQNqSqH0O0KshfZPUfyqz4kHWMNgOqsilkSnLtPksXn0KVnr4oupqRab7CBO
J0iZB8yIjsMereIEPTaTbyssYlSvECoHeBYcSKzfVmjbaGtGT79NyaFSVbDUkh2Fj7walBLzNmcU
lKzT8mUzKLSutEbTw+OP1k69Un4SXjfDNWJIw++Sk82tQA3Uk5zrdpxz7VNPtROcSkuw+JW7XkqN
nhm8VU/WQLLmimIwyq5RIPi3nTj24+wBW5FS8GAocQqjSbV0+bmWAWW5dmHwksNQQ9akY8iLWiUY
TgcmvK6e2KG/Ll5I40vefpZiCh75wahgG191nQNkkplLwJzObEVA2xkk3dcZlvjNE30V0jWG6HtI
a+2t0x/uWvj6ts8UIsEAVenT0y/6HZsBrgLPdopppE83Ugp3yktDilcyYdo3cf1MMK+1KS1Na2Sq
qL32ixAa5+ZIYXM1Iot6W4/xVRz4Y0Z+ATxn4TQkF5eUs1bSpRQt777GIiOts72cUavZf2q6LPKQ
qSCIatLEVmwu3/6fU0E+0cYnIvBoGDobgtcZ4zYCUr1TqNm3xCOv6F6ylnkut5Mq0ElVu60dj3Ej
+FrQUIY6qow46VWJEY9u0OYy7Jz8wZNqxaSMoD9FosidIdvHjHnp05dhhD6VLdV4lSIGfDRZV/b0
4YVx4qv33tKgZccz1jlQb1bmooeMgXTf4n6nOFTxU8Ecb4oS9TMIJjyxiQ17DlbSFwPNQeGwLkTK
09y3ZT2BRh+Ik2NirWzmzjw77qOExzlS4g152LzeNq0GJZQfo9bjP9yq2SMMhRLYGH01dprqRar6
9jRH9PJ9fheukTEEszQkqzGT/EGc2hsVUyv1hm9uhqBHhg2LV+P9J8ScBNJzAwgaHE5OvbM+6PdT
Z5TW4YUr7OMWDgO1QV+o/REn26rPk0tHvK784PO00JYOtnwJS50B4ESLTvrIR5pRQ1Uu9e7ToN9E
McyZh2JIDKjNLlfrOnv5JPq2r4l0+WuWkUXkIiBwIOU+oZf6EU3+5HujJrdDI4mPmTLXT3W+LL+w
WZ3qOPVu0qD8nRDIaSkw1fZRqiR3sYMjBZffZQT9qdM/ZhzQLetOMZ8XHFz5Em0j8miafF360wvU
e9tUKl36chKTy8zi6O/y/IbDOYlsLycYsZk9btPBr12R4BjxEAd5DVl6U2k4+lzLVjrI3GXoYzwB
wT/EZuzLvQDOKYImjT+ZaVcVjBqxRdtm16hDdhOguYYTqeBPhtHEcxA1RkOYNql2ThCzNOniWqvE
xWSia0qRHx0haIuHWPhMAJPiaAMvM1kX7nTkNPSfKAOdgrz+oxKfmaSUpIgIG3JH4+iU8sxIru94
yXTe57xsCqZtjWf3jV0vdbQIjIalX0BdFqnjNaUKlWyzIjpQCH+NihJjLff43xrN+MZZyr08fH+t
dwO1fU/H4qeVqiTnaMSFtM20GIUVp2UfhMKGHu/rLrVKS/0R7Hm2HpzijOgusrgwqPZcv9zTldTW
EkZNKgyAQlZoFl3bBQykI/M/qAuzkkRgQlBV3+H+VGuBs9gJ7SWupA33J9iuYBRLns8k2NhGAOKA
EG1Pctg+AmmPPM2vhX4hLqBK4rXIMLEfCjF3bj1qkrqOAvunsQDLcrRGzffodrbCDoBcsVKoSv1n
eBEFPTm/wWzlxTL0V9JQx1GkyvYzmQ7EF+nXBsGbvQtqlNgRKUqxeOFle7/65vSA8zsu9At8A+ye
ueIMUvBOwNMaJczn2itI7+y2X1EscQ4vPVgKq8Gb2F28klIk8TANT6k+UlggWFhOetfdYwlavUxl
fi+H0pthrvNesLKhlwedxobgJ975oAphZ6FD6Z83MnIaYa50Ru2SWAJ6BqHUwbahTyZDmLKBS3sV
AWXYVMvdsPocZXQuIpeRw+7IJdafSYRaChzCwFx89kSSBMrqoRoMF5U/pCUgV5ILAGHOdzyXzSRf
PiMPx1IooB80R98y4vBeiKox3k1x4cMHASdkVMVNr8aAg/vmNiXFizDO2ZNvWEbhWmQpzm6KIKrt
Lf6SEsmY+L+n4+J0FeLXwNg1b1CSzDPt0VKbtoXe6EobIpTrUUKp4Uxl5mdX/mBhkOeTHmqKfYGG
JOnza5s03b1vE+3TDV0UZbdJ2SpV+RZ/LB9LYblTO31jPDMW1IKVLiwPPIY0VLFHoR3+xs62PMLj
dyWu+VFKLysyHN9smj6pqA5ggVeDnl2xGIt196A802O8E92QYrlczOtOZgDZ4r4L7Ve0bHaZsaRy
auzT5Ros+mBbPaK69yk9cR/u1JqD9w0TudfWSmzLx9OlDbbuqtcqROOJAbYiS7rYnWExo5tjoaxp
Lr6Ls3yUolfdkJADkMRDKkq4ZIDlUHoCAZ2v40Fi81dDJDUln3jNtvxtdaiIwMSdl8FKoVBIWU35
GQ8i1bpy37WdN9fZY+pMEOcVrJdlM8nhdM4BYB/NjsHL9DwRPJGZ05Tqn44fUEIwqb8YzFNgMfWx
7HSGH+oEgqDUXDrB4Hn/NC7FArAzrKsKFKnfCwDlpEy+YieReDFwiOHfeicXOgssOejpdbtmZz4x
eetx1wubth8Y1gnvhehD8+vceMgRj4Z6xb2xPum53uYx59zSmD0dg2+9oN2L1kNs88x1+aZeLkO+
N2ZBxi4fyCNN8/1iqIUjqFDoN6ggNK3hetMmsYugUEy0GmwoGrHj5k5AaaC3xUt4GyetxS91+dJf
9z0Srqe1pkxKyfetZ6t1m/XWaLzPU4FP5f8STxNuvPKtgUI3Mu1Vo2+v6A4ansTkVMbwWdRKVuKZ
S7IbCg1Ln8ZZL+eseQc/nlfKmkAkBUfAD5azVqtJOUDsle7UFY8hTcxLBO5TDqDTxS30aZjLZYrE
PKADrW9xUccbhHjXZGaJRlmYuO2OWFWxRifavQH4l5O6tOQ8hxiu1baMRMhSGIb13FOAy9lOxOjT
UHYZzaJ2YUhv3Iy1iPQouD3x1+wBMGrVXCtBmrkdHBD278zV+N+YcQOhnRaJ57l4YTDpuHwfdJKh
/VeqnAShpwHqz4ydrcYrDRCW/xjzw5cnFJAbWLKyQtBPlJEX61jH3656F9OhLsoD7/6a0X1jsIzH
RPoMTRh0E5iUlcc7z3nfy7BeFZ/k3JOnDbJI39uDv64WeaR+vd3krQ4f/U91Y8Nx3cZasIjfGfhq
fqSOoqkvOdPqmK6oYWImoEMPNFIg7Edzn4m08lAaE21VwC83Xo0vaTgoAuTNQLeIs+TfzveieAlL
h59acFNgNyZiKyZVGxzwWhYxxzu8eIFbRbwuDKOYYJT5S2zVABsrJCIt5ezw09a5ftsXuFHdbTWY
N7o0jxtv2RErSE7dRyAL8Dz1q5nlNitMhX0outUgQZpNj2kIOQIdtfaPKp3reF8wsdzWcf+t8Q2C
D+UKUp6QwtnTFbY3KpftHuZqbjgZVFSve+MpNiUG9NQADAZijqTr/hVGYXRAvqGlNzfX3ga1mp9r
TSJFnSNAr32CqzK6cN6QF262awtpnBF2YvWN718c1UPacJO/Dp8yyRXXmoSkLCPhvYDXQ/90GrZA
AlvIHiFeHKgBiwE9UHGCc+uTZWoXBdgUd44U/vvJV5vEcKJYQBi4c84ELjlJpxOI57s/XtZOHW8J
SscLfhaxJOJklA46u5hW/P7c8ibuwn5Dsj4/RBDa83VDkVom3A/eJKRzsss4PEv43Z2O3Lk4qvT/
XnS0dKgKEF4Zl8J4AZd8Kpp/QQfB729t49jHGCl4TMU3rXZoM8qVD07AmRTdXoiG+bR1kgOqYal+
73FeLh5VwY5c6VewEpF/Bk/8XcQKv3/fR1CVYdd+SSb/Tm6tm7u87slbTno1wfYARr2/hfbQ2f3t
L9EuUW4oIpQ70YnsfOiYZOtEQcq3Tm92Ovgr0GcaXXrs1WpvZkZlpQ81xonl2imOQuHv5gouvvzD
kv1U+0+iuCAVH2p05TDuvqzULU8+4TpZXWr0paGb00MN4XCW/JM+c6ajEhnC0C5r7uFERjSczvr7
HDV1QKzmQyukqnna8X/SviTtcsmk0IBNMLu3S75VzHTJSeR8ZUZQ2RMsu2ZfqNjFh5rxoS7v27E1
X+v31oYfCDcAZRhM+IZxsT6euhoU0x6+7EW89YMPXwkDlkbsPCdsNHMVX3P4p4N2iRQOPEP2740G
8ke3mLyKofsYqnG4OBrMZm26XmXrRUA7cAKhewAfZ3krf70QfLlYb+eth+1iftvBhknRrK+MRlqf
zhaIuXGoKJhL/6CeMocP2g+IDblnlLNCl5F1rA1lPIfskIH+y5ujY+Ludz95zhql7pA/oFH4c97V
QdGGdFkpgYA8haKB6iXBEEjkDLpnVAtj6rPv4ShOJ3E/5Ku/3u7g9bz9ETHeslyouCJf6T0Bt2cS
rHmtoDvoArElgEGYuNL9UKQSAUhGwdDZKFruj29d4u87nh/smzoljpv3FcO4jlcEcH3Ton4NVIfn
xR8d7kBnjCVT63vj0ITD2e7F0KOO6m1gjjHv8o5zoU8l1M8qowT3O9rRsH39qx1FFnNjQssCfRIA
DbUETnW1pwfdxixN5ELMm/lbiFO1110DSPNOHgvtfV0pC43pEcyg57oXwooPUbK+UYIKJm8z5B+R
sqdq8FHgUfvtyPEDbE2ZhsV+paJxOiK6zvLRU+tE20Yw2qjDiaGWxc+K69mh/fPSfQt1Hy4q5WFP
2bYqlO3nX0fwJbDbgP51Zxcd4eUrtbno/YKCGuWI4URbpSp7HX8h7sF45/pFqmy6uCe81shAFRtb
YN+9F8eb50gaJ0fTG6SmlMia6wNRWxhg21bBrOdP9id0XVav1vbrtH0x1HvxajMQKekrCkt7bMQF
ydY88MYCRmhUaZ3kN+uvs/4Ik5mGDETbU6PHqezlZ6HSGYYdpCAKlsL2S7uge7hEmSqA47SaoOE3
riSFqK0hJG2sb/zp1b/qxzphYvjgxpvJuZsMvckLzXyThtC6VojWzYaabchFm776yj4pX0J9mawW
K/Sl4xMAwK63LDyIQJGx9ISQnvBpbRhcykoa+6RwNg5wz1w/ANsJbicjfwlDdnpvDQAwf4FD4Oyr
En8aGaGSY5yw4V0+pmWY/5oDY6xThkRT3NHG1+8cprqSCX2a2lvUbVOlXG/gvpawFmxqUxgnfWMf
gSTK8xO+YoGtgte/Yq5NM4qcY4lhmlB01H1tIFAxnFXzXmQ7mK1pj0yrWEpZ50NPDuvXbG35MALy
BaLCBbQL6H2OGAXDmpXYgDQjUb60MZZI+pK9BWNZFxKTCDY/e2KqH0d5+qnT6u483Op4ZS93t3Ad
F2N0XYr5yrE/EXnVy6fVb14twsQpYYZGLx53EXuZ1ZST3dbzlzh9UyGNpOWxeWD/MwhddyNPTRph
eSZS4Aryn7o8Zn4q9AiAJ43b2l0wa+H8OQkQbl4ZUjzrL3nWwHqdimsb3626PHY8CkNEKCefc7Vn
B5BqDABMRmHs3KuvZ/3tgJHGXguYDvhYK4d8SOz3i4WL10wiT2KwdufViGSh251qdch1vIdsotF3
093UJexbdEYwqb0JLuEkPsKQT65Ex5uZf/j0fYHv8EregPSR5f3is0vryeHt7KPbClSvEbw3GK/i
nT+Q4FRzE+4DLQ9W/d/qMoYLH/zwCxiL4bfH9rg3eGnXMMhFuRtzMe8+6glSASrPVxRH7etvW9wQ
Q3IvBUWDhCnzw8eNSzTOshyRWI/iAcGokDW4kWjnOE3lSCFgx0TICpa0IqUxM2ZmbXLONJ1Zjxk2
Wqs9gCKjUPIh0kqY0SfsnNCcMFuxXhdvCpai5WIVTfr+MCLLAy8Z9o7oygUUGGJkLuno8wS71G3o
bbjb7GFA9hp4fhoBJgrsMOpcGHfzTH9yhNS1MYRzIlXLtLhJISdgKSXjTsMuJw4d2UA0O0aDRYFY
yVc5QkEGnwMGfJ8jWzotPRAvAcxl5uS0V3zc4hEYJgy+/0PtOXi3bwQng4VBL0xujCE+8emfzHvG
IByxM9t8FUcEKab7L8oURpLwlxQ/7XSA160mrxx4t6UB0Alb1/oOeinh3kiNSuqu4DWaMsCr9zAx
qKdG5P2uh/SA2zG9L8NEdayPwHt2zu6jBbeFEsg8aO7vfFwKLxX5XFakL7zuu5w6ka9gGn/UC9YC
Yljq11rQm1utAJ4MAfaxX4l1Uq6EQ8Z7j4zbNkbDSJu4lyYzYql+J0TIVq9eDxuV1DgIybft0tCS
b23UdfD6FarXPdF10+ex9JSjMRd5VMKamrPiqTwG19dOpxo1HTRTnQITjiQh5QUE6X5hVQBgwhNT
DBOAz0cMyanSHyXe1mX/8y4Wod8IizT3SszPUMVDROC4tZTCIiirNCd9XHM65MMXTqh+ho0bxfC4
KGqUXVQci7a0YpeRqTILfCyTyWKS3H/tYEVXQ1B+Djre28FgbQMXkt1/hQLuzcRl2iokI9EKMKtV
cnLXiahS9wuiepOh8XpY0BQYxe0a8sH0OizNmZpz7+QBFCBWCDCaGJml6VlNXJ3VrTYC+EBQEewX
/4AMO0zQR8aR+vqQ048/h5SGx8VWzcFWxhwP8LbvFCBdksVZv2BiSCRlRLU71a8sau9ofr1XE4aa
4KDoNFRK8163o8iBUFQzoI4LGEOpgf79TilJMD/c2IpHbyEN7LR07Q4rWi7hRfAR9Ea7K6mQg5s6
1YrKsv9SG48Wyi+hh9hoLsL8+/jiqwlyhvylSOhMnM3ZG4bZLreWjyXSAccveTLArVX6dlMLUd4j
McdrIfaRrAw5sysKFY+OkdOdQgzIjECiryB9W8neGCmLr5A3WsGKNm4OG4Hc9/7D2drW6pCPKdR9
GyznK9aLfvyk64jGY2lcUN7rM6T20gLEhfHO8xYBqZN9H3268ElPCUshmAw3JXIdN7tL9GqWmVWT
JLwSShfX9yHn9GRvw6LEj/XMEFcN+9WskwbiV/Dn8B/9UZsyOsNvQP1fud/nmHy6COANHKIRETwz
pB0dJDXqXX+Xk9zcZzqFFqgZ5RVSsKIeVggIrGp8u6lWnFo+YVwafE4bEWp2Mv+Qox5H4kNc0jUS
6tQHdBeozpM2VFYuhC1VNUNgVOCnXYmg9z4GMwERyWUdLHsPPJ2iJKNhCUoPfgcyERQYy8FxEr2m
OccgyonUSia63ohyxNrbycBX6dLHZ8LyUDlA3UmU/LVWN+g+VZJDWpYZNKNAxaKL85dQm8N83rcB
Y9nVsAUFG23lQdbTD0RuJWuNEiZYS5u98LauEWq59lwjuOSDhEIHAfYOrlT+YdGyHuwiG3/KFK7y
Dhep48BHiZVXZ7EfN8R2UGiIbZrdD7xTSA6mHXkYtq/4D8UxduVm7FzisQo1W3pLbdst7hpZF2BI
Yb85puz+L9eKOSUr4zjTxqL2VGeDZk7SbvuzSeEMB1PRVkr5yI1NLWEjRKhKQXucvQquJ3bxov4J
UK9n/ZlSHznhTAF+AEeWXp8YaMDFzEtZKmhgq6Mgld1qu8kF1kbJITn+oVvjVFOSDjWs0PcvfbbL
TvIEWvY4tQ2N9xMXkqP0SyGa8V9/pKvB/4pWRhdAiyUqF0S902tR5SNm9CxEM/6aq0Kxo7lvBBsr
iz7JmeofApfNZTiflG9EusCZ7fRsNDsa9dL9YYniYQr9j016WZ5likEXJAkapt0spuhVeXTikbev
hqMiddupGSf7Vyk23D+qMomcjkMF13yD3+GmC1feme6PzbU6TnsI+MY7yVdigng1YYr4Bm5vcxMn
BbXabwSMdg1+oWZs2pZ88coyQ/QslNGkX1v7Wf3C27K8tGHdY5rZrYWGbooFkJ99Yj5aeU+QgctI
D6fhyfzd0Pe5oe0269BJ4sk8MEAbLjXd603S1titLXGKHhBJcuAVPI6kgE5PNRTDbp0s8Agy4QBE
8iWWZoMnB7us8ZFtE7C8qMh+qE0jwe0TsuNlie2aAi1ssGdPIPbcKGnUSPRH1Gxwsw5PWKAr9Rkn
zD/I3Ops6p9gRDOM2KyIkxBpmsBRAN5m5RxT1CdbCevQ7lZN13MkUX0Juj15m8du6qJHpre4X6ix
+OI3Aa+mRpZ01fmd+zZFpbydUtShp2WJAycoCXr4oRGbhKrkGpyeSmtfR+4LfQNQpzYvHyOH0ajS
UH/CzX84TAxoY8koCyQpdCrMZrBSOCcSQyMRr58HPfzgk390jd9QNc3brUwDWACRv9VjprPGPXup
fx3/M2QOAFRsPIqPjTraMD5O8WQzPl0oaq+h3Z0CUi1rO7lnIXA3+t7BQXRToSOYylC8MjRVk0Or
T8MBR3hxofRNO9da3On7N7vu8+fLqL0VNYk0n58dKGrSd2goquQKoyRS4ndupmRQtyHhwsOZM6d9
GWevYRoGyjVZspMv5GjT2yOkxlG6kXRu4D/SeBTSvNFjgHXbn8oY/U5C4ZjMHniiOOcTnVMFr4di
quD+GDp2gZm8FvPeIvzBBBfrLRDJ+APZkEWTt2EltCfq47VhU0m4e2d+eCrw0Ci6i9WxevZlO12B
ULNjdNqvXLhy0aIs/A6Ylk78ZrRqYil9UfPGMSlqMQoYiF7vWl6M62KjhIxV43ajYSYSZkucVJmU
aNR6nHQf8FlG7YBhGCMkYRi1Qo1M/fZkOhZclAo8ZyPO8pgmFUD8J5lqTD/F/nlRcoH83gn00IeA
b7OTiXfTq7PZjkBoShlqWm5uwWixhNjy1mHFJFvdALtFhTKwyTRcYySK836khrpckz0lA96Qe0CD
8OdjOYsWQ5X9AHib+APWxdsZXCOdZd/eSl0Iuage3ZRyZBUdnVjMvrTjMr8m6H/C3suD+JCqb02u
yF8SIo9xUZzKiy04RSIgn2u9WOA36GPUIKTXO3oIMpYmhAt1fF5wzb6oBN/rpBGKdy44DFwLlpxo
NwbNNbwuK5zjTOcKuaternPAQK7Jwn9NP4mFeVI8FEa9eb6N/vEN7JjU/JkNCh6jMfUQlncrXeNu
b6cCgNrVrU59hCQogTVc1QS5a3D/CFZsy3sNCXgiaswHVsG+NKvbv/R+QkcpQlAJB8F6NX4Htz1Z
zuS9Kue7mMv03k2o4rWQ9c1chRV4rEkPFCKIPYaDsM4yXz9dasVjoBiRCXNNq6mVtcC6rcqFcIDb
LlBqLUFsydAg4ID3vGCRfe96YZr/TpZhZ2TIMcjaY8I0c++oY069s8lKnOZCcjthYJ5vB7XJsNw6
`protect end_protected
