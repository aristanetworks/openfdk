--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
iQ6HLmEeAOT53hNdxPECLJfK/YMJC8OPhh9VVCBW48154DuslmI0XCrv0HaCvTfWtmYgspCpTXCB
LszkRBFWnNozGtUGuZizad5MM2Nq0xiU1rUjDKU+f2Uz3Cl63NXzGSJgToPJbfpkiK/iH1q/4w9h
6gX2D0JHrmw5BU+TGyl8ALk/KPQv2d2qC7urb3EZ+z4s/PShujZLrrvVkSb5vH3WLFSXv7VKF9Xk
I70JGUSjTAMEUtQSY7dTUjAVVkIHPEawaajFgQBs5iaoGHihkyRxH5qsmmcyccMOFA+bDP4O0/Ov
DrHNBs21gcN+E1F1Gej3sC1ut6SiNHOMVaazYQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="UEovArl+lv1jmEIudwoMq6ZExH9NkveSO7biWSBHHMo="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
jQBUfjNX/j4cOLv+SnQjb155QLA2CMVEm3du4CQOWDq3AuIaTicbdrj0A8saCCQ2TQUGrFOyesyG
8t1XOdFUUyOKXw9JjpgDsU8NMdjUn7OQJFN/WltmrS/Ynz/NSaCbmsmhLyZQrKGmNFXL9WFxNx+k
2UTnQVlf0beuZZugCgpingfrVtNDZioqUuFLVVgY0K5nlW+gDUt3DVQXCMziSD6qpLfRWZSBePRU
ndtLDI3vL6ZDI/Ng5BXkMR3dsu3P5vznro1RlfYGNHcyeNtYt9P1yfnxSqPCZle8x9DWvY37iJpe
pWZqYUx+rBK04bxI6/Q68ABNeYA76Qfshv2mIA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="hHoPNA78+OpgCzAyDPbc+WwqxxOrlGnNTll/d3HxeK0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
2pC6253s+fGMxlnXwng87xC4xgeZf8/f+ebSZWZ9wVPN3llbUqp+R8+karNAMQcnVxlqWHYMRD67
+AYuV7Gd1+lfYS6Fp2nGjBvnDOKXoX6dTGfm/4Q+zveLENmH49hQB9QUkOmV+kQ7TVCwEo0WL+37
mZZh232xBL4QOD3j0yIDOK6g/UNqJNj57SPi+AifxH3+igvVEliiZ7FB4cX6vE+6H6rBQacmtJZk
NIQlAwv2K85NVONas8bElLkoCdOWhHLy4goaq4um0qRjCsKRQYTbwNHYzy9E3CyjspOdKGCSqKzu
VCaZXvgvAINDe7RNTGn7O2yzyTEERMbs+fpHEuIL3vxKoi320Kdn3LPBuBobMwfXXSRGhR0TNM/+
MTLVNUu0xD6ZjpWI05MY/dVmccZru07hFFrhmTbIiDb1Mj6gEjzOxYlioqFXAm+MqV9wPkas4+iP
idEu4L6YT/JP9A5HGR48O89vlJMZ7iyGFlIwcBKKsV7mQqQRjcAu2qoWT2a+p7b0x/xUPJuSW9sx
w940lER4zevpWaZquE+cpomRNGdEQnimC2KObG7HsgMTZdXh4LVqo0srJXxYi+DgFeMFVPW6sWUK
dABzq1r2UW/kPMp0vU5qyuZPMmB8wNaHPguqAlFhRXby557szruLP7trW88YAl5vU1y/IvE3TPpD
Uxox1R36I1afPh3lCg6wHhrC/t/2GlkzpUs7n3t5TvOesQl+BKOo0d/OFB29Phusyt40ugig4hNS
rQu4r1NupE3agecjG0i7hwN4SvmGDHSGzk3pgmMrPw+enEo7kesRJKY2SrcGQhfG0JUIAcuy30Xa
jOtmrVflwm28tSx1NgiabOEJUmrgYY2WcpdZamaZtzSr44tZc0XPFTin8UogzfLVf4cqGfm6olKK
+I1KEVYpvLlOXxK/m73jZzkh48Oerj5Md8gS72FY2IXCHE3/ls3p96JMbjMahWYE1uXX6BCtOCMm
9FRqTYNvyIDuxwpVObGSIMUZK1G/i3cqvEdna2rzxlqfotReqRLLz7f50Ikp3IUIADNU6eXdEj7J
rXDA6sK3sqs7R6KcuBPwFwaj+xaJ9UUBWJGMvU4Z3TTTaU08CkAPX0eCRNR+YlhfaabR026XISpe
j4yGEMBAMQRIJE9eGJ8YccxDcnJWFdPbNkT3rQL3y5pSmb4y9nboV3V29vY6nsElMLlPoGCshToG
TPjkCXwGw8uvVN6SM+8sWMkGbeqUrDmshJSWeHAE8BZktiZIbclphCR9xyR1l0AzVGsNXHTeUFaq
vTYVjg4p0e2UFQfbN4+znvxZ7YWMcKoPg6Uoh9DdCqBTUoEt2cO64wqwSYU/7Jj+HHvkvwezYpQ7
oDpvQstvsfaNmeZdEQOG1Elr0gnKreHKwSTuRGBiZCPVyaEq+W/6+R3wy85nXvvbslUr3zyGpbi+
OAeFFJaDMOc+J6e31wA3fsvJpeSrh8ut1UBjtjBOjPovH0titJS615wsDhWlQufcl3WeUDZbSqoW
OjXPIR4Jf70dugDieD3nKAF7uzEGCIDo0kuFKYKGgPI5HFDH1sUt0KHEtLDbPrbyz4Z50/SaOO2q
iq/fdgJ6L61LqvhVX6Gj+WtdfhUz+DYgMEl9lXfOLkwX+R5tRFKRndWp9/3iXnKblg/8K0yfKdIe
eS9IZ5wrvxeumbfhBJBwzUXmnnk3cYOrOsbvB33b57LDpbrWJqd0df8kwzWJIPKAghQZdMuvJqER
LzBSuxuSKgF0nRxXjibQ+gZsIJg8/Olnqa4apLVjLXQgBtK8WbCxUmlhrggUx79VyDpmo1bPnN7z
9pz4SmXJZVbTEtNO0W7VBy+v96xnBZMZtgAqZiCaexoL+JDVn3qABwc6woG8IBXBhgobYdx9mWjo
gQLCH0XCZqfjWRTvzUuCOhluwV33JbYv7Htn+i2FmUw2EP8V51vDIXFXdJPBjl3g92I3FXoII1DS
CE0vUam6xURlwDip2FROqyFyoGA+QOHfinT7/ITOqTnYfZpXIEU4FfgUs+2kgBREp7i/C9pxle5E
tesT+BEus8a6wamcFqbWCilowpMyNgO2ApqF4GZkvdbl0+9t14sOJnAx+nlHiKFnJoqLFveTSTgy
dh4cfQ+7gRQ/s9ohHZCCNJVDBJrJGRQca49HCtJQtkuHAk5+wQdR0zvgkfflAxcL3ej3k+b+wNDD
P7hp08VHhScwkHglvTBquTiK90Eu2twBoH0n46H70XnXwgoEsOSV5syIiLbV73VtS/rC/j/YkH5Y
PcJBUn347T+vmvfWBns7G/NgnbvY1FJF/2cnFvhYov/OubCb+4behJWICT3WR67EJdmQsblLMTW2
TLPfDc6QprzyJ+tN2N7y/hKa9WPr+fYUvM/bItBq6ytmmQcUwIZ6S/4ZrD/VnUnsDZ5S5TzrX26e
GT0dpb1SGqMCaOltJK7M2B70BPkWkc788MLB3QIZx//AOnSfpla8dQTOSEHbKtqOnJ57EuR0T+aY
dLdj8m1DZl1BHBzNi2rPwT30JByvtTvY3Fpbsm2wnglitASVKex5whihr/X4QGkpkX+wueHYfadH
w07vZZNjO2rPvhehlQXGgMeWRIShoBWfEzNnXyXV+KkGeHksNPg3vWK/lpJ+VUClbh6Ty6DOrPO0
3uE45wqOmTZOHNB61JgjACnHqnKxNFYIDBnBOtDTP7NTGOS5aS3xJuZUS/R7GmVwuDD/SzZZ+n/Y
DMfsbhuzDs/L61pR343NVO+wHCQo64nIlNl+jwGORZe7u3QgcsGiJLDuohrb0WSVdeLfR+4YVmGY
31wvP/CyxcHKvjuwcuT3Ol8xH34m0KtVsYYUOQSoCSWxgxlomnQAriheqljSZ3m2rOgKUv9Qubi7
BAbn3n1ENU2bdYtPrttfxWRdOXmKQ9KbJ/wci9RfgHdhZbg7ZJSyALGV3eeqW3Kuw3vr2tR8/KAv
jHgqhofojcqotmJkUBAPUplM+VskeVovDW5dOqDONjWlpH648Op4sKeQApCZYJQ9/6e7Dqt9SmK8
OXdmzrMWFhn/k+kXGkb9ZPztlJ3dzFOsLICpbZKvuyWaZldgKYfEVmWI20EY+KK0EeD7c2aPGoKI
3qIUrBpQrJxpGAfix4AasB/67xdQ1knsvhvjbCLB18/U7Fj2UChTNmonzfMIB8O4x3pkyB9mgN5e
VRDg8BY/Rmht+fuh+BLRNFWaufczjN+TbMCpp9yGrlz5qE7rQVdiQZO3ASzhgo6X0y5KSlkJyiTw
U4kNn2eJCDDAcEMBiIZv4UxEwHS5GDB8oaHvdLB1jDEwHtQBzVyvU74kU0eNg4QPNVWHMV2+funX
rSxcaKWwsQBrsV7SfKQHIu+UWIxWiRwlpg6DM7RMslH2L3/uOH+uZ53I8ekLuU6/+0Dgq4XpR8x9
ve9K1AfBE5hcXps0fEDRkk6BPuNpnBf0TuPBRlbFTKxBbtCtfmbxmJ5i8A9W+GUaiJ4CoqeQFH03
XKTvmflqCjq0QwuSWxG3+bSvI5XqzmhCnPOJmPFJMY8NJ4f5/IMZ2mrwO/y8d+VWQHFT4iyOu6f5
qxM09uViZ1fvKxLE+Da9xx8aqRcAOHXEZ03VyQ8dV6Sma5x+S7VSnwcbbctWLpRQXeWYW45aapz6
wHYg9yu1LuSXlgjguCfVmYR8/XiFFOf568QgCutwGtVlp3bZIS63oe+C5d6hggJcihF50C5wnv12
EOP3xZMoRaG7+YK9BDKje0DrurLOI1GKGOL1bcVBhbkOk21awTk1p01ipSslejPAM88/Ya7Ppijx
NCyYbS7Rtwy4tIOd09S3U8zlCywERyUONa9mPjOBg8F6YaAWgCnUz7ATZrOqSFeLNUPF07xr/UmP
l/de0+pCslfHh4IcUl+ubU9nYjDmeVqZWEa9AzAS+1pqwhn4AmTe4CtzcMd/Dt0rMOwn2xh8Amrc
3UUBiGnUky8jJAk9wddM105TAcwEoQeKDJdwFBxoJNP735aHsPiF2Z1okPAowyASN/3JAvkzGfIk
27b5gUiEFoUv/nohwbZkgiFVwlNEfiorYhU5lmvh4/2OC165eZ/ZxArzbCyZFSAwhDVRM63Lt/JH
mLBLLTfvopcwquBkKX7xyZU4fkA0XC5kgIgpBfunqt9ZtX3w8mFbYOnPZlX+DFvvezxaq9NIGTig
ifmNJXZJBJihAUgegDjsZVk7pA2z0aolpaHoegyqYilAupXPgN6lk/JpI8BofSECZxdO9ysH6i9m
OLy81HnQ510/ReFzm844BLdKU0fYcsCjRpplRHOJB0vrX3gUFdtmztibgcTzWmo94pUtr7MprfPE
AOPuKhoHGzWgJ5yxYBrXby+FNOzluUx644KyRHZNIOGSekzgLJQsTbW3kBqXQPNNHP76SL+/lfyf
ipt1WoH43rhQ8D4M7s2ho5+c0hgJV1/u6Us+W3Es+UaaSgWEX5KPXzl6TFZ4woySkI6+6hfVcIOy
BgyQKP8IlpSmcPFZUwQPxUCARUj/MI8eJTL6zgzoDcKVz8/5QByNgijyrj4xxoHaPNyAaSB1peme
AnHl4AWZdS2nQ1vSkqcZ71QyDAVHIbyXxurERFygGeX3yUC88hhaVTyBUfEtZIeepD83Nz4vaURP
1IBsDf9Rc6jP/WKRyh+/DS2WfiBkQTQym/5maOVak4FQPCe8pGgBxbujkWNX8H/eOyeXDiR855Ij
gts6cLXjPFkrrRMI0MNKZJsLebjvSYNF4vJX9pS2K/J5We42zRBdhj+DyO2EILeS1WC06HmAqtp8
MkG4Cdb3mdJ/gqHp8r5u7QwjYIMw2mWftNfokqyPKz4x18JMWYXvmOre/SpJBhl62L9DBFsPp+bd
seIpPWTytNAeMHeN+tF7VzjUiOVzW2SOGdS2ND/18at8/YfNXi4wxIbXGTpCkiFcqt9IWr1QEivo
BXrfklnxaV05Y09LBPB98EY07qkadY03ZP99eConabwkd8nXN+7fWc+5xCTfGAB4qOshGfrjFTVA
QoiVYK+4TjaHvgx5A9wJyHoq+TEXBOnRWm5lm9i/MNPg0To6+0qrH96mypj1TkybHzbTY812ReSj
E3DdLcYOM3XM9vR199KPOsmDscMrXgsSRvXfG4Kfr8Oty89TGp5XKX4KLyJmRoy6wyZXtC9brB7M
5Vwgzq+Z3jkSKTvG4WijSpgJqzRw7ay5qeUHwjoPbj0oRuFMUxNKqOEIlmFXKgm8Rdza+ksw79O+
ky5Oq8KS/xmMAAgQ6I9kKMgElJW1/Zu939ZGKqKT7qXr4Ouo8Z1inbDT43yUKsN8cDiCV3k5XxYC
jm+ClhYvxNgXPqIP/82ruIZ512yRncNnZj1Phl/qvuxZKC4vH+cT/8Ay1JLYoj72SSjxseRJPTb9
TerrlVFEETk9AyWYJYGPFPTQTyqhMxaPpkqO45jSGBSdifxpSMkLznKzai1HlK5N1rpLuo836843
WF+/LmS0FJkn07Cyhk+3F2EAexscDgu4sPChuXWcmkiVy+JadrOylkiheeLMir1HaEt8bGe1ePdd
lyDRBQsM0g0SRYsqUKXr3hwJi0akKIuhUMIZ0k4DJSeVjxcmLuHXEaNr83NteGAi9uNCANKBJy9+
nxou56jMD3iYYBvNFl8VZ/ike2TOenvaqVJeKTGho2Krez3jYSa0S/rKSW+K37fRtTrk3xQI+q4b
QZ7agZU7cF0NcCQzuhEbcx9adnB4mSNOTVRILbnE6Loo6ht1EtRTuV8fmVXVeCUPV589XAVgRJJB
4Fsd6T5HxiN2hglR4oMmJD1nQsLkSW3jeg+QcYK1yVbMihRH1OIuI0hZWqB7zggJxJHbbBzNw1lC
Cv19AMZNoCXeEXTbMwzZfiet3MA6kqf8pq5ZZYr3vz5mRrbvXWQfa/FovpYe1lGrBv1vWg3gyRzZ
dTXglcfuxqQY2jIuuZUcZbLcs58KXk0MyoccYuaGPidXxSoTrrsLe4mwy3duVPBf0hHV5Z/ar2q5
nwC9QqQtJccPC5mmxedF5HhNMOHBP7JVA+CBA/wU9FnURDyv8K3EiXfp9R6p2ZFJQCNKsbG4Z/dz
CpqWfW4p4wCoyKoQZ3bpiYXDdRMeqbA53XVVY0ccMAuuI/icz7mUXEwktOCiQ8WE773EwBrYBuZF
O2VE2hMxk++QaCVkwBFDDueRk8Dk+qSlmaloKQ8E4ZQYKIL345hDrRp0HajrVj0Vv3BT7AGsM+IZ
NAYbvwNwZI+xz79wiXkebUzS7YZH0zqvRNwhpqFEEXtKkYe0g06XmNR+LYOThloCJKBXIXkmwLRl
RJgSlaHFP9k3eDH6obNUV8j+VwzKXoYgT9wy3wGGhukZBkMFCdai1HWGSlY/a2O36XAj6doIUNu2
np6s06o0dgyKgbsV6/o9yJCveofYC8AIiySEGEu1tHxVqiHH4U+fG88IkallI6US0Z+At5FszP6N
wYquf6CBoNmowiuaooTuMTWnltWwR5UGBl5Ouhqsusk9xEJZEnBgo12AK6tD23DSky2qcgrXfIZk
AhwSveAuH92PPZurX8EbOZJ4sKcygYAgcH2mT9DrBxN/DnhvAHf6MVLFcSzAt5UnZGIuEMRv5ePd
obiMHeyAsIjdH48oyJSM3S5qh/sUvKKrh6wKyOvNbb8DOT7Jg7EnkFsk+nTZWaZgCMbdjDnxvl2b
4H/nLw/kZ/aJaqFQHqofy8U5877R+DfV2zq6Mday8Ns5HOsnkXqA1dCraSm+egqpGm9wHZ4UHrlT
QxT+Asw6guvRYfMfZqk5f4f6A+MWuVKLSc9nNMQxwcv//VNowBuiYfXmLVy5vbBa/Z4RNFjZ3ja7
yxPBl/YyydEQ3FGErgi3S5+eNbPmALdLBpZH7DJvXHIY9EPuIcrGvnEOD/AHJQitE8i4wpg+6L1k
Oni5wR9Kd6/dfOlZfn+O9KcfmtBFdaqleX3tS2xiSMZBVdcbzaehf3OX1l86wNciqZ1gyZFLH7Hj
zvJZZVCApyD65TK4+sssfhDfPs/GTnKHuRwDVNa1DTMlTcjIjeRodW8Zi/JNhkypJdN7xdyHU3ZL
g/rXpWCktYa1yoU=
`protect end_protected
