--------------------------------------------------------------------------------
-- Copyright (c) 2025 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
HNk1ILmlrSj7O2W65cNvP7+batah9XYhqpd9vdnmdskMKXm+niWPdOCWy7mUTXI6TFeuqr2Jm5Nu
taHVz+HTGQz97/QGnYf0kEnJO/XnltuC4bmIwteQbNtFSTEkfOw8yAZetBRMJ7ZxgFuKSyBDgBVX
i9HkzQVWPnP2gtuKu09qnUu393JyJ59iMLMk9hpm9Fvli1rgXTDJUzdlnJNOxhGjZMeaTA1SCE0o
0vnwkq4TZg0DNCTLuEyebguZurlfuvHJ7hApf1i/HmwJoyD43vIbDM+9bqbKQblGfRNWvH7sz1Af
g7Sff7KA8Gl7qXA0szdSrZ3jJb+6qAMOt9Vbyg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="7cxMIMZ0UmdS71EjyomSC5uCM3xQfgueC6xPywJF2Dc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
oXVYiWGNwxEoiYtE6pvdhtxSzSHr8bOsL9aIUM8sQdclqlV69V//Few8aaisqTtJNZrlIgNuwP4R
fwHVT/oeqhLyGJjnopscDzmuY9sJH+YdytrNSlHSPzOn6WOfyTW7g6rxLGMqONfBGVfuZzrt3TgG
nFjjmKF6QPZZlQGfDM3nufa1nA84lpkOlDtFw4yvQxQmf/A3e9nWyaCLugBC6xYGkXeZbYAPTE98
ZDAicaG5UT5YtaloEWZHK+iNUSab5UihqI3s5KyKhoArYp0bObK7lV1EbYzzNT0GtEMuOoN7ykDX
/D/X6whpJlq2iSIR2q7AdQVTlI6aXZCZiTWrGg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="yRILSNyUuOYoHUedD/55A7FKYXSVZWMeoTsS8y5rvHg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21216)
`protect data_block
sFsNh9Yp+vsK025XsZyZty63N54ddldn3g7gD+N+WXcd+4v2G9BNSjgioPogB7RNlPF3ezepl5cw
mE6TLDHbGEeB/dhjwfoz+0M7TcO2mA2mYW1H2kSNV5KW8MAiyrTjZNXV1qN9dI0FVp/y2fWVpZOF
Ga/VUv+WxceU1D0L+2gLyY1R5nc2BlPeKXV29sbQKIwO9hhtmDQdJMc30a8C/OdgbgLaWC3f+m+x
BMGE3ZRg14oES7XJh8P3qSHqBiOXSyA8vuGgFQYlMH2byqvfRvRr4pXJksFysg8SHzyODXIzVrBV
uMhkl+WeKJpMY24jV2xpl3VE0zUaz5uYfnCd7dXBCwIW7i1iD9R7JKQlNXKJ1IeobtS6XXSbRuzM
E1BKaHEJyDepm/s4bqMfjuGLWrqeB9anU1ntrFFj2675CTGBvi5HuWmFcZGTdXILMiA49xp2nMNG
mCXSuP+Vs3vgs+2JDI3pxgOPZTxrFBeyxLXrP0AmWvjZEhvLefj2GqAUKW/wn7ptvSl2XO+mHOsG
2vSCotvILSSNDeUeMf49CCSzBlLqUvEWYRk8axGFcqoWaHjRLjcAL5Hx0fV0mcVG0fvkUojTgpCx
ZeFAG5zhlHgoxPe9EzNgbuv7aAUuI9dCxCC+o3rm0Y71s97Uce29O3Lri+6jfv6UKFMiS2tDYrtA
2FyJ/GgeIgenRacN20A2M6lCgCJjcSiXZitXcFgJYnGe7U2LjtRr657aIHsyjx7JEPRPb+uypUW6
85KAOdkj7nQXFvKiLIOnflUh0LCVsabRjuelCGsMC1TXpdNuPdMsgN/2j8CEWsRfWUpk5MZzGnVO
em4ZWNLm6Y7RikT72Xn7CAX91DEgNWXXrUNj9kUycC4ff3TpbgSk8mQQ2ZydMk66bVpCN3z1yi8X
yEdz1qtk5KqgIe4Y2I5Eqw3yR0jZ1SNekjW3+GXEZ7s1RFgLm98IYbIh30TJNuJE6+WdSw3EaSUh
fUSLMYq59BuP5ZlL9pRE3tcNifYGL4QNpMUEhI4tk+buHTil3HTCNUJ00OqFkcbuJh0YfbCqceVt
rjHUJdPBCFNS9TGnYvcl2XhZp0wMeZyW3+vTVyzCFdqcB6D7w6Ygpws6Suzk8eFgnO2+3sH08/ko
/VxqGnzECJyEuFiYODfOHaru3+ivWDLAvaydw2hCLZQTu7X4Ip8241fx6Xzik6ql75Ddb6hjl7Ov
aLItf3/9jb0lc84905GQga586e/+dkkULy0yTJC/bKgLSXM0GMWl9ryTyxUGJttzR1ZJF4ccsyaU
OpXsg3iEc49rmAabHWSrGpzBV2YwukQ7mh0wLvzW7W7KZaUomXbA+S5EfA+sUXtEJRpZUju6seap
DZdLsGbZPCY+fmPp+F8/AeDLCII1pg5BF/y0HXYKRhSvnmsfNWdj2GM3Ki3oKQ6ebyjOawRmL+ll
qRQ/r0b4GgXYBrYOLLScpyB0bv/W85SKkheAcbR8uzTU2wUCOE5tnQjW6pMz9E482E2CbW0SRBqT
oySJYoNWUfb6vx0Zz18L+mORj7t1ve95zS+yoBEnamcyNyglB+P9aqZoKEEeczqW+9G4WhV+8evz
1Q882ESLy85mWaKu5ebVTs9gipSBzTeQMvzqyjRJtLT/BKXLN8OpI7QTXvHgN1fcSb759vZfAShj
tqEoBZJXEYDV5gIb1d5WCm7kR4N33LYUMqb02wm31Vur509eP9z2kusk8+9QPsXuHbelYtnXPRJx
b37eX23CQKgUYjjl/EtMNhnginsD4Jrve5JkmkzmPaQCLuBVYX7yiqNyrzCfz8CICtYeYwyMVbjp
X0kU56+MrSgmF2/tCwpt9XntHMjw1imRd2C2tk6/i8wkI7C8Xj7P3p09FJYzy+RNNTCCxWBtgnW7
3l9rbLoqSYLU+eFC2rzTbUcGiV6vnqaRv7a/Xt/MshUkV7F1ewgs8GU+lppVDNRj7UDNN9rchDwM
ec+6vbbJCh4dna3nhsatyjyi5MV5oW72hXHHq8w571V61pfpZWUQuRFv9GYLvAx+qSCPZw+2n563
6eEcw3ZdbJiVEKJo+xh6JWu1udb5NxlZGcIf2gS+hnQuMNQmEUtm3zSk3PY9QNqxqQoM0oGP7JnK
AUV6gm7q8I6JzR58i6/SkYX+53wzlYP02TvP64fR18nES0kYUuUTUvisHv7nSE/cRJZSpTKV54d/
hQaWjKbioun7srfoKTjy7+vVa6o114Xi41frIjKatt8kkudCPD/xK25eeIAKTrUMcVo+encsJmwL
7g8d1hmIalCGyUptghj41QIYAZ5iXURGQQUgK0LsIk3DUnk87ta45L3WGlijFKTFeLWeHYpD7W2M
cE3Q6pRfZyLSarAcRqrA3z/Nrrusrbd6gIxxhHu1st/DvUoFMp3d8Fw9ChqwTqkAh9YSrnbrc0WA
9c0ZTzLPYIg8Au4d4rVfcAtvYtnHE0vj/Gsnifxq9ofw8OAtHb/ZOfEVtROwCCBw87xGMJFvRHiM
fL5YpqzTdOSmw3+L6RIHr9lNGhCQnq0hvjQ+KEPbvp6VK45ConcC1DmJ/3Le2a8M+eX79yqDrMVa
YPI+qqmkKsXJy5yMBYYMU8vnrIfHWxsBiNg8O/+MsXPWEuxzdy2pjEF0nq8o85uzzmbvUUjXk4aI
r3DycohwXbHE4dEHABnPQ8M2nDVp+rXKmVBKh/NnGxTWtFkRHEJdjGPQ8pm3075dl00uWWuXbyNg
piQ8lB9w9oq3s2fDnNVeqwRhbGfB4ZO1mzVD8iAcX+PlslgKp9Au6Uf3gCClsPxfSgJOe3SEfB+3
gVSXXHXvNoy+Na7zArbipY5L8Z8wf2IFjuDT+A5uYSeVz9HoXq30L8hGUStQbhBpoLOvuN9ocnE8
izSVyXRB4XrH38jIZtnF2pjz479EMxMYdFbwosgAZURR6lu3UGUq3/c0oigm19Yek1QJStWbxTa7
Y6N4pn0FMfRUngxq4c+zf5WUbT6BX3e270Fw0k9Xrqs5wyUlaore3mkePcjW0S36Pbc1EfxtQD/A
7iM7CtgbQ/OhfOy23ruWwp+2kSC3Nx26m+lXGfqF+GuAz8dkAJR6U1Z1SX1KKP5/rEX0QmwWu607
7iC3c7RgjAzGFopXdKJSxLpi0uFZ7bFyF1zDumC6iyEon36pRk0NexTR8SOibowsndvRU77RDDUl
F7I+YxQwhOTWkNyreWc+MwO7GMqgMc/94YtafCbAy/vUdfh3S6UWWsgBHKDlPVyVVUy5guEfzqUP
ozAdSZ3lecP2W2Rjeuo/NEZBenu+tb2/4VcU9IGpWwJw8sn0TOSzTuxlBHPBQsLAdfMH4l+dNgJ1
l7NVhU2eAZFv7GU1gNwPd9JPDzjOOmyf6TLFDkE0LsG2XqR+oss8nzqKWGqk2LCGqOuBycjbBIby
j+glojpF0T5BrLq8AoM+ABVaQE/ZGCmah2E/CNJWaXdPyGWX3V8ie6yNJ9qLHMAYPAB1JEkw0sIm
QC5+B1EDSEo1kWTMZHydfVn24KAah9fXaTUiDmXXFn2/bGuO9jW8hdNT2N38KsLJ+WrZ3EyN/4E8
ZXhJfo5tRaoCe6yuHApimcEsl667VZ2qL0t6YtyW0zqUd/9GT7uAdzbSAYvnTYonCJrG9TD2efrE
UxYRSwhAsbbhue3fk73b6EodXcMm8wcQMgHYtHRyxUzXzzwTTqfIhgY8W5eT5eICTwqMuuXR3NUf
00LO6N6GgeiwrM5Oe42Rgzczm56Ja6b5gKunbipZweVbEeyGid5LCUI5Yg+50zR02MGfk4nr7JTK
RAe9l6EMJQ/jFZoM1h9SEm+rbvA/9lLZ3W9nq9cDHk4LVHtdB1O/HW1nqUdSXLcawigylsKhgOXo
FOU5GJmmOAU9a8FezI8SEYJW8UeDU3hXgOnxxTC/16RAa4UbQoRPcEOVX1KO0Xb2ahVXOJSvG3Uq
hBDQ3xfTA9gAQVIuLVJ5oJQ7b+6U4omsbwEtPgvNluRXtV0ZrvCaPTEmQovvD9TUBJeltg2UvVKp
C7BDqBcjjkEwfbMAxA5klm7+iQkQhp8c+YPlcvSlWB9BeRDqd0/YArit0YIA4IpWT73yTEZz6dbK
eOqQCcg9Pmov4wDLYdxTsEr21Siz51wwjSejT72k3cilVV8fqmRd7PgRinGdAtI1bbVc2mETRnai
8aimEUtajMA5OKEzr0DMfFIHZFw5NW1CPoH1MrZ3XejyeTbPSJGOUSipqZDHgxoD2y1V+1KS565C
n/3SHflesEHnGO+au+TiRqYzE4SYJdQHDI/m1jIDrYBiHXacReNuIaKeca5wqAFZ6SxOptOfDhLD
YwNrjVdfAjaSnlhJzxlcnphy8G4S+0aRuudpwuSxZnpCe/MCLrBZ2r7AvasfFax8uhYYOjSw9IYb
lrYPrCpDh6wcR1GsPFMh/Zah7csBAZ6LsbbRC1iSlRX1BB/yRh2cI8nejI/DL2gUchINVr6DNgms
IbzASn5+zl3dYHjlDy9iSO7xsFyOZgNy5a7pExBU7cYsb6tLh4N9j4ZOzAelaE3KFOhNjK/FqKKF
7J58VelTEu4NDbdtAw7ifRMwfqAWCmHh36YNMliPEw9BSpm4IJCUceJfVEsqIT5cADXautOKBlQi
nAAFN3n8ndB+XF8vO3p2QsxXouRZAX9B8lpkRz5QTA4AaKtlxXmofoERc0uW5iBUE/DMhLvpdkEe
ME1pnwVdytpJzgjSumaTz0KeaTP9QQMsKF5ApqdDvNsm/esm4qjmRDqj84ZV8hUs+dy0LP7DJnNs
N4gcFRbTIV99iWylqK0iq62qeDB3xqQHC1AbPMGLblQLRACp2JwYNixZdnio6RxcjwUOizHVKofy
hgz8KM6LyPnqU01MKesjXb3O2yIvfoeCCW+t9r0ZlmvDOVbf8NGkZBTgVI66MzcbrPGqrFvUzV55
ftH8VKde/DKUbagrHkWQi3uYk/DUzIuV6E/xT2QmTVefeIv8zQ14FM4WTHRg+n7FHTGQaysGQKiQ
wDzu4cjX1ViVmh4PzYdQRJFS5WgHszXEUlpuV+xP32P1dThkYSpcTKCT0CcYrA9dQYanLaOgrT84
L2OspLpHyvf+T0E+/uJwZ/tj3JWM8aggoNsKNlB+myg8WUx1OaRGcizPDDkFT7zr1xUEJDJmU26J
q5wkDYePy4/nWJ70Cmag8dFjLKWuBrBuvyIwzUy1DCixrLk23+6hPoXMzGp2yyXKYy3BdYVBDgj/
uxcnc7LEJUi1IGCKckfKtcdLU30H6YCz6nYpaW772W3I8YtLz1MANVmB/5onZJGFc7Z9GRcXC9Mh
N080vNWhueZeRxygJ20QZm4EPN74OpMRgMMOJ3/uC0q35o9ZccsgrPJJaF5HO4xBQSw4thlGSwGb
ptJ4Ro+aPOIh9dOcy9roXH3hl/qHtjzEmsAoylRzpfhVB/KiteU1mTdACDVdyti7HqIp89oD7SXX
UmAZmbFEYJ1G5y2ybaSWUnS4rDUn+8HvGwaH7pf3UMwOfknHsQeq9wPV5pQSxd5Io4dJFozNNRgu
FHLhkaXC89UPBbYPKxONAiL79jTvigo4dpIRX62vH3Zekywb7O2Dz7rIgJORkrHFVRVQjkFdDwdS
U/2hALMmJibE4d/nzUVZJB+nD8wOW6fKFclxdbpNgrq8eBrI8/XQipq4wZb7hHuNqN2w3U7PqF66
pdiv9XB8Jgbn8d0SIH7MkjUI1uk8DXMnYcAH3cxCSoR/1GIvPeEI3GaquA+/UGA0So+id7DAUWiL
u+uzeiC37ulHaiHWBdQKU/2v4yllnsJOKnA4/UHgvqB4AMCDes793u+zfBHkuA41DMaZvgaconIv
+VG4dxdl2DjpjBRxk9lqSU7V9sqfEYoJc6o/ZAXyoi4THR2/haBTaIDrjSd5MteKFN8JQanRwGjD
3Ix2auEXo6WWzROkmdXqHCAPraDDV3RSrLpiWcqcpsLMxGrNkJ/d6XAMk6yzOsckCzwsmbxueB8q
YCQNGfXr28B+/v9zjz8ZjYD3tSUtmb7DHdo0js0yXqydnyBEdGoFQRxRNgDBTIpUrlV2dLCoeVAV
OnnWYxFnH/gduIhNKWmmUidEQkYnv4OQ4EFzHRkjNaUQW6qyPvS+63/txCqfO2JWStJCZJgkWwOr
Dwy+yAkyztZBwWJFsejTjp+3QmvDIETLpRGvW1Qm4crtQBv1UNbMrtoh9NmsXBf+PO2cEkuCdFRy
hmKFFujPw6wdFJzgu3sjE00lqUCjbJDZm9a5eiWTflehJjRrn9avJyls3xTL/Tnj/QoPq/xmPvx5
4GdPk0rJPB71ytX2fGI8P6fTPNuVJNCz5PHdeQJh0YTH3zWrLiBgJ91LWttsG50gOgMAiUXRfl9k
/KC0Lq8xL97CIgp8q8AfWzhqMQDlbSFRhpp9H48zV9S4/GiZSY5DQURtvnaHA8mHlBle+Ge/e8sQ
DPzhU+jcumvqyFwdOMOO3p5yhPuwn0AIuH5taJEFmrn0pQNGdAQG17Ip6fGjVKuh6+BNsTaICF0F
xXI3ulIcTbt28/yVenfp4HTlbURooyCruXSLV3kv0cutH1esxJ8X+JG6eq4tddlZ1ka0JPEFnSWG
6FNdW5m8CAmUPyJTMoRdpxa7GYuUEXOp1zFx+WmLS5YaVuRe4YC4MsOa8sQqR3CP5owt00lfDGga
Ydx87aCZE0hzBuxAdnkx/xRyFotnNbsTQis27BxX15fWSCE7cVkoOaCx7iPfDKn887uuEXhX/dZ/
6laKaBBnU0+V4MjrpuidCGoGLhwAiSvjhX3dIX2lut6thVWChMzFavPZEiD3Q6AMF+KUg7sPcMn9
IBym4XLyIPsG3q/0AFbtYVxjC/hdZRiyf9WTY8dWc/pSeN/Uf0NYWuKMMWB8M4ZXhNaTOrzdrOkw
SnjpfGPUpZiwZY14iZt1nE+xQHp5TOnn2fTquloGmv9tnNp4K6vX6TlEdO5kyrWFTcC9yPg0RxgP
pppPuyGb4qJTgBaEk39JvMoH8DMQE0vx5m7tNMm+NFhgNqYds1Xv+g7Px6DJGYseUtU7RjmD9Axx
LpqeA5ZDlAseW9hIFJc4ApI0H7alGdUpHdXZdfwSVr9eUGNFFclGZfH2OHj1vDZBotrngKx5a0V4
aFOUjLfevTkppVJu5SlTFcDhjSUyF+XUFqHEx5OBKJT5IF7VXYzc31fYFSrdKMmxFThFgGa5th/2
aPvuAhlvvegkut/qbYYXCComtJc0jH2UgfBBNLeeCkhd1VzsuBH/AXJ8y9teJko/TikMr2xPmlfA
cxCFkb5+goTPrEmKyeWFumJ7l51eghJTERx3ymAoOTAK7h1h2pCHKmkqL1APBh+Sz2xEaJUhfY/B
VmqdzCbrs7x26Szju9aRzPpIl9XCKaZKS9cmGPQnqieyRFYRc9IKEPF5xkpYc7EUPVYMOSw9QRi4
q56k8m3DoH0g3gwdCia+n23i+VfBbQpqQhOoOkBf74WI2eLRqGfPQ5pTU40Edv5dyXfemjzqsZyh
jMklWb5hH+l/jTEo9d8+M5BoI0UtQ/6CthKIaw/UFOpnXoOFJoP+MZQsCiFhIhAbKxrFYZszyDIF
/ICdr6SZkmv/8AYCpLYkgfaTt1rAfp5gFxaX33iIq5aRdUGBzFDPPOWT9+v+gluiRmJOW94Xjqkn
i51RCUFgsJn26RKgorjuqipTe0f0lDrgg80oAkzYM3izt1CQKpQ499UnhBT++SyQ7mRca+a19d81
YlzLpYRE+7PvEYmlf/3IvRNika5B8nGSTiGcZ8lq3cp/tgD+ztF8oxca877WjYW15BgzhSC+LVhX
M4lxqzp31NCa0PYmWhe8se+mNGKjuKe78ligHi9Wx48hX5QHpb8sWgQSP3dG6VLeK1TqOquL+z5F
sska5I/RIdNmQGOSabn9NNSOwzc9ISB9fQjO2sGYjb4GnSvPsaixd2vDmdU8mcsRXU3XEU9A7e9W
MRnAAu1pri3pBKppqV6HoWiC1zQ+/Kn6SGKeWLaTSwRbqAkZolyneIsKEbGqLJz/eleAWlHbKJfl
N7Ea6lUyMB6bQ6e+Is0/90/OSvo9c/SvY8PUiq2ySvXd9pOmgRJJmTj39y1JoN0eU5EMeggX0ckN
R+CrvIoIz+BFaANmltxgIIUM6g22omU4YcrAzIDw5FQKi9/TzokaaXmWTMA7pwwvQe7O8RnhXQjY
1E1SCernAcltSeRvqpUJJYJYyi33nUzKFQ7DcaLYCalnu9ZkZ3Ca2mYwMaiKAmijJGewAd271pMK
E1zSKqzmk/vf+JPyfwi6401iiSCHsGMrGjT+N/Zs84ZkQ57e+ek0wOTCJR3szeIzhahPwyQJXRIT
pplw/3Zg8ViasB0TBzYO/K3o7iUeqW2yLaAGJgZRT/+E96wKC3I/BVHNCKoXeDscQ1K7FYuE+iPo
yq99Y73tHkgvCMjZgWTLdPUBrkV+COpx/tOiGDdTvioOOq2t0gKl7ayvqqUGDNREkD4CHejuK25k
XEQwGjPEIR78DWoIchNq6dE2idGPAsCG8vaw7DUm2jFH9y2Q4qaaZgyuBkwcneDWAvqCZBSk7T7m
b3Pa3pOcg8xx3CmFlPBgQF8Wkt7m/oNG4jA6bec20MSFSkS/gsdPKsq2gG91vn79KMYz3GljqcS1
DPutANcATlsD+8iHtV8Eo1y9FaGePsWyadZUIecl37/EGJwpPwjvDCugdc6CAlzM/RJdMdOAcA1B
RE0bGiE3dsa86cjciUqmjS1iceV8RU4Nx5gid/tzxLQaqUxYMGWgYtx54HM8QRnlOggH7c9up1T/
zfK34n3kMeYPxCgSDlKiYudu2lEjKT0tFhXTaohG3ytW3OyLNlPBw0NEScH1UHYZuDTMT+pig3oL
jPlS2bZX5MzgPSmW/sWqlB+qDQi8e+K3vmVQvv9tP8UvxzYtJ4cTIkJyKkt32vf+9+TsrP4pU1Ts
V4NTdKDIXmu8EdvQQRUs7WBc1aYjqZW6lFnMvB5odkCDQJSxbkY1GcuAOjskYHA+csfkrwUm6bGs
tTCvnVlY8YpH0jPMD/dHbpzml4Z+TknNnrmo506f2HZVaibWqR6xJptFi5hn5GDj2kzR2fYwOM3c
/MltaiTZlmPKO/RhfHhs8bgpDZi9tPchRIIqgIq3951nv9nFl52vsc2wOqfCAOiP3ikN+bt1nKAF
SwEUfoSXJBqRjqBCOH0SZbq4chq9CHCqy8rJztXVHxmC8lQBpuUsGk8xiQEUy9PjZS0TvAgowF8/
ySvNAjtAW67WY1jDw0kFrdQGgB8GFKP2uS3Vq1jBPfCXOGyKw45Rfh7a18STW3hOdWqO3vL4IW4V
HNhQh4+QUTze23PG01t4X1336dXaYVyt6rX891X7s+DND0BF9/gbBzCLFiMvc6/+AfHAUyyWkKFf
cm6sWGmUBl2audCUuD9gEGrXo/FdIHJza1zRLPU80puiyDSvCJ08oN05Apqxj7BLDS0sZgYI2m/g
EJ0hMThxdf0IoPJjyd5Gx8p9WPr5kYT5+vVl0Abd9L0Kkt5FblV9VCrZjIenMcfFEfA6vrwuqJXf
EFEFMTcUf7REmzSVN26Kkskowyv20eWEF7uGo2vtvyMUMLBGNd2akkIG23q8mxHjIrBOAPj3ZNok
V4UPqSS/46FZnX5wulXRUvI4PzhW4BQMzmDUI/obQgSA1pG7Jld94HcsOnaO10KBMe/oQcbu9AZd
z/ARbylgE/qRWsWCY+UJoNbHWOlxUg0nitaoDNaDCX57nlC/PETerjoBUamkTNsAoGRAjlmLpm49
8wUcXJwCCNXMS5GJ6rqivUmtFmq5Fvq73yIJWgYSZ23xiiqAaBbTHV3cbJ6nmAGKK4mxgXSLdTOb
8cEWGB7PBvPeeVuwcpvO7EfY+1xH453j7MQqnym9lQHw5Szsquhzn8u2ioiXIPhubtbBBfIl4tgy
gvDtAz0yJAs9K2AgDU56D4wwhuPBM6Ld3jLcCNzMbqs3/XT6ayg3lXdE6SOwhmlCZeXuklhlvRuf
6NFYXgJJq3rhhag380xpp6zrwE6bg/5LzFtScvdmnzXFFduHJou/mc7N8LyksJDm+7aep2ENs3bh
LKEzNd9ETD1d0DMXOZS3074oHJ/eGy6urYnacjyDAknYr6ENA8WAg1bqcs7CttQaGua9Eq4TCnDy
W1yJfuWRK6O9GPx9aM9J8q3buN9vvB7TZ0a1+W0pgynm0Cp2s4UDwjVPdc4RSR+hXSjhJfyaViQK
dNhyBKTrY5N9ldnSAlj55aWnJktKJk4TFLzc7ipuHjnJvb3gFzIWns13sbNtvhqvsNRcwvFX87XQ
AX3gj5hPw6OFExHU425NafxLncbN1CG81O98W+12XYSC8MxUDYjdlCXFVgX+tyj90YXQNGpIkayO
h+OHZpxXsllgN5NdNCkQE/VcjUD41mgjuLYFMWIjSdVFuliivpB+JiuKM3h+bUiWZyD4NTp2aEF0
Yl0JtJvnIWTFurEwE6hFRmFSR7ifkGKOJPjLAgjoTEbap0SoCXnWayoI6C/GGIog0FmneLTD3xEB
aR6y/BcP4SH3BOal3onDm6ga4d4xflKN+WctxTWnfXGvXicUoPyPsRpU0roGDYnulLlEG+ey/brd
rTHZ7qX1vum6FEOMShODdYiW4l4uDb2tRt3iVqDwT3R88iWAO5sj9EoaAQWoDElhW/Cvx8GM7nP5
1lx9cRNcTq9ywFVpuRg2sKaeOc2gNbttt0QgVxAyGU2ucMlAZzT2IecvPeaB9u5XpGjvey/4QA22
aNq7KLckBtgv1aM7mtKaXHi+SKyeHSebHeGjQHDOl8DiPXohUvLZ3nr9KyV9fFlJmJ0QzeIGVruK
hjH6qLQLIbIHlDX+AkXvtepGBwKH6uJXsXgQxjkP0/2L8SIunYVy64cXhaz+/D+UpBnWplszC8ek
rhqKRuVFWxMlBD4HbBHDvyRnV4Yqx9+aeUV0lmYUWDqCYFEwiP3rzXX9A9VqckpV7/7WdWXRRqmD
10cgqBqrnQWKCzixaeDRGt2j187Y/jx8m12Dp/VNRtFsho5Cx+/viCOelIl466fjLCUS05Zd6Boy
O3JkMsM24gbyhqMqTWnPeKFWOyRmhannjN0cxdQMCDl6qUkm6dIiNp6EQkYAWtv9IX08H1ij6fJD
YfUOw2y5Sh+SkI/hYYdfugDeI11vfy7Q1ygGwYP/D2KxjXNTNOWlxJic3ShwY+mSox73L7b92KJJ
Vy7GQovKtAOOe+bLzgXebE8uTy8sIHR19a6ekMCfrPMZdK1XRUu1rNBWGq8hvioBX0ISgLtQ/uy2
kOxGykVb12AdisKppbVG8Yj96Z1Snzifg9T8U1G7Z6ftl2EDnyglDfF6WAd738Xap6CMSlpOWscF
8msmoV9Bg6uWUGDBxaaPV7MszkEydAxalCDLOzcGMhkHl1MpgGEOFDatXg0B9/bMVBlhVBCOkFML
BRzpnkV5MX/BCk7BBvl1///YF0PLTDD6z8hU5BO5znm32/jcjD9T4hJRo854evKSwVj6XUxdQONI
BazVMx9ZZ0i+GnxLm81dllNQwxY17df+nnVjyCEAU3AqNHCyQ2bvFTHkMvdl2R5vd0sTNavE5bU3
bTcr97SPWjHyu+TOSXYevEtT9LmL039S1V3iE2u3ETnBiFZCAK3iisgPu+U74cHKiUkO85qcP4hk
pJr854EqHkm1l+y06SOTnWsRyDLM82PGgIvstj1xUXbcR+nm3S33lLR0Xn0qZCf2Pc7m+/M0ZxPv
b9y7rFi5hUoR7Yh/Vzmg3Rlzky9DSRJrLvSxmAyw2aVPYRJnJcp46iYq4fEjoxFc4QM7w0PiHYpO
R/rk75d1FWdiDcp0FxrVtnTALLMTsM5ArORefCOXSapP/hDi30/GmeMmiVv2VOR4p729oGqTI6Uh
avjf6nZC6QW/Zc72xPBA8zZMZ3/ku/q1MVCUlsrwnLh92CbQPcWgllX/7w7FpWkmVwZnMWPSvJDy
I+Mu58Fy8jiyf8+nRJs/43ZuArwT/JM72eztyFnpVJhMgHthEV8YxvFwMIcPdmzovzUdSnEbCZ8O
1Y2omPOqtqYDJTr3RFNd22rFrXbq4+ORDsVtRFWR6QW3DQ7VokYuObWqFw4cvYUi4KQmPzOAsQEG
IdclQ6iB4Ux+3JhoPOCsQbE3j4O2X8k8MjW5bdlDQaNNPmvGC4diJ9dCjnIsvDkTYzzdepSzzgVQ
SKZH+W07z+HjL1SINOJNtcwdYgRa+l3M1qefFHC9cbnpl4J8CeDMJC2AiJG7Ae/rCtN9J8G4ORHr
H6JOd8hVzQq7RkwJF/9Ybethdhl0u5R1RQ7J8YRCjeqkXLX3zr27f/G1Jw7P5zliDLcDqbyvg84f
q3MvfX8izidVBlRQdvv2GBEZNbW2xkV+NZ3Q5Durks361lSp39fapS8YZtYhYcJcVWYlveFq3NMN
KJWfoGdhv8k9Vp+p/B0py1g5V7RJIs0t0Aip1lAg8roQK8rYYZbrUFXZ6FG6k7c2KPCH6bO4EEVN
F0xs6Nr7hJqX/4yRWKS8pIbRzE5kf0UrQ+OJN+86gUC0oDODtQvR5oH1higglB8bZqK+mjslUwpc
bdyju0DEpP1ZBdXW8B0zRpIBSiMoVHWTdQCtfMpF4l8CuDtWAuVyzYfJe+MW6r1r5VSQUaAqV3g+
Cy/jc7W5w5rMK6hlM6oit340tIEVpz8Bp3QjQao6NTGIJAdCtjgVwTZnnRVxLeO9KdpUa7MCiHKh
kZ0R4O8F/CCRPzYXJZ/QUyzcf5nTzLPUMEZAOCpnELTipdBqwuDmkz/pHbSkkctjFLmJVfzHUlIs
Qsn3b7f4OLmgpb6DZLvGDAWtGZ0LIN1LL1GCMTL/nuZvKi3DwNMNbYQpK9Kx0W/g9EyzoQeboI0E
c4Cf8F1YeG6x/9pGVhG+JrYogVNXoXWBX3a0Kmkh2mX8nwhSuhOQ+CSgFaAW9qHHiLZriYZxd1H0
eCmektH82x/OELY5j/fK2Z/Ab2OrNH/u3OA48iDsT5Js+CBzQG9juK1kA+pT/v9AyoMN3oiIQ3FY
mpEemQlNpKl3J/SgIzMiZ88RS5kC6Svz3Er2fdrHQRnZVWPnBKq+X+gt1GwwsQs5ri1G7f3BU567
GvK3O+01BwBgxf1QDudX7k4WEoRJHx0WWllxswvW1jC/H6JVMQm6W8M1uKkirRC86v758ClMwtfS
LUmPYy0QUDOEpk5oe0k3PjLMpyRBrdmoG0+Z86EAPgB6kZ7+TJeYYW/9+GfWYTu1vPj/e4H1eDub
vnCE5t3UQWSjg5MaxxFHzQWY3xgKb3/GCtKyCUC1UzELEvmrh+25rwDMqTou3Ka//dTRrYNZvXtt
9MmhIPeCHyfYU6k5HUJCOVhkH/ZGEBwVjIiEgca/yCOa+fHj7QC8KRta+BWs5lbX+JG/pZlJvh2v
pAKue5NpL12Pv3UAdEqHXCWaFZeMf5IuKmdSBQUR/Ln1FCuXNlWpfvruZEWWjAEchxTlQR9yU+Yy
cBI2ME5SDuwFachetfgyMheVgawtKZKEjZ+wHuXSkUsOJHWSzmDKqwhBnaIZtuVa9AMSpjPO2vp5
RVpapIAX5d0CcOQjxFV9htMIke86hx0s+pYxgP1y/d1YQ/rZAbmqszcABHrcXBDaXk95GbTxUUFf
pKxT6prFlctdzty9VyFSbN/xfA3CkFFXPogEN/OSQw2d6yRypx3HwW+dDetUdEXmuEHLn6cu12w8
0GivOApHoBa0GVy60DM+svR6uqvtLyNBe8mlNOTArjgWEPjq7LMMZ7IwIHJno+QGDUOY6U5IgI4K
L9IzPUfNbIWoE+PS/OhYaxP7yFaKtve2sV5pDobkKNWglcbkgC7f92SrbSJQscohJkNxEF75jUxi
4C6JAc70RqA7x5zJCVJHVDazyOQGgcr7hIgU06k0RErROwnApmKwC0JDYWPMkymIkImn7fiaqfac
6P0c/X/jhF0760NVfxwMC7+fzU2/5EMH6uqXxn8MptKgdQodW3OrciZ7Ucrk2jSvqkIzOsGlGYxj
kn5VjRzrPsCi4hmj98VYC/hmkN0kW1DAmqbyLiyCCZ/MVCr1X1fJK6k0ix2bZCGyHbhhjXGw+AZR
UXyOHGDaVB5JylWaMAl8eXdJ3X331cWiYfTFUEa2WtoprmeIpgjBGfchbnno1krm0qfzzB59UC4t
SJybJ1q3f+LzaXpBnipQyXCcSMaXnkCVZdZvZ+/RsB6T6OjVrw4ghYtHYdOJBVY7xaFTIAGmDESQ
GeiM09obaWv1HAbn90nSK4rmLvNcOWNj2OShtuv1pFo1X6HSwai0ycKIcHczh/Pz2gUnCUdRKIWf
GxsYL3o3XrdljYlABd/CDteslgxC7voWlmGS5dr/cR5MSSOfoKONKrF0L8KbFe/cBVHx5J3OFGOM
SKCAmmDR6Hg5Va8U4GI9IxKTDKmXdppfrz2Suk97UhJPQ7hfhz7YJAZexTeVqDdf8hF52ohCQiKy
YOiHZl5rF0Pi/K5g1U7JwDfmDSsGrmHOEnmqyWbh3vfQ7pv+M8EinazdCUyI7YfsRyOqjDRyh3Vq
5DzFXmtlElJwkqIUKhwadHhjR/U+ZgiP2bo0+YzEIKkYhGbREQfSWTQ6d7rQSftrBZirjFB/15pG
fKulyddcc8GCwL2cee2d9y6eri1sHp8gV4epWwvYmthXPilBmVsaSxJhlbj4vl/r6CdrDsygt/SW
2lSOirlNQ5RQMdNGASGfNHCGDnujI6szLeZkS70zpV6w7dLESV/InE0Q1izBYkZKqObu6B5VjDb5
kS9vJ52jYu0wf5JvojyyLOBVn2Tt4xf+z4QRimByatwShpui1aE/EJk32DnVBi2w9/DIVk41izTs
Z0ajE1AiOq0/6iva8aC7kftVkPJPIAaWX4G2XVdB10Hv2Ekt68jtiFIbNH1XjpC7G5XvD0/ipmli
fpRv7irw99TILS/L8TlV0OAABeKWDcJ5JrFim28u6WoNRWBd7toVM0zZmmiRvEdKWZPPcxkYly/y
Q0pemEUGQTdHimsYpeOs/qjqhpKTy4s21YkOFKFaVZslGbl66K2jI2G/N1JLvOFdRzWMvvRB85PE
v1rauXgxhSki9kXOFscVsU5/fD/SgN1ZyqZLRcD6/XdBV5mw6gGf0x3fCeELMytleQmTzcag8WA8
oUBOLDfMF7CFF/DQTi4C20O3EhGK/asB0xQC1LrNidvJck+5FlhMeq7bElxWtW4RBiUqJAP8xI2q
vg010VPajUDA3sEzndVXh46mEekDD5YklXuvsPTCpnFGgAmjH6sGx7CXBQCqrZJat/wxodcS3AH6
eCO1n2TR6nqBzNxemiAzDbu+3lUf/rJ3xRQx9Cq3y1UJugyui8h2CGKwKhuVqtdBcCKM6xLYSTgG
6pBovYIi6I0F365Iu1zc4X3xpqE5zFQ5lB4hLMvuiVbEjTQA/2Xxexh7lqXnyDJ6dkjX+DGI27/f
bLvth+MHhNvCb71k0gvKwKDIRx6Cxb4ZMNbC5nh47il5TCGQDuNMGm1QFu8oYc1bWGH3FkSVmbAr
1q4+6Wx7h38fGJKzrAZJ7n26AOMYjbNUiD3/ZLXuA+LVD/w+DMroQxrsGjpOv6Qkqz6Zd7ih7lix
8iWwJ+G3OTH8jsGwL8ghGQyKWvDH5bQuSksoEYFH8nobbCKUB2/vFyyNEM5ZQzgui2JE6V5E5RcB
FDEGUgFqDk4UuqpTGpSn9YsMqRc96ec1IW2nxx2kydc6xrIFmvE9w6ndiQ5Y2yWLsrMTA9pZOzon
BPdSvF/nCnic6DF3J0SJr+Xya9MiwkNQSTNx6WFnSyt4EnslxEDpaDKFsX5xC6u3xE32c0liLkrk
DS4UZ6W0odXIjGRnIGHheWW0K+VANgtnNVEX+iWjm3rcP1tQqdkLbfAZWce/bdEh6i9Vn0Af4RkJ
BKwSDWXLmOJvLtomS8Xn/vGGxpcR72nECjCkJuJchesTHZhDm9rpLyVrxuOIRpP8QN1fg5Wl5z9I
aLWz5wYmlQKRjNHiHnEr5FBIKHw9JOGTlLjU5DnFaCBSo26R9xL0z8wZ+efyrC2wK0dYrxjcgKRF
Y3SK5MBrBLvKrLFS4UXLRLn19XvBzIQ+TXQsqh7IwR7reJGth7lluIHVEegOuzzFOt4GbkPbQIhd
jQjPEIGyMOO2JCOPIW+BF5AQY9k8nl+K+F2Tba4DDgMadWZP3pdz8J8eQcdt9qaSLSR2U3hYP65a
R0rv/B6Ol8HvWtpgmVdDEKRo1TcI19Q7W/0kJIPwkePREtapNYejxKfsVbWhTHeM425nr2W0XbY0
ESiXX2t/35FBxLXmmLCYUzsQQtwo1dL2O/uO6rWT1FxBUU1xxDiCHAoc2GiEe+xdsmGhnTCtCETb
Wmv0MhPjo4GqqSZkRm42BYYQrMn9X7FHb2qK9sPh7iQU75NQU4nKDJ0ZUjVTMG63v5611jE2XsLZ
TgMyPWgY0uyC5aRMmDRpn4YLp4kZBnnukgZVitYi7x+uxtulKQVpiuUAJXHLFPPpe4eMLe9ROJww
hYMjCKcb4XQvpcPsE35rqg4YiTY6B2OYMonDFTT7nhkxgLFd+nYyxP7FRElxiPKOpg2u8MTpoTOd
xsOtb2jLDAGwFSGM916lR/GHo4lK7uPatfYoAVCEqMfaKQwltAxV8QFtE2fowrNO0PELtxMEepfg
8MAOT3H1lMyrhtsZOZg8wfqxahzX5blOH/lVtzVqJ3JBE51vXGItd8alWkJJypMfuyyHQsoFyrM4
JX1oZzefLkvYoxNNm76CIhChg/kWzk/Rd+Cw9XDzOjhhHj+qYxCVvuurmVGr8En70YZwHhwYpUzt
jzpPQlWQVzcns0cfIQI8W/CqV+F3uqOVvNcEsLGLbyWUsCtbDYKGEKatoSbDWcO9hBX1wUXyoYVM
mpoMi3O61xbnwd/xdkM+FT4qt36v5oRkmrGzK4LQpBJy+aQuFZPd+mynMitWs9g67qof821qnTN8
uig6ipsL3ki7v+bzSum+H02zWuvKhKgMf/YEGijHuGLU7hM94JeON1Fi99tvrjQvkT8PydFXnni1
JSjy6NGEGSrn+GyW2IdH/jyLnXezWVE+6DUJ1nwJpEGjdft3FtySNL6XbRn+R67uGDbxEre7erbC
gVaNHyCHRz451sCTvLz/SmaCgDzXVKAqIUW9Amk+gJkXUjl8YoK6ORIMqLsIgULOqO7iWf2gcRuS
iEGVKIxlv5HUPUuhOGh6XxC1G77liojqldyHSR7FzNsTieXhqbU1IPub+OZP3R3Na/ytNLF5fHVd
pVnne97U/Z7S4ATeILNuwH5/ZeTe1KPQnCqTAvBqciOBBOFVaErCd3sKDoE7h9iMrOAfLUQlG0n8
jpI2EfSD94MVW+Pgf3CWUpyotNNAlDWt8c8Pj/80L+jZhCflDDi//Om6hsOgnjamMFS+Dbj74MxU
b3PVxUPgFYPE7afAyfMnY30fYW1aRnZysL270ZiGDEHnExmSN0/sR1Yw2wQiWzhwRF76loS1Z9jU
C2STmYsPDaNnKGc9g3JU1yIP6vvzaFdjoMIfZsaAkEzFTiAGo6t+9P6D6MruiPFWz1LY/szfOBdW
66Kyo/omtfhuAj12xzJkCA0ENP0IfTvQlIRPXBS245xyURAtLr8HdEo2Ktytvh6ZXPcEhSgTgj9W
Qz7zDRd5n6+BFIAMHEwe8UZ0jSa8ttNOJlYRM6EJalXlOA9E4aDJV1rt6DLEFQ64opiasbdasGPy
q867UE3cixPtHKuwQH1qI3jEdSPngHv9OSoICTr8FCuNkuMai/By8m7wWmR8IUGrMkcbnmyU4yvt
lxYKNrgGOgOZyap3WuJyJHFUGJ1jEyKHcyIDZDG+goGMKf8GbvsYjVrw6tjg7YwS97VQQiszcxLH
2u1N2oJo0deQ6gSkuKO5z5hGlvqhveZfDycxmYRsv0RJR9A2Ruk0lPZzTjacpEH7YoTebVo9i0Kk
PNVA5L+pErzGEKzelMCk5QECYukRdBj6C44GpIboJdXbp3JkNTZSLUGqP6rdxtOAgiQFRgY4bxBQ
KPwFc2T0/d62JkEPd6pRiuznrSaExaUUHy47fSL8yYqKcmMqQCCXlM5p/XDmDsXZsgrQQDRa0iS+
daqG3uDCXKYfnfVFhzVieO+zLH9GSDh1zAI+GZP98kAOxwbXtcm6xNogrWcV9wj+r0fnACOndK4z
TYWJOLfl9SZAuBMcSTMqKbs7+gpP4oNIpOTCRZRWyi4MzQL1hQKekUerm/1OLRl9hDiLwCyvWo4O
ay2LVxRZPT+LeJ9xcUqD8jEpbUZqrQtcLxyjJEoSnCyWc60v4dnCtehzfqyv5DKpNEBbzEfwoNBI
BQ0m3VM1R/XZRbA64bJk2CHjx22Y3ep3bkszFhzaNReiMv/buiOYp53YTHuI3R9V/wgBV/qyz6f9
g3FTMoVurfGyL+s2p8LTCE/kBKmQHIB6pVJKrOdWHWrUpw/Oiv+hBkxgDzZ1dSED2LuSUaZFqhZB
NucU0Op6WpIBGDFH9pnA90wtKKds7X0j2hNpO84kTXtyrR9B5vO5CXLmMqJBQLIAqfn7vkjzEEfB
CTwinKiEHWPFrVxQF0p2aMWDTwJvgAvrbWzCBT0bU35CKN+C4xiMRSYqNZzqovHz8DjjIMzansQ+
3FJMYmDeLcxuy8QYVyLd42KAukukIxMxtn0dqUeCxS0b8VyiROLfzOCSECr6SRFGOV3VHC40rTlP
kfH5cir3XVJJ19nsUx4U1TIkRF16zt9HNUwwzUj2gg8uJxFPZpl8xa8OcFHmcMt9hjpzle11N8Iv
ubCispC4Q97M3/v3ZLQg3Mu536zA5VUg5I9H+z4HfHfBBPVGNWrmDab2qwUvsnDob+KlK5vAa09O
TuWxexqn1CPH2FIH/E68QgTKagiDGGKxmyQ5VfMWx2Opd/pHgq7ZL6YOp1aCt/ajqqvYvWcnW/1Q
6VRNlNdSSkn/lhsjkrnQ4FCEifLDCr6EDEQaA1zKGOqZGX9VdUFr/jC3TBqAH321mbEhCpulToNx
412bFSMSI9Ww12SxSGO2k6c1ZdMqiT/PS6YwRoQtkc2erZO7CbLY6vjso1bD3O3sEtdn04I9YoJ6
DS6CmCWPq+Z02T6DQduMYAIMwyNtPD5mloSeLsFCcJmTSmjljtmo0BxHhdHlAu9rLWQe2qegR9mH
Ik2f1ZNBwXv6Ys/eDiXe5OCqHK8pt+lWlO74/gqjotQzNS8s8982V24P4al3OsslOShyDT+yFSJE
c2wdE4dp7qJ3YX8q1lOyqhP4P9Nk2AEuHROoNf4UhjToGMxiDqLwjMQvHtEmBy2K0BnDk6xR9zlD
IZ0f9wNvPovXKibQypwWQrtJuGS6/WjggCa8fYFkh2uKilSpDitV7rEFdBvk8bfM0dOWSFWG28I9
mD6eeG5eNohfwFW/dkQCdoWwbCZVVed7u3e2M+ZEIkbLpT2LWw+ZtDKcSuBOXpE9In6H/Wn+KimI
MYDbGRweiCmBN5bLrLF7FtKFOcFvrf4Q/w0coRP8nWNqBD8dhPXszd28u4ukQfz5gt6QjBBCglFY
9fb2woPaeAGvJZIfM8+nU74wrVJlh+HOebnLmd7+3HDSVHBweE35SK/xlG7lx6FmcmUI7g42r+fJ
pICZ2iLZXWRD82D1JTMU9pUf9rgegbF+43VP8/Lh4hvnNlXkAMcIneuDNNrcueRxQJsg1dU6YzLc
y1+8WOrZZtCKlyiPB6qxX/sYc/FLNj1aePom4zz1S+j91GV4ozW4+xZ0W1r7k21WNUj8zuDcLcfr
+k37QZI2KbnCn3A/NJilMVIr7uW1JN+IrbCofC5dRmNUL+I2XJHs5zUk8DCYOcjfxRuhzn+Jaar9
Uf1y9plq4gWJWS+ZYmPgweKl7h3JAF73gXyv4tLxDGI/QGAyczEIY4XvZJqmfpXVOnUxsSMNh6b+
j8G2U13cqu1u8mIEqH2YmYIpIQz/z0PLiwQAaHZaGVyuLKW6Nh5h4wpqnO80uNJp8pGhjpCf9mmJ
ln30K6o7ePJSlwUhCcijkdUoBPIs8+zxJSYQq4e2l0SuY27fiQ7EngeT2BbFlsAuaWbKm7o7GiKA
i1A/kRexbiLLPPqhjsyYQ3lMeK5qW+7f6WucmddfEBN/3P/dHmLmvy8OvF+cuWkSJgwzmmXr84bR
lz3ncpIDYFA6jzECUZALhLypxaGBnynSu3gzEEBeiHgh/qumVLyxhHacMPg4GPwf8OsTUBhC/ptZ
OrmBxhTB9jAB5WvrLUobhsmiv5sbUe09GOVpYWBnGn1N0xaU46wEZWVEh4BbSE3ojcaksusPKv/0
PlC6zpI4uUaLrsI/eNlvMH8aSAPqBMpLkuXOeUr/5Rk43xnuu0nRZQzMPiUt0CTeRhygsYmTmXza
xis8ONxGSDF3OI6d78YDKB5Mpfar1kfaOgTRKusbJEk18TthjosCJjXBR8KjddzEqjHcmmVIUtkv
xiT3qAMtd1kjEZ/wDuZlw2ePUP853PI/98oTAIf5rCanqeCFRb2ruVuVT1MFggCiGlpSN5NtDKhN
p8AQAyovfq9p1H3bndLLAu+ueQNgqpBUIutSDHwVYeaZ7UlLlhzBOTIpMEs4B9xc1RCLn1CN8xtO
XASyyXzmk6+vhlovMmQzYLwAoCH+ZFv3kYn/aEMjYB7H1wJh8iAeknvaBvjIlYYFjKqGo5ovip88
jT6Zhw/4lBPOLug1RzA5qgKJI40/Is3sUWvmizcw4JAlCIy0tX4jpX/j5LMo7MJ67RwVEk6EoCpD
lnX29rBpkTihDwmOUWmLUcLJmqFsTlnQ7qkq/zaFutxv0zX1VqowjSwfGnHdH/eqvjzZ8l7QAWSj
+rdlXMsa20vzyQAdwR5J7UL6IwHVrCO2igwj1gneyYc1KDZvhXejA+LwTqsWL/XWrSnizmGB+hod
/VEFPTTmqKBz3TM2CQeEN0iiJSsQ6yFemusqSsg2KHydEAWT65mEkqX/53ncj3QdWGbcRiShmFf/
Walk2udEEOrMOn0TmL/EHKIWq4hbQmhfOkdalTwz05WbvxzaK8Roap536SeP0hT+9NH1pRpEa6Jk
kylSZt+WrTiFtxkWwdQVXoy1LUgaCn/HYpt1glrE2DM04GGPt6sy53KUr0ABf08Naio4e5h0Cv2o
AV5zLMjgw3J3oHcY3WWNrb1Yxx1Afe4NnEKT9LCprHBfsco6qX+vybU+RWfQnYQuwJCk1m2Swm1W
WHxvtTsB6J0TElZy3kF3oJ4xXnBmy4B6M2uLgwV8PSa2PtxgIrN97/uUF71n0PAUrNAfXPt9yoey
EXYUzzUNyEWkL+COpT/BygVcz6rt6ZNED1cBT9gJJMG6DXWtvao0imi98mQGwltklIVhbmDbKKn9
kDG9WTEqkVanIRrBTObis12TRUi8eMEY8nW3OtKjIJF+XqDorqmK9akKzIUmxD83RfpkybuwXPLL
LziE9DmY6STnWuoivHlGtv44/nDCD2r9PetMZhJTq0Jvc6ApIIhz5Hwg9DHwWRuxYNczo2n0hVzw
XM+9sIUY+RFJ4Iwfg74KRTqK4J3fW1CsUpj4FDUml5wTTqwnzql4olX4pc0DKuvTbov6uQoxfOl0
lX0HS9liuuEMPdDeA5/rIrqmmU++Yb+vJX5nAXK6eERvNBbba2ggCAfuB+n5K09Ih/S2Bv6ASLLs
RXJlL+cJjh3hTNe4bimk6m3M8YwF3iq1PWTQGOjgxOwb2iCSZveZ1lS9xVZZfCO6/UotvCDoFw8J
l2RLl5E7BptX9f8w66y999B+DA/QaP9ZY8L1Q1umjALWM+/F0K/uvBcu++AE1M12g3hxoFa+szgw
T4Cq4tdQwdyVB/fvyaGZt0bIxq/X7eIGELJjFdw5bkP2P82ItN5FgdRoTwT3hevLywln2Z2st2DA
TTt0XOT3mZI9BzIsz6hEUi9YSbVe37mvdlQXKVgux9fNo0VJBbr153hN1JMCpOkhVURSF2KdrBOt
3mrf/ljfVGFh4c9hX3WlJxOVITfmtAHXlhEetH9ZpfdbNRhbNItlo/Z7yPfFyVj6rPSnyvSAkAJ8
2Q8jxg4MJG6B/M4lrlFLi2ohMD9P9xw/Uu9INq3nzImf4CmL/AxUnWcTyrFfb3XfbLOikxxzOPCs
kPpaxoGox0UkL++PIlSf5rmMMPRMKQw6xeM/Qkf4dBl6RJbJlwO5DMQQahZIq3hbAxum1W3TU0jO
bUaetEJoBea54PEw+ivT7pxPyWPO6DiafN90L5+eHCXLIlYrlMnqRthIs9ojatYgLx/Cjood9uj5
NiDvZdLgvS3qg4/Qa6D62/e/oQuB4F7UvACMKJFj18TxwNTPsOWd0U8AuqCW5QhzXy4Bxohjqz/f
VzqDIjds2AvnvtQyKvowJ3SEN/CpxgTtuHJNXdpzXDMMCS+oCCAHtHGR13fyDN35gb7dYuj9uB2Z
mdWolu/avlzm12Z5JPdC+qsumNKWOUw1d3vT3a4rB+URXhKdcd5vbZ5lvRPIAjZOf2w04Czw82nQ
Zgy/h3dhguYl/FHZE6K37wrqwbb+RqiWvnR5D7JbfKwTnW3SyD1oxRHfNM5iMnhaXSGAfBD97wmA
78tn6hFT42SJQy4tWv5kFlLtEvup6vQgEco1lb7SSFTSL1y5CLkJ2dJXdg7RjVvGekfhRIIb2Cpc
Rbn4lUOTa+3/rjEzTd94/idOFFafE8j/95jZAljeB2ARK/N6vq8/Z1DoNvp8MpGsYDqHA8Yxu/+B
dEOTe88iT73f5riBrqVUWU84cvJQJ7K09jNCqc9cPpac+GCuVAjMD1NMDznqNhBDWqHHa6atJuGj
q3et6nB0DlDjwZP4FJOR3ljsEisUrN9sTeVNkwt9oO7sP/1CLPaHfYeDzmFYAgPwnr8TfAzfukzZ
lOEZU2HMugE7YlELcxhNq1OviBgwzxCr4c9dwxmWCeinndSzNjgjpB4ZrOwIT+S3I/e9GNBS7ETu
q+LbkjzN9z2R7gQc/gmoNJfcdhKYcxXBloRZo6Kss8gIK/09yH6yALbp54kyojmdo5PVT0lyC4Yy
ZUfV/U2qAYWuRl/Cy+6P3X4n81Q/QOhN6GyH0Z2EAbOQFN6RFKLK+Unx1xj56iChuDCIlD9gU5rB
DqveRWBzVBV4h49yO40FrOHLY7bJ1Y4JpB95uaH4abfhSgGoD8/ujlC5mIESug+E3QmveB/MODLO
vPKmH2UqP3yLK8eWqLYsOYKxlb8tOhfi8H74QjkAe01z269dfcIVvvy4BH/5Z3/UTFgurN1FkgGT
25NsXMcCXmMNW9U2p8nBNziI/HD81ZbYL/v1j+N9a0shbEo6g7sN/A9QMPHPQDBFcxiaMF2VaxSv
v6QuDyZ9jzZKNl/fWmbglzsNEwdqP7I5RaSmhWksj7cAjHmx9voB9NgUnuChZcqnPEvegsaRNTyz
LrjS/1ln1Liz+vzQ1dEh9yomK+xgQuD9OODdvUs8xEXK+1e4dcrcJHZAyuxi7egUcUlWixlOfl2v
NIZdt5ilNoWOIBHyqiUjvXqXx6LEji24ixMfW2w9SwXEANldfgSB/Bd6Bvhi3VUth4n0oOVm8y8r
3tgiOzpO4Mv3YByO9YN+tpT6xNZMHefKS5C8tb6Ty3F0SHHLHL4wlIMWdYWpQM5599P1IrJz7Pv1
dNYEdWxT9puO+S6ahbMmkY713u1JR8NH2rXlWoWx11nAZGkr/Yv23Ujpt1u2EoFxvUGS0jypErry
7WtddVpMni2lVmH7gJbSF/VqEa57sLnLp3I/hn+DgMKmJ2Mrj+JVYuMmPovriw7Lrgnat5q/Zurh
qdyigsi7pMZOH0nbMJUFsDqK7LKa5nGyv34XDwsGWCDOTvhfQm0f15v9TIRN7+uIgO6DUIhoD0if
RD+GpeXtU24UlHHg9R9JNIei7VEM70Nv35/222UkET+alOXqmohFeYi3vD8oK3AzmQS+NP3dsqfx
c6ycEpsy+L80Y3AXt+BH19x+JgIW6A6jVkw5oMn+59I6qwFAp43deJ32Nxsl7CBIowGGKQeAGfjU
qzY4pCCYN99yTRshAuzSm4VYzd//JMA58IfD98Pzf1K6oycGbOg1xlhEphIXM6QMx+JvwLt6tO3p
kCy22hkpbj8bT1kLt7sr+fVINStoRVzphAZW1IzNCIYisPr4PS3K9MR9iEH5VDlMYte5XXUxWh0D
YvAfd9XLFsEl98zwr5wWacNrCJen2R1+14nEU+M/xOd0w/b/5O050VeYcAhousfbKm9Q0VulIM/N
AGavxuywAL1OkFg15idrSGsEk0sMaGuXqn5Wmv8Tv5khS+zd8zCHCHqPcmTVPtumMFKL45bzTPjJ
a+zDTV2DrQt/Q82WtRqo+cSZDW4InscdN36ELpCsoDkWNBcyzqXGhTLDVSSOZv2hyIGFqGUdADdL
KZSlCx8ZMfKDcPLrZDklZjfU/w7PwwzedtsAV1t5FBEn6I30xrI/b1aInLBL0ZbeAB+6JzRbqElX
N3Ao89XrVFf7u+4VNSn3T+nB5pHgXi15e1CdKsK5MfocXFIruHxXqecYUtVLRjysNdIxsUEssEsP
C3W1jKVBkS8DbMekKNRoWUBiL7oucnXr0SQyd4OSMc8ZjUsZzIjAkYbmXHc1J2cAmaWmzfW+i+8q
BgPPnb/6+p9gcRlGq+fS9N/flDPcUXcWi3QCXTppDEB2jsztD8QkXIF6U19Mp31wnHy5ZC08Gpeb
OFntfl8gqTeXLLehtqMkX6MAAf3tQ0Cfi+/hl8eHCBzJVvnp6Y/pf25ln3qGrXeOiilGgRDVbNN6
K6nKrEfLSzSUWce0QZ55QMw5Z3fdssEhQjo4xRTboKLntywwG4CdVlgbqkzBUtrzLesH6IAXT/F0
i5v510fDlzRNfk9lzMqEvfT94wDtXVeKqJqJ561/sP5dBs/evDZ84KKpUJbWqGy2hjFLT6mqENAl
qM9an7hmlMauFyZEq4qAlUsiSZYdyeaXZ8o+McBSZiYRRxNGFZyUY4DWb3O7WDLMH1C+qcISPJK9
LrxZAKlS+1ZT3sOPld20iFcRdb4mKwidM0kCviIpn/AA7ML06HQzKN8oD5xYZYJzSBKP/KxsQame
wsXhhgpo3jPzES5ej7YGv8XMANl2ZQLMIoPYIlTiILu+K+/AO7BqlaDHKz7i4j3onKNTFJAf5hB6
l9hb1S5J/4Rg5CRi6y2GtyhSjJ0E2jAp7AUz8VNRvKFZwgHWoPZjitL+LWV06ruCsbQV+XK49eL8
kA+HYDaHdkFah+SDcRJ5IZuRXSXUIMSYYGc0XCc8kiL0O4UTsiF1bQ7/Cijc+92Cte6Bbb8jY4H5
nlbkjRFanAsyDtp7bPB+qqKkaBbbg0huAgI1SneA15RQE01nukYFyWnUykt7hw84B7UnhozQovCd
HldoFPryJKO8DhasNfL9Nae5Hxb8CP63sTp2O/B56K1moQBIU19U7YGnuHO/OyYNyucXOqsnbzuq
6D+X54QPtqVdvKi+XMoWOrUrfHukEBsUZavwG/Tv5GE632NtZ1ZC8RuUMSaFjab34LsgzMA587zT
UlvlrYNTTlacNKsINQskad/PJRLIdfewPa14GkvIkrvz6/rBYw7vGd2YQl006yUVGp2u0g7Kjqo8
gfRpRhKaUKIkSP/OSvAHUkcvnDcXf2JQeDw0WA4hFnrUf7BOkT87GzYZD18XcOB4QpEoazkU7bp1
ix4KNLhM91pjHsv5KTn3vXw7bprkv4hhiayVSw8KgwPEmXa9P6xzZbvn8QYuuAWDZpoUkO22JeJw
FxECX//wipT2J8WxCnAZeZDPEpL2p+bE4w0W55P8RweYS7rUpAAgok1I49k1g9uk+2/5Z1OQ5DQ2
PNQQhgF5+eIFN8GBDNuvrKwZrXkm6MQsAkuhYooO6fB7WCLqU5todShBgGacMnhyLCJFOPhuq4nS
xPbtIqMnGNHOgqwr35NVaTL6exXDlYP9c290gZCmFS9GUm9aDpVo/a6LVuC9DouEAA4xIwMd4Den
yo4oUWoKP4kMq6XxfWtcf3L5dTlHoinWczSFAEQWAE+z3nbpP8nHdqgmAw1BSQNgvqCQcwoP0by9
as4OGzDhJK48BiAlEEkNF42lS6M8mxSnoorgLMLyAQHOMZgSkKYI8bVlQYNbwYyxPx1eVxry9+YY
tNLSS0N1YQoNLs8w+FPWFJdrTQ9jweLEljzTb5lYF5sIaxW+62SGg8rPXWkzR9RU45JPACDZ7LsX
rPgr7I4Yk4BosnHzaDBe5y36xsRhlCyderEqg9MBDnhmBMjuE1AtcKUe3zQ/qPT8GE5M7exeDUP9
qQ8lS+eQSoYrIssOUuRVRz/dX0rgcpFO4aumZ3Gq4m7jNzdMcJSm3edXmj6mKg3//Y7/lHpVDqWg
bu8udM7NzxCNvYIVSs3QChrC38Y9XIDUq3f6ArxHXj8M0ZZG9aJSsvzwMa7Vj8k10uZwFkBN9GIp
qGnIqvtdWhVDW88YVBRe8/WAtkGwne+mZS6QNbFfpLW1ikdDVUQ6XlkTKdfAUIBDxnT5Y8yYK8kz
nOw8+sbj/Do39f/Zi75z/0/jKqDE2kcCR7M3B6vHDV2bipFE5C2dKWidvveOr3ItoJ+rtsClQuqp
THk2D59JA8VTrAtmEPDuFErPN8Tc1ps2T0zCTuP8UdBr+JqpOwKOLQ33slGZXCwjobCrD+XTIZJe
iTOLBtFEkJGg0twgFe/wSeYKDZ203JS32dT6Kd/LBFZqxGY9j5PMV4aCZi/sZEhQUlajvP4UM7bm
ANELKOThjoMNAqLwouBimHacj4pdkJAuKjnIZfXJEuoS5HSGBFkdjBS9+gk9tkA0kW/+Qd21noEs
0jqvfEOhnfWLqboHISlu+S0jA5MbmpzQaBr8zsDigDWip2BavtH8aiKgFmpxaBQRWPRGYOllxmnX
+E7aGxj2juxxqSYf3CRysnB4+3zyi/Hazb6V0Sq037rgwHeyq0tawFBOgqMO1UibmnStSBeImLrR
VOnNFF2GkuaW8kBsKZaIC1ePN0T+V9RCfzATZaYoJ8Vx3ARv7ql2fZdpVFOGn9yHOw89Ykq3eLQv
XQ7ruOUZi6ddXBzT0MerEGwDpTsXIjpJI6MGXm+tKa8ehH0+IP47ZF25IZQokNjM+siDEn29SNDp
fgKdvbSIT8mt0L97fmYsmmzS1S+C8qhWU2HLT2w+y1w8wBkCOo2htCGbGnBIFbFOb32AtIor4Ick
jGTktrBbsmO58yYluaKeAVEmx6osEz61MTHZgl2VZFTCpXkW3WhiXzZgQsOMEu8pB/YniwIQgDoL
XbAh6a7gySQgquoBQdj7VgeV7W4OsDjDmHja18haYmyfEnfoe3ypBSqdCRBC/13ameY02I2MdhvB
K4eZJj2dGcF/TV23kHtVsB0svYWniqGbOsPxvbAMdKPIYE25jpNLILUP6GBW7+NMZNMQb45Fb8rv
o6x+5sdRAwI5v3oZ6pOTMgOqDLH2YcSX+VDRF4L1dwWFBos/1kHsFXjY52xS5bsS3ni7WP23JCK2
V0c8TT2m8T/LOJ/67hmBr24uARY5l/vuZ55gKMNWlwlzx56sU+50q3eED823OTI73uRoNURTkkbf
3pk7NAtV0sjC9aRDTEJQsSuTQjiztnKMW1MoQu+40qsr/a8tWMC3sMG+xYg+dwwSRV1Ws6rzcrDc
nFCDJk2fjXox29KtcIdNA1Sa4g+hbAx+LrpV01mgV+sdvtdnD80uHREIJtIVjx8D24iER7kKzk1f
j8DPCZnGRs1a1Qm7GQCqTrJUH8Q+f1vqrqmJiU2ecyPB2NY7+ssrQ2i6EiYwFuK9A3hoWVePH3mn
IfMSQjJOpvgoFz6DT/LF8eH/FAGtP2CA5kh6OUa6bw5v3i5NVrmRYqRD5LJirytJWyZ1EZ3o6rAP
wJuvomRc4QwV1tgDfGnOoFN+QnRHbWSIjGxmOIO+Js+Imnd65CfiCjm9xrWaUmw+ZoWfrn3ocZx9
mgT2AU39FHJMu2FZEZrHS0DsygBdRKMvo9Rw6/z3/MmbYnpHv+p9/cO71orbgK2ps7PHEHrcndn0
BOo4yvEG9NwTMvzJ/Pv4LHHiQyfe9ApOvfzGTE4ZGjhUdH+nQgbIm/rXiFUwLUHppff7XS3GNbcV
HEbDrZQPHjITD3M3HayUc2PMf0vmp7wPn9HNDMcy/1kvHctMA3mPbDHGQidvAesqT2pcKblbffcq
icW1gTbPtz5bJtaP
`protect end_protected
