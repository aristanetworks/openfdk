--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
mx8VKiKc7M1Q8irOZqDIoT4IJ9QKrekvV4E0TUo+kxw2WwkE/FSK1Zgkt6MYngLqaeAJi+iIM1V/
AiY1pCY+ccKnHqnQO+N43CmCWRu91R2iGHhTrgwy7nT4CBj7J5I/a+LPFu8PU6a9/W3jSKdl1IIi
TiZUif9Cn0UdPfOHZDByNDQzm+JhC+Z/S28lGwNFK0lHIkfF0Fns4FTVZ31L1AdGRnTTSnGg2esa
lC9YiUDOCbRkjc53IoVIR46Tpu2fimvp+0ZkVNOEX4QJppP3fxZ1z3ytPNBz8d2qFXXn+KEmWbpe
UU3/Ru8Znbw7KdoA41EQAn3MFojdtZ+XYdfSUQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="GhJTYnuVe6tHjjBws3AxtXG7OKAcNZSEH0/tZ646JNw="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
niy3ZE6FgStyWkhViDEvCTI+UeBxT+Ztm6clKQw82KOiRA80BsKpyQLFOwRF3qwkLgqipAFKk+wk
xQuqYkMOgq0HVgDpqxIAWWvhBbNa45Vhv850a7te5qD8JxvdtmJkyEV81ojTHaFAaXY1mg/FAqJt
vTKVi9DDk7E/J1rhFkzbs9dzbrtSV0/Lu/gFrvWQFGAYUk0Lnr8h83DzfURfkp/zoyNQ2AQ5ThON
c00UX+hdVYHhdjU1r9/0Mr1GSR1dFaP8JG1l1G/wEujeOpPoTufRQy2euq+e5/TTCh5KQ65uN8B1
rM0baWLK1eZb3e4Bp85CJxMoNMjh7Kbs0Ktmng==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="Xcdw7ComiR+0kR9G195Dmc/NbTAolMWbOcXhHrIujkQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4672)
`protect data_block
X1XJR1IWLnbTooytFxYMN2DPX3A95q76oUCpcXvyNJtRWXlSCL4Voi2BVrrfOGFkvPfpYBQ66EsW
Pn6iY/6A16ElaXqLsiC1Oyw6p94iND2AhiMD/xkMLC2+z6M+eofrsyWv17C6+cniLq9oG5BNVh9Y
RBNr+PSLHSLSGLAFdPrNKQwBdeEUiPzrKe194oq9gT8GHPFtIUwUb2SzXLx6yz/1ss9gLo2uCSTt
vBGluQtGk8TG+IjnS11GSnysF9KTBHdlV64/qV1KoDLNOLwl3w8vt36/2m+Gc3hpbJmEga5zwLIH
9NO3R39vYZJ3RjQpymnj6JeR8tUufK52iajTcTtnUiw51r2E8wjOneHsac0N2poi3vVW/QXsM1sg
u03XXhJ3zNuwPExYmtvc5WCkcs1ih1P4CJWUV5rj1RDyZT3aBrjZ5wHNWhXkd2dR6yE3zP6Ixh3T
LJRvZUkUn5q4n1kDXx/GadAMtqJ2wnfapfwxxiKFT37cWgO6gA+vScro7AkKcZfOu6fYnvpSXD9B
ggq8NKC+Kek1v4RDoYUQEawudWwjibQ29gr275oJ1ekQ9mWGbmldrUVmWfj+vw0coy94/msWwaWh
rGbhBTRCoQoiznp/EDesh5enQVt2B+69coMqn9WtB4rSF83PulTcmHcK5nana1bLt7T9hVcWQ6MK
2r/IimP2xKebxnM7QlAWPYoC0W2fEvZvzAb5lGpnMSFAkQ18a6ARvIo9LKtxan5fPKPBZk+IVZ1x
74qCECr2C+nQalqonEw5yN+OJNRjR3r9OsYFS1ZK7okixdBDIjzHCW70ZWYGln2l+drYmw8pw0Wb
w7duyxC9dtJCULqKIRFxrmfEob/5tN/CYeFV1/cjSY1HXAzNWCPQQkZcWraqJOr/6fifdrQDav7n
M8JG33q1PFB29cxGkW9dIN3xwDH25n55Q6V5l0vtIMoV6slv4UZ11OFFuf1ga0Aj0tIbPgHzwmrB
IqKndDPcmTXYVgtPuHjotYwC5rdRlbMRkMRC/0yTjFCSQE3KVHYtLSlWSz60q0Srd+YsY2nNBpVV
Bra6MPAMlWhZY+O0Fqu+ENGdl6QubqAFufcpWrKLSOkwdPoQv2QrdE8APJzGs4+hWLtiEYkbbRBm
pJV/TLoVSLD1miOOcu6NCHoRzRspnIq6jWfIRuFNgjRgvNB0tjJP6ChQ5NnuaUoOdSRcRLoHYQf3
av6uFw14ZbwTe6riCiNB4s6QUjgkNRSY4yyDdkyFuEGdLId5XTYn2pE9tiOXsQvM1CLgrHp68Kx7
tJNiPy7jF3zZDB+nhOJM7CZUQg02VW+MEtYz2HVTCB8EgmIaMw6waokzwHXWNDPnYhRY8xUz2e0t
wc2ot702gwDvtlQjeAw2D7As3lCqxFoLjEpj8Qmj41xKsd1Nspn4cXI9Bk++SPYa5Ot50aqQuYET
xqhagOr17A+BC2ihrr2vPV+ZOtiRsEsRbnMpZ+3w88U/7DKx88FRWBBxPipjIzaimyBilSGf/u3i
XXjn2dC6FsmsyqWkXdvs8/gBTEJpFGMrOJFnjZRWvveom59cqqTjzz7yJhxyHiH0T0mgAY1ABLim
4Pm5aE4IX9YBly4qs85VRTbhZr3jAiXM/MOouVqhQnEJVidX3A/zElQlCK7oqnivzuQ3t3b9PLOb
ZPzs1uh3AUq3D19w7YiSbFmCDc7TGBmEnHNhG8cdwQwCz6VyZMEJHdYEQ5/sNawRpTD2LLZqF5hw
iGgyqFqaIyYpZWWoilpQ1jKeC6XuSz5Sfu6UynG+A7/wsoyAK3+nciesSigbmuqVE/2ks0+XnANm
kuL3+TSeRAluaTxe4uHNlnJ0O73QWUdZDOKaCUUM4xuGQyu1nHAuyKPyqf3s2LDRfWk9HEcUchMe
TvDLeAuKpysV3+YMw7MVb+aWyVU7LVKS2mO45pvPoKmQE3FVMUIDSEoHWnkAN+eoi7u7BKg7K3Q6
6WyUqVthPRzqw1h8InufzoDDTvRPZMkbbvBVCnjwvgR8hm+umv+gfLBHkS7sXiYsOOnenIpD0Qo0
oH2pY9638ZD+d7sydWpJnh68td1ElnIYvGD5j207HglL6uqGAI7B6400C3RcWvrMkvaL0/IWwQex
ScThlAoX+H5Y9Neg5n8JIHaSrLViCE28ZgotGU+EIDekGbihXbUPvM5WL/04optjUFgS+Am2rCuL
bXLKAsQcpQlmeLvtJ7w2Pm2Bqj+M4+QwfqFdzpoDP51tzZqWlrHMQD2Qv+7Du3FeNMOPiIpvj9pa
lmgM1NJYvhk0Ac8/UVfncSIryTo+KO/mh0jpyqvQKsUuvusAOGouom0KV+VPVXT3Bxtb6jTU+PZJ
I4e13IPogWIEToWwPbjuCN9XJYQck0BHmvb14KTdBq96H8BQQGmsCN314k/l6najhi5ayraP0YHj
cMMkZ5AFnq9WhrQEyg3xC+56YaavBVALzj0cuv3zJcLBCcw9sG+XiinCzPWY8ECWBXJ8zOZ2tNCP
VDU8RgXrL4R6HHTxKft/3eIDvO96iq689gWI+r75KHYJykdJc4AafNbTVAfzr6cUOecT9J0eT8ZI
T/afKMyipqLfy6sVUUUrbVixaGFwTZIQvWK82INiFv3YWH6CIs0kOjMRiDKAdKeYb4ynJVlem1jK
HWnL86+/gC6I/pQs3ztP5qYVg/Hemate89jbynczYTjDjIwRTHSjDnSm2jFsmjLecdC+NI+Xefir
nhhK4RDVP06hmaKmZG+Cg6zCBa4NA0Don9BYrRF9syLa9V4kxRMdpMMeCYBSKDguzHDR9exauacj
vIO+fsjwbKQEQ3wfoAV9je0BZThV2SiSuyLpS0kCnuZPcTGMnCj8U9sPVmMJdXhB6ZLqWdXfrmOd
ICCpm+nBbCqlgCGfCTSTSl++vaQMMT1LBzJH/HtWFRyCIsS3xz/fhl2bwe7U5rTcxgj/ccLLlqjf
0ebDXflFAded1P1b+OR/gwngNvLO+jU8B2SOkiyBRGClX6PTwInSVfyiaIQoSo5eTBi/ucabjlOB
8dh70vb3cepOfzsHofhYNWsXM1oqv3RAGNhYTb48nuGNBnZnbUBFIdBcdrA2C9Ex2V8X1uuYUn32
Pm3v7sI6GpMIs4XZhvf16yt/4q85qTX7iZUKomG2qY20bGUx1wHXJgMEsPRgDnPvkXiJsbKMfENq
ppphCNNVZLNuFPsQacoQkFXBxzN5zq3cdPEjbqPpbBhqH6mQKqRHW0mx00HpUODMfNmiYUk1ETif
iJUO9amV7cd3Tr/d3QQVUQB8psT4OPQe4nXvEbeWmex7PpbiAZnWceA8oDXl0RmOxoKEeeB7HrPW
dgdiEdRvYHSsv+Mdu7ToCf7warWjXDDXkDQo0RxcL/lu0prWtxo9LjIucrJe1PJW65sQhwSnQhtz
U2f1svz4Nn3RrgL2jhuquEqnfd1pe2Hjk02DEIrVZm274iCbHfQEJZdKzcEZeUulwjROVm3dJi4I
XKUE60VhQiwrXbM1gVCGHOxH3lAO4wtgh4sKDhnUAVupjwu7Jp7/OK8ldkEMwM8UH2jJ9TWbWC57
fRy71ZXq1smP4J972y6r9iWK2TgFnVCTqCIPlc4beHJIh26FwqJ5IxrEoGlG//llySC4EOL9BfML
ub+MwoToUHzXMR51BfbQZR8gkER+7oVcwqPn6ZHgFIPRzXq3vCO4accwm3vZYLGLYNcT+p/LZViO
MaffOpeoTVJxJ3Zive/g2V7BGRqO2gxSkV6gnlqknplaRk60q5nu1bc7PH2xXrB69EEZ9L4rRYas
XlF/huRYL7+tKmQYhCcvzKkJJFwSC+yIsniaLl/1RTFOnQ03BZr5bU3m8g+9rI2iSTeEt16RUOeX
CeRMD7T+G6VObBRfFwFbF1mEH2XYKbIfCY8ief6TurQgiwMZfrqd25SAtTMV0WBH5g0BjjuW0LoM
hR6dwfQeqly2oFmcio7jWG44VKEzP/OodRfD06UScLCf3Nv6vVCvj+BSs6fxtzf0GO9iDXD+v+1A
ugQfwsEYaQuT3cAtcrG9spNvHzIDAPdbimYw9EchqAHlc7PWBTS6UtoEkAaFc5l4OR5w2JWaXHE/
AAyyd22lOMAqHBysz83vDONDhoMllPlnQAxc36p96A4UZPIs1gCUKYLFBxjPXDLXiQj0MdvDCmpw
tGXHsCs2TxOEYzTDLDD1r/+LC5pzEpDZjTmXlI8bW4BHqVRl3+a30otDUIpFpklmZd9WvAgdS0b3
VlCCRzt8VMzUfqKvEFS3bk8hAY83Z7JfGVTBCIZQMrudyDx+T1ApuLtn3o0qXFGbS2qMmfjgHmgD
RjJhoOFMi+aFOOOMtlpaLb2Nl7E8xEYyNJBoGMsp9FQp6GahnG2YXXjlxxTrewkf6XnvL7QX9DQL
2tzsEE8hQsWjn4wZcGcWOoQCezdkydwqmmH3lnxohi/7RixGFg7gpvhuFq/OgmXrqR0WKSdlg7Ud
W+B7qDwQh48M3Q6Jz2t/jp4yzNiquR8TF9haQyYSD5N1Gdbb/iTTMkJniAotiVH9HOkvyS3jmzai
ApRiJqoUl6B88yzjm2jonTSqZ3nx5IcYAYHNyj9LJNqashyt1Z9DJEt2BIi8YPcKhP2Of1JTTW9w
B9CKJfMKEh5mE3t0KTSBJ00LMLqjc1bO1KT89RXpDWPUPBb+Dvs1vVcmRLuFZLiLWJ8vmluk0RTL
lzOdV1zDNlVqTHE34O7UnIpxvTtRWQIvEQMI6x9RHLqVRq9Ukol7XzTQHOTI00QNHu/AuDoWMcT/
AycNIvFI9IhyzVfcmog5JKtxsJ1T3oBQ9SVvMiuX3gdbprsEh+gVtqMiCNiRVGWX6YC0komuS11a
5y79IpOLxRv94gwtO+O+FCdl75yeYlXiHsMtEx6etnQsa7y1G5ylnaffjGYDi6IpQugtuV+/pk+E
xoABye2uQPq6pAcSNW2XrGqGDlVRgDa6ovKkEysRqSj08/fKm7QHoYoKbpPCKkAhMDJ2edc0JM6F
QGNYIMv/7ArNeWFvWwKI83bh7ves9jd894nHpgvHNqGawo0R9yoAzD8sUPEULINotFLTTndblq/x
MNa7wfAMFI5Th6mkt14KZ87LFpGeASLhjANfTn30KBi3atBBQI+tVIgyPTKYzgqLz1IDRBBTFweY
IaaEswi2A8I2LLje8l82naxZf1v/aSsiZTmscOdb5oUBFSNNSmGSupnu++3q9RX+4TXs/NqRHYjQ
eJEiQL0hEAwwNNUY6gQuKtOcxAwvsBJj2bo3RfYWjpaFswtI9xlKakwN8PLM/qJ2QXBxmNxye5N5
/HAAj9yq3B6eNOLROMTN0vBV7i7l9tzfbN7kG5Wu127S0Er3aNMt/KJF7mLWmHkk0P7yc1aTz1O9
xRklTBec/NU/Inz9GQPonWNfo3O6bxS7AOJ0YyG7n/+yqQCcj6mGvroTtWMlQaFMY1+WpTjVzD2o
IIemxyZBO17iQPlh2bvYXkK2e75B+vxsWZFjnMmyByR9BGaXxqSChssJJH3Gcp2Ua35l9t/GDE43
I8gE3G3+kAEtvv1M9l05VQeVX3MErs+mab5BRsIEW5bVoCW2FVTZJx9kLFNbzeEY2Jxg0JkNqSKO
USffg7jkaRiSYSWcCikz3n5icyJyQ/rWu5QjEfSy2cSQ9x4UiheyVhTF/xdMlJHADLA8X7O2l/wQ
2cD2lwUAL/k/Mv2vm+Pc4Os/mr8SptOEewLBJOaiQIadmIrPDMKC0N03rRDVvzmG2tMkl7wAOdO3
ilbfiZyoaq/aUYgd6mzXNICUpJlQ7j+0Q/EneEyMb8LB5so6sCnV8lbopiZSh7/AW7pYFYqKuig5
iZ6mCom4iO93k1xNxMjmmiKXXopu9RgODR0YaKcPFUoxQew9t1OdiWIwyj31yOjBZJCOBs9JCdmU
RNCPHH8hHBkuYgx1qgFKPIDDV4vbHCRPg50MUgqpQ59yTjYuHzttyjjkdqDl7p66VIacrQeLDRXG
53PYWgvUG6sNkmxixZ3CVFCI9CPDIwGDtauKQfx3a34rvfkBe+pQ9lSyJL07uuNE+byMDOYqYHt4
1ylo48DwZyLuPl6B27dMrc1Y90/pgii3CKm+xAg4uALf3+7XDO7ccRRYV7BmsPtzLN8IQ+8kQfJa
6qKmoEQMMOG3mBorKKoEwW3DDw2pTfHq4jmfr8n0P/Jdcvtl/5bOPgecrWRqdfFozQbP9AwLew==
`protect end_protected
