--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
LiBSwu1dVdOnzx8jQYCb/wQvVYGBAT8W+3FDG02iDHRotnW3NOXuBf54GdZsg45+UxDKlXfM99+h
vO1nMToCaly1D38Q8QAOcWDy1GBGQvmfE3igHyTN80aftrGZr5drZzcj/4RwizJzMP5oCD9RsI6W
DjVCU47+6GMeuVP91pnQciFdFNf5L+Va/8YkA8pkXdAoUPxi6l3XifkRm733XoVxDSUylKvXXPn5
XURzVa8XoiWvOC9VZDNruEwhbRGI/UhgnxBDE5IpHj9Dg8eK4mj6oQxMWC9O5HcIO4o+SYxTSQqX
9/IFQxpSZVFm/ePQRetBiEwrzUCGo/wBkx6Plg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="JplOrkUs4L2tuzeA6E54W45IwfdszfoRftrv9wHJRT4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
RtR4hkm0fJahBc84hav/u8pHQr7XGoPgSA+q7kxH2zHHUHRhl1OwmYajQpsKMbUKnxj5miYkf0TP
V1/WQpd4BIT3mbmbDxRTc3fpjVUuuUErOQqB4xKPUXfOvg3260cAUG40NNpXHPQfXGwtECL8R2f7
/th2/v+RwtgXGhLyPZPS3cOwGqdmRmaIiwy5b6BibAUEgvZHhHrWg+OAOuUrigzu1+IhShodfnpt
eBqpn7buripLYx9C6WHN4teQvKWKRmsjP8OQsewPTMQuQ7JXwgEhhzYGA/8/vZAL/EHMTaIyj568
888gTocwKeqSCwQeZ3DsJ71ZIJb6Ybe+WZnUfg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="j7jtZG5NhJiXPEoLKGZpiK3FTG3+I6S7a3L75mcgPOw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4480)
`protect data_block
DVpIfTAk1bk3T6HXM/0Xd86VScT0MMLyaim5Y0HdjqRVZ6UBQt/kPOw9PqV7wllFo9HY9XVei8oN
x3gWAbJ60MHO8j6I4AuY6/DSBcbOgb30j5mWa4PjtpXBgz3xIxLX4Y/mZnwvbSDuLdNHSPmqHcZ4
hbFBMGYEiB/CbYQlJ2dt5yhsMBZK9llBw7f4pStGVr0qQ6JAxJ2qKInAjACwpexYqtcOqFv8quKM
jftBbmF/9xu8s/Gw9iUDvKP9KZ1+O6sQSQ9nKzodwR97Ovwy72KfV/jYJA+z4lVVu8Ywa93B6eVr
WVKPD/6pd+5RGySF5G44yIoVBumL7kAcCuUhG/8o+QFoAraDLOstpJP3LMBnlKhJz2xseAz5yncn
O3cOJ6FRzr+B1r5G0NhO+iZNasDzPWx4kgeO9yviS/Yb87JRzVExZXScp0+YCaDiXjZAnkmvIf+b
qqBZHWMMgPCigLy9yAjBNiiAkHmUmjfg+9JLB+QjNttMwMLWchqn898zkSr9VI6FVJKfcYC3o+rt
A+eR+KJhNSIaof/GN2eWJOtWWVb0wLExvzc+krEe6mJFzGeI+zUgkxdRSfuUbew6L/UZ7pUo44UW
8F8qkTBYJdC66kygd6sVJQfJkMZjdXy+RXfVBkVtEoQGIXeKdI56QmuD/H8KKtsReevrAhW0G3Ck
EVixDAA8MSe8wsd/rPJLdG/1XrWTv/fzRw3h1eMwXGQtucVwlokcE0//Jn7Igwg1yi9vsW/OoHzG
Pfg/P/lE8++aqW54tMgdhgUtgZlkxAY1IUG8K2B7cvcJPanmhO4ybh8wr5kzeeHX3zkwv8K088Ep
ToBs+VhysJViYNtY8ZaZOkJEB0CpAAkXRPLkXbO/TTy+Ehmb6jdXZkjFAxPrLpnAzkZVcoOQYPiu
hGty+HOay9TMHO2fUgGTu3HCxt+VlibEmFQdDB1A6FHNc9eprdR3c2JoCFmN1nGiH0Q/gUH576go
CCtsgv1W6yfGvVKtY1KsCLvGshdJpyErHaqF/zyBt4aYt+k2/hPhGzgUUGMAc2Gr06cxhH4Bk0Z/
8AHynVjgjzd9tRDL7HKp+vuqHveyDHN/ra7gIE2NFQe2J7BiHp3ng6vDNsTS/gAAaBITXF1nHJ1M
1FQBb3tUVT+UMnWwrReV9SYmvLpCp0JzU0Q/7743vJzLuLidv4/pZNFjYxj+q5E11K8ZaAAkR10o
0usK/PRF1QPrelLUnMS5sG6da3ATIFFNZjpWqJzpwWZIfT+gIgOUzlvK5H1oDlKt7mumnl+vo09Q
/OJpj4dRGZQT7i98DV5eOMtzehAj6zZyyAglKjmxfAWh3wjuYoVPOrFY0WFNRjmC0xWA6/Fy0dYG
cVzvG9pMOD2+hp0ObliDf1AeC1wdcxj62WfoeTOMHnSgh1gBEzUAVPlbkjKkFnbsj1qszgHqxdd7
gPtH3/PvQKMgaih1cvYWsjb6UjZLBSZ1YfW0aLR+cbr8X9Vsga+cVPNrlLJ+6hQkc97v3k8KJHKW
Ww1q3bbCv5xixTuv9gzyztdr8rnBlil+aQ5FIbtbmg7tUAxuF6e2YRR2IOspeKEanscyTEYUciRK
ZR5tFanYX9v+9r9hU2GTySBNiQuom5ZmdVbNS3ymUXr1JojJsaGquvhM/1qc3vNwZnxhFmoe7B3W
/hww5EwLWtJKwqHxRubfdVNAUfyMcgaDwUcYti+z4wYrE1uucSVLJbT5Gc+bbW9C7KCk/3v3/v0X
K8PctQSierMn4AzOH8syQXowD0WeApxeIE71h6ADzJDoDOR0koW5B8a+11Br6tLeqsuFN0Xhb7oP
dVzCxscPPEF6Gx/dLKLOO4e/sPkyyH3ay1vBEztYA7QXQzAlReZAWXdiOogrUy3xC9jXBDvbwvZa
HhZgm8NBZzjKt/7w1++wg/USq96fdTx02iUMb6SQUnD+xZteXbcZoI7CHpo8uOng+wcJ7xY2lajX
G83ynBHGlyb9Rx8+yYTPc9+WIezAd6HK4I1vLrCcqgpavrWTVwrmQj85a4yedzltLpKbD/AVx8zF
vrqwfCswVAVhZg+I2DTTgB1ZlQhB9d295iBDZInpFk55e1NELDBPFvObs6+ADhTHb+zuFkgn//AR
/2apFHKS+u7FyqmPHmpyPF56JTpO1l4l+vhh8CIV8+ju6oLsCFrnQ7PgOJstgfjTWCmNMSZGHIAp
wcb4k28vsxQ5c+clgoxtAZv2QDfqUaBFbinUj/TtWzt/LnJcTnYeoWX45+bIQtqe219RLeVwbWrv
BAKAi4gvTc4Q4p8GhmHcR+oZK8pcftSmwhJqBRCsHeMyMGxV9Mrig6K4wucbAnFlSt9u9hkHCt5M
OH/Tb2n9+rNrj+j+Bb3MSGb7dRZdDm0UsoCrNA0POugGDPSojLDBWFQPwfvZT3r6IzUzV3PaDmwB
QNUPxPnrck47GFEtFp0dGN6vALwt7RN+r0J2pX0jQ9KWP9UP96fHpLXCVy8P3v8ZV7Jh/K4dImyM
wMEakSkPTcVKVuIzEyPvZDJomRKIfp+3BUrvkzDuFV6HrZVlXYy0/zAB49hGK0E+DHavNTNtUg9d
zsTAtcLlou8H/0HY7PgR88oQTykpADrWjdzNJLyThXPxH19yUBWX6P/wfTHG4IqswmHtuSZ1rI4Y
J27i71JchXM4UUJa/OCw7sKv3Fiaj12FBcPDQ17ZQI1qkjQnx/N27rBVEgdduUFYTmjID5NhDyCU
UgApsqoLyESqX8UxgSenTfZCPVRr6UKsVEkcXOfmfYpeov8VfNOYIt0rj96OQsryq8o7GGNwtGwA
hItJmtxk75Ymmf+RL0jFCpWWPjwClz+fgyoDsNRIc1iWSHnfQdJ5ChVa/R+S5plUcFg/hmmdS9gu
G3WtT4b4plmnLvcZzFOZZr1pIoZ380ZbgQUBuZRaTMStHActmSGkWHphEWf22E99sMW+AfZgOeRf
ny2WeeMMhM/q6yttEZwy5nAUtdeOVsG+X53eUiFvYwCZT9ZkAsbUXiNgZ2vbDRnwDz9rZdcTrEpi
PG+/MqTG1Hr88mTgI5lHOxMkbexkCue4A5MMZOSRtAuCEYyWMvzaUXK5i8ScC3XD7ww8d4TPR/uW
/wZw6a6JdAXJCfuYp7tXq20Su35WfxOKMufnpYKauH0ST/gd/7wVhgs6tQeqNYtJvau+FZ2Q4nFn
+r8k7GAXumaGm65xaeCOBaqOCjS7ZVueIHyCFIUmMdyAxeQxRwiFEQYZ181i678gYjrlNlIPJVMB
pp4zfmRC1qWhYg239PAMDD6Yk4ICSTrU6yJFtaKgBs97VmqDtRFu8nuhW21LzfkPYzYSJEwfhf5S
JmWcXL94E6QH38WNx//YVFW5t+YnST4/VaJWG6kAlFPOisuugShS76fcOz1fCNuW+7n+aGXArJI5
j3N+Vw9DheeKPkazTLTN+BXSOQzyp9PVdvmZAJ13WX934n6pYE8PVlAPhBcsWPq6bhgdDYK7caDF
L/ufXVDtOuBjqt+k6ewwNZapdjeOfbZMQwml+igkx/cy2JWG2XPPoL012hIGP1dtio/T0eNqB40F
5kQeZp/hHl0cPjgLx6dtR06Sj/25q3R62inlDVmNo8Q+FSQeejVqbbEIaoSNneFEATwQJCDhxkNl
EKCwrKWPGGU4QMEpoP6/upEFoPkpX1EYCmRO9c7i1UpbN3rM7muByOW9nC45kRL3ewPz3JFUrKxV
8M+1Pfrs/e+Owzv70NakaE1V0Kdai0mderoL7RyriuMYTe5NZfsv5S/OmA83oSKX4TN4/Cj7UZ9b
/84YjdoCdv4/3Qn2CYfju8vrU2d8Vnckpfw+KH0u56j6/C/WoZSu40pXY6rLuK1GcntR0hG3pdU0
AXVjl6YOe5lgqyzoBucxNQHIUEDihIEMe0UyeM0MOl8DQXJ9xn/aV32reWgWxc/yG02JL/Az86Dd
rLa6dqxWvjJ0HE0ZU8SWXyH1kyVjlEZmhElSHxbnZGY4olqw/KanNzwDYFod2TlX8DC+1B/i9fXW
qs3Ayyn7ElDbeMqIxYi4KuCddGXh2bXniqHA6pJy0/YJiI27eYq4AXk7Gkft+EiCLdEOHXYlJYF5
frlAYA4E7Y+Q4GXofBkxtNB5VxkVY389PbBTgCBbYC0/2KnLmgONMyl0MruUdl4WLEAkkyZXa+UD
hEZOmvm9X6Afjx7J5K8puHG42mbTUrmZkE6eVS2yNeM8MZcSIw1vy+dtngEy9CVGAjOieg0dEaO5
yaqkbayiHSkAOq+0Fk8wqmsgJqKJAbihRj8+ivSrKORVlj3qBxYNO04sI1EHhpmpJmWGf24q6Vrb
Hhxi0FWIMSD/N9El9rdNRM/wIjUaq8F3Q3ds878QMZbz2rZobUghrQUQ1sCHp5fCWhr+Reg7axYf
AAyQGcmd3URBeKlEnCv7k6x6V4K7obanxSfU+DvXEoi+8NzTW503FrcIxCmrEu9b8CEH80vr0j/v
pRtVvpnhG4DUdYWVsnvD4RP0+0ubDeK8vFGWsc75AVHiNLwO5FbyeNCYONc8Zgl7Di34m6h+cdhv
kSF3PA8t4Y/lNmaqeYENHhGC0vDXaW9qi1D42KzUI9FU4mWyLQIyKTIqF5xqt8DhhOf+ptC8Jjr6
GTvYOBpeTBxW89mfopK1in00WHBa/nH9y2jWbLGpfMs06Ld4vcHHn6tVA8WdECfbhtXPYmHifMHW
WFWvByj3wl2A6rJ/LbL2DEVphSwoMNMIKzc/0uAiQ38puFrtIGy/4V/+doSp8s0AsS+8fnA8/2cE
t7LkAWO+EbTjqH2RuBvX6/N9N6ObNMxNq5xgw5XSq/KSg+Bn9JvAbHZgG2Wi93l/1i5J6nHee7EA
s5Tt16JvsAbFmceBoYJV0/BXc0Ag2YIepeyXXebRoCBBU0FanddPEX67MqJ93xEIIdrPVFngBm7Y
cuDR4r42KLxEadrMpDOkf1WpE0eTeEkPb1DC88Kl6kSuRd/iObjeuvpY1ZHtLiFSHOeAr+fBy4gM
7B09asRsurLOA+UGVTndEIlgIir8e0eXYy8soF/3+zcNbirt/D043/DUYJDKfZkIbVGzRlJELyuy
6NaomUcWEmjte9RzSrLqXb+JNQAAUvQdC81Zi+zkrCTron+DhBZj3QYITSN9TibI2Qs6IOOk8Z3d
/kLTW3ArOEhRv/ZR4kiHc/pndSzYG1+9mUBV0UhXp8r+E+mopQwAZ7kQwPj+PKAoLTTdNGy3j6aS
q518iK1XtlY/RBF181kb8OyjJRxhS+vz0vBm9Ml0eKXfw8etL9pyIbrApCtKaybPhhI0lnce5zZH
nIAmquA0Wo6RDLMmb0Po+PafjbqUnhYJep46TIBZe1FItXiAIocYqoz4HmEYzUjPuPTYIvvnhhgD
x28Gj5cRtMz3G3xXVeGMSuxiwK+/NGYKE28KVCZgAES3rojPcFVv0eVVcDbfaJN2w66/GWMfHTky
wAy3wLzGI08KyndZ+PXQpi4E9QmF3Kyl68mH9JJtPD6SRwjNxsJoLGZsbS96gi7xKJk6u6JNRcLH
dq5nkAGL/SkQ4EBQhnOhf1ahIG4ZGHH+l/BXsx4IV4TpQm1gZs8+QlNc0ZyMaSmc3SAjE2+5KDLh
AcpLQX1CDca2fWBGbGd67HYIBtylGaDKcFmgHgQOnuFSNBeTY7iXRAV4dSO4s4b8shmWlqjnaxdV
SGeFy0G1LiduKip0enY2FbcArId+fMT58lL+Tht8sXO8yYnDZnFdOF1TEfsLTRIKZcI/fyyon29x
iouGxVkD9V+7L/LHUxvLln69O4C2NFCswiKpJVkDVINAX2k0YHm1N4Y/V6v1WTFBAI+bTGlI4fn6
3phDT7CFhzO8LTPgePDvkrHcJkSUsBzZSB4m0IeSbQm1MQhdCky/T9OFdI4EulzUXpSSPAdH+DYn
Revo9gojCA+Eoiy6/aMw5U8f367B+CiJ9ezQU/SZfaJA+A==
`protect end_protected
