--------------------------------------------------------------------------------
-- Copyright (c) 2024 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Maintainers:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
bYQavKblBYmgPQ2EVILmZ7q6xIRUyXxAG1Wswzlf8zG/Czbf6QkBb0UKlIItc7BOa6zZnGPlr4pc
mlYH+TKZrYA39gjEnkxuHsWaGIpbzvb1263ye26WluA4YuX/vUutoc3sgx4Gai8WCvRv/EcvrWog
DaMTtOhVhDrnMF1StLpq/Ji6WyQTjpS2unm3BsMQOl8Oi8M5jCNqeZTJ3wPRqzOPU5lx09mGja+G
I2zL5wblMD577XQT7l9fyfN6NzUMcRJQ4AvN5KnFn+jjrd98bgU9rqXdjxdPSYVvjYrKB+oTkYpT
xURGIKaDILL7byIjJboxG2EgZmW0Zapg1vK0gg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="ALuynaY1UbJELErKGKH0Hyx8KnK2v8suoM7UHmsIavc="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
E/WgiZQvaWKKn36315lkSbA+0HboneJSOCgInYMmAk2EOMCgD6u5FFkzkcvEz6Zf69Ec5dmFlAb/
JVn22q5LnmkcbgkIv+I4ewUAhLxnRffX6ldm7swLNPXj/KAHNlNps6PLEEJCRfOVjyE5DrxXrzLe
GHQ0qVprjpunPjJ0ISckC7bHbd+qt2osRpZ0r867IAgm/uHjOsphhbhTO/v0oR3qG3paw53hEhbp
HuLn6bxVtSFSN874phyU/Xv0gj2bDJhODH64XSbkvCl2TkQz0b0czE6COaumvAZWlfy+3SrSJRgw
du6aWGGpWDzcOm3NHceFAEnVTZV/kY5wvCMhhQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="w9qd0Yy7QKEesZGZmbAS+4npmKq5P++SToZwg1IxrrM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3968)
`protect data_block
hcQduJ55dCsfCAYeVipq6M13Di/TqGZ+yl1NnTp0O+yZAIbsVQORG4zRG224cQbpgRbl2e8zrGBL
qkul5sQbz355kjYbfjT06jCIFJvSOOLdb6ZqtAj2eDwdM9FA1yFklpkxaZV8xCJHBCFxEXRupNQQ
82yO4L7do/t1J2E97sEwp43GbLExGv3cnrOUiKBTmy58v8vuknRKlC8U+MJzw0uKP9g4p7zu7MJZ
VIQV5AZIVnebGt4Bt6KhnfQoV3zFgN4cHzCugvwMuQRjGMoSKtD6D7r5zOatrXjtpEcbVzbMRLuk
pLtFv6Ibh5MyiJ4NoxajwGkiImQ8pqUSUcLk/Wg1dqERtszC0/tiAuBbkC9vATnTMN3KAZT2cO8V
pb/DVR6ZxgJdFRsmUQOI7IJgRwmHg0/lqLc3rhtt7zx3fjUdA9BS/3VnTuMKpXoyGGnWtZrjw12N
xfzA46VTOUJzPtovzgbCL4oKd2nrfI/cGxz/OM/2+1CtaeSAbUWF9h0ea2bxMjP/WMFKh0lqeLW7
Yns8RN/K1JGnl4NCOqK+VJ48ppjckluc5DZswdLUhioN13Pqxoo/Gk9uzBayZ8gvjLuuo1Im4NUn
o6l/PaOYPiWC6C0jpz5WOQsUDyths5tCOIjv1Yn4SGqQsVzBYHYUnSHwUombw/Kp9DAAqQySaZrh
ucMNK5yKHWldmZyfrFeIaYRVXCP+Cr7u/2Gx9F6m0dMYZPUuiOSWKLGmQhvFSSbTAWpApIoXe8/n
tH++jiRTxYPbpqAB0ZhO+XW25OePvjqbBJ4/OWOkahCVmpKaDlO9Xj/AkpFzp2AbCOEGrUsVbVfS
cL+7urCl9+EHWgIiQPSWVHTlF1MPmFh13JBQwmF5s2+l7MbJyKmLdiUojW/YtYEb/nufmykcw9UN
DoF8M5zZ+CE26ojOGY0b9Wk44/1c/8fB/7BIdjprs3hB2SPZzDepKHUbNP2RdXolNksOPymnt68r
VbD31E72ds5jG+NKfTne4AVZI41ACbF6PAGZp036RoCbRtgyifEgtn+diwjWCi0F5IcmLaHz5fi3
g+oLb7sWGm6T12i6TwY6DWezdAkloEqplfL2Q4aOVlAt9NdJw22/vglNfJ1kKTVIqO07f5ayOXQa
+AxVYO1kYkDdQG0wS8noEcv2quRBPZ9vx8Km8WIwN7hy162iGt0GU1Nm4vBKASWWOk0QEi6qni+e
3dxIn9rw6itxtulrw3eAVDwHDYWGQ7KQZ6pG/ZIMsouNXK+Cn73F1CSoIdlcBddD7MH4iADx4IWK
aVsfVPqZLpWeFlReiO+05zFuNHFoyn6XJfQvQrbAOGnVdfADr0/AW19gdK0cLlMl6sGG67nDTaNv
CpWpWugFdjCMqiJfbuJw1y4hsoiLZV8Y1sCYsqb6CaiPZX/j1DOT5IERYYFz06V+yfB++ZjsXchY
WslBoXQQMCd8mgbSm/tK3rrclUPOtT6pv1QDF3tGFIs53gRJ+f2+5NIa/zZCqFJOknLHMZndrVky
4bVqAVgxsrI2s5Qs9yF6E5u00DNv0Nq02kWHvq6KEs8UBhdqNa0A9Lj+oJWjC3k4IfdO4atCn5JT
oCW+IpHs6xcL3gnbmkHQyppoKnqCO364gzGH+S3V8hPQo+KlCVfILdGkrKep/z7Z2q0DGLKp/uzT
12Ai0ZhqT8GFyXENffuaWTTQ8XEXUBNVIW6boNMpDbrI7MgfbI+9bO/rff1MLMsFWOCOv4KuFuEb
RcXjcYxNSsf1ukPsvfRe7V6jbKs8d5iUvb5OV3DN21msYr2rcuTzRgddHoIx/3CwFSEsxOCWP/Ux
WagI2Z9jbeI55ii3kL96Aj3zI+2vgGdHwDShxU2si7MHyq32CLgtJLt5zOyfKCvxSUF2XmSc84wL
/owb4iyUrix9ibxWf8fGm8g+dK3n3yXqGQh4KoffSbtJyqJBAOFIcGX0FNumIDLVTKn3qqbEqiAQ
4xjRpPgDW/MsTJsBxVdDo5wfG2OPYecMSoYidZ7m+430d+W1NUvPQ+jTUX2Ed82XCmBoiBBw3mnY
FIHZrDwbxJNrDifD6bu54Zdl/QW7pgR4Atquj5N3/HluhTFEQU4+2UvLxqMwiM09ZPl6yMgoN8XU
d76EKvrK1EKWQzFoJMDaKOzuDCgDWSJVoWeuZn90e9ay29HFDGohi2YWjcV4CIzxzIB7K/s+GY3k
fFkRLc8zNk2UK2c3T/RFLiMuN+MauGEZV+u3XyCLyQLS4SoyXj1N/o/FjJVQWTiHeURryoMhMSS5
QM0/oi4mF5VVdMYwjVg4dvR+EFCgbbzwFiH5Dku494YEd2EJYxGMCsUShS+4Qs3mHl2iOJG1BbR4
fB8nsQsbOht/Xyomn6YdcnyXdvYmBJb5ooW+T2lS92Vu5AWBvmx0cM0//s6Uwh3IZMmUmi7Eavec
6ldANBLOMyQ07OjLnlYJGNbLVuqSUvWlMOqhqKMjimth8pXZbWaA/SUqqsGMbOkIWrIr4XyHHXrP
H/Yxc5puIM6CyeJJkAPEUg86b2GfoDid0dWSX81vsN6yxsVimlPlxiCCfkLng1+LYhqmC6SIb3Wn
c+dKfgx0yJvfzongpdO+bw3sNDXICH3TPzhwVHh3YVuhApa56cm85rQ6z6tF0wuCucx6ry1csEJC
85kaNCjFpHpRMdlpO2DAtjSQ3GbgowAC1XFAWDAuIJrwq+lO4apYckM6YSMirbqJXotJDlZaXjFt
t5p6hNi2LNSR9yA0iZa+Hr0dKrFbF1EDst/u5Pkx4iTZP6LBcKH5HhXiMok1ITzdcxxEPc7ow/wq
3YdEHiLEtpS40YOhtdO8VABxYkoH3q4/T7EICB1NJlpcaYHa8TZB5E9FI/ysLStK4B41cTI4mR4k
B1HT4d28yCgQd/EmJC5uDfR7Teu1O6f4KGAPkPHT99oVO0n/QGdi75vY9fTqdeYKER1bXKiWJKCd
WiypvzSXI3NbZ9A/J0Xof+qFrCg0l5ZHcEgs0m8cQ6r6/IlA6xae4jn7BdNNAebfMpKQp3fygOG2
dFaZ/r4P81j4jBuTZH6Z0KdWpsBwM6HBYbqKCQgA5K5qBqmV6V4pmDr7JdzHU2ViMpztH2S39zhw
Qzugzo0LWiQI7+JMp7yNQao0AmgiQWPdB2vSHxvrtDGyk68JG4NS/VjyueloePGqrLfbfN00uqQ7
yv+GpcgrVADpwrLbApupAuvqJpMDBxWWPT22y+Eti5up9UyCjTEqfP2gBT5zeHlcJBALakYcG0C3
xHp/QLADf2GA1u9voCA06TG6vFd0BmkpTLiBEk0YYVCX1+DlGTDHKfwLHxB/7Y8++zuVhPz5Zy0l
y98q8+bGnbvMKlvw3c7UtENd3MMP79fJ04KYX5yz/ZMtK2txuExLY6QikKyOFHZHeTcmg3yQI1qd
nzeFST3w7vK95/3tDH6hCbe8A22NfIXsWiG/iggvv5/3/DuuabDhbAOL0YHY26xj0h7bKYlYQmob
kRtUbsHO59u/fssUmdmTEQkisAa9WOzTwnITT+a0UyOUc8SUQn/n2ej9e+4PrDgy2W0pTke54gjK
IJnQCPUa4ih0/Wm59qtt7H7e4lDQ4R+U3RCW1Bgc7c9+z9A6jqsaEo9HJ+rj/4JPpvs6WIanoVoD
TnVa5UcxOUDsUpGsrWqNfWpKxb7HiGrNsFYhDjISRXM60gc6BM4+gHwWjOH9sjL76fhooqaPOwZb
IPMkRPbSt8PzQ5Kpwy4sjeBFGVSE34dbPpfPZqhQkVPJuvpNVrFHQuN5A4cegps9U/2wBFfTdOpZ
sF+Q+BUpQlxjteCsxm6E80X8leEO9WDUXDZNSNZ7vuuKOlnA5yTdau5KZJusmABRScVb590QQieZ
J//JkiTiLxUVcvQgLWbXR+V4ZqVqCkIYSoRdmOcj/TRXuYYQHf/NpIAFVdSIkKF9/oa07+M91nd6
z/BkTYa0mO3ZwzbNylmUadGvP0VhyeMpJu1CI1Nb3ZByRwAGGRpoETYhduYlKxdynLjxb6ne/gAG
8pdNHm3Lm3ovFYRhdx0W8NVJHh298v8hkTSRo6nZkBKAbwGgBc0JssM0i1uSO/5FLJafF3Pl1OIF
d5W5tmjNesjB/pcjvl1MOEw1d+yCllhzn37Z1ILTO0KewUglHvbKMQeCw7YLjHHWzwWtEMIk9pXy
k9xnG9W0TpjXNMel+B5k/PYvFavuESRx3Tc1MHIP33Evp8t8qc3yzXk+30rBxEcBKOKSmrk5+7Fe
/+oFLFbmVch+upa7rlAqfy4R3yP7Ccx2qwEYpMFq6nppnpSmGtouO62x78DU6dEHbTBJSXM9MpVG
WyMfDnKnk2O8Q2y7YOtAnw/O/DJT/bdzntlNSWonfx4lNdIuzA8liYthHUlwKftCB35nxzj40ntF
08PGeeX27pj7Uv0QWEh8kldIBeYCiARShTt48FyOBMrdVwrFQQVwjvcZ/iqtWaEeo+8auPg+KlSG
Ig7l44q2T4g0Yqt/zrQqjIrDVJ19nNQcXdCzG2fEIaRgNb8vY8JDPcyjvK2FIAgo0ALF23MDkLCJ
MaH6P+dSkpJXiAVOW4jwYzxoMfrH8v7wBuV2GW9raa3nmp7CbH8V6P2rZUW1lSmXt1DrUBa7QLC5
Zm4GGuwCEDODuOPddEbWo+WEUt987pmVUFVmQPD3cL2jRBjNSLHyBWlYll/OkmxHGt+tNPEXT7Uk
c0zBlnDQjglexhiLg7w/UAaitv7ZxvFaOlR1V8nfEbgdattyug3qd4Y/CvZ7x1GfHNEsVhMSY3YK
yiyKtGhjEBnpPxBJtzZfIuv8SLAItD0vEhVt/4cvM1a/OrMZEhqLH4eVElKl9HY6fx9XK5x7P8BG
JqzI9Lt0NGMz9Odu3fzs02Ffb5Xc8Hu6O2o9Yi8u+sObEdaPlAdffiS/VsGKovPqvceNfG1EnBuR
YtOTWsnDJobb+t31SqHKmcGECctoxt5ty2mQCwzY0nZoZjoQLfKJHE7XmPNZVBHb2ygKzoAYkwAD
KccPRrPA920V99P5c0OHJbWvuX+/9fGladQVizMVH870mV6RnhYroABQuYeDtAetpcv0oo3wKYN9
3vrRx2dVE+HBo0OBWm1Moe8sHqLyUJ0y57oXn7G9OFnkqyRSS8NBZk3tMeukHc4ZtSVm/7UCRjt0
ibMpoOrgYEfNoQ2b+/zCcSPvFJFZ1BO4UvYs6p3O5oLXVz5WxTR9f8yv+dmIEIdvywMizbNZvzso
o6It4HgTm9clvTXdop4K3Mi7o7B0tDunfEbbdQi4xu1qOZ4=
`protect end_protected
