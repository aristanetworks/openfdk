--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
SKPigo291Ddnzn4v+4TmbQ6iNS10hjpK2wLYpx8Mf8pYVgViBJaAu9a5k514gaPLMWFBLGz1T4oU
8XTVBNQGdpct2We6yAYuIliDX74MEQfkio8fBck0cgJkSxeF6SVELU2KxJKmXC06aJQf8fdFybzF
wZ9D8LmRjZiBBd8FZXUhaYCaGwBwLdo+KHHkvRKCvBJmIJXudQ13eqrDSkJJiLCkhOT6vIByRqCL
ocWVtx2kAWRMjiwDuOgGAfrDV0hdpVNEmq39+DzimuAcy0UTmLi+OFO4G2Fh7ZlGYFidW9YAW2d8
8AYpdpTOvTpOeUbvWewG9gUwnIWOIpM91wkSoQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="N5kn/Gg3neZvbdf0sFdVSzPwWiJPtz8pPJ3yhqrrhio="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
oM/k2d/Vqkx2eV6gRmZk02IRaHY0k9kZ01X0Ymn3alCQbz+wP9rCRiMB5WIj1Bv23sIID8QnB1/X
vHo2d/Dgag4z7fAWKp/+tv7UZZxfXpLtrlB1RkKxufvjx6oHoL6QJkjLzeaS0TKcQypYpqtzL/9c
UvNlTPqY4agMr1LKEa+HV9kIgy6hcVN5470mKvvUdpzDJpQAX2tB3hAQ5IebYs1SPjdmxk4+uATt
xRGoNGrOK3uBlqPhkMkz0KPV0MZZaTIwRKvgiCzAQ8cgwmw9Y/tkBwB6WNyXiiDpujZHLZuphxMF
h9eoYECHRJJ0D5atwQ/hBCW9pBaOQUoenDWGww==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="dt0aGq/PlDDPOAUdlCiqw9YnBmLOEyAd+IBZkskSZGw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 29600)
`protect data_block
0huQCIiW+3CtiX8FBAqytzTNxHmi2X/4iBCdHECB3SIAcAlbZdOui7Eg2Ljjipwbv8H1m4k2roCl
POm/lZBwpHjenU/FxKfcPa3cGCP9KQnmveG7x5HP9Hdyptym2wCI2CVAPPGxVHpCAiky1Z5Mw+/g
SwjdEo1kaOnsBWTlbi4+39PMZm5+rzm8WaNTCBvMKZSi8gzjk27JyE5SS7ojx48drrxFahLIeX/O
/Fla27iHgJfr8BQuw1m2O19GBZcBMCiCnneqqccX/rlOK4XYRLFm5lkeeZMeH/aCcsceYzW6rlwl
gm2AkyjxT6IEDHuwgEVqTsuDCxZP849/d1uOJHiAqdT6wxW5GYEt5CFxlC5EfcHiw3PsQw7imzFH
AlH0PzQ8Dc6CKl5xOPD4H3q64oKmnV7U6GDZLTEYEwbWFfn1lQu8Iu+7sGPnA3Rgn2G8pDvnZSXU
G0XaeS2mdwrTeQat8M7ua8N2jshCo50UZFhwkhN4WX/FCbTZNa2j/7NJ36ViSO+sbYNeh0nIiSvI
JuERtI68A1hixjX8BgA3Dh3qEtb0MI1JDTL/vJ8ICflqvATVjcZ8fkP2OOFgEWW0S2YF/LpBlrnA
tISV7OTqembURioUjrakRIoiFIMI2GRUKIPyOhDJQXNGKoIHtcl5hmUtwWHklILt3MPMcLG1DMTm
swVSUhw+mrpUPQ9zzq5AFECeh36Pw/heC7cXWmOkfmCcJSqCcSDxLVqqXqvnUGyPYsZe3QqPZmxF
njR14MbfVK8kFPPqg/c69fQGRy4Ggb+Mit5henLfyZGFG9eTFAkOCrlrn+Gwn2LATlAjcLL2m5dq
3WHKiVOcGkM0zZhT1ztFwGtLH8Cs9LdCjmVcVYXiUJs6VI3tWnRgU5Lpl9PzRRvwdU9n6slXLbqd
i3le2+JhNtoEWEE8lYEQjSqfcKyPkOzt/ipH1RaDWPS4BNOdDhCYtnvkFIR58yy3JyWJ9u/e2dbi
ShCXe7p8bjvpbPEFVJBHmwcmKPOC+byF3t2PQB4IDmQzXrjIHIZR2lHywOz45dikOXZ9ARXCSU9J
t7qY9PfTZltfKpe28QLn5qbzvwbaowPzTM4/+lhuK70pH6q76ZzkCh8Y7MvWYNhqvDGA8DXidsMS
smo8+ZhBqzFwQFPmWqQfZNmDAdORg1tf3pIkzpvk4Y0fewqOBRMznJPXWL1O3k3KIqh2T59bqsjE
ygKz3CoOz/67rugxzxadVhTSZAafHzrUKT52736SRGAbRd9sCrpc2WPHoRQI2SOCXSloJUSqWZS/
V/ScdI6bpLNL8gynhcWBacODadkKs55VusAxQjM2jr8aaioU7jvE1nLSiHk2L8VOXJMG0qg7so3c
7Qqqo1mzC64Xbx0Bb7uv6gNk6/UBzk6zhIQX5HWR+tCcl6xWSEnZZXHi43nHc8aCdzobvd+/JoVe
DUQ/oUlF0LFl1oTdQXw89gBX+vexWI8cB0dy7R+dnI8zcYER3509KcmYN6eZ1yhxamQJ4W/YRvld
+HX3HuZYIfhZe0Wj+gE8+zPyIdvXdmBipWBSE85tZIEGxqKtbD5Ers9Gqie/6IJ7GxLW0fTNALgA
uidYCbOW09iuFtu2zOZKqFhqs8aP0X+gk9VHUCwY07lf1a11agaY0uOjcOMi6R04kHacpsQ/WsrX
PslRweDzh/Hw1Jdswe0DYlJOMkgBrtSPDgd9BWSFfu5Sg0Qey4iccPTPr7PFxZT3KV4+kbqcA6fT
I6oLyF4kHvsdlPwhowOClxotMcjCDqE9uKibvzdk7vOP4ZHxa9sI0/Ra4z6qlaB9+ddam4QqZJ2O
Q5wImshyABhuJFMBYpePC+JR7jchYcWQsC+O7ntv17PNM5yThARC9SoOZxy/vhLb6vk/5tZ8wQg1
HeQY17LH+1xAxz/VwCOv1/SBj1oATTbKAKbQfH7s98reMff3MnfSAyTEBH2EQHtVsVRWa6Q5njEr
5BqhX4FhOB5mZV2XwY/epb3g0Tr3Tr9xwKKk7CecTolSICpvFiyhx7bsJo+2mEgohXec6RvznAUv
o24xhPZ5txjLuA1zP6f0dww2mYTGIabo57SOLjEhfajUW24AuAAqGgmZ+UGyIjRbqNM+zjhNChMr
iG1CF4zIYl8HGwZgLUMRGxAciA4PkUoCCmaXAuCpguiw5S8v+BQ6YzlGV/AwWBw9SgNsFdoV+fm2
53iKzvy3sx1OhhpASU9lBIQvx1RSTGYy4xTTaST3kweO4zORh5mH0xmqsBzIvGsxB3ZO1AIfxDN/
eDabLCYTqy7ju9xBh5o0jun8Mm53uRizbLw15Hb0y13QmrChXkW0S16YvrnYN6vIb50X6C4qcKK/
FBv3hmAbAKdCkEQNU7lOfchc770CNvKh8ktkYTDYDK4K8lrJ+b5XoQsJH5XW0xTnHJFgwezRcI8B
Cg0eip6EGzlmSaKrbXnvK/Q66AAWrrad1feyUTrC7aJq+SmhimGDgjYQsjhgMBvXebpqv60Rw5yG
a0/LQKz7jVlSpYdi22Pp/CO3Vcoj8JPwbn2MLKSJFrq5F2Tna5tQXNJnR2Ac2I8LvKW3LACuubUK
P0ug7oDlTk+BJKhE9R5gts5ecT85l4US7+YjAP44GNzwYrCEQMAnyVgmVni766pxn2Zsa+tgcx3k
Y2JFmwD3ZqbYmbHGA59s+00DDvCoLuQM63YbX6b87xjS3FvkG4hbvc5NTxUputPf7Vm7KOvS5+PK
HLnipP0YKZjJqP/ipZroViCZnVhDkm8kkLABB55LjYzz0jkgoGWDnW6JM30LCdOeEZZxVtQyRl0D
4YDggs/Vj98DX7cEpclQ5mxuJQtA684g96uZS9/UwERaihHYNuRNridz2tdVNwBgigvYCgs2yfaz
A4G+pJlrJNk9Vdz4C94GwaqC2vNTfnDacdyymdMfR8cFBxsvRuVTBqKQsv1mFcxCckqSq6phwMOk
siYAE5z8NxUCwpKJ+KBIOYOSAYJ393dyzOG54gxrRF8tMoBj6u4IaDFrBI0EH7UQnlavRI/GG/z9
SA+rGW0mFJriw6Z90FPz4AqIOip0LiHA6nRF519BbSQeXhYb0Ey/uf5H9lmUfb8qszBcB5TtJQSz
6WBTLXURIUQr2u2idpcssBAm6latz6Go222G3+EiQbGa7QKzi/5TCWCui6NZBU2s1jLGyuzpX/x9
L8qKGoI+rUkCJK0aWo+er0hV7Hhn88oGdB6wLrOaVlE+pIpHXbDUzZNImKl+ptoqBu1HP4aprhdw
dFqPRQQjyJPKGSu3t8vRHY6DX4qUejnmRVE7k2mpeQt331qMjxA76TmEf6GH8FbXTivlRqba8weu
MnrVP4VeSQXaZES0dKgK2VCl3tGrcJE0ZjDVgZ0OByBhDLFn3C4DsDN8hNlYZySCGW3SCV5pH89g
Izg9u07gxVDiT8EWQMg9fvd9HEHwIWxOnE7voh0veUvGM8tRil4mC5yHkFXRBckYPSK1XbrrmsK0
4p8OKjKXWVreMlW31/klcu4IF3dDtbSTOFtTCOnBvOFXEJC/mNt6tF0Y/xT1il3P5jAflS5bdJc7
7p4eOAAba8zSI2RNnJ71SBN9rN5No5WtBOjITOnLRZylzp/O4Ha+sLR0eQ6sGqUoLPKHsbtOQD79
gQobdzCE0McZDucIAiqSIE5UZm+eU+Ys5In7bcDAurdZLBmHrggCQb6/oE2FOUVch+6y40wkMrlG
htF1lUlxPCCUL2VKOSUMDmeN3vAEZRqHuzotJVX8yS0KjQLdMPfA3OawCXPa15yM0cfLHMrTi7p1
MdArGTOAI7EJyf9N+EyfN9B3b1XlrvRizws7qlR8ulF+Yk4mm58CvhkTErIlIQLNHcHnQE34Cea4
qCMdof0SRDzTOHDXBpLDATPNoFB6yfG2mVVSO2MkB5bnOKouy8pXG6vHAOWftxCkfUzMXicOz9yV
BS+f4evyb53BcSzcG6HZYKGrMnanrzMFPMkTBJFq9O3ADdLfQ8rE8mX+zGlMQEOrOmiW0GNQoTwR
Q+/fRnCmGHe6+0G+wAeIDF1jZiNClXG8RTJgc/ThKo5nVoOmXMlFx5/0iydQ13ryRQ2418llVkW3
C9E7LJznlzLdFgT2nofSesM+hCM+Yk73GbdtzGfSWnw4z4s9phqmVcrbT2B4dwuMJOlnvLLbH7sZ
XgYZWaiz3gnXQ/AHDKVY5Os0ebh6UYGcWVgjlI69oHSH8a/1B05Y80XInfjLtgGNKD5URRlRZUde
LUI0+6hC2oEjIASEpyCK2TQ37vSGjp01dFElfVKdlr170+fLUen5htkMLziOOe9jOPv48jp4tojJ
jju0/gfWK76tpGKqrNnukx0qzO2cZof59Rtg4xcpwpjupD1GAA452nMcbts3IiJnSNtchIzFAfAg
bI9ZuHUHzS5Jwo59O39CUw5YucW9wKiQbQV+a8UZkbQRGb+PXbGcOES3ocX4TiDahi9yX3MIQxqa
/oF9Z3DMDbtI8tbQChzPoWmrXmUDVefE1fMBpbGm37xXXyWCbjsf+MQkf5MjMTx5reE06tpmkc4U
RkJE2KqgcMmhhQZn++8i5523uQdCvdaP7+hm2B7PMf7Fj91L6vwU8Ncmv7t1AD4W+zSUOvZRpPkG
a283WWkLqrPFZSaDX96DFH0IUYt3gYq7EBMe9BzJHqXN7to9eVWZECCFKFi5RL1PrxZWenqjLqAr
opudReEA4k9QK0g25UbfGWWj6Ddey/bwXmgxEkU3OT4ozkWUVM7ba76U+IgV0TL+XTSdhT1xfzsK
CYvefje76POUpTYy+sACOfsy34QsgyR2+QrX2ARqpHkzZ1ns08hXP+k7oEbJjBP3y9alh1So8cHh
m0tWTMxO+VsImysJC4yU77qZxyf6/TmoN+CmdOeYMcd7BSg1/Da/Ca+J8rImfy0NRmabFVTu3xuO
80J+/17VJDyGxIvXUBsHZLa6bmStsD0jY2RQBZKKoej2Y0jqmxHfolgcv83U0+6DtkDw+K6YaVj3
PX8oixS7I63pSe/XSCLSmfOyweegrXsk/bglh7Ph1z4LvCJXd2qua5Pb3WZHT2iPRHOdH5UDVWUG
+1J1o3UdyHeOiKMOsyCkqyrI3XkxZpv229Xmy6mlNG8I5VH6DXjS6UwuMYiX77nw8Zuou/t0r4nx
G9TPyJrfDRe0VrM8l2kd4T4CwfjoEfZcYSfMejWvYgzys6IiLK6oYRoqUKFh6o9CYQ95tEbokLCJ
U9NSAopv+JkWDTtSdwPgev8Bpz7F378T7RKan2WABbd1mYuHSy6T4EcccvJItiqpH11tZvat/C1u
hIKWtd7k2onKSyR0cMqADfotU+fp+qWNGhn0F7DO2nPS7ryROdfIa2ImfeJXbvB5FPH4uGU/tS0M
jmlVwAGogbDA8HVh1/t6ZJkMcq8hKhXDwjiC2HOBsg86gS4G+yshZ6GOh1HLKjqtQrYhuAxDXRhQ
ECllqu2ZOE+6twpub8nKeXWgbm/iASeHXtDeWOo9DtUNDCMVeNbkR5udmQUMkignEifJeeXv3SOC
8HWNuA4hvVJ8Z6NzHFcmfyhCnyr4eDgfxsjhHM/3gmfNkHNvoHsexb6Z79nyuzcH97JAb4qU6IaY
H7aC7WWzOBMNWIB+90GHEP5FiVPr9gym02mutFYdkUjYGr2jUjzxiIPO99OS8IaoEz7kooLJaq6i
M/aavgTySAYBqRrIvVJOph0WmRCRjUR1nTvd2XWZHP5rg8EPu+bwUXaBE+urWqq/ROI7b/sZP9vM
UZuDxfCysXd1EE7IDd7Hh+ILTpJo/87L4pEr/wMlQgt29zXlToLvItjce54ecVdANGOlXLh4//Do
zqbsIds1+7Wp3+MiWxTuTrQsf5MFrrNyjj6QX04Rw2RyjBfAWnlq1yoByjSZXL71SH0jZ5+s1/5x
ooWOby+4YoENBkA7rsz7X7Pe9ab/HbAMvDdjQ4yF4dRLi+9zpdoiCS8GJj0FK87cL4AF4+MJfuqv
P9lS/ginHmvOm9xg59Y67Xp4uquFZ7KcP7gmiOKEI33Bm1qf6NEFjHEuU0TWm9y95K+lOWGY9qaD
Cl5CD96UL/2BCdzw9NjfwIJUDjksb3QbNt8Rw5z1nu5aJkXr9QdSH0B7J+o5KfHSo/xKXIHWDpI5
T80oOYfv/lbLuF/nfSoxptBqkc5ZF11zxHVV09O6do4Q65j6zCr8dBj1ewkhJpq39mcKtDLiq7yc
w8j3w2jEishAeR5phakvTf/YRPWMIuxWBahI06iF4sBcCOISrcOjIC1eDX6zi6Q8LFFZ9cCnO+L8
4OuClEDxtF0k1kvdZ6na0U8wHqszSasHuKmDUWSwx0sFaO7MAcd/l+b2DItZulrU8YbLXNug0TFr
UL3C4vG9F+fsIGZTv1kPaDIIv+EjNzq2IGrD+HuY5VGFUx5KXKm1FZoEA2f/9dwVIzOKAcv8Ougg
Xn3DNN6rHugscNFKmcZ1mlRGAC0L7EF7OXtsX8LncGYZqRNJTypFqkAK4wE4HeeZcJucBJgUK3vZ
fkFWlLTwD0b2zZH/CM5Z3Id8hGgi7Tpqx46YIu17wkMbuOUV6f1Sr2XMOGxJTwytVxyNJwHn4hIy
eJmJsxem6YsBbhtHSWPXfvJyqRaqXw+aJqfl+WvLHdbzjYpsgkIjtva51oT7aS7DM3BFqfcmJ7UI
R+Na9dXRBmELO/MVtUxy7NEVsmwKkQHWhxBoGgwjPKZ1uXuWYMKdgvwwJy+nckIQkRH7ZEhk9zEc
otkM4n9T84k0j7L4YOR35LcwFZG7BkvaeCHVSKptV99GILyhADhNKQsj2iMlDLB0M+/WOzR0zZuB
ZeL4lDIMVWJfZoBk8ICQWDzdzbgfPwfCbv+GKUwc5hJfCmdGKf6LNn2ox5G8Utdipk6/yGaZpLY1
w1SXDx7j8H/kJz5O/PNJ/HVXx2tfuqwc1yg0+PkejZBbNVgFkZw7DmybLuGejS1lnHDJg1cLc/zR
bDZgxfO3+JRhaQLbwisSCfr+8qiSLNlL7hk68EoaTssGOLhTDPKlhtW8LpJMiQfqw8ZBxCK7qtnM
NKcntGRu7DxmyTxbPkz79mRdr0U25WQNCeLBKOCJW2IKByuIU1jEJ8QziI7s9UfB45vQznRiuKSI
B7hflx3FpsHjpsvudoSLIgjEK8KuwxEHnXqMrphIiD3CIK3rCcEHff6IxPnAkJAmO5NtviONcb7U
hbJebnAzJSU0IajQJXRMNo5kyhLKqXzYGlGizRlymyK816vPnKlgKTnOiMgKs+Cfsxm7ZxLNLiTo
/y6YuAkUtvH3m3LUjK+sqiOlUv0lR5ookhR7vQU+Gm9X8ZKNozNaETAia5Ml9CtuiY5DHbgNnPW0
ZxN5EUwyVuloQVtTXKhwD4EchUeNJ8cAU0jktUCBy/PR7p+T0uFsMdOQ/KQA11+JgQkAjaTsOa0H
Gd2xn1yd8SA0kX8749g7yaxr0+yxVYEgvq+Xy3ucSSMRvQmCMQf9nJMamjkQBZ11vS1B0PNnCWB6
54AofeKmV52/NS2m/czJUD2wrN8XxFAf4RrFECSPzo4H1pAxujveugWbaFOFMD/RnhHevWomLJTm
MErrtFjVzP7ZEXYb8pOUBi73wc3dhjtQi1hdLF227KQ0iIvswBGv56tbpaYHKyxgm9fSDVbZkKW7
S4x4mAfM8WqSZw+fNCzpH7Is6EnOeocQTfHm0700YBkayqUEfM3a+3jjfHaeeJWiVaRZ0rj8Be0R
UzSSKuVpkeOqq80eyP3b1/x8CKTt/YcHJaFxiTKTfprkw3cdG95GIR2ev6M3ihzhb8rSvgdaYdQk
w1nKSw6JhVENs5xkXz8BdiMLuHMI7E1KFRlumQj2x5S06a+4fKuG8bkUnwe8lIpabSO0+3fBQ/1c
AjQO3b9GZ9LrNK3PFpxKMjFYu1K0SwUs7i/Ks+Lp+jCsg9phCw0h9KjKv9tSGrfp8E7RiSAcXak+
9UKkltQXffUI0UnTf3wQCRAlKxmp6Ef9Z3IqH+ywu5V8faiZnrDAK4FRbFX82Uz7rBUeAnSOV2dN
qYodiBW99WyLSRHrKm26a21UdByEVnokCy1fAezGbPhS1ubvg0xxjhgRFbQBviISAC88vE3inApO
9fbStVE/tGTHdmhGtn9gjdoQF0GnkWi4Bq0IBRuMHOK85blAlDo74gTkkeBOXLlBFCqBaCZNHudt
/UBzfmL2MMaHtKNfNpsWOSO6J6Gg3jCAKqeKTHv/QRZqBszR3rFUimog3U6ze4om+PFZdeYtpehe
ANP2m7N33qw3NdOkbC/kYpv4TZma2hDGqqSon8kmvDGbXe9c23KQbF8V0SOLViIXoFR9mBsuh04F
bjak9OxKCR3VJ/cq8yYV7KgcRBN3VlpABK2qUlLIikLwyx8LeuaZRXj+Et/95l1GfgAs0vFnP3kQ
DsLUteL/Gt4MLW3LdVcaN2vZd4nDiP8WfSMqbJswgGckoXXWCchxKcjhtelSxPCdlJS1EBC/JpDx
buPJ6AFhbms/upIp5XDJkio//atXH6mwlIuaXdJ0yYiBgLjVOY1dyQQYJQdctI27zziI8MiD/Cj2
t/3ioX02RdmOmq9WgjtdNxu7LSphJVlri6FVuypWpaDqT95Y2TA3MAtJseswCmeENa3Vu8ndekkA
3hGAOUfU9YdYnmmg56Qtc2jM2ktvVHQzpW1RoyZl9Kc9CRcklZV3ctQLxAVLDKFQchf96PTiRNi4
RuM0Y9tRFbGS47/KfNUJzmCriCiAlMAaQsLv1F5cdf8Sl2vm2bMJnQ/riOZYirEanPvBpw2R/xS3
yXa9ldc3agP4ty9JUtHvZkBujMw6PH0DXvUwE6DVcSfDXL91aebqhp9sTpv6Jjl0jU2fSr9FwuvS
gs0lkVgogSnl+aWkERibUdqzC6ERDwKxtzMXsBSVjYU4/rg/FRWufKVv552AJszNCpAuVz4hKA1t
Y84iQ4+uXqYwC+L++BKCUKF1SEq5XmSE2qYRvS1kAcbzyELBHB/7Xq0MwKiec70V9c5J2GUS851R
7YYKYOvuIeMhZZdg4WVN8j2LwnK2f/EslQxGh/V7ua303A7lJxB3rdQmrr3BGko5XTAMad/iWihs
yAogx845/ZJUxBYpq0n6DtJZIusPCOMXK/zz7kPEr96UZhYEe/65UNxd62/1Z9/t7xkKNyvAVsfK
MSs3YyjMaH8rWx5C8trQ9fK4hz2UNU9tnV7/J+R3WJzxcz8r/FmVxlslHghfjXio9rnv7I7UuZEV
Un2A0GPppgohsQilrAUMjsW6NEFtYpi8qS1Guif8wvdzXV9VLmdbBIDRsWT8lsCfJIfUkI0iGr1p
I/ZXE9j0olP8UjKjucM5Ndbg5TCsjdkfeLjg76GSN7mWUSCnjRoKTyw8toiO1n594JULMxRuzczA
daSvTdAo3hhS6ZHPZwFuzEv8wN1wm+6C0LElLQwaMtDvOUrNJ9fq4iG6OYleaxawKULyu9k+wZKO
C/Xw5BINR1nSgBhiOX5qGchRfKOejupg6xFnSrJgfztPBHtMbKN/coNiCOpupOPn8ilLx1qFd7QT
n//Saxn4s0FZc64FWGMIazE1k2omGEQqDFa7cC1AC2iwFRqvU7PBrfYxGnpSULpLtCU9qzP8mjWm
ZeCEt/MxdypknZR/+PEgDDg6IOHYaOJU6YTjuQlIJKqaYQbmvNk9m7AbQ6AvJhNpOCjXgdCXnldr
JHHipEJkW71As1aTyj8aEkI1RxM86S0nBqWeY59OaPevrUrXF5atpFW4vw33JtR5pTCupYSG/4HG
CFF+HqY1isMW3sAqcTuG0AXy+4RaD/TfYDoF72mXYIMq4rEGi0CbMtqzRI+lI21K7Bx+rrau5fb3
NUabg6RW4AvrSfUBAylmaeRvI1Hx+bBoeE2o3NKxdnjUn+81eBcYDoVkxq2gZaa6h461AXlybg8i
5ekODQaPmlHqxvJ1wLbjWeg8ybQKIBbXTZJ+IoJw9hYDQCEtl852OhLsh/H0pgzZ3bYxOdBq3PUV
3DFUTtaBR0KwRXXsgakXfpNsG7Zz0JmDnYEQSfeyjUR1bePa3j/8uqdMBVTu0EF6NPhOksDHWc4T
7M+jFyvJMl3GLGCeSK0VIISxZOgL3oOn5HsUg8CgwAbcDcbP2CASUbHoHAECsedyMzO5DbbjzqTK
Juf50iIQFBpOU7UqXdYzF2WIej2R78aLM7H7U75arc+OwxsOskClbRYR4PJDSzBwYuKlq0j+ZKV/
BbFIjwc4+tfI5QELucNOFPbI8rec4L4ZOGpxXrOG15GIKq0CGgSXE8rYXkyC4FiQee2ZwbJ0VoB0
ZgL+XaDqQjDsizLNDk35h8pQe1Q0+EwKR+b79u/GEfctgO1N8d5xEWmJLP/3CpsxhGsCvofGVI/P
BlFus3dHz7F1QN+a4iS0XMbYbii+LZvG03QYp/NGh/klkjVAZi5biAfTgQxO642iMP3jJ2Ktu1BX
ajgQD/1lKKPsrTt7gjopOxtXE4Uozs9VkbdecD924b45pqfqzGchrCmzB4tYyKQ3tDuUVLtO/nQH
rsfa5Pf+qmDBjmPayi362ymLZ/njL2/xmvJFP3JFAkwDi7/RjWkFZN6rWe2hIi5VxBdDH9qFCTRw
MFNyugjtr0HL3ee1typvq4NEOjoZ0bqrrTIVrJCqo0AkWoOSV1/z4Xv+isPDFVOpOKqmysu/i08J
xblcm+tZxhwWgCMhnU66GCtt3fM2dqb3IhyVNHRCDHq8d4gm3GMjYRyupJMejK97j7wgsJ4Fuvwl
SZVUEUOsS0CDX+D6l9PH15Mu7rjTiBWQs6/R21bggvKdQ5HOR/O/OEDNwSxXTDngKw1NfG+rdmsz
oOL4LhJFFXYPJFQiFBeYY8HvqatQvA8meAkHHvDFjXADD3FoN+m7qn4RfbQr25dEzbSewYVoi4hr
w5oBs6VYIxsVDcljW/Jn3uDtzSKJJ/KhcsufVCdKXr4ut3N7iOteqV74GNOd2t+NjBZMVZNRtVUs
enhGO/t/JJaiJ1JZoS3WbJKqd3PjDBNpg8rkErHmsqcUhvfmiFNmnA3d9kUKXzosT4vrrSLfF3an
FVfszbvLWNkScrJM09Cd/FAeohltlgPtvbM0e4YapuJ8vKGWedTWDuU6mlVMCwmxeoqRUW2jqt/s
hKr0PchBmqWxZmWaCholBPJkxFhMVbabng+b+Xau0MEElXvzVOq2rUp797bxVpqr76wNeJd6lV4j
LupSdwXUieT/EiBliOgWJFB3qNon/kz8E/tdi2s5SiCa14fN0SuGeOiTfMZyD5J32QSHPWXmf/xy
YFvaT2BjqUpIZyzXKGMVVXZNA5BKPvaph/2FXHOPmXRQ2gI5rHjnREx/KDMQVM0ffa++r7pnkBw+
s1iCuvfuXb/3T9WhBIvKqMJScxqicq79w0ZBTiS/Td1i/A573DAqn1bfKCpZB6GfnfwnheTLZa0K
M/9F8dod98L6cIift6GofBlD2mk5p+GkDJMD2vGf7mITE2X2udxmAkpZE4N0Rc/NB5mPwkBeUWup
jPJi80U3lGivyGzoj5vWs55JXIri6pLHqWQtDnuRMcOwgF0jklZViy2i7meMcJNLLV4DurzK1tKD
r3r/kZvglspu794s+U/c9iu++YLG81OVrVswDGMX9U5SWWe5EJQMoUSuonZElHjxwGHNPaIiiSgw
jnn2H5ON9eVSzjIpHUpDYfrWl2YSN5SwwCZwfQJXTXToK4Axy8Z/rwNERuCuVLpHx9oBJANYSXIv
RvY5McoG9UnQEFrrMKA4H0HuWEN89SEs177/cDfIMUUkqX89cykIxbfCzhIBe4jzZ1mCnMjIQ5Fs
h8FXYthx1P9Vh2ozMSFW+Xvpfov8nSL2c+DW6xmz3mQHNqea/g6RjM1c1b7LyRE8S2T3o32A+WBU
OjE8xtg8XntCQ2JPOMcd2/HokllxEr7SzYUlbkWm+T6LNh3huq/EIp/iQZSm/ScNMCwzIbJEGhFn
HBtO69ruHUp9TYTATvBoPpLL/q99kiimQFvZAnltoKoqd3OucMksjg+GapEoOuoDAxe1YCjEE+Vk
lPqqYz/T5OM7+hLBb7GGqSRSG/k47ySfP6XeKQxCI4aMt6vV4OyvTC2+HBDAQjwWibqUQneL/6Dm
Yrefnu83SqkKtAn9SShVYZfHTS+IejFmkD2cjlDZkxbtMQKwrDSUt8/Fxwx+76IxBROZml+GOQRq
dIczuhSeiWJBy2Yk3YEd1TbI9OvzbO0MVJ45O2qWFWeIOQm14RQvt25mHlbMg1RES1HE9JxtIlcl
ty66I5Yp65A6kqrMxql9sORyOONErL1w9xO9v3waSoiWnNulcRxNCpv6pQPqLjyyNOSY4bhT30+D
EQfFJGArr3hf5gOmrGXRI11vM/qZwRcW1carfYR8nunlEPVYF8nOZG1lZLrQVoXTdXWBCGu8gG9u
rFOaeC8LRDk8ERadRgASnVop+S5XcgLctJsu2SRdSfF6uV1eifOutTnVih/+5qXlrhWlv03NX9go
l3R1c765YATwPfUWIL8y2dFKxO0sXo5ZNso+sFg+34KvvhpUa0kp3HsoZY5lGur9NAznNobvqWfq
f65Cj0htwMlSQ6IoWVAAtNTcWGlhsxw7gOBgHresbaiyNPFubO2kgLwm+0spRo/m+NZoXPxC7Ld2
r0QVxLfzI/mDIRHn8jPNyhVy7QfkY3NNWpPYKs3j3Hfnv3+si9QDcscmvqH4lqHawM1W4c54+QJ8
V0VkxjV476Xx0MaE8v6qcqnZEbjHRN3+tSiIQjcZ/KKX/SQhG57RUoxscb2hOJwf+dQi6E63CNzC
Jn+8vsR7GIJjXEcg2rKk2I4EKm3kV41Z620yNF0AGh8lhY17dgsdg+ao7GCVuVJJcjTG9vCXjWLM
BGtLix8yOazbBAIZPGP3vbHjdbaC2bgObDhqdA4P5PRIofJ67kxN7g6uEVxJGQM643BuG4/vVxr5
+Fy8j84Yhu4E+CiQPTH3qAP+HmMZypIXR2/ZeIBggBon1A2TmWd+KynBtRl1K5W0k7z6vVQjOEzg
O8f7LEs0nHRkaXRJr/RapociJn02gjt3UPHX+VwKG0rZ9uBPf/ig9MRS7sjSyS7PLYiZBcalphfa
ua5ugGOLShY+eN8w2++yt6TSOCGXMH6P5GmeSB0ulzrz6X5pFk2+lY6WokfQj+kbmdcGBbtUPHdk
pCyQ/k5bYJOo8fgEePjpM1P2+zC+P8gmpvQ09geHmiC05hyVc6JGF/6lXf24Tgb3LisWx9kY/JqK
6lwtNENQ4rCdKY4LWZPwTf7lBlMc6EAQuIHBRQ9r3Cb7A8IuXJfg5xaWp/9Hubm3Mxe3/Ocm1uSL
iKYoY5GcqXDbEDI0D/SqRFvV7Yj/VE/NBFcDdy2TLO2gVmGkXgk3qqVp8VWyKe3x2eupXHU7xJxU
MGyzxSCHqFVXTAGopnsuQl0Q7UbUFVq8TiPW0PyLto5lTDRzpsyCYmdgjiITlQVRbJxCJaPukKmh
QoY6blmRDhXE7K940H+9QuCZkTc5wr9J9VWtsxQ7/j76Bm16l2Qxdd6Pni38aUcI2oCqI6RPc4+s
26KGQiWYlvX4DN47fKD26NsNX8jlwUShFDtMHuFD3xW11DOh1Ztfl9TH8O+XLlidC1U3snwheCq3
pEEJeon35N9vTlD/UOqyNpNjzhRkAWcl16jNDxJxzgJx5fFD9yU6zG0ly72Oc3nAY3UzS2C5eW8V
sK2mPgi7OIfVSEI4Vxl5rOCCrmH2lOkjWzWPCjr96AoCccUpLMsDZJww/nqzlyE+0Yz3f6DfOa0c
wwxTI4EcDaWedsTApIv5hVGrY7h4z93Duwvm0bmdWCS0CyYl4jcyV93Tk5PD6Og/prXYCJ2Uec7K
yuf4xdAD1onEzryMxV0CGaE7sUwUg/5NDn4GovKeVdM0nvbmx8QLhkRfRC0vbuO2Kxz0EGTbrAuf
D5/xPBNExcsKEfkw0LVwg1Dxw0+R3yq6UsCJbRUlRR7SoATvfyROcV+gcJlmyM0n9HDWzTrnAyDM
ANJNWrpRbE8CDfvU1m4wq6iiUgxDJVjtQpaaWYlDOZDllvBFSxTa0paD3NeVmy4mxPz9+fboIOoC
gO3FGkX7nrUd8MDk0EG034vmFJhWKSmZasp7jF1SkT3ROITw2yxmdYSCndRBbkd2VrQNy4USacZq
8/xlp2b6l3HGI5ULD0faCIUBp62IUGZ01eLjMaPvPysmbH6iSGvyOsdL7PBd4mJ55wRX/WF/e80O
tV7Q1gv1K0NGvbW//u8vfInysFsJ9hxHzbJcQ3ehwMY0tV3Rr8TpP6EnzSNLywno0PmkM2AfNdop
7NAUBFU0tBS/Q4334JhIn8BMFU1aPetylBDhIH9lGjs40QxEtg1UUA3moQAYmsSn4ntkCD04uOVC
8Ge3AZ1W+zwZ2N1QVjuApzf6GW6o6i9XTDqRzqMmz//9iWjxG5chpgTKOzBezONtpH87yr58gOBb
GmKr4qCW/1arylrui0G/kfBsxfzx6f1K4yEfuwxq96mwbaulL/pdH9HHvh700uMfHK2Hc6ITEXE8
HjFBordRhz2ugv9rTQCAIvQseogyqACfQ7Dh1QHhhxCS8X1p7quZGhsFt7rcbLWE+fUzqO46vEGV
KlyYdeAAGFhtilfVevKL7wok4I8S6DtjLoV0tOpXuN4vWUL21SkE4IbYwz/M9yD+dGsObD4ufKal
9yubgygraZNLvshVVM5AxmCE/A5vrncGZDCGtD72NkIxTnGtM5CFIt2KG1nAYHBUl4QmP9MxDmwr
DUZGzuAwrEh+82HMTAogfcCcdiE+1pcq9aPQhzqdBP05sS076q8fDv3yQkvWYqR+L1FoIE6oHBAT
K8vpKIxHyXeEKjr1//BA/5hRqoKtbOo+NwOhSVnGWgjl4DUbEnZs3GrpsbO102SHEI4liFz8uBKU
Qj7WeQ8RolxM/UrkvIvFNmbbiYxQqMgh/z4rPHtfQw9PkCOMOxmIWXGjW7cobIWGkl5KzQM8EOXr
eGKmovv8Zrxxg32JB2pm5Ay5rklghAesQDWRH1TbmMbfgcStQa5bk2dwQj1lfNFSqrCp8iLQvfUC
d7sq1H4gk8thaSfjBX2Wdb+AKDCcXE+ZkY7hcZ0/kRcyRhPsqwEwLYbpf2ruV/v7ODRT5zNfhCOP
L4Tqa4F3yl2CBeHia3ZCzyEKOsIts1r8RmpyRSZd4aBOwWdTOff2h94bjwPZIjuGZqVMCFZlTUJ3
wqVOx/ft6mFL2TvrI+e5Ui1yeSvrWp9p+4ZA/T7x0GP+vIQCki2zhyx4GhqKc53ueGTMEWNhLMac
1ru8qbWnznEtjEezgf5XsH6aOzdBP1PrxjS3XkBXjYbkIrQ/j60gWqM+2t/3roA5zvP7zYEj7GHk
YfJWrg95GmeCV+Z1byx4ka988+JhgTfJizCxwFYbFjbFTgHjaYoVwcneDebZZTqIy5KTlOjOeoUA
4owANbUU0+8Z0xB6PHa9efrYGfv6RgClhbYFHI6lpuXV5BvRvbVdo5nNlAFqrT/Y8LEY6K/0PxfM
6WWiVxsYV5DJLt3aYtoZyIz9oQO6wBDlKKsNkgbmaZx2ntjkclqIwNkdDoJ1BZ5bL14v5PO7vyrr
IDS0yYzh4ewwBVnG2ZwgZi5JvKRGKGBZNtPwYcYuE9DuJsxA09wsGgYVe2qekklSQSNBT0hSy6bC
qvcCtxCtIZvVGis9sJRgrBJ3siSfm6TFYZ0i9h9IeI4vH9H75N/bW0tvotyvsNkTRgYqkSsF1IvK
ZdxpslodwqoqWMwQttZy4HLg9Bxa3cTkEsMNucbIeUrd7ESaIEqRmgimrS7YtvIGeE7N8sePUOOf
7it5KOey5TAmZCJ7czkgZLHXz64Js0tkwO5xdnZC7jySQ8CIn+nB1mEMx1nfhPiMN04gyYWnhoBv
iZxzS54BBga379W6VIJD0n8jp9P8sRWDZG8rkmQjLU91zf6cCMvEIvJTvAJby9Eb3cgEtTxhtOS4
r4qBwG+QN43Is9tV8t9CfG0Qoz6dNUvI83L7L7R4xadH4wS8SpEgCgIc+BAndG8UZ+MGZVHW08rE
RSXkcQ5Wa9XtNv1+8LgO8+yJFAD+dgdyj6uaOFEkieMjQwe02ssb4HtE8yJ3OLZXeKYyX5Te1xIF
yOk7ENnNMoNe6kRAFnFWGfkTMG5j5OvjRfQOPQPu7Gzu5ocNQtdbOVL5AXIFvxNtViG3LfZ2VbsD
b/WucBfAM+LqXpq4lHDmmbqPbcHaItL2xtoZgNJFcUh9Cm9PU5q8hEgzM5HKdL5ytdQ805kvoAbW
XCI13A8HEkZ/oReJsiq4UWC85Zcfwmrna7QafYw6MA2ezPwok68Uslwt3qLq9BtzxXki38qyYLbF
VfhrXE+nU21x1DGjPXhAqMa1WSgTiLk6caSTuSWvc808g5v3AX1w/Dck/g9W5A0B/zplaPZfAaHS
ZmkA839x7ap5CtGtadzym5FvplPoCstAS/zbz8Wqfk4S391+b1pjRfqQK7TU6ePuZtXAShXZibul
0Bpx6p0ZMacOhKKBrmv7r17JBFem7UBJnaTiflpJaO49Z2tAtWEhemb1SS3lOLhwUZ/gf2jH5+Q6
KiomUV+k1PtHrZuTFhHb447PpRcIg1wFxk+oIWIgIO/khCXuSHJiMGVi4gAR+Gzzw4O57dkzSwJX
UwPE7yRUIBatALzZ8nnJmG2VnE/GuTITSIPZZ9dPg88sUjJMF2ACtl6AdSDEotvohKP9RmLtyh0Y
dU91uc4H8MtuXdZHH3eLEcKAjbaHc7ABasF6S5AGipL7b+DZ0GsKSM/xUSdDsZ4u6BNEMrbVjApY
sV0AMgUgiRbT6ZEoxKRP8MfYLiW48885KiieIY1+yrnZZoP/mVcxkePpktTpN3grwOUwOB7SdGPI
NSuid5rUw3dhSMELFikt0JF4YhAezO5xy3OGRqAh/TGyiG4PQ2N7GA1qIFSxVJ6NofaBhuo2OF5V
WPfnDQV5LYeo63n0lZa4/Z/HDMylNneNDAeoCSqDdmWi8oTHJ4SL8lCtt+ALpZLRuTiIDg1hDX7g
0jJP4Z4A2c0xhBzDL1Sc0Jl0sPWoGwkOxBvTfv/YWExo5B3r9Z/JeMz2SS2IZpB37N9SWvWkMaqj
BPCRdqZHoKYw4i6VI2RnAhyPMNaiyhhx4E4LbjFIBgdIXjcq0YnOzjFXkgpY/wcsKjpGgcZ1Zsdx
IkpyctvOZbLFBK9xAr50/z8xBnbccSckRdHSzP5sW5ImxGCqwmV6QbGFQeora/Ac7CeVAqDAZV0k
rUhIgJq4/NOZOftbrNud55btVyCPrRZ7pd85T6Kh7rOIeVw5IXE+Ybshm2L3lkJfiAkyWgKDx+Yh
CEqKDE1I3YgHs99RWYabCV3Wb8MVenZ2vaR/ChZJy3SDdvaQMsKFvnIJjxIoENuIyH/pfM9EQWf2
J2AEzbYHyHQ6vJFJ5PWwRn1XmOvc9IO/qObvG7S/vGyc3Si7i4hMAglV0AlT9SSuDYxVqhHpug/x
tGU5aarjpZO9JXO3uvamO2xtTcwvo2JUQAd5bcdkEyIMqxsL8vpbOharBmQSqxORG5FtIcLOaziq
zmepVv6nM+7Q3aL0eqqSsV1Bc2ZYNmqaFxYOtLg62I8vGNs/bDBtCK5fGprMjbmOJwUk3HHW9Qvk
V7QCpAMKNi8UsdE2o79Dm8uFiAMMTaeirfe7o/K+JnCK7S1uuDSr5D+aIB7Dfh90FIqXwJ7gAEyI
GtJMb3EsNl+yVZtu3ABDYsFR2fYfPhK4pQdw3aZ+NHAaC/3dNMicP9sHjO1H8QNy51GF0j20WgZt
STvpOG73uoGp9GrEsMyt95FT6Wje+u+kBHwKUacmghDhrfpY4fogRcJu98ra/jm0ZBT49H5nDJOe
cI+5bQkVAvDuaIYJLUbvz4/TNgL2qApLebdavp0HAlRDCYW3Shu1nZUBd4juBfmqShpmgCh1thCP
Mn8BgfP9EgDGcbhQc4jqFAfFx+po4ByWpWQalyika6rdD2gk8MNZVlXAqCgDwD6fUf0O4yaGciYk
8NWixo6YMiCUiy3w1i/7mTcG9Gefkn8J5lafQZtWGuQZs8UDmXnavHL1m7aYee5UheqTrNOCGDft
3lKwxxKyrZRDYB+BpG1O8x0qhCiHt1BVab6WrsUV2kSlWy04lDXXGodL57FIahcYu43lBdGuneV4
rUqWgvWPqpQ3GewrwnGalyk/abuLqXG94JC4PYAClq5N+wt/YnpjLQPieAMS+tygy7Y5wPxPBraN
Cq8d/papGpiFD3wfW31p5IoYUsOsZ7nBHsmIf4bsNUwt0YaPGn0A7ndHQBVl378kEFUgvdB4jRTN
SNs0+LrP7Qoh9IePxUW9WWQPbczFiz2/BRhs37AfhVv5mvr6mzAA9CKknNCS3TbLuEN8MrC1qWoF
LNGzUdYGPnGYuvZfapbgLi4axQHDLCkmI7dsNbtKQrL8ARzS4rG4rGS2P/G/rSOfMi15SN1sgQxK
Ytir4mYhDgb8ivISa9DBgsI1K5g7vHkfTny345+oSSrE7GjIPHquhGdmy2AQFNxfxV+2xeDkooQn
imZWqZ6u5A4Ad1ku/+qzGiameir/H6fewG9oq5RAitxgLiIAg6e6HBuOBccgmtXVULYzQahSmS1c
sfr9iF40vgvWaK5O57AwzAmK9bHlju3o+ZI4vulesHOc9dHwIRXyWcr3gVn1eLwe2YaBh8cWPXks
Cm9+WIMpP/oLdIJfON8hxeUlKsh4frsbjlE98SKP817NOP68KIZkBBTybTusP4rWklw/qt/OA7Jo
bL5KFGaDn6kpjMVae4lpeynJ1PaPM3BIrOvKh1lSwhMqv1golhYz4D2bNUFndOVzkPVmxVvV3uCn
FZdrg38i8NWh91UXUZag3BYEC4/FNhX56XG9AK5xNFSOI265n/EqzmBpknK2fo21GdhoAej89KCn
y7fVfo/euNCnhvUX+PhtAqfcP2UhYx3UtcnE/yb3wLshNMEPDhP66Xl23O7mR+Mr9xnxdx0U7smC
XEOV+99RnFxIIwDcnCL24NmLNcn76MAbEGbuNaLacKdekqV70fT8TYYL6MDVFAsRluW+TgsII+cJ
gGRHADI1BGVo96oL5TUjIlr9dIKICZ46oo/PdLuIM5quvuKJclJZkpKYgMdpTxOMXOdiGq0JPXn+
a+/KDMyCgxh+CZ2lxgLI/uUu2lIxdzHiLQu2ZzHWmiCPt3Iixfh9iGsY6/eYYh+w0rr7asc9hf8H
CWMWOpYqzpFnqgv2m8AMbkuOMA0jNIekCjnaGwNI4YHndbvmMAAb8KsxyFif6wXOiMfpRE+eMXq9
Kx22SQMiOpIdM2GIK2Rv/YeHTd8+2ktONgwgCQJr8sQePuNNTFYcKTTQXJlo0NbaSH1VUwMulEOj
rTHZJvCNno84siOMqELLZNd2za9cMybaYlX62y1k8eRYZZkvwQa38Jwv+GvQs2BigNqQOU6H6spX
yWIBb0cLMuNzfWvKmuG2exz+PATbwcjzKK/Pq9S2Bkhi5ZAYUplO7ouShrubLOPQO4xTnEiNiJLe
mok0cq0uHe+qhl+5JxpKCqxaYQ6TRyMs6NgXiLoWMP2EWTBalGMGmQQtRTvOZRsK12vU7bJoWBwM
I/j/Vv/TZCpaDORUi8CUGZFbtvpk1LeYNny3Rqm2/5vXoqIjcRRHiPxwYN69Lk2Pml6V2OVC6MaB
TEK/Q5RZ+d5ONAmor7ye/othRSFuZGbuJrbNxwvHsRtKOG6PQOBFpCWC7kafKoZdWxAuNMm7d5nU
YK89gaHBuFvGp3piGKGWLMnlF7941Usn7bgw8x5Zl+IWTS9S9RLr/P8EC1OaLmKvtwRCjYMQwGuG
o9SR4l+W4l2hKxnGnFcjsxaKEIkcy6qVbtRCVQOgIbX6t7c3TAEWz36v/67a6TmuuznnKFHY+rxO
YhdnPxYMIlaja1rw79AqdTOAzDX7nP50Gx9bzR4XY19P4zVipGJYz/cfbEpW4X0GpT3yOfxVpah3
zt+5SoNWnLFy3K38kWNZnVzc9nM3JJsLEXpojs8qTPXc6eAGrgLn4v0S5GKJzRrOb7S51LsXl//1
m+ehz6H96ribduF6lg4g/2ElehpKBNQGF/246kkMKaW0Lv4FWwzKHf+fkUXPNxRtWr3rTu4NA6Os
jWkQnmplTOE8AOIZxlpqEtDv8g4H5lKVFflocRfWTW9l9/cfbm+rKeg9yIa3aMO0Ezk+h3ua+Ay+
Tl1M/GS3UH9Ccytj7E+Un1hl8+WHxd4Hxi3j5nNNVbS0G1WkJvqK0qwIpsrqfJGd76rFr5LvQKBu
6A7XsPnZCo9WK6FqccYX6ay/t5WOHP+WVMjtR8H8mYyi+PSbsjLnPrqJiWe3YgXkRGXupq2z5f9R
Zw/jMeEe4TQdKps+ES5/aUlpfJVtDuzzRUeeB8bH/SZ4OMbKCzsRAf/VubScpDAhI63QYHQmuXlF
ECIRdnqMrUqDY+5rgJW0hPLbM7TdXAwRUm7fyIE9zl7vqfXg+MRetmu+UZGNJUSbRFGVY4Td2Rpx
YMv0CHL0HGo3vX00GP77NwUl2sNF8ANs0t0RM//CcSEUihoqh9811NET6LdHE8G6NiK13AvMSAxW
M9Da8g5e1rdqymbM8BmaLWVaTH9TzU+ol4Fj/59dfNcjFsYIki5/BOWU0c21FYnh8mYXWFEvumfQ
GUV9+VK5WA8Dmqg7qe8Bw5ZYkHMDd0yghs5p7e68LcZ/Q/AX1P9SmytuPi9D4++T1utv1PaEvhGb
ugTlG9diyOdSjoLsuehPYbwnLlsqobtwZuwTmwZDPsPiAvlh93KbirEJhncC2ddPEPKuiKuE9/de
cNahB4MsbPKwLkYCCjR22iIKHA+0BmtpC2lYvnX/VhCuVVtT/GSNozxeVrskNsvpuFf/SPVFjJ/c
w3dQrmGeVuNE9WmGUPYWstKgFXPVCbdhseAF/HHPvD3uC+rApCBC/+wsobA2Xi/cJs7Cjme5ECAK
gTDH/tyQgUW+1OZRS99Zd2axdtkoDmBvpPvDCxLU/iwejDQ7tqZs3SdHlxWhOYjImzI8cvF09zK9
kTlLacardaH6p1yWCHJFsh3e2oSHmqVIWCYRIGLHXBcdz9oHzjKgbdIdw0xOismiHBfu5vLJr4e4
9xu5cgXrf0gDlaHDxLhLSpgs394P585fkVp4DLYnEqCWV+thqo6+cGjpiJlANx/x1AoMm9l4rzEM
7If64bjHW2sdsYxRKR7fsG9AUqziXZSbu+M0ZNUj5mnBxMXogas0j+VUtoUDAuzronqx/Zp2dCor
nFxL25PKZEPDKoPfhnmiqfCfOfF6JMFi34Ab7J3lNUoxr01KJuTu3SPOpbg6HwNknQnYrg+hYSSc
qci/EhpUnAWmRn2seqTrFqH301lo1ixtc4kJQK1/1YCd2G12ZuwAzpMJa6pAQ8FxW1OTZ/yjU/JA
6cU2BEn0h6qvpw4S7MOAgu6gk5iehxE19dGQM69WzfBAjiQ9l5LLBYXnKiy0QOROXe/2HSPlwQ7b
OKvd8oCATVJGoHGpTMbzerkhgXbvz7W3XiT7xMpSz4Fy6MeY3Bf/UgJjAnINFh7NhFEqTie2j7XX
NZAJF6T8bDpNTRJVYiON++Y8rK81wnViVVG2nDAhmUYoOg40ICyMwcotWUNY1Vb6bCXHmg82aUFO
3qsG2QKSLWX6Q5lOs0ncFPxRzS6OIGls4piZcpyXaz7VzLm1kjZG259p8Nqxlh+PaeEiSxazmvMC
tiKGlcHXcHOerZj9uIgaac9greOGPuWkYHV331Bo5vw7nq9ZBGM6A5kMsFFggKcDyZdDy+vdE2KE
aV/8ye0xnRCT0Ys/+Qd1a0aKOT0pybej+YbJlJ9YPYTf6i+7cRArn3B2sQvv9kH+dXGV8y8lNjE0
dHeTjHX57oOvsvp7E+WNYIonZK92sMmMMc/y2I7YoN6pCuxj69kBZJGV4sPViALsHKkw2VjXqgGZ
7xCcuxjTbUG//s/it8x6gjFtUUeuEY3DJgk5FG2Xs6lgSYsSM0DnRyVpHpEtfnnv7cfd1Rng9C5K
ZsISsk4IPIeMTK8VtITk1AH65PhR2psjO0qc3/QhscEHSO0L/WQJDH5Nj3B2wRtQMopHvqBNmr4K
Q7E+VQS+yIMa+7JEQcJg9Bh1eQAc2LzxXArJ1m+ThAHUnMkPr6GQ9E1G7TjYBYEGh4wSck6IBfNQ
LjQBt+wQ9PeIV4/8n1Up9hfQraQpdjrsHcrobZmY0kS5AG+W8DOw92pvWwtX592/J0LaVzxqVUpV
ArxKXeH3FV0jJfaA+JzoqzqrzDauPCm3mcKToOnVhBWoEQ/Oj3raWrte4f2owUctkGdZoAY4U2pw
I2MvRDaPb0WQ6+lFTi1gSM7P90U5unZBc/TT6CuY3/gKx4FGrG7sOoh5wuyhZai7zSYOILkZ1sTC
eM0ITHVgh/Q9RdmtjNvFqxCxZJ2HZu/EvzI9AFhZoryh6pAKxJ1rUxRklaSWbDyKVCzEAVwzirw2
6US9cnlCEc+d9y2YlkVX+jMnH1AB3dF9tNeioOgRa252Qznc1+nt8Anh5ddoNF28KQhXPSO8Pv1D
tOCZi1kM7JdWVvOtL0hgMnnF5l5n+IZ7uYOBDH/fSdHOjHRfaue5+P/7ozbeRK9aEeEvPUtjrMFF
kkECj4EAnppP7qrpXRXcfG+xJPZIF8YpNk9SqcKFZ+G8fjABNFrifmjQkaDCb1EPkt4zI1WLX2wy
vxNRdftIC2pMrrS4Acukj5H5s7J2bYQ5hzi2K1stlpoRL9kKWVqCEn3VST3yZ6pEiepVOGAnj+39
kt0pQv1TJqlyk3siIYg+lKcpr3WGJmm83Tm67z+IGnEdM5Hky8YsAyWhtLsiZLfueTnQwC2jjIlu
lZcbh+u+zSENXKjJXpVhVjxEfAx2xoXK3bZ6n93sXTDQP4o+p8rUubwkZjB+OyIQOx8kLl9f53Mx
hm+65QMYQYLvzchX8cTmTuHaFm4qKJSJOsq2c9qpK3zL9V7k8JUTEtIw8UohQfWW5kDYqMBvZgOg
vbCFiq4aCQzK8EVqPN3heO5DY+acOtYrk+ZIoBJlzEy5Ds+UT4CvxanRpix/RwFAg51OI4nwOuGC
2Fs7TOFoGClzd8/nVN5wsRDrLSzK8RhelgdqYsQQ2/ipiLFJ1PvMcje/v1OmVSnwYDin/Pp3lDZ4
g9qcsdOeCH4LFhTDm1P96mde2sSQwQn5vyRRh7loJOuUU/nPLa/7QmMm7mP1aBYAU7gWW7PUwqWu
h2z9M2uqAJZVdtFo021q5bE76inhflzyOad31H4WzaPWcDgj2XdAEAO4plcg8gVVFVX+04SjY3Bo
nuCYdy41BTQtT4p+zThTsj+8C1bUhabu9Y+XCZ9smEX0dfb6jqgZWxr0RWP2w2XWIVvc0fONIWLF
JZcPHjM7PIwqiQzlDGyEqSzPY+QM0JozTjmHGyffrPsAfI1wvLzXMWd+mkxjXaop+3xpjVhDxoNh
DKyx2Oxl7UJuNs5K+A3qydsjbDouJEcHBgh7Od3uE1USZL8Y8zjqchT1VkY4FmfoFyMCmCIbUZ8p
i2djF0Iy8NOI5Jf7kdrYS1iX51C+QlEjvM0iDU3yufAxSOHCCT/35wKIXdXOlgqqyxfd7BikPotT
7UPuEx1NTi15IihRqVKQBs74JrIjNxggs6KmKZaxB1KW38B/tGzv/q9egZHWPZ8RrWqBISX4GI2L
mU5bQ+8KcH1A8KXZxRf6Pd1Oj9J5PwE71p5HaU3IO8r5nHFVURSlKkqxiKePFXaVRcoLv7wU7xki
vIyVnN4gVz/ZHvTT8Q6KdYNFO3z4UShd+q7GzeEr4r+Y6pwcot312BNKinHwTjkv6txnNW+jUo1E
GVzKrzH7mHRVQOqUQE62tFhkgNOgC023mVpbNBWQn70m5PFwwxvHt2yJiNsOa2S7tghrm3+EVEBP
zLNQqbcQ/LW80C1uC5ntE4CNx+mw4hk+h/d73YmutEqNZri/OTM2qz0bCF2XVEto0bNIex6PjQWz
YDivPberVkg7lRVGO3rnohVX3OEYr1tB/9t8GXvkJusogACP47THr4JlCouo3hurpgf3hOPeqm3x
xEckWYcSXMxQj4IbFxSMTu38a4n2I96VPA3JWyh3opXsew6vqEaXS7x78YwGf8Tuiv22ptVFgWRn
mx0hcJStIq+JKzlEeXVLJP+Ubz8ScvHngZz30lwZzlEdOlgQ0QybX0a8hIO0ZjKEekIVOOzwB1yH
pK+V35eJHP7mXIVTYtIZkIo4kCHrgZW0tYjhlozy3QJBzkJ4YlJbORRL/YUUM9o/1Ev9aZ7oDdBG
K4oA0VWdxazrF+LM102n8ThVPd3iDNKUapKbDAONobsTKJo6ZKPYho28xXPNupyl3LI/ajeDdLXE
f7Sybg4Qs2XVLDMwYuCFEuZxuENhYwpkRFYGMf1HYv+I0CCVEPOpYTrkZFkR2+PD4BFgzjR1Ft1O
01tSu27lsRK/ZvCaXa05V2XWgaomnWVQO500ZK5rJvrx6elumLP8aw5UFpbTUvqMd8wb+09FnIP1
HLrLf6gB7Ixe0aPE/sBJGbUh/lZstBKVuzkhojYCwEagCmIVKb+h5FRSqtu/VPQtjb0okJh2Tsva
P3hIGd0yhc0CYHlM06OkWRpeS8w51M/Z7sZEXbbIj/X2ST1lKZvLge8gQXzh0UdmeXL3Lr2ffPrP
sCh5jrL09/o86x994YA8FVgS1tPuVCdVlNgCFNCRZV0mh2Y/5lM7V7iVsrTJRzlHaXGLBAhlvaMO
9euUsKrhsnPyT/4PlEIz4bh0Xb1Z81yt5UA1ykJdUJgkt6GG3add/Fq3CrqxtbTLxfZrnxMOJaOZ
bjm2+LM3IxFHfMQt/8VI/rRkn/sK1WCcXjzj2bpJoiS5DpBT9paW6L5obSl7obESPjLLOs9/3rYe
IuiwPS+krGFos3jIxeFcys6U4fwhyB0WP3Yq9rnIpM9WFx8rfoM7XvY/2LtWfQ6qjhuelbZG/5D+
7sFf5WmXq43tn+15dwE4h8JMwsNkf2X7k1QHtK91fmLpGl5fBSRPAN0VG3+zQpJ3FZRwdnDn5Yrp
LW7igiRYonk3RA/PavLhhEIl+90+ehH1mLQrxzA3FLa3xFmTLiPj0CkTNPjbD67lBccs6tZQ5tjI
3Kf8eTexTKfEQFm4oYL28ZbawSNlkeiU8YPrHIT+A1MmeUl2pJlixCAY+QUJ6cAPlJiW075y3jq8
TLyTX2guriAOWsrAZHj7X2ys+k4gkdO41zbaqapSqtkw3q0JeKw5LqCLsmi+79nMcZLPn8XBalBK
L8z7kAUs2f7xvB6T+zKML7IpsxasFlEMsNAAwkUk5PQ5e/dzNS8qXqJs7ayMi4rSvXM2dgAiOLJA
rBeqcemprweB8KgXuwrT4Anms6Cw1HMU9zoKecbhh6s5pfYp1b56J3sEzFT/8ao613nO/GaTCvob
JBezneZh8/EGwPTeN4hKCDkgCCRKw+t9TkLQiMZVkfDdGdKsDuGjUmRHvJNPC4c+FgtvlhRg9chg
XGKqTjgiNI3OF0EyWSP6MnLFvX2B4oe2uurkgl9fXIgXx3wsIplIqn2WO2llhWNrTNQ8+uUVf1k5
/3WD9dEVc1KIuXu3Hqt4bFGjrdj9CcR510F7x3+2pbIHnKzFfXvUjv7y08lA52RZalRjynr/DI32
7DIJlOxhC7561SNPKGcVu7SKS3g/dLwWHwBXXEYLvjumJ5y1SUYfvVet94Wk7oITfWoaeC7StC1x
aYIAQZIdRbYL1Tpydc/RjSuJuOm/1Q/+sEJENcOBte7VmmED8k9vBgH6iwo35L7gXyKXcm3ZWgk4
C0MlRGasmDvcrnRiHTt089XElLjECVkGUGZ/BKlNLbZYjKXtVYoRxzoKQxY1ti2NCz05Xl8dZ40r
gLaxu4Q/gGEEBmocNzSFpwPUpLFO8Tf8C4U9lB0OaLvGx6uWXm0D7lLUvbcwalSipRI+PbD8zgQm
/PCEEp37+FcmfykTHrZwP0sy38Vw/6ni5HDuy8DHFXzNos3lFv2RWRKim2lu7vMqwQFq6mOLiYjf
xqHcsbYaI/cUfncpNt8gjs5fn6zewUcKmjRsHzi117PNPaS9M8Do3qt0BxlDNHZJJ/eaBkhgpIHG
e6ARDZVfAOLYzkCzgs0vyCOqfF2xrzR9MZrVDko9uoZgmSWHXSvf5PiesGWsiud8HXhYSMQD/4wO
bneFJ1czz3DeptrqY09JRF2VhY1XBv/n1avJZSwBj1vAbDeCmGQNKEQqPodEQa+F/k39hQmEeOu/
bS+aG0IcltNnNyVVVAjMVBbpjxQxVdRYC+jr8WCOcKfBCDS0P8OM1WCbNcRrbYOhGqcDGlbx3qsJ
sj122FRqsEbgZdeTRKk7TVVLj4i8oqz1tVtgoscZW7DvRs3XKQu2R8PQenCpTnvGHymgDfiUj+He
GerQdgkSGFauOiPWgZ7e9rolRCPGNExj9MIO1r96hq5Y5JSrkslp2Do54iCuzIxBSd9ZVCo21k5Q
M4uXsRyWg7IC66gBm14ANsOZhbGhq+/GjHPyiaEoS1lgazBhjGWv4OORaLujwT6tMo1sFIibLlzY
l8JEGkS0T7VEtrCFKoB3XMbJj7cWZ/v+vXRyRbdRrSgvgoitQ1I58gEsVTai1uVELPBuKh+rDs6u
KG7BG5SADXoJABnUHqEmmH4/U/NmL14NQbyvmvAq3G0e37PnTdBPWoFXXTtdhpp2ybeHosJpJrYB
JLFyqtVoslyqY/p17QpvohGIfXo2/CiigQ/GRPmNYd5z+8p8vTv+9iX7solVmVCIYMzH1QI1/lL6
V3AJFa37i0exBUCu1CiIXGUkMXMR2+WFaPOrkCUT22WhN5n4FYIkXD+JAD3g698gx/LvqEfQHKpI
FCjQTZyYrT1AaUGE7g6dkK9aoAcpHafFoGX0sVaBItelOTO2JoUTX+FKTLNIsqHR58ZdGaX03iVw
rTj6vISfQNJB7BRNQ37QBa1pNO/4k90du/2S+hidTQXtDk5+aK4fPOaKhyyrFfr7mTKVgeMO4FGP
HaZPW0UKERLh/lonEtTS3EHQBNDHB6X9xYbf2ymmT0e4gWCYbeiK8aRK19q+qHwJuXu953BJeyzc
OqQVznBg6per9wUXgWPDyMTkJinEaA2R9gS218T0GJmugTrOF9nyBSaBsATmd/BUh3VqWQ69d5BX
h7c9Sirm1nry1FvLszcZqo8l5Hfac2aBgj4XWojGO3j+wvO/5sOhsIBKWe5CvRGQ/4q09E/Fa82f
sEbN8jDuvDM/ThlWkdJQM5O6uoPKlB/cWZPq5OMPWlhwBlYXubGxOotl+zsm8x+X6ljmGJvTEZMR
uj6MkpupA2fEbZnF411GnqP8LON1V190UAZshmIQWADONQsOcSGC1bA0ePdUXBgDIQWH1VOZt8QV
+V8yjHMfgFEJ4CkRcdXE16e7+0ex+39UvjkdUbzdyqGw+XeuhVHi7puS+lJ1/lDhh36KUfKOn0OC
rilTSjwH4QBZq+GbuZjrk/xaNVzle/0nqiCo1gjlp04vYP+RPxNJOXj1HaDU7JOGISZi9MPnW5zr
Vk78qdHGIINyNOpDz1dTcI0OWU7rD1KCMwmeC1XUD4WlskpHHRsghYgZdEkKYoBab7HOwY59qH7S
fvQ6N2aWdb94xYs7uTbiq3g3mXGdHKvpYcXv66O3N4oezB7nE5XLxkg9ArdE9kArWdLmeXkic91x
M0aPrmbHkaxgtclw8hgUp+o6ut53r84BHwFank7CfM7D+sVVK+Cde6J4PE8YQWZuLJZPT+7wG+EJ
gSL1jLgm8wXE80wt383a7xM8720PcNAlmKWarkj/7VhzPHNOs0fHgOulLTYWGyEHtK80tZ2rS6Ll
X+H+eHZAD7fJEa/V3QwWrksDtyxQJNbrQOdp6qRylSJ0jkRvhlUphbWItNaX2pdHfY+ad7niY5Kt
F28BI5b2oDGFDJv8aFDmrKW12/Fyr3Ghp+Cb0NQ+dniXqMn2dfUlEq/r++WfBuOZSx1VRen4m8+w
RWdQT2HAUJFPFTN6RcPuuN8GDOglgnfUbv5qlMZH+7RfyYOW5JVsCkngJmHDtWzyTOcm+ijljwsu
8lN9YV94vfVA74QEzPBtTsldTXF+wXMjxQ7ZuB/hc0cHlwtRQieBjsKpYyf64t+Nf6HU7A81vt1H
ID3Fx2wkbB41QRNHTO7p5+jIwoL6wlpPeYJ4/CFc+AO78wCYR2lVyFaWZsEy28qaf/MMV4zbe8hv
ldCOzX1KZ7BsEylVDryFIaCEv/Wf0hOceshQGyHvQilIn4G8xxzXn39napSAmyz4RN8VSUksrTqe
SSfVV3jrvNVrCE0Ay23tvXRbTV751wfIQVZjVu42+f0hZTu5489VQhHNO2kzmT4I/5wQbalft1ev
nMHFFaNnL+K/ZyP6wK4N7hhlaWFYupz/dP9dnIP7Pd31UwGIrLwwbUZQj0Ql5k5aAIl3DarLDY/s
qTfBEHroN/Y7B17u3giOy/WzMgegx17gjWRNlXKoWxEmyFNDWA74H0QVdnWM0whYN5ZXMF5NG6PS
5RsU5qxq0MhmCzXnqR9AXm2DLeKWyBwGNETt7kGE5cBjpJwrOnAPycpVg0FmEbnJpWIZZ2Pz8zCk
OZ8wAI24mu+E9S21clQVTzjphFrrqEHpfjgGxg1lPFAcDBRx8vUNaw6o+REUMtkRpYXmv4kSgUvB
gUBoN+1EiEr8PIHX1mn5mqBAcPTueGszAxuEx94qeAG4FqFgEakwZbFCVBoWkADMjXZQoIXbCsyL
XWXDM+4q+lm6Ms6yEo2VQJ1+XkbpH5+F54Im63xqGjLkpA++DwU/m0f/4KDIY7pzLHGGoRnC10H/
hgQW/71NiDvS9Xa+OU+c9oY3d04yQ0+AuHgGRYta40QtrEJxsThz0hiCa5Y0MUAfy+CbjBbZafBQ
xsYwvif4dz2lIVJVpaOivRkoHtRGk4ko8AMy9czk3iX/wtlNJYkGL346xkHpIqdj2aB+WMp4Aymm
ResB7MikfHXn2QBiL6YMNL3HzzZkYigLP+87s6Mo7Xbo0aR3f31d1bJlY2HD4NfNF86dXgUS5nfl
j9yzJkKWobg0EG1lVrnj9xzm/5Ro9Hu3c9OTPBBv5Ulc/umJUHmUKgRwKi1y131ZJ5zH4OdjzFvm
JpmiTNogTgriMZa4FhHQn37ima5qRpNkMjAm3FVvkv8zHC1U0kIvVZ6+V2CVq+tWmTZqetVUuz9+
o3rrOPhkjKztXszLRXhR/B3x3/GhiQQdaCa9WHu5vzhm3JYcck4vtOAWxu0gWor4S1HwsIN7L/zX
dJvS6U18DoPkbT6DeHGZgcX8hoZyit29MktoS4lmV9Vm3qGctTY5eK7YhMBQnvEwnA9UbgFLd3jb
AgxyF8kSqOKSNnznF6nHgsGNtwSl5CP/mq5vQMzXx938JGx4nvNpY7LPSbmXxXk2fvJg4AIQQKG+
JVsyu6gpfe0k6OYOzZUqdiRUitvnjMu3sb2DHtGjYvXQhBhIoXcqXjJBo/4P7Yr7Cu1/vtkRIb+F
vqnQFc9Kmc627ElSUxb2sZiC8AMbm4QYUXa2+lCmOAZlKlAdtwKgpcT9OOZrgvCM/0MvUk4EKpnh
YrFkPjP+PbDZAq79kt5asikeFCylwxklsX0hEyp2gG1IP1WcHeWnziJtVfv73qYDI5uwZO8z0zgZ
r/8sLKDbB32hYYgCBqCV9Z77DCMWyXKvujS3cZteiSSLTlCOkc32DaPO5UIhGZOW62aSnjvc93eD
6ssPaOIBvFeE+TQQ/orRaZkCsjcwkUQrzWSCaSB/NOzlJAwEPfJrlIPYSAqn2zTQ3YN92wJ+Lg1Z
HNYJcXcoMDQeViysBrF1N1u9KOG5Ex9Lt3dOTXmFmFbIgGjuKMtDfFzUjtjJJP68wCGs/45Lbzgl
xP+/QNSI/X3+36S+Cx19nhZHFAvh5pgwr55oAaGz3WPcOLlEuzj4eK6N+cw1O7VOn4U2XnvmcJHT
EUSJnZqGekj+MziU/grG0/767/E/simJmjcGRJY2tfYhC1R53puRxtRW6oBGFPlZBZV/vBRPP2EL
da1H3SqRnhlSyhIV3Q/Mgd9rqTllropc40S8ztvK0kjaaRCdqjQrzZwnvLfFH7xIGHfdVqEiHA1G
b+Sb1qJiwta2hKhIG2k1GyjRE9p3IjFMsn0L38whaq9MGcbHDAxvnZyqfMDtHKte8UUO0tra00ON
mWS7kwT2j4L5+Ivv9G8KiYjJsHtOhevegcw4+dNBhb6yCmUQrzUne1x4ibHukloHoFYU98zsw11i
CWuT8vsunT25t9deJ9Nid0uTsoZQ1gTfyBaETzUujIbAkVtFGzkN/hty0JHwIi97g/SfKx1uXTIa
LLj/TNQwspLdoNJgUKLWULw5Oqgik0RuLm5lKP20h/Q3TvL8TCr54otu2nQTgbalntGG3sc9BdGI
HrmGs9bJk0yKfiWlwqZXBdxFe4jemf8hSytgaaHfE0rC9yxiYmJkXP2lUHPxQl0Zyd7j86VlewLu
RL+UrNbjYD030Dy8x9fKT7ePxUBeriFr4f/IruectuDqg5kVPTvE4rjecVjzheRo4T85XvreNGNS
PKiKqyq7DAxORniP9P93egrd5wXELiXUNqIIBDYt+SpSNkR3boZea8plyAzKs6QW2ugeMv8h+xhm
B4v8b+lRjQGd78zuPqe9WtkkqUJx9BV+sQbYl+0GyhnxyHj8CItkFw6BjwggQ+xXvQvkgDvbw64b
kkwG3E60E42lY+SZIUvkgHrEGDL2FXMTdexfZTM9nQYZNFlk/XNHCmpaI5U9J6hJebLD+kxUzE9d
HS7JlhUXOzcUI2x+Xh2m9H+uH2oxUIdfsgHF8Mc+YS8PnjBCrT2MwsLGG0PfrVlRRW0agxY+JOHU
N4s3w6OryuvAx/DSzVrKvzJztFQ2xTewKJ+vh+u47h7fMaHJ1uR7Sv/Qmo86XMMqM7hjke8Dcs8o
tKWmArxs62NxtP6GOoMrUwDZ8fHrg+1e+9sWPhU0jQ7MrVnHmcWJxVNLG7ddvPoVJcddFQwXOuSy
ab8lRpxurK0Bo8qw30MmjXEXF2QGF291tvAAm+ObIFMmNDUmrsaxT2cNn6BjGS6V7p+CfHpCRW+Z
fkaUhAugUSE7l7y87Uax0kNIV5bJEoi/t/uBma8MMhkrEAQMhnZHY5Oy96fvGVe/5O85eMrH7Rnv
CftRy/p0PXJ8pQz5n5Ul7T8Kir1s11nBTCFkNrDC/PXUrbidCHZT/O0RQRUWHfl5ZYinUQAJtr4l
4HPA6jwndNmZf7p+Ry2ZSFAJAUa6+hRYkvvIIUg4liKtp2GZCrgWMs1GzQUCdS/gVpSNiR98wSMD
NerpccK5Rr/RQPXjw/9tzXKXQWBpEAyG0qST3i1TCJI6OPCgvrZAqIYf3ny9vqDDBfb5cNxQx2DA
4qrCEsvRkS/8xE/vswfwWUmpPZfm7/IwQ6WH4zkbEjJHbsLPS+YaFRSsRRb7D+dj97nfUyFlHoqm
x3vy8aKAm7Acq6jnSxwvRlmQp4GGkYew346mLD7k8fKKWB8r86+Rj0CFsz/GN0mU+zUbuT4ZnE2w
akkvsVYC02HZAChS9MO+/taDuapEQdkMzLzEC5OVum+JMBbm8EBgfcnIx4iGneUBCrM7958bnBC1
8+DcDS220dPMjx3EzWqUPfx9BoMc9MobR7DfSInAELs5tv5EQG6h+n3nwpO0RhyOMKSctOSuG3ky
/eWdmgdDtOcXaiQUt9j/F21W07WZD+hXowovip044yc59hCSDDluJJF9+a9vjVVcaxKrzwKhCSPo
nkTAHxN3jgdvtqvj9cvLfEVGUBrO5IwMB/MXq00C7cl5eiAsC7PgBslpmyO9E9DlodhQfZ2s1JNy
ud8QMXm4GQ20PMS9vgbkAvqdODT1SMDhenoZVjbLxzwOE7xG9yaG2pfXmO6LL92WkB1a7h90hxUt
MsLahJJNB4vsqV41exhH9a7OeY5C6N7wikHDAnh1rELmga4xvosFWUoBrYUqUmHy3+WisrOYl54W
Wf54BEGITigdlY7BE5eOM5zM/wvih6OmbuuVwvJOcL49E/ZqBwXlUKcWXAC6zPKiaouU915BvotX
wBh4qxnpbksE36RLd5D11FDQ2QZGYth1sDZETcFyGD7tHi9IBVSHMmHOBQoVd8TvlZIUvwHgVpZk
exsk/R4cITfSyITN2W67LrmbVSWCO6rWOst+bklUbWwq2jrxvRNSJAQ0bn5h6f5quFJY8bsFIUeY
xctl8ZeZinBp+lY3adCGSTiMObBNQ1WtmG+fGUkts5A4UOELoj/vsg/lCseHtkM8R/YgfFHe+hJJ
Sjn6F9CQdC70iczSGOTH4+RfqSJFXMcNee+tJ68HwxKMD94Cg5XlmZJoBj58nrTOCMswIjK2Js3w
5GhwKyeIzEf6i6J+iqbWBqb0yu7I/YIK+XeyErA2zFCzf1sRZJf2eP8da/KjSPmUebTghZ+ZcJG4
Cgy/CXKFVeRM1BRBhXBDLK5fej6TjfoqrNBsxi2B5gGFt2AL5wRmjqGdbyvBt7g4PHthieJLKyji
po+fLJK3uYH30PiqvlLp48UzudmAXrrF1jvED5uMy3UQAHK4qGUVKPNTguGtI4b4sqCKcYfBS/hw
IvroCAziJBVpbCdOXf21Z0+96j3lY+PgH3NXSFkUeC3l6BqtJmv2TsB5mVbhzagzZlN/449E5txl
sLov3A36zYbaZwGRS/to+LHJ8aXgxZOVydp2ZV+hPuEm1KkcEzu9J4Nxg2qQsOtVlOf54e6Uq1eX
rtwaGMgeG+JnnrBbAWEKtM8C2CB2FQKzxYu82kFJqfSkNjjMXt+bn1TQfQ26S1q6dupWcKCSHenb
LVJHKBmB9uIds9J8KtkC61Guu0WvlMHcB3DRHjyiJgwW2hSX0+ZJKq7eQ5yRwnP3lwZlJ9NH2Isf
ZD4NFdA6KRinLIdnZL8gwvFo5ckgXsoajbjBuE2im+zSe8SNhh3GOtdnUjMCSkQwbbbykykqIOQ7
RhFf/D7MlyzVnIy6PZy9hCf0Ze2ZMIh4T6fkxH6zEPV/5qXfSQnumOZIpgZt2wIDVWnASPl4Pmu7
huYzOjvW44TxWiysxu51n73M8DvnB5DCUbjy8vWUwg7K1fcmtylNxrMYpKG185XpBXhA9ZX2QgFm
7TgJio/YfAvD+D9klwfkdtw1HWFZJvsE0qYBK/X5FFeanzypTXXGgjyb2+NvtRu0G9cCS1rbtu9P
fZiYVtRPYGQPVdhnH8/Y30T37kFXtJIrhmxxu6HYgrtRrNSQ1KkR6WeuzzmwtbXLIqpIv4sBf7qO
EpaXV9rgZBGyubZ/ccqQpTVIOvK6b6pWDus7XhUMKMHP6Y1lndvbUIrPUx8OawHSQjJymoxHriCk
Kxu+dt3NsHvVdtbadO8Hz6M5+JU5ht9w8QbmcRVrxSQXqHvlsxxWGc2Y5q+bmqJ9lLYCTRIJ9XjH
SNao4RmkG/oqfnxbQoVkZDXwTnCTIvcx8eUFQ0aRgCQ+mbL9Yi6L3etkneH1OaEGndZRtRVvp4Ae
ujVW7LNuDTOSKPdsEN08sy3W1HX5ZdzoUwZWiPdbc+EQgiAZ/ukx7WSw04ao0ZDhShRQkAkjDFsH
bUhIos5o5621Xr5NhMQm5WwsaYcesSM7HaR5dBFzcYANKl1d09QeURj4Jsv0Jdp+mM6NpJrODqBd
jNs4z0NnQgVxzQVf4Ks9xXJ7f8NS55g3uGe4tlOYGD1FfFL+UEnMsluFovGIQY8UDtYFpcgPLXQi
h0ONSII54qObXHCAB5vXp5dsOyRmcYe4sCZyzkQxM8XZKkLwa3YqGjRhxcgozuasP2uqQp4my0J4
5yAiJpZYCzYaOXcyYdWsxD4a0JdC/jIpUCqn4+r+VB0BVUirwozu/9Xl7WFwoQbiN9FiH5aauW2l
E0AwsHzYSDtcDOdML5mUNKkcH8YqOu91OrVpNpOiEr2aTp68GOlFKQ0si/dWfwvvsmQxf/qcbgQ0
ftx3+0O/nIGeLESzC9KhihuNL5pUGWMLwr89IvQo6zbE30sGYgzDfbpZ+xe1wF1RpQU1FlVfzqq+
ctXSIiCpRMF2fwtA1zCxbPXDjTewTPVFbf3Acg1YArVfHFrV0QEG5WUQhWTsvhffO5St2ST83Zm1
uLahsdfE8ejMvd+/3ycU7D4YgKOUDTryXQX+xAPtlp2HKnUAPw7evIwYI9uf3bjyl7+x5vNqNU6j
sVm9ImJYeA08TadBKILLm2tq8RDqjEKa2ZlDlt6X4neCCuepetRkIAQ1jcCxY/zhl4JZH2HGSrtW
reeRh64Zg7uA5yUm8eeDAil8PCCCigP8WwakMSB9MS6krtQSA5UPf6gpwiEKh/TOwfYzd2+QoS1g
Gntw7XTCLgkYi/D/oKh4pc+MOpz6E7moFQk6QGBl2K8um14fRTkWGX+1bM3jceQ1YsgpIfxfoMTZ
z/quiSnkdELKxYVP1cLXqgd/Xfis8b8ZHgr3aGeycvYvWkrFtas9eu2hRanpIwJnWTxpRi+pSwLw
FeL2xjt3cXJApS/DYYv9mTaJK1r0nVX+f26+cGGXPXuWfrYDvu1/G3xyWQi2oxZ3vmq2RWb2+Ljs
Sh6JqHxJ4gPPRsdYJ/tqUsGmI+ficpazm3aa5/XGItUr6m9O3NozaTUs6YCW80GWOIjG69mWyo0a
0v57udYtHEeoiDdx7iKPr3JQEPKdmkXw4InTiIFeecRcH12tJRnYdL5CtNYkfbnP2acC4LYNqk6m
9JF6R5XVo/Vut/eDMHjwntMx3Gh5tlEMsBjsipUTo6kdaIWCQd1frWktHa1351gWyfFIsIeBmidN
bsWFSYIFpRV3OrQkzagxl3/Yf4duqbSS6oHGO8xwJqcNgZd9C/wuapJt+7Njk6ZvnPTO8LY1Jutw
N852De0wLiUuezSMfIpMfB2Ma9kovjMuxRcO+eJfIaoT9QjC0ylnOmI4l29tysAsnOW3EeSa7nhU
5fAf4yenM3t0V/T7Xy/+sxnDxYn9c1FiKgzHMwuTpTtryvYwFhMBcmhLBwi91oeSmpWZE3mwnSwR
VcXpidGGr0D45DwpeteNnkD4DCoPQ01l3KTA9F1wvUlGz3bcDguC4MRTfJQyN+jLjn9i6TivEd6/
kmKTK3aLw0bdzLwYc2BMHalgGNeFG+6o3QbIq9HsELnaSKjSw4XS2CUr7YEWNbyrN8Oiu3A51I1K
NRdmuirmKRs9GyScSIE8+IcqwNzuTASYFcqPiumLbl/a6xfXhreNE/0MBGO1cBqZMNu4OyUI3lYj
HTJ9IAccqyn2CwxdIw3cqNnwQlaDq7qWcipQ1tO/2jgmaREj3UXLCttb5kbXiPCm19oUYcaNOaUW
3zfUs/SfI9qvV9GX+37L/0DaGP5liZxDKtxnX9J1P+gZbt4E/dC/2FcAvSawgRtVckYPChA++TQi
FGv2FhiPnRy/6SPdv5o1XvBp9DdfXAmnkYhv1weUIptAr/6yu+IXBC7OohoiJYmpPLTIF/YBUSLE
07Ueayh7gkc41VqL/zM2kIvpjYPsy6kWW91OQWgBE4oS2Q8w5kbg0gidf6rIpGs0hXLVhU63HXs3
KTAJQLgjYkZiHx+M8f2iE6r5k3FCtCue82R8vBy44pvZ1wOdGg/R5ebN6we6+o9DIwdeI3/DfId6
0BGjIIPnQltZwg95c74pRUXhSv0yf0EP7zWdz5Ipwl0xzqv4ghA9vnPPUAJ4gsHFT52ggnw6pglo
faf56T3ZwXTaXOqlxD1ZSYmVLgr+E1p7CwJn48S43Es88XF67whTQZPJlDi9v8GEx0uc65u8uffK
PiQUshYC/65OPer3Uh2vZJ0Vwc0ZpgZ6dlJtrNkcIJFXORFN9cKpZ2dWfFXdeTc4UC6Zqk60iw0D
COQB1ED80aE+iGuQ5xIzsdxVfSVTa12duvJBheLv06A0Mwg5zOYd11hksgow6iQ/vl/dEyPCGpYw
khVhHyxDvG6Du5svKvVvurfRQFtIMFCSQuErYoLtVTF4wA2ONQXgWLOq9wG2eagicY5JDqPFB9jl
U9xqcOXabvsG2ap0h+37coPCiBAke8WkBf5cEoi8rYXWTmIewRr9UI+pR2+S1/rm/LVin8G8ESKi
PXkduvm88OsGgmYNGMpdinpZab/OS0ZTGMAUhY3TUknTjvXR+YQ4u6Q6C7Q5OAKR1BkJhaik0oru
UWZw9uDnNJ91rrgJUaDnmR+yyWRJ0xDIsHovKRp41wEAHeowzkaqjrpIn9W79D5y1UgiDWSKzIUl
soQHp1lEH2EHlVgqgER5B5sn8LZAPreeoACCQKxe5N0aNV/uROkyevxe21Koa4A6IpZBcit2L4KM
u3TUsfpRaTcDaoxjoBcKAtT86bshtU3S5K4SzpJx2zH3MS4dqPaMpGbJK3ivrySdNAU3xxS7QoEg
CLbSy5enuJpWlwb08E5GzrTj8jqr3FX/++GGL8Vn81bI/J433jFS60bDaMhpmAyxJu6JXNFXb9Na
8DkH2EevA16JAKnUy6+lQqiD+ofb8PxI09JQlmyh9dX1Af3Fe/YbjpUc+DDqsv5mP2WoF5g8X7SK
if7oK2F2jcDZgpxp3oeJrBKRhFT/7q6oPKNjTTJOsIyhBPVslQyZ9+HgLLXEawlHt0rBUCB8mSgP
IJg6aO4n5+8V/yV1/MwzeCeEW+rLUM2mZ48xmIGGUF0l1/V9vxTFbnOSnIAEH4hkkra09X7a5IOM
dzPYd149zc5/IOJrynFgz39urTtrFRz/HU/TCWev+GaZCereJwlITrZyK3Rkr0K4oABC+YZkdwI8
KHfk5y3a5ZoYr7sk8Kqw5ucNf3L1KcfPMF/laE9dvcq1mhgo4Q1lroBFwJac7/q5FVP6AMU0vFX/
NP//7biwWAxlhw6tDuhREShP0H1jXvb285/Ze6+fqNM6tS7+kvnBpbUX2pU5yfBGKGjx2mvj4n23
GRHros6aKmxJ9TqyQTi7l4h92iPHFrcW0+hyw3Wi6pg8mhyXydnkG3qVAQVbARLraAE3Y4c01wbR
oGwLv1JmSGTXOwuuYH3I4Zc0w5RpTlFpctL8yqnnETz7ut6V9PI0TDf7fXSue+70c9Rs0TflhG9L
l7vTSOmKszSQQel7Cl87QCI6JH6bWFVgHuJYfx8vzs2JnrNgxWTsulW2WP+sR0gfAxdfsmsbVAER
9+QYtdhRcyPuHr4h0M9Eq/upiBnfuE6WOM/vkaxITdV91KU8gPFQVHuk/RL4HCXeZ8gw5il117Yx
fDhdyCYccvB5yHpOaVarPiVcx5qaZe7nwul9Em7WmPOa+yBF5aJxJruDCcZx51Bv5AtkbvAFHChH
rwO/1XXIK0tsJxe8Jx1uJFf1xNcFWNSmo3Nk4MaVdkLfu1jfrvuhIBHp0SWUvka4o2dvz+Cfac0/
ttNyc6A1IdezkGRO3/3/YrRe5e+1xc54fvSznOAVqD/DjwP5xGH9LvFcGqgh73xegLySbaXw2WJD
aYB/25z/r1YBvHVrUPgSO5ty4Pf31PWuDxiVplK6IMik1FE1k2U84JBjxa8FrFWn1Z4x7W8955Bl
FQmo8oN8sQos+PslKTi9gHLiDVLshpJ6H5NvRHbHTFgI2dUp+CvTUTFRL6YcR5gob9KvJ4F1dtrx
nKk7r5Lr2RUHqVe47c73kJx4HbUHVBnNDyD0KH1043LKuGxux3KNaVWl8CIbfkejjZu3rqNUUFON
CUE05JsrwIwURQFefJkhNhg3xxNJ8q7eXVeb55TorEMz0qfmuAf+8Ns380rsGYvTrY6EeYukjBaf
96TVPlxsyEOxuXvi/3YJwoc2/+2ztReygdVj46QNKgUNOT27DCc1TUUTXtN1ZtCq41VzUDXeX7yq
+Snpwttwuw8/r9vGrnVCSASQsUQOZEJIjQLSJY0u7blDT3Q1EkS43dO2CmcsLbj14TEKs1ZhN7qq
moDiLomUqnLApdKHMnDPjQdUWDxxsMmiceSeMuO48AxTF42TJKGu1QCnxpSpG0XZlLoL1Cl8vfUx
uTH6oSSlXP3CyHXazFgqNacByycbkSk94XZfolTQV0DyHjaVacQ5hq40L2gYaEjAex+aK/Gxo9n9
LJFvBtVbioTFwpp65UPBnP+a20XkBFqOEDMKRGhlKRwuvz3/XQuX97muz7ZObPggQ0t69vqE6AeM
Oc4DNA9IHIY56nmdI0Hlisp8nyITWUPp73hKiKUTKQes4IammxYPpEtcwl4ldG4yUB0uxL3hlGZv
s6XQYXs1HbFfTK8YLW3+oyBEZJt09r72bQ5xvwME4ig1TAURdXf8A4zTlpRf3RWrgNRljM57e2UD
PHTk5wE4aWSdOcW0Acvka3SQ4rUAFl/9WQovY9ItFxUiWnUNjqwvjJ3WnKlbAB8wXGO2N2UAiKtz
zZHRhEgN7X/6JBKtHaR4msw/D77tYDc9NZhD7ZGBZX0W1NhwbjVj+ZGCnIXdi7VgxadCQv71BxU8
YTRNSuYLZ72BsTaYKgOxKh+cXA6W8gzkUiW7DEvudZip8WsAPDTw/ZBWo1r+2fuhyvBxhYDX0zsY
KiUi/JOgm8UyixlgpJS+E7NiPGZunT5JaJzka8+W+MNXdgn6JQTHq0duIgA5FUmfYFvcSh5yLtci
urRUrlDXttKaRz0hR880iczd24s5yrgz+Ckpo1vD9NLgs9ip/bdgjVMNsBRYdqj0QxdU8pz5qoTX
fKdysOETnOK0GTUGj969p+ZNacHSbL3yMfz3g62fmYJh9onio5Y+Cb9/ISdDazEbzawrF4Q9rV55
USwSvtuRuxWR5IfjrX/WK2+8Hk1WaejZloRW+srFh7Njl5inGK6Tq/c2qPpjvcCIziE365K5ja6t
9FuT7mL44jwAnRmqjda8pbqbhosd70uoI78nbkifwECv8Jv4QGUBeauzGPsgOszPRa5yZcA3xSA9
Dn7SaxFjk3P2lDAOr3/R+9ZBHbOrFPTbvtMiWgWy/JMl9AYZ+sAPa9kptq7CR1kRobjGp4Yr8qYy
5zqczCkrVh8zPWiPhpB6cMyTrUo1mdXci3cwhBL/sYiVsHprPdSMQJJwVb0VsAsgT3/CCuOUyNcJ
YTOBe4ui3WA2xNQf9Rpqo3v5UrEIW+NJDdU+JpHNae3IJWRj6G5Kh5SLkgtn7WVUEc6aRePOVcnU
YAtJ93NXWzIQepAhmfByzytz554cXAunedz2IKlc60LTIkyhUuBGWXVfBVSEzD6I2mwvpcKoI4vC
yiw8ZKzOOhLBPhZXAXvQ5Rs7DxfY2LQpaLQCcf5LFf6yEHVAXAJcfE9MtWWSqV+f9jH/rbuzHH8R
/39R4Ggco+4ErYzhqokRoz0=
`protect end_protected
