--------------------------------------------------------------------------------
-- Copyright (c) 2023 Arista Networks, Inc. All rights reserved.
--------------------------------------------------------------------------------
-- Author:
--   fdk-support@arista.com
--
-- Description:
--   Encrypted file.
--
-- Tags:
--   license-arista-fdk-agreement
--   license-bsd-3-clause
--
--------------------------------------------------------------------------------
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
cDYKsWz72KPaEITecTsL/72H4qNUP/2hl5fQqphvlqncmh7KaaqN8lDcv3CuqVNXKF1+VAYcB0Ft
uJRAPZ4w3Kf39Eomv4RKBDZM1Bgi7naw228Hp52WLTJUQqctJsxIqOfs8xqsG8OU9EvegI3Q31Zs
T3+iAdDhs3aVzMMhv/gLqWX3ng+oxzvrRyc8Y8gBDnfIfo//N8N0sIKhAvFrwy7bJzdnjO1t0K2V
7oCirL2llaoQ/gBsjLiUeJf4Kf4IAGf9G4B67miA+ttalSBhG4GTJQ6cSQadxt6xdMyNpe3gMeaU
SleGFj15xyjMCEUv0665/IHuC8WCGDdJTSRKZw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="8B92CVDmQlpBSltVNYMzHAGD7jghyd78kF5zqZrLAtY="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method="rsa", key_block
bqm29kRbnaLPKQT+1f3p0RPFibOOP1FYOgWFFe5HTf0LGipz/1aU31+50ZOoBNLDwISTU/W6FFD1
wZVAgUiwpnY3AphxSgyJwINrS9YV/JtS9f4/7xezYxmQvhN4i0N3rFbt3S2X3RadDGUqh80jKEWF
YpjxWmz6UHEeQqMXhsoAb5lmCQic0VkqmZY0q/vkVFq6/jbjgVzrM3XO++89v9/kGel3N2YJB1tG
wU6nlRNMs2UXOrSGdxRuO8IRQ9PYv4hsmlaOTDcvLwvnw9D+ZyhLKw7c/woaeMHSjTOUhmSbjfgJ
4JbHlVLGmT6LsUSvzg5DnBvvl9Mv5+1zT0a22g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="sTVXfAq7d3dA1/GHphpmd13Kc6n2151PtHFiaaDlxSI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3888)
`protect data_block
P7q9XXOLxn/ry5BCV7R/ghak0N1qjj0F3PgWluFszz4qzZfp2AJhEH8IQ7lXEnl6jqVNFDlns8h+
TVtfQosE/iQ+0+BnZjVDhSPtVF5czJO6rqL7JidQfPC5eaLQv0fR4bQnM2rEv+3rSQi69Y4r26vt
+k8I0pAfD20nCgyuSDUhyvxEvt0HbI2VvdoM2luEUXjHf/kz1JVURy5ULZ6cKRIo8+8XoC0f9zMY
Ui/3l0VEYEbLlpH3W4wXYbcANvdhskICFIKtfZYCJDaMo2sLtsWflze9kumvjLv1d6jIeyJeZZPQ
LN04ri65UNvFjYiajq8oo0pu44Vfz7UAzRjdsVkVB2bQZmHLIDgxQJLI2FzoggDyLGsx7sLqfbx0
GzZoQzXkVO0Q2UakiyZdWmAwhrmTTm/UbnXL4nLMPF0gomVmBQoxPilLnLBZ2hx5lPC/AJeKqWg/
tRcKigcWFZX69Lxle16O2I4EBYjYT/X5Ip1t9iU2Mbqdr98L2yhsC/eVpF3jOrQWpK65nysPx5q0
KG7SqfwiPcxIwtjQgWroPoQ3tPdqgEjHqEn8b681T8Ov8i8z52lERkzHftvGeiKKmRHrAYRAfa0G
SRAtGT6EtOwn50dbJublkYmFls0x2a5Sf9C0zTS6cuKOG2Cura03+SSDv5OwJ1SKc2w6GxMrtdId
pT+6K7FkmylvV06cDE6tsR9dnbDlL+pTs9aKAxIUeOFcZiG8vSJgDjBpl8FuTfHYIXvpwKBBW7aI
QgwWPo3pvMDAwCTn5cUpM1FYRoNZnOODEn/IYCIf8x7zr632LE7THankDDdvxNEQbsLmvRYWc6t9
y3a+AIxyKQIPxhPUN99vbvyRGtCneo/fEBWFKEA+gl4spwWRaUvwU7+i5n48P5aVZUF873Bf1f9R
YcHzQvK9YbbtN8vKR/6Lypa4gFyHlB9w++PrUD1p1hFzGjeaYQ7CR87+HiP+tQQr1ybzVj8HFLF7
57IjAoyT17T4Ig6UgZHMfEQ5GZ3mv27SXiEEo6hOhQ2m8BveptixViVxCjYNu1543nYJdUHtlFUV
c+VlNO0l3c1u+0xIAR2fcde4Zp9gjgZGOx0M1a8QL9kisSTZIFAMSEgoJ8LQ2Ld4wo3qMrF0BeKa
DaDY9iGAvlZ18nB3qiopElsg8vDdAsbvg/nd3gkZMGdwRxCKNLy4Nv0TKVwKfFZ6san8qP0VsPrL
4gglFRdRrLfEWT7ZNl7OJRdLE0OqDWtcMEDz555Gs/hOtU9Y/3s0qPRIvLH7dN6IjsYf6BIqwWpV
Web/mU+xgRex7qNGlphwZscdzALuptSBYtJuLndevkD4uqQWZVAAu/WV2/NuJ3fyURc8DXd4WX+s
0vU4jNK2BYuZ5w9nhZZQSwb5AE+XdQh8HBpoDEiT7zO5mp+niIoaodZXeosTmIUDJ87ai5gaNCbU
OrXzXspctQYtQfOjqdbPa1YEYXK2IsGAsFUBT2ZTXWCQzuS6Z3LHMpqei/iGgyqERjPfNPhmlAkA
dLzDQHCWSbu2EwIaajmhSgK6unpQzh6XUuN03IeNElAQysQixnKghe2h+D0ZIA6lIL4md1udh4+3
2G48rua4k+fUrurKLFe4X0tDOyFGNbiy0i8U6ce/6bRwWKssFA6gZhWFAabyfcD2JKLZlvHsDGfB
eOXuI/xQ1rHmnbEVSQf24IPteXnaTJU+PMbDk5SqrHLLYuqKlKAlPT69t0F99ZhybpJUeqIFfOpI
GP7Rp+53dpMx5xOEY+cfUHYSMPjedIqCx8wOc20etBglkdhqA9RQArezerMgP6jbPdjaEMAqlDGY
NJbx6tfoMAiO+dphKfQk7431Pl2i9f2M8ZOIreNa4GkFjzfThai9esPi6x0lx4hvVTvlgKba+gGh
O9yA0fOunVKQ22Jf9hkoHp8zMKQQIZbhl/VP5ZoCo/bx78pL+C019Y+SR6PhuyHVYqZLiFZRvQ6r
XBJEPPMQCBSpS8/afhjhHR7/v/kbG/i2JeqFdYqT6LCx83m4ZYGS6f1rkuVudNzP1mBpb73V5MC7
3KSDGIsjXBBwmrdqYjAy/M+CDqc5RBxRJd7TYEmz+eTp68iOu/1GvihJsjA8YV+w6No3VIkQM6il
/4B/2bUaV0D4u9mum0OY94BOlogumP88IvobeBwBh0G0BCZpML88yqmkTUPs0aqczHFcpk1moosG
2ejBMxdDNT99tRSqPAADgSCCxSoYRHFXeeG1TdW2bUF2UucF75gNzDPKJmpkz/iM4h6yTX9aEazd
Xf7I1aIiZuY6qw0ad99cjG2/wZ927NfbBmbAasa9ZLa96GFwY6XlO+GQbZtz+nod/Imk8cPZm9QX
blubErQynjY9rHns78yoyoUk/1CHBFlG5mIVSVSmVTlQaB+PQyMrz06rRFoiRIQtYBg53ceoQKt8
SE7oHtHyAX/rd076FuGcB69FRnzHF0A6EH0+dHrsJKbA+2ka0KBL/Zva6SqlmUOH+QQamR9BU12k
1WlCeTE5F83shHsk+M4vCVuisQXQLC8MRIUi7AqUVkDQEXD8wwQ96XJX/k5iGzCr1Dq0om/W++4H
SyeP2zl3Rtp6g60fcem/eRX/nGb6/QKFfY0+XM5GLMdBh3f17Chx+crYm4DhON33dQ1/Evo7uP9W
N4kXkqoKFngFOrBC+STpvkHFBfpiS2WDTYbFQ682bn7kFpbVh2RYCSlyNr7kqvKteRftsAgVmW9w
tCmt0OE+1qMeJgiJleLh0nli8swRRVLFFlMaQKYCn/Fg65iU4vQqFeWwd7Ft3eChxC6D4UKOMpL8
Mq47Q5oVAB9p9UFvMCOz9wVab5oEKu45ei9eipEzFRM4rTXO/vdr9rzlE1cfh95MxiLUc0fBTNX0
u3etHXfkSCva/tPQfp4EZBEhXxmN5JIwOox+prIzGVY8xgrZ3PPFL+udcRzFPJsP9TBWdDR2pZWh
0kxtPcQDsTpWxigGdYypAH+SD4je5OBw2ZyHzHZ1dSj7+Q39VpFh/hjxRF3UAnJUGGZh9ZAOnlpg
PaofcrDO9pNVVvEr5abs9v4kkNX+gb+2pRKyV6IwZMZHrEj85G60w0mwWGETwZwlok3YMR4tN6VU
6lGQkbMs033VNO89ydP3QEKkJ1ugfd8FoTyWKY2i9x7f11WUT4hQ2LX16lfW5GYD9RWf2VsPRGIv
84xGp44jN+Bg/sm8OXPGu++3/+pH0McATYLO+fXbPI7BboMdes7C7Sy2I4xMgQsM4+wA5kOLYvOk
aJBmRY7EkfTM+N+KBNyUeQhk6kj/VleBtfzVo7z00IwNg/dOwkV2ggOT88YHA6NfYXi65+2sGyRW
5eKH6zsePjPehPVrexeAR8qwj1KgcYKbNN/4mNtnrj/SKjBYgby9XoddFQm54Gu3zZuic8eCwsXq
PJrPfwVtg0nGNf/ZDZzbQFK3M8KpTBZacqEM97fKaSAR/F9R/rFIzzU6m1TiiqVkFw5TljZ1BYNR
hZ7z64sp2ZEbFFjlRHi6kHvsmZeW8ORtA0RCFgjkVSQQQfaCVIikleesQSu62tfJEwp+xkNNLU5C
WaIjolSOpM6wUoK/9fYM3feOnsEa5Zmk4RSlzxRXyL9t6U5+clNbELwVMzLzcqlbuatI72k9jqMn
KwDGDuWxHd71lzU0CpmY7iSUnTVoCtYryTjbX6NvwJovDPMQHCRcJmYi6PMYi44XYRdwu1GMOgs9
aOM8S7EOJdfatFnKkkGRaqlv0mgj3j9cnIqK4gUmXzSM5v77MeL8mnz8I575pcYFHS3J68AbTH27
zuZ5Q8mjv84b3DOHoYn8aRWhKyWzss3f1JjrrWpCZDmmjsitWzoE6KObnySXi/A9Y5y/wn+8TdLW
6BlOT1lqMLbV8yKowRd/kWRLxeUJx6B6oap0iiRj6jC0sWEcOlIIqmXqPcjqlvdlWD/46rUsVwN/
tlpnTLHLwHVkRc/PYjs3nZ++vQXx8m0GnX+JlTI1GKHLxS/MDxhpcezfO0lhbw+DQs8rFDpW2qpa
8Pq7nBzIarf9eoDtWorSmfgNbjd2jg4nuNn1mi3tgxVvYjnRvPSnXhYuFArbBTpEuEzs0EPOUAed
hYWfoi8IprvHSmq1N6E5C2WZyFizJJeI3vTGMC84jk1Ox++e0JR7aphXoxDKWQ+eQ1FLEY3DXShF
FLY/8cQrGLYqlj3ZkDveClisdEnZGM+bNO2m7ZA97eVy2VKl0SrVrp7onVo8iz1UgJHPjnaax5u7
srqlChzB+/RH6l+zNQWBUigkbl753v9cc/qe89uFbCpD5vkd+egIzl9VgqagFhhAHGp+Boa65oNi
pGMC3gzfFQW/ph/Ybqm8IuVL8EGXo9A1VDtTsmmcgDvqHZGMjAPJy802GroD/baKU9K/GaG/RzE/
QO9wmSsStmAGqeyKgNB6j2VqxGflzrtrbvfteUr8zX7RkO527tH5dIDJQCJo6VCxPkexBQmq9FZx
xhhZmXPo9ZkcID8W9l7n1u2o6Ltif0Q6/YHck8ggQr3y0BWBhQ8uT0jbWM1JOvgWN5E0NSDcoPB7
lR/UrtKEDVkRTycQBUPNwOFG7fuInCaLyJF15lsriPvkbGWasmLMMdQFoP3aBAXVy3B5VLrwbDIw
a9szv12VGZ+pASYp9gmIncn+L+P6zdEIcVKw2MxRKM7+zQEVQL4wOkn2x11bCYSV1d6wSgHHGelK
QDia4cQLAPHDQcqUXgqJwQWX6vCY75zLYeLsnEynpbBZlDzAUJEU70yQFuX+J+Z1tlwADFIQrLqc
I+R1/72jMQYmKn1BN1Du1a4wfKOofMeBE32cU08Mig/V9fQozcyEwYBIOYP72Hk3HE69Y56XFDeE
14Fpnf1Fdf845OedVWqSKJjOelHYVGZ/7PkKTFXAczSZSyInrfWTqdddkY//JWRQ1TnET0uWrzeA
l3CUv6ugmBnnpkFsFh5QG0wKIcM+jl6SDTP8mqfJ9wrrKn0v8wZgdUnu8kYlpqrPBBzmYHqCIhF6
JcHU6pt3rHFx51iYQMOeDEbFKU2zWRdZYW7i48tss0AWqrZmrCReHhqwJ+XKIl0UliQU8lxpoZq7
Ymku9XyQ+dXUCiJ+mWxusR9GwPklpNqO3E3w02NQWendACOJvvq8awCCzykEvSFBQiKXnuV9lmfo
QA8ZYanwBWI40tyB
`protect end_protected
